module basic_1500_15000_2000_3_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10005,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10046,N_10047,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10127,N_10128,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10145,N_10147,N_10148,N_10150,N_10152,N_10153,N_10154,N_10156,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10171,N_10172,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10192,N_10193,N_10194,N_10195,N_10196,N_10198,N_10199,N_10200,N_10201,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10212,N_10213,N_10217,N_10219,N_10220,N_10222,N_10224,N_10226,N_10227,N_10229,N_10231,N_10232,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10257,N_10258,N_10259,N_10260,N_10261,N_10264,N_10265,N_10266,N_10267,N_10268,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10282,N_10283,N_10285,N_10286,N_10287,N_10290,N_10292,N_10293,N_10294,N_10295,N_10297,N_10298,N_10299,N_10302,N_10303,N_10305,N_10306,N_10307,N_10308,N_10309,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10319,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10340,N_10341,N_10342,N_10343,N_10344,N_10346,N_10347,N_10348,N_10351,N_10352,N_10353,N_10354,N_10356,N_10357,N_10358,N_10360,N_10361,N_10363,N_10364,N_10366,N_10367,N_10368,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10387,N_10389,N_10390,N_10391,N_10393,N_10394,N_10395,N_10397,N_10399,N_10400,N_10401,N_10405,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10420,N_10421,N_10422,N_10423,N_10425,N_10429,N_10431,N_10432,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10447,N_10448,N_10449,N_10450,N_10453,N_10455,N_10456,N_10459,N_10461,N_10462,N_10463,N_10464,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10481,N_10482,N_10483,N_10485,N_10486,N_10488,N_10489,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10501,N_10502,N_10503,N_10505,N_10506,N_10507,N_10508,N_10509,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10523,N_10526,N_10527,N_10528,N_10529,N_10532,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10547,N_10548,N_10549,N_10550,N_10552,N_10555,N_10557,N_10558,N_10559,N_10561,N_10562,N_10563,N_10564,N_10567,N_10570,N_10571,N_10572,N_10573,N_10575,N_10576,N_10577,N_10578,N_10579,N_10581,N_10583,N_10584,N_10585,N_10586,N_10587,N_10589,N_10590,N_10591,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10603,N_10604,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10634,N_10635,N_10636,N_10637,N_10639,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10681,N_10684,N_10686,N_10687,N_10689,N_10691,N_10693,N_10694,N_10695,N_10697,N_10699,N_10700,N_10701,N_10702,N_10703,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10721,N_10722,N_10723,N_10724,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10733,N_10734,N_10735,N_10737,N_10738,N_10739,N_10740,N_10741,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10783,N_10784,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10799,N_10801,N_10802,N_10804,N_10805,N_10806,N_10807,N_10808,N_10810,N_10811,N_10812,N_10813,N_10818,N_10820,N_10822,N_10823,N_10824,N_10827,N_10828,N_10829,N_10830,N_10832,N_10833,N_10834,N_10835,N_10837,N_10838,N_10839,N_10840,N_10841,N_10843,N_10844,N_10846,N_10847,N_10848,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10862,N_10863,N_10864,N_10866,N_10867,N_10868,N_10869,N_10870,N_10872,N_10873,N_10874,N_10875,N_10876,N_10878,N_10879,N_10880,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10903,N_10904,N_10905,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10917,N_10918,N_10919,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10930,N_10932,N_10933,N_10934,N_10935,N_10937,N_10938,N_10939,N_10942,N_10943,N_10946,N_10947,N_10949,N_10950,N_10951,N_10952,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10981,N_10982,N_10983,N_10984,N_10985,N_10987,N_10988,N_10989,N_10990,N_10991,N_10993,N_10994,N_10995,N_10997,N_10998,N_11000,N_11004,N_11005,N_11006,N_11007,N_11009,N_11011,N_11012,N_11014,N_11015,N_11016,N_11018,N_11019,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11030,N_11031,N_11032,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11043,N_11046,N_11047,N_11049,N_11050,N_11051,N_11052,N_11054,N_11055,N_11056,N_11057,N_11059,N_11060,N_11061,N_11062,N_11064,N_11068,N_11069,N_11070,N_11072,N_11073,N_11074,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11086,N_11088,N_11089,N_11090,N_11091,N_11093,N_11094,N_11095,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11128,N_11130,N_11131,N_11132,N_11134,N_11136,N_11137,N_11138,N_11141,N_11142,N_11143,N_11144,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11171,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11181,N_11182,N_11183,N_11184,N_11185,N_11187,N_11188,N_11189,N_11191,N_11192,N_11193,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11236,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11259,N_11261,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11279,N_11280,N_11282,N_11286,N_11287,N_11288,N_11291,N_11293,N_11294,N_11295,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11318,N_11320,N_11321,N_11322,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11335,N_11336,N_11337,N_11338,N_11339,N_11341,N_11342,N_11344,N_11346,N_11347,N_11348,N_11350,N_11351,N_11352,N_11354,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11365,N_11366,N_11368,N_11371,N_11372,N_11374,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11415,N_11416,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11443,N_11444,N_11445,N_11446,N_11447,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11472,N_11474,N_11475,N_11476,N_11478,N_11479,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11498,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11507,N_11509,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11526,N_11527,N_11528,N_11530,N_11534,N_11535,N_11538,N_11540,N_11541,N_11542,N_11543,N_11544,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11568,N_11569,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11588,N_11590,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11599,N_11601,N_11602,N_11604,N_11606,N_11607,N_11610,N_11611,N_11612,N_11613,N_11615,N_11616,N_11617,N_11618,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11628,N_11630,N_11631,N_11632,N_11633,N_11634,N_11636,N_11638,N_11639,N_11640,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11655,N_11656,N_11657,N_11658,N_11660,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11675,N_11676,N_11677,N_11679,N_11681,N_11682,N_11683,N_11685,N_11686,N_11688,N_11689,N_11690,N_11691,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11710,N_11712,N_11713,N_11714,N_11715,N_11716,N_11718,N_11719,N_11720,N_11722,N_11723,N_11725,N_11726,N_11728,N_11730,N_11731,N_11732,N_11733,N_11735,N_11737,N_11739,N_11740,N_11741,N_11742,N_11743,N_11745,N_11746,N_11748,N_11749,N_11750,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11769,N_11770,N_11771,N_11772,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11784,N_11785,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11803,N_11804,N_11805,N_11806,N_11807,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11827,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11840,N_11842,N_11843,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11884,N_11885,N_11886,N_11888,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11943,N_11944,N_11945,N_11946,N_11947,N_11950,N_11951,N_11952,N_11954,N_11956,N_11957,N_11958,N_11960,N_11961,N_11962,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11976,N_11977,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12045,N_12046,N_12048,N_12049,N_12053,N_12054,N_12055,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12065,N_12066,N_12067,N_12068,N_12070,N_12071,N_12073,N_12075,N_12076,N_12078,N_12080,N_12082,N_12083,N_12085,N_12087,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12096,N_12097,N_12098,N_12099,N_12101,N_12102,N_12103,N_12105,N_12107,N_12109,N_12110,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12119,N_12120,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12134,N_12135,N_12137,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12167,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12182,N_12185,N_12187,N_12189,N_12190,N_12191,N_12192,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12212,N_12214,N_12215,N_12217,N_12218,N_12220,N_12221,N_12224,N_12225,N_12227,N_12228,N_12229,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12258,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12274,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12323,N_12324,N_12325,N_12326,N_12327,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12341,N_12342,N_12343,N_12345,N_12347,N_12349,N_12350,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12432,N_12434,N_12435,N_12439,N_12440,N_12441,N_12442,N_12443,N_12445,N_12446,N_12447,N_12448,N_12450,N_12451,N_12452,N_12454,N_12455,N_12456,N_12458,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12469,N_12470,N_12471,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12494,N_12495,N_12496,N_12497,N_12500,N_12503,N_12504,N_12506,N_12507,N_12508,N_12509,N_12510,N_12513,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12527,N_12529,N_12531,N_12533,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12548,N_12549,N_12550,N_12551,N_12553,N_12554,N_12555,N_12556,N_12558,N_12559,N_12560,N_12561,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12580,N_12581,N_12582,N_12583,N_12584,N_12586,N_12588,N_12589,N_12590,N_12591,N_12592,N_12594,N_12595,N_12596,N_12598,N_12599,N_12600,N_12601,N_12602,N_12604,N_12610,N_12612,N_12613,N_12615,N_12617,N_12620,N_12622,N_12623,N_12624,N_12625,N_12627,N_12630,N_12631,N_12632,N_12633,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12647,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12667,N_12668,N_12669,N_12670,N_12672,N_12673,N_12674,N_12675,N_12676,N_12678,N_12679,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12691,N_12692,N_12694,N_12695,N_12696,N_12697,N_12698,N_12700,N_12701,N_12702,N_12704,N_12705,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12724,N_12725,N_12726,N_12728,N_12730,N_12731,N_12732,N_12734,N_12735,N_12736,N_12737,N_12739,N_12740,N_12741,N_12742,N_12745,N_12746,N_12749,N_12750,N_12752,N_12754,N_12755,N_12756,N_12757,N_12759,N_12760,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12772,N_12774,N_12775,N_12776,N_12778,N_12779,N_12780,N_12782,N_12783,N_12784,N_12785,N_12787,N_12791,N_12792,N_12793,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12832,N_12833,N_12834,N_12835,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12867,N_12868,N_12869,N_12870,N_12871,N_12874,N_12875,N_12876,N_12878,N_12879,N_12880,N_12881,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12895,N_12897,N_12898,N_12899,N_12902,N_12903,N_12904,N_12905,N_12906,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12925,N_12926,N_12930,N_12931,N_12932,N_12933,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12958,N_12959,N_12960,N_12962,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12974,N_12975,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12989,N_12990,N_12991,N_12993,N_12995,N_12997,N_12998,N_13000,N_13001,N_13002,N_13005,N_13007,N_13008,N_13009,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13028,N_13029,N_13030,N_13031,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13042,N_13043,N_13044,N_13045,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13066,N_13068,N_13069,N_13070,N_13072,N_13074,N_13077,N_13080,N_13081,N_13082,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13128,N_13129,N_13130,N_13131,N_13132,N_13134,N_13135,N_13136,N_13137,N_13138,N_13140,N_13141,N_13143,N_13144,N_13145,N_13146,N_13148,N_13149,N_13151,N_13153,N_13154,N_13156,N_13157,N_13158,N_13160,N_13161,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13172,N_13173,N_13176,N_13177,N_13178,N_13179,N_13180,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13202,N_13203,N_13204,N_13205,N_13206,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13218,N_13220,N_13221,N_13223,N_13224,N_13225,N_13226,N_13227,N_13229,N_13230,N_13231,N_13232,N_13233,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13248,N_13249,N_13250,N_13251,N_13253,N_13254,N_13255,N_13256,N_13258,N_13259,N_13260,N_13261,N_13263,N_13264,N_13265,N_13267,N_13268,N_13270,N_13272,N_13274,N_13275,N_13276,N_13277,N_13280,N_13281,N_13282,N_13285,N_13287,N_13288,N_13289,N_13290,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13309,N_13312,N_13314,N_13315,N_13317,N_13318,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13328,N_13329,N_13332,N_13333,N_13334,N_13335,N_13336,N_13338,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13417,N_13418,N_13419,N_13420,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13432,N_13433,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13490,N_13491,N_13492,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13527,N_13528,N_13530,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13548,N_13549,N_13551,N_13553,N_13555,N_13557,N_13559,N_13561,N_13562,N_13563,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13577,N_13578,N_13581,N_13582,N_13583,N_13584,N_13586,N_13587,N_13588,N_13589,N_13591,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13604,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13617,N_13618,N_13619,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13628,N_13630,N_13631,N_13632,N_13633,N_13635,N_13637,N_13638,N_13639,N_13641,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13670,N_13671,N_13672,N_13673,N_13674,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13690,N_13692,N_13693,N_13698,N_13700,N_13701,N_13702,N_13703,N_13704,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13715,N_13716,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13746,N_13747,N_13750,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13762,N_13763,N_13764,N_13766,N_13767,N_13768,N_13770,N_13771,N_13773,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13822,N_13824,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13847,N_13848,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13858,N_13860,N_13862,N_13863,N_13865,N_13866,N_13868,N_13870,N_13872,N_13874,N_13875,N_13876,N_13878,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13889,N_13893,N_13894,N_13896,N_13897,N_13898,N_13899,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13928,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13954,N_13955,N_13956,N_13958,N_13959,N_13960,N_13961,N_13963,N_13965,N_13966,N_13967,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13990,N_13991,N_13992,N_13993,N_13994,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14021,N_14022,N_14023,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14040,N_14041,N_14042,N_14043,N_14044,N_14046,N_14047,N_14048,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14065,N_14066,N_14067,N_14069,N_14070,N_14071,N_14072,N_14075,N_14076,N_14077,N_14078,N_14080,N_14081,N_14082,N_14084,N_14085,N_14086,N_14087,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14102,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14114,N_14115,N_14116,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14125,N_14127,N_14128,N_14129,N_14130,N_14131,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14141,N_14142,N_14144,N_14145,N_14147,N_14148,N_14150,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14193,N_14194,N_14195,N_14197,N_14198,N_14200,N_14201,N_14202,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14212,N_14213,N_14214,N_14215,N_14216,N_14221,N_14223,N_14225,N_14228,N_14230,N_14231,N_14232,N_14233,N_14235,N_14236,N_14237,N_14238,N_14239,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14275,N_14277,N_14278,N_14279,N_14281,N_14283,N_14284,N_14285,N_14286,N_14287,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14331,N_14332,N_14333,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14342,N_14344,N_14345,N_14346,N_14350,N_14351,N_14352,N_14354,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14383,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14394,N_14395,N_14396,N_14397,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14429,N_14430,N_14431,N_14432,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14450,N_14451,N_14452,N_14453,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14462,N_14463,N_14464,N_14465,N_14467,N_14469,N_14471,N_14472,N_14474,N_14476,N_14477,N_14478,N_14479,N_14480,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14492,N_14493,N_14494,N_14496,N_14497,N_14498,N_14499,N_14500,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14517,N_14518,N_14519,N_14520,N_14521,N_14523,N_14524,N_14525,N_14527,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14543,N_14544,N_14545,N_14546,N_14547,N_14549,N_14550,N_14552,N_14553,N_14554,N_14555,N_14558,N_14560,N_14561,N_14563,N_14564,N_14565,N_14566,N_14568,N_14569,N_14570,N_14571,N_14572,N_14574,N_14575,N_14576,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14592,N_14594,N_14595,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14608,N_14609,N_14611,N_14612,N_14613,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14622,N_14623,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14639,N_14640,N_14641,N_14643,N_14644,N_14645,N_14646,N_14648,N_14649,N_14650,N_14652,N_14653,N_14654,N_14655,N_14657,N_14658,N_14660,N_14662,N_14663,N_14664,N_14666,N_14667,N_14668,N_14669,N_14671,N_14673,N_14674,N_14676,N_14678,N_14679,N_14680,N_14682,N_14683,N_14684,N_14685,N_14687,N_14688,N_14692,N_14693,N_14694,N_14695,N_14696,N_14698,N_14699,N_14700,N_14702,N_14705,N_14707,N_14708,N_14710,N_14711,N_14713,N_14714,N_14716,N_14717,N_14719,N_14721,N_14722,N_14723,N_14725,N_14726,N_14728,N_14729,N_14730,N_14732,N_14733,N_14734,N_14735,N_14736,N_14738,N_14739,N_14741,N_14742,N_14743,N_14744,N_14746,N_14747,N_14748,N_14750,N_14751,N_14752,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14773,N_14774,N_14775,N_14776,N_14777,N_14780,N_14782,N_14783,N_14784,N_14785,N_14787,N_14788,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14800,N_14801,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14811,N_14812,N_14814,N_14816,N_14817,N_14819,N_14821,N_14822,N_14825,N_14827,N_14828,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14870,N_14872,N_14873,N_14874,N_14875,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14889,N_14890,N_14891,N_14892,N_14893,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14915,N_14916,N_14917,N_14918,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14934,N_14935,N_14936,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14947,N_14948,N_14949,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14978,N_14979,N_14981,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998;
nand U0 (N_0,In_143,In_1238);
and U1 (N_1,In_416,In_764);
nand U2 (N_2,In_732,In_369);
xnor U3 (N_3,In_1168,In_1391);
or U4 (N_4,In_1,In_1453);
nand U5 (N_5,In_1184,In_623);
xnor U6 (N_6,In_1167,In_527);
or U7 (N_7,In_858,In_718);
nand U8 (N_8,In_550,In_429);
nand U9 (N_9,In_535,In_1328);
nor U10 (N_10,In_1215,In_90);
nand U11 (N_11,In_455,In_350);
and U12 (N_12,In_354,In_525);
or U13 (N_13,In_1091,In_456);
nand U14 (N_14,In_1400,In_1025);
xor U15 (N_15,In_1191,In_421);
and U16 (N_16,In_131,In_607);
nor U17 (N_17,In_1422,In_1231);
nand U18 (N_18,In_646,In_290);
or U19 (N_19,In_1244,In_577);
and U20 (N_20,In_393,In_1409);
xnor U21 (N_21,In_804,In_287);
or U22 (N_22,In_534,In_20);
xnor U23 (N_23,In_793,In_845);
and U24 (N_24,In_466,In_1175);
or U25 (N_25,In_89,In_282);
nor U26 (N_26,In_836,In_1476);
and U27 (N_27,In_1348,In_400);
nor U28 (N_28,In_986,In_553);
and U29 (N_29,In_1013,In_460);
and U30 (N_30,In_620,In_451);
xnor U31 (N_31,In_798,In_932);
xnor U32 (N_32,In_925,In_885);
nor U33 (N_33,In_255,In_486);
nor U34 (N_34,In_690,In_1464);
nand U35 (N_35,In_1102,In_1380);
nand U36 (N_36,In_1412,In_961);
and U37 (N_37,In_361,In_839);
and U38 (N_38,In_803,In_491);
nor U39 (N_39,In_9,In_928);
nor U40 (N_40,In_973,In_1126);
and U41 (N_41,In_1265,In_1252);
xnor U42 (N_42,In_907,In_568);
nor U43 (N_43,In_745,In_1301);
xor U44 (N_44,In_63,In_1163);
xnor U45 (N_45,In_992,In_502);
nor U46 (N_46,In_1200,In_1003);
xnor U47 (N_47,In_834,In_729);
and U48 (N_48,In_1250,In_373);
nor U49 (N_49,In_903,In_709);
nor U50 (N_50,In_326,In_641);
or U51 (N_51,In_999,In_711);
xor U52 (N_52,In_603,In_28);
xnor U53 (N_53,In_1179,In_1406);
or U54 (N_54,In_410,In_840);
or U55 (N_55,In_167,In_1486);
or U56 (N_56,In_450,In_128);
xnor U57 (N_57,In_1302,In_1341);
xnor U58 (N_58,In_1274,In_497);
and U59 (N_59,In_206,In_750);
xnor U60 (N_60,In_755,In_723);
xor U61 (N_61,In_774,In_257);
nor U62 (N_62,In_650,In_107);
or U63 (N_63,In_375,In_1236);
or U64 (N_64,In_125,In_526);
xnor U65 (N_65,In_698,In_906);
nand U66 (N_66,In_1034,In_913);
and U67 (N_67,In_1012,In_610);
and U68 (N_68,In_148,In_974);
and U69 (N_69,In_1386,In_1482);
and U70 (N_70,In_112,In_880);
xor U71 (N_71,In_580,In_504);
and U72 (N_72,In_1376,In_1128);
or U73 (N_73,In_675,In_1454);
nand U74 (N_74,In_592,In_1022);
nand U75 (N_75,In_949,In_1402);
nand U76 (N_76,In_1357,In_94);
xor U77 (N_77,In_1189,In_1460);
nor U78 (N_78,In_1450,In_1254);
nor U79 (N_79,In_1044,In_513);
nand U80 (N_80,In_588,In_1279);
and U81 (N_81,In_1067,In_707);
nand U82 (N_82,In_981,In_262);
nand U83 (N_83,In_1349,In_1056);
and U84 (N_84,In_1307,In_216);
xor U85 (N_85,In_1467,In_693);
xor U86 (N_86,In_1105,In_1240);
nor U87 (N_87,In_682,In_970);
or U88 (N_88,In_498,In_377);
or U89 (N_89,In_897,In_565);
or U90 (N_90,In_205,In_123);
nor U91 (N_91,In_780,In_855);
nand U92 (N_92,In_1408,In_226);
xor U93 (N_93,In_1288,In_298);
and U94 (N_94,In_976,In_1283);
nor U95 (N_95,In_1031,In_426);
and U96 (N_96,In_166,In_1083);
nor U97 (N_97,In_1473,In_895);
and U98 (N_98,In_1130,In_4);
nand U99 (N_99,In_557,In_862);
and U100 (N_100,In_637,In_263);
nand U101 (N_101,In_83,In_242);
nand U102 (N_102,In_408,In_1465);
xor U103 (N_103,In_1439,In_1181);
nand U104 (N_104,In_31,In_245);
or U105 (N_105,In_987,In_322);
nor U106 (N_106,In_86,In_1135);
or U107 (N_107,In_1077,In_315);
nand U108 (N_108,In_1227,In_339);
nand U109 (N_109,In_878,In_1214);
nand U110 (N_110,In_401,In_399);
nand U111 (N_111,In_622,In_1363);
nor U112 (N_112,In_26,In_964);
nand U113 (N_113,In_582,In_473);
nand U114 (N_114,In_1498,In_149);
nor U115 (N_115,In_1143,In_998);
or U116 (N_116,In_52,In_859);
nand U117 (N_117,In_10,In_267);
nand U118 (N_118,In_1293,In_448);
nand U119 (N_119,In_1272,In_1196);
and U120 (N_120,In_499,In_76);
nor U121 (N_121,In_307,In_1441);
or U122 (N_122,In_864,In_816);
or U123 (N_123,In_822,In_278);
nand U124 (N_124,In_389,In_1392);
or U125 (N_125,In_27,In_1037);
and U126 (N_126,In_630,In_1212);
xor U127 (N_127,In_1120,In_1187);
xnor U128 (N_128,In_746,In_922);
xor U129 (N_129,In_464,In_483);
nor U130 (N_130,In_276,In_967);
xnor U131 (N_131,In_501,In_585);
or U132 (N_132,In_1074,In_325);
and U133 (N_133,In_977,In_1309);
xnor U134 (N_134,In_405,In_1149);
nand U135 (N_135,In_178,In_666);
nor U136 (N_136,In_1193,In_1417);
xor U137 (N_137,In_576,In_457);
nor U138 (N_138,In_789,In_215);
and U139 (N_139,In_1389,In_1388);
xnor U140 (N_140,In_1308,In_902);
nor U141 (N_141,In_312,In_1014);
xnor U142 (N_142,In_1242,In_681);
xnor U143 (N_143,In_1041,In_1033);
xnor U144 (N_144,In_697,In_289);
xnor U145 (N_145,In_657,In_514);
nand U146 (N_146,In_861,In_1073);
nand U147 (N_147,In_1321,In_760);
nor U148 (N_148,In_1269,In_911);
nor U149 (N_149,In_940,In_296);
nor U150 (N_150,In_1222,In_614);
and U151 (N_151,In_715,In_1375);
nor U152 (N_152,In_643,In_1239);
and U153 (N_153,In_119,In_394);
nor U154 (N_154,In_1451,In_459);
or U155 (N_155,In_13,In_1416);
xnor U156 (N_156,In_108,In_220);
xnor U157 (N_157,In_97,In_1413);
xnor U158 (N_158,In_1267,In_265);
nand U159 (N_159,In_32,In_333);
nor U160 (N_160,In_351,In_190);
or U161 (N_161,In_484,In_806);
nor U162 (N_162,In_856,In_705);
and U163 (N_163,In_712,In_1371);
xor U164 (N_164,In_628,In_635);
xor U165 (N_165,In_590,In_1355);
nor U166 (N_166,In_342,In_285);
xor U167 (N_167,In_1468,In_113);
and U168 (N_168,In_275,In_213);
xnor U169 (N_169,In_1090,In_1327);
or U170 (N_170,In_587,In_560);
xnor U171 (N_171,In_1496,In_337);
nor U172 (N_172,In_863,In_321);
and U173 (N_173,In_1393,In_1069);
nand U174 (N_174,In_161,In_243);
or U175 (N_175,In_1347,In_765);
or U176 (N_176,In_1049,In_184);
nand U177 (N_177,In_417,In_567);
and U178 (N_178,In_1230,In_367);
nor U179 (N_179,In_739,In_1206);
xor U180 (N_180,In_602,In_432);
and U181 (N_181,In_1152,In_777);
or U182 (N_182,In_923,In_554);
xor U183 (N_183,In_542,In_909);
and U184 (N_184,In_1286,In_236);
nand U185 (N_185,In_1436,In_500);
xnor U186 (N_186,In_615,In_1491);
nand U187 (N_187,In_562,In_767);
xor U188 (N_188,In_1334,In_831);
and U189 (N_189,In_629,In_713);
or U190 (N_190,In_1195,In_42);
nor U191 (N_191,In_1499,In_966);
or U192 (N_192,In_202,In_430);
nand U193 (N_193,In_1338,In_155);
xnor U194 (N_194,In_843,In_1111);
nand U195 (N_195,In_176,In_479);
and U196 (N_196,In_523,In_933);
xor U197 (N_197,In_211,In_978);
xor U198 (N_198,In_934,In_868);
or U199 (N_199,In_191,In_838);
xnor U200 (N_200,In_329,In_980);
and U201 (N_201,In_876,In_704);
xor U202 (N_202,In_120,In_1125);
xor U203 (N_203,In_382,In_1364);
and U204 (N_204,In_726,In_84);
nor U205 (N_205,In_154,In_699);
nor U206 (N_206,In_1407,In_1373);
and U207 (N_207,In_496,In_511);
nand U208 (N_208,In_355,In_638);
nand U209 (N_209,In_1018,In_81);
nand U210 (N_210,In_422,In_660);
xor U211 (N_211,In_988,In_334);
or U212 (N_212,In_1114,In_208);
and U213 (N_213,In_538,In_25);
or U214 (N_214,In_1220,In_468);
and U215 (N_215,In_1146,In_30);
nor U216 (N_216,In_366,In_872);
nor U217 (N_217,In_33,In_1352);
and U218 (N_218,In_174,In_1054);
nand U219 (N_219,In_1161,In_67);
or U220 (N_220,In_280,In_1367);
nor U221 (N_221,In_311,In_809);
nand U222 (N_222,In_165,In_345);
nor U223 (N_223,In_1124,In_291);
and U224 (N_224,In_412,In_874);
xnor U225 (N_225,In_207,In_1481);
or U226 (N_226,In_331,In_1160);
nand U227 (N_227,In_1428,In_571);
and U228 (N_228,In_655,In_1194);
nor U229 (N_229,In_153,In_871);
or U230 (N_230,In_23,In_182);
xor U231 (N_231,In_805,In_1213);
nor U232 (N_232,In_595,In_1462);
xor U233 (N_233,In_1285,In_1109);
nand U234 (N_234,In_1106,In_505);
or U235 (N_235,In_49,In_1245);
nor U236 (N_236,In_714,In_304);
xor U237 (N_237,In_229,In_17);
nand U238 (N_238,In_972,In_672);
nor U239 (N_239,In_144,In_293);
nand U240 (N_240,In_75,In_54);
nand U241 (N_241,In_1058,In_1035);
xnor U242 (N_242,In_270,In_612);
or U243 (N_243,In_1081,In_995);
or U244 (N_244,In_440,In_792);
or U245 (N_245,In_277,In_135);
xor U246 (N_246,In_1387,In_1221);
xor U247 (N_247,In_1353,In_685);
nor U248 (N_248,In_1061,In_71);
and U249 (N_249,In_1317,In_730);
or U250 (N_250,In_258,In_1336);
and U251 (N_251,In_1397,In_198);
nand U252 (N_252,In_1438,In_1185);
xnor U253 (N_253,In_230,In_536);
or U254 (N_254,In_575,In_1472);
nand U255 (N_255,In_41,In_636);
and U256 (N_256,In_555,In_124);
and U257 (N_257,In_520,In_844);
and U258 (N_258,In_842,In_1243);
nor U259 (N_259,In_45,In_1378);
nor U260 (N_260,In_952,In_327);
nand U261 (N_261,In_316,In_1010);
nor U262 (N_262,In_37,In_80);
nor U263 (N_263,In_398,In_1411);
nor U264 (N_264,In_702,In_1000);
nand U265 (N_265,In_100,In_461);
or U266 (N_266,In_1414,In_983);
xor U267 (N_267,In_1396,In_317);
nand U268 (N_268,In_1095,In_1237);
nor U269 (N_269,In_383,In_644);
and U270 (N_270,In_1419,In_971);
nand U271 (N_271,In_1026,In_683);
nor U272 (N_272,In_887,In_181);
and U273 (N_273,In_1062,In_252);
xnor U274 (N_274,In_259,In_1088);
nand U275 (N_275,In_727,In_943);
or U276 (N_276,In_541,In_938);
nor U277 (N_277,In_708,In_662);
nor U278 (N_278,In_810,In_665);
and U279 (N_279,In_1270,In_543);
nor U280 (N_280,In_1110,In_1322);
nand U281 (N_281,In_1326,In_141);
nor U282 (N_282,In_1350,In_801);
or U283 (N_283,In_766,In_1379);
and U284 (N_284,In_458,In_990);
xnor U285 (N_285,In_1292,In_758);
nor U286 (N_286,In_893,In_435);
nand U287 (N_287,In_668,In_982);
xnor U288 (N_288,In_589,In_60);
xor U289 (N_289,In_378,In_892);
nor U290 (N_290,In_508,In_1178);
and U291 (N_291,In_1123,In_619);
nor U292 (N_292,In_101,In_177);
xnor U293 (N_293,In_867,In_1115);
and U294 (N_294,In_1209,In_748);
xor U295 (N_295,In_1192,In_1471);
nand U296 (N_296,In_1296,In_658);
and U297 (N_297,In_1087,In_1147);
nor U298 (N_298,In_1346,In_480);
nor U299 (N_299,In_1268,In_1188);
or U300 (N_300,In_1040,In_1430);
xnor U301 (N_301,In_1009,In_487);
nor U302 (N_302,In_1100,In_1289);
nor U303 (N_303,In_688,In_736);
xor U304 (N_304,In_656,In_1199);
or U305 (N_305,In_1170,In_340);
and U306 (N_306,In_370,In_1097);
and U307 (N_307,In_5,In_21);
nor U308 (N_308,In_437,In_96);
nand U309 (N_309,In_545,In_443);
nand U310 (N_310,In_808,In_826);
nand U311 (N_311,In_376,In_477);
nor U312 (N_312,In_139,In_667);
and U313 (N_313,In_731,In_881);
or U314 (N_314,In_427,In_406);
nand U315 (N_315,In_1071,In_1226);
nand U316 (N_316,In_882,In_1306);
nor U317 (N_317,In_1131,In_960);
xnor U318 (N_318,In_1197,In_953);
nand U319 (N_319,In_824,In_1136);
or U320 (N_320,In_1113,In_414);
and U321 (N_321,In_899,In_817);
or U322 (N_322,In_1039,In_652);
xnor U323 (N_323,In_770,In_795);
xnor U324 (N_324,In_36,In_1461);
xnor U325 (N_325,In_1314,In_55);
nor U326 (N_326,In_945,In_719);
and U327 (N_327,In_146,In_95);
nor U328 (N_328,In_627,In_1047);
xor U329 (N_329,In_1165,In_546);
and U330 (N_330,In_1258,In_1052);
and U331 (N_331,In_330,In_1162);
xor U332 (N_332,In_740,In_110);
and U333 (N_333,In_1080,In_1445);
xnor U334 (N_334,In_1356,In_734);
or U335 (N_335,In_875,In_446);
and U336 (N_336,In_559,In_1219);
nor U337 (N_337,In_1410,In_1281);
or U338 (N_338,In_651,In_386);
nor U339 (N_339,In_1351,In_939);
nand U340 (N_340,In_196,In_156);
and U341 (N_341,In_916,In_232);
nand U342 (N_342,In_782,In_659);
xor U343 (N_343,In_528,In_762);
xnor U344 (N_344,In_1019,In_1365);
and U345 (N_345,In_14,In_1201);
xor U346 (N_346,In_185,In_495);
nand U347 (N_347,In_947,In_193);
nor U348 (N_348,In_465,In_424);
or U349 (N_349,In_1093,In_1133);
and U350 (N_350,In_1354,In_1295);
nor U351 (N_351,In_138,In_1028);
xnor U352 (N_352,In_1488,In_653);
xor U353 (N_353,In_1169,In_600);
xnor U354 (N_354,In_132,In_444);
and U355 (N_355,In_754,In_827);
xor U356 (N_356,In_954,In_1104);
and U357 (N_357,In_274,In_142);
nand U358 (N_358,In_791,In_975);
nor U359 (N_359,In_724,In_105);
nor U360 (N_360,In_1094,In_962);
and U361 (N_361,In_109,In_441);
or U362 (N_362,In_227,In_516);
nand U363 (N_363,In_1297,In_250);
nand U364 (N_364,In_811,In_905);
nor U365 (N_365,In_931,In_362);
or U366 (N_366,In_807,In_1177);
or U367 (N_367,In_1001,In_173);
and U368 (N_368,In_1493,In_1068);
nand U369 (N_369,In_187,In_676);
xor U370 (N_370,In_613,In_616);
nor U371 (N_371,In_941,In_771);
or U372 (N_372,In_1248,In_503);
or U373 (N_373,In_512,In_233);
or U374 (N_374,In_896,In_201);
xnor U375 (N_375,In_159,In_551);
xnor U376 (N_376,In_910,In_716);
or U377 (N_377,In_639,In_122);
nand U378 (N_378,In_833,In_515);
nor U379 (N_379,In_991,In_1429);
nor U380 (N_380,In_984,In_492);
and U381 (N_381,In_209,In_873);
nor U382 (N_382,In_56,In_244);
nor U383 (N_383,In_1036,In_162);
xor U384 (N_384,In_1256,In_157);
or U385 (N_385,In_749,In_283);
and U386 (N_386,In_929,In_1435);
and U387 (N_387,In_7,In_348);
or U388 (N_388,In_46,In_1275);
or U389 (N_389,In_419,In_15);
nand U390 (N_390,In_314,In_677);
or U391 (N_391,In_415,In_1107);
xor U392 (N_392,In_829,In_788);
and U393 (N_393,In_781,In_175);
nand U394 (N_394,In_832,In_1086);
nor U395 (N_395,In_609,In_372);
nor U396 (N_396,In_761,In_1372);
nand U397 (N_397,In_103,In_823);
and U398 (N_398,In_865,In_469);
xnor U399 (N_399,In_169,In_720);
or U400 (N_400,In_735,In_1335);
and U401 (N_401,In_1051,In_1023);
and U402 (N_402,In_1207,In_957);
nor U403 (N_403,In_336,In_747);
nor U404 (N_404,In_308,In_320);
or U405 (N_405,In_583,In_790);
nand U406 (N_406,In_219,In_1385);
or U407 (N_407,In_1190,In_1315);
or U408 (N_408,In_1112,In_106);
and U409 (N_409,In_737,In_578);
or U410 (N_410,In_261,In_87);
xnor U411 (N_411,In_203,In_886);
and U412 (N_412,In_59,In_1145);
and U413 (N_413,In_249,In_671);
or U414 (N_414,In_194,In_847);
nor U415 (N_415,In_150,In_349);
xor U416 (N_416,In_381,In_848);
xor U417 (N_417,In_489,In_596);
nand U418 (N_418,In_1029,In_379);
nor U419 (N_419,In_359,In_454);
xnor U420 (N_420,In_1487,In_1440);
or U421 (N_421,In_294,In_347);
or U422 (N_422,In_1134,In_1017);
or U423 (N_423,In_684,In_1007);
or U424 (N_424,In_920,In_2);
nor U425 (N_425,In_1173,In_1470);
nand U426 (N_426,In_1452,In_524);
or U427 (N_427,In_830,In_130);
nand U428 (N_428,In_396,In_1273);
or U429 (N_429,In_1425,In_1316);
nor U430 (N_430,In_212,In_1057);
xnor U431 (N_431,In_1300,In_1304);
nor U432 (N_432,In_621,In_670);
xnor U433 (N_433,In_678,In_915);
nor U434 (N_434,In_384,In_338);
nand U435 (N_435,In_1024,In_218);
nand U436 (N_436,In_140,In_1280);
xor U437 (N_437,In_266,In_1381);
and U438 (N_438,In_738,In_1103);
or U439 (N_439,In_1490,In_279);
and U440 (N_440,In_1427,In_281);
or U441 (N_441,In_11,In_1497);
or U442 (N_442,In_703,In_579);
nor U443 (N_443,In_195,In_968);
or U444 (N_444,In_1426,In_428);
or U445 (N_445,In_323,In_1383);
nor U446 (N_446,In_357,In_1132);
nor U447 (N_447,In_1478,In_1159);
or U448 (N_448,In_433,In_1183);
nor U449 (N_449,In_180,In_784);
or U450 (N_450,In_1455,In_70);
nor U451 (N_451,In_111,In_204);
or U452 (N_452,In_1064,In_318);
nand U453 (N_453,In_365,In_701);
or U454 (N_454,In_721,In_57);
or U455 (N_455,In_533,In_1443);
nor U456 (N_456,In_1399,In_385);
and U457 (N_457,In_127,In_388);
or U458 (N_458,In_1305,In_888);
and U459 (N_459,In_1101,In_946);
xor U460 (N_460,In_1072,In_134);
and U461 (N_461,In_1198,In_1089);
and U462 (N_462,In_854,In_300);
nor U463 (N_463,In_796,In_183);
nand U464 (N_464,In_558,In_241);
or U465 (N_465,In_402,In_1078);
and U466 (N_466,In_210,In_114);
or U467 (N_467,In_605,In_692);
and U468 (N_468,In_825,In_772);
nand U469 (N_469,In_392,In_246);
nor U470 (N_470,In_1144,In_403);
nand U471 (N_471,In_695,In_1312);
or U472 (N_472,In_472,In_1202);
nand U473 (N_473,In_358,In_1311);
nor U474 (N_474,In_1475,In_1489);
and U475 (N_475,In_561,In_442);
xnor U476 (N_476,In_1483,In_564);
nand U477 (N_477,In_380,In_769);
or U478 (N_478,In_591,In_1290);
xnor U479 (N_479,In_189,In_1480);
or U480 (N_480,In_1318,In_1038);
or U481 (N_481,In_937,In_908);
nand U482 (N_482,In_794,In_663);
nor U483 (N_483,In_725,In_785);
or U484 (N_484,In_1232,In_1186);
nor U485 (N_485,In_186,In_518);
nor U486 (N_486,In_238,In_260);
or U487 (N_487,In_69,In_813);
and U488 (N_488,In_919,In_481);
and U489 (N_489,In_1447,In_673);
and U490 (N_490,In_1148,In_642);
nand U491 (N_491,In_231,In_664);
nand U492 (N_492,In_1053,In_951);
xnor U493 (N_493,In_625,In_253);
nor U494 (N_494,In_1449,In_118);
nand U495 (N_495,In_1362,In_1174);
xnor U496 (N_496,In_1127,In_530);
and U497 (N_497,In_507,In_835);
or U498 (N_498,In_1154,In_356);
xnor U499 (N_499,In_1431,In_99);
and U500 (N_500,In_1359,In_1138);
and U501 (N_501,In_470,In_640);
nand U502 (N_502,In_164,In_759);
or U503 (N_503,In_857,In_1405);
or U504 (N_504,In_1343,In_1377);
or U505 (N_505,In_741,In_395);
xor U506 (N_506,In_462,In_237);
and U507 (N_507,In_818,In_234);
and U508 (N_508,In_171,In_837);
xor U509 (N_509,In_299,In_1277);
xor U510 (N_510,In_420,In_1298);
or U511 (N_511,In_1050,In_319);
or U512 (N_512,In_944,In_531);
or U513 (N_513,In_669,In_1070);
and U514 (N_514,In_593,In_1004);
or U515 (N_515,In_846,In_1055);
nand U516 (N_516,In_1218,In_1263);
and U517 (N_517,In_1344,In_1259);
xnor U518 (N_518,In_1276,In_1329);
and U519 (N_519,In_522,In_490);
xor U520 (N_520,In_851,In_529);
nand U521 (N_521,In_1030,In_269);
xnor U522 (N_522,In_1457,In_996);
nand U523 (N_523,In_1182,In_1437);
or U524 (N_524,In_544,In_1368);
nand U525 (N_525,In_256,In_918);
nor U526 (N_526,In_66,In_1108);
or U527 (N_527,In_264,In_295);
nand U528 (N_528,In_517,In_390);
nor U529 (N_529,In_869,In_573);
and U530 (N_530,In_624,In_598);
xor U531 (N_531,In_1217,In_1361);
nor U532 (N_532,In_301,In_43);
nand U533 (N_533,In_661,In_92);
xnor U534 (N_534,In_137,In_1158);
or U535 (N_535,In_305,In_1032);
and U536 (N_536,In_223,In_1059);
xnor U537 (N_537,In_849,In_1261);
nor U538 (N_538,In_548,In_228);
nor U539 (N_539,In_1172,In_439);
nand U540 (N_540,In_284,In_78);
and U541 (N_541,In_29,In_547);
nor U542 (N_542,In_1176,In_1085);
xor U543 (N_543,In_993,In_493);
and U544 (N_544,In_1210,In_1042);
xnor U545 (N_545,In_800,In_799);
or U546 (N_546,In_292,In_574);
nor U547 (N_547,In_434,In_956);
nor U548 (N_548,In_958,In_654);
or U549 (N_549,In_1117,In_1271);
xor U550 (N_550,In_1291,In_597);
nand U551 (N_551,In_1092,In_1096);
and U552 (N_552,In_1456,In_728);
and U553 (N_553,In_1313,In_706);
xnor U554 (N_554,In_1398,In_942);
or U555 (N_555,In_853,In_1339);
xor U556 (N_556,In_632,In_1079);
xor U557 (N_557,In_617,In_51);
nand U558 (N_558,In_891,In_1224);
nand U559 (N_559,In_40,In_532);
or U560 (N_560,In_634,In_1142);
and U561 (N_561,In_1141,In_1340);
xnor U562 (N_562,In_1332,In_53);
nor U563 (N_563,In_775,In_569);
and U564 (N_564,In_452,In_570);
xor U565 (N_565,In_313,In_6);
nand U566 (N_566,In_647,In_586);
nand U567 (N_567,In_539,In_18);
nand U568 (N_568,In_1229,In_552);
and U569 (N_569,In_352,In_332);
or U570 (N_570,In_158,In_116);
and U571 (N_571,In_324,In_776);
and U572 (N_572,In_763,In_900);
xnor U573 (N_573,In_1404,In_1374);
nor U574 (N_574,In_1204,In_303);
xor U575 (N_575,In_1171,In_679);
or U576 (N_576,In_271,In_841);
and U577 (N_577,In_965,In_815);
or U578 (N_578,In_1005,In_272);
nand U579 (N_579,In_540,In_1046);
and U580 (N_580,In_969,In_884);
xnor U581 (N_581,In_91,In_409);
and U582 (N_582,In_779,In_773);
or U583 (N_583,In_268,In_914);
and U584 (N_584,In_733,In_1099);
and U585 (N_585,In_22,In_1423);
and U586 (N_586,In_1045,In_136);
nor U587 (N_587,In_1401,In_626);
nor U588 (N_588,In_618,In_1211);
nor U589 (N_589,In_72,In_449);
or U590 (N_590,In_168,In_1284);
nor U591 (N_591,In_1260,In_0);
or U592 (N_592,In_753,In_649);
xor U593 (N_593,In_648,In_1234);
xor U594 (N_594,In_1008,In_1485);
nor U595 (N_595,In_1139,In_1157);
or U596 (N_596,In_1390,In_1325);
nor U597 (N_597,In_1477,In_133);
nand U598 (N_598,In_1394,In_752);
and U599 (N_599,In_254,In_935);
and U600 (N_600,In_1180,In_1006);
nor U601 (N_601,In_1249,In_286);
nor U602 (N_602,In_475,In_147);
nor U603 (N_603,In_1156,In_1333);
and U604 (N_604,In_47,In_68);
or U605 (N_605,In_1384,In_1303);
xor U606 (N_606,In_963,In_488);
or U607 (N_607,In_368,In_1420);
nor U608 (N_608,In_64,In_494);
or U609 (N_609,In_606,In_870);
nor U610 (N_610,In_221,In_1122);
or U611 (N_611,In_1282,In_537);
nand U612 (N_612,In_1233,In_1076);
nor U613 (N_613,In_199,In_904);
nand U614 (N_614,In_1366,In_1016);
xnor U615 (N_615,In_756,In_1020);
or U616 (N_616,In_1002,In_757);
or U617 (N_617,In_877,In_674);
nor U618 (N_618,In_1137,In_1063);
nor U619 (N_619,In_599,In_1255);
or U620 (N_620,In_611,In_431);
and U621 (N_621,In_35,In_438);
nand U622 (N_622,In_482,In_251);
xnor U623 (N_623,In_222,In_572);
or U624 (N_624,In_411,In_344);
nand U625 (N_625,In_88,In_1494);
and U626 (N_626,In_1021,In_549);
or U627 (N_627,In_73,In_1320);
nor U628 (N_628,In_820,In_170);
or U629 (N_629,In_476,In_364);
and U630 (N_630,In_200,In_104);
nor U631 (N_631,In_48,In_12);
and U632 (N_632,In_997,In_288);
and U633 (N_633,In_802,In_85);
nor U634 (N_634,In_1205,In_1246);
xnor U635 (N_635,In_328,In_61);
xor U636 (N_636,In_160,In_994);
or U637 (N_637,In_1319,In_1415);
nand U638 (N_638,In_1082,In_584);
nor U639 (N_639,In_1121,In_423);
and U640 (N_640,In_79,In_1264);
and U641 (N_641,In_297,In_407);
nand U642 (N_642,In_926,In_1155);
and U643 (N_643,In_787,In_1424);
xnor U644 (N_644,In_1358,In_744);
xnor U645 (N_645,In_302,In_510);
nor U646 (N_646,In_687,In_1474);
nor U647 (N_647,In_273,In_1075);
xnor U648 (N_648,In_927,In_235);
nand U649 (N_649,In_74,In_786);
or U650 (N_650,In_1098,In_1382);
nor U651 (N_651,In_117,In_309);
nor U652 (N_652,In_601,In_239);
nand U653 (N_653,In_8,In_34);
or U654 (N_654,In_192,In_989);
and U655 (N_655,In_115,In_604);
nand U656 (N_656,In_645,In_3);
nor U657 (N_657,In_306,In_743);
nor U658 (N_658,In_519,In_1043);
nand U659 (N_659,In_1466,In_224);
or U660 (N_660,In_1418,In_371);
nor U661 (N_661,In_39,In_485);
xor U662 (N_662,In_1403,In_563);
xnor U663 (N_663,In_1360,In_797);
or U664 (N_664,In_1262,In_509);
or U665 (N_665,In_360,In_581);
and U666 (N_666,In_247,In_248);
nand U667 (N_667,In_812,In_948);
or U668 (N_668,In_889,In_121);
xor U669 (N_669,In_310,In_1266);
nor U670 (N_670,In_850,In_1150);
or U671 (N_671,In_346,In_917);
or U672 (N_672,In_1370,In_1287);
xor U673 (N_673,In_1208,In_413);
and U674 (N_674,In_1065,In_1469);
and U675 (N_675,In_24,In_1444);
xnor U676 (N_676,In_391,In_1310);
nor U677 (N_677,In_1060,In_1048);
or U678 (N_678,In_343,In_1432);
and U679 (N_679,In_1223,In_852);
or U680 (N_680,In_1324,In_521);
or U681 (N_681,In_1299,In_710);
nand U682 (N_682,In_985,In_751);
or U683 (N_683,In_1369,In_374);
nor U684 (N_684,In_879,In_633);
or U685 (N_685,In_631,In_930);
nor U686 (N_686,In_172,In_921);
and U687 (N_687,In_463,In_1084);
nand U688 (N_688,In_1458,In_717);
xnor U689 (N_689,In_38,In_680);
and U690 (N_690,In_694,In_1479);
or U691 (N_691,In_608,In_474);
nor U692 (N_692,In_1342,In_197);
nand U693 (N_693,In_1294,In_1119);
and U694 (N_694,In_467,In_447);
or U695 (N_695,In_1434,In_1164);
nand U696 (N_696,In_1446,In_1241);
nand U697 (N_697,In_151,In_1323);
or U698 (N_698,In_936,In_397);
nand U699 (N_699,In_890,In_866);
xor U700 (N_700,In_1151,In_217);
nand U701 (N_701,In_179,In_1216);
or U702 (N_702,In_979,In_418);
xnor U703 (N_703,In_686,In_959);
and U704 (N_704,In_82,In_445);
and U705 (N_705,In_506,In_912);
or U706 (N_706,In_1166,In_924);
nor U707 (N_707,In_1484,In_1463);
and U708 (N_708,In_1459,In_1253);
and U709 (N_709,In_1395,In_1448);
nand U710 (N_710,In_901,In_335);
and U711 (N_711,In_353,In_188);
xnor U712 (N_712,In_1337,In_387);
nand U713 (N_713,In_1235,In_955);
nor U714 (N_714,In_819,In_768);
nor U715 (N_715,In_1153,In_828);
nor U716 (N_716,In_145,In_742);
nor U717 (N_717,In_152,In_65);
and U718 (N_718,In_58,In_240);
or U719 (N_719,In_814,In_126);
nand U720 (N_720,In_566,In_594);
or U721 (N_721,In_1251,In_883);
and U722 (N_722,In_1278,In_556);
nand U723 (N_723,In_950,In_16);
nand U724 (N_724,In_1345,In_77);
or U725 (N_725,In_689,In_1433);
xor U726 (N_726,In_860,In_696);
nor U727 (N_727,In_1331,In_214);
and U728 (N_728,In_894,In_436);
nand U729 (N_729,In_1027,In_1140);
nor U730 (N_730,In_62,In_341);
nor U731 (N_731,In_1129,In_471);
xor U732 (N_732,In_1492,In_1011);
xnor U733 (N_733,In_129,In_691);
nand U734 (N_734,In_1118,In_1330);
xnor U735 (N_735,In_1495,In_1203);
xnor U736 (N_736,In_98,In_425);
or U737 (N_737,In_1442,In_93);
nor U738 (N_738,In_404,In_44);
or U739 (N_739,In_19,In_783);
nand U740 (N_740,In_102,In_778);
or U741 (N_741,In_722,In_1066);
and U742 (N_742,In_478,In_821);
and U743 (N_743,In_363,In_898);
or U744 (N_744,In_1225,In_225);
nor U745 (N_745,In_1015,In_1247);
nor U746 (N_746,In_163,In_1228);
and U747 (N_747,In_1257,In_1116);
and U748 (N_748,In_1421,In_50);
or U749 (N_749,In_453,In_700);
or U750 (N_750,In_316,In_1079);
or U751 (N_751,In_51,In_750);
xor U752 (N_752,In_350,In_996);
and U753 (N_753,In_673,In_1352);
nand U754 (N_754,In_1206,In_471);
nand U755 (N_755,In_166,In_519);
nand U756 (N_756,In_487,In_636);
xnor U757 (N_757,In_1444,In_121);
nand U758 (N_758,In_300,In_1008);
and U759 (N_759,In_273,In_1353);
xor U760 (N_760,In_491,In_515);
nor U761 (N_761,In_974,In_1417);
nor U762 (N_762,In_173,In_586);
nor U763 (N_763,In_561,In_30);
or U764 (N_764,In_212,In_336);
or U765 (N_765,In_842,In_1478);
nand U766 (N_766,In_1082,In_1352);
nor U767 (N_767,In_1050,In_624);
nand U768 (N_768,In_179,In_456);
and U769 (N_769,In_1006,In_669);
or U770 (N_770,In_884,In_965);
nor U771 (N_771,In_200,In_618);
xnor U772 (N_772,In_1411,In_659);
nand U773 (N_773,In_853,In_342);
nor U774 (N_774,In_609,In_499);
nand U775 (N_775,In_338,In_716);
nor U776 (N_776,In_669,In_468);
or U777 (N_777,In_1341,In_665);
nand U778 (N_778,In_55,In_417);
xor U779 (N_779,In_210,In_1436);
xnor U780 (N_780,In_74,In_114);
nand U781 (N_781,In_678,In_753);
xnor U782 (N_782,In_90,In_448);
or U783 (N_783,In_429,In_1334);
nor U784 (N_784,In_577,In_884);
and U785 (N_785,In_912,In_1411);
nand U786 (N_786,In_662,In_1430);
nor U787 (N_787,In_618,In_1015);
nand U788 (N_788,In_147,In_1453);
and U789 (N_789,In_1201,In_1489);
nor U790 (N_790,In_572,In_1144);
or U791 (N_791,In_97,In_621);
or U792 (N_792,In_181,In_298);
or U793 (N_793,In_193,In_218);
nand U794 (N_794,In_1463,In_626);
and U795 (N_795,In_888,In_122);
or U796 (N_796,In_621,In_1315);
nand U797 (N_797,In_192,In_23);
nor U798 (N_798,In_651,In_523);
nand U799 (N_799,In_1242,In_1257);
nor U800 (N_800,In_551,In_4);
and U801 (N_801,In_649,In_930);
nand U802 (N_802,In_647,In_765);
xor U803 (N_803,In_1301,In_889);
and U804 (N_804,In_672,In_382);
xnor U805 (N_805,In_260,In_1305);
or U806 (N_806,In_993,In_1070);
nor U807 (N_807,In_1115,In_863);
nor U808 (N_808,In_1137,In_1222);
nor U809 (N_809,In_1190,In_268);
nand U810 (N_810,In_334,In_788);
or U811 (N_811,In_788,In_1063);
nand U812 (N_812,In_561,In_168);
or U813 (N_813,In_1188,In_906);
xor U814 (N_814,In_694,In_600);
nand U815 (N_815,In_427,In_714);
and U816 (N_816,In_1239,In_1334);
or U817 (N_817,In_136,In_607);
nor U818 (N_818,In_1368,In_1299);
nand U819 (N_819,In_459,In_721);
nand U820 (N_820,In_989,In_366);
nor U821 (N_821,In_103,In_417);
xor U822 (N_822,In_396,In_1374);
nand U823 (N_823,In_739,In_538);
or U824 (N_824,In_114,In_1420);
xor U825 (N_825,In_345,In_1178);
nand U826 (N_826,In_580,In_942);
nand U827 (N_827,In_316,In_965);
or U828 (N_828,In_194,In_647);
nor U829 (N_829,In_644,In_440);
nand U830 (N_830,In_842,In_980);
xor U831 (N_831,In_819,In_1372);
or U832 (N_832,In_569,In_572);
xor U833 (N_833,In_81,In_536);
xnor U834 (N_834,In_361,In_472);
xor U835 (N_835,In_120,In_738);
xnor U836 (N_836,In_1083,In_411);
nand U837 (N_837,In_878,In_1222);
nand U838 (N_838,In_1218,In_1286);
or U839 (N_839,In_1311,In_1450);
nor U840 (N_840,In_852,In_1112);
nor U841 (N_841,In_337,In_945);
nor U842 (N_842,In_1261,In_901);
or U843 (N_843,In_1304,In_1418);
xor U844 (N_844,In_368,In_1463);
nor U845 (N_845,In_75,In_680);
and U846 (N_846,In_1149,In_991);
xnor U847 (N_847,In_1338,In_953);
nand U848 (N_848,In_863,In_360);
xnor U849 (N_849,In_6,In_981);
nand U850 (N_850,In_278,In_191);
and U851 (N_851,In_104,In_916);
nand U852 (N_852,In_992,In_1034);
xnor U853 (N_853,In_1478,In_424);
xnor U854 (N_854,In_747,In_149);
xnor U855 (N_855,In_1076,In_1362);
or U856 (N_856,In_412,In_1003);
or U857 (N_857,In_1024,In_674);
or U858 (N_858,In_1418,In_1310);
nor U859 (N_859,In_717,In_752);
nor U860 (N_860,In_303,In_575);
or U861 (N_861,In_211,In_1482);
xnor U862 (N_862,In_715,In_283);
nor U863 (N_863,In_1475,In_983);
and U864 (N_864,In_868,In_309);
xnor U865 (N_865,In_1440,In_54);
or U866 (N_866,In_177,In_1407);
and U867 (N_867,In_1102,In_632);
or U868 (N_868,In_1135,In_119);
xor U869 (N_869,In_616,In_1123);
nand U870 (N_870,In_280,In_491);
nand U871 (N_871,In_766,In_1469);
and U872 (N_872,In_282,In_1160);
or U873 (N_873,In_1124,In_225);
xnor U874 (N_874,In_325,In_1092);
nand U875 (N_875,In_1134,In_1404);
nor U876 (N_876,In_1316,In_589);
nor U877 (N_877,In_863,In_1017);
nand U878 (N_878,In_370,In_1063);
nand U879 (N_879,In_142,In_685);
xnor U880 (N_880,In_760,In_65);
and U881 (N_881,In_678,In_1242);
xor U882 (N_882,In_284,In_475);
xnor U883 (N_883,In_382,In_885);
nor U884 (N_884,In_1205,In_1184);
nor U885 (N_885,In_45,In_1193);
nand U886 (N_886,In_557,In_642);
nor U887 (N_887,In_780,In_749);
nor U888 (N_888,In_97,In_1309);
and U889 (N_889,In_502,In_917);
and U890 (N_890,In_365,In_1056);
nand U891 (N_891,In_808,In_101);
nand U892 (N_892,In_745,In_987);
nand U893 (N_893,In_105,In_1038);
nor U894 (N_894,In_1152,In_1072);
nand U895 (N_895,In_313,In_64);
xnor U896 (N_896,In_866,In_11);
or U897 (N_897,In_1153,In_24);
xor U898 (N_898,In_1183,In_987);
nand U899 (N_899,In_230,In_236);
and U900 (N_900,In_456,In_269);
nand U901 (N_901,In_335,In_1244);
or U902 (N_902,In_1408,In_69);
nand U903 (N_903,In_1237,In_512);
nand U904 (N_904,In_672,In_499);
or U905 (N_905,In_628,In_887);
nand U906 (N_906,In_870,In_1320);
nand U907 (N_907,In_1096,In_123);
nand U908 (N_908,In_67,In_1057);
nor U909 (N_909,In_385,In_1058);
xnor U910 (N_910,In_861,In_782);
and U911 (N_911,In_843,In_1104);
nand U912 (N_912,In_842,In_1359);
or U913 (N_913,In_811,In_884);
and U914 (N_914,In_206,In_330);
nor U915 (N_915,In_189,In_666);
xor U916 (N_916,In_567,In_217);
or U917 (N_917,In_1070,In_624);
or U918 (N_918,In_1354,In_254);
and U919 (N_919,In_1048,In_244);
xnor U920 (N_920,In_710,In_34);
or U921 (N_921,In_1430,In_320);
or U922 (N_922,In_382,In_517);
and U923 (N_923,In_848,In_499);
and U924 (N_924,In_727,In_1374);
nor U925 (N_925,In_20,In_49);
nand U926 (N_926,In_76,In_1316);
nand U927 (N_927,In_1082,In_1081);
xor U928 (N_928,In_1208,In_1243);
or U929 (N_929,In_1362,In_639);
nand U930 (N_930,In_694,In_909);
xnor U931 (N_931,In_606,In_412);
nor U932 (N_932,In_202,In_1486);
or U933 (N_933,In_1065,In_73);
or U934 (N_934,In_1323,In_1393);
xnor U935 (N_935,In_1256,In_141);
and U936 (N_936,In_38,In_874);
nand U937 (N_937,In_586,In_328);
nor U938 (N_938,In_1094,In_1246);
or U939 (N_939,In_42,In_155);
nor U940 (N_940,In_220,In_692);
and U941 (N_941,In_836,In_615);
nand U942 (N_942,In_1181,In_155);
nor U943 (N_943,In_498,In_1194);
xor U944 (N_944,In_351,In_329);
or U945 (N_945,In_961,In_339);
or U946 (N_946,In_764,In_513);
xnor U947 (N_947,In_614,In_1260);
nand U948 (N_948,In_277,In_1352);
nand U949 (N_949,In_1266,In_1289);
or U950 (N_950,In_707,In_921);
or U951 (N_951,In_510,In_1404);
nor U952 (N_952,In_1073,In_850);
or U953 (N_953,In_173,In_279);
nand U954 (N_954,In_656,In_1099);
xnor U955 (N_955,In_447,In_733);
and U956 (N_956,In_140,In_805);
xor U957 (N_957,In_100,In_1183);
xnor U958 (N_958,In_861,In_1304);
nor U959 (N_959,In_1160,In_193);
nor U960 (N_960,In_342,In_936);
and U961 (N_961,In_389,In_1462);
and U962 (N_962,In_1130,In_6);
xnor U963 (N_963,In_966,In_948);
xor U964 (N_964,In_373,In_1113);
nor U965 (N_965,In_70,In_211);
and U966 (N_966,In_1291,In_62);
and U967 (N_967,In_1196,In_827);
and U968 (N_968,In_510,In_832);
nand U969 (N_969,In_1210,In_1148);
nand U970 (N_970,In_377,In_651);
xor U971 (N_971,In_729,In_1359);
nand U972 (N_972,In_1496,In_198);
xnor U973 (N_973,In_95,In_832);
or U974 (N_974,In_996,In_142);
xnor U975 (N_975,In_538,In_574);
nand U976 (N_976,In_466,In_1126);
nand U977 (N_977,In_138,In_172);
and U978 (N_978,In_76,In_854);
or U979 (N_979,In_1082,In_105);
or U980 (N_980,In_500,In_215);
nor U981 (N_981,In_1178,In_1153);
nor U982 (N_982,In_1088,In_701);
nor U983 (N_983,In_188,In_311);
nand U984 (N_984,In_219,In_1171);
xnor U985 (N_985,In_233,In_911);
nand U986 (N_986,In_1474,In_1040);
or U987 (N_987,In_1250,In_1436);
nor U988 (N_988,In_481,In_25);
and U989 (N_989,In_129,In_952);
xnor U990 (N_990,In_1397,In_651);
nor U991 (N_991,In_695,In_1268);
nand U992 (N_992,In_339,In_1412);
or U993 (N_993,In_587,In_869);
nor U994 (N_994,In_601,In_752);
and U995 (N_995,In_1325,In_179);
xnor U996 (N_996,In_39,In_1101);
nand U997 (N_997,In_1415,In_1436);
nand U998 (N_998,In_87,In_565);
and U999 (N_999,In_782,In_1023);
nand U1000 (N_1000,In_1399,In_1488);
and U1001 (N_1001,In_699,In_87);
nor U1002 (N_1002,In_689,In_913);
nor U1003 (N_1003,In_1323,In_272);
and U1004 (N_1004,In_480,In_93);
xor U1005 (N_1005,In_850,In_958);
nor U1006 (N_1006,In_1071,In_1129);
nand U1007 (N_1007,In_413,In_1298);
and U1008 (N_1008,In_1042,In_1325);
nand U1009 (N_1009,In_246,In_1084);
nor U1010 (N_1010,In_1490,In_926);
or U1011 (N_1011,In_364,In_1215);
or U1012 (N_1012,In_1275,In_1287);
or U1013 (N_1013,In_718,In_388);
xor U1014 (N_1014,In_642,In_1183);
xnor U1015 (N_1015,In_256,In_702);
xnor U1016 (N_1016,In_102,In_433);
and U1017 (N_1017,In_1147,In_928);
nand U1018 (N_1018,In_83,In_21);
nor U1019 (N_1019,In_952,In_87);
and U1020 (N_1020,In_428,In_353);
xor U1021 (N_1021,In_215,In_43);
xnor U1022 (N_1022,In_1270,In_1140);
xor U1023 (N_1023,In_846,In_717);
nand U1024 (N_1024,In_785,In_1102);
nand U1025 (N_1025,In_351,In_1204);
and U1026 (N_1026,In_794,In_1496);
nor U1027 (N_1027,In_411,In_1086);
or U1028 (N_1028,In_422,In_1014);
or U1029 (N_1029,In_1157,In_979);
nor U1030 (N_1030,In_1181,In_858);
xnor U1031 (N_1031,In_1166,In_1149);
nor U1032 (N_1032,In_1096,In_497);
xnor U1033 (N_1033,In_420,In_1256);
xor U1034 (N_1034,In_829,In_1464);
nand U1035 (N_1035,In_677,In_1318);
or U1036 (N_1036,In_1207,In_647);
xor U1037 (N_1037,In_702,In_910);
or U1038 (N_1038,In_645,In_1242);
nand U1039 (N_1039,In_1025,In_365);
or U1040 (N_1040,In_1007,In_1032);
nor U1041 (N_1041,In_1252,In_789);
nor U1042 (N_1042,In_1152,In_602);
xnor U1043 (N_1043,In_164,In_11);
or U1044 (N_1044,In_800,In_1030);
nor U1045 (N_1045,In_382,In_1149);
xnor U1046 (N_1046,In_1329,In_1326);
nand U1047 (N_1047,In_1415,In_341);
xor U1048 (N_1048,In_12,In_584);
nor U1049 (N_1049,In_1269,In_1131);
nand U1050 (N_1050,In_296,In_366);
xor U1051 (N_1051,In_308,In_453);
or U1052 (N_1052,In_812,In_1310);
and U1053 (N_1053,In_91,In_25);
and U1054 (N_1054,In_1204,In_77);
nand U1055 (N_1055,In_1060,In_1494);
nand U1056 (N_1056,In_72,In_291);
or U1057 (N_1057,In_866,In_611);
nand U1058 (N_1058,In_778,In_78);
nand U1059 (N_1059,In_376,In_192);
or U1060 (N_1060,In_981,In_1460);
or U1061 (N_1061,In_231,In_1413);
and U1062 (N_1062,In_100,In_306);
nand U1063 (N_1063,In_238,In_1082);
and U1064 (N_1064,In_818,In_961);
nor U1065 (N_1065,In_195,In_1432);
or U1066 (N_1066,In_758,In_447);
nor U1067 (N_1067,In_1115,In_933);
nand U1068 (N_1068,In_583,In_656);
nor U1069 (N_1069,In_529,In_972);
xnor U1070 (N_1070,In_1307,In_876);
and U1071 (N_1071,In_998,In_833);
nand U1072 (N_1072,In_648,In_1220);
xnor U1073 (N_1073,In_532,In_404);
nand U1074 (N_1074,In_714,In_1245);
nand U1075 (N_1075,In_1342,In_947);
nor U1076 (N_1076,In_17,In_1406);
nand U1077 (N_1077,In_1066,In_238);
and U1078 (N_1078,In_1325,In_373);
xor U1079 (N_1079,In_1411,In_642);
or U1080 (N_1080,In_1239,In_525);
xnor U1081 (N_1081,In_1331,In_953);
or U1082 (N_1082,In_829,In_319);
and U1083 (N_1083,In_522,In_248);
nand U1084 (N_1084,In_796,In_1361);
nor U1085 (N_1085,In_1219,In_1290);
and U1086 (N_1086,In_553,In_815);
or U1087 (N_1087,In_911,In_1299);
xnor U1088 (N_1088,In_1264,In_957);
xor U1089 (N_1089,In_351,In_1320);
xor U1090 (N_1090,In_1055,In_237);
nor U1091 (N_1091,In_814,In_1114);
nor U1092 (N_1092,In_150,In_1139);
and U1093 (N_1093,In_518,In_475);
and U1094 (N_1094,In_683,In_127);
nor U1095 (N_1095,In_392,In_1208);
xnor U1096 (N_1096,In_766,In_310);
or U1097 (N_1097,In_358,In_455);
and U1098 (N_1098,In_61,In_1470);
or U1099 (N_1099,In_336,In_415);
nor U1100 (N_1100,In_76,In_1324);
or U1101 (N_1101,In_614,In_379);
xor U1102 (N_1102,In_1258,In_729);
xnor U1103 (N_1103,In_357,In_880);
or U1104 (N_1104,In_20,In_872);
xnor U1105 (N_1105,In_337,In_1121);
nor U1106 (N_1106,In_848,In_1319);
and U1107 (N_1107,In_95,In_1096);
or U1108 (N_1108,In_1349,In_1057);
xnor U1109 (N_1109,In_657,In_182);
nor U1110 (N_1110,In_517,In_800);
xor U1111 (N_1111,In_1179,In_1171);
nor U1112 (N_1112,In_1106,In_908);
xnor U1113 (N_1113,In_208,In_472);
nor U1114 (N_1114,In_1428,In_1079);
or U1115 (N_1115,In_892,In_1278);
xnor U1116 (N_1116,In_1456,In_79);
nand U1117 (N_1117,In_242,In_983);
xor U1118 (N_1118,In_898,In_659);
and U1119 (N_1119,In_522,In_879);
or U1120 (N_1120,In_975,In_1230);
nand U1121 (N_1121,In_99,In_30);
nor U1122 (N_1122,In_379,In_1461);
nor U1123 (N_1123,In_179,In_1086);
xnor U1124 (N_1124,In_672,In_1109);
and U1125 (N_1125,In_239,In_1419);
xnor U1126 (N_1126,In_206,In_661);
xnor U1127 (N_1127,In_1083,In_1105);
and U1128 (N_1128,In_804,In_1070);
nor U1129 (N_1129,In_1154,In_1397);
xnor U1130 (N_1130,In_1069,In_1196);
nand U1131 (N_1131,In_1079,In_1131);
nand U1132 (N_1132,In_255,In_87);
nand U1133 (N_1133,In_458,In_43);
and U1134 (N_1134,In_856,In_1394);
and U1135 (N_1135,In_1467,In_383);
xor U1136 (N_1136,In_955,In_878);
or U1137 (N_1137,In_1044,In_264);
or U1138 (N_1138,In_840,In_205);
or U1139 (N_1139,In_1066,In_130);
xor U1140 (N_1140,In_1271,In_87);
and U1141 (N_1141,In_1097,In_499);
and U1142 (N_1142,In_22,In_989);
nand U1143 (N_1143,In_1085,In_643);
xor U1144 (N_1144,In_44,In_222);
and U1145 (N_1145,In_940,In_1387);
nand U1146 (N_1146,In_1305,In_699);
and U1147 (N_1147,In_1472,In_1106);
or U1148 (N_1148,In_1214,In_1275);
xor U1149 (N_1149,In_942,In_789);
nand U1150 (N_1150,In_1202,In_1076);
nand U1151 (N_1151,In_491,In_1208);
xnor U1152 (N_1152,In_1136,In_535);
xnor U1153 (N_1153,In_408,In_393);
xor U1154 (N_1154,In_1047,In_1255);
and U1155 (N_1155,In_954,In_816);
and U1156 (N_1156,In_1315,In_789);
or U1157 (N_1157,In_100,In_1414);
and U1158 (N_1158,In_513,In_636);
and U1159 (N_1159,In_569,In_1058);
and U1160 (N_1160,In_674,In_185);
nand U1161 (N_1161,In_1318,In_964);
xor U1162 (N_1162,In_97,In_870);
nand U1163 (N_1163,In_382,In_417);
nor U1164 (N_1164,In_363,In_5);
or U1165 (N_1165,In_434,In_688);
or U1166 (N_1166,In_812,In_377);
nor U1167 (N_1167,In_734,In_758);
xnor U1168 (N_1168,In_578,In_796);
nor U1169 (N_1169,In_1309,In_248);
nor U1170 (N_1170,In_534,In_605);
nor U1171 (N_1171,In_12,In_462);
xor U1172 (N_1172,In_802,In_656);
or U1173 (N_1173,In_733,In_594);
nor U1174 (N_1174,In_861,In_308);
and U1175 (N_1175,In_1212,In_213);
and U1176 (N_1176,In_1110,In_109);
and U1177 (N_1177,In_1016,In_523);
and U1178 (N_1178,In_932,In_562);
and U1179 (N_1179,In_843,In_66);
xnor U1180 (N_1180,In_580,In_1259);
xor U1181 (N_1181,In_1292,In_1403);
or U1182 (N_1182,In_1456,In_578);
nor U1183 (N_1183,In_1013,In_1468);
or U1184 (N_1184,In_155,In_466);
xor U1185 (N_1185,In_1024,In_1357);
nand U1186 (N_1186,In_867,In_536);
or U1187 (N_1187,In_1454,In_1256);
and U1188 (N_1188,In_1428,In_579);
nand U1189 (N_1189,In_21,In_1394);
xnor U1190 (N_1190,In_631,In_718);
nor U1191 (N_1191,In_31,In_1005);
nand U1192 (N_1192,In_208,In_1071);
or U1193 (N_1193,In_779,In_934);
and U1194 (N_1194,In_1492,In_74);
nand U1195 (N_1195,In_506,In_661);
xor U1196 (N_1196,In_588,In_632);
nor U1197 (N_1197,In_943,In_1485);
nor U1198 (N_1198,In_550,In_1188);
and U1199 (N_1199,In_832,In_1247);
and U1200 (N_1200,In_565,In_1371);
or U1201 (N_1201,In_423,In_65);
xor U1202 (N_1202,In_103,In_949);
or U1203 (N_1203,In_170,In_836);
and U1204 (N_1204,In_1411,In_431);
nand U1205 (N_1205,In_1160,In_1080);
and U1206 (N_1206,In_1119,In_1132);
nor U1207 (N_1207,In_850,In_864);
or U1208 (N_1208,In_43,In_1341);
or U1209 (N_1209,In_1299,In_932);
and U1210 (N_1210,In_1146,In_354);
nor U1211 (N_1211,In_618,In_148);
or U1212 (N_1212,In_1253,In_104);
and U1213 (N_1213,In_642,In_423);
nand U1214 (N_1214,In_232,In_36);
xnor U1215 (N_1215,In_1031,In_888);
and U1216 (N_1216,In_1481,In_575);
or U1217 (N_1217,In_557,In_708);
nand U1218 (N_1218,In_768,In_518);
nand U1219 (N_1219,In_1286,In_531);
xnor U1220 (N_1220,In_200,In_983);
nand U1221 (N_1221,In_810,In_421);
and U1222 (N_1222,In_1196,In_1283);
or U1223 (N_1223,In_950,In_1296);
or U1224 (N_1224,In_1262,In_517);
and U1225 (N_1225,In_1050,In_606);
and U1226 (N_1226,In_656,In_594);
or U1227 (N_1227,In_1058,In_560);
nand U1228 (N_1228,In_337,In_555);
or U1229 (N_1229,In_1113,In_452);
and U1230 (N_1230,In_631,In_129);
nor U1231 (N_1231,In_315,In_410);
or U1232 (N_1232,In_1429,In_1312);
or U1233 (N_1233,In_337,In_1201);
and U1234 (N_1234,In_453,In_715);
nand U1235 (N_1235,In_73,In_1489);
or U1236 (N_1236,In_18,In_212);
and U1237 (N_1237,In_957,In_402);
nand U1238 (N_1238,In_1439,In_629);
nor U1239 (N_1239,In_1156,In_1397);
xor U1240 (N_1240,In_509,In_357);
and U1241 (N_1241,In_735,In_1027);
nor U1242 (N_1242,In_1424,In_1337);
xor U1243 (N_1243,In_74,In_813);
and U1244 (N_1244,In_252,In_1095);
nand U1245 (N_1245,In_661,In_1117);
nor U1246 (N_1246,In_295,In_1126);
nand U1247 (N_1247,In_884,In_433);
xor U1248 (N_1248,In_1039,In_742);
nand U1249 (N_1249,In_1455,In_937);
and U1250 (N_1250,In_1123,In_229);
nor U1251 (N_1251,In_981,In_1292);
nor U1252 (N_1252,In_297,In_671);
nor U1253 (N_1253,In_1250,In_582);
xor U1254 (N_1254,In_799,In_1207);
nand U1255 (N_1255,In_70,In_295);
and U1256 (N_1256,In_804,In_1419);
or U1257 (N_1257,In_1460,In_1494);
nor U1258 (N_1258,In_116,In_1331);
or U1259 (N_1259,In_855,In_1419);
nor U1260 (N_1260,In_292,In_430);
nor U1261 (N_1261,In_125,In_1331);
or U1262 (N_1262,In_1010,In_11);
and U1263 (N_1263,In_1007,In_1446);
and U1264 (N_1264,In_1258,In_681);
or U1265 (N_1265,In_176,In_708);
xnor U1266 (N_1266,In_1248,In_1053);
or U1267 (N_1267,In_1404,In_1162);
and U1268 (N_1268,In_1464,In_354);
or U1269 (N_1269,In_1031,In_421);
nand U1270 (N_1270,In_1202,In_1166);
or U1271 (N_1271,In_1064,In_480);
and U1272 (N_1272,In_173,In_1103);
xor U1273 (N_1273,In_211,In_1075);
nand U1274 (N_1274,In_1219,In_182);
xor U1275 (N_1275,In_212,In_712);
nand U1276 (N_1276,In_915,In_704);
or U1277 (N_1277,In_1262,In_1143);
or U1278 (N_1278,In_960,In_1201);
or U1279 (N_1279,In_17,In_442);
or U1280 (N_1280,In_771,In_1283);
and U1281 (N_1281,In_685,In_540);
nor U1282 (N_1282,In_941,In_1102);
and U1283 (N_1283,In_777,In_1061);
xnor U1284 (N_1284,In_573,In_1148);
or U1285 (N_1285,In_438,In_590);
xnor U1286 (N_1286,In_539,In_80);
nand U1287 (N_1287,In_49,In_987);
and U1288 (N_1288,In_606,In_155);
or U1289 (N_1289,In_1075,In_1383);
and U1290 (N_1290,In_626,In_851);
or U1291 (N_1291,In_888,In_295);
xnor U1292 (N_1292,In_567,In_129);
nor U1293 (N_1293,In_742,In_609);
and U1294 (N_1294,In_172,In_315);
nor U1295 (N_1295,In_1480,In_1347);
or U1296 (N_1296,In_1460,In_356);
xor U1297 (N_1297,In_1278,In_491);
nand U1298 (N_1298,In_1317,In_288);
nand U1299 (N_1299,In_1338,In_660);
and U1300 (N_1300,In_573,In_444);
or U1301 (N_1301,In_1004,In_374);
nand U1302 (N_1302,In_1036,In_740);
and U1303 (N_1303,In_256,In_677);
nor U1304 (N_1304,In_702,In_698);
nand U1305 (N_1305,In_587,In_313);
nor U1306 (N_1306,In_520,In_680);
xnor U1307 (N_1307,In_1183,In_1034);
nand U1308 (N_1308,In_20,In_1471);
nand U1309 (N_1309,In_488,In_492);
nand U1310 (N_1310,In_928,In_735);
xor U1311 (N_1311,In_1321,In_1027);
and U1312 (N_1312,In_1420,In_84);
nand U1313 (N_1313,In_314,In_252);
and U1314 (N_1314,In_1025,In_1055);
nand U1315 (N_1315,In_1005,In_931);
nand U1316 (N_1316,In_1114,In_1280);
nor U1317 (N_1317,In_1004,In_1184);
nor U1318 (N_1318,In_726,In_950);
nor U1319 (N_1319,In_162,In_958);
xnor U1320 (N_1320,In_386,In_492);
and U1321 (N_1321,In_134,In_1340);
xor U1322 (N_1322,In_595,In_286);
nand U1323 (N_1323,In_972,In_166);
nand U1324 (N_1324,In_3,In_357);
nor U1325 (N_1325,In_840,In_46);
xnor U1326 (N_1326,In_1491,In_319);
nand U1327 (N_1327,In_584,In_1339);
and U1328 (N_1328,In_836,In_448);
nand U1329 (N_1329,In_554,In_210);
xnor U1330 (N_1330,In_730,In_584);
and U1331 (N_1331,In_839,In_505);
nor U1332 (N_1332,In_142,In_826);
nand U1333 (N_1333,In_1158,In_512);
or U1334 (N_1334,In_859,In_24);
or U1335 (N_1335,In_108,In_804);
nor U1336 (N_1336,In_502,In_953);
and U1337 (N_1337,In_723,In_1117);
nor U1338 (N_1338,In_621,In_143);
or U1339 (N_1339,In_385,In_1045);
or U1340 (N_1340,In_697,In_173);
nand U1341 (N_1341,In_720,In_775);
nand U1342 (N_1342,In_67,In_735);
nor U1343 (N_1343,In_1297,In_1129);
nor U1344 (N_1344,In_781,In_1003);
and U1345 (N_1345,In_1018,In_1182);
and U1346 (N_1346,In_810,In_1051);
and U1347 (N_1347,In_586,In_853);
nand U1348 (N_1348,In_259,In_916);
nor U1349 (N_1349,In_484,In_214);
nor U1350 (N_1350,In_59,In_465);
nor U1351 (N_1351,In_65,In_370);
nor U1352 (N_1352,In_825,In_1428);
and U1353 (N_1353,In_544,In_261);
nand U1354 (N_1354,In_1393,In_1316);
nor U1355 (N_1355,In_657,In_604);
nor U1356 (N_1356,In_1298,In_731);
nand U1357 (N_1357,In_120,In_1197);
nand U1358 (N_1358,In_470,In_150);
or U1359 (N_1359,In_762,In_1427);
nand U1360 (N_1360,In_504,In_942);
or U1361 (N_1361,In_1265,In_442);
nand U1362 (N_1362,In_664,In_773);
xor U1363 (N_1363,In_206,In_667);
nor U1364 (N_1364,In_1452,In_221);
nand U1365 (N_1365,In_1165,In_190);
xor U1366 (N_1366,In_273,In_28);
xnor U1367 (N_1367,In_160,In_518);
and U1368 (N_1368,In_743,In_1124);
or U1369 (N_1369,In_465,In_748);
xor U1370 (N_1370,In_651,In_360);
nor U1371 (N_1371,In_1060,In_1468);
and U1372 (N_1372,In_1405,In_1471);
or U1373 (N_1373,In_988,In_1317);
xor U1374 (N_1374,In_58,In_211);
and U1375 (N_1375,In_858,In_848);
nor U1376 (N_1376,In_1056,In_260);
or U1377 (N_1377,In_1360,In_473);
nand U1378 (N_1378,In_1183,In_880);
nand U1379 (N_1379,In_1072,In_1490);
and U1380 (N_1380,In_245,In_1187);
xor U1381 (N_1381,In_694,In_149);
nand U1382 (N_1382,In_1350,In_1241);
nand U1383 (N_1383,In_763,In_381);
nand U1384 (N_1384,In_902,In_1375);
xor U1385 (N_1385,In_1394,In_1173);
nand U1386 (N_1386,In_251,In_486);
or U1387 (N_1387,In_1097,In_648);
and U1388 (N_1388,In_1153,In_42);
and U1389 (N_1389,In_548,In_234);
xor U1390 (N_1390,In_53,In_1244);
or U1391 (N_1391,In_339,In_1002);
or U1392 (N_1392,In_873,In_838);
nand U1393 (N_1393,In_1239,In_822);
or U1394 (N_1394,In_1459,In_1409);
nor U1395 (N_1395,In_1243,In_306);
and U1396 (N_1396,In_1475,In_361);
nand U1397 (N_1397,In_253,In_359);
nor U1398 (N_1398,In_357,In_1278);
xnor U1399 (N_1399,In_995,In_70);
nor U1400 (N_1400,In_803,In_64);
nand U1401 (N_1401,In_1171,In_212);
nor U1402 (N_1402,In_295,In_44);
nand U1403 (N_1403,In_902,In_253);
nor U1404 (N_1404,In_1297,In_980);
and U1405 (N_1405,In_1431,In_949);
xnor U1406 (N_1406,In_957,In_1458);
and U1407 (N_1407,In_805,In_71);
or U1408 (N_1408,In_310,In_1391);
xnor U1409 (N_1409,In_140,In_819);
xor U1410 (N_1410,In_709,In_1219);
nor U1411 (N_1411,In_1190,In_1271);
nand U1412 (N_1412,In_351,In_863);
xor U1413 (N_1413,In_598,In_122);
nor U1414 (N_1414,In_699,In_28);
nand U1415 (N_1415,In_928,In_1371);
and U1416 (N_1416,In_744,In_357);
nor U1417 (N_1417,In_928,In_516);
xor U1418 (N_1418,In_151,In_244);
nand U1419 (N_1419,In_742,In_141);
xnor U1420 (N_1420,In_1231,In_207);
or U1421 (N_1421,In_62,In_90);
xnor U1422 (N_1422,In_1148,In_192);
and U1423 (N_1423,In_592,In_896);
or U1424 (N_1424,In_988,In_558);
nor U1425 (N_1425,In_1454,In_430);
nor U1426 (N_1426,In_650,In_1265);
nor U1427 (N_1427,In_589,In_200);
nand U1428 (N_1428,In_998,In_848);
nand U1429 (N_1429,In_841,In_1194);
or U1430 (N_1430,In_143,In_1042);
and U1431 (N_1431,In_36,In_303);
nand U1432 (N_1432,In_846,In_1197);
and U1433 (N_1433,In_1160,In_614);
and U1434 (N_1434,In_1298,In_1099);
or U1435 (N_1435,In_874,In_449);
nor U1436 (N_1436,In_462,In_1036);
nor U1437 (N_1437,In_480,In_1191);
nor U1438 (N_1438,In_834,In_915);
xor U1439 (N_1439,In_591,In_1241);
nand U1440 (N_1440,In_877,In_1378);
xnor U1441 (N_1441,In_23,In_1035);
xnor U1442 (N_1442,In_1228,In_775);
nand U1443 (N_1443,In_795,In_831);
xnor U1444 (N_1444,In_1455,In_575);
nor U1445 (N_1445,In_1335,In_1037);
nor U1446 (N_1446,In_904,In_323);
nand U1447 (N_1447,In_1373,In_193);
nor U1448 (N_1448,In_752,In_788);
xnor U1449 (N_1449,In_507,In_191);
nor U1450 (N_1450,In_1192,In_468);
nand U1451 (N_1451,In_413,In_511);
xnor U1452 (N_1452,In_1066,In_159);
nor U1453 (N_1453,In_811,In_1025);
xor U1454 (N_1454,In_785,In_1492);
and U1455 (N_1455,In_1353,In_293);
nand U1456 (N_1456,In_1260,In_1261);
or U1457 (N_1457,In_784,In_271);
nor U1458 (N_1458,In_1107,In_346);
and U1459 (N_1459,In_98,In_38);
or U1460 (N_1460,In_1196,In_967);
nand U1461 (N_1461,In_667,In_224);
nor U1462 (N_1462,In_901,In_457);
and U1463 (N_1463,In_471,In_1214);
nand U1464 (N_1464,In_441,In_538);
or U1465 (N_1465,In_939,In_652);
or U1466 (N_1466,In_112,In_354);
nand U1467 (N_1467,In_13,In_1244);
or U1468 (N_1468,In_626,In_675);
nor U1469 (N_1469,In_188,In_1155);
nor U1470 (N_1470,In_1031,In_1082);
nor U1471 (N_1471,In_748,In_419);
or U1472 (N_1472,In_891,In_1225);
and U1473 (N_1473,In_1105,In_918);
or U1474 (N_1474,In_1400,In_373);
nand U1475 (N_1475,In_168,In_638);
and U1476 (N_1476,In_1426,In_90);
and U1477 (N_1477,In_25,In_43);
nand U1478 (N_1478,In_974,In_635);
and U1479 (N_1479,In_697,In_821);
and U1480 (N_1480,In_122,In_1429);
and U1481 (N_1481,In_357,In_423);
xnor U1482 (N_1482,In_895,In_258);
and U1483 (N_1483,In_722,In_792);
nor U1484 (N_1484,In_462,In_350);
and U1485 (N_1485,In_246,In_36);
xor U1486 (N_1486,In_1101,In_222);
nor U1487 (N_1487,In_1012,In_1487);
nand U1488 (N_1488,In_1289,In_666);
and U1489 (N_1489,In_940,In_499);
nand U1490 (N_1490,In_1042,In_111);
nand U1491 (N_1491,In_353,In_928);
and U1492 (N_1492,In_1066,In_1037);
nand U1493 (N_1493,In_341,In_72);
and U1494 (N_1494,In_1033,In_183);
and U1495 (N_1495,In_43,In_1465);
and U1496 (N_1496,In_990,In_659);
xor U1497 (N_1497,In_871,In_1360);
nand U1498 (N_1498,In_1112,In_557);
xor U1499 (N_1499,In_779,In_1469);
or U1500 (N_1500,In_361,In_1466);
nor U1501 (N_1501,In_676,In_638);
or U1502 (N_1502,In_1190,In_587);
or U1503 (N_1503,In_960,In_900);
xnor U1504 (N_1504,In_1271,In_748);
nand U1505 (N_1505,In_11,In_1235);
nor U1506 (N_1506,In_518,In_1294);
nor U1507 (N_1507,In_131,In_477);
nand U1508 (N_1508,In_1386,In_967);
nand U1509 (N_1509,In_1432,In_739);
and U1510 (N_1510,In_1423,In_1271);
nand U1511 (N_1511,In_1380,In_994);
xor U1512 (N_1512,In_679,In_291);
or U1513 (N_1513,In_1476,In_164);
nor U1514 (N_1514,In_69,In_722);
nand U1515 (N_1515,In_193,In_1315);
and U1516 (N_1516,In_1322,In_282);
xnor U1517 (N_1517,In_803,In_1473);
nor U1518 (N_1518,In_521,In_386);
xor U1519 (N_1519,In_931,In_1446);
nor U1520 (N_1520,In_857,In_53);
nand U1521 (N_1521,In_973,In_1136);
nor U1522 (N_1522,In_346,In_43);
nand U1523 (N_1523,In_817,In_371);
xor U1524 (N_1524,In_724,In_344);
nor U1525 (N_1525,In_1160,In_374);
nand U1526 (N_1526,In_1363,In_255);
nand U1527 (N_1527,In_461,In_706);
and U1528 (N_1528,In_557,In_374);
xor U1529 (N_1529,In_1150,In_1322);
or U1530 (N_1530,In_639,In_620);
nor U1531 (N_1531,In_1401,In_839);
nand U1532 (N_1532,In_1470,In_1262);
and U1533 (N_1533,In_407,In_341);
xor U1534 (N_1534,In_966,In_813);
or U1535 (N_1535,In_472,In_635);
nand U1536 (N_1536,In_860,In_52);
or U1537 (N_1537,In_1071,In_405);
or U1538 (N_1538,In_82,In_414);
nand U1539 (N_1539,In_1128,In_939);
xnor U1540 (N_1540,In_103,In_272);
and U1541 (N_1541,In_1235,In_422);
or U1542 (N_1542,In_578,In_840);
xnor U1543 (N_1543,In_1311,In_842);
or U1544 (N_1544,In_1187,In_444);
xor U1545 (N_1545,In_92,In_1023);
or U1546 (N_1546,In_1425,In_132);
or U1547 (N_1547,In_432,In_555);
nor U1548 (N_1548,In_201,In_411);
or U1549 (N_1549,In_4,In_1362);
nor U1550 (N_1550,In_471,In_649);
or U1551 (N_1551,In_1171,In_1346);
xor U1552 (N_1552,In_973,In_1176);
nand U1553 (N_1553,In_1489,In_323);
and U1554 (N_1554,In_1329,In_1067);
xor U1555 (N_1555,In_181,In_72);
nand U1556 (N_1556,In_493,In_86);
or U1557 (N_1557,In_147,In_1158);
xor U1558 (N_1558,In_934,In_29);
nand U1559 (N_1559,In_434,In_927);
or U1560 (N_1560,In_163,In_1338);
nor U1561 (N_1561,In_698,In_1495);
nor U1562 (N_1562,In_858,In_753);
and U1563 (N_1563,In_1247,In_669);
nand U1564 (N_1564,In_188,In_286);
nor U1565 (N_1565,In_410,In_725);
nor U1566 (N_1566,In_715,In_1202);
or U1567 (N_1567,In_450,In_134);
or U1568 (N_1568,In_520,In_468);
nor U1569 (N_1569,In_1260,In_1021);
nor U1570 (N_1570,In_204,In_213);
or U1571 (N_1571,In_501,In_331);
nand U1572 (N_1572,In_1160,In_1457);
nor U1573 (N_1573,In_1397,In_53);
or U1574 (N_1574,In_1158,In_1304);
and U1575 (N_1575,In_629,In_814);
xor U1576 (N_1576,In_448,In_153);
and U1577 (N_1577,In_142,In_802);
or U1578 (N_1578,In_1174,In_1031);
or U1579 (N_1579,In_315,In_339);
nand U1580 (N_1580,In_1178,In_947);
xnor U1581 (N_1581,In_351,In_483);
xor U1582 (N_1582,In_140,In_962);
and U1583 (N_1583,In_780,In_1010);
nand U1584 (N_1584,In_1072,In_417);
or U1585 (N_1585,In_424,In_843);
nand U1586 (N_1586,In_373,In_1175);
nor U1587 (N_1587,In_1088,In_747);
or U1588 (N_1588,In_153,In_839);
xnor U1589 (N_1589,In_473,In_803);
and U1590 (N_1590,In_461,In_597);
nand U1591 (N_1591,In_235,In_599);
or U1592 (N_1592,In_446,In_1259);
nand U1593 (N_1593,In_544,In_308);
xor U1594 (N_1594,In_1311,In_824);
or U1595 (N_1595,In_698,In_231);
and U1596 (N_1596,In_757,In_1484);
xnor U1597 (N_1597,In_28,In_931);
nor U1598 (N_1598,In_30,In_35);
or U1599 (N_1599,In_837,In_597);
and U1600 (N_1600,In_828,In_137);
nor U1601 (N_1601,In_1438,In_1148);
nor U1602 (N_1602,In_216,In_701);
nand U1603 (N_1603,In_211,In_1208);
nand U1604 (N_1604,In_1308,In_1026);
nand U1605 (N_1605,In_888,In_1050);
nor U1606 (N_1606,In_920,In_1154);
and U1607 (N_1607,In_547,In_596);
nand U1608 (N_1608,In_121,In_704);
and U1609 (N_1609,In_739,In_8);
nand U1610 (N_1610,In_1123,In_984);
nand U1611 (N_1611,In_1289,In_672);
nand U1612 (N_1612,In_83,In_1346);
or U1613 (N_1613,In_909,In_1301);
nor U1614 (N_1614,In_41,In_1269);
nand U1615 (N_1615,In_1340,In_573);
or U1616 (N_1616,In_333,In_178);
nor U1617 (N_1617,In_94,In_708);
or U1618 (N_1618,In_1006,In_3);
and U1619 (N_1619,In_287,In_940);
xor U1620 (N_1620,In_799,In_731);
and U1621 (N_1621,In_1239,In_113);
nor U1622 (N_1622,In_289,In_1459);
xnor U1623 (N_1623,In_1060,In_337);
or U1624 (N_1624,In_1346,In_195);
nand U1625 (N_1625,In_520,In_875);
xor U1626 (N_1626,In_187,In_257);
xnor U1627 (N_1627,In_1384,In_323);
and U1628 (N_1628,In_228,In_1499);
nand U1629 (N_1629,In_1477,In_754);
and U1630 (N_1630,In_845,In_193);
or U1631 (N_1631,In_1179,In_1265);
nor U1632 (N_1632,In_1219,In_931);
nor U1633 (N_1633,In_1488,In_1365);
or U1634 (N_1634,In_731,In_730);
nand U1635 (N_1635,In_1331,In_489);
and U1636 (N_1636,In_613,In_791);
nor U1637 (N_1637,In_1408,In_1410);
and U1638 (N_1638,In_545,In_988);
and U1639 (N_1639,In_608,In_958);
and U1640 (N_1640,In_51,In_1280);
nand U1641 (N_1641,In_1497,In_1203);
nor U1642 (N_1642,In_703,In_303);
nand U1643 (N_1643,In_269,In_1296);
xor U1644 (N_1644,In_79,In_338);
or U1645 (N_1645,In_1434,In_1287);
or U1646 (N_1646,In_463,In_648);
nand U1647 (N_1647,In_784,In_172);
or U1648 (N_1648,In_1180,In_761);
nand U1649 (N_1649,In_735,In_739);
nand U1650 (N_1650,In_978,In_456);
nor U1651 (N_1651,In_1490,In_113);
xnor U1652 (N_1652,In_1439,In_593);
nand U1653 (N_1653,In_78,In_175);
and U1654 (N_1654,In_955,In_448);
nor U1655 (N_1655,In_975,In_1075);
nand U1656 (N_1656,In_885,In_175);
or U1657 (N_1657,In_955,In_661);
and U1658 (N_1658,In_155,In_487);
and U1659 (N_1659,In_916,In_519);
and U1660 (N_1660,In_818,In_1011);
nand U1661 (N_1661,In_649,In_778);
and U1662 (N_1662,In_64,In_414);
or U1663 (N_1663,In_1320,In_936);
or U1664 (N_1664,In_223,In_1365);
nand U1665 (N_1665,In_1267,In_541);
or U1666 (N_1666,In_698,In_41);
and U1667 (N_1667,In_1141,In_629);
or U1668 (N_1668,In_459,In_585);
and U1669 (N_1669,In_171,In_168);
nand U1670 (N_1670,In_281,In_808);
xor U1671 (N_1671,In_1001,In_1110);
xor U1672 (N_1672,In_188,In_342);
nor U1673 (N_1673,In_117,In_592);
and U1674 (N_1674,In_1077,In_252);
nor U1675 (N_1675,In_845,In_1009);
xor U1676 (N_1676,In_787,In_40);
or U1677 (N_1677,In_92,In_840);
or U1678 (N_1678,In_388,In_1496);
xor U1679 (N_1679,In_130,In_266);
and U1680 (N_1680,In_952,In_281);
and U1681 (N_1681,In_1262,In_1290);
or U1682 (N_1682,In_1178,In_945);
nor U1683 (N_1683,In_1327,In_1224);
or U1684 (N_1684,In_268,In_841);
and U1685 (N_1685,In_1219,In_1442);
or U1686 (N_1686,In_584,In_439);
and U1687 (N_1687,In_745,In_786);
nor U1688 (N_1688,In_1426,In_937);
or U1689 (N_1689,In_1389,In_264);
and U1690 (N_1690,In_1214,In_78);
xnor U1691 (N_1691,In_819,In_454);
and U1692 (N_1692,In_431,In_143);
or U1693 (N_1693,In_255,In_36);
or U1694 (N_1694,In_1481,In_115);
and U1695 (N_1695,In_391,In_461);
or U1696 (N_1696,In_44,In_337);
nand U1697 (N_1697,In_1290,In_600);
and U1698 (N_1698,In_1128,In_95);
nand U1699 (N_1699,In_269,In_1155);
nor U1700 (N_1700,In_297,In_1391);
or U1701 (N_1701,In_694,In_969);
xnor U1702 (N_1702,In_944,In_584);
nor U1703 (N_1703,In_1386,In_282);
or U1704 (N_1704,In_229,In_513);
or U1705 (N_1705,In_1446,In_971);
and U1706 (N_1706,In_235,In_1327);
nor U1707 (N_1707,In_672,In_323);
or U1708 (N_1708,In_67,In_1460);
and U1709 (N_1709,In_834,In_1146);
xor U1710 (N_1710,In_359,In_364);
and U1711 (N_1711,In_863,In_476);
or U1712 (N_1712,In_874,In_111);
and U1713 (N_1713,In_1075,In_552);
xor U1714 (N_1714,In_1447,In_1369);
nor U1715 (N_1715,In_555,In_1184);
and U1716 (N_1716,In_828,In_1172);
and U1717 (N_1717,In_1293,In_230);
nor U1718 (N_1718,In_671,In_428);
xnor U1719 (N_1719,In_814,In_720);
nand U1720 (N_1720,In_1285,In_154);
nand U1721 (N_1721,In_1023,In_1031);
or U1722 (N_1722,In_404,In_1244);
nor U1723 (N_1723,In_1487,In_412);
or U1724 (N_1724,In_393,In_252);
and U1725 (N_1725,In_1189,In_382);
nor U1726 (N_1726,In_243,In_1309);
or U1727 (N_1727,In_190,In_1136);
and U1728 (N_1728,In_345,In_271);
xor U1729 (N_1729,In_1146,In_225);
nor U1730 (N_1730,In_493,In_1323);
and U1731 (N_1731,In_483,In_1350);
and U1732 (N_1732,In_434,In_992);
xor U1733 (N_1733,In_1377,In_802);
and U1734 (N_1734,In_144,In_632);
nor U1735 (N_1735,In_926,In_786);
nand U1736 (N_1736,In_1370,In_635);
and U1737 (N_1737,In_1361,In_1011);
nor U1738 (N_1738,In_1055,In_666);
and U1739 (N_1739,In_446,In_695);
nor U1740 (N_1740,In_1102,In_1188);
xnor U1741 (N_1741,In_115,In_1280);
xor U1742 (N_1742,In_229,In_531);
or U1743 (N_1743,In_759,In_47);
xor U1744 (N_1744,In_1394,In_12);
nand U1745 (N_1745,In_954,In_1245);
and U1746 (N_1746,In_634,In_38);
nor U1747 (N_1747,In_28,In_31);
xnor U1748 (N_1748,In_818,In_1465);
or U1749 (N_1749,In_54,In_1176);
nor U1750 (N_1750,In_166,In_1137);
nor U1751 (N_1751,In_1096,In_1233);
nand U1752 (N_1752,In_872,In_349);
nand U1753 (N_1753,In_28,In_831);
or U1754 (N_1754,In_842,In_362);
and U1755 (N_1755,In_21,In_352);
and U1756 (N_1756,In_1074,In_1038);
xor U1757 (N_1757,In_103,In_1104);
nand U1758 (N_1758,In_1282,In_625);
nand U1759 (N_1759,In_1089,In_1334);
nor U1760 (N_1760,In_1244,In_623);
nand U1761 (N_1761,In_821,In_224);
xor U1762 (N_1762,In_414,In_90);
nor U1763 (N_1763,In_255,In_1200);
or U1764 (N_1764,In_1153,In_1172);
nand U1765 (N_1765,In_234,In_1439);
or U1766 (N_1766,In_1015,In_154);
nor U1767 (N_1767,In_1261,In_1216);
nand U1768 (N_1768,In_1312,In_671);
nor U1769 (N_1769,In_34,In_205);
and U1770 (N_1770,In_45,In_43);
or U1771 (N_1771,In_1491,In_240);
or U1772 (N_1772,In_792,In_1385);
or U1773 (N_1773,In_964,In_1131);
and U1774 (N_1774,In_1133,In_610);
nor U1775 (N_1775,In_1259,In_388);
and U1776 (N_1776,In_1241,In_652);
xnor U1777 (N_1777,In_428,In_113);
or U1778 (N_1778,In_1079,In_1391);
and U1779 (N_1779,In_1417,In_1174);
nor U1780 (N_1780,In_1024,In_849);
xnor U1781 (N_1781,In_275,In_1438);
xnor U1782 (N_1782,In_667,In_1092);
nor U1783 (N_1783,In_906,In_673);
nand U1784 (N_1784,In_1143,In_1482);
and U1785 (N_1785,In_1299,In_684);
nor U1786 (N_1786,In_1334,In_561);
xnor U1787 (N_1787,In_1329,In_1405);
and U1788 (N_1788,In_710,In_44);
or U1789 (N_1789,In_941,In_1383);
and U1790 (N_1790,In_586,In_263);
xor U1791 (N_1791,In_856,In_7);
xor U1792 (N_1792,In_328,In_1224);
or U1793 (N_1793,In_68,In_1364);
xor U1794 (N_1794,In_1113,In_820);
or U1795 (N_1795,In_104,In_959);
or U1796 (N_1796,In_58,In_700);
xor U1797 (N_1797,In_945,In_54);
xnor U1798 (N_1798,In_1351,In_75);
or U1799 (N_1799,In_1165,In_1050);
and U1800 (N_1800,In_392,In_1113);
nand U1801 (N_1801,In_455,In_1055);
nand U1802 (N_1802,In_660,In_594);
xor U1803 (N_1803,In_1402,In_884);
nand U1804 (N_1804,In_841,In_72);
nand U1805 (N_1805,In_444,In_421);
nor U1806 (N_1806,In_559,In_982);
or U1807 (N_1807,In_321,In_301);
and U1808 (N_1808,In_1269,In_167);
xnor U1809 (N_1809,In_148,In_43);
and U1810 (N_1810,In_755,In_955);
xnor U1811 (N_1811,In_940,In_1174);
nor U1812 (N_1812,In_138,In_1266);
xor U1813 (N_1813,In_443,In_343);
or U1814 (N_1814,In_1249,In_912);
nor U1815 (N_1815,In_340,In_1072);
xnor U1816 (N_1816,In_954,In_1378);
and U1817 (N_1817,In_375,In_1114);
or U1818 (N_1818,In_1003,In_1089);
xnor U1819 (N_1819,In_201,In_277);
and U1820 (N_1820,In_216,In_647);
nand U1821 (N_1821,In_1219,In_1418);
nand U1822 (N_1822,In_199,In_145);
nor U1823 (N_1823,In_792,In_978);
nand U1824 (N_1824,In_885,In_956);
and U1825 (N_1825,In_1459,In_109);
nor U1826 (N_1826,In_1054,In_1483);
nand U1827 (N_1827,In_90,In_707);
nor U1828 (N_1828,In_1371,In_1086);
nand U1829 (N_1829,In_1144,In_385);
and U1830 (N_1830,In_703,In_1344);
xnor U1831 (N_1831,In_1222,In_458);
nand U1832 (N_1832,In_280,In_1349);
and U1833 (N_1833,In_1016,In_271);
and U1834 (N_1834,In_1345,In_945);
nand U1835 (N_1835,In_1268,In_1224);
nor U1836 (N_1836,In_930,In_203);
and U1837 (N_1837,In_1098,In_711);
or U1838 (N_1838,In_697,In_392);
xnor U1839 (N_1839,In_1230,In_1070);
and U1840 (N_1840,In_983,In_1343);
and U1841 (N_1841,In_862,In_1192);
xor U1842 (N_1842,In_1091,In_578);
and U1843 (N_1843,In_54,In_791);
nor U1844 (N_1844,In_860,In_245);
xnor U1845 (N_1845,In_598,In_212);
or U1846 (N_1846,In_693,In_622);
xnor U1847 (N_1847,In_1175,In_50);
xor U1848 (N_1848,In_816,In_944);
nor U1849 (N_1849,In_355,In_345);
nor U1850 (N_1850,In_1362,In_1236);
nand U1851 (N_1851,In_139,In_695);
nor U1852 (N_1852,In_1427,In_178);
nor U1853 (N_1853,In_404,In_698);
and U1854 (N_1854,In_960,In_896);
or U1855 (N_1855,In_1448,In_1062);
nor U1856 (N_1856,In_1338,In_1387);
xnor U1857 (N_1857,In_916,In_951);
nor U1858 (N_1858,In_970,In_162);
or U1859 (N_1859,In_842,In_13);
or U1860 (N_1860,In_960,In_1489);
and U1861 (N_1861,In_1485,In_275);
xor U1862 (N_1862,In_413,In_10);
and U1863 (N_1863,In_491,In_928);
nor U1864 (N_1864,In_144,In_15);
or U1865 (N_1865,In_765,In_1309);
or U1866 (N_1866,In_1012,In_1133);
and U1867 (N_1867,In_474,In_445);
nor U1868 (N_1868,In_853,In_870);
or U1869 (N_1869,In_1329,In_201);
nor U1870 (N_1870,In_833,In_592);
xor U1871 (N_1871,In_1224,In_7);
nand U1872 (N_1872,In_686,In_380);
nor U1873 (N_1873,In_268,In_956);
nor U1874 (N_1874,In_705,In_40);
or U1875 (N_1875,In_1257,In_1481);
xor U1876 (N_1876,In_1481,In_1492);
nand U1877 (N_1877,In_691,In_1141);
xnor U1878 (N_1878,In_449,In_1376);
nor U1879 (N_1879,In_1236,In_1127);
nor U1880 (N_1880,In_1496,In_73);
xnor U1881 (N_1881,In_1475,In_238);
nor U1882 (N_1882,In_959,In_91);
xor U1883 (N_1883,In_518,In_579);
or U1884 (N_1884,In_988,In_641);
nand U1885 (N_1885,In_1437,In_374);
or U1886 (N_1886,In_1042,In_501);
xor U1887 (N_1887,In_735,In_610);
or U1888 (N_1888,In_569,In_599);
or U1889 (N_1889,In_929,In_1199);
nor U1890 (N_1890,In_960,In_1350);
xor U1891 (N_1891,In_1123,In_1462);
nand U1892 (N_1892,In_166,In_1077);
and U1893 (N_1893,In_1453,In_595);
nand U1894 (N_1894,In_596,In_371);
nand U1895 (N_1895,In_437,In_1413);
or U1896 (N_1896,In_781,In_997);
and U1897 (N_1897,In_836,In_1182);
and U1898 (N_1898,In_750,In_741);
xnor U1899 (N_1899,In_1160,In_929);
xor U1900 (N_1900,In_144,In_530);
or U1901 (N_1901,In_439,In_300);
nand U1902 (N_1902,In_364,In_350);
xor U1903 (N_1903,In_1019,In_548);
xnor U1904 (N_1904,In_352,In_24);
or U1905 (N_1905,In_171,In_210);
xor U1906 (N_1906,In_1208,In_325);
or U1907 (N_1907,In_96,In_1037);
and U1908 (N_1908,In_1344,In_396);
nand U1909 (N_1909,In_146,In_1254);
nand U1910 (N_1910,In_1238,In_1324);
or U1911 (N_1911,In_1270,In_47);
and U1912 (N_1912,In_25,In_1014);
xor U1913 (N_1913,In_247,In_172);
nand U1914 (N_1914,In_683,In_329);
nand U1915 (N_1915,In_178,In_753);
or U1916 (N_1916,In_18,In_140);
nor U1917 (N_1917,In_148,In_374);
and U1918 (N_1918,In_808,In_382);
xor U1919 (N_1919,In_1075,In_671);
nor U1920 (N_1920,In_500,In_895);
nor U1921 (N_1921,In_1455,In_722);
and U1922 (N_1922,In_1451,In_1477);
and U1923 (N_1923,In_376,In_1201);
or U1924 (N_1924,In_184,In_1112);
and U1925 (N_1925,In_868,In_839);
xnor U1926 (N_1926,In_520,In_225);
or U1927 (N_1927,In_906,In_612);
nor U1928 (N_1928,In_145,In_511);
and U1929 (N_1929,In_1369,In_1);
nand U1930 (N_1930,In_1024,In_1351);
xnor U1931 (N_1931,In_795,In_1357);
or U1932 (N_1932,In_537,In_1350);
or U1933 (N_1933,In_461,In_846);
or U1934 (N_1934,In_96,In_1175);
xor U1935 (N_1935,In_304,In_1363);
xnor U1936 (N_1936,In_221,In_487);
nand U1937 (N_1937,In_377,In_1190);
nand U1938 (N_1938,In_722,In_100);
or U1939 (N_1939,In_1144,In_1025);
nand U1940 (N_1940,In_835,In_1308);
or U1941 (N_1941,In_1211,In_490);
and U1942 (N_1942,In_1153,In_819);
and U1943 (N_1943,In_272,In_245);
nor U1944 (N_1944,In_870,In_1031);
nor U1945 (N_1945,In_922,In_204);
nand U1946 (N_1946,In_1441,In_1185);
or U1947 (N_1947,In_1117,In_651);
and U1948 (N_1948,In_1012,In_821);
nor U1949 (N_1949,In_1386,In_900);
xnor U1950 (N_1950,In_994,In_976);
or U1951 (N_1951,In_1101,In_1310);
and U1952 (N_1952,In_1403,In_296);
and U1953 (N_1953,In_1198,In_1144);
and U1954 (N_1954,In_1122,In_865);
or U1955 (N_1955,In_1313,In_1301);
and U1956 (N_1956,In_1361,In_175);
xor U1957 (N_1957,In_825,In_427);
nand U1958 (N_1958,In_1479,In_1417);
nor U1959 (N_1959,In_1141,In_1317);
nor U1960 (N_1960,In_297,In_1458);
or U1961 (N_1961,In_360,In_1152);
xor U1962 (N_1962,In_445,In_613);
and U1963 (N_1963,In_318,In_323);
or U1964 (N_1964,In_1197,In_939);
and U1965 (N_1965,In_752,In_735);
or U1966 (N_1966,In_1284,In_520);
nor U1967 (N_1967,In_433,In_748);
nor U1968 (N_1968,In_1397,In_672);
nand U1969 (N_1969,In_66,In_1330);
nand U1970 (N_1970,In_296,In_844);
xnor U1971 (N_1971,In_232,In_1485);
nand U1972 (N_1972,In_1267,In_954);
nor U1973 (N_1973,In_1051,In_711);
or U1974 (N_1974,In_236,In_943);
or U1975 (N_1975,In_138,In_641);
xnor U1976 (N_1976,In_1420,In_629);
or U1977 (N_1977,In_1475,In_356);
xnor U1978 (N_1978,In_1297,In_1368);
or U1979 (N_1979,In_565,In_1185);
nand U1980 (N_1980,In_223,In_1338);
nand U1981 (N_1981,In_272,In_1278);
or U1982 (N_1982,In_144,In_209);
xor U1983 (N_1983,In_157,In_591);
xor U1984 (N_1984,In_343,In_185);
xnor U1985 (N_1985,In_64,In_192);
nand U1986 (N_1986,In_670,In_656);
nor U1987 (N_1987,In_1471,In_1478);
nand U1988 (N_1988,In_225,In_375);
nor U1989 (N_1989,In_479,In_677);
nor U1990 (N_1990,In_1169,In_1228);
nand U1991 (N_1991,In_233,In_618);
or U1992 (N_1992,In_734,In_926);
and U1993 (N_1993,In_385,In_770);
and U1994 (N_1994,In_1252,In_255);
and U1995 (N_1995,In_1457,In_227);
xnor U1996 (N_1996,In_158,In_1205);
nor U1997 (N_1997,In_193,In_1155);
or U1998 (N_1998,In_604,In_1341);
or U1999 (N_1999,In_1153,In_945);
and U2000 (N_2000,In_995,In_629);
nand U2001 (N_2001,In_142,In_1058);
nor U2002 (N_2002,In_1139,In_1064);
xor U2003 (N_2003,In_877,In_858);
xnor U2004 (N_2004,In_687,In_1360);
xor U2005 (N_2005,In_1245,In_274);
nand U2006 (N_2006,In_1058,In_405);
or U2007 (N_2007,In_400,In_170);
or U2008 (N_2008,In_298,In_1183);
and U2009 (N_2009,In_812,In_110);
nor U2010 (N_2010,In_734,In_1363);
and U2011 (N_2011,In_771,In_284);
nand U2012 (N_2012,In_726,In_1434);
xor U2013 (N_2013,In_1252,In_55);
or U2014 (N_2014,In_767,In_567);
nand U2015 (N_2015,In_247,In_179);
xnor U2016 (N_2016,In_27,In_272);
and U2017 (N_2017,In_1138,In_996);
and U2018 (N_2018,In_58,In_105);
and U2019 (N_2019,In_1392,In_814);
and U2020 (N_2020,In_1208,In_437);
xor U2021 (N_2021,In_1212,In_1042);
or U2022 (N_2022,In_316,In_1358);
nor U2023 (N_2023,In_944,In_1438);
nand U2024 (N_2024,In_916,In_440);
or U2025 (N_2025,In_1131,In_312);
nand U2026 (N_2026,In_1025,In_315);
nand U2027 (N_2027,In_491,In_955);
and U2028 (N_2028,In_204,In_602);
nand U2029 (N_2029,In_589,In_1022);
or U2030 (N_2030,In_1396,In_1442);
and U2031 (N_2031,In_309,In_695);
nand U2032 (N_2032,In_590,In_1318);
and U2033 (N_2033,In_294,In_715);
or U2034 (N_2034,In_1095,In_296);
nand U2035 (N_2035,In_570,In_427);
xnor U2036 (N_2036,In_1117,In_140);
nand U2037 (N_2037,In_626,In_928);
xnor U2038 (N_2038,In_670,In_1186);
xor U2039 (N_2039,In_1310,In_1085);
xnor U2040 (N_2040,In_767,In_615);
and U2041 (N_2041,In_624,In_642);
nor U2042 (N_2042,In_1324,In_334);
and U2043 (N_2043,In_1386,In_276);
and U2044 (N_2044,In_1268,In_895);
or U2045 (N_2045,In_109,In_246);
and U2046 (N_2046,In_866,In_339);
or U2047 (N_2047,In_532,In_306);
xor U2048 (N_2048,In_881,In_563);
or U2049 (N_2049,In_888,In_1447);
and U2050 (N_2050,In_903,In_586);
or U2051 (N_2051,In_730,In_463);
or U2052 (N_2052,In_158,In_1102);
and U2053 (N_2053,In_1453,In_1142);
xor U2054 (N_2054,In_1262,In_1169);
xor U2055 (N_2055,In_1189,In_750);
nor U2056 (N_2056,In_769,In_1335);
or U2057 (N_2057,In_963,In_138);
or U2058 (N_2058,In_703,In_869);
xor U2059 (N_2059,In_77,In_503);
or U2060 (N_2060,In_1045,In_352);
xnor U2061 (N_2061,In_979,In_1411);
or U2062 (N_2062,In_1170,In_616);
nor U2063 (N_2063,In_191,In_884);
nand U2064 (N_2064,In_533,In_342);
xor U2065 (N_2065,In_1254,In_303);
or U2066 (N_2066,In_176,In_543);
nand U2067 (N_2067,In_391,In_714);
nor U2068 (N_2068,In_776,In_767);
or U2069 (N_2069,In_425,In_293);
or U2070 (N_2070,In_342,In_571);
and U2071 (N_2071,In_1092,In_75);
nor U2072 (N_2072,In_421,In_1288);
xnor U2073 (N_2073,In_316,In_599);
xor U2074 (N_2074,In_714,In_95);
nor U2075 (N_2075,In_1462,In_118);
xor U2076 (N_2076,In_838,In_694);
xor U2077 (N_2077,In_150,In_4);
and U2078 (N_2078,In_1149,In_858);
or U2079 (N_2079,In_194,In_324);
and U2080 (N_2080,In_805,In_949);
xor U2081 (N_2081,In_779,In_800);
nand U2082 (N_2082,In_932,In_530);
and U2083 (N_2083,In_151,In_1031);
xor U2084 (N_2084,In_620,In_467);
and U2085 (N_2085,In_640,In_946);
xor U2086 (N_2086,In_1473,In_769);
xnor U2087 (N_2087,In_871,In_251);
xor U2088 (N_2088,In_306,In_334);
nand U2089 (N_2089,In_1030,In_1308);
nor U2090 (N_2090,In_716,In_504);
nand U2091 (N_2091,In_1106,In_1345);
xor U2092 (N_2092,In_281,In_1093);
nand U2093 (N_2093,In_741,In_1034);
nand U2094 (N_2094,In_439,In_158);
xor U2095 (N_2095,In_76,In_172);
nand U2096 (N_2096,In_1177,In_300);
nor U2097 (N_2097,In_1038,In_140);
nor U2098 (N_2098,In_935,In_457);
nand U2099 (N_2099,In_1152,In_293);
nand U2100 (N_2100,In_729,In_899);
xnor U2101 (N_2101,In_132,In_223);
nor U2102 (N_2102,In_393,In_563);
nor U2103 (N_2103,In_1392,In_34);
nor U2104 (N_2104,In_1244,In_670);
xor U2105 (N_2105,In_1164,In_271);
and U2106 (N_2106,In_690,In_362);
nand U2107 (N_2107,In_651,In_318);
or U2108 (N_2108,In_498,In_1431);
or U2109 (N_2109,In_4,In_938);
and U2110 (N_2110,In_948,In_1420);
or U2111 (N_2111,In_773,In_930);
xor U2112 (N_2112,In_1340,In_448);
nor U2113 (N_2113,In_99,In_1456);
nand U2114 (N_2114,In_652,In_1184);
nor U2115 (N_2115,In_725,In_1265);
nand U2116 (N_2116,In_327,In_98);
nor U2117 (N_2117,In_273,In_112);
nor U2118 (N_2118,In_1053,In_593);
or U2119 (N_2119,In_488,In_833);
xor U2120 (N_2120,In_590,In_413);
xnor U2121 (N_2121,In_1137,In_1321);
nor U2122 (N_2122,In_1459,In_893);
or U2123 (N_2123,In_94,In_328);
nor U2124 (N_2124,In_495,In_746);
and U2125 (N_2125,In_495,In_1372);
nand U2126 (N_2126,In_192,In_830);
xor U2127 (N_2127,In_989,In_380);
xor U2128 (N_2128,In_484,In_1161);
or U2129 (N_2129,In_173,In_1081);
nor U2130 (N_2130,In_437,In_1044);
and U2131 (N_2131,In_29,In_1375);
and U2132 (N_2132,In_887,In_283);
xor U2133 (N_2133,In_1392,In_248);
and U2134 (N_2134,In_1277,In_1187);
nor U2135 (N_2135,In_1241,In_1202);
xor U2136 (N_2136,In_965,In_925);
and U2137 (N_2137,In_1378,In_40);
and U2138 (N_2138,In_1077,In_819);
xor U2139 (N_2139,In_474,In_96);
nand U2140 (N_2140,In_977,In_1064);
or U2141 (N_2141,In_666,In_742);
or U2142 (N_2142,In_998,In_114);
and U2143 (N_2143,In_943,In_535);
or U2144 (N_2144,In_746,In_836);
nor U2145 (N_2145,In_960,In_74);
nor U2146 (N_2146,In_772,In_82);
and U2147 (N_2147,In_76,In_430);
or U2148 (N_2148,In_162,In_332);
xnor U2149 (N_2149,In_727,In_1062);
xor U2150 (N_2150,In_509,In_104);
or U2151 (N_2151,In_1117,In_958);
nand U2152 (N_2152,In_135,In_264);
xor U2153 (N_2153,In_1193,In_904);
nor U2154 (N_2154,In_221,In_176);
nand U2155 (N_2155,In_801,In_788);
nand U2156 (N_2156,In_1352,In_462);
xnor U2157 (N_2157,In_722,In_589);
nor U2158 (N_2158,In_472,In_1476);
or U2159 (N_2159,In_216,In_1251);
or U2160 (N_2160,In_962,In_1156);
and U2161 (N_2161,In_1325,In_1125);
or U2162 (N_2162,In_730,In_842);
xor U2163 (N_2163,In_1466,In_1021);
nand U2164 (N_2164,In_124,In_723);
nand U2165 (N_2165,In_776,In_842);
nor U2166 (N_2166,In_524,In_948);
nand U2167 (N_2167,In_64,In_524);
xnor U2168 (N_2168,In_320,In_1270);
nand U2169 (N_2169,In_848,In_1195);
or U2170 (N_2170,In_896,In_679);
nand U2171 (N_2171,In_147,In_1475);
and U2172 (N_2172,In_889,In_546);
or U2173 (N_2173,In_810,In_781);
or U2174 (N_2174,In_1449,In_885);
xor U2175 (N_2175,In_560,In_119);
or U2176 (N_2176,In_589,In_1378);
nand U2177 (N_2177,In_1144,In_671);
nor U2178 (N_2178,In_1348,In_230);
nor U2179 (N_2179,In_801,In_140);
nand U2180 (N_2180,In_1018,In_439);
and U2181 (N_2181,In_1428,In_189);
nand U2182 (N_2182,In_891,In_1013);
or U2183 (N_2183,In_916,In_1237);
nand U2184 (N_2184,In_63,In_151);
nand U2185 (N_2185,In_1043,In_910);
or U2186 (N_2186,In_337,In_798);
and U2187 (N_2187,In_1021,In_1153);
and U2188 (N_2188,In_159,In_1169);
nand U2189 (N_2189,In_1222,In_803);
xor U2190 (N_2190,In_244,In_1186);
nand U2191 (N_2191,In_924,In_59);
nor U2192 (N_2192,In_1065,In_36);
nor U2193 (N_2193,In_1359,In_495);
nor U2194 (N_2194,In_352,In_73);
nor U2195 (N_2195,In_876,In_940);
nor U2196 (N_2196,In_272,In_456);
nor U2197 (N_2197,In_381,In_230);
nand U2198 (N_2198,In_670,In_584);
nand U2199 (N_2199,In_1342,In_470);
xnor U2200 (N_2200,In_756,In_516);
xnor U2201 (N_2201,In_1148,In_231);
nand U2202 (N_2202,In_552,In_1152);
nor U2203 (N_2203,In_680,In_551);
or U2204 (N_2204,In_404,In_1390);
nor U2205 (N_2205,In_1455,In_1412);
and U2206 (N_2206,In_894,In_1376);
xnor U2207 (N_2207,In_88,In_556);
xnor U2208 (N_2208,In_1136,In_678);
nand U2209 (N_2209,In_909,In_993);
nand U2210 (N_2210,In_727,In_774);
nand U2211 (N_2211,In_1157,In_834);
nor U2212 (N_2212,In_1217,In_164);
nor U2213 (N_2213,In_1068,In_477);
and U2214 (N_2214,In_1154,In_784);
nand U2215 (N_2215,In_1418,In_833);
or U2216 (N_2216,In_504,In_278);
and U2217 (N_2217,In_1081,In_1294);
and U2218 (N_2218,In_196,In_1482);
xor U2219 (N_2219,In_117,In_72);
or U2220 (N_2220,In_1090,In_54);
and U2221 (N_2221,In_861,In_1372);
nor U2222 (N_2222,In_867,In_654);
nor U2223 (N_2223,In_440,In_252);
xnor U2224 (N_2224,In_1427,In_1125);
and U2225 (N_2225,In_454,In_1198);
xor U2226 (N_2226,In_1359,In_816);
xnor U2227 (N_2227,In_665,In_863);
nor U2228 (N_2228,In_663,In_871);
and U2229 (N_2229,In_823,In_294);
nor U2230 (N_2230,In_1453,In_5);
and U2231 (N_2231,In_558,In_74);
and U2232 (N_2232,In_20,In_979);
or U2233 (N_2233,In_991,In_821);
nor U2234 (N_2234,In_1275,In_414);
xor U2235 (N_2235,In_913,In_1142);
and U2236 (N_2236,In_471,In_767);
xnor U2237 (N_2237,In_133,In_508);
nor U2238 (N_2238,In_41,In_920);
nor U2239 (N_2239,In_268,In_903);
nand U2240 (N_2240,In_432,In_756);
nand U2241 (N_2241,In_212,In_920);
nor U2242 (N_2242,In_332,In_1288);
nor U2243 (N_2243,In_437,In_1424);
and U2244 (N_2244,In_901,In_338);
nand U2245 (N_2245,In_1067,In_364);
nor U2246 (N_2246,In_843,In_253);
or U2247 (N_2247,In_837,In_242);
or U2248 (N_2248,In_1304,In_911);
and U2249 (N_2249,In_41,In_821);
nor U2250 (N_2250,In_239,In_1324);
nand U2251 (N_2251,In_104,In_108);
xnor U2252 (N_2252,In_1410,In_762);
xor U2253 (N_2253,In_1061,In_441);
nand U2254 (N_2254,In_953,In_305);
nor U2255 (N_2255,In_331,In_270);
or U2256 (N_2256,In_237,In_1120);
and U2257 (N_2257,In_720,In_1260);
xor U2258 (N_2258,In_304,In_1054);
xnor U2259 (N_2259,In_303,In_1267);
xnor U2260 (N_2260,In_197,In_73);
nand U2261 (N_2261,In_59,In_921);
nand U2262 (N_2262,In_737,In_63);
xnor U2263 (N_2263,In_98,In_583);
nor U2264 (N_2264,In_1476,In_317);
nand U2265 (N_2265,In_1168,In_618);
nor U2266 (N_2266,In_1361,In_772);
nand U2267 (N_2267,In_69,In_43);
nand U2268 (N_2268,In_617,In_109);
nand U2269 (N_2269,In_560,In_993);
or U2270 (N_2270,In_297,In_744);
and U2271 (N_2271,In_689,In_1225);
nand U2272 (N_2272,In_94,In_663);
nand U2273 (N_2273,In_372,In_129);
xnor U2274 (N_2274,In_1478,In_838);
and U2275 (N_2275,In_931,In_1322);
or U2276 (N_2276,In_1208,In_1345);
xor U2277 (N_2277,In_1056,In_80);
nand U2278 (N_2278,In_1013,In_1201);
or U2279 (N_2279,In_122,In_626);
and U2280 (N_2280,In_811,In_1026);
nand U2281 (N_2281,In_176,In_610);
nand U2282 (N_2282,In_1110,In_1206);
nand U2283 (N_2283,In_123,In_1118);
nor U2284 (N_2284,In_250,In_669);
xor U2285 (N_2285,In_1209,In_694);
nand U2286 (N_2286,In_63,In_741);
xor U2287 (N_2287,In_182,In_459);
and U2288 (N_2288,In_1255,In_1209);
nor U2289 (N_2289,In_1080,In_231);
xnor U2290 (N_2290,In_279,In_1185);
nand U2291 (N_2291,In_736,In_1275);
nand U2292 (N_2292,In_415,In_74);
or U2293 (N_2293,In_194,In_937);
nor U2294 (N_2294,In_1361,In_865);
and U2295 (N_2295,In_900,In_67);
nor U2296 (N_2296,In_634,In_970);
nor U2297 (N_2297,In_390,In_88);
and U2298 (N_2298,In_515,In_42);
nand U2299 (N_2299,In_1235,In_435);
nor U2300 (N_2300,In_1064,In_228);
xor U2301 (N_2301,In_1144,In_456);
nand U2302 (N_2302,In_670,In_221);
nand U2303 (N_2303,In_1030,In_1126);
nand U2304 (N_2304,In_1359,In_501);
nand U2305 (N_2305,In_720,In_890);
nand U2306 (N_2306,In_1098,In_770);
nor U2307 (N_2307,In_247,In_923);
or U2308 (N_2308,In_78,In_135);
nor U2309 (N_2309,In_284,In_706);
and U2310 (N_2310,In_309,In_306);
or U2311 (N_2311,In_416,In_522);
and U2312 (N_2312,In_127,In_232);
nor U2313 (N_2313,In_739,In_533);
nand U2314 (N_2314,In_1221,In_330);
nor U2315 (N_2315,In_1182,In_18);
nor U2316 (N_2316,In_246,In_515);
and U2317 (N_2317,In_1104,In_703);
xor U2318 (N_2318,In_299,In_1451);
nand U2319 (N_2319,In_1180,In_1403);
and U2320 (N_2320,In_435,In_791);
xor U2321 (N_2321,In_813,In_360);
nor U2322 (N_2322,In_996,In_209);
and U2323 (N_2323,In_642,In_1124);
nor U2324 (N_2324,In_92,In_1070);
and U2325 (N_2325,In_759,In_1181);
or U2326 (N_2326,In_752,In_799);
or U2327 (N_2327,In_110,In_290);
or U2328 (N_2328,In_1132,In_486);
and U2329 (N_2329,In_1063,In_283);
or U2330 (N_2330,In_162,In_700);
xnor U2331 (N_2331,In_232,In_792);
or U2332 (N_2332,In_1399,In_1191);
or U2333 (N_2333,In_1335,In_1230);
and U2334 (N_2334,In_1392,In_833);
nand U2335 (N_2335,In_584,In_1152);
nand U2336 (N_2336,In_18,In_700);
nand U2337 (N_2337,In_1145,In_25);
xnor U2338 (N_2338,In_1004,In_786);
or U2339 (N_2339,In_468,In_498);
or U2340 (N_2340,In_647,In_296);
nand U2341 (N_2341,In_792,In_265);
nand U2342 (N_2342,In_482,In_324);
xor U2343 (N_2343,In_5,In_349);
nand U2344 (N_2344,In_1457,In_880);
or U2345 (N_2345,In_153,In_1409);
or U2346 (N_2346,In_625,In_249);
nand U2347 (N_2347,In_818,In_1202);
xor U2348 (N_2348,In_909,In_144);
or U2349 (N_2349,In_599,In_561);
or U2350 (N_2350,In_1309,In_407);
or U2351 (N_2351,In_256,In_47);
nand U2352 (N_2352,In_1308,In_113);
and U2353 (N_2353,In_1147,In_229);
xor U2354 (N_2354,In_301,In_251);
or U2355 (N_2355,In_249,In_1458);
or U2356 (N_2356,In_558,In_1399);
and U2357 (N_2357,In_24,In_48);
or U2358 (N_2358,In_1075,In_1191);
and U2359 (N_2359,In_716,In_257);
or U2360 (N_2360,In_1183,In_999);
xnor U2361 (N_2361,In_805,In_559);
and U2362 (N_2362,In_1221,In_1125);
and U2363 (N_2363,In_204,In_551);
nor U2364 (N_2364,In_1019,In_583);
nand U2365 (N_2365,In_41,In_155);
and U2366 (N_2366,In_744,In_5);
and U2367 (N_2367,In_499,In_1468);
nor U2368 (N_2368,In_257,In_79);
nor U2369 (N_2369,In_1076,In_396);
nand U2370 (N_2370,In_949,In_177);
or U2371 (N_2371,In_325,In_278);
nand U2372 (N_2372,In_19,In_480);
xor U2373 (N_2373,In_70,In_740);
xor U2374 (N_2374,In_257,In_1377);
xnor U2375 (N_2375,In_1053,In_574);
or U2376 (N_2376,In_584,In_874);
nor U2377 (N_2377,In_511,In_1452);
and U2378 (N_2378,In_869,In_1176);
nand U2379 (N_2379,In_330,In_1071);
and U2380 (N_2380,In_974,In_485);
xor U2381 (N_2381,In_1119,In_394);
or U2382 (N_2382,In_1367,In_1176);
nand U2383 (N_2383,In_1334,In_555);
nand U2384 (N_2384,In_611,In_130);
xnor U2385 (N_2385,In_833,In_76);
nor U2386 (N_2386,In_438,In_229);
xor U2387 (N_2387,In_73,In_663);
xnor U2388 (N_2388,In_290,In_1462);
nor U2389 (N_2389,In_200,In_644);
or U2390 (N_2390,In_1057,In_1424);
nand U2391 (N_2391,In_916,In_158);
or U2392 (N_2392,In_781,In_664);
xnor U2393 (N_2393,In_1367,In_690);
nor U2394 (N_2394,In_382,In_866);
xnor U2395 (N_2395,In_722,In_1209);
xor U2396 (N_2396,In_1416,In_364);
nor U2397 (N_2397,In_1424,In_747);
and U2398 (N_2398,In_299,In_92);
and U2399 (N_2399,In_653,In_387);
nand U2400 (N_2400,In_470,In_648);
xor U2401 (N_2401,In_906,In_471);
xnor U2402 (N_2402,In_408,In_91);
nand U2403 (N_2403,In_765,In_924);
xor U2404 (N_2404,In_22,In_635);
nand U2405 (N_2405,In_525,In_158);
or U2406 (N_2406,In_798,In_1088);
xor U2407 (N_2407,In_588,In_571);
nor U2408 (N_2408,In_1035,In_1393);
xor U2409 (N_2409,In_708,In_1291);
nand U2410 (N_2410,In_1130,In_1100);
nor U2411 (N_2411,In_1348,In_97);
xor U2412 (N_2412,In_1188,In_984);
and U2413 (N_2413,In_644,In_109);
or U2414 (N_2414,In_721,In_668);
or U2415 (N_2415,In_752,In_10);
xnor U2416 (N_2416,In_142,In_832);
nand U2417 (N_2417,In_393,In_517);
nor U2418 (N_2418,In_1135,In_69);
nor U2419 (N_2419,In_1125,In_1257);
nor U2420 (N_2420,In_1445,In_1335);
and U2421 (N_2421,In_929,In_765);
and U2422 (N_2422,In_402,In_1278);
or U2423 (N_2423,In_359,In_1459);
xnor U2424 (N_2424,In_653,In_556);
nor U2425 (N_2425,In_374,In_170);
and U2426 (N_2426,In_385,In_719);
nand U2427 (N_2427,In_931,In_831);
xnor U2428 (N_2428,In_339,In_1069);
xor U2429 (N_2429,In_996,In_993);
and U2430 (N_2430,In_1351,In_1447);
nor U2431 (N_2431,In_404,In_311);
and U2432 (N_2432,In_96,In_315);
nor U2433 (N_2433,In_1132,In_689);
or U2434 (N_2434,In_1238,In_1385);
nor U2435 (N_2435,In_659,In_4);
xnor U2436 (N_2436,In_1065,In_1278);
xnor U2437 (N_2437,In_534,In_1197);
nand U2438 (N_2438,In_288,In_196);
nand U2439 (N_2439,In_31,In_271);
nor U2440 (N_2440,In_706,In_384);
or U2441 (N_2441,In_1233,In_1061);
nor U2442 (N_2442,In_1455,In_1034);
or U2443 (N_2443,In_360,In_30);
and U2444 (N_2444,In_190,In_1350);
nor U2445 (N_2445,In_856,In_626);
nor U2446 (N_2446,In_435,In_601);
xnor U2447 (N_2447,In_827,In_987);
xnor U2448 (N_2448,In_729,In_635);
xnor U2449 (N_2449,In_1171,In_729);
nand U2450 (N_2450,In_1414,In_636);
nor U2451 (N_2451,In_922,In_235);
nand U2452 (N_2452,In_601,In_13);
nand U2453 (N_2453,In_948,In_757);
and U2454 (N_2454,In_64,In_311);
nor U2455 (N_2455,In_1161,In_172);
nand U2456 (N_2456,In_133,In_1352);
and U2457 (N_2457,In_30,In_1494);
nor U2458 (N_2458,In_88,In_464);
or U2459 (N_2459,In_95,In_1487);
xor U2460 (N_2460,In_1315,In_912);
and U2461 (N_2461,In_1394,In_1186);
and U2462 (N_2462,In_980,In_744);
or U2463 (N_2463,In_952,In_990);
nor U2464 (N_2464,In_826,In_1462);
xor U2465 (N_2465,In_1160,In_617);
nand U2466 (N_2466,In_47,In_1068);
and U2467 (N_2467,In_290,In_745);
and U2468 (N_2468,In_474,In_1242);
xnor U2469 (N_2469,In_195,In_159);
or U2470 (N_2470,In_1448,In_297);
xor U2471 (N_2471,In_975,In_762);
xnor U2472 (N_2472,In_1423,In_1288);
or U2473 (N_2473,In_813,In_372);
and U2474 (N_2474,In_1276,In_707);
and U2475 (N_2475,In_834,In_543);
or U2476 (N_2476,In_57,In_193);
nand U2477 (N_2477,In_610,In_652);
xor U2478 (N_2478,In_642,In_1100);
xor U2479 (N_2479,In_6,In_470);
or U2480 (N_2480,In_1330,In_120);
nor U2481 (N_2481,In_675,In_973);
nor U2482 (N_2482,In_384,In_389);
nand U2483 (N_2483,In_800,In_1308);
nor U2484 (N_2484,In_233,In_480);
and U2485 (N_2485,In_739,In_1083);
nand U2486 (N_2486,In_778,In_760);
and U2487 (N_2487,In_1100,In_1184);
xor U2488 (N_2488,In_1164,In_940);
xor U2489 (N_2489,In_839,In_1272);
nand U2490 (N_2490,In_1471,In_1356);
xnor U2491 (N_2491,In_1007,In_449);
nand U2492 (N_2492,In_1183,In_1315);
and U2493 (N_2493,In_96,In_44);
nand U2494 (N_2494,In_710,In_1083);
xor U2495 (N_2495,In_150,In_1126);
and U2496 (N_2496,In_1197,In_1372);
nor U2497 (N_2497,In_1288,In_407);
xnor U2498 (N_2498,In_273,In_886);
or U2499 (N_2499,In_387,In_825);
nand U2500 (N_2500,In_951,In_30);
and U2501 (N_2501,In_71,In_905);
xnor U2502 (N_2502,In_413,In_661);
nand U2503 (N_2503,In_502,In_160);
nand U2504 (N_2504,In_1171,In_1365);
or U2505 (N_2505,In_817,In_114);
and U2506 (N_2506,In_1322,In_370);
and U2507 (N_2507,In_1434,In_648);
or U2508 (N_2508,In_699,In_192);
and U2509 (N_2509,In_866,In_1032);
and U2510 (N_2510,In_46,In_209);
or U2511 (N_2511,In_1485,In_474);
nor U2512 (N_2512,In_901,In_1360);
and U2513 (N_2513,In_187,In_537);
and U2514 (N_2514,In_1267,In_823);
and U2515 (N_2515,In_926,In_653);
and U2516 (N_2516,In_1310,In_162);
and U2517 (N_2517,In_292,In_637);
nand U2518 (N_2518,In_430,In_374);
xor U2519 (N_2519,In_904,In_1324);
nor U2520 (N_2520,In_1337,In_1297);
or U2521 (N_2521,In_854,In_801);
nor U2522 (N_2522,In_1053,In_737);
nand U2523 (N_2523,In_740,In_304);
or U2524 (N_2524,In_274,In_613);
nand U2525 (N_2525,In_140,In_1326);
nand U2526 (N_2526,In_699,In_40);
or U2527 (N_2527,In_732,In_397);
or U2528 (N_2528,In_959,In_685);
nand U2529 (N_2529,In_1404,In_1367);
or U2530 (N_2530,In_1026,In_1015);
and U2531 (N_2531,In_284,In_1346);
xnor U2532 (N_2532,In_1084,In_1289);
or U2533 (N_2533,In_874,In_1192);
xor U2534 (N_2534,In_249,In_765);
nor U2535 (N_2535,In_517,In_145);
and U2536 (N_2536,In_100,In_1272);
or U2537 (N_2537,In_1485,In_818);
or U2538 (N_2538,In_1277,In_551);
or U2539 (N_2539,In_397,In_1313);
nor U2540 (N_2540,In_273,In_539);
and U2541 (N_2541,In_703,In_1157);
or U2542 (N_2542,In_1087,In_1159);
nand U2543 (N_2543,In_944,In_382);
or U2544 (N_2544,In_960,In_1289);
nand U2545 (N_2545,In_1000,In_1031);
or U2546 (N_2546,In_81,In_507);
and U2547 (N_2547,In_1429,In_786);
xor U2548 (N_2548,In_1027,In_662);
nor U2549 (N_2549,In_675,In_1207);
xnor U2550 (N_2550,In_1205,In_1227);
and U2551 (N_2551,In_282,In_529);
or U2552 (N_2552,In_574,In_1238);
nand U2553 (N_2553,In_1173,In_1162);
xor U2554 (N_2554,In_743,In_421);
or U2555 (N_2555,In_461,In_514);
nor U2556 (N_2556,In_1283,In_621);
or U2557 (N_2557,In_1400,In_1276);
xnor U2558 (N_2558,In_570,In_44);
and U2559 (N_2559,In_708,In_1427);
nand U2560 (N_2560,In_86,In_254);
nor U2561 (N_2561,In_260,In_517);
nor U2562 (N_2562,In_1199,In_1013);
and U2563 (N_2563,In_374,In_951);
nor U2564 (N_2564,In_603,In_77);
xor U2565 (N_2565,In_1490,In_434);
nand U2566 (N_2566,In_162,In_78);
nor U2567 (N_2567,In_1405,In_1012);
xor U2568 (N_2568,In_1421,In_951);
or U2569 (N_2569,In_128,In_870);
xnor U2570 (N_2570,In_638,In_74);
nor U2571 (N_2571,In_832,In_825);
xnor U2572 (N_2572,In_124,In_1353);
nand U2573 (N_2573,In_375,In_525);
nor U2574 (N_2574,In_609,In_1060);
nor U2575 (N_2575,In_59,In_1007);
nand U2576 (N_2576,In_719,In_111);
nor U2577 (N_2577,In_665,In_1171);
and U2578 (N_2578,In_1002,In_598);
or U2579 (N_2579,In_128,In_1491);
nand U2580 (N_2580,In_692,In_716);
nand U2581 (N_2581,In_1128,In_1375);
xor U2582 (N_2582,In_687,In_1131);
nor U2583 (N_2583,In_278,In_505);
nor U2584 (N_2584,In_1483,In_1233);
and U2585 (N_2585,In_1209,In_1380);
or U2586 (N_2586,In_826,In_1466);
xnor U2587 (N_2587,In_356,In_959);
xnor U2588 (N_2588,In_400,In_452);
or U2589 (N_2589,In_1405,In_1353);
nor U2590 (N_2590,In_1007,In_1439);
nand U2591 (N_2591,In_224,In_1147);
or U2592 (N_2592,In_960,In_1058);
nand U2593 (N_2593,In_868,In_1136);
and U2594 (N_2594,In_633,In_1257);
and U2595 (N_2595,In_1139,In_568);
nand U2596 (N_2596,In_1363,In_630);
nor U2597 (N_2597,In_492,In_933);
nand U2598 (N_2598,In_176,In_787);
and U2599 (N_2599,In_77,In_270);
xor U2600 (N_2600,In_1133,In_22);
nand U2601 (N_2601,In_1150,In_934);
nand U2602 (N_2602,In_710,In_1388);
nand U2603 (N_2603,In_1446,In_90);
nand U2604 (N_2604,In_1364,In_971);
or U2605 (N_2605,In_613,In_628);
nor U2606 (N_2606,In_1130,In_225);
and U2607 (N_2607,In_519,In_281);
nor U2608 (N_2608,In_629,In_750);
nand U2609 (N_2609,In_677,In_734);
nand U2610 (N_2610,In_123,In_1069);
nor U2611 (N_2611,In_431,In_618);
nor U2612 (N_2612,In_606,In_119);
nor U2613 (N_2613,In_369,In_614);
and U2614 (N_2614,In_101,In_541);
xnor U2615 (N_2615,In_141,In_44);
nor U2616 (N_2616,In_838,In_463);
and U2617 (N_2617,In_1283,In_1248);
nand U2618 (N_2618,In_388,In_218);
nand U2619 (N_2619,In_904,In_776);
nor U2620 (N_2620,In_184,In_272);
nand U2621 (N_2621,In_1,In_436);
and U2622 (N_2622,In_569,In_535);
and U2623 (N_2623,In_1373,In_558);
and U2624 (N_2624,In_1076,In_217);
xor U2625 (N_2625,In_586,In_912);
and U2626 (N_2626,In_667,In_877);
nand U2627 (N_2627,In_803,In_692);
nand U2628 (N_2628,In_832,In_770);
or U2629 (N_2629,In_366,In_388);
nor U2630 (N_2630,In_251,In_1289);
xnor U2631 (N_2631,In_982,In_674);
nor U2632 (N_2632,In_615,In_1025);
nor U2633 (N_2633,In_1417,In_1363);
nand U2634 (N_2634,In_283,In_234);
nor U2635 (N_2635,In_544,In_618);
xnor U2636 (N_2636,In_1422,In_578);
nor U2637 (N_2637,In_1066,In_885);
nor U2638 (N_2638,In_326,In_559);
nand U2639 (N_2639,In_32,In_1149);
xor U2640 (N_2640,In_1116,In_376);
and U2641 (N_2641,In_1275,In_1277);
nand U2642 (N_2642,In_870,In_389);
xnor U2643 (N_2643,In_1245,In_279);
and U2644 (N_2644,In_344,In_1494);
and U2645 (N_2645,In_1443,In_686);
nor U2646 (N_2646,In_1271,In_168);
xor U2647 (N_2647,In_676,In_644);
xor U2648 (N_2648,In_935,In_1273);
xnor U2649 (N_2649,In_247,In_1024);
nand U2650 (N_2650,In_1058,In_1201);
nand U2651 (N_2651,In_1001,In_594);
or U2652 (N_2652,In_258,In_1326);
or U2653 (N_2653,In_1005,In_1279);
xor U2654 (N_2654,In_364,In_1382);
or U2655 (N_2655,In_301,In_935);
xnor U2656 (N_2656,In_1081,In_1454);
nand U2657 (N_2657,In_160,In_444);
nor U2658 (N_2658,In_1270,In_83);
xnor U2659 (N_2659,In_101,In_1476);
nand U2660 (N_2660,In_1494,In_45);
nand U2661 (N_2661,In_165,In_188);
nand U2662 (N_2662,In_812,In_918);
nand U2663 (N_2663,In_655,In_1315);
or U2664 (N_2664,In_1157,In_1301);
xor U2665 (N_2665,In_571,In_1414);
and U2666 (N_2666,In_1481,In_1316);
or U2667 (N_2667,In_1301,In_37);
nor U2668 (N_2668,In_1112,In_368);
and U2669 (N_2669,In_1018,In_998);
nor U2670 (N_2670,In_830,In_689);
xnor U2671 (N_2671,In_1359,In_275);
nor U2672 (N_2672,In_960,In_995);
nor U2673 (N_2673,In_1015,In_1346);
and U2674 (N_2674,In_69,In_1213);
nand U2675 (N_2675,In_395,In_774);
or U2676 (N_2676,In_847,In_260);
or U2677 (N_2677,In_185,In_861);
xnor U2678 (N_2678,In_76,In_495);
nand U2679 (N_2679,In_1471,In_807);
nand U2680 (N_2680,In_522,In_456);
nand U2681 (N_2681,In_190,In_579);
xor U2682 (N_2682,In_643,In_1051);
nand U2683 (N_2683,In_1418,In_986);
xor U2684 (N_2684,In_66,In_871);
nand U2685 (N_2685,In_1126,In_1040);
or U2686 (N_2686,In_1246,In_1086);
xnor U2687 (N_2687,In_1139,In_157);
nand U2688 (N_2688,In_938,In_700);
xnor U2689 (N_2689,In_914,In_1315);
nor U2690 (N_2690,In_7,In_504);
and U2691 (N_2691,In_529,In_1384);
or U2692 (N_2692,In_1467,In_324);
and U2693 (N_2693,In_1451,In_121);
or U2694 (N_2694,In_904,In_659);
and U2695 (N_2695,In_1012,In_98);
and U2696 (N_2696,In_262,In_510);
nand U2697 (N_2697,In_667,In_708);
and U2698 (N_2698,In_619,In_194);
xor U2699 (N_2699,In_971,In_256);
xnor U2700 (N_2700,In_753,In_1390);
nand U2701 (N_2701,In_937,In_346);
or U2702 (N_2702,In_329,In_348);
nand U2703 (N_2703,In_1220,In_1071);
nand U2704 (N_2704,In_1401,In_1345);
or U2705 (N_2705,In_581,In_963);
or U2706 (N_2706,In_1152,In_742);
and U2707 (N_2707,In_747,In_361);
nand U2708 (N_2708,In_636,In_48);
nand U2709 (N_2709,In_419,In_972);
and U2710 (N_2710,In_1239,In_870);
and U2711 (N_2711,In_1017,In_353);
or U2712 (N_2712,In_224,In_44);
nor U2713 (N_2713,In_594,In_1263);
nand U2714 (N_2714,In_663,In_1313);
and U2715 (N_2715,In_1231,In_466);
xor U2716 (N_2716,In_490,In_421);
nor U2717 (N_2717,In_927,In_830);
nand U2718 (N_2718,In_14,In_1117);
nor U2719 (N_2719,In_1218,In_1089);
nor U2720 (N_2720,In_1228,In_674);
or U2721 (N_2721,In_500,In_31);
nand U2722 (N_2722,In_551,In_776);
or U2723 (N_2723,In_399,In_1497);
xor U2724 (N_2724,In_1153,In_341);
and U2725 (N_2725,In_1055,In_390);
xnor U2726 (N_2726,In_15,In_683);
nand U2727 (N_2727,In_312,In_132);
or U2728 (N_2728,In_959,In_458);
nor U2729 (N_2729,In_290,In_1085);
xor U2730 (N_2730,In_1395,In_180);
xor U2731 (N_2731,In_227,In_748);
nand U2732 (N_2732,In_193,In_1287);
or U2733 (N_2733,In_307,In_390);
nand U2734 (N_2734,In_234,In_1331);
and U2735 (N_2735,In_1091,In_974);
nor U2736 (N_2736,In_1008,In_1007);
xnor U2737 (N_2737,In_355,In_928);
nand U2738 (N_2738,In_800,In_1398);
and U2739 (N_2739,In_1497,In_929);
nand U2740 (N_2740,In_1141,In_111);
and U2741 (N_2741,In_1222,In_1498);
nand U2742 (N_2742,In_1284,In_1076);
nor U2743 (N_2743,In_1374,In_830);
xnor U2744 (N_2744,In_650,In_22);
xor U2745 (N_2745,In_163,In_210);
or U2746 (N_2746,In_724,In_202);
nand U2747 (N_2747,In_1254,In_1337);
nand U2748 (N_2748,In_1347,In_295);
nor U2749 (N_2749,In_1035,In_1448);
and U2750 (N_2750,In_1465,In_1433);
xor U2751 (N_2751,In_610,In_977);
nor U2752 (N_2752,In_109,In_148);
nand U2753 (N_2753,In_1235,In_1437);
nor U2754 (N_2754,In_795,In_17);
nand U2755 (N_2755,In_255,In_65);
nand U2756 (N_2756,In_1012,In_402);
and U2757 (N_2757,In_1412,In_1199);
or U2758 (N_2758,In_486,In_228);
or U2759 (N_2759,In_487,In_594);
or U2760 (N_2760,In_1218,In_65);
or U2761 (N_2761,In_574,In_1185);
xnor U2762 (N_2762,In_887,In_15);
xnor U2763 (N_2763,In_143,In_810);
and U2764 (N_2764,In_1230,In_1406);
xnor U2765 (N_2765,In_1186,In_345);
xor U2766 (N_2766,In_1059,In_907);
and U2767 (N_2767,In_17,In_366);
nand U2768 (N_2768,In_932,In_727);
or U2769 (N_2769,In_1441,In_1160);
nand U2770 (N_2770,In_640,In_728);
and U2771 (N_2771,In_17,In_346);
nand U2772 (N_2772,In_1420,In_526);
nand U2773 (N_2773,In_305,In_1395);
nor U2774 (N_2774,In_1368,In_979);
nand U2775 (N_2775,In_869,In_1464);
xnor U2776 (N_2776,In_1209,In_635);
nand U2777 (N_2777,In_917,In_21);
and U2778 (N_2778,In_1029,In_263);
xnor U2779 (N_2779,In_1262,In_423);
nand U2780 (N_2780,In_1313,In_84);
nand U2781 (N_2781,In_198,In_453);
nand U2782 (N_2782,In_151,In_661);
nand U2783 (N_2783,In_714,In_841);
nor U2784 (N_2784,In_751,In_1393);
nor U2785 (N_2785,In_127,In_112);
nor U2786 (N_2786,In_744,In_1467);
nand U2787 (N_2787,In_941,In_1005);
nand U2788 (N_2788,In_52,In_1050);
nand U2789 (N_2789,In_744,In_1479);
or U2790 (N_2790,In_217,In_194);
and U2791 (N_2791,In_207,In_1050);
nor U2792 (N_2792,In_1370,In_1309);
nand U2793 (N_2793,In_766,In_426);
nand U2794 (N_2794,In_1264,In_704);
or U2795 (N_2795,In_869,In_1237);
and U2796 (N_2796,In_422,In_307);
nand U2797 (N_2797,In_1396,In_163);
and U2798 (N_2798,In_779,In_1240);
nand U2799 (N_2799,In_925,In_224);
nand U2800 (N_2800,In_293,In_617);
xnor U2801 (N_2801,In_590,In_440);
xnor U2802 (N_2802,In_282,In_467);
nor U2803 (N_2803,In_662,In_348);
nor U2804 (N_2804,In_1378,In_1141);
nand U2805 (N_2805,In_1139,In_752);
or U2806 (N_2806,In_1018,In_120);
xnor U2807 (N_2807,In_1385,In_1218);
xor U2808 (N_2808,In_64,In_1033);
nand U2809 (N_2809,In_754,In_513);
and U2810 (N_2810,In_390,In_650);
or U2811 (N_2811,In_1224,In_373);
or U2812 (N_2812,In_289,In_464);
xor U2813 (N_2813,In_93,In_1445);
nor U2814 (N_2814,In_889,In_468);
nand U2815 (N_2815,In_108,In_844);
nor U2816 (N_2816,In_471,In_256);
nand U2817 (N_2817,In_292,In_675);
or U2818 (N_2818,In_724,In_692);
nor U2819 (N_2819,In_400,In_1002);
xor U2820 (N_2820,In_716,In_427);
xor U2821 (N_2821,In_1075,In_369);
and U2822 (N_2822,In_475,In_1324);
xor U2823 (N_2823,In_1386,In_149);
nor U2824 (N_2824,In_1094,In_1319);
xnor U2825 (N_2825,In_218,In_674);
nand U2826 (N_2826,In_1123,In_439);
nor U2827 (N_2827,In_54,In_350);
and U2828 (N_2828,In_1300,In_1193);
nor U2829 (N_2829,In_375,In_566);
nand U2830 (N_2830,In_1134,In_1491);
xor U2831 (N_2831,In_188,In_244);
or U2832 (N_2832,In_1448,In_279);
xnor U2833 (N_2833,In_553,In_150);
nor U2834 (N_2834,In_79,In_46);
and U2835 (N_2835,In_66,In_537);
nor U2836 (N_2836,In_1355,In_290);
nor U2837 (N_2837,In_841,In_343);
or U2838 (N_2838,In_1239,In_219);
and U2839 (N_2839,In_1057,In_320);
or U2840 (N_2840,In_916,In_723);
or U2841 (N_2841,In_46,In_219);
nor U2842 (N_2842,In_93,In_734);
nand U2843 (N_2843,In_1200,In_81);
and U2844 (N_2844,In_837,In_682);
xnor U2845 (N_2845,In_533,In_1054);
nand U2846 (N_2846,In_44,In_480);
xor U2847 (N_2847,In_1408,In_184);
or U2848 (N_2848,In_406,In_1494);
nand U2849 (N_2849,In_1125,In_1422);
or U2850 (N_2850,In_1049,In_973);
nand U2851 (N_2851,In_356,In_646);
and U2852 (N_2852,In_1437,In_1394);
and U2853 (N_2853,In_513,In_749);
and U2854 (N_2854,In_496,In_40);
nor U2855 (N_2855,In_1372,In_1133);
or U2856 (N_2856,In_544,In_1360);
nand U2857 (N_2857,In_1462,In_657);
nor U2858 (N_2858,In_17,In_422);
and U2859 (N_2859,In_147,In_444);
or U2860 (N_2860,In_958,In_24);
nor U2861 (N_2861,In_1224,In_1453);
xor U2862 (N_2862,In_1239,In_83);
and U2863 (N_2863,In_1100,In_1128);
nand U2864 (N_2864,In_1258,In_742);
nand U2865 (N_2865,In_561,In_861);
or U2866 (N_2866,In_530,In_0);
or U2867 (N_2867,In_1398,In_29);
nand U2868 (N_2868,In_176,In_234);
and U2869 (N_2869,In_521,In_68);
nor U2870 (N_2870,In_844,In_705);
nor U2871 (N_2871,In_801,In_620);
and U2872 (N_2872,In_139,In_751);
and U2873 (N_2873,In_237,In_1074);
nand U2874 (N_2874,In_262,In_381);
xor U2875 (N_2875,In_339,In_202);
or U2876 (N_2876,In_496,In_642);
and U2877 (N_2877,In_352,In_674);
nand U2878 (N_2878,In_858,In_1136);
or U2879 (N_2879,In_975,In_24);
nor U2880 (N_2880,In_1267,In_648);
xnor U2881 (N_2881,In_1497,In_473);
xnor U2882 (N_2882,In_1407,In_741);
nor U2883 (N_2883,In_548,In_96);
xnor U2884 (N_2884,In_1161,In_788);
and U2885 (N_2885,In_209,In_1184);
nor U2886 (N_2886,In_868,In_956);
nor U2887 (N_2887,In_640,In_559);
nor U2888 (N_2888,In_1348,In_1465);
or U2889 (N_2889,In_526,In_1465);
xor U2890 (N_2890,In_111,In_112);
nand U2891 (N_2891,In_818,In_146);
nand U2892 (N_2892,In_813,In_186);
and U2893 (N_2893,In_722,In_366);
nand U2894 (N_2894,In_758,In_533);
nor U2895 (N_2895,In_616,In_454);
xnor U2896 (N_2896,In_499,In_919);
nor U2897 (N_2897,In_590,In_1073);
xnor U2898 (N_2898,In_727,In_930);
nand U2899 (N_2899,In_838,In_457);
nand U2900 (N_2900,In_861,In_326);
nand U2901 (N_2901,In_199,In_35);
nand U2902 (N_2902,In_220,In_117);
or U2903 (N_2903,In_813,In_431);
or U2904 (N_2904,In_773,In_334);
and U2905 (N_2905,In_860,In_950);
and U2906 (N_2906,In_213,In_1068);
or U2907 (N_2907,In_1179,In_1108);
nor U2908 (N_2908,In_1194,In_321);
nand U2909 (N_2909,In_1185,In_146);
nand U2910 (N_2910,In_1107,In_29);
xor U2911 (N_2911,In_1454,In_311);
and U2912 (N_2912,In_1062,In_1163);
nand U2913 (N_2913,In_326,In_311);
or U2914 (N_2914,In_979,In_329);
and U2915 (N_2915,In_1408,In_836);
nor U2916 (N_2916,In_111,In_612);
and U2917 (N_2917,In_446,In_1305);
nor U2918 (N_2918,In_1224,In_798);
nand U2919 (N_2919,In_53,In_1369);
nand U2920 (N_2920,In_142,In_269);
nand U2921 (N_2921,In_963,In_39);
or U2922 (N_2922,In_1443,In_1294);
or U2923 (N_2923,In_409,In_840);
and U2924 (N_2924,In_829,In_100);
and U2925 (N_2925,In_891,In_1127);
or U2926 (N_2926,In_1251,In_333);
xor U2927 (N_2927,In_374,In_1479);
and U2928 (N_2928,In_208,In_601);
and U2929 (N_2929,In_1031,In_1369);
nand U2930 (N_2930,In_772,In_1345);
xnor U2931 (N_2931,In_1230,In_744);
nor U2932 (N_2932,In_1048,In_809);
xor U2933 (N_2933,In_50,In_181);
nor U2934 (N_2934,In_431,In_354);
nor U2935 (N_2935,In_1451,In_758);
and U2936 (N_2936,In_120,In_1165);
or U2937 (N_2937,In_644,In_1466);
nor U2938 (N_2938,In_607,In_1210);
nand U2939 (N_2939,In_1473,In_698);
xnor U2940 (N_2940,In_1111,In_1143);
and U2941 (N_2941,In_1282,In_254);
or U2942 (N_2942,In_1413,In_1064);
nor U2943 (N_2943,In_1085,In_1439);
or U2944 (N_2944,In_951,In_1183);
xor U2945 (N_2945,In_897,In_1073);
or U2946 (N_2946,In_279,In_109);
and U2947 (N_2947,In_516,In_915);
and U2948 (N_2948,In_575,In_1486);
or U2949 (N_2949,In_587,In_951);
xnor U2950 (N_2950,In_981,In_1126);
nor U2951 (N_2951,In_810,In_395);
or U2952 (N_2952,In_262,In_499);
nand U2953 (N_2953,In_163,In_336);
xor U2954 (N_2954,In_880,In_807);
and U2955 (N_2955,In_558,In_889);
and U2956 (N_2956,In_877,In_1144);
nand U2957 (N_2957,In_990,In_187);
nor U2958 (N_2958,In_1348,In_804);
xor U2959 (N_2959,In_176,In_131);
and U2960 (N_2960,In_937,In_1497);
nand U2961 (N_2961,In_1284,In_162);
or U2962 (N_2962,In_1012,In_791);
and U2963 (N_2963,In_1045,In_270);
or U2964 (N_2964,In_1253,In_964);
nor U2965 (N_2965,In_213,In_117);
nand U2966 (N_2966,In_1308,In_43);
nand U2967 (N_2967,In_1198,In_544);
or U2968 (N_2968,In_559,In_297);
nand U2969 (N_2969,In_1271,In_606);
nor U2970 (N_2970,In_1363,In_1313);
or U2971 (N_2971,In_563,In_1319);
nand U2972 (N_2972,In_685,In_849);
and U2973 (N_2973,In_298,In_686);
xor U2974 (N_2974,In_805,In_80);
nor U2975 (N_2975,In_884,In_523);
nand U2976 (N_2976,In_242,In_1322);
xor U2977 (N_2977,In_1352,In_839);
nand U2978 (N_2978,In_63,In_1378);
nor U2979 (N_2979,In_32,In_158);
nor U2980 (N_2980,In_1269,In_145);
nor U2981 (N_2981,In_395,In_1060);
xor U2982 (N_2982,In_505,In_483);
nor U2983 (N_2983,In_1182,In_133);
or U2984 (N_2984,In_1489,In_1280);
xnor U2985 (N_2985,In_774,In_233);
nor U2986 (N_2986,In_636,In_1025);
and U2987 (N_2987,In_606,In_354);
nor U2988 (N_2988,In_868,In_893);
nand U2989 (N_2989,In_825,In_638);
and U2990 (N_2990,In_232,In_1423);
and U2991 (N_2991,In_1045,In_827);
or U2992 (N_2992,In_71,In_1475);
xor U2993 (N_2993,In_886,In_1364);
xnor U2994 (N_2994,In_747,In_1078);
xor U2995 (N_2995,In_1433,In_571);
and U2996 (N_2996,In_531,In_332);
xnor U2997 (N_2997,In_922,In_512);
and U2998 (N_2998,In_551,In_1228);
xor U2999 (N_2999,In_1481,In_953);
xor U3000 (N_3000,In_734,In_1355);
or U3001 (N_3001,In_76,In_359);
xor U3002 (N_3002,In_1112,In_1452);
nand U3003 (N_3003,In_1152,In_863);
or U3004 (N_3004,In_78,In_788);
nand U3005 (N_3005,In_157,In_1258);
or U3006 (N_3006,In_1430,In_1128);
and U3007 (N_3007,In_1451,In_162);
nand U3008 (N_3008,In_905,In_1492);
nand U3009 (N_3009,In_145,In_123);
nand U3010 (N_3010,In_241,In_1063);
xor U3011 (N_3011,In_1191,In_546);
or U3012 (N_3012,In_1041,In_313);
or U3013 (N_3013,In_1142,In_334);
or U3014 (N_3014,In_672,In_865);
and U3015 (N_3015,In_514,In_143);
xor U3016 (N_3016,In_412,In_1409);
nand U3017 (N_3017,In_697,In_646);
nand U3018 (N_3018,In_1099,In_804);
or U3019 (N_3019,In_168,In_384);
xnor U3020 (N_3020,In_1315,In_684);
and U3021 (N_3021,In_310,In_874);
and U3022 (N_3022,In_1407,In_527);
xnor U3023 (N_3023,In_1419,In_177);
xor U3024 (N_3024,In_1041,In_793);
xor U3025 (N_3025,In_352,In_1375);
and U3026 (N_3026,In_1130,In_867);
or U3027 (N_3027,In_1315,In_1215);
or U3028 (N_3028,In_1424,In_351);
xor U3029 (N_3029,In_743,In_266);
nor U3030 (N_3030,In_1266,In_588);
nand U3031 (N_3031,In_1498,In_1366);
nand U3032 (N_3032,In_578,In_266);
nor U3033 (N_3033,In_849,In_843);
or U3034 (N_3034,In_1340,In_739);
xor U3035 (N_3035,In_1228,In_985);
and U3036 (N_3036,In_1493,In_186);
and U3037 (N_3037,In_1265,In_743);
or U3038 (N_3038,In_652,In_769);
or U3039 (N_3039,In_452,In_405);
nor U3040 (N_3040,In_774,In_1029);
or U3041 (N_3041,In_75,In_660);
nand U3042 (N_3042,In_849,In_792);
and U3043 (N_3043,In_1422,In_725);
or U3044 (N_3044,In_1065,In_1081);
or U3045 (N_3045,In_37,In_608);
nor U3046 (N_3046,In_1480,In_1103);
nor U3047 (N_3047,In_793,In_1195);
nor U3048 (N_3048,In_1124,In_1215);
or U3049 (N_3049,In_412,In_343);
xor U3050 (N_3050,In_516,In_934);
and U3051 (N_3051,In_878,In_584);
or U3052 (N_3052,In_785,In_94);
nor U3053 (N_3053,In_668,In_650);
nor U3054 (N_3054,In_140,In_274);
xnor U3055 (N_3055,In_94,In_908);
and U3056 (N_3056,In_1130,In_420);
nor U3057 (N_3057,In_950,In_1483);
xnor U3058 (N_3058,In_1014,In_674);
nand U3059 (N_3059,In_165,In_1124);
and U3060 (N_3060,In_62,In_1306);
xor U3061 (N_3061,In_227,In_357);
or U3062 (N_3062,In_251,In_0);
or U3063 (N_3063,In_198,In_111);
or U3064 (N_3064,In_1497,In_889);
nor U3065 (N_3065,In_1199,In_1361);
nor U3066 (N_3066,In_989,In_494);
or U3067 (N_3067,In_1422,In_498);
and U3068 (N_3068,In_222,In_755);
nor U3069 (N_3069,In_40,In_620);
nor U3070 (N_3070,In_386,In_1314);
nor U3071 (N_3071,In_258,In_1464);
and U3072 (N_3072,In_1456,In_1361);
nor U3073 (N_3073,In_232,In_1041);
xnor U3074 (N_3074,In_1214,In_953);
nor U3075 (N_3075,In_1425,In_863);
nand U3076 (N_3076,In_1084,In_634);
nor U3077 (N_3077,In_661,In_1233);
and U3078 (N_3078,In_921,In_1186);
and U3079 (N_3079,In_551,In_435);
and U3080 (N_3080,In_968,In_496);
and U3081 (N_3081,In_810,In_990);
xnor U3082 (N_3082,In_25,In_1467);
nand U3083 (N_3083,In_249,In_978);
and U3084 (N_3084,In_214,In_1226);
nor U3085 (N_3085,In_635,In_1218);
or U3086 (N_3086,In_672,In_1124);
nor U3087 (N_3087,In_1375,In_515);
nand U3088 (N_3088,In_611,In_0);
or U3089 (N_3089,In_468,In_188);
and U3090 (N_3090,In_1322,In_1083);
nand U3091 (N_3091,In_1345,In_1256);
or U3092 (N_3092,In_667,In_1066);
and U3093 (N_3093,In_543,In_1219);
nor U3094 (N_3094,In_285,In_1114);
or U3095 (N_3095,In_1176,In_1253);
nor U3096 (N_3096,In_505,In_5);
nand U3097 (N_3097,In_1473,In_325);
xor U3098 (N_3098,In_953,In_429);
nand U3099 (N_3099,In_58,In_1068);
nand U3100 (N_3100,In_1447,In_614);
nand U3101 (N_3101,In_839,In_1313);
xor U3102 (N_3102,In_396,In_1452);
nand U3103 (N_3103,In_181,In_1375);
nor U3104 (N_3104,In_436,In_229);
or U3105 (N_3105,In_1393,In_276);
or U3106 (N_3106,In_462,In_489);
xnor U3107 (N_3107,In_965,In_370);
or U3108 (N_3108,In_1489,In_71);
nor U3109 (N_3109,In_1085,In_826);
and U3110 (N_3110,In_971,In_503);
xor U3111 (N_3111,In_1107,In_255);
or U3112 (N_3112,In_1269,In_1049);
and U3113 (N_3113,In_1055,In_1043);
xor U3114 (N_3114,In_692,In_846);
or U3115 (N_3115,In_643,In_1398);
xnor U3116 (N_3116,In_789,In_1417);
nand U3117 (N_3117,In_1029,In_55);
xor U3118 (N_3118,In_1332,In_923);
or U3119 (N_3119,In_1006,In_893);
and U3120 (N_3120,In_30,In_552);
or U3121 (N_3121,In_489,In_1361);
nor U3122 (N_3122,In_296,In_1024);
xor U3123 (N_3123,In_551,In_1244);
nor U3124 (N_3124,In_106,In_1050);
and U3125 (N_3125,In_898,In_985);
nand U3126 (N_3126,In_1079,In_168);
or U3127 (N_3127,In_41,In_569);
xnor U3128 (N_3128,In_419,In_914);
nor U3129 (N_3129,In_554,In_1071);
nor U3130 (N_3130,In_277,In_1405);
and U3131 (N_3131,In_782,In_1353);
nand U3132 (N_3132,In_516,In_135);
nand U3133 (N_3133,In_202,In_19);
and U3134 (N_3134,In_1247,In_1091);
nand U3135 (N_3135,In_351,In_1484);
xor U3136 (N_3136,In_709,In_1404);
or U3137 (N_3137,In_1353,In_1286);
or U3138 (N_3138,In_952,In_1237);
nor U3139 (N_3139,In_1171,In_911);
nor U3140 (N_3140,In_140,In_250);
or U3141 (N_3141,In_482,In_541);
nand U3142 (N_3142,In_1450,In_214);
or U3143 (N_3143,In_1216,In_502);
or U3144 (N_3144,In_97,In_863);
nand U3145 (N_3145,In_46,In_6);
or U3146 (N_3146,In_256,In_1157);
and U3147 (N_3147,In_1275,In_597);
xor U3148 (N_3148,In_1352,In_869);
nor U3149 (N_3149,In_860,In_889);
and U3150 (N_3150,In_264,In_983);
and U3151 (N_3151,In_1054,In_1410);
nand U3152 (N_3152,In_807,In_1487);
and U3153 (N_3153,In_610,In_590);
nor U3154 (N_3154,In_183,In_1269);
nor U3155 (N_3155,In_939,In_714);
and U3156 (N_3156,In_1227,In_1258);
and U3157 (N_3157,In_107,In_26);
nor U3158 (N_3158,In_678,In_1475);
xor U3159 (N_3159,In_464,In_6);
and U3160 (N_3160,In_484,In_51);
nor U3161 (N_3161,In_954,In_457);
xor U3162 (N_3162,In_758,In_126);
or U3163 (N_3163,In_1183,In_624);
or U3164 (N_3164,In_215,In_230);
nor U3165 (N_3165,In_624,In_984);
nor U3166 (N_3166,In_161,In_1187);
xnor U3167 (N_3167,In_559,In_1388);
nor U3168 (N_3168,In_704,In_1494);
and U3169 (N_3169,In_1261,In_624);
xnor U3170 (N_3170,In_1348,In_37);
or U3171 (N_3171,In_659,In_1134);
and U3172 (N_3172,In_1018,In_603);
and U3173 (N_3173,In_940,In_762);
nor U3174 (N_3174,In_1200,In_332);
and U3175 (N_3175,In_1326,In_227);
xnor U3176 (N_3176,In_1207,In_629);
nor U3177 (N_3177,In_1484,In_1056);
or U3178 (N_3178,In_45,In_1250);
nor U3179 (N_3179,In_1014,In_795);
nor U3180 (N_3180,In_641,In_714);
xnor U3181 (N_3181,In_890,In_729);
and U3182 (N_3182,In_1111,In_742);
nand U3183 (N_3183,In_452,In_1023);
xor U3184 (N_3184,In_1397,In_349);
and U3185 (N_3185,In_1190,In_1119);
and U3186 (N_3186,In_604,In_695);
and U3187 (N_3187,In_121,In_946);
and U3188 (N_3188,In_3,In_415);
nand U3189 (N_3189,In_778,In_1018);
nand U3190 (N_3190,In_1412,In_1141);
xor U3191 (N_3191,In_1347,In_1402);
nand U3192 (N_3192,In_888,In_1153);
nor U3193 (N_3193,In_1046,In_536);
xor U3194 (N_3194,In_586,In_726);
nor U3195 (N_3195,In_433,In_301);
nand U3196 (N_3196,In_758,In_624);
nand U3197 (N_3197,In_1272,In_15);
or U3198 (N_3198,In_36,In_1209);
or U3199 (N_3199,In_109,In_1362);
nor U3200 (N_3200,In_25,In_690);
xor U3201 (N_3201,In_858,In_19);
nor U3202 (N_3202,In_1309,In_860);
nand U3203 (N_3203,In_443,In_1416);
and U3204 (N_3204,In_241,In_1466);
nor U3205 (N_3205,In_1438,In_1003);
xnor U3206 (N_3206,In_1383,In_1148);
and U3207 (N_3207,In_1148,In_1107);
nand U3208 (N_3208,In_1164,In_1242);
and U3209 (N_3209,In_701,In_378);
xor U3210 (N_3210,In_35,In_250);
xnor U3211 (N_3211,In_231,In_191);
and U3212 (N_3212,In_28,In_814);
xnor U3213 (N_3213,In_869,In_1302);
and U3214 (N_3214,In_399,In_589);
or U3215 (N_3215,In_881,In_1456);
or U3216 (N_3216,In_722,In_583);
nor U3217 (N_3217,In_766,In_539);
or U3218 (N_3218,In_294,In_1277);
xnor U3219 (N_3219,In_1296,In_1222);
nand U3220 (N_3220,In_508,In_1253);
xnor U3221 (N_3221,In_1055,In_1292);
nand U3222 (N_3222,In_1076,In_844);
nor U3223 (N_3223,In_718,In_328);
and U3224 (N_3224,In_174,In_227);
and U3225 (N_3225,In_1424,In_28);
or U3226 (N_3226,In_441,In_799);
nor U3227 (N_3227,In_667,In_197);
or U3228 (N_3228,In_783,In_731);
nand U3229 (N_3229,In_855,In_1368);
nor U3230 (N_3230,In_75,In_103);
xor U3231 (N_3231,In_1141,In_236);
xnor U3232 (N_3232,In_501,In_346);
or U3233 (N_3233,In_751,In_1120);
nor U3234 (N_3234,In_197,In_241);
or U3235 (N_3235,In_152,In_515);
or U3236 (N_3236,In_1269,In_156);
nor U3237 (N_3237,In_273,In_318);
nand U3238 (N_3238,In_985,In_94);
or U3239 (N_3239,In_809,In_135);
nor U3240 (N_3240,In_742,In_163);
and U3241 (N_3241,In_354,In_1173);
xnor U3242 (N_3242,In_786,In_1149);
xor U3243 (N_3243,In_1309,In_598);
nand U3244 (N_3244,In_1490,In_953);
and U3245 (N_3245,In_255,In_970);
nor U3246 (N_3246,In_273,In_528);
nor U3247 (N_3247,In_193,In_753);
xor U3248 (N_3248,In_1304,In_1320);
nor U3249 (N_3249,In_574,In_416);
nor U3250 (N_3250,In_217,In_385);
or U3251 (N_3251,In_1496,In_715);
xor U3252 (N_3252,In_533,In_125);
nor U3253 (N_3253,In_18,In_1442);
nand U3254 (N_3254,In_202,In_124);
xor U3255 (N_3255,In_1078,In_1158);
and U3256 (N_3256,In_881,In_504);
and U3257 (N_3257,In_393,In_1153);
nand U3258 (N_3258,In_783,In_378);
xnor U3259 (N_3259,In_396,In_1101);
or U3260 (N_3260,In_1462,In_832);
nor U3261 (N_3261,In_493,In_317);
nor U3262 (N_3262,In_231,In_489);
xnor U3263 (N_3263,In_667,In_1034);
or U3264 (N_3264,In_84,In_469);
nor U3265 (N_3265,In_412,In_1236);
xnor U3266 (N_3266,In_127,In_574);
nor U3267 (N_3267,In_1468,In_498);
xnor U3268 (N_3268,In_1495,In_1277);
nand U3269 (N_3269,In_1309,In_318);
or U3270 (N_3270,In_614,In_510);
xor U3271 (N_3271,In_142,In_382);
or U3272 (N_3272,In_1292,In_1249);
nor U3273 (N_3273,In_1174,In_800);
nor U3274 (N_3274,In_482,In_760);
nand U3275 (N_3275,In_184,In_1212);
or U3276 (N_3276,In_341,In_778);
xnor U3277 (N_3277,In_207,In_141);
xnor U3278 (N_3278,In_361,In_729);
and U3279 (N_3279,In_444,In_1150);
or U3280 (N_3280,In_584,In_396);
or U3281 (N_3281,In_602,In_1313);
nor U3282 (N_3282,In_873,In_965);
and U3283 (N_3283,In_512,In_1469);
and U3284 (N_3284,In_209,In_179);
xnor U3285 (N_3285,In_694,In_1391);
nor U3286 (N_3286,In_777,In_800);
nand U3287 (N_3287,In_475,In_836);
and U3288 (N_3288,In_819,In_903);
xor U3289 (N_3289,In_1466,In_14);
nor U3290 (N_3290,In_816,In_21);
xnor U3291 (N_3291,In_973,In_504);
nand U3292 (N_3292,In_1452,In_1352);
xor U3293 (N_3293,In_1123,In_489);
nor U3294 (N_3294,In_602,In_575);
xnor U3295 (N_3295,In_1368,In_399);
xor U3296 (N_3296,In_449,In_489);
nor U3297 (N_3297,In_1332,In_281);
nand U3298 (N_3298,In_1101,In_1008);
and U3299 (N_3299,In_179,In_1497);
nand U3300 (N_3300,In_997,In_1468);
nand U3301 (N_3301,In_951,In_2);
and U3302 (N_3302,In_951,In_11);
nand U3303 (N_3303,In_503,In_585);
nor U3304 (N_3304,In_218,In_1422);
nand U3305 (N_3305,In_1472,In_985);
nand U3306 (N_3306,In_485,In_510);
xor U3307 (N_3307,In_1266,In_177);
xor U3308 (N_3308,In_94,In_1092);
xnor U3309 (N_3309,In_1322,In_435);
and U3310 (N_3310,In_225,In_601);
nor U3311 (N_3311,In_498,In_385);
nand U3312 (N_3312,In_123,In_372);
and U3313 (N_3313,In_231,In_278);
and U3314 (N_3314,In_730,In_265);
xnor U3315 (N_3315,In_719,In_617);
or U3316 (N_3316,In_311,In_1034);
nor U3317 (N_3317,In_747,In_183);
or U3318 (N_3318,In_1132,In_928);
or U3319 (N_3319,In_1103,In_601);
nor U3320 (N_3320,In_996,In_1251);
nor U3321 (N_3321,In_1222,In_496);
or U3322 (N_3322,In_1286,In_45);
nand U3323 (N_3323,In_627,In_1035);
nand U3324 (N_3324,In_425,In_1123);
xnor U3325 (N_3325,In_802,In_816);
nor U3326 (N_3326,In_921,In_371);
nand U3327 (N_3327,In_272,In_1153);
nand U3328 (N_3328,In_2,In_1229);
and U3329 (N_3329,In_765,In_825);
xor U3330 (N_3330,In_1345,In_940);
nor U3331 (N_3331,In_387,In_1139);
or U3332 (N_3332,In_986,In_466);
nand U3333 (N_3333,In_143,In_256);
nand U3334 (N_3334,In_1385,In_416);
or U3335 (N_3335,In_259,In_828);
or U3336 (N_3336,In_162,In_1070);
nand U3337 (N_3337,In_184,In_475);
xnor U3338 (N_3338,In_964,In_62);
nand U3339 (N_3339,In_781,In_760);
nand U3340 (N_3340,In_1034,In_1083);
nand U3341 (N_3341,In_1441,In_1493);
or U3342 (N_3342,In_1479,In_140);
or U3343 (N_3343,In_965,In_728);
nor U3344 (N_3344,In_864,In_523);
nand U3345 (N_3345,In_1025,In_1359);
or U3346 (N_3346,In_1006,In_1244);
nor U3347 (N_3347,In_419,In_266);
xnor U3348 (N_3348,In_481,In_805);
or U3349 (N_3349,In_21,In_287);
and U3350 (N_3350,In_677,In_1198);
and U3351 (N_3351,In_728,In_1220);
and U3352 (N_3352,In_1355,In_1495);
nand U3353 (N_3353,In_139,In_655);
nor U3354 (N_3354,In_1170,In_335);
and U3355 (N_3355,In_276,In_1351);
nor U3356 (N_3356,In_69,In_600);
or U3357 (N_3357,In_133,In_189);
xnor U3358 (N_3358,In_1243,In_27);
xor U3359 (N_3359,In_221,In_287);
xnor U3360 (N_3360,In_451,In_565);
or U3361 (N_3361,In_157,In_767);
and U3362 (N_3362,In_112,In_962);
and U3363 (N_3363,In_728,In_1072);
xnor U3364 (N_3364,In_1274,In_464);
xnor U3365 (N_3365,In_607,In_1355);
xor U3366 (N_3366,In_1006,In_665);
nor U3367 (N_3367,In_504,In_558);
xnor U3368 (N_3368,In_1378,In_1455);
nand U3369 (N_3369,In_610,In_230);
nor U3370 (N_3370,In_810,In_981);
and U3371 (N_3371,In_1094,In_428);
nand U3372 (N_3372,In_656,In_1016);
nand U3373 (N_3373,In_647,In_222);
xor U3374 (N_3374,In_1496,In_542);
or U3375 (N_3375,In_654,In_1073);
or U3376 (N_3376,In_301,In_1499);
nand U3377 (N_3377,In_767,In_410);
and U3378 (N_3378,In_847,In_1313);
nand U3379 (N_3379,In_1248,In_303);
xor U3380 (N_3380,In_563,In_1100);
xor U3381 (N_3381,In_708,In_857);
nor U3382 (N_3382,In_343,In_1156);
nand U3383 (N_3383,In_756,In_676);
xnor U3384 (N_3384,In_874,In_1041);
and U3385 (N_3385,In_610,In_1298);
and U3386 (N_3386,In_1357,In_1141);
nor U3387 (N_3387,In_1246,In_953);
and U3388 (N_3388,In_327,In_617);
nand U3389 (N_3389,In_1291,In_358);
and U3390 (N_3390,In_358,In_378);
nor U3391 (N_3391,In_1281,In_1027);
xor U3392 (N_3392,In_101,In_308);
nand U3393 (N_3393,In_522,In_842);
nand U3394 (N_3394,In_1131,In_1229);
xnor U3395 (N_3395,In_282,In_505);
xnor U3396 (N_3396,In_637,In_660);
xnor U3397 (N_3397,In_589,In_36);
nand U3398 (N_3398,In_759,In_1117);
nand U3399 (N_3399,In_966,In_1320);
xor U3400 (N_3400,In_456,In_1317);
nand U3401 (N_3401,In_1202,In_1455);
and U3402 (N_3402,In_1102,In_946);
nand U3403 (N_3403,In_731,In_53);
nand U3404 (N_3404,In_1251,In_332);
nand U3405 (N_3405,In_1444,In_1303);
or U3406 (N_3406,In_628,In_832);
and U3407 (N_3407,In_149,In_706);
and U3408 (N_3408,In_578,In_1381);
and U3409 (N_3409,In_1312,In_1488);
and U3410 (N_3410,In_457,In_138);
nand U3411 (N_3411,In_1120,In_367);
nand U3412 (N_3412,In_871,In_244);
nand U3413 (N_3413,In_1046,In_707);
nand U3414 (N_3414,In_763,In_494);
nor U3415 (N_3415,In_138,In_1036);
nor U3416 (N_3416,In_1315,In_1230);
xor U3417 (N_3417,In_486,In_344);
and U3418 (N_3418,In_1274,In_847);
or U3419 (N_3419,In_323,In_1461);
nand U3420 (N_3420,In_694,In_1390);
nor U3421 (N_3421,In_371,In_225);
xor U3422 (N_3422,In_1427,In_96);
or U3423 (N_3423,In_880,In_647);
nand U3424 (N_3424,In_589,In_1440);
or U3425 (N_3425,In_709,In_373);
and U3426 (N_3426,In_611,In_649);
nor U3427 (N_3427,In_1328,In_689);
xor U3428 (N_3428,In_942,In_1433);
xor U3429 (N_3429,In_402,In_286);
nand U3430 (N_3430,In_986,In_327);
nor U3431 (N_3431,In_259,In_1469);
nand U3432 (N_3432,In_815,In_683);
or U3433 (N_3433,In_269,In_1252);
and U3434 (N_3434,In_405,In_657);
nor U3435 (N_3435,In_1211,In_1066);
nand U3436 (N_3436,In_1385,In_79);
and U3437 (N_3437,In_91,In_1085);
and U3438 (N_3438,In_1145,In_788);
or U3439 (N_3439,In_1356,In_359);
nand U3440 (N_3440,In_980,In_938);
nor U3441 (N_3441,In_1074,In_434);
xor U3442 (N_3442,In_1123,In_1416);
nand U3443 (N_3443,In_566,In_1437);
or U3444 (N_3444,In_835,In_594);
and U3445 (N_3445,In_818,In_180);
nor U3446 (N_3446,In_513,In_928);
nand U3447 (N_3447,In_810,In_33);
or U3448 (N_3448,In_992,In_1238);
xor U3449 (N_3449,In_582,In_1343);
or U3450 (N_3450,In_727,In_498);
and U3451 (N_3451,In_154,In_381);
and U3452 (N_3452,In_677,In_207);
nand U3453 (N_3453,In_107,In_542);
nand U3454 (N_3454,In_1382,In_635);
nor U3455 (N_3455,In_1038,In_1295);
or U3456 (N_3456,In_31,In_152);
xnor U3457 (N_3457,In_485,In_337);
or U3458 (N_3458,In_88,In_1044);
nand U3459 (N_3459,In_391,In_140);
nand U3460 (N_3460,In_418,In_78);
xnor U3461 (N_3461,In_1403,In_1041);
nor U3462 (N_3462,In_684,In_816);
or U3463 (N_3463,In_705,In_765);
or U3464 (N_3464,In_596,In_52);
nor U3465 (N_3465,In_1065,In_437);
and U3466 (N_3466,In_979,In_1022);
nor U3467 (N_3467,In_1003,In_1273);
and U3468 (N_3468,In_641,In_982);
and U3469 (N_3469,In_1068,In_1059);
nand U3470 (N_3470,In_126,In_1109);
xor U3471 (N_3471,In_1354,In_478);
or U3472 (N_3472,In_1378,In_225);
and U3473 (N_3473,In_530,In_374);
xnor U3474 (N_3474,In_289,In_1104);
nand U3475 (N_3475,In_958,In_1007);
nand U3476 (N_3476,In_1034,In_326);
and U3477 (N_3477,In_617,In_895);
or U3478 (N_3478,In_903,In_423);
and U3479 (N_3479,In_853,In_103);
nand U3480 (N_3480,In_1033,In_413);
nand U3481 (N_3481,In_263,In_420);
nand U3482 (N_3482,In_1274,In_119);
or U3483 (N_3483,In_1409,In_918);
xnor U3484 (N_3484,In_919,In_848);
nand U3485 (N_3485,In_808,In_1195);
and U3486 (N_3486,In_1191,In_893);
nor U3487 (N_3487,In_1017,In_1076);
xnor U3488 (N_3488,In_1476,In_132);
and U3489 (N_3489,In_1093,In_670);
xor U3490 (N_3490,In_1398,In_344);
nand U3491 (N_3491,In_1250,In_221);
nor U3492 (N_3492,In_70,In_10);
and U3493 (N_3493,In_341,In_836);
nor U3494 (N_3494,In_509,In_116);
or U3495 (N_3495,In_1152,In_1153);
xnor U3496 (N_3496,In_1488,In_1480);
nand U3497 (N_3497,In_282,In_261);
or U3498 (N_3498,In_415,In_599);
nor U3499 (N_3499,In_947,In_1431);
nor U3500 (N_3500,In_705,In_1032);
xor U3501 (N_3501,In_431,In_1010);
nor U3502 (N_3502,In_1026,In_1147);
nor U3503 (N_3503,In_981,In_361);
nand U3504 (N_3504,In_532,In_319);
xnor U3505 (N_3505,In_446,In_821);
or U3506 (N_3506,In_661,In_329);
xnor U3507 (N_3507,In_418,In_556);
nand U3508 (N_3508,In_241,In_44);
and U3509 (N_3509,In_95,In_822);
and U3510 (N_3510,In_710,In_368);
and U3511 (N_3511,In_1343,In_1073);
nor U3512 (N_3512,In_1340,In_176);
and U3513 (N_3513,In_392,In_169);
and U3514 (N_3514,In_1388,In_861);
nand U3515 (N_3515,In_1254,In_308);
nand U3516 (N_3516,In_6,In_897);
nor U3517 (N_3517,In_1198,In_547);
nor U3518 (N_3518,In_435,In_398);
or U3519 (N_3519,In_1117,In_308);
xnor U3520 (N_3520,In_1487,In_1007);
and U3521 (N_3521,In_167,In_319);
nand U3522 (N_3522,In_223,In_870);
nor U3523 (N_3523,In_20,In_1259);
nor U3524 (N_3524,In_130,In_1025);
or U3525 (N_3525,In_226,In_582);
nor U3526 (N_3526,In_658,In_253);
and U3527 (N_3527,In_1295,In_1266);
nand U3528 (N_3528,In_142,In_36);
nand U3529 (N_3529,In_1472,In_540);
nand U3530 (N_3530,In_697,In_1325);
or U3531 (N_3531,In_763,In_42);
and U3532 (N_3532,In_668,In_1487);
xnor U3533 (N_3533,In_1494,In_26);
nand U3534 (N_3534,In_247,In_1097);
nor U3535 (N_3535,In_446,In_838);
xor U3536 (N_3536,In_132,In_1216);
and U3537 (N_3537,In_1401,In_268);
xnor U3538 (N_3538,In_210,In_246);
and U3539 (N_3539,In_1094,In_759);
and U3540 (N_3540,In_130,In_1327);
or U3541 (N_3541,In_1221,In_1005);
nor U3542 (N_3542,In_904,In_805);
nand U3543 (N_3543,In_1234,In_1022);
nor U3544 (N_3544,In_580,In_1160);
xor U3545 (N_3545,In_1053,In_684);
and U3546 (N_3546,In_646,In_230);
and U3547 (N_3547,In_755,In_871);
nand U3548 (N_3548,In_808,In_1445);
or U3549 (N_3549,In_1476,In_1178);
nor U3550 (N_3550,In_515,In_995);
nand U3551 (N_3551,In_107,In_705);
and U3552 (N_3552,In_751,In_165);
nand U3553 (N_3553,In_1495,In_313);
and U3554 (N_3554,In_123,In_1089);
or U3555 (N_3555,In_1194,In_200);
or U3556 (N_3556,In_19,In_1137);
nor U3557 (N_3557,In_291,In_1376);
xor U3558 (N_3558,In_18,In_1363);
nand U3559 (N_3559,In_1123,In_1285);
and U3560 (N_3560,In_39,In_261);
nand U3561 (N_3561,In_627,In_263);
nor U3562 (N_3562,In_13,In_1040);
and U3563 (N_3563,In_842,In_773);
or U3564 (N_3564,In_601,In_881);
nand U3565 (N_3565,In_658,In_1152);
and U3566 (N_3566,In_1222,In_585);
xnor U3567 (N_3567,In_732,In_619);
nand U3568 (N_3568,In_1302,In_128);
xnor U3569 (N_3569,In_300,In_182);
and U3570 (N_3570,In_18,In_1381);
xor U3571 (N_3571,In_478,In_697);
and U3572 (N_3572,In_632,In_1196);
xor U3573 (N_3573,In_432,In_548);
nor U3574 (N_3574,In_692,In_986);
and U3575 (N_3575,In_236,In_189);
nand U3576 (N_3576,In_1319,In_372);
nor U3577 (N_3577,In_32,In_85);
nand U3578 (N_3578,In_1360,In_930);
nor U3579 (N_3579,In_605,In_979);
xnor U3580 (N_3580,In_288,In_190);
and U3581 (N_3581,In_300,In_1186);
nand U3582 (N_3582,In_1185,In_1406);
xnor U3583 (N_3583,In_1241,In_1083);
xnor U3584 (N_3584,In_295,In_179);
xor U3585 (N_3585,In_926,In_28);
nor U3586 (N_3586,In_193,In_948);
nand U3587 (N_3587,In_437,In_551);
and U3588 (N_3588,In_1378,In_1076);
nand U3589 (N_3589,In_1023,In_1241);
nor U3590 (N_3590,In_1023,In_1253);
and U3591 (N_3591,In_1052,In_492);
xor U3592 (N_3592,In_452,In_1343);
nor U3593 (N_3593,In_166,In_70);
or U3594 (N_3594,In_77,In_830);
or U3595 (N_3595,In_501,In_1349);
and U3596 (N_3596,In_157,In_695);
nor U3597 (N_3597,In_1174,In_303);
nor U3598 (N_3598,In_1469,In_1331);
nor U3599 (N_3599,In_334,In_8);
nor U3600 (N_3600,In_760,In_156);
nand U3601 (N_3601,In_272,In_168);
nand U3602 (N_3602,In_89,In_907);
or U3603 (N_3603,In_704,In_550);
or U3604 (N_3604,In_919,In_861);
or U3605 (N_3605,In_971,In_1231);
or U3606 (N_3606,In_993,In_484);
and U3607 (N_3607,In_1063,In_1049);
nor U3608 (N_3608,In_798,In_1018);
xor U3609 (N_3609,In_285,In_286);
or U3610 (N_3610,In_1234,In_125);
and U3611 (N_3611,In_1145,In_1230);
xor U3612 (N_3612,In_654,In_1476);
or U3613 (N_3613,In_1316,In_578);
xnor U3614 (N_3614,In_225,In_881);
and U3615 (N_3615,In_554,In_789);
nor U3616 (N_3616,In_622,In_222);
nor U3617 (N_3617,In_544,In_1229);
or U3618 (N_3618,In_102,In_465);
xnor U3619 (N_3619,In_807,In_174);
xnor U3620 (N_3620,In_24,In_1203);
or U3621 (N_3621,In_561,In_899);
nand U3622 (N_3622,In_1028,In_600);
nor U3623 (N_3623,In_986,In_1403);
or U3624 (N_3624,In_548,In_787);
or U3625 (N_3625,In_524,In_1186);
and U3626 (N_3626,In_872,In_974);
and U3627 (N_3627,In_808,In_853);
or U3628 (N_3628,In_1276,In_148);
nand U3629 (N_3629,In_277,In_592);
or U3630 (N_3630,In_35,In_552);
xnor U3631 (N_3631,In_55,In_1400);
xnor U3632 (N_3632,In_1337,In_581);
nor U3633 (N_3633,In_982,In_1465);
or U3634 (N_3634,In_271,In_406);
or U3635 (N_3635,In_1324,In_345);
xor U3636 (N_3636,In_26,In_1213);
xnor U3637 (N_3637,In_1216,In_574);
nor U3638 (N_3638,In_1130,In_1325);
and U3639 (N_3639,In_510,In_1490);
or U3640 (N_3640,In_425,In_119);
nand U3641 (N_3641,In_959,In_1295);
nor U3642 (N_3642,In_1150,In_339);
and U3643 (N_3643,In_1461,In_1336);
nand U3644 (N_3644,In_331,In_716);
xnor U3645 (N_3645,In_1362,In_1400);
and U3646 (N_3646,In_294,In_477);
or U3647 (N_3647,In_553,In_1267);
nand U3648 (N_3648,In_1496,In_62);
nor U3649 (N_3649,In_276,In_573);
nand U3650 (N_3650,In_1141,In_334);
nor U3651 (N_3651,In_459,In_370);
and U3652 (N_3652,In_611,In_890);
nor U3653 (N_3653,In_1172,In_664);
xor U3654 (N_3654,In_701,In_890);
nor U3655 (N_3655,In_509,In_1064);
nand U3656 (N_3656,In_833,In_296);
or U3657 (N_3657,In_1065,In_399);
xor U3658 (N_3658,In_1454,In_504);
xnor U3659 (N_3659,In_205,In_730);
nand U3660 (N_3660,In_1069,In_868);
xor U3661 (N_3661,In_1289,In_266);
nand U3662 (N_3662,In_197,In_472);
xor U3663 (N_3663,In_427,In_404);
and U3664 (N_3664,In_1246,In_468);
xor U3665 (N_3665,In_996,In_1099);
and U3666 (N_3666,In_502,In_1311);
nand U3667 (N_3667,In_388,In_1129);
nand U3668 (N_3668,In_928,In_168);
nand U3669 (N_3669,In_1394,In_923);
xnor U3670 (N_3670,In_403,In_107);
xnor U3671 (N_3671,In_909,In_398);
or U3672 (N_3672,In_701,In_1395);
xnor U3673 (N_3673,In_76,In_293);
or U3674 (N_3674,In_1284,In_894);
xor U3675 (N_3675,In_1449,In_136);
nor U3676 (N_3676,In_878,In_977);
xnor U3677 (N_3677,In_178,In_1472);
or U3678 (N_3678,In_1435,In_1018);
or U3679 (N_3679,In_56,In_1329);
nand U3680 (N_3680,In_611,In_387);
or U3681 (N_3681,In_1129,In_358);
and U3682 (N_3682,In_66,In_998);
nand U3683 (N_3683,In_416,In_1382);
xnor U3684 (N_3684,In_33,In_456);
or U3685 (N_3685,In_216,In_556);
xnor U3686 (N_3686,In_750,In_491);
nand U3687 (N_3687,In_334,In_1206);
nand U3688 (N_3688,In_390,In_1212);
nor U3689 (N_3689,In_1115,In_564);
and U3690 (N_3690,In_1354,In_1022);
and U3691 (N_3691,In_1424,In_412);
nor U3692 (N_3692,In_1426,In_199);
xor U3693 (N_3693,In_785,In_1331);
xnor U3694 (N_3694,In_633,In_274);
nor U3695 (N_3695,In_319,In_68);
nand U3696 (N_3696,In_930,In_508);
nor U3697 (N_3697,In_1101,In_97);
xor U3698 (N_3698,In_116,In_1273);
xor U3699 (N_3699,In_300,In_330);
and U3700 (N_3700,In_1357,In_434);
nand U3701 (N_3701,In_160,In_29);
and U3702 (N_3702,In_206,In_538);
or U3703 (N_3703,In_133,In_512);
or U3704 (N_3704,In_775,In_783);
or U3705 (N_3705,In_702,In_1295);
or U3706 (N_3706,In_477,In_666);
and U3707 (N_3707,In_1284,In_920);
nand U3708 (N_3708,In_902,In_1365);
nor U3709 (N_3709,In_655,In_257);
xor U3710 (N_3710,In_313,In_1094);
or U3711 (N_3711,In_736,In_1379);
nand U3712 (N_3712,In_1472,In_147);
xor U3713 (N_3713,In_161,In_661);
nand U3714 (N_3714,In_370,In_1245);
and U3715 (N_3715,In_1117,In_864);
nand U3716 (N_3716,In_1024,In_921);
nand U3717 (N_3717,In_127,In_247);
xor U3718 (N_3718,In_619,In_299);
xnor U3719 (N_3719,In_533,In_523);
xnor U3720 (N_3720,In_316,In_82);
nand U3721 (N_3721,In_1428,In_1191);
or U3722 (N_3722,In_303,In_3);
nand U3723 (N_3723,In_1479,In_1026);
or U3724 (N_3724,In_1263,In_644);
nor U3725 (N_3725,In_599,In_661);
or U3726 (N_3726,In_877,In_1079);
or U3727 (N_3727,In_746,In_525);
and U3728 (N_3728,In_473,In_1435);
or U3729 (N_3729,In_1120,In_613);
nor U3730 (N_3730,In_1466,In_813);
or U3731 (N_3731,In_1411,In_1281);
or U3732 (N_3732,In_188,In_24);
nand U3733 (N_3733,In_1302,In_265);
nand U3734 (N_3734,In_398,In_1087);
nand U3735 (N_3735,In_1080,In_1373);
or U3736 (N_3736,In_915,In_1203);
nand U3737 (N_3737,In_188,In_158);
xnor U3738 (N_3738,In_1063,In_1385);
or U3739 (N_3739,In_87,In_574);
xor U3740 (N_3740,In_1478,In_1066);
or U3741 (N_3741,In_1037,In_490);
and U3742 (N_3742,In_276,In_1375);
nand U3743 (N_3743,In_1187,In_1180);
nand U3744 (N_3744,In_1114,In_697);
nor U3745 (N_3745,In_150,In_1124);
xnor U3746 (N_3746,In_136,In_578);
xor U3747 (N_3747,In_1340,In_1385);
nor U3748 (N_3748,In_741,In_1123);
and U3749 (N_3749,In_346,In_1130);
or U3750 (N_3750,In_1361,In_1177);
xnor U3751 (N_3751,In_230,In_451);
and U3752 (N_3752,In_741,In_687);
and U3753 (N_3753,In_1224,In_109);
nand U3754 (N_3754,In_1127,In_358);
nand U3755 (N_3755,In_502,In_1471);
and U3756 (N_3756,In_446,In_760);
and U3757 (N_3757,In_853,In_594);
nor U3758 (N_3758,In_387,In_1130);
nor U3759 (N_3759,In_463,In_13);
nor U3760 (N_3760,In_1271,In_1236);
xor U3761 (N_3761,In_849,In_253);
and U3762 (N_3762,In_1377,In_552);
and U3763 (N_3763,In_1271,In_1110);
and U3764 (N_3764,In_398,In_1059);
nor U3765 (N_3765,In_609,In_503);
nor U3766 (N_3766,In_578,In_282);
nor U3767 (N_3767,In_406,In_125);
or U3768 (N_3768,In_1037,In_1443);
or U3769 (N_3769,In_705,In_958);
nand U3770 (N_3770,In_143,In_1176);
or U3771 (N_3771,In_1402,In_1237);
xor U3772 (N_3772,In_236,In_1013);
or U3773 (N_3773,In_1075,In_1323);
xnor U3774 (N_3774,In_203,In_896);
nand U3775 (N_3775,In_481,In_630);
xor U3776 (N_3776,In_73,In_860);
and U3777 (N_3777,In_1453,In_84);
nor U3778 (N_3778,In_1037,In_516);
or U3779 (N_3779,In_1411,In_52);
or U3780 (N_3780,In_230,In_1175);
xnor U3781 (N_3781,In_1031,In_1387);
and U3782 (N_3782,In_326,In_1311);
nor U3783 (N_3783,In_1126,In_1100);
and U3784 (N_3784,In_1002,In_560);
nor U3785 (N_3785,In_601,In_1005);
nand U3786 (N_3786,In_754,In_412);
xor U3787 (N_3787,In_888,In_281);
xnor U3788 (N_3788,In_1093,In_238);
or U3789 (N_3789,In_988,In_393);
or U3790 (N_3790,In_424,In_987);
or U3791 (N_3791,In_258,In_1291);
nor U3792 (N_3792,In_86,In_710);
nor U3793 (N_3793,In_972,In_1318);
xor U3794 (N_3794,In_1193,In_840);
or U3795 (N_3795,In_181,In_1345);
xnor U3796 (N_3796,In_533,In_852);
and U3797 (N_3797,In_267,In_75);
nor U3798 (N_3798,In_1327,In_1028);
xnor U3799 (N_3799,In_64,In_283);
nand U3800 (N_3800,In_1315,In_894);
nand U3801 (N_3801,In_1032,In_1413);
nor U3802 (N_3802,In_1381,In_1267);
nand U3803 (N_3803,In_1119,In_1017);
nor U3804 (N_3804,In_218,In_1327);
nor U3805 (N_3805,In_880,In_998);
or U3806 (N_3806,In_1236,In_645);
nand U3807 (N_3807,In_382,In_968);
nor U3808 (N_3808,In_155,In_1366);
xor U3809 (N_3809,In_214,In_387);
or U3810 (N_3810,In_398,In_899);
nor U3811 (N_3811,In_309,In_930);
and U3812 (N_3812,In_698,In_44);
nand U3813 (N_3813,In_312,In_17);
nand U3814 (N_3814,In_1068,In_1193);
nand U3815 (N_3815,In_233,In_684);
or U3816 (N_3816,In_1327,In_1216);
nor U3817 (N_3817,In_1278,In_749);
nand U3818 (N_3818,In_1479,In_360);
or U3819 (N_3819,In_1290,In_1251);
nand U3820 (N_3820,In_747,In_514);
nand U3821 (N_3821,In_9,In_1166);
nand U3822 (N_3822,In_879,In_447);
xor U3823 (N_3823,In_990,In_1357);
nand U3824 (N_3824,In_1442,In_457);
nor U3825 (N_3825,In_464,In_562);
and U3826 (N_3826,In_1248,In_1137);
xnor U3827 (N_3827,In_143,In_1154);
nand U3828 (N_3828,In_702,In_1023);
and U3829 (N_3829,In_1036,In_691);
or U3830 (N_3830,In_1314,In_166);
nor U3831 (N_3831,In_1195,In_823);
nand U3832 (N_3832,In_77,In_1430);
nor U3833 (N_3833,In_726,In_646);
xnor U3834 (N_3834,In_166,In_1260);
xnor U3835 (N_3835,In_580,In_947);
and U3836 (N_3836,In_557,In_1437);
and U3837 (N_3837,In_276,In_1089);
xor U3838 (N_3838,In_103,In_1025);
nor U3839 (N_3839,In_485,In_81);
nand U3840 (N_3840,In_634,In_645);
xnor U3841 (N_3841,In_553,In_789);
and U3842 (N_3842,In_1088,In_966);
or U3843 (N_3843,In_635,In_1048);
and U3844 (N_3844,In_529,In_911);
xor U3845 (N_3845,In_218,In_563);
nor U3846 (N_3846,In_83,In_1212);
and U3847 (N_3847,In_1469,In_541);
or U3848 (N_3848,In_700,In_285);
and U3849 (N_3849,In_826,In_772);
xor U3850 (N_3850,In_1454,In_820);
xnor U3851 (N_3851,In_549,In_51);
nor U3852 (N_3852,In_1153,In_637);
nand U3853 (N_3853,In_177,In_498);
xor U3854 (N_3854,In_37,In_1109);
xor U3855 (N_3855,In_1308,In_1064);
nor U3856 (N_3856,In_1074,In_856);
or U3857 (N_3857,In_1380,In_339);
nand U3858 (N_3858,In_1386,In_862);
xor U3859 (N_3859,In_231,In_764);
and U3860 (N_3860,In_1273,In_42);
and U3861 (N_3861,In_995,In_1161);
nand U3862 (N_3862,In_1472,In_610);
nor U3863 (N_3863,In_227,In_375);
or U3864 (N_3864,In_270,In_304);
or U3865 (N_3865,In_1396,In_1419);
xnor U3866 (N_3866,In_307,In_116);
and U3867 (N_3867,In_1074,In_1290);
xnor U3868 (N_3868,In_1150,In_586);
nor U3869 (N_3869,In_1200,In_121);
nor U3870 (N_3870,In_738,In_1161);
nor U3871 (N_3871,In_312,In_1302);
and U3872 (N_3872,In_688,In_865);
or U3873 (N_3873,In_1345,In_180);
or U3874 (N_3874,In_366,In_841);
and U3875 (N_3875,In_1174,In_850);
or U3876 (N_3876,In_64,In_698);
or U3877 (N_3877,In_548,In_156);
or U3878 (N_3878,In_1098,In_1317);
and U3879 (N_3879,In_431,In_1184);
xor U3880 (N_3880,In_288,In_59);
nor U3881 (N_3881,In_316,In_1410);
nand U3882 (N_3882,In_1086,In_1074);
xor U3883 (N_3883,In_121,In_1164);
nor U3884 (N_3884,In_473,In_100);
nand U3885 (N_3885,In_901,In_399);
and U3886 (N_3886,In_1003,In_342);
nor U3887 (N_3887,In_730,In_122);
and U3888 (N_3888,In_131,In_564);
nor U3889 (N_3889,In_247,In_1359);
or U3890 (N_3890,In_912,In_762);
or U3891 (N_3891,In_154,In_915);
or U3892 (N_3892,In_354,In_582);
nand U3893 (N_3893,In_632,In_1319);
nor U3894 (N_3894,In_588,In_1230);
and U3895 (N_3895,In_403,In_1296);
and U3896 (N_3896,In_1394,In_329);
and U3897 (N_3897,In_1216,In_1480);
and U3898 (N_3898,In_359,In_879);
or U3899 (N_3899,In_174,In_329);
nand U3900 (N_3900,In_903,In_1498);
nor U3901 (N_3901,In_557,In_812);
nand U3902 (N_3902,In_1199,In_856);
xnor U3903 (N_3903,In_1462,In_504);
xor U3904 (N_3904,In_1476,In_1201);
nand U3905 (N_3905,In_90,In_1069);
and U3906 (N_3906,In_1148,In_619);
and U3907 (N_3907,In_664,In_317);
or U3908 (N_3908,In_752,In_1360);
or U3909 (N_3909,In_1260,In_548);
nor U3910 (N_3910,In_911,In_231);
nand U3911 (N_3911,In_541,In_1177);
nor U3912 (N_3912,In_138,In_1143);
xnor U3913 (N_3913,In_714,In_852);
nor U3914 (N_3914,In_99,In_857);
or U3915 (N_3915,In_133,In_150);
or U3916 (N_3916,In_306,In_1226);
and U3917 (N_3917,In_1472,In_950);
nand U3918 (N_3918,In_667,In_311);
or U3919 (N_3919,In_502,In_1383);
xnor U3920 (N_3920,In_130,In_1257);
and U3921 (N_3921,In_1337,In_815);
nor U3922 (N_3922,In_1329,In_966);
and U3923 (N_3923,In_416,In_284);
and U3924 (N_3924,In_54,In_1463);
and U3925 (N_3925,In_273,In_1251);
xnor U3926 (N_3926,In_959,In_657);
nor U3927 (N_3927,In_557,In_956);
and U3928 (N_3928,In_257,In_1495);
nand U3929 (N_3929,In_487,In_426);
and U3930 (N_3930,In_1216,In_1137);
nand U3931 (N_3931,In_1193,In_629);
nand U3932 (N_3932,In_920,In_1183);
and U3933 (N_3933,In_143,In_278);
or U3934 (N_3934,In_753,In_673);
nand U3935 (N_3935,In_1224,In_314);
and U3936 (N_3936,In_1447,In_753);
or U3937 (N_3937,In_1250,In_1237);
nor U3938 (N_3938,In_200,In_287);
nor U3939 (N_3939,In_122,In_119);
or U3940 (N_3940,In_1186,In_478);
and U3941 (N_3941,In_1250,In_914);
or U3942 (N_3942,In_1343,In_1196);
nand U3943 (N_3943,In_1278,In_162);
or U3944 (N_3944,In_512,In_105);
nand U3945 (N_3945,In_859,In_433);
xnor U3946 (N_3946,In_796,In_966);
and U3947 (N_3947,In_1033,In_864);
xor U3948 (N_3948,In_160,In_56);
or U3949 (N_3949,In_573,In_6);
or U3950 (N_3950,In_900,In_1036);
nand U3951 (N_3951,In_724,In_766);
nand U3952 (N_3952,In_676,In_752);
xnor U3953 (N_3953,In_525,In_428);
xor U3954 (N_3954,In_106,In_378);
xnor U3955 (N_3955,In_240,In_200);
nand U3956 (N_3956,In_1023,In_1357);
xor U3957 (N_3957,In_898,In_1255);
and U3958 (N_3958,In_291,In_1374);
or U3959 (N_3959,In_1426,In_1339);
and U3960 (N_3960,In_991,In_570);
nand U3961 (N_3961,In_1471,In_898);
xor U3962 (N_3962,In_884,In_136);
xor U3963 (N_3963,In_136,In_657);
xnor U3964 (N_3964,In_133,In_995);
and U3965 (N_3965,In_1130,In_206);
xnor U3966 (N_3966,In_1042,In_521);
and U3967 (N_3967,In_1118,In_612);
nand U3968 (N_3968,In_289,In_192);
nor U3969 (N_3969,In_1172,In_536);
nor U3970 (N_3970,In_1154,In_581);
nor U3971 (N_3971,In_810,In_615);
nor U3972 (N_3972,In_186,In_1415);
nand U3973 (N_3973,In_1219,In_624);
nand U3974 (N_3974,In_242,In_48);
nand U3975 (N_3975,In_1054,In_453);
or U3976 (N_3976,In_386,In_144);
or U3977 (N_3977,In_1038,In_1416);
and U3978 (N_3978,In_403,In_915);
xnor U3979 (N_3979,In_1065,In_562);
or U3980 (N_3980,In_1496,In_835);
xnor U3981 (N_3981,In_903,In_1258);
xnor U3982 (N_3982,In_1325,In_1197);
nor U3983 (N_3983,In_1278,In_977);
or U3984 (N_3984,In_863,In_502);
and U3985 (N_3985,In_398,In_835);
nor U3986 (N_3986,In_237,In_1498);
nor U3987 (N_3987,In_1423,In_833);
or U3988 (N_3988,In_1303,In_13);
xor U3989 (N_3989,In_748,In_302);
nand U3990 (N_3990,In_1437,In_977);
or U3991 (N_3991,In_610,In_1151);
and U3992 (N_3992,In_444,In_606);
nand U3993 (N_3993,In_45,In_1055);
nand U3994 (N_3994,In_1343,In_656);
xor U3995 (N_3995,In_7,In_625);
xnor U3996 (N_3996,In_1406,In_487);
and U3997 (N_3997,In_1119,In_335);
and U3998 (N_3998,In_617,In_1291);
and U3999 (N_3999,In_367,In_1462);
nor U4000 (N_4000,In_990,In_658);
or U4001 (N_4001,In_171,In_368);
nor U4002 (N_4002,In_547,In_178);
nor U4003 (N_4003,In_397,In_600);
nand U4004 (N_4004,In_1138,In_1026);
or U4005 (N_4005,In_503,In_174);
and U4006 (N_4006,In_717,In_179);
nor U4007 (N_4007,In_191,In_627);
or U4008 (N_4008,In_78,In_44);
nor U4009 (N_4009,In_1403,In_945);
or U4010 (N_4010,In_957,In_156);
nand U4011 (N_4011,In_924,In_899);
nor U4012 (N_4012,In_33,In_219);
or U4013 (N_4013,In_1289,In_1369);
nand U4014 (N_4014,In_1348,In_1379);
nor U4015 (N_4015,In_626,In_1470);
or U4016 (N_4016,In_891,In_1189);
nand U4017 (N_4017,In_679,In_335);
or U4018 (N_4018,In_709,In_202);
or U4019 (N_4019,In_1381,In_849);
nor U4020 (N_4020,In_828,In_1404);
nor U4021 (N_4021,In_1007,In_691);
xor U4022 (N_4022,In_696,In_1349);
xnor U4023 (N_4023,In_940,In_1468);
and U4024 (N_4024,In_251,In_1451);
nor U4025 (N_4025,In_519,In_1294);
nand U4026 (N_4026,In_51,In_1305);
or U4027 (N_4027,In_641,In_136);
nand U4028 (N_4028,In_878,In_1257);
nor U4029 (N_4029,In_52,In_1433);
xor U4030 (N_4030,In_106,In_479);
nand U4031 (N_4031,In_982,In_865);
nor U4032 (N_4032,In_846,In_1456);
or U4033 (N_4033,In_685,In_1425);
xor U4034 (N_4034,In_318,In_14);
xnor U4035 (N_4035,In_809,In_153);
nor U4036 (N_4036,In_1177,In_814);
or U4037 (N_4037,In_1076,In_1237);
and U4038 (N_4038,In_146,In_1417);
nor U4039 (N_4039,In_418,In_464);
or U4040 (N_4040,In_70,In_280);
or U4041 (N_4041,In_750,In_464);
nor U4042 (N_4042,In_968,In_1124);
or U4043 (N_4043,In_1155,In_187);
nand U4044 (N_4044,In_260,In_1312);
and U4045 (N_4045,In_516,In_691);
or U4046 (N_4046,In_171,In_1255);
nand U4047 (N_4047,In_1491,In_719);
nand U4048 (N_4048,In_542,In_8);
nor U4049 (N_4049,In_1480,In_804);
nand U4050 (N_4050,In_802,In_1283);
xor U4051 (N_4051,In_1489,In_1216);
or U4052 (N_4052,In_422,In_904);
nand U4053 (N_4053,In_1441,In_710);
nand U4054 (N_4054,In_1382,In_663);
and U4055 (N_4055,In_888,In_135);
or U4056 (N_4056,In_394,In_1152);
xnor U4057 (N_4057,In_916,In_655);
and U4058 (N_4058,In_117,In_52);
nand U4059 (N_4059,In_930,In_1269);
xor U4060 (N_4060,In_137,In_899);
nand U4061 (N_4061,In_63,In_126);
or U4062 (N_4062,In_177,In_518);
xor U4063 (N_4063,In_1409,In_911);
and U4064 (N_4064,In_1280,In_224);
nor U4065 (N_4065,In_1419,In_1079);
or U4066 (N_4066,In_373,In_1427);
or U4067 (N_4067,In_1066,In_1162);
and U4068 (N_4068,In_328,In_724);
nand U4069 (N_4069,In_1434,In_460);
or U4070 (N_4070,In_574,In_440);
nand U4071 (N_4071,In_85,In_718);
and U4072 (N_4072,In_108,In_271);
xnor U4073 (N_4073,In_1251,In_59);
or U4074 (N_4074,In_723,In_63);
xnor U4075 (N_4075,In_952,In_492);
and U4076 (N_4076,In_435,In_224);
and U4077 (N_4077,In_1263,In_451);
or U4078 (N_4078,In_531,In_279);
nor U4079 (N_4079,In_194,In_1040);
or U4080 (N_4080,In_110,In_318);
or U4081 (N_4081,In_841,In_1473);
nor U4082 (N_4082,In_623,In_1288);
xor U4083 (N_4083,In_664,In_989);
and U4084 (N_4084,In_308,In_480);
xnor U4085 (N_4085,In_559,In_1171);
or U4086 (N_4086,In_1029,In_356);
nor U4087 (N_4087,In_564,In_48);
and U4088 (N_4088,In_1027,In_507);
and U4089 (N_4089,In_1455,In_1352);
and U4090 (N_4090,In_964,In_132);
nor U4091 (N_4091,In_438,In_626);
and U4092 (N_4092,In_117,In_315);
and U4093 (N_4093,In_1427,In_691);
nand U4094 (N_4094,In_473,In_680);
and U4095 (N_4095,In_1235,In_764);
nor U4096 (N_4096,In_192,In_428);
and U4097 (N_4097,In_198,In_1483);
and U4098 (N_4098,In_857,In_910);
nor U4099 (N_4099,In_1198,In_201);
nand U4100 (N_4100,In_1224,In_1175);
xnor U4101 (N_4101,In_700,In_381);
nor U4102 (N_4102,In_426,In_606);
or U4103 (N_4103,In_1390,In_295);
nand U4104 (N_4104,In_805,In_518);
and U4105 (N_4105,In_1431,In_71);
nand U4106 (N_4106,In_171,In_997);
or U4107 (N_4107,In_55,In_615);
or U4108 (N_4108,In_1478,In_859);
nand U4109 (N_4109,In_285,In_770);
nor U4110 (N_4110,In_1166,In_1306);
or U4111 (N_4111,In_1297,In_1469);
and U4112 (N_4112,In_665,In_528);
nand U4113 (N_4113,In_1286,In_1142);
nor U4114 (N_4114,In_1287,In_684);
nor U4115 (N_4115,In_612,In_616);
or U4116 (N_4116,In_617,In_1200);
xor U4117 (N_4117,In_1021,In_554);
xor U4118 (N_4118,In_1363,In_1142);
nor U4119 (N_4119,In_1417,In_1405);
or U4120 (N_4120,In_1482,In_725);
or U4121 (N_4121,In_343,In_360);
and U4122 (N_4122,In_131,In_1288);
or U4123 (N_4123,In_1292,In_56);
or U4124 (N_4124,In_564,In_1344);
or U4125 (N_4125,In_1236,In_914);
nor U4126 (N_4126,In_1077,In_1352);
nand U4127 (N_4127,In_310,In_835);
or U4128 (N_4128,In_90,In_1123);
xor U4129 (N_4129,In_282,In_1289);
or U4130 (N_4130,In_1465,In_70);
xor U4131 (N_4131,In_516,In_724);
and U4132 (N_4132,In_1208,In_128);
nand U4133 (N_4133,In_1491,In_806);
or U4134 (N_4134,In_761,In_890);
xor U4135 (N_4135,In_820,In_556);
and U4136 (N_4136,In_1295,In_648);
nand U4137 (N_4137,In_1154,In_1014);
nor U4138 (N_4138,In_892,In_295);
and U4139 (N_4139,In_772,In_1087);
xnor U4140 (N_4140,In_278,In_320);
nor U4141 (N_4141,In_1232,In_248);
nand U4142 (N_4142,In_784,In_315);
xnor U4143 (N_4143,In_1080,In_422);
nand U4144 (N_4144,In_808,In_1420);
or U4145 (N_4145,In_1073,In_647);
nor U4146 (N_4146,In_811,In_384);
xnor U4147 (N_4147,In_499,In_120);
or U4148 (N_4148,In_1080,In_309);
nor U4149 (N_4149,In_626,In_145);
or U4150 (N_4150,In_1305,In_212);
nand U4151 (N_4151,In_158,In_29);
nor U4152 (N_4152,In_871,In_840);
or U4153 (N_4153,In_775,In_631);
nor U4154 (N_4154,In_235,In_1489);
or U4155 (N_4155,In_590,In_242);
and U4156 (N_4156,In_1407,In_1366);
nor U4157 (N_4157,In_996,In_390);
nor U4158 (N_4158,In_990,In_937);
or U4159 (N_4159,In_576,In_836);
and U4160 (N_4160,In_1240,In_799);
xnor U4161 (N_4161,In_15,In_36);
or U4162 (N_4162,In_108,In_1286);
nand U4163 (N_4163,In_833,In_576);
nand U4164 (N_4164,In_835,In_863);
or U4165 (N_4165,In_120,In_1382);
and U4166 (N_4166,In_297,In_696);
nor U4167 (N_4167,In_25,In_531);
nor U4168 (N_4168,In_1315,In_1070);
xnor U4169 (N_4169,In_166,In_1339);
xnor U4170 (N_4170,In_589,In_54);
xor U4171 (N_4171,In_766,In_136);
nand U4172 (N_4172,In_66,In_1416);
nand U4173 (N_4173,In_870,In_843);
and U4174 (N_4174,In_676,In_877);
nor U4175 (N_4175,In_1319,In_528);
nand U4176 (N_4176,In_1338,In_726);
nor U4177 (N_4177,In_271,In_1288);
or U4178 (N_4178,In_1313,In_179);
and U4179 (N_4179,In_248,In_434);
xor U4180 (N_4180,In_146,In_333);
nand U4181 (N_4181,In_889,In_394);
nor U4182 (N_4182,In_989,In_632);
nor U4183 (N_4183,In_1332,In_1477);
nand U4184 (N_4184,In_675,In_655);
and U4185 (N_4185,In_316,In_669);
nor U4186 (N_4186,In_1315,In_238);
and U4187 (N_4187,In_163,In_1038);
or U4188 (N_4188,In_1119,In_459);
nand U4189 (N_4189,In_1209,In_204);
nor U4190 (N_4190,In_239,In_1003);
or U4191 (N_4191,In_661,In_1214);
nand U4192 (N_4192,In_1295,In_113);
xnor U4193 (N_4193,In_1166,In_1064);
nand U4194 (N_4194,In_979,In_1382);
nand U4195 (N_4195,In_560,In_441);
nor U4196 (N_4196,In_675,In_432);
nand U4197 (N_4197,In_473,In_993);
nand U4198 (N_4198,In_1165,In_439);
xor U4199 (N_4199,In_579,In_1215);
nor U4200 (N_4200,In_564,In_395);
and U4201 (N_4201,In_412,In_1347);
xor U4202 (N_4202,In_456,In_859);
or U4203 (N_4203,In_716,In_1302);
nand U4204 (N_4204,In_12,In_536);
and U4205 (N_4205,In_686,In_156);
nor U4206 (N_4206,In_746,In_433);
or U4207 (N_4207,In_1413,In_176);
xor U4208 (N_4208,In_252,In_747);
nor U4209 (N_4209,In_824,In_267);
nor U4210 (N_4210,In_246,In_89);
or U4211 (N_4211,In_1091,In_9);
or U4212 (N_4212,In_1239,In_936);
or U4213 (N_4213,In_712,In_585);
or U4214 (N_4214,In_152,In_354);
and U4215 (N_4215,In_588,In_1174);
nor U4216 (N_4216,In_477,In_349);
or U4217 (N_4217,In_178,In_921);
xnor U4218 (N_4218,In_248,In_1305);
nand U4219 (N_4219,In_941,In_714);
or U4220 (N_4220,In_1486,In_1464);
and U4221 (N_4221,In_158,In_184);
xnor U4222 (N_4222,In_152,In_1091);
nor U4223 (N_4223,In_379,In_580);
nand U4224 (N_4224,In_698,In_1364);
and U4225 (N_4225,In_1151,In_1426);
and U4226 (N_4226,In_323,In_458);
or U4227 (N_4227,In_1465,In_62);
xnor U4228 (N_4228,In_1062,In_162);
and U4229 (N_4229,In_85,In_627);
nand U4230 (N_4230,In_1393,In_1280);
nand U4231 (N_4231,In_1395,In_700);
and U4232 (N_4232,In_1267,In_861);
xor U4233 (N_4233,In_1078,In_661);
or U4234 (N_4234,In_495,In_680);
or U4235 (N_4235,In_759,In_1392);
nand U4236 (N_4236,In_1351,In_298);
nand U4237 (N_4237,In_1429,In_540);
nand U4238 (N_4238,In_932,In_1078);
and U4239 (N_4239,In_1300,In_930);
nor U4240 (N_4240,In_273,In_1058);
and U4241 (N_4241,In_721,In_270);
and U4242 (N_4242,In_750,In_1271);
nand U4243 (N_4243,In_467,In_197);
nor U4244 (N_4244,In_422,In_871);
or U4245 (N_4245,In_1012,In_1119);
or U4246 (N_4246,In_716,In_981);
or U4247 (N_4247,In_252,In_518);
nor U4248 (N_4248,In_447,In_419);
nand U4249 (N_4249,In_1142,In_1320);
nand U4250 (N_4250,In_1052,In_1487);
nand U4251 (N_4251,In_178,In_977);
and U4252 (N_4252,In_220,In_364);
nand U4253 (N_4253,In_1296,In_641);
nor U4254 (N_4254,In_1332,In_26);
nor U4255 (N_4255,In_1168,In_982);
nor U4256 (N_4256,In_883,In_1489);
xnor U4257 (N_4257,In_292,In_314);
or U4258 (N_4258,In_1031,In_452);
xor U4259 (N_4259,In_607,In_225);
and U4260 (N_4260,In_212,In_777);
and U4261 (N_4261,In_602,In_275);
and U4262 (N_4262,In_1129,In_474);
and U4263 (N_4263,In_376,In_948);
and U4264 (N_4264,In_1417,In_1137);
nand U4265 (N_4265,In_1203,In_223);
nand U4266 (N_4266,In_816,In_745);
and U4267 (N_4267,In_136,In_1165);
nor U4268 (N_4268,In_1365,In_503);
xor U4269 (N_4269,In_1388,In_1098);
nand U4270 (N_4270,In_643,In_210);
and U4271 (N_4271,In_678,In_550);
or U4272 (N_4272,In_1426,In_184);
nor U4273 (N_4273,In_1410,In_528);
and U4274 (N_4274,In_329,In_246);
nor U4275 (N_4275,In_538,In_1067);
nand U4276 (N_4276,In_6,In_35);
nand U4277 (N_4277,In_1408,In_7);
nor U4278 (N_4278,In_234,In_1324);
and U4279 (N_4279,In_1368,In_1265);
xor U4280 (N_4280,In_527,In_618);
or U4281 (N_4281,In_1166,In_1154);
nand U4282 (N_4282,In_821,In_383);
or U4283 (N_4283,In_1106,In_979);
and U4284 (N_4284,In_1281,In_335);
nand U4285 (N_4285,In_747,In_974);
nand U4286 (N_4286,In_420,In_530);
nand U4287 (N_4287,In_993,In_890);
or U4288 (N_4288,In_329,In_538);
nor U4289 (N_4289,In_301,In_1038);
nor U4290 (N_4290,In_1220,In_312);
nand U4291 (N_4291,In_792,In_695);
or U4292 (N_4292,In_669,In_1120);
nand U4293 (N_4293,In_969,In_1104);
nor U4294 (N_4294,In_403,In_627);
nor U4295 (N_4295,In_688,In_966);
nor U4296 (N_4296,In_931,In_599);
nor U4297 (N_4297,In_1429,In_1139);
nand U4298 (N_4298,In_280,In_1350);
xor U4299 (N_4299,In_670,In_1124);
and U4300 (N_4300,In_647,In_990);
or U4301 (N_4301,In_902,In_1322);
or U4302 (N_4302,In_654,In_1387);
xor U4303 (N_4303,In_1094,In_843);
nand U4304 (N_4304,In_377,In_598);
xnor U4305 (N_4305,In_480,In_707);
nor U4306 (N_4306,In_1423,In_1308);
and U4307 (N_4307,In_1172,In_260);
nor U4308 (N_4308,In_369,In_66);
and U4309 (N_4309,In_1027,In_572);
nor U4310 (N_4310,In_954,In_410);
nor U4311 (N_4311,In_673,In_1395);
nand U4312 (N_4312,In_1320,In_976);
nand U4313 (N_4313,In_1329,In_935);
nand U4314 (N_4314,In_6,In_1499);
xnor U4315 (N_4315,In_111,In_227);
nor U4316 (N_4316,In_1449,In_485);
nor U4317 (N_4317,In_478,In_1158);
xnor U4318 (N_4318,In_1018,In_635);
nand U4319 (N_4319,In_19,In_664);
or U4320 (N_4320,In_947,In_254);
nand U4321 (N_4321,In_1009,In_569);
and U4322 (N_4322,In_1161,In_325);
nor U4323 (N_4323,In_169,In_822);
nor U4324 (N_4324,In_247,In_450);
nor U4325 (N_4325,In_252,In_1303);
nor U4326 (N_4326,In_648,In_995);
and U4327 (N_4327,In_540,In_763);
xnor U4328 (N_4328,In_127,In_66);
xnor U4329 (N_4329,In_1385,In_1030);
nand U4330 (N_4330,In_196,In_741);
or U4331 (N_4331,In_341,In_101);
or U4332 (N_4332,In_1200,In_880);
or U4333 (N_4333,In_112,In_1199);
nand U4334 (N_4334,In_1343,In_238);
nand U4335 (N_4335,In_783,In_1148);
nand U4336 (N_4336,In_1286,In_1109);
nor U4337 (N_4337,In_645,In_815);
nand U4338 (N_4338,In_286,In_1029);
or U4339 (N_4339,In_1174,In_187);
xor U4340 (N_4340,In_108,In_1359);
or U4341 (N_4341,In_1327,In_504);
nor U4342 (N_4342,In_840,In_279);
and U4343 (N_4343,In_426,In_508);
and U4344 (N_4344,In_208,In_1392);
nor U4345 (N_4345,In_1082,In_363);
nor U4346 (N_4346,In_171,In_1410);
and U4347 (N_4347,In_621,In_418);
xor U4348 (N_4348,In_229,In_1256);
nand U4349 (N_4349,In_1288,In_1362);
or U4350 (N_4350,In_336,In_647);
xor U4351 (N_4351,In_1248,In_1453);
nand U4352 (N_4352,In_670,In_728);
nand U4353 (N_4353,In_92,In_1331);
nand U4354 (N_4354,In_1046,In_1216);
xnor U4355 (N_4355,In_742,In_1232);
nor U4356 (N_4356,In_1456,In_413);
nor U4357 (N_4357,In_623,In_1398);
and U4358 (N_4358,In_927,In_408);
nand U4359 (N_4359,In_678,In_565);
nor U4360 (N_4360,In_992,In_579);
nand U4361 (N_4361,In_580,In_1375);
or U4362 (N_4362,In_759,In_420);
xor U4363 (N_4363,In_367,In_630);
nand U4364 (N_4364,In_630,In_980);
or U4365 (N_4365,In_68,In_332);
nand U4366 (N_4366,In_767,In_919);
nor U4367 (N_4367,In_715,In_676);
nor U4368 (N_4368,In_1186,In_539);
nand U4369 (N_4369,In_1120,In_73);
xnor U4370 (N_4370,In_93,In_1036);
nor U4371 (N_4371,In_59,In_1298);
and U4372 (N_4372,In_778,In_439);
xnor U4373 (N_4373,In_860,In_1089);
nor U4374 (N_4374,In_121,In_58);
nand U4375 (N_4375,In_1058,In_968);
nand U4376 (N_4376,In_670,In_1219);
xnor U4377 (N_4377,In_2,In_568);
xnor U4378 (N_4378,In_701,In_724);
or U4379 (N_4379,In_965,In_1433);
and U4380 (N_4380,In_347,In_815);
and U4381 (N_4381,In_458,In_834);
nand U4382 (N_4382,In_1364,In_692);
and U4383 (N_4383,In_1266,In_1021);
or U4384 (N_4384,In_1133,In_954);
or U4385 (N_4385,In_1015,In_1072);
nor U4386 (N_4386,In_556,In_1226);
nor U4387 (N_4387,In_4,In_473);
nand U4388 (N_4388,In_1387,In_387);
xnor U4389 (N_4389,In_119,In_1393);
and U4390 (N_4390,In_916,In_839);
nor U4391 (N_4391,In_1495,In_605);
or U4392 (N_4392,In_1227,In_212);
xor U4393 (N_4393,In_1015,In_621);
xor U4394 (N_4394,In_16,In_249);
or U4395 (N_4395,In_659,In_62);
and U4396 (N_4396,In_1063,In_879);
or U4397 (N_4397,In_800,In_353);
and U4398 (N_4398,In_1298,In_342);
xnor U4399 (N_4399,In_878,In_352);
xor U4400 (N_4400,In_893,In_704);
or U4401 (N_4401,In_1127,In_746);
nor U4402 (N_4402,In_949,In_942);
and U4403 (N_4403,In_1202,In_389);
nand U4404 (N_4404,In_14,In_540);
and U4405 (N_4405,In_1167,In_495);
xnor U4406 (N_4406,In_1167,In_912);
and U4407 (N_4407,In_682,In_1148);
nand U4408 (N_4408,In_1050,In_1096);
nand U4409 (N_4409,In_619,In_104);
or U4410 (N_4410,In_1202,In_163);
nor U4411 (N_4411,In_593,In_951);
xor U4412 (N_4412,In_1304,In_257);
or U4413 (N_4413,In_930,In_249);
nor U4414 (N_4414,In_1079,In_1137);
nand U4415 (N_4415,In_114,In_653);
nor U4416 (N_4416,In_274,In_558);
or U4417 (N_4417,In_206,In_588);
nor U4418 (N_4418,In_310,In_1202);
nor U4419 (N_4419,In_596,In_906);
nand U4420 (N_4420,In_80,In_1289);
and U4421 (N_4421,In_151,In_648);
or U4422 (N_4422,In_1152,In_600);
nor U4423 (N_4423,In_512,In_974);
nor U4424 (N_4424,In_1333,In_760);
xnor U4425 (N_4425,In_741,In_554);
nand U4426 (N_4426,In_577,In_675);
and U4427 (N_4427,In_1467,In_1305);
or U4428 (N_4428,In_1409,In_974);
nor U4429 (N_4429,In_1041,In_949);
nor U4430 (N_4430,In_669,In_897);
and U4431 (N_4431,In_1469,In_1144);
nor U4432 (N_4432,In_1238,In_175);
or U4433 (N_4433,In_1406,In_1367);
xor U4434 (N_4434,In_923,In_852);
or U4435 (N_4435,In_1099,In_1056);
xor U4436 (N_4436,In_180,In_1458);
and U4437 (N_4437,In_334,In_1199);
nand U4438 (N_4438,In_467,In_1220);
nand U4439 (N_4439,In_792,In_830);
nor U4440 (N_4440,In_1280,In_1095);
and U4441 (N_4441,In_1353,In_858);
xor U4442 (N_4442,In_451,In_58);
nor U4443 (N_4443,In_1262,In_885);
nand U4444 (N_4444,In_1496,In_220);
nand U4445 (N_4445,In_218,In_548);
nor U4446 (N_4446,In_1173,In_999);
and U4447 (N_4447,In_876,In_141);
xor U4448 (N_4448,In_86,In_523);
xnor U4449 (N_4449,In_909,In_450);
nor U4450 (N_4450,In_785,In_1341);
nand U4451 (N_4451,In_332,In_554);
nor U4452 (N_4452,In_841,In_1285);
nor U4453 (N_4453,In_478,In_923);
nand U4454 (N_4454,In_619,In_1119);
nand U4455 (N_4455,In_1098,In_637);
nor U4456 (N_4456,In_913,In_1401);
nor U4457 (N_4457,In_661,In_1209);
xnor U4458 (N_4458,In_41,In_297);
nor U4459 (N_4459,In_529,In_151);
nor U4460 (N_4460,In_468,In_88);
nor U4461 (N_4461,In_547,In_176);
or U4462 (N_4462,In_600,In_833);
nor U4463 (N_4463,In_250,In_1494);
xnor U4464 (N_4464,In_2,In_841);
nor U4465 (N_4465,In_125,In_115);
and U4466 (N_4466,In_336,In_738);
nor U4467 (N_4467,In_1009,In_940);
xor U4468 (N_4468,In_357,In_721);
nand U4469 (N_4469,In_603,In_103);
nor U4470 (N_4470,In_1109,In_944);
nor U4471 (N_4471,In_1072,In_1458);
nor U4472 (N_4472,In_974,In_86);
and U4473 (N_4473,In_702,In_892);
or U4474 (N_4474,In_1426,In_1252);
nand U4475 (N_4475,In_124,In_1034);
and U4476 (N_4476,In_43,In_1000);
xor U4477 (N_4477,In_1140,In_914);
and U4478 (N_4478,In_538,In_761);
nand U4479 (N_4479,In_1389,In_421);
xnor U4480 (N_4480,In_1272,In_1032);
nor U4481 (N_4481,In_33,In_2);
or U4482 (N_4482,In_1125,In_180);
nand U4483 (N_4483,In_407,In_1469);
nand U4484 (N_4484,In_1361,In_416);
xnor U4485 (N_4485,In_1287,In_772);
nor U4486 (N_4486,In_783,In_674);
and U4487 (N_4487,In_1327,In_697);
nand U4488 (N_4488,In_401,In_1345);
xnor U4489 (N_4489,In_178,In_480);
or U4490 (N_4490,In_187,In_1165);
xnor U4491 (N_4491,In_1338,In_662);
nor U4492 (N_4492,In_471,In_772);
nand U4493 (N_4493,In_1323,In_1141);
and U4494 (N_4494,In_165,In_82);
nand U4495 (N_4495,In_137,In_973);
and U4496 (N_4496,In_769,In_1143);
or U4497 (N_4497,In_130,In_525);
or U4498 (N_4498,In_426,In_999);
xnor U4499 (N_4499,In_1119,In_67);
or U4500 (N_4500,In_999,In_592);
and U4501 (N_4501,In_536,In_229);
or U4502 (N_4502,In_109,In_58);
nor U4503 (N_4503,In_943,In_1146);
xnor U4504 (N_4504,In_1089,In_414);
xnor U4505 (N_4505,In_775,In_745);
or U4506 (N_4506,In_871,In_1311);
or U4507 (N_4507,In_97,In_55);
xor U4508 (N_4508,In_584,In_76);
xor U4509 (N_4509,In_855,In_58);
and U4510 (N_4510,In_825,In_562);
xor U4511 (N_4511,In_96,In_779);
or U4512 (N_4512,In_780,In_864);
nor U4513 (N_4513,In_151,In_1061);
and U4514 (N_4514,In_948,In_242);
or U4515 (N_4515,In_874,In_248);
xnor U4516 (N_4516,In_2,In_764);
and U4517 (N_4517,In_1468,In_1360);
nor U4518 (N_4518,In_1327,In_1333);
nand U4519 (N_4519,In_1331,In_761);
xnor U4520 (N_4520,In_979,In_247);
nor U4521 (N_4521,In_580,In_1390);
or U4522 (N_4522,In_788,In_407);
nand U4523 (N_4523,In_1125,In_1487);
or U4524 (N_4524,In_43,In_466);
nand U4525 (N_4525,In_957,In_144);
and U4526 (N_4526,In_685,In_1012);
or U4527 (N_4527,In_484,In_1156);
or U4528 (N_4528,In_1451,In_753);
xnor U4529 (N_4529,In_461,In_748);
and U4530 (N_4530,In_797,In_336);
xnor U4531 (N_4531,In_1036,In_1087);
and U4532 (N_4532,In_390,In_1486);
nand U4533 (N_4533,In_129,In_672);
xor U4534 (N_4534,In_269,In_886);
and U4535 (N_4535,In_641,In_669);
nor U4536 (N_4536,In_94,In_1071);
xnor U4537 (N_4537,In_1379,In_796);
and U4538 (N_4538,In_440,In_250);
or U4539 (N_4539,In_87,In_210);
xor U4540 (N_4540,In_4,In_888);
or U4541 (N_4541,In_380,In_887);
nor U4542 (N_4542,In_74,In_226);
nand U4543 (N_4543,In_1182,In_910);
nor U4544 (N_4544,In_527,In_991);
and U4545 (N_4545,In_158,In_1327);
nor U4546 (N_4546,In_111,In_917);
xnor U4547 (N_4547,In_1088,In_1433);
nand U4548 (N_4548,In_832,In_673);
nor U4549 (N_4549,In_1360,In_222);
nor U4550 (N_4550,In_34,In_1211);
nor U4551 (N_4551,In_364,In_1042);
xnor U4552 (N_4552,In_837,In_1473);
nor U4553 (N_4553,In_81,In_572);
and U4554 (N_4554,In_1176,In_37);
nand U4555 (N_4555,In_235,In_1465);
nand U4556 (N_4556,In_1410,In_13);
xnor U4557 (N_4557,In_144,In_739);
nor U4558 (N_4558,In_722,In_921);
or U4559 (N_4559,In_1317,In_809);
and U4560 (N_4560,In_410,In_77);
and U4561 (N_4561,In_878,In_873);
and U4562 (N_4562,In_1299,In_437);
and U4563 (N_4563,In_860,In_35);
nand U4564 (N_4564,In_386,In_888);
or U4565 (N_4565,In_1138,In_273);
and U4566 (N_4566,In_426,In_967);
nor U4567 (N_4567,In_858,In_390);
nor U4568 (N_4568,In_546,In_789);
and U4569 (N_4569,In_553,In_1206);
and U4570 (N_4570,In_739,In_52);
nor U4571 (N_4571,In_1434,In_593);
xnor U4572 (N_4572,In_44,In_75);
or U4573 (N_4573,In_187,In_1164);
nand U4574 (N_4574,In_382,In_489);
nand U4575 (N_4575,In_42,In_1043);
or U4576 (N_4576,In_963,In_275);
xnor U4577 (N_4577,In_516,In_600);
nor U4578 (N_4578,In_901,In_111);
or U4579 (N_4579,In_1488,In_966);
nand U4580 (N_4580,In_1132,In_924);
nand U4581 (N_4581,In_1126,In_100);
and U4582 (N_4582,In_794,In_803);
nand U4583 (N_4583,In_825,In_798);
xor U4584 (N_4584,In_815,In_1381);
xnor U4585 (N_4585,In_770,In_341);
or U4586 (N_4586,In_1346,In_204);
nor U4587 (N_4587,In_783,In_912);
or U4588 (N_4588,In_686,In_245);
nand U4589 (N_4589,In_416,In_417);
nor U4590 (N_4590,In_693,In_920);
and U4591 (N_4591,In_508,In_86);
xor U4592 (N_4592,In_705,In_678);
xnor U4593 (N_4593,In_769,In_1318);
xor U4594 (N_4594,In_842,In_955);
xnor U4595 (N_4595,In_313,In_1096);
nand U4596 (N_4596,In_126,In_461);
or U4597 (N_4597,In_781,In_774);
or U4598 (N_4598,In_414,In_126);
or U4599 (N_4599,In_213,In_1145);
and U4600 (N_4600,In_1302,In_35);
xor U4601 (N_4601,In_576,In_720);
nand U4602 (N_4602,In_1450,In_1148);
nor U4603 (N_4603,In_889,In_494);
nand U4604 (N_4604,In_39,In_353);
nor U4605 (N_4605,In_1457,In_1337);
nand U4606 (N_4606,In_316,In_346);
nand U4607 (N_4607,In_655,In_1449);
nor U4608 (N_4608,In_1328,In_562);
nor U4609 (N_4609,In_1207,In_662);
nor U4610 (N_4610,In_663,In_924);
and U4611 (N_4611,In_923,In_223);
and U4612 (N_4612,In_463,In_460);
xor U4613 (N_4613,In_1327,In_674);
and U4614 (N_4614,In_466,In_459);
or U4615 (N_4615,In_348,In_309);
nand U4616 (N_4616,In_662,In_770);
xnor U4617 (N_4617,In_1017,In_203);
or U4618 (N_4618,In_1374,In_483);
nor U4619 (N_4619,In_1393,In_396);
or U4620 (N_4620,In_1188,In_149);
nor U4621 (N_4621,In_1095,In_1305);
nand U4622 (N_4622,In_1461,In_1453);
or U4623 (N_4623,In_1382,In_96);
or U4624 (N_4624,In_463,In_1378);
xnor U4625 (N_4625,In_207,In_695);
nor U4626 (N_4626,In_121,In_1402);
xor U4627 (N_4627,In_1349,In_457);
or U4628 (N_4628,In_1007,In_706);
xor U4629 (N_4629,In_669,In_1375);
nand U4630 (N_4630,In_1176,In_1289);
nand U4631 (N_4631,In_154,In_1111);
xor U4632 (N_4632,In_1215,In_810);
nor U4633 (N_4633,In_1302,In_40);
or U4634 (N_4634,In_1452,In_1480);
xnor U4635 (N_4635,In_814,In_992);
nor U4636 (N_4636,In_14,In_118);
nand U4637 (N_4637,In_820,In_1172);
nor U4638 (N_4638,In_1263,In_1284);
nand U4639 (N_4639,In_555,In_795);
xor U4640 (N_4640,In_486,In_648);
nand U4641 (N_4641,In_611,In_815);
nand U4642 (N_4642,In_936,In_611);
or U4643 (N_4643,In_465,In_1306);
nand U4644 (N_4644,In_666,In_796);
nand U4645 (N_4645,In_618,In_613);
or U4646 (N_4646,In_999,In_469);
nand U4647 (N_4647,In_151,In_817);
nor U4648 (N_4648,In_647,In_459);
and U4649 (N_4649,In_57,In_1383);
xor U4650 (N_4650,In_473,In_1130);
nor U4651 (N_4651,In_1151,In_922);
or U4652 (N_4652,In_1229,In_664);
nor U4653 (N_4653,In_735,In_881);
or U4654 (N_4654,In_566,In_782);
and U4655 (N_4655,In_186,In_1457);
nor U4656 (N_4656,In_1093,In_190);
nand U4657 (N_4657,In_378,In_903);
nand U4658 (N_4658,In_1094,In_417);
xnor U4659 (N_4659,In_1442,In_775);
nor U4660 (N_4660,In_809,In_929);
and U4661 (N_4661,In_371,In_417);
and U4662 (N_4662,In_117,In_1252);
nand U4663 (N_4663,In_1489,In_241);
and U4664 (N_4664,In_1312,In_872);
xor U4665 (N_4665,In_1442,In_200);
or U4666 (N_4666,In_772,In_723);
nand U4667 (N_4667,In_184,In_282);
or U4668 (N_4668,In_812,In_211);
nor U4669 (N_4669,In_56,In_565);
nand U4670 (N_4670,In_509,In_1093);
nor U4671 (N_4671,In_124,In_130);
xor U4672 (N_4672,In_778,In_473);
nand U4673 (N_4673,In_1004,In_1401);
or U4674 (N_4674,In_560,In_489);
or U4675 (N_4675,In_1112,In_151);
or U4676 (N_4676,In_307,In_276);
and U4677 (N_4677,In_607,In_661);
nor U4678 (N_4678,In_1073,In_808);
and U4679 (N_4679,In_585,In_1150);
nand U4680 (N_4680,In_627,In_1127);
xor U4681 (N_4681,In_447,In_118);
nand U4682 (N_4682,In_1439,In_933);
and U4683 (N_4683,In_1075,In_1359);
or U4684 (N_4684,In_718,In_665);
or U4685 (N_4685,In_1396,In_509);
nor U4686 (N_4686,In_1417,In_445);
nor U4687 (N_4687,In_726,In_982);
xor U4688 (N_4688,In_1429,In_197);
nand U4689 (N_4689,In_1229,In_1418);
xor U4690 (N_4690,In_563,In_1389);
nand U4691 (N_4691,In_190,In_1173);
nand U4692 (N_4692,In_332,In_24);
nand U4693 (N_4693,In_573,In_1195);
nand U4694 (N_4694,In_858,In_1410);
xnor U4695 (N_4695,In_1355,In_539);
xnor U4696 (N_4696,In_965,In_1316);
nand U4697 (N_4697,In_587,In_1279);
nor U4698 (N_4698,In_1393,In_1032);
xor U4699 (N_4699,In_1387,In_370);
xnor U4700 (N_4700,In_1174,In_1196);
nand U4701 (N_4701,In_1343,In_1459);
nor U4702 (N_4702,In_544,In_843);
xor U4703 (N_4703,In_1371,In_572);
nand U4704 (N_4704,In_80,In_445);
nand U4705 (N_4705,In_1345,In_1402);
nor U4706 (N_4706,In_1435,In_660);
nor U4707 (N_4707,In_431,In_1000);
nand U4708 (N_4708,In_312,In_1488);
nor U4709 (N_4709,In_1307,In_18);
or U4710 (N_4710,In_1400,In_897);
xor U4711 (N_4711,In_29,In_319);
or U4712 (N_4712,In_449,In_192);
and U4713 (N_4713,In_613,In_854);
nor U4714 (N_4714,In_806,In_820);
and U4715 (N_4715,In_364,In_68);
nor U4716 (N_4716,In_97,In_815);
xnor U4717 (N_4717,In_1287,In_1437);
or U4718 (N_4718,In_1247,In_1451);
and U4719 (N_4719,In_872,In_951);
nand U4720 (N_4720,In_658,In_507);
or U4721 (N_4721,In_1337,In_1497);
or U4722 (N_4722,In_746,In_500);
nor U4723 (N_4723,In_494,In_1435);
or U4724 (N_4724,In_463,In_636);
xor U4725 (N_4725,In_422,In_198);
nor U4726 (N_4726,In_1445,In_1292);
xor U4727 (N_4727,In_973,In_654);
nand U4728 (N_4728,In_402,In_624);
xnor U4729 (N_4729,In_1047,In_462);
or U4730 (N_4730,In_305,In_120);
or U4731 (N_4731,In_1098,In_400);
or U4732 (N_4732,In_1337,In_1102);
nor U4733 (N_4733,In_991,In_104);
xor U4734 (N_4734,In_1394,In_13);
and U4735 (N_4735,In_587,In_757);
nand U4736 (N_4736,In_207,In_1388);
nor U4737 (N_4737,In_1003,In_727);
and U4738 (N_4738,In_263,In_95);
nand U4739 (N_4739,In_1490,In_721);
nor U4740 (N_4740,In_733,In_1122);
or U4741 (N_4741,In_1233,In_1188);
and U4742 (N_4742,In_551,In_221);
nand U4743 (N_4743,In_29,In_61);
and U4744 (N_4744,In_916,In_577);
nand U4745 (N_4745,In_320,In_383);
or U4746 (N_4746,In_942,In_1048);
nand U4747 (N_4747,In_113,In_169);
nand U4748 (N_4748,In_1046,In_466);
and U4749 (N_4749,In_713,In_1046);
and U4750 (N_4750,In_114,In_1317);
xor U4751 (N_4751,In_230,In_50);
nor U4752 (N_4752,In_269,In_147);
nand U4753 (N_4753,In_814,In_1262);
nand U4754 (N_4754,In_779,In_452);
or U4755 (N_4755,In_1205,In_20);
nand U4756 (N_4756,In_801,In_1296);
nor U4757 (N_4757,In_1306,In_887);
nand U4758 (N_4758,In_283,In_1243);
or U4759 (N_4759,In_359,In_1252);
or U4760 (N_4760,In_1496,In_235);
xor U4761 (N_4761,In_479,In_1213);
nand U4762 (N_4762,In_1309,In_501);
nand U4763 (N_4763,In_1453,In_481);
nand U4764 (N_4764,In_486,In_965);
nand U4765 (N_4765,In_804,In_1115);
and U4766 (N_4766,In_237,In_330);
nor U4767 (N_4767,In_628,In_1122);
nor U4768 (N_4768,In_192,In_1457);
nand U4769 (N_4769,In_1472,In_10);
or U4770 (N_4770,In_1236,In_1067);
nor U4771 (N_4771,In_711,In_1162);
nand U4772 (N_4772,In_728,In_560);
or U4773 (N_4773,In_1240,In_1367);
and U4774 (N_4774,In_12,In_400);
xnor U4775 (N_4775,In_867,In_1060);
nor U4776 (N_4776,In_539,In_583);
nor U4777 (N_4777,In_177,In_1112);
xor U4778 (N_4778,In_803,In_200);
and U4779 (N_4779,In_10,In_1236);
or U4780 (N_4780,In_10,In_704);
nor U4781 (N_4781,In_822,In_1056);
xor U4782 (N_4782,In_1478,In_138);
and U4783 (N_4783,In_681,In_202);
xor U4784 (N_4784,In_1046,In_935);
and U4785 (N_4785,In_1317,In_1090);
nand U4786 (N_4786,In_967,In_666);
and U4787 (N_4787,In_887,In_71);
nand U4788 (N_4788,In_739,In_782);
nand U4789 (N_4789,In_136,In_993);
or U4790 (N_4790,In_194,In_1476);
nor U4791 (N_4791,In_1227,In_841);
and U4792 (N_4792,In_1232,In_749);
and U4793 (N_4793,In_563,In_178);
or U4794 (N_4794,In_86,In_31);
nor U4795 (N_4795,In_791,In_851);
nor U4796 (N_4796,In_1144,In_1178);
and U4797 (N_4797,In_845,In_914);
nand U4798 (N_4798,In_1269,In_1126);
nand U4799 (N_4799,In_580,In_867);
and U4800 (N_4800,In_231,In_1188);
or U4801 (N_4801,In_1235,In_175);
xor U4802 (N_4802,In_848,In_1133);
and U4803 (N_4803,In_353,In_573);
or U4804 (N_4804,In_507,In_647);
or U4805 (N_4805,In_828,In_1301);
nor U4806 (N_4806,In_79,In_1322);
or U4807 (N_4807,In_426,In_896);
and U4808 (N_4808,In_741,In_1317);
and U4809 (N_4809,In_509,In_305);
nand U4810 (N_4810,In_1217,In_997);
nand U4811 (N_4811,In_603,In_119);
nor U4812 (N_4812,In_1414,In_732);
and U4813 (N_4813,In_612,In_848);
nand U4814 (N_4814,In_138,In_989);
nor U4815 (N_4815,In_12,In_217);
and U4816 (N_4816,In_1030,In_1003);
nand U4817 (N_4817,In_779,In_990);
nor U4818 (N_4818,In_889,In_499);
nand U4819 (N_4819,In_1170,In_1387);
nor U4820 (N_4820,In_631,In_1170);
nand U4821 (N_4821,In_2,In_1161);
or U4822 (N_4822,In_1076,In_1145);
and U4823 (N_4823,In_1487,In_870);
nor U4824 (N_4824,In_1138,In_900);
xor U4825 (N_4825,In_721,In_950);
nand U4826 (N_4826,In_1156,In_244);
nor U4827 (N_4827,In_692,In_141);
xor U4828 (N_4828,In_931,In_3);
nor U4829 (N_4829,In_763,In_276);
and U4830 (N_4830,In_482,In_817);
and U4831 (N_4831,In_1099,In_1124);
or U4832 (N_4832,In_603,In_1034);
and U4833 (N_4833,In_671,In_419);
xor U4834 (N_4834,In_1152,In_1268);
nor U4835 (N_4835,In_769,In_1493);
nor U4836 (N_4836,In_86,In_47);
or U4837 (N_4837,In_474,In_1384);
and U4838 (N_4838,In_10,In_619);
xnor U4839 (N_4839,In_490,In_1039);
xor U4840 (N_4840,In_1053,In_1377);
xnor U4841 (N_4841,In_909,In_288);
or U4842 (N_4842,In_1418,In_1186);
nor U4843 (N_4843,In_557,In_846);
nand U4844 (N_4844,In_1379,In_1109);
xnor U4845 (N_4845,In_1380,In_102);
nor U4846 (N_4846,In_502,In_110);
and U4847 (N_4847,In_1187,In_916);
nand U4848 (N_4848,In_73,In_1453);
and U4849 (N_4849,In_1425,In_16);
xnor U4850 (N_4850,In_1402,In_15);
and U4851 (N_4851,In_1019,In_192);
xor U4852 (N_4852,In_683,In_561);
and U4853 (N_4853,In_338,In_163);
and U4854 (N_4854,In_149,In_237);
or U4855 (N_4855,In_1126,In_8);
xor U4856 (N_4856,In_314,In_1110);
or U4857 (N_4857,In_849,In_1424);
and U4858 (N_4858,In_73,In_360);
nor U4859 (N_4859,In_1447,In_339);
xor U4860 (N_4860,In_51,In_417);
and U4861 (N_4861,In_1235,In_1361);
nor U4862 (N_4862,In_101,In_1192);
xor U4863 (N_4863,In_244,In_1248);
nand U4864 (N_4864,In_657,In_1403);
or U4865 (N_4865,In_520,In_1264);
and U4866 (N_4866,In_750,In_461);
and U4867 (N_4867,In_1077,In_1309);
xor U4868 (N_4868,In_582,In_541);
nand U4869 (N_4869,In_115,In_740);
nor U4870 (N_4870,In_1290,In_764);
xnor U4871 (N_4871,In_435,In_341);
nand U4872 (N_4872,In_1127,In_825);
and U4873 (N_4873,In_135,In_1091);
nand U4874 (N_4874,In_34,In_1168);
or U4875 (N_4875,In_367,In_74);
xnor U4876 (N_4876,In_248,In_135);
or U4877 (N_4877,In_1045,In_1299);
nand U4878 (N_4878,In_1049,In_603);
and U4879 (N_4879,In_144,In_282);
xor U4880 (N_4880,In_1285,In_27);
xnor U4881 (N_4881,In_277,In_564);
or U4882 (N_4882,In_1440,In_1091);
and U4883 (N_4883,In_664,In_29);
nand U4884 (N_4884,In_860,In_666);
nor U4885 (N_4885,In_668,In_682);
xnor U4886 (N_4886,In_348,In_1096);
xnor U4887 (N_4887,In_126,In_22);
and U4888 (N_4888,In_91,In_634);
or U4889 (N_4889,In_1105,In_1014);
nand U4890 (N_4890,In_1290,In_1137);
nand U4891 (N_4891,In_107,In_584);
xnor U4892 (N_4892,In_1436,In_1471);
or U4893 (N_4893,In_819,In_1462);
nor U4894 (N_4894,In_532,In_41);
and U4895 (N_4895,In_875,In_464);
nand U4896 (N_4896,In_1291,In_184);
nor U4897 (N_4897,In_1290,In_491);
nand U4898 (N_4898,In_1388,In_665);
or U4899 (N_4899,In_871,In_757);
xor U4900 (N_4900,In_1051,In_434);
nor U4901 (N_4901,In_1348,In_496);
nor U4902 (N_4902,In_327,In_543);
and U4903 (N_4903,In_1444,In_1468);
or U4904 (N_4904,In_303,In_164);
or U4905 (N_4905,In_692,In_350);
nor U4906 (N_4906,In_969,In_1082);
nor U4907 (N_4907,In_104,In_844);
or U4908 (N_4908,In_1425,In_39);
and U4909 (N_4909,In_764,In_208);
xnor U4910 (N_4910,In_1167,In_17);
or U4911 (N_4911,In_647,In_736);
nand U4912 (N_4912,In_1250,In_24);
nor U4913 (N_4913,In_1463,In_772);
nor U4914 (N_4914,In_208,In_257);
and U4915 (N_4915,In_398,In_1383);
and U4916 (N_4916,In_639,In_56);
nand U4917 (N_4917,In_1129,In_430);
and U4918 (N_4918,In_302,In_1079);
xor U4919 (N_4919,In_1371,In_1464);
and U4920 (N_4920,In_642,In_1474);
xnor U4921 (N_4921,In_1443,In_1464);
nor U4922 (N_4922,In_1336,In_152);
and U4923 (N_4923,In_1246,In_240);
and U4924 (N_4924,In_1387,In_833);
nand U4925 (N_4925,In_1260,In_1268);
and U4926 (N_4926,In_1094,In_1261);
or U4927 (N_4927,In_105,In_615);
or U4928 (N_4928,In_1325,In_762);
or U4929 (N_4929,In_1279,In_70);
nand U4930 (N_4930,In_257,In_1155);
and U4931 (N_4931,In_279,In_964);
xnor U4932 (N_4932,In_865,In_760);
xnor U4933 (N_4933,In_827,In_859);
nand U4934 (N_4934,In_14,In_1072);
and U4935 (N_4935,In_1233,In_535);
nand U4936 (N_4936,In_953,In_173);
xnor U4937 (N_4937,In_349,In_208);
nor U4938 (N_4938,In_189,In_1170);
nand U4939 (N_4939,In_352,In_303);
nand U4940 (N_4940,In_1335,In_567);
nor U4941 (N_4941,In_1384,In_1283);
nand U4942 (N_4942,In_244,In_581);
and U4943 (N_4943,In_965,In_31);
nor U4944 (N_4944,In_581,In_1329);
nor U4945 (N_4945,In_882,In_1110);
or U4946 (N_4946,In_385,In_850);
nor U4947 (N_4947,In_1334,In_811);
nand U4948 (N_4948,In_896,In_1145);
and U4949 (N_4949,In_670,In_137);
and U4950 (N_4950,In_1455,In_17);
xnor U4951 (N_4951,In_1028,In_1220);
or U4952 (N_4952,In_932,In_550);
xnor U4953 (N_4953,In_142,In_202);
nand U4954 (N_4954,In_761,In_478);
nor U4955 (N_4955,In_817,In_1061);
xnor U4956 (N_4956,In_659,In_634);
or U4957 (N_4957,In_897,In_1338);
or U4958 (N_4958,In_784,In_255);
nor U4959 (N_4959,In_681,In_508);
xor U4960 (N_4960,In_778,In_739);
nor U4961 (N_4961,In_1430,In_399);
or U4962 (N_4962,In_724,In_395);
and U4963 (N_4963,In_1016,In_185);
xnor U4964 (N_4964,In_188,In_1141);
and U4965 (N_4965,In_116,In_664);
nand U4966 (N_4966,In_398,In_4);
nor U4967 (N_4967,In_740,In_1367);
nor U4968 (N_4968,In_1099,In_252);
nor U4969 (N_4969,In_462,In_324);
and U4970 (N_4970,In_1228,In_724);
and U4971 (N_4971,In_132,In_1382);
xnor U4972 (N_4972,In_82,In_1295);
nor U4973 (N_4973,In_1254,In_1145);
nand U4974 (N_4974,In_362,In_1078);
xor U4975 (N_4975,In_761,In_102);
xnor U4976 (N_4976,In_854,In_210);
nand U4977 (N_4977,In_274,In_1198);
nand U4978 (N_4978,In_1354,In_627);
nand U4979 (N_4979,In_1078,In_1437);
nand U4980 (N_4980,In_823,In_625);
or U4981 (N_4981,In_598,In_1152);
nand U4982 (N_4982,In_1289,In_845);
and U4983 (N_4983,In_964,In_1341);
nand U4984 (N_4984,In_758,In_1246);
xnor U4985 (N_4985,In_102,In_1434);
or U4986 (N_4986,In_1138,In_1174);
nor U4987 (N_4987,In_544,In_1219);
xnor U4988 (N_4988,In_1367,In_157);
nor U4989 (N_4989,In_480,In_755);
xnor U4990 (N_4990,In_361,In_1136);
xor U4991 (N_4991,In_276,In_1499);
and U4992 (N_4992,In_1028,In_1230);
nand U4993 (N_4993,In_64,In_1365);
nand U4994 (N_4994,In_265,In_21);
nand U4995 (N_4995,In_917,In_935);
xnor U4996 (N_4996,In_948,In_9);
nor U4997 (N_4997,In_479,In_1259);
nor U4998 (N_4998,In_453,In_1200);
and U4999 (N_4999,In_12,In_1413);
nand U5000 (N_5000,N_2533,N_1745);
nor U5001 (N_5001,N_3666,N_460);
and U5002 (N_5002,N_2180,N_2541);
xor U5003 (N_5003,N_3137,N_3990);
or U5004 (N_5004,N_2364,N_3986);
or U5005 (N_5005,N_4572,N_4246);
nand U5006 (N_5006,N_682,N_3842);
or U5007 (N_5007,N_2860,N_4501);
xnor U5008 (N_5008,N_4297,N_858);
and U5009 (N_5009,N_2523,N_3275);
nand U5010 (N_5010,N_1471,N_398);
nor U5011 (N_5011,N_4015,N_66);
nor U5012 (N_5012,N_4870,N_2203);
nor U5013 (N_5013,N_463,N_227);
nor U5014 (N_5014,N_2782,N_334);
nand U5015 (N_5015,N_4684,N_4177);
and U5016 (N_5016,N_3680,N_3557);
nand U5017 (N_5017,N_4304,N_1419);
and U5018 (N_5018,N_4247,N_63);
and U5019 (N_5019,N_2023,N_915);
nor U5020 (N_5020,N_3399,N_2935);
and U5021 (N_5021,N_2504,N_2751);
nand U5022 (N_5022,N_532,N_1006);
nor U5023 (N_5023,N_2578,N_4701);
nor U5024 (N_5024,N_1063,N_3594);
xor U5025 (N_5025,N_3466,N_4775);
nand U5026 (N_5026,N_827,N_589);
nand U5027 (N_5027,N_4402,N_4351);
xor U5028 (N_5028,N_3372,N_1695);
or U5029 (N_5029,N_1603,N_3858);
or U5030 (N_5030,N_1691,N_4742);
or U5031 (N_5031,N_3463,N_4592);
nor U5032 (N_5032,N_3365,N_1384);
xor U5033 (N_5033,N_3462,N_4957);
nor U5034 (N_5034,N_4013,N_4662);
or U5035 (N_5035,N_2387,N_4685);
and U5036 (N_5036,N_3994,N_253);
or U5037 (N_5037,N_4654,N_1953);
xor U5038 (N_5038,N_4837,N_1360);
nor U5039 (N_5039,N_2419,N_466);
and U5040 (N_5040,N_780,N_618);
or U5041 (N_5041,N_1078,N_1388);
xor U5042 (N_5042,N_1511,N_1267);
nand U5043 (N_5043,N_1067,N_345);
nor U5044 (N_5044,N_3004,N_2526);
xor U5045 (N_5045,N_4976,N_1568);
or U5046 (N_5046,N_1940,N_162);
or U5047 (N_5047,N_3014,N_4365);
and U5048 (N_5048,N_1706,N_1948);
and U5049 (N_5049,N_2110,N_2626);
nand U5050 (N_5050,N_1024,N_945);
nor U5051 (N_5051,N_1076,N_2564);
and U5052 (N_5052,N_1802,N_2257);
or U5053 (N_5053,N_4869,N_4471);
or U5054 (N_5054,N_2147,N_431);
nor U5055 (N_5055,N_2583,N_3498);
or U5056 (N_5056,N_1469,N_2801);
or U5057 (N_5057,N_1122,N_4280);
nor U5058 (N_5058,N_1109,N_1100);
xor U5059 (N_5059,N_4787,N_1824);
nand U5060 (N_5060,N_904,N_3022);
or U5061 (N_5061,N_2947,N_1052);
xor U5062 (N_5062,N_1607,N_4300);
xor U5063 (N_5063,N_4108,N_4340);
and U5064 (N_5064,N_1296,N_3811);
xor U5065 (N_5065,N_2622,N_2666);
xnor U5066 (N_5066,N_4192,N_4476);
and U5067 (N_5067,N_1212,N_2448);
or U5068 (N_5068,N_2765,N_2356);
or U5069 (N_5069,N_1647,N_4276);
and U5070 (N_5070,N_3813,N_4499);
or U5071 (N_5071,N_1938,N_4479);
and U5072 (N_5072,N_1924,N_987);
nand U5073 (N_5073,N_3917,N_734);
xnor U5074 (N_5074,N_2657,N_685);
or U5075 (N_5075,N_1997,N_2922);
or U5076 (N_5076,N_4496,N_579);
nor U5077 (N_5077,N_4872,N_4797);
nor U5078 (N_5078,N_1001,N_2787);
or U5079 (N_5079,N_3102,N_4709);
nand U5080 (N_5080,N_2471,N_3565);
nor U5081 (N_5081,N_625,N_4871);
nand U5082 (N_5082,N_946,N_3091);
xnor U5083 (N_5083,N_424,N_886);
and U5084 (N_5084,N_2795,N_4689);
or U5085 (N_5085,N_1759,N_2334);
nor U5086 (N_5086,N_1071,N_1239);
nor U5087 (N_5087,N_1884,N_3590);
and U5088 (N_5088,N_2789,N_655);
nor U5089 (N_5089,N_909,N_2825);
nor U5090 (N_5090,N_4708,N_1875);
nand U5091 (N_5091,N_2444,N_1032);
xnor U5092 (N_5092,N_3177,N_3244);
nor U5093 (N_5093,N_2640,N_4289);
or U5094 (N_5094,N_73,N_4101);
nand U5095 (N_5095,N_2446,N_1379);
and U5096 (N_5096,N_916,N_4268);
xor U5097 (N_5097,N_479,N_2404);
nor U5098 (N_5098,N_3288,N_1519);
nand U5099 (N_5099,N_2510,N_1630);
xor U5100 (N_5100,N_3510,N_49);
xnor U5101 (N_5101,N_2687,N_748);
and U5102 (N_5102,N_4604,N_3097);
nor U5103 (N_5103,N_4676,N_3657);
nand U5104 (N_5104,N_1628,N_1265);
xor U5105 (N_5105,N_2136,N_660);
or U5106 (N_5106,N_3896,N_2024);
nand U5107 (N_5107,N_4643,N_3732);
or U5108 (N_5108,N_2405,N_3684);
nand U5109 (N_5109,N_1900,N_4745);
or U5110 (N_5110,N_4190,N_4919);
and U5111 (N_5111,N_2407,N_3052);
and U5112 (N_5112,N_1242,N_3330);
xor U5113 (N_5113,N_17,N_928);
nor U5114 (N_5114,N_3856,N_2366);
nand U5115 (N_5115,N_4765,N_2171);
and U5116 (N_5116,N_1530,N_1999);
and U5117 (N_5117,N_3017,N_4687);
or U5118 (N_5118,N_178,N_2007);
xnor U5119 (N_5119,N_1275,N_668);
nand U5120 (N_5120,N_4830,N_1372);
nand U5121 (N_5121,N_3563,N_645);
nand U5122 (N_5122,N_4645,N_3534);
or U5123 (N_5123,N_765,N_1725);
xnor U5124 (N_5124,N_1505,N_3524);
nand U5125 (N_5125,N_4714,N_2450);
nand U5126 (N_5126,N_4959,N_3519);
and U5127 (N_5127,N_4374,N_3297);
nor U5128 (N_5128,N_1373,N_3350);
or U5129 (N_5129,N_3380,N_4366);
nor U5130 (N_5130,N_1359,N_3092);
xor U5131 (N_5131,N_4807,N_12);
and U5132 (N_5132,N_3737,N_2679);
xor U5133 (N_5133,N_3391,N_937);
xor U5134 (N_5134,N_247,N_1522);
and U5135 (N_5135,N_2096,N_271);
or U5136 (N_5136,N_4978,N_174);
xnor U5137 (N_5137,N_4311,N_1363);
or U5138 (N_5138,N_2411,N_4914);
nor U5139 (N_5139,N_4903,N_2664);
xor U5140 (N_5140,N_4860,N_4754);
xor U5141 (N_5141,N_1793,N_245);
xnor U5142 (N_5142,N_1623,N_4142);
and U5143 (N_5143,N_590,N_2309);
nor U5144 (N_5144,N_4600,N_1143);
and U5145 (N_5145,N_449,N_4831);
nand U5146 (N_5146,N_3998,N_3315);
xnor U5147 (N_5147,N_974,N_2527);
or U5148 (N_5148,N_1182,N_2519);
nand U5149 (N_5149,N_3769,N_414);
and U5150 (N_5150,N_3311,N_3833);
nand U5151 (N_5151,N_3224,N_2443);
xor U5152 (N_5152,N_1258,N_3505);
or U5153 (N_5153,N_2712,N_3509);
nand U5154 (N_5154,N_2777,N_2037);
nor U5155 (N_5155,N_230,N_3474);
xnor U5156 (N_5156,N_1104,N_3772);
nor U5157 (N_5157,N_1529,N_752);
and U5158 (N_5158,N_2833,N_1491);
or U5159 (N_5159,N_1166,N_1184);
or U5160 (N_5160,N_4740,N_803);
nor U5161 (N_5161,N_3384,N_3877);
nand U5162 (N_5162,N_1035,N_1240);
nor U5163 (N_5163,N_4290,N_4703);
nor U5164 (N_5164,N_4805,N_1847);
nor U5165 (N_5165,N_4545,N_336);
xor U5166 (N_5166,N_365,N_2853);
xnor U5167 (N_5167,N_1936,N_3446);
nor U5168 (N_5168,N_416,N_328);
xor U5169 (N_5169,N_98,N_2786);
or U5170 (N_5170,N_243,N_2127);
xnor U5171 (N_5171,N_4429,N_3001);
xor U5172 (N_5172,N_234,N_591);
xnor U5173 (N_5173,N_2951,N_817);
nand U5174 (N_5174,N_2476,N_3490);
nor U5175 (N_5175,N_1825,N_979);
and U5176 (N_5176,N_705,N_3464);
and U5177 (N_5177,N_1831,N_2872);
or U5178 (N_5178,N_4343,N_282);
or U5179 (N_5179,N_1674,N_4704);
xnor U5180 (N_5180,N_3265,N_448);
and U5181 (N_5181,N_4691,N_795);
or U5182 (N_5182,N_2067,N_2149);
and U5183 (N_5183,N_4760,N_2633);
nor U5184 (N_5184,N_4046,N_1541);
nand U5185 (N_5185,N_2612,N_1701);
nor U5186 (N_5186,N_1190,N_866);
nand U5187 (N_5187,N_2974,N_1444);
nor U5188 (N_5188,N_742,N_1846);
and U5189 (N_5189,N_469,N_1783);
nor U5190 (N_5190,N_1806,N_4673);
xnor U5191 (N_5191,N_4639,N_4780);
and U5192 (N_5192,N_1921,N_3974);
xor U5193 (N_5193,N_2324,N_4436);
and U5194 (N_5194,N_4183,N_4763);
xnor U5195 (N_5195,N_3072,N_3724);
nand U5196 (N_5196,N_2039,N_4347);
nand U5197 (N_5197,N_3483,N_3438);
nand U5198 (N_5198,N_1513,N_3236);
nor U5199 (N_5199,N_788,N_4212);
or U5200 (N_5200,N_1199,N_4737);
xor U5201 (N_5201,N_1913,N_458);
or U5202 (N_5202,N_2472,N_1711);
xnor U5203 (N_5203,N_4725,N_329);
nor U5204 (N_5204,N_353,N_4900);
xor U5205 (N_5205,N_2827,N_3422);
nand U5206 (N_5206,N_4532,N_4517);
or U5207 (N_5207,N_4521,N_735);
nor U5208 (N_5208,N_2621,N_257);
and U5209 (N_5209,N_4448,N_4886);
or U5210 (N_5210,N_4424,N_1061);
nand U5211 (N_5211,N_4195,N_4204);
and U5212 (N_5212,N_1082,N_1315);
xnor U5213 (N_5213,N_2807,N_1213);
xnor U5214 (N_5214,N_2959,N_4659);
or U5215 (N_5215,N_507,N_4980);
xnor U5216 (N_5216,N_199,N_1778);
nor U5217 (N_5217,N_549,N_3303);
nor U5218 (N_5218,N_3306,N_3941);
or U5219 (N_5219,N_1099,N_959);
and U5220 (N_5220,N_3271,N_4842);
nor U5221 (N_5221,N_2018,N_2650);
nor U5222 (N_5222,N_501,N_2874);
nand U5223 (N_5223,N_1713,N_2544);
nand U5224 (N_5224,N_2454,N_955);
xnor U5225 (N_5225,N_2248,N_4984);
nor U5226 (N_5226,N_1776,N_2511);
nor U5227 (N_5227,N_1720,N_286);
nand U5228 (N_5228,N_2912,N_2080);
xor U5229 (N_5229,N_993,N_369);
nand U5230 (N_5230,N_1993,N_759);
and U5231 (N_5231,N_2477,N_3132);
xnor U5232 (N_5232,N_1362,N_1739);
xor U5233 (N_5233,N_2514,N_2655);
and U5234 (N_5234,N_1228,N_1738);
nand U5235 (N_5235,N_447,N_3797);
nor U5236 (N_5236,N_3909,N_4857);
or U5237 (N_5237,N_2464,N_914);
nor U5238 (N_5238,N_4974,N_2185);
or U5239 (N_5239,N_3736,N_4112);
nor U5240 (N_5240,N_985,N_3564);
xnor U5241 (N_5241,N_3526,N_3226);
nor U5242 (N_5242,N_1968,N_3454);
nor U5243 (N_5243,N_4925,N_2071);
nand U5244 (N_5244,N_1866,N_333);
nand U5245 (N_5245,N_1317,N_1876);
nand U5246 (N_5246,N_698,N_31);
or U5247 (N_5247,N_4337,N_4197);
and U5248 (N_5248,N_2266,N_325);
or U5249 (N_5249,N_4313,N_906);
nand U5250 (N_5250,N_623,N_1430);
nor U5251 (N_5251,N_4145,N_2545);
or U5252 (N_5252,N_1659,N_3748);
nor U5253 (N_5253,N_833,N_2372);
nor U5254 (N_5254,N_4938,N_2848);
or U5255 (N_5255,N_1966,N_2627);
xnor U5256 (N_5256,N_1238,N_3926);
or U5257 (N_5257,N_2099,N_1905);
nand U5258 (N_5258,N_384,N_2701);
nor U5259 (N_5259,N_3600,N_4833);
xor U5260 (N_5260,N_2887,N_1934);
or U5261 (N_5261,N_4893,N_889);
nand U5262 (N_5262,N_2841,N_4997);
nand U5263 (N_5263,N_1902,N_1343);
and U5264 (N_5264,N_3370,N_2822);
and U5265 (N_5265,N_4922,N_4789);
nor U5266 (N_5266,N_2652,N_2619);
nor U5267 (N_5267,N_4353,N_3368);
nor U5268 (N_5268,N_989,N_542);
xnor U5269 (N_5269,N_3079,N_2600);
nand U5270 (N_5270,N_714,N_617);
xor U5271 (N_5271,N_4683,N_1262);
and U5272 (N_5272,N_2562,N_343);
or U5273 (N_5273,N_3827,N_4410);
nand U5274 (N_5274,N_710,N_1269);
nor U5275 (N_5275,N_3119,N_4827);
and U5276 (N_5276,N_413,N_3961);
or U5277 (N_5277,N_931,N_4111);
or U5278 (N_5278,N_636,N_4868);
or U5279 (N_5279,N_1323,N_3693);
or U5280 (N_5280,N_2749,N_2191);
nor U5281 (N_5281,N_4864,N_2215);
nor U5282 (N_5282,N_605,N_2349);
nor U5283 (N_5283,N_4030,N_4758);
and U5284 (N_5284,N_2550,N_1815);
or U5285 (N_5285,N_610,N_4883);
and U5286 (N_5286,N_972,N_338);
nand U5287 (N_5287,N_786,N_2499);
xor U5288 (N_5288,N_2288,N_1030);
xor U5289 (N_5289,N_129,N_2552);
or U5290 (N_5290,N_1889,N_2416);
xor U5291 (N_5291,N_1324,N_4070);
nor U5292 (N_5292,N_1551,N_1730);
or U5293 (N_5293,N_4722,N_4273);
xor U5294 (N_5294,N_2985,N_2660);
or U5295 (N_5295,N_794,N_707);
nor U5296 (N_5296,N_3547,N_4442);
nor U5297 (N_5297,N_2576,N_1668);
nor U5298 (N_5298,N_3646,N_732);
nand U5299 (N_5299,N_3404,N_2549);
nor U5300 (N_5300,N_1803,N_4487);
xnor U5301 (N_5301,N_2316,N_4008);
and U5302 (N_5302,N_4587,N_2540);
xnor U5303 (N_5303,N_4393,N_1536);
and U5304 (N_5304,N_303,N_4207);
nand U5305 (N_5305,N_1334,N_4681);
or U5306 (N_5306,N_4288,N_3395);
nand U5307 (N_5307,N_4854,N_1615);
and U5308 (N_5308,N_4164,N_3569);
or U5309 (N_5309,N_1991,N_1163);
and U5310 (N_5310,N_538,N_1435);
xor U5311 (N_5311,N_3445,N_3672);
and U5312 (N_5312,N_497,N_4004);
nor U5313 (N_5313,N_4115,N_2321);
or U5314 (N_5314,N_4027,N_3338);
nand U5315 (N_5315,N_2704,N_1681);
nand U5316 (N_5316,N_544,N_2132);
xor U5317 (N_5317,N_2513,N_1042);
or U5318 (N_5318,N_1886,N_3792);
and U5319 (N_5319,N_473,N_2251);
or U5320 (N_5320,N_3810,N_3383);
and U5321 (N_5321,N_173,N_4753);
xnor U5322 (N_5322,N_997,N_4417);
nand U5323 (N_5323,N_1466,N_4061);
nor U5324 (N_5324,N_2586,N_1500);
or U5325 (N_5325,N_3747,N_1402);
and U5326 (N_5326,N_1205,N_3754);
nand U5327 (N_5327,N_1613,N_2351);
nand U5328 (N_5328,N_4165,N_1186);
nand U5329 (N_5329,N_2894,N_3901);
and U5330 (N_5330,N_1479,N_1506);
nand U5331 (N_5331,N_4235,N_1308);
xor U5332 (N_5332,N_4269,N_2598);
and U5333 (N_5333,N_155,N_411);
or U5334 (N_5334,N_4158,N_2802);
xnor U5335 (N_5335,N_3249,N_1047);
nand U5336 (N_5336,N_4814,N_1004);
or U5337 (N_5337,N_720,N_276);
and U5338 (N_5338,N_1396,N_269);
nor U5339 (N_5339,N_2669,N_4841);
nor U5340 (N_5340,N_1351,N_2681);
nand U5341 (N_5341,N_4981,N_2012);
xnor U5342 (N_5342,N_516,N_3013);
nor U5343 (N_5343,N_1394,N_4493);
nor U5344 (N_5344,N_1677,N_1418);
nand U5345 (N_5345,N_2214,N_3277);
or U5346 (N_5346,N_1784,N_4649);
and U5347 (N_5347,N_3607,N_1679);
and U5348 (N_5348,N_639,N_4218);
xnor U5349 (N_5349,N_2972,N_326);
nand U5350 (N_5350,N_4364,N_528);
nor U5351 (N_5351,N_4163,N_3020);
xnor U5352 (N_5352,N_3550,N_3702);
nor U5353 (N_5353,N_2468,N_1589);
and U5354 (N_5354,N_4071,N_683);
and U5355 (N_5355,N_2968,N_2914);
nor U5356 (N_5356,N_3453,N_366);
nor U5357 (N_5357,N_1959,N_390);
or U5358 (N_5358,N_1879,N_1462);
xor U5359 (N_5359,N_408,N_4921);
and U5360 (N_5360,N_4932,N_3613);
nor U5361 (N_5361,N_2873,N_419);
and U5362 (N_5362,N_3387,N_3228);
nor U5363 (N_5363,N_2409,N_894);
or U5364 (N_5364,N_2547,N_4862);
or U5365 (N_5365,N_171,N_3397);
xnor U5366 (N_5366,N_1245,N_1405);
xor U5367 (N_5367,N_1237,N_1731);
or U5368 (N_5368,N_4427,N_3947);
or U5369 (N_5369,N_1477,N_1292);
and U5370 (N_5370,N_4695,N_1977);
nor U5371 (N_5371,N_4063,N_1287);
or U5372 (N_5372,N_3417,N_132);
or U5373 (N_5373,N_3798,N_4042);
nand U5374 (N_5374,N_2695,N_3134);
nand U5375 (N_5375,N_317,N_1367);
nor U5376 (N_5376,N_3603,N_1031);
nand U5377 (N_5377,N_711,N_3329);
nor U5378 (N_5378,N_2269,N_890);
xnor U5379 (N_5379,N_236,N_3279);
nand U5380 (N_5380,N_130,N_4942);
nor U5381 (N_5381,N_2756,N_4840);
xnor U5382 (N_5382,N_4102,N_2665);
xor U5383 (N_5383,N_4182,N_1152);
nand U5384 (N_5384,N_4711,N_4598);
or U5385 (N_5385,N_996,N_4955);
xor U5386 (N_5386,N_4001,N_2608);
xor U5387 (N_5387,N_3596,N_3301);
nor U5388 (N_5388,N_4650,N_2249);
and U5389 (N_5389,N_135,N_2521);
nor U5390 (N_5390,N_3706,N_3041);
nand U5391 (N_5391,N_3496,N_1582);
or U5392 (N_5392,N_2834,N_1107);
nand U5393 (N_5393,N_4706,N_3973);
or U5394 (N_5394,N_1655,N_4250);
and U5395 (N_5395,N_1638,N_2899);
nand U5396 (N_5396,N_963,N_3394);
nor U5397 (N_5397,N_396,N_1676);
xnor U5398 (N_5398,N_4021,N_2141);
and U5399 (N_5399,N_1765,N_3407);
or U5400 (N_5400,N_3421,N_1303);
xnor U5401 (N_5401,N_2696,N_1557);
and U5402 (N_5402,N_4880,N_3932);
nand U5403 (N_5403,N_4091,N_1064);
and U5404 (N_5404,N_3839,N_106);
xor U5405 (N_5405,N_4469,N_2989);
nor U5406 (N_5406,N_2967,N_2001);
xnor U5407 (N_5407,N_2698,N_940);
or U5408 (N_5408,N_1310,N_3439);
and U5409 (N_5409,N_4432,N_3559);
or U5410 (N_5410,N_1176,N_2710);
nand U5411 (N_5411,N_4206,N_4597);
and U5412 (N_5412,N_1428,N_4119);
and U5413 (N_5413,N_638,N_1743);
nand U5414 (N_5414,N_674,N_485);
xnor U5415 (N_5415,N_2859,N_1312);
xnor U5416 (N_5416,N_871,N_2281);
nand U5417 (N_5417,N_3674,N_4750);
or U5418 (N_5418,N_4563,N_4324);
nor U5419 (N_5419,N_837,N_1087);
and U5420 (N_5420,N_4629,N_3103);
nor U5421 (N_5421,N_2566,N_1389);
nor U5422 (N_5422,N_2119,N_440);
nor U5423 (N_5423,N_3843,N_4982);
or U5424 (N_5424,N_1456,N_681);
or U5425 (N_5425,N_4510,N_265);
or U5426 (N_5426,N_4610,N_3220);
and U5427 (N_5427,N_2623,N_4638);
nor U5428 (N_5428,N_653,N_922);
nand U5429 (N_5429,N_4672,N_1943);
nand U5430 (N_5430,N_2982,N_2729);
and U5431 (N_5431,N_1896,N_3819);
nand U5432 (N_5432,N_2418,N_2159);
nand U5433 (N_5433,N_117,N_4294);
nor U5434 (N_5434,N_2166,N_266);
nor U5435 (N_5435,N_4669,N_1660);
xnor U5436 (N_5436,N_1740,N_263);
nor U5437 (N_5437,N_1947,N_4511);
xnor U5438 (N_5438,N_3632,N_4998);
nor U5439 (N_5439,N_629,N_4799);
nand U5440 (N_5440,N_1138,N_3187);
or U5441 (N_5441,N_4249,N_4964);
or U5442 (N_5442,N_3434,N_1062);
nand U5443 (N_5443,N_3900,N_3316);
or U5444 (N_5444,N_1273,N_1982);
xnor U5445 (N_5445,N_1653,N_4136);
or U5446 (N_5446,N_3518,N_2788);
nor U5447 (N_5447,N_644,N_1020);
and U5448 (N_5448,N_2206,N_86);
nor U5449 (N_5449,N_496,N_4320);
xor U5450 (N_5450,N_715,N_4362);
and U5451 (N_5451,N_2579,N_1483);
or U5452 (N_5452,N_4892,N_2285);
or U5453 (N_5453,N_3012,N_920);
nor U5454 (N_5454,N_700,N_3919);
xor U5455 (N_5455,N_2651,N_1207);
xnor U5456 (N_5456,N_71,N_1233);
or U5457 (N_5457,N_3837,N_1620);
xor U5458 (N_5458,N_1344,N_392);
nor U5459 (N_5459,N_3806,N_756);
nand U5460 (N_5460,N_3356,N_4051);
xnor U5461 (N_5461,N_4512,N_1856);
nor U5462 (N_5462,N_283,N_572);
nand U5463 (N_5463,N_843,N_2174);
nand U5464 (N_5464,N_19,N_2925);
nor U5465 (N_5465,N_3222,N_4352);
or U5466 (N_5466,N_1480,N_4037);
and U5467 (N_5467,N_4636,N_2525);
or U5468 (N_5468,N_2135,N_105);
xor U5469 (N_5469,N_4576,N_2052);
or U5470 (N_5470,N_3211,N_2447);
and U5471 (N_5471,N_1295,N_179);
and U5472 (N_5472,N_2158,N_1680);
xnor U5473 (N_5473,N_3785,N_52);
and U5474 (N_5474,N_1413,N_2903);
nor U5475 (N_5475,N_1658,N_4256);
or U5476 (N_5476,N_3848,N_1039);
nor U5477 (N_5477,N_3219,N_4898);
nand U5478 (N_5478,N_802,N_4159);
xor U5479 (N_5479,N_3667,N_1449);
nand U5480 (N_5480,N_2307,N_2897);
xor U5481 (N_5481,N_1807,N_3411);
nand U5482 (N_5482,N_4590,N_438);
and U5483 (N_5483,N_2758,N_3174);
nor U5484 (N_5484,N_1306,N_1549);
nand U5485 (N_5485,N_1828,N_520);
nand U5486 (N_5486,N_4335,N_3351);
and U5487 (N_5487,N_607,N_1559);
and U5488 (N_5488,N_1037,N_693);
xnor U5489 (N_5489,N_1484,N_2192);
nand U5490 (N_5490,N_101,N_4334);
xor U5491 (N_5491,N_4009,N_254);
or U5492 (N_5492,N_2332,N_1486);
xor U5493 (N_5493,N_3728,N_1387);
nor U5494 (N_5494,N_4141,N_335);
xor U5495 (N_5495,N_1327,N_2329);
and U5496 (N_5496,N_4093,N_1050);
and U5497 (N_5497,N_3449,N_3078);
nor U5498 (N_5498,N_441,N_1542);
xnor U5499 (N_5499,N_3199,N_14);
nand U5500 (N_5500,N_4449,N_509);
nand U5501 (N_5501,N_3887,N_3953);
nor U5502 (N_5502,N_1594,N_564);
or U5503 (N_5503,N_1395,N_717);
or U5504 (N_5504,N_3451,N_1450);
nand U5505 (N_5505,N_897,N_467);
and U5506 (N_5506,N_2716,N_4223);
xnor U5507 (N_5507,N_1423,N_2581);
and U5508 (N_5508,N_3247,N_1642);
and U5509 (N_5509,N_4867,N_2979);
nand U5510 (N_5510,N_4302,N_2051);
nor U5511 (N_5511,N_701,N_1626);
nor U5512 (N_5512,N_3274,N_1540);
and U5513 (N_5513,N_1504,N_2855);
xnor U5514 (N_5514,N_3957,N_1116);
xnor U5515 (N_5515,N_472,N_2204);
nand U5516 (N_5516,N_4342,N_2938);
or U5517 (N_5517,N_812,N_4891);
xnor U5518 (N_5518,N_523,N_2530);
xor U5519 (N_5519,N_2303,N_733);
or U5520 (N_5520,N_4227,N_3125);
nand U5521 (N_5521,N_3694,N_3535);
or U5522 (N_5522,N_1377,N_1572);
nand U5523 (N_5523,N_4041,N_2978);
nand U5524 (N_5524,N_3139,N_4381);
nand U5525 (N_5525,N_1685,N_3396);
nor U5526 (N_5526,N_4140,N_4966);
xor U5527 (N_5527,N_3808,N_846);
and U5528 (N_5528,N_315,N_2246);
xor U5529 (N_5529,N_2318,N_3478);
xnor U5530 (N_5530,N_508,N_797);
and U5531 (N_5531,N_2924,N_2768);
nand U5532 (N_5532,N_1044,N_1251);
or U5533 (N_5533,N_2105,N_1045);
nor U5534 (N_5534,N_4878,N_729);
xor U5535 (N_5535,N_3830,N_2599);
or U5536 (N_5536,N_741,N_4287);
xnor U5537 (N_5537,N_954,N_4884);
or U5538 (N_5538,N_3800,N_3160);
nand U5539 (N_5539,N_2224,N_1929);
or U5540 (N_5540,N_3150,N_3776);
or U5541 (N_5541,N_4482,N_3624);
xnor U5542 (N_5542,N_4723,N_3783);
or U5543 (N_5543,N_4961,N_4734);
and U5544 (N_5544,N_2004,N_3841);
and U5545 (N_5545,N_646,N_3371);
nor U5546 (N_5546,N_793,N_1165);
xor U5547 (N_5547,N_3323,N_4771);
or U5548 (N_5548,N_3130,N_4317);
and U5549 (N_5549,N_1012,N_4178);
xor U5550 (N_5550,N_4029,N_534);
nand U5551 (N_5551,N_1422,N_1195);
and U5552 (N_5552,N_3005,N_2568);
xnor U5553 (N_5553,N_2759,N_4620);
nor U5554 (N_5554,N_115,N_2429);
and U5555 (N_5555,N_1465,N_3935);
and U5556 (N_5556,N_768,N_3047);
nor U5557 (N_5557,N_1663,N_3376);
or U5558 (N_5558,N_1887,N_1501);
nor U5559 (N_5559,N_3031,N_1957);
xnor U5560 (N_5560,N_856,N_4881);
or U5561 (N_5561,N_1733,N_747);
or U5562 (N_5562,N_1616,N_2676);
nand U5563 (N_5563,N_4917,N_2272);
xnor U5564 (N_5564,N_965,N_2531);
nor U5565 (N_5565,N_2352,N_3683);
nand U5566 (N_5566,N_2178,N_2849);
xnor U5567 (N_5567,N_3513,N_455);
nor U5568 (N_5568,N_3061,N_1839);
nand U5569 (N_5569,N_2907,N_3230);
or U5570 (N_5570,N_2487,N_4185);
xor U5571 (N_5571,N_3690,N_1742);
or U5572 (N_5572,N_773,N_4808);
xor U5573 (N_5573,N_4621,N_2913);
and U5574 (N_5574,N_910,N_3141);
or U5575 (N_5575,N_164,N_3958);
and U5576 (N_5576,N_4243,N_3214);
or U5577 (N_5577,N_1918,N_184);
nand U5578 (N_5578,N_4356,N_1494);
and U5579 (N_5579,N_3580,N_1569);
and U5580 (N_5580,N_2891,N_1651);
nand U5581 (N_5581,N_32,N_1162);
or U5582 (N_5582,N_133,N_4623);
nor U5583 (N_5583,N_4570,N_2678);
or U5584 (N_5584,N_3871,N_203);
xnor U5585 (N_5585,N_4224,N_4896);
xnor U5586 (N_5586,N_4945,N_4048);
and U5587 (N_5587,N_1285,N_4390);
and U5588 (N_5588,N_2864,N_2036);
or U5589 (N_5589,N_1812,N_2850);
nand U5590 (N_5590,N_3198,N_3414);
nand U5591 (N_5591,N_4023,N_1191);
xnor U5592 (N_5592,N_4525,N_4067);
xor U5593 (N_5593,N_2143,N_1442);
or U5594 (N_5594,N_1843,N_136);
nand U5595 (N_5595,N_1124,N_3987);
and U5596 (N_5596,N_1768,N_1133);
and U5597 (N_5597,N_1333,N_565);
xnor U5598 (N_5598,N_1782,N_4617);
or U5599 (N_5599,N_1931,N_883);
or U5600 (N_5600,N_4019,N_4355);
nand U5601 (N_5601,N_3701,N_923);
and U5602 (N_5602,N_4376,N_1632);
or U5603 (N_5603,N_3098,N_782);
nand U5604 (N_5604,N_2870,N_2647);
and U5605 (N_5605,N_982,N_3595);
and U5606 (N_5606,N_3458,N_950);
nand U5607 (N_5607,N_3671,N_962);
nor U5608 (N_5608,N_807,N_284);
or U5609 (N_5609,N_1944,N_3309);
and U5610 (N_5610,N_4120,N_2555);
nor U5611 (N_5611,N_3071,N_1758);
nand U5612 (N_5612,N_746,N_2910);
and U5613 (N_5613,N_2575,N_4044);
nand U5614 (N_5614,N_215,N_1635);
and U5615 (N_5615,N_2398,N_1618);
xor U5616 (N_5616,N_1211,N_112);
nand U5617 (N_5617,N_1714,N_3593);
and U5618 (N_5618,N_3620,N_2255);
nand U5619 (N_5619,N_2361,N_1411);
xor U5620 (N_5620,N_805,N_879);
xor U5621 (N_5621,N_3528,N_2699);
xor U5622 (N_5622,N_2718,N_322);
and U5623 (N_5623,N_1527,N_69);
or U5624 (N_5624,N_358,N_499);
and U5625 (N_5625,N_3193,N_1872);
nand U5626 (N_5626,N_1951,N_4873);
or U5627 (N_5627,N_4796,N_670);
nand U5628 (N_5628,N_3032,N_4279);
xnor U5629 (N_5629,N_1975,N_4693);
nor U5630 (N_5630,N_3362,N_2455);
xnor U5631 (N_5631,N_2536,N_1586);
nand U5632 (N_5632,N_3003,N_2779);
nand U5633 (N_5633,N_2715,N_4916);
nor U5634 (N_5634,N_1898,N_4242);
or U5635 (N_5635,N_4199,N_1532);
nand U5636 (N_5636,N_4385,N_144);
xnor U5637 (N_5637,N_4129,N_35);
nand U5638 (N_5638,N_1170,N_1535);
xor U5639 (N_5639,N_1916,N_1041);
nor U5640 (N_5640,N_1764,N_2195);
or U5641 (N_5641,N_361,N_4451);
or U5642 (N_5642,N_1490,N_775);
nor U5643 (N_5643,N_493,N_3485);
xor U5644 (N_5644,N_1855,N_2428);
nand U5645 (N_5645,N_2557,N_1656);
and U5646 (N_5646,N_731,N_3805);
and U5647 (N_5647,N_4173,N_474);
nor U5648 (N_5648,N_2112,N_4679);
xnor U5649 (N_5649,N_4543,N_1756);
nand U5650 (N_5650,N_2686,N_3952);
and U5651 (N_5651,N_3173,N_1103);
or U5652 (N_5652,N_841,N_1788);
nand U5653 (N_5653,N_1065,N_3538);
nor U5654 (N_5654,N_1369,N_2074);
nand U5655 (N_5655,N_4370,N_3618);
nand U5656 (N_5656,N_4518,N_4489);
nand U5657 (N_5657,N_2607,N_3491);
and U5658 (N_5658,N_4909,N_2929);
or U5659 (N_5659,N_4962,N_569);
nand U5660 (N_5660,N_864,N_2173);
nor U5661 (N_5661,N_1019,N_1596);
nor U5662 (N_5662,N_1096,N_2565);
and U5663 (N_5663,N_139,N_1664);
and U5664 (N_5664,N_1852,N_2535);
xnor U5665 (N_5665,N_4107,N_4359);
xor U5666 (N_5666,N_3202,N_568);
xnor U5667 (N_5667,N_1154,N_43);
nor U5668 (N_5668,N_2328,N_1332);
or U5669 (N_5669,N_4772,N_3764);
and U5670 (N_5670,N_2302,N_2011);
nor U5671 (N_5671,N_992,N_26);
or U5672 (N_5672,N_1137,N_4531);
and U5673 (N_5673,N_3553,N_97);
xor U5674 (N_5674,N_4316,N_4210);
nand U5675 (N_5675,N_3291,N_4910);
nor U5676 (N_5676,N_3037,N_207);
xnor U5677 (N_5677,N_2996,N_3241);
nand U5678 (N_5678,N_4074,N_1591);
nor U5679 (N_5679,N_1290,N_2601);
nand U5680 (N_5680,N_574,N_2572);
nor U5681 (N_5681,N_4990,N_312);
xnor U5682 (N_5682,N_2262,N_4080);
xor U5683 (N_5683,N_3359,N_2824);
nand U5684 (N_5684,N_1429,N_222);
nand U5685 (N_5685,N_4123,N_2767);
nand U5686 (N_5686,N_3059,N_409);
or U5687 (N_5687,N_2053,N_4321);
nand U5688 (N_5688,N_3920,N_2939);
nor U5689 (N_5689,N_3983,N_3746);
xor U5690 (N_5690,N_4099,N_650);
and U5691 (N_5691,N_1923,N_3344);
xor U5692 (N_5692,N_744,N_2675);
nor U5693 (N_5693,N_1754,N_3649);
xnor U5694 (N_5694,N_4,N_2928);
and U5695 (N_5695,N_561,N_4712);
or U5696 (N_5696,N_2187,N_166);
and U5697 (N_5697,N_1260,N_4038);
xor U5698 (N_5698,N_400,N_4105);
and U5699 (N_5699,N_4373,N_522);
xnor U5700 (N_5700,N_2958,N_2179);
xnor U5701 (N_5701,N_3379,N_3794);
xnor U5702 (N_5702,N_2606,N_2636);
xnor U5703 (N_5703,N_4686,N_868);
or U5704 (N_5704,N_1888,N_1606);
and U5705 (N_5705,N_2046,N_2799);
and U5706 (N_5706,N_4812,N_1398);
or U5707 (N_5707,N_4467,N_761);
nand U5708 (N_5708,N_2437,N_407);
and U5709 (N_5709,N_4319,N_1272);
xnor U5710 (N_5710,N_3204,N_1487);
xnor U5711 (N_5711,N_3766,N_3054);
nand U5712 (N_5712,N_1346,N_1830);
nand U5713 (N_5713,N_2064,N_4828);
xnor U5714 (N_5714,N_3302,N_1734);
xnor U5715 (N_5715,N_3578,N_694);
nor U5716 (N_5716,N_902,N_4804);
or U5717 (N_5717,N_2697,N_2305);
and U5718 (N_5718,N_2021,N_4267);
or U5719 (N_5719,N_873,N_3727);
xor U5720 (N_5720,N_1827,N_1578);
and U5721 (N_5721,N_1646,N_116);
and U5722 (N_5722,N_2311,N_2901);
and U5723 (N_5723,N_505,N_2946);
xor U5724 (N_5724,N_4005,N_4568);
nand U5725 (N_5725,N_2746,N_3633);
nor U5726 (N_5726,N_2100,N_925);
xnor U5727 (N_5727,N_4544,N_3902);
or U5728 (N_5728,N_4124,N_4546);
and U5729 (N_5729,N_3602,N_675);
nand U5730 (N_5730,N_3738,N_4776);
xor U5731 (N_5731,N_2275,N_2911);
and U5732 (N_5732,N_4970,N_3717);
or U5733 (N_5733,N_4398,N_4694);
nor U5734 (N_5734,N_481,N_2120);
or U5735 (N_5735,N_1645,N_3412);
or U5736 (N_5736,N_107,N_4825);
and U5737 (N_5737,N_4731,N_1320);
xor U5738 (N_5738,N_1453,N_3849);
or U5739 (N_5739,N_1654,N_3517);
or U5740 (N_5740,N_4428,N_3579);
nand U5741 (N_5741,N_4457,N_3777);
xor U5742 (N_5742,N_4494,N_2926);
nor U5743 (N_5743,N_1729,N_3850);
xor U5744 (N_5744,N_4465,N_3734);
nor U5745 (N_5745,N_3943,N_4006);
nor U5746 (N_5746,N_2126,N_464);
and U5747 (N_5747,N_2986,N_1766);
or U5748 (N_5748,N_4582,N_2200);
xor U5749 (N_5749,N_1859,N_1917);
nor U5750 (N_5750,N_3616,N_867);
or U5751 (N_5751,N_429,N_678);
or U5752 (N_5752,N_3730,N_4996);
xor U5753 (N_5753,N_3537,N_1058);
xnor U5754 (N_5754,N_1197,N_2796);
xnor U5755 (N_5755,N_180,N_1289);
nand U5756 (N_5756,N_3117,N_2331);
nor U5757 (N_5757,N_2003,N_480);
nand U5758 (N_5758,N_1051,N_3677);
xnor U5759 (N_5759,N_2374,N_281);
nor U5760 (N_5760,N_4378,N_4947);
nor U5761 (N_5761,N_3700,N_3691);
xnor U5762 (N_5762,N_216,N_2091);
xnor U5763 (N_5763,N_4214,N_1008);
nor U5764 (N_5764,N_4823,N_4139);
or U5765 (N_5765,N_3287,N_4456);
or U5766 (N_5766,N_2617,N_2376);
and U5767 (N_5767,N_3322,N_2820);
nor U5768 (N_5768,N_3907,N_486);
and U5769 (N_5769,N_1003,N_4113);
and U5770 (N_5770,N_810,N_4550);
or U5771 (N_5771,N_4272,N_330);
or U5772 (N_5772,N_258,N_4371);
nand U5773 (N_5773,N_3209,N_4160);
xor U5774 (N_5774,N_4281,N_1814);
or U5775 (N_5775,N_2054,N_2017);
and U5776 (N_5776,N_1811,N_706);
xor U5777 (N_5777,N_170,N_2056);
and U5778 (N_5778,N_202,N_1089);
and U5779 (N_5779,N_3502,N_4800);
or U5780 (N_5780,N_2632,N_4547);
nand U5781 (N_5781,N_506,N_809);
or U5782 (N_5782,N_2854,N_4874);
xnor U5783 (N_5783,N_3661,N_2063);
nand U5784 (N_5784,N_1371,N_4791);
nor U5785 (N_5785,N_308,N_10);
nor U5786 (N_5786,N_4565,N_4713);
xor U5787 (N_5787,N_4162,N_1531);
xor U5788 (N_5788,N_1229,N_1585);
nand U5789 (N_5789,N_3324,N_401);
or U5790 (N_5790,N_160,N_4834);
and U5791 (N_5791,N_3456,N_1792);
or U5792 (N_5792,N_755,N_3804);
and U5793 (N_5793,N_4408,N_2390);
nor U5794 (N_5794,N_47,N_4154);
nand U5795 (N_5795,N_494,N_4179);
or U5796 (N_5796,N_1526,N_3081);
nor U5797 (N_5797,N_1567,N_3196);
xor U5798 (N_5798,N_2635,N_4897);
or U5799 (N_5799,N_4170,N_3729);
or U5800 (N_5800,N_512,N_1457);
and U5801 (N_5801,N_1777,N_908);
nor U5802 (N_5802,N_4783,N_1499);
and U5803 (N_5803,N_2475,N_4631);
or U5804 (N_5804,N_2345,N_2181);
xor U5805 (N_5805,N_2900,N_781);
and U5806 (N_5806,N_3975,N_4863);
and U5807 (N_5807,N_1507,N_3972);
nand U5808 (N_5808,N_2236,N_3642);
nand U5809 (N_5809,N_2066,N_899);
and U5810 (N_5810,N_2165,N_2748);
xor U5811 (N_5811,N_3908,N_2714);
and U5812 (N_5812,N_3200,N_3494);
nor U5813 (N_5813,N_4801,N_1048);
nor U5814 (N_5814,N_648,N_4664);
nand U5815 (N_5815,N_3331,N_3861);
xnor U5816 (N_5816,N_4882,N_2529);
nand U5817 (N_5817,N_1562,N_4727);
nor U5818 (N_5818,N_3782,N_1482);
and U5819 (N_5819,N_4252,N_531);
nor U5820 (N_5820,N_4702,N_1027);
and U5821 (N_5821,N_304,N_2567);
nor U5822 (N_5822,N_1698,N_1106);
nand U5823 (N_5823,N_1688,N_4541);
nor U5824 (N_5824,N_1034,N_4759);
nand U5825 (N_5825,N_1796,N_1716);
or U5826 (N_5826,N_1194,N_4480);
xnor U5827 (N_5827,N_4992,N_4509);
nor U5828 (N_5828,N_2223,N_4400);
xor U5829 (N_5829,N_3131,N_3194);
nand U5830 (N_5830,N_4533,N_292);
nor U5831 (N_5831,N_1514,N_175);
or U5832 (N_5832,N_3087,N_4034);
xnor U5833 (N_5833,N_1090,N_4485);
nor U5834 (N_5834,N_4901,N_2320);
or U5835 (N_5835,N_1322,N_3066);
xor U5836 (N_5836,N_4228,N_1848);
xor U5837 (N_5837,N_4188,N_2084);
or U5838 (N_5838,N_1577,N_2239);
xnor U5839 (N_5839,N_380,N_3934);
nand U5840 (N_5840,N_652,N_998);
and U5841 (N_5841,N_2271,N_383);
and U5842 (N_5842,N_4696,N_3077);
or U5843 (N_5843,N_4599,N_938);
xnor U5844 (N_5844,N_1675,N_2639);
xnor U5845 (N_5845,N_3183,N_3847);
or U5846 (N_5846,N_1621,N_1622);
nand U5847 (N_5847,N_3481,N_4262);
or U5848 (N_5848,N_4716,N_677);
nand U5849 (N_5849,N_4946,N_4153);
xor U5850 (N_5850,N_2070,N_3057);
nand U5851 (N_5851,N_2424,N_2116);
nand U5852 (N_5852,N_2493,N_1189);
nand U5853 (N_5853,N_206,N_3191);
xnor U5854 (N_5854,N_2964,N_3243);
or U5855 (N_5855,N_4586,N_4251);
nor U5856 (N_5856,N_2886,N_4392);
or U5857 (N_5857,N_2892,N_1503);
xor U5858 (N_5858,N_1518,N_2106);
nand U5859 (N_5859,N_291,N_592);
and U5860 (N_5860,N_2484,N_4025);
nand U5861 (N_5861,N_4677,N_4468);
nand U5862 (N_5862,N_4850,N_4028);
nor U5863 (N_5863,N_3834,N_2378);
nor U5864 (N_5864,N_1967,N_3339);
or U5865 (N_5865,N_3448,N_826);
nand U5866 (N_5866,N_3911,N_679);
xor U5867 (N_5867,N_150,N_3227);
xnor U5868 (N_5868,N_3879,N_2920);
nand U5869 (N_5869,N_3854,N_885);
and U5870 (N_5870,N_3767,N_1391);
nor U5871 (N_5871,N_2644,N_4059);
nor U5872 (N_5872,N_2837,N_4049);
or U5873 (N_5873,N_3929,N_2121);
nand U5874 (N_5874,N_3899,N_4058);
and U5875 (N_5875,N_3285,N_4062);
or U5876 (N_5876,N_3874,N_792);
nand U5877 (N_5877,N_688,N_4887);
nand U5878 (N_5878,N_4078,N_2379);
or U5879 (N_5879,N_3529,N_4089);
and U5880 (N_5880,N_1583,N_2588);
and U5881 (N_5881,N_3375,N_1241);
nand U5882 (N_5882,N_3489,N_1563);
xor U5883 (N_5883,N_4611,N_3479);
nand U5884 (N_5884,N_872,N_4953);
or U5885 (N_5885,N_53,N_332);
nand U5886 (N_5886,N_81,N_832);
or U5887 (N_5887,N_1800,N_4022);
xnor U5888 (N_5888,N_3960,N_4741);
or U5889 (N_5889,N_3266,N_990);
xnor U5890 (N_5890,N_3318,N_2517);
nand U5891 (N_5891,N_2877,N_2161);
and U5892 (N_5892,N_772,N_659);
or U5893 (N_5893,N_4394,N_3965);
and U5894 (N_5894,N_3844,N_738);
or U5895 (N_5895,N_1910,N_3656);
xor U5896 (N_5896,N_3039,N_2093);
or U5897 (N_5897,N_1804,N_3662);
nand U5898 (N_5898,N_791,N_61);
or U5899 (N_5899,N_4295,N_4668);
or U5900 (N_5900,N_3298,N_2038);
xor U5901 (N_5901,N_3991,N_576);
xor U5902 (N_5902,N_3731,N_4902);
xor U5903 (N_5903,N_3687,N_4088);
nand U5904 (N_5904,N_4375,N_4680);
nor U5905 (N_5905,N_417,N_2630);
xor U5906 (N_5906,N_297,N_3345);
nand U5907 (N_5907,N_3863,N_3857);
nor U5908 (N_5908,N_2732,N_3790);
xnor U5909 (N_5909,N_854,N_4360);
or U5910 (N_5910,N_1349,N_4198);
nand U5911 (N_5911,N_560,N_3964);
nor U5912 (N_5912,N_3561,N_4819);
nor U5913 (N_5913,N_1266,N_543);
or U5914 (N_5914,N_436,N_4338);
and U5915 (N_5915,N_3562,N_1546);
nor U5916 (N_5916,N_1304,N_2014);
nand U5917 (N_5917,N_126,N_3477);
and U5918 (N_5918,N_783,N_699);
and U5919 (N_5919,N_2009,N_3923);
nand U5920 (N_5920,N_3400,N_296);
and U5921 (N_5921,N_4146,N_944);
nand U5922 (N_5922,N_4633,N_3034);
xor U5923 (N_5923,N_1408,N_2047);
nand U5924 (N_5924,N_2738,N_4756);
nand U5925 (N_5925,N_1703,N_2340);
nand U5926 (N_5926,N_2337,N_4332);
nand U5927 (N_5927,N_3889,N_3765);
and U5928 (N_5928,N_949,N_4632);
or U5929 (N_5929,N_2377,N_4630);
or U5930 (N_5930,N_3292,N_3231);
nand U5931 (N_5931,N_1066,N_2284);
and U5932 (N_5932,N_726,N_1552);
nor U5933 (N_5933,N_2720,N_4296);
xor U5934 (N_5934,N_816,N_3914);
nand U5935 (N_5935,N_1834,N_1410);
nand U5936 (N_5936,N_1473,N_2258);
and U5937 (N_5937,N_4913,N_435);
nor U5938 (N_5938,N_385,N_391);
nor U5939 (N_5939,N_238,N_4836);
nand U5940 (N_5940,N_4073,N_4717);
xnor U5941 (N_5941,N_3832,N_1631);
or U5942 (N_5942,N_1780,N_2862);
or U5943 (N_5943,N_4665,N_2277);
xnor U5944 (N_5944,N_2427,N_3284);
xor U5945 (N_5945,N_3623,N_1819);
nand U5946 (N_5946,N_3460,N_2797);
and U5947 (N_5947,N_2750,N_244);
or U5948 (N_5948,N_3470,N_3733);
nor U5949 (N_5949,N_1995,N_2290);
nor U5950 (N_5950,N_2144,N_4504);
xnor U5951 (N_5951,N_2785,N_4127);
nand U5952 (N_5952,N_3676,N_2584);
nand U5953 (N_5953,N_3252,N_147);
xnor U5954 (N_5954,N_1954,N_3577);
nand U5955 (N_5955,N_4203,N_488);
or U5956 (N_5956,N_4682,N_2957);
nor U5957 (N_5957,N_4109,N_1074);
nand U5958 (N_5958,N_2819,N_1156);
nor U5959 (N_5959,N_4122,N_1206);
and U5960 (N_5960,N_3281,N_1427);
nand U5961 (N_5961,N_477,N_1860);
nor U5962 (N_5962,N_616,N_609);
and U5963 (N_5963,N_3637,N_4380);
or U5964 (N_5964,N_2702,N_323);
nand U5965 (N_5965,N_4733,N_4167);
nor U5966 (N_5966,N_2292,N_785);
or U5967 (N_5967,N_2615,N_2417);
xor U5968 (N_5968,N_3922,N_1140);
xor U5969 (N_5969,N_1537,N_3866);
and U5970 (N_5970,N_2172,N_835);
xnor U5971 (N_5971,N_4045,N_2491);
nor U5972 (N_5972,N_2098,N_2497);
or U5973 (N_5973,N_318,N_2280);
and U5974 (N_5974,N_3556,N_1283);
nand U5975 (N_5975,N_3053,N_1858);
or U5976 (N_5976,N_740,N_3);
or U5977 (N_5977,N_1579,N_1920);
or U5978 (N_5978,N_1038,N_4068);
and U5979 (N_5979,N_3995,N_672);
xnor U5980 (N_5980,N_1151,N_2000);
nand U5981 (N_5981,N_2232,N_510);
xnor U5982 (N_5982,N_1690,N_445);
or U5983 (N_5983,N_4894,N_3369);
or U5984 (N_5984,N_3627,N_4244);
xnor U5985 (N_5985,N_3090,N_4635);
nor U5986 (N_5986,N_4561,N_4103);
nor U5987 (N_5987,N_4690,N_3042);
xor U5988 (N_5988,N_4075,N_4895);
and U5989 (N_5989,N_888,N_3099);
nand U5990 (N_5990,N_163,N_250);
or U5991 (N_5991,N_103,N_2482);
nor U5992 (N_5992,N_4743,N_127);
xnor U5993 (N_5993,N_4435,N_3109);
nor U5994 (N_5994,N_2591,N_4278);
nor U5995 (N_5995,N_3650,N_193);
nand U5996 (N_5996,N_1892,N_3726);
and U5997 (N_5997,N_432,N_3615);
nand U5998 (N_5998,N_217,N_1707);
nor U5999 (N_5999,N_4912,N_4003);
nor U6000 (N_6000,N_3360,N_1816);
nor U6001 (N_6001,N_667,N_4020);
nand U6002 (N_6002,N_2134,N_1164);
nor U6003 (N_6003,N_3942,N_3025);
nand U6004 (N_6004,N_3504,N_2300);
or U6005 (N_6005,N_1704,N_3872);
nor U6006 (N_6006,N_1637,N_3045);
xor U6007 (N_6007,N_4849,N_1818);
nand U6008 (N_6008,N_16,N_1693);
xnor U6009 (N_6009,N_2421,N_4528);
and U6010 (N_6010,N_743,N_613);
nor U6011 (N_6011,N_1553,N_2993);
and U6012 (N_6012,N_443,N_3910);
nand U6013 (N_6013,N_4534,N_3904);
nor U6014 (N_6014,N_4189,N_4995);
xnor U6015 (N_6015,N_4488,N_1515);
and U6016 (N_6016,N_1376,N_3982);
xor U6017 (N_6017,N_2692,N_811);
and U6018 (N_6018,N_3708,N_1919);
and U6019 (N_6019,N_3937,N_1439);
and U6020 (N_6020,N_138,N_2741);
nor U6021 (N_6021,N_4958,N_3459);
or U6022 (N_6022,N_3891,N_1722);
and U6023 (N_6023,N_294,N_146);
nor U6024 (N_6024,N_4907,N_3773);
nor U6025 (N_6025,N_4537,N_298);
or U6026 (N_6026,N_1299,N_1790);
nor U6027 (N_6027,N_4994,N_4085);
and U6028 (N_6028,N_2596,N_4418);
and U6029 (N_6029,N_2879,N_327);
xor U6030 (N_6030,N_4450,N_4641);
and U6031 (N_6031,N_725,N_1670);
xnor U6032 (N_6032,N_2537,N_4084);
and U6033 (N_6033,N_4991,N_2518);
or U6034 (N_6034,N_1749,N_3488);
nand U6035 (N_6035,N_2327,N_2594);
or U6036 (N_6036,N_2852,N_3822);
or U6037 (N_6037,N_3660,N_2662);
or U6038 (N_6038,N_1735,N_8);
or U6039 (N_6039,N_1330,N_3212);
xor U6040 (N_6040,N_4802,N_1710);
nor U6041 (N_6041,N_2044,N_1561);
or U6042 (N_6042,N_2885,N_3619);
or U6043 (N_6043,N_3497,N_4735);
or U6044 (N_6044,N_1256,N_167);
xnor U6045 (N_6045,N_2766,N_728);
nand U6046 (N_6046,N_3023,N_2736);
nand U6047 (N_6047,N_887,N_3148);
nor U6048 (N_6048,N_3864,N_4520);
nand U6049 (N_6049,N_3312,N_1906);
or U6050 (N_6050,N_293,N_4506);
xnor U6051 (N_6051,N_3450,N_1187);
nand U6052 (N_6052,N_2156,N_2059);
nor U6053 (N_6053,N_1539,N_2415);
nand U6054 (N_6054,N_2089,N_1686);
nor U6055 (N_6055,N_2432,N_3235);
nor U6056 (N_6056,N_4622,N_2196);
xor U6057 (N_6057,N_3572,N_28);
nand U6058 (N_6058,N_4264,N_3326);
nand U6059 (N_6059,N_4168,N_24);
or U6060 (N_6060,N_3588,N_3763);
or U6061 (N_6061,N_3638,N_82);
nor U6062 (N_6062,N_524,N_2917);
and U6063 (N_6063,N_3898,N_633);
and U6064 (N_6064,N_2073,N_2830);
and U6065 (N_6065,N_4667,N_4705);
nor U6066 (N_6066,N_3336,N_6);
or U6067 (N_6067,N_3190,N_767);
or U6068 (N_6068,N_1960,N_76);
xnor U6069 (N_6069,N_567,N_2723);
and U6070 (N_6070,N_3949,N_4331);
nand U6071 (N_6071,N_4675,N_1772);
or U6072 (N_6072,N_3308,N_1294);
and U6073 (N_6073,N_3233,N_984);
xor U6074 (N_6074,N_2780,N_1767);
nor U6075 (N_6075,N_3255,N_3867);
nor U6076 (N_6076,N_4116,N_3242);
nor U6077 (N_6077,N_3433,N_1253);
xnor U6078 (N_6078,N_2991,N_223);
nand U6079 (N_6079,N_3104,N_3217);
nand U6080 (N_6080,N_3890,N_2394);
xor U6081 (N_6081,N_3645,N_519);
nand U6082 (N_6082,N_1925,N_1013);
nand U6083 (N_6083,N_4865,N_1128);
and U6084 (N_6084,N_2546,N_1416);
nor U6085 (N_6085,N_1248,N_2490);
and U6086 (N_6086,N_4033,N_1098);
xnor U6087 (N_6087,N_1481,N_4100);
nor U6088 (N_6088,N_4312,N_142);
and U6089 (N_6089,N_1605,N_2420);
nand U6090 (N_6090,N_3711,N_1095);
or U6091 (N_6091,N_2385,N_3888);
nand U6092 (N_6092,N_1988,N_3401);
or U6093 (N_6093,N_2040,N_2384);
and U6094 (N_6094,N_1773,N_2326);
nor U6095 (N_6095,N_844,N_2784);
and U6096 (N_6096,N_4258,N_892);
or U6097 (N_6097,N_2313,N_1657);
or U6098 (N_6098,N_2298,N_3327);
nand U6099 (N_6099,N_143,N_666);
nor U6100 (N_6100,N_4133,N_3924);
or U6101 (N_6101,N_2072,N_3523);
or U6102 (N_6102,N_2775,N_1478);
xor U6103 (N_6103,N_1432,N_4186);
or U6104 (N_6104,N_4395,N_641);
xnor U6105 (N_6105,N_1386,N_251);
or U6106 (N_6106,N_2082,N_2587);
nor U6107 (N_6107,N_3862,N_4238);
or U6108 (N_6108,N_393,N_3101);
nand U6109 (N_6109,N_2201,N_704);
xor U6110 (N_6110,N_3382,N_4229);
nand U6111 (N_6111,N_663,N_2722);
nand U6112 (N_6112,N_331,N_3629);
xnor U6113 (N_6113,N_3413,N_4118);
xnor U6114 (N_6114,N_2895,N_4646);
nand U6115 (N_6115,N_3129,N_2190);
or U6116 (N_6116,N_4558,N_1276);
xnor U6117 (N_6117,N_4285,N_3128);
or U6118 (N_6118,N_620,N_2520);
xnor U6119 (N_6119,N_804,N_382);
nor U6120 (N_6120,N_50,N_2507);
and U6121 (N_6121,N_3779,N_2727);
nor U6122 (N_6122,N_2994,N_1571);
nor U6123 (N_6123,N_1118,N_1282);
nand U6124 (N_6124,N_1989,N_2649);
xnor U6125 (N_6125,N_2189,N_852);
or U6126 (N_6126,N_3426,N_540);
and U6127 (N_6127,N_891,N_2693);
and U6128 (N_6128,N_4644,N_120);
and U6129 (N_6129,N_799,N_4655);
and U6130 (N_6130,N_1566,N_4637);
or U6131 (N_6131,N_1922,N_3778);
nor U6132 (N_6132,N_4971,N_3002);
xnor U6133 (N_6133,N_1264,N_3355);
nand U6134 (N_6134,N_4614,N_1565);
and U6135 (N_6135,N_2198,N_3539);
nor U6136 (N_6136,N_454,N_3290);
xnor U6137 (N_6137,N_2139,N_1897);
nor U6138 (N_6138,N_4571,N_2353);
and U6139 (N_6139,N_3272,N_2595);
nor U6140 (N_6140,N_2095,N_1625);
or U6141 (N_6141,N_1072,N_1794);
and U6142 (N_6142,N_3679,N_3238);
nand U6143 (N_6143,N_3989,N_4233);
or U6144 (N_6144,N_3793,N_360);
nor U6145 (N_6145,N_4475,N_3111);
or U6146 (N_6146,N_2916,N_1221);
xor U6147 (N_6147,N_619,N_123);
nor U6148 (N_6148,N_4419,N_498);
and U6149 (N_6149,N_1564,N_3106);
xnor U6150 (N_6150,N_3870,N_3455);
xor U6151 (N_6151,N_1870,N_4383);
or U6152 (N_6152,N_3589,N_4739);
nor U6153 (N_6153,N_188,N_3704);
and U6154 (N_6154,N_834,N_1130);
nor U6155 (N_6155,N_1470,N_3575);
xnor U6156 (N_6156,N_1813,N_2160);
and U6157 (N_6157,N_1939,N_878);
xor U6158 (N_6158,N_4943,N_3113);
nor U6159 (N_6159,N_1885,N_1005);
or U6160 (N_6160,N_1097,N_4815);
nand U6161 (N_6161,N_882,N_2057);
or U6162 (N_6162,N_373,N_2048);
and U6163 (N_6163,N_771,N_3408);
and U6164 (N_6164,N_1592,N_1857);
nand U6165 (N_6165,N_1871,N_1307);
nor U6166 (N_6166,N_1741,N_1581);
nor U6167 (N_6167,N_3625,N_3869);
or U6168 (N_6168,N_2956,N_1838);
xor U6169 (N_6169,N_4726,N_1108);
or U6170 (N_6170,N_4110,N_1443);
and U6171 (N_6171,N_3635,N_13);
nor U6172 (N_6172,N_1142,N_2470);
xnor U6173 (N_6173,N_4421,N_3967);
and U6174 (N_6174,N_845,N_1414);
nor U6175 (N_6175,N_2569,N_2495);
xor U6176 (N_6176,N_3374,N_581);
or U6177 (N_6177,N_1375,N_580);
nand U6178 (N_6178,N_2431,N_573);
and U6179 (N_6179,N_1000,N_3851);
or U6180 (N_6180,N_2685,N_2589);
and U6181 (N_6181,N_3440,N_4889);
and U6182 (N_6182,N_1928,N_3770);
xor U6183 (N_6183,N_4403,N_2933);
and U6184 (N_6184,N_787,N_3317);
and U6185 (N_6185,N_4508,N_4821);
xor U6186 (N_6186,N_2502,N_4017);
xnor U6187 (N_6187,N_3927,N_3313);
and U6188 (N_6188,N_4585,N_4578);
and U6189 (N_6189,N_4769,N_1809);
or U6190 (N_6190,N_4357,N_2688);
nand U6191 (N_6191,N_3546,N_724);
nor U6192 (N_6192,N_828,N_2002);
and U6193 (N_6193,N_2034,N_1883);
and U6194 (N_6194,N_3695,N_3745);
nor U6195 (N_6195,N_3346,N_195);
xor U6196 (N_6196,N_3658,N_2659);
nor U6197 (N_6197,N_2508,N_3969);
nor U6198 (N_6198,N_2609,N_4205);
nand U6199 (N_6199,N_2838,N_3406);
xor U6200 (N_6200,N_3118,N_2342);
or U6201 (N_6201,N_1437,N_4937);
and U6202 (N_6202,N_2731,N_287);
nor U6203 (N_6203,N_2403,N_4117);
or U6204 (N_6204,N_1196,N_1750);
nand U6205 (N_6205,N_4926,N_550);
or U6206 (N_6206,N_3976,N_1842);
nand U6207 (N_6207,N_2276,N_4138);
and U6208 (N_6208,N_2291,N_3420);
nand U6209 (N_6209,N_995,N_231);
xnor U6210 (N_6210,N_4774,N_669);
and U6211 (N_6211,N_3149,N_2642);
nand U6212 (N_6212,N_981,N_1015);
or U6213 (N_6213,N_665,N_1390);
nor U6214 (N_6214,N_4257,N_4274);
nand U6215 (N_6215,N_757,N_1769);
xor U6216 (N_6216,N_3145,N_3597);
xnor U6217 (N_6217,N_4176,N_3361);
nand U6218 (N_6218,N_1040,N_2909);
nand U6219 (N_6219,N_2212,N_3492);
nand U6220 (N_6220,N_239,N_824);
and U6221 (N_6221,N_3718,N_475);
xor U6222 (N_6222,N_2952,N_137);
or U6223 (N_6223,N_489,N_224);
and U6224 (N_6224,N_2150,N_1785);
nor U6225 (N_6225,N_2730,N_3644);
or U6226 (N_6226,N_356,N_1510);
xnor U6227 (N_6227,N_4858,N_1234);
nor U6228 (N_6228,N_4416,N_1448);
nor U6229 (N_6229,N_241,N_3340);
xor U6230 (N_6230,N_930,N_2175);
nand U6231 (N_6231,N_3192,N_912);
or U6232 (N_6232,N_3573,N_2998);
nor U6233 (N_6233,N_1181,N_4239);
and U6234 (N_6234,N_158,N_690);
and U6235 (N_6235,N_2486,N_3940);
and U6236 (N_6236,N_651,N_1345);
xor U6237 (N_6237,N_736,N_530);
nor U6238 (N_6238,N_2435,N_4773);
or U6239 (N_6239,N_70,N_4425);
and U6240 (N_6240,N_4018,N_3999);
and U6241 (N_6241,N_77,N_4788);
nand U6242 (N_6242,N_4920,N_1634);
nand U6243 (N_6243,N_3026,N_716);
nand U6244 (N_6244,N_4877,N_621);
nand U6245 (N_6245,N_4354,N_3089);
nand U6246 (N_6246,N_3067,N_3669);
xor U6247 (N_6247,N_4437,N_3820);
and U6248 (N_6248,N_1864,N_4507);
and U6249 (N_6249,N_4593,N_2868);
xor U6250 (N_6250,N_3985,N_4039);
and U6251 (N_6251,N_3925,N_4985);
and U6252 (N_6252,N_4036,N_4455);
and U6253 (N_6253,N_277,N_2845);
nor U6254 (N_6254,N_4171,N_3601);
xor U6255 (N_6255,N_65,N_4462);
nand U6256 (N_6256,N_3761,N_671);
and U6257 (N_6257,N_2503,N_1908);
xor U6258 (N_6258,N_749,N_1348);
and U6259 (N_6259,N_4453,N_3261);
xor U6260 (N_6260,N_702,N_4180);
xnor U6261 (N_6261,N_4562,N_1909);
nand U6262 (N_6262,N_2433,N_3799);
nor U6263 (N_6263,N_604,N_3180);
xnor U6264 (N_6264,N_2335,N_104);
xor U6265 (N_6265,N_1996,N_1598);
nor U6266 (N_6266,N_3681,N_662);
nor U6267 (N_6267,N_527,N_2905);
nor U6268 (N_6268,N_4624,N_4446);
nor U6269 (N_6269,N_2194,N_2083);
and U6270 (N_6270,N_2689,N_3075);
and U6271 (N_6271,N_2800,N_3640);
nand U6272 (N_6272,N_495,N_4464);
nor U6273 (N_6273,N_627,N_2528);
and U6274 (N_6274,N_4944,N_554);
and U6275 (N_6275,N_3651,N_2231);
nor U6276 (N_6276,N_1972,N_1224);
and U6277 (N_6277,N_2301,N_2512);
nor U6278 (N_6278,N_2380,N_822);
and U6279 (N_6279,N_3755,N_4184);
and U6280 (N_6280,N_2794,N_1421);
or U6281 (N_6281,N_1339,N_2904);
nor U6282 (N_6282,N_221,N_4879);
nor U6283 (N_6283,N_4764,N_3263);
nor U6284 (N_6284,N_1341,N_1962);
nor U6285 (N_6285,N_2462,N_1770);
xor U6286 (N_6286,N_966,N_4514);
or U6287 (N_6287,N_1927,N_1520);
nor U6288 (N_6288,N_2253,N_3367);
xor U6289 (N_6289,N_2115,N_1779);
xor U6290 (N_6290,N_4908,N_1235);
xor U6291 (N_6291,N_2637,N_1696);
nor U6292 (N_6292,N_3852,N_2244);
xnor U6293 (N_6293,N_2208,N_1301);
nor U6294 (N_6294,N_2585,N_3259);
nand U6295 (N_6295,N_4618,N_614);
and U6296 (N_6296,N_3757,N_4710);
nor U6297 (N_6297,N_2449,N_113);
xor U6298 (N_6298,N_211,N_3609);
or U6299 (N_6299,N_4438,N_3945);
or U6300 (N_6300,N_721,N_3043);
and U6301 (N_6301,N_434,N_2703);
nand U6302 (N_6302,N_461,N_45);
and U6303 (N_6303,N_3784,N_546);
nor U6304 (N_6304,N_1640,N_898);
nor U6305 (N_6305,N_2333,N_377);
or U6306 (N_6306,N_1337,N_3416);
nand U6307 (N_6307,N_3668,N_2358);
or U6308 (N_6308,N_4790,N_1854);
nand U6309 (N_6309,N_2965,N_1259);
nor U6310 (N_6310,N_1958,N_395);
nand U6311 (N_6311,N_4785,N_4859);
nor U6312 (N_6312,N_2961,N_1113);
and U6313 (N_6313,N_3427,N_3508);
nor U6314 (N_6314,N_2131,N_4326);
nor U6315 (N_6315,N_578,N_969);
or U6316 (N_6316,N_2319,N_2890);
or U6317 (N_6317,N_34,N_2921);
xor U6318 (N_6318,N_973,N_157);
nand U6319 (N_6319,N_3735,N_2953);
and U6320 (N_6320,N_4470,N_3392);
and U6321 (N_6321,N_3714,N_4906);
and U6322 (N_6322,N_3648,N_1523);
nand U6323 (N_6323,N_4261,N_712);
nand U6324 (N_6324,N_4024,N_1604);
nor U6325 (N_6325,N_3465,N_2162);
xnor U6326 (N_6326,N_3321,N_762);
xor U6327 (N_6327,N_1964,N_1318);
and U6328 (N_6328,N_4369,N_176);
or U6329 (N_6329,N_3215,N_3918);
or U6330 (N_6330,N_1865,N_3154);
nand U6331 (N_6331,N_4202,N_4838);
or U6332 (N_6332,N_41,N_3080);
and U6333 (N_6333,N_4549,N_1787);
nor U6334 (N_6334,N_1412,N_1175);
nor U6335 (N_6335,N_3686,N_3506);
and U6336 (N_6336,N_2867,N_368);
xor U6337 (N_6337,N_1077,N_2821);
nor U6338 (N_6338,N_983,N_2856);
nand U6339 (N_6339,N_4720,N_2726);
nand U6340 (N_6340,N_2122,N_1085);
nand U6341 (N_6341,N_583,N_3682);
nor U6342 (N_6342,N_4384,N_140);
nand U6343 (N_6343,N_1721,N_2506);
xnor U6344 (N_6344,N_3011,N_2816);
nand U6345 (N_6345,N_3516,N_1056);
nor U6346 (N_6346,N_4899,N_3294);
nor U6347 (N_6347,N_437,N_2556);
nand U6348 (N_6348,N_2029,N_1263);
nor U6349 (N_6349,N_148,N_3471);
nor U6350 (N_6350,N_4473,N_1661);
nor U6351 (N_6351,N_4299,N_3245);
nor U6352 (N_6352,N_2164,N_2908);
and U6353 (N_6353,N_3206,N_1662);
and U6354 (N_6354,N_3611,N_570);
nor U6355 (N_6355,N_2534,N_4309);
and U6356 (N_6356,N_1495,N_4095);
and U6357 (N_6357,N_111,N_2554);
xnor U6358 (N_6358,N_3802,N_2092);
nand U6359 (N_6359,N_548,N_2461);
nor U6360 (N_6360,N_208,N_1937);
or U6361 (N_6361,N_2357,N_2279);
nor U6362 (N_6362,N_1279,N_161);
nand U6363 (N_6363,N_2592,N_1230);
or U6364 (N_6364,N_3715,N_829);
nor U6365 (N_6365,N_615,N_4924);
nor U6366 (N_6366,N_1763,N_131);
or U6367 (N_6367,N_3036,N_422);
xnor U6368 (N_6368,N_680,N_3541);
and U6369 (N_6369,N_4271,N_3289);
xnor U6370 (N_6370,N_4461,N_3083);
or U6371 (N_6371,N_84,N_2124);
nor U6372 (N_6372,N_2896,N_4553);
nand U6373 (N_6373,N_2509,N_1516);
nand U6374 (N_6374,N_692,N_727);
xnor U6375 (N_6375,N_21,N_4002);
nor U6376 (N_6376,N_2469,N_0);
or U6377 (N_6377,N_3617,N_2744);
nor U6378 (N_6378,N_4012,N_753);
and U6379 (N_6379,N_367,N_4144);
nand U6380 (N_6380,N_1115,N_1841);
and U6381 (N_6381,N_3670,N_739);
and U6382 (N_6382,N_3903,N_3612);
nor U6383 (N_6383,N_513,N_1400);
xnor U6384 (N_6384,N_3768,N_4560);
xor U6385 (N_6385,N_2242,N_1029);
and U6386 (N_6386,N_4866,N_4625);
and U6387 (N_6387,N_4330,N_737);
nor U6388 (N_6388,N_988,N_2620);
xnor U6389 (N_6389,N_4194,N_2875);
and U6390 (N_6390,N_1210,N_4522);
xor U6391 (N_6391,N_968,N_2129);
or U6392 (N_6392,N_4732,N_1911);
nor U6393 (N_6393,N_3189,N_1833);
nor U6394 (N_6394,N_4500,N_92);
xnor U6395 (N_6395,N_2022,N_4174);
xor U6396 (N_6396,N_2625,N_798);
xor U6397 (N_6397,N_2401,N_2426);
nor U6398 (N_6398,N_504,N_197);
nand U6399 (N_6399,N_2843,N_4208);
and U6400 (N_6400,N_2205,N_1141);
nand U6401 (N_6401,N_1667,N_3621);
and U6402 (N_6402,N_3654,N_2414);
nor U6403 (N_6403,N_2494,N_3628);
nor U6404 (N_6404,N_975,N_4098);
xnor U6405 (N_6405,N_4415,N_2762);
nand U6406 (N_6406,N_3073,N_3552);
or U6407 (N_6407,N_1945,N_1517);
xor U6408 (N_6408,N_1180,N_1650);
and U6409 (N_6409,N_3527,N_4305);
nand U6410 (N_6410,N_1002,N_2383);
nor U6411 (N_6411,N_1392,N_1877);
xor U6412 (N_6412,N_4491,N_635);
xnor U6413 (N_6413,N_3576,N_4423);
nor U6414 (N_6414,N_2574,N_2806);
and U6415 (N_6415,N_3363,N_2445);
xnor U6416 (N_6416,N_3162,N_4260);
xnor U6417 (N_6417,N_4230,N_3697);
nand U6418 (N_6418,N_2015,N_1183);
and U6419 (N_6419,N_2406,N_4226);
nor U6420 (N_6420,N_2229,N_2742);
or U6421 (N_6421,N_1014,N_3126);
or U6422 (N_6422,N_1018,N_1278);
xor U6423 (N_6423,N_1026,N_349);
and U6424 (N_6424,N_4803,N_1629);
xor U6425 (N_6425,N_3207,N_4940);
nand U6426 (N_6426,N_2146,N_2250);
nand U6427 (N_6427,N_2516,N_2949);
nor U6428 (N_6428,N_1126,N_4851);
nor U6429 (N_6429,N_4822,N_3040);
xnor U6430 (N_6430,N_1643,N_1227);
nor U6431 (N_6431,N_4904,N_3592);
or U6432 (N_6432,N_751,N_4777);
nor U6433 (N_6433,N_1687,N_1558);
and U6434 (N_6434,N_3931,N_1017);
nand U6435 (N_6435,N_2138,N_4979);
and U6436 (N_6436,N_2365,N_1832);
or U6437 (N_6437,N_2771,N_3257);
or U6438 (N_6438,N_994,N_4729);
nor U6439 (N_6439,N_1985,N_536);
or U6440 (N_6440,N_2148,N_3136);
xnor U6441 (N_6441,N_2522,N_1601);
or U6442 (N_6442,N_2931,N_4768);
nand U6443 (N_6443,N_4540,N_2500);
or U6444 (N_6444,N_2683,N_588);
xor U6445 (N_6445,N_3610,N_4934);
or U6446 (N_6446,N_2653,N_3514);
or U6447 (N_6447,N_4844,N_2761);
or U6448 (N_6448,N_54,N_3475);
and U6449 (N_6449,N_2478,N_3507);
and U6450 (N_6450,N_4056,N_1990);
nand U6451 (N_6451,N_4156,N_1930);
nand U6452 (N_6452,N_2760,N_1075);
xor U6453 (N_6453,N_2102,N_3305);
nor U6454 (N_6454,N_1123,N_708);
or U6455 (N_6455,N_3016,N_4502);
nand U6456 (N_6456,N_1682,N_4661);
xnor U6457 (N_6457,N_48,N_4530);
and U6458 (N_6458,N_1575,N_1043);
xor U6459 (N_6459,N_314,N_2);
and U6460 (N_6460,N_2682,N_2496);
or U6461 (N_6461,N_3739,N_2708);
and U6462 (N_6462,N_4151,N_3069);
or U6463 (N_6463,N_754,N_3855);
or U6464 (N_6464,N_2674,N_4845);
or U6465 (N_6465,N_183,N_2025);
and U6466 (N_6466,N_4724,N_2079);
and U6467 (N_6467,N_4339,N_2058);
and U6468 (N_6468,N_348,N_4216);
or U6469 (N_6469,N_3873,N_220);
nand U6470 (N_6470,N_1121,N_4748);
nor U6471 (N_6471,N_279,N_2278);
nand U6472 (N_6472,N_4634,N_2709);
nand U6473 (N_6473,N_3250,N_1835);
and U6474 (N_6474,N_602,N_2918);
and U6475 (N_6475,N_2880,N_2711);
nand U6476 (N_6476,N_2314,N_1117);
or U6477 (N_6477,N_608,N_4969);
xor U6478 (N_6478,N_1092,N_4513);
or U6479 (N_6479,N_2725,N_3751);
nand U6480 (N_6480,N_2866,N_3968);
nand U6481 (N_6481,N_1127,N_3251);
and U6482 (N_6482,N_89,N_3809);
xnor U6483 (N_6483,N_1895,N_4846);
xor U6484 (N_6484,N_27,N_2747);
xnor U6485 (N_6485,N_3893,N_2350);
xor U6486 (N_6486,N_789,N_3085);
xor U6487 (N_6487,N_3147,N_654);
xnor U6488 (N_6488,N_1652,N_1709);
nor U6489 (N_6489,N_3343,N_3254);
or U6490 (N_6490,N_4241,N_1381);
nor U6491 (N_6491,N_3258,N_750);
nand U6492 (N_6492,N_256,N_637);
or U6493 (N_6493,N_3883,N_2460);
and U6494 (N_6494,N_347,N_2219);
xnor U6495 (N_6495,N_1059,N_1458);
and U6496 (N_6496,N_4538,N_2238);
and U6497 (N_6497,N_3548,N_3210);
xnor U6498 (N_6498,N_1903,N_2256);
nor U6499 (N_6499,N_2252,N_1555);
and U6500 (N_6500,N_3146,N_2561);
xor U6501 (N_6501,N_3335,N_537);
nor U6502 (N_6502,N_2422,N_2987);
nor U6503 (N_6503,N_3753,N_4097);
and U6504 (N_6504,N_2481,N_3709);
xor U6505 (N_6505,N_2808,N_3143);
and U6506 (N_6506,N_1105,N_59);
and U6507 (N_6507,N_4286,N_935);
and U6508 (N_6508,N_4930,N_4459);
and U6509 (N_6509,N_2667,N_4965);
xor U6510 (N_6510,N_929,N_4322);
or U6511 (N_6511,N_410,N_3065);
nand U6512 (N_6512,N_1358,N_836);
nand U6513 (N_6513,N_4843,N_2225);
xor U6514 (N_6514,N_1409,N_3791);
nor U6515 (N_6515,N_487,N_357);
or U6516 (N_6516,N_1406,N_1726);
and U6517 (N_6517,N_439,N_1781);
nand U6518 (N_6518,N_3846,N_957);
nand U6519 (N_6519,N_248,N_3688);
and U6520 (N_6520,N_1712,N_290);
or U6521 (N_6521,N_4292,N_1208);
nor U6522 (N_6522,N_459,N_4699);
and U6523 (N_6523,N_4929,N_4700);
nand U6524 (N_6524,N_3431,N_1853);
nor U6525 (N_6525,N_2425,N_2684);
xnor U6526 (N_6526,N_643,N_563);
xor U6527 (N_6527,N_153,N_3807);
xnor U6528 (N_6528,N_4993,N_2104);
xor U6529 (N_6529,N_3435,N_2028);
nand U6530 (N_6530,N_2783,N_4781);
nand U6531 (N_6531,N_4181,N_1595);
and U6532 (N_6532,N_2573,N_4303);
or U6533 (N_6533,N_3756,N_4388);
nor U6534 (N_6534,N_1146,N_1311);
xnor U6535 (N_6535,N_212,N_134);
nand U6536 (N_6536,N_684,N_2755);
nor U6537 (N_6537,N_1385,N_2459);
and U6538 (N_6538,N_2006,N_4307);
or U6539 (N_6539,N_1692,N_405);
xnor U6540 (N_6540,N_2975,N_4397);
and U6541 (N_6541,N_943,N_2336);
xor U6542 (N_6542,N_758,N_3443);
nor U6543 (N_6543,N_2769,N_880);
nor U6544 (N_6544,N_246,N_1974);
xnor U6545 (N_6545,N_2563,N_1313);
or U6546 (N_6546,N_4318,N_4000);
or U6547 (N_6547,N_2010,N_3801);
or U6548 (N_6548,N_3347,N_3276);
nor U6549 (N_6549,N_1083,N_1352);
nand U6550 (N_6550,N_2764,N_1185);
or U6551 (N_6551,N_3218,N_1321);
and U6552 (N_6552,N_3429,N_2094);
nor U6553 (N_6553,N_3630,N_603);
nor U6554 (N_6554,N_2081,N_2423);
or U6555 (N_6555,N_3486,N_1508);
or U6556 (N_6556,N_2582,N_3095);
nor U6557 (N_6557,N_1364,N_953);
or U6558 (N_6558,N_2927,N_2940);
nand U6559 (N_6559,N_4248,N_3643);
and U6560 (N_6560,N_2560,N_960);
nand U6561 (N_6561,N_4076,N_1633);
nand U6562 (N_6562,N_2265,N_2888);
or U6563 (N_6563,N_1114,N_446);
or U6564 (N_6564,N_1702,N_4172);
or U6565 (N_6565,N_3469,N_374);
or U6566 (N_6566,N_3282,N_1525);
or U6567 (N_6567,N_30,N_3468);
or U6568 (N_6568,N_4032,N_2883);
and U6569 (N_6569,N_1425,N_79);
xnor U6570 (N_6570,N_1393,N_1455);
nor U6571 (N_6571,N_1863,N_3696);
xor U6572 (N_6572,N_4915,N_3076);
and U6573 (N_6573,N_4660,N_3608);
or U6574 (N_6574,N_2551,N_85);
xor U6575 (N_6575,N_2045,N_1612);
and U6576 (N_6576,N_4169,N_2019);
xnor U6577 (N_6577,N_2101,N_4770);
xnor U6578 (N_6578,N_4463,N_1451);
nor U6579 (N_6579,N_2086,N_2168);
nor U6580 (N_6580,N_3153,N_1817);
and U6581 (N_6581,N_2846,N_2153);
or U6582 (N_6582,N_2293,N_29);
nor U6583 (N_6583,N_2295,N_3722);
or U6584 (N_6584,N_1257,N_2955);
nor U6585 (N_6585,N_4346,N_4358);
and U6586 (N_6586,N_877,N_3405);
nor U6587 (N_6587,N_4121,N_3221);
or U6588 (N_6588,N_3678,N_2570);
nor U6589 (N_6589,N_3044,N_1192);
nand U6590 (N_6590,N_2962,N_2152);
nor U6591 (N_6591,N_4209,N_1648);
or U6592 (N_6592,N_4277,N_1399);
nor U6593 (N_6593,N_1436,N_1331);
and U6594 (N_6594,N_1452,N_3614);
xor U6595 (N_6595,N_4778,N_2828);
or U6596 (N_6596,N_2915,N_3962);
or U6597 (N_6597,N_4341,N_4616);
xnor U6598 (N_6598,N_4811,N_2078);
nor U6599 (N_6599,N_2145,N_3540);
or U6600 (N_6600,N_3390,N_3979);
xor U6601 (N_6601,N_3758,N_4412);
xor U6602 (N_6602,N_4697,N_695);
xor U6603 (N_6603,N_2532,N_3006);
xor U6604 (N_6604,N_1054,N_4835);
xnor U6605 (N_6605,N_25,N_2363);
xor U6606 (N_6606,N_4653,N_1602);
xor U6607 (N_6607,N_3158,N_2268);
nor U6608 (N_6608,N_3876,N_4315);
or U6609 (N_6609,N_301,N_1708);
nor U6610 (N_6610,N_3544,N_4529);
and U6611 (N_6611,N_3461,N_289);
and U6612 (N_6612,N_4584,N_2643);
and U6613 (N_6613,N_1201,N_3430);
nor U6614 (N_6614,N_4923,N_971);
nor U6615 (N_6615,N_4466,N_2367);
nand U6616 (N_6616,N_3319,N_3088);
and U6617 (N_6617,N_3015,N_626);
and U6618 (N_6618,N_1160,N_1155);
nand U6619 (N_6619,N_4792,N_2663);
xnor U6620 (N_6620,N_2228,N_3170);
nand U6621 (N_6621,N_4757,N_2884);
or U6622 (N_6622,N_3300,N_1255);
xor U6623 (N_6623,N_3208,N_108);
nand U6624 (N_6624,N_3155,N_1669);
xor U6625 (N_6625,N_2049,N_1370);
xnor U6626 (N_6626,N_2032,N_403);
or U6627 (N_6627,N_321,N_3897);
nand U6628 (N_6628,N_1699,N_1144);
nor U6629 (N_6629,N_1965,N_978);
and U6630 (N_6630,N_555,N_3774);
xor U6631 (N_6631,N_766,N_1823);
or U6632 (N_6632,N_3108,N_790);
or U6633 (N_6633,N_1033,N_1158);
and U6634 (N_6634,N_492,N_3836);
nand U6635 (N_6635,N_1079,N_3056);
xnor U6636 (N_6636,N_2438,N_1492);
and U6637 (N_6637,N_3184,N_673);
xnor U6638 (N_6638,N_1023,N_2706);
nand U6639 (N_6639,N_2603,N_278);
nand U6640 (N_6640,N_2259,N_2717);
xnor U6641 (N_6641,N_456,N_1340);
xnor U6642 (N_6642,N_3916,N_1609);
and U6643 (N_6643,N_1383,N_4043);
nor U6644 (N_6644,N_1534,N_4126);
and U6645 (N_6645,N_2050,N_559);
or U6646 (N_6646,N_273,N_2479);
or U6647 (N_6647,N_4516,N_1366);
and U6648 (N_6648,N_235,N_4762);
nor U6649 (N_6649,N_359,N_3354);
or U6650 (N_6650,N_4526,N_859);
nor U6651 (N_6651,N_774,N_295);
nor U6652 (N_6652,N_2308,N_3787);
and U6653 (N_6653,N_310,N_3515);
nand U6654 (N_6654,N_3930,N_941);
or U6655 (N_6655,N_2501,N_64);
nand U6656 (N_6656,N_2634,N_3915);
xnor U6657 (N_6657,N_93,N_3996);
or U6658 (N_6658,N_4647,N_2234);
and U6659 (N_6659,N_4114,N_585);
nor U6660 (N_6660,N_1036,N_1286);
xnor U6661 (N_6661,N_1284,N_3348);
and U6662 (N_6662,N_1978,N_267);
or U6663 (N_6663,N_967,N_2992);
and U6664 (N_6664,N_4478,N_2826);
and U6665 (N_6665,N_539,N_3168);
xnor U6666 (N_6666,N_2668,N_4839);
nor U6667 (N_6667,N_4221,N_1719);
xnor U6668 (N_6668,N_1610,N_406);
and U6669 (N_6669,N_2451,N_4935);
nand U6670 (N_6670,N_4066,N_1874);
and U6671 (N_6671,N_2177,N_2857);
and U6672 (N_6672,N_2033,N_1244);
and U6673 (N_6673,N_3159,N_2498);
nor U6674 (N_6674,N_121,N_2613);
nand U6675 (N_6675,N_2781,N_2041);
xnor U6676 (N_6676,N_1046,N_2130);
nand U6677 (N_6677,N_3328,N_490);
or U6678 (N_6678,N_502,N_3185);
or U6679 (N_6679,N_3409,N_364);
nor U6680 (N_6680,N_3436,N_1544);
xor U6681 (N_6681,N_4231,N_1101);
xnor U6682 (N_6682,N_4856,N_3503);
nor U6683 (N_6683,N_3120,N_4795);
nand U6684 (N_6684,N_2062,N_3725);
or U6685 (N_6685,N_4736,N_3626);
xnor U6686 (N_6686,N_299,N_4609);
and U6687 (N_6687,N_1829,N_901);
xnor U6688 (N_6688,N_3142,N_1353);
and U6689 (N_6689,N_2193,N_2369);
nand U6690 (N_6690,N_2402,N_4053);
nand U6691 (N_6691,N_691,N_1338);
nand U6692 (N_6692,N_777,N_3933);
nor U6693 (N_6693,N_4007,N_1246);
or U6694 (N_6694,N_2932,N_1700);
nor U6695 (N_6695,N_2343,N_3944);
or U6696 (N_6696,N_3583,N_1588);
and U6697 (N_6697,N_3712,N_4497);
xnor U6698 (N_6698,N_2542,N_285);
or U6699 (N_6699,N_4786,N_350);
nand U6700 (N_6700,N_1867,N_1415);
and U6701 (N_6701,N_22,N_4325);
or U6702 (N_6702,N_2323,N_1502);
nor U6703 (N_6703,N_4426,N_172);
xnor U6704 (N_6704,N_1178,N_1200);
xnor U6705 (N_6705,N_2876,N_2359);
nand U6706 (N_6706,N_2705,N_4333);
nor U6707 (N_6707,N_601,N_4367);
nand U6708 (N_6708,N_1217,N_1851);
or U6709 (N_6709,N_3533,N_4072);
nor U6710 (N_6710,N_2362,N_15);
and U6711 (N_6711,N_779,N_319);
xnor U6712 (N_6712,N_2389,N_181);
and U6713 (N_6713,N_3997,N_1666);
xnor U6714 (N_6714,N_1357,N_3123);
xor U6715 (N_6715,N_3692,N_869);
xnor U6716 (N_6716,N_1243,N_2216);
or U6717 (N_6717,N_4149,N_1808);
and U6718 (N_6718,N_2772,N_2434);
or U6719 (N_6719,N_4219,N_2005);
nand U6720 (N_6720,N_1837,N_3816);
nor U6721 (N_6721,N_769,N_3905);
or U6722 (N_6722,N_1135,N_1932);
or U6723 (N_6723,N_168,N_3840);
xnor U6724 (N_6724,N_1560,N_2169);
nor U6725 (N_6725,N_763,N_1454);
or U6726 (N_6726,N_1587,N_3357);
and U6727 (N_6727,N_1554,N_640);
and U6728 (N_6728,N_109,N_4628);
xor U6729 (N_6729,N_1125,N_870);
nor U6730 (N_6730,N_4328,N_3500);
nand U6731 (N_6731,N_3663,N_3939);
xnor U6732 (N_6732,N_1060,N_4368);
or U6733 (N_6733,N_4606,N_2283);
xor U6734 (N_6734,N_3639,N_1747);
and U6735 (N_6735,N_83,N_1132);
xor U6736 (N_6736,N_1446,N_1198);
and U6737 (N_6737,N_1342,N_2439);
nor U6738 (N_6738,N_1624,N_4627);
xnor U6739 (N_6739,N_2030,N_2035);
xnor U6740 (N_6740,N_2966,N_1850);
or U6741 (N_6741,N_3948,N_4950);
or U6742 (N_6742,N_4016,N_2677);
nor U6743 (N_6743,N_4422,N_1580);
xor U6744 (N_6744,N_470,N_2792);
nand U6745 (N_6745,N_3140,N_20);
or U6746 (N_6746,N_3262,N_2368);
nand U6747 (N_6747,N_4663,N_1757);
nand U6748 (N_6748,N_3167,N_4196);
and U6749 (N_6749,N_1220,N_4766);
nand U6750 (N_6750,N_2114,N_3182);
or U6751 (N_6751,N_2457,N_11);
nor U6752 (N_6752,N_4747,N_4253);
or U6753 (N_6753,N_586,N_1188);
and U6754 (N_6754,N_1440,N_3082);
nand U6755 (N_6755,N_1407,N_1204);
or U6756 (N_6756,N_124,N_3021);
xnor U6757 (N_6757,N_194,N_3875);
xnor U6758 (N_6758,N_2754,N_2882);
or U6759 (N_6759,N_1799,N_918);
nor U6760 (N_6760,N_1401,N_228);
or U6761 (N_6761,N_857,N_1550);
and U6762 (N_6762,N_415,N_339);
and U6763 (N_6763,N_3237,N_4191);
xor U6764 (N_6764,N_2263,N_214);
nand U6765 (N_6765,N_1775,N_2170);
or U6766 (N_6766,N_1737,N_808);
and U6767 (N_6767,N_630,N_2088);
xnor U6768 (N_6768,N_3499,N_4888);
nand U6769 (N_6769,N_4349,N_2202);
or U6770 (N_6770,N_2413,N_4608);
and U6771 (N_6771,N_1270,N_2832);
nor U6772 (N_6772,N_3385,N_96);
and U6773 (N_6773,N_1080,N_4977);
xnor U6774 (N_6774,N_3062,N_3744);
and U6775 (N_6775,N_939,N_2604);
or U6776 (N_6776,N_38,N_2347);
and U6777 (N_6777,N_3225,N_2842);
xor U6778 (N_6778,N_2984,N_2981);
nor U6779 (N_6779,N_156,N_596);
xor U6780 (N_6780,N_1417,N_3151);
nand U6781 (N_6781,N_110,N_3762);
or U6782 (N_6782,N_4715,N_2055);
or U6783 (N_6783,N_4809,N_2858);
xor U6784 (N_6784,N_3364,N_1463);
xnor U6785 (N_6785,N_2430,N_842);
and U6786 (N_6786,N_3293,N_800);
xor U6787 (N_6787,N_3007,N_634);
or U6788 (N_6788,N_275,N_4596);
nand U6789 (N_6789,N_4806,N_3978);
or U6790 (N_6790,N_2344,N_3585);
xnor U6791 (N_6791,N_3826,N_255);
and U6792 (N_6792,N_632,N_3373);
or U6793 (N_6793,N_2700,N_696);
nand U6794 (N_6794,N_201,N_2077);
nand U6795 (N_6795,N_268,N_1404);
nor U6796 (N_6796,N_2811,N_1672);
xor U6797 (N_6797,N_4477,N_4539);
nand U6798 (N_6798,N_1961,N_514);
nand U6799 (N_6799,N_4389,N_2943);
or U6800 (N_6800,N_1493,N_926);
or U6801 (N_6801,N_4193,N_4648);
nor U6802 (N_6802,N_4344,N_3452);
xnor U6803 (N_6803,N_4941,N_4490);
and U6804 (N_6804,N_7,N_471);
nand U6805 (N_6805,N_2871,N_703);
or U6806 (N_6806,N_4481,N_457);
nand U6807 (N_6807,N_2658,N_1316);
nor U6808 (N_6808,N_3105,N_4954);
nor U6809 (N_6809,N_4719,N_3955);
or U6810 (N_6810,N_961,N_252);
or U6811 (N_6811,N_387,N_3304);
nand U6812 (N_6812,N_18,N_3278);
xnor U6813 (N_6813,N_423,N_4082);
or U6814 (N_6814,N_4948,N_2818);
or U6815 (N_6815,N_2997,N_4363);
nand U6816 (N_6816,N_3581,N_316);
nand U6817 (N_6817,N_388,N_2061);
nor U6818 (N_6818,N_4810,N_3423);
or U6819 (N_6819,N_1485,N_4152);
and U6820 (N_6820,N_3531,N_3719);
nor U6821 (N_6821,N_3178,N_3653);
or U6822 (N_6822,N_4936,N_3859);
nor U6823 (N_6823,N_3352,N_1955);
nand U6824 (N_6824,N_427,N_3853);
nand U6825 (N_6825,N_2919,N_622);
or U6826 (N_6826,N_4454,N_4474);
nor U6827 (N_6827,N_3689,N_2373);
or U6828 (N_6828,N_1445,N_2237);
xor U6829 (N_6829,N_2176,N_2339);
or U6830 (N_6830,N_4861,N_4401);
nand U6831 (N_6831,N_2815,N_533);
and U6832 (N_6832,N_3740,N_815);
nor U6833 (N_6833,N_3084,N_4928);
or U6834 (N_6834,N_1820,N_452);
nor U6835 (N_6835,N_3325,N_1468);
xor U6836 (N_6836,N_4853,N_1901);
nand U6837 (N_6837,N_352,N_3008);
nor U6838 (N_6838,N_4077,N_149);
and U6839 (N_6839,N_3970,N_210);
or U6840 (N_6840,N_4055,N_4730);
nor U6841 (N_6841,N_1891,N_307);
nor U6842 (N_6842,N_3046,N_1915);
xnor U6843 (N_6843,N_4987,N_1826);
or U6844 (N_6844,N_921,N_4310);
nor U6845 (N_6845,N_1728,N_1021);
or U6846 (N_6846,N_1011,N_3138);
and U6847 (N_6847,N_2103,N_4348);
nand U6848 (N_6848,N_612,N_801);
and U6849 (N_6849,N_1068,N_3152);
xor U6850 (N_6850,N_1593,N_430);
or U6851 (N_6851,N_1148,N_1147);
nand U6852 (N_6852,N_999,N_1214);
and U6853 (N_6853,N_1361,N_3197);
xnor U6854 (N_6854,N_2031,N_1438);
xor U6855 (N_6855,N_2618,N_386);
and U6856 (N_6856,N_2948,N_3000);
nand U6857 (N_6857,N_770,N_2463);
or U6858 (N_6858,N_4382,N_33);
or U6859 (N_6859,N_425,N_402);
and U6860 (N_6860,N_2128,N_3549);
nor U6861 (N_6861,N_9,N_4215);
nor U6862 (N_6862,N_3341,N_2043);
nor U6863 (N_6863,N_4443,N_376);
xnor U6864 (N_6864,N_3116,N_3993);
nor U6865 (N_6865,N_4875,N_4575);
and U6866 (N_6866,N_3936,N_1069);
nor U6867 (N_6867,N_3698,N_1512);
or U6868 (N_6868,N_849,N_1420);
nand U6869 (N_6869,N_1461,N_3027);
nor U6870 (N_6870,N_3512,N_100);
nand U6871 (N_6871,N_4933,N_2543);
nor U6872 (N_6872,N_3114,N_3951);
or U6873 (N_6873,N_4413,N_4535);
xor U6874 (N_6874,N_3164,N_1216);
nor U6875 (N_6875,N_2386,N_3240);
xnor U6876 (N_6876,N_3403,N_2739);
xnor U6877 (N_6877,N_2763,N_4301);
and U6878 (N_6878,N_2898,N_2691);
and U6879 (N_6879,N_4505,N_556);
and U6880 (N_6880,N_3060,N_3966);
or U6881 (N_6881,N_2790,N_3055);
or U6882 (N_6882,N_1614,N_951);
or U6883 (N_6883,N_2183,N_2629);
and U6884 (N_6884,N_1890,N_3213);
nor U6885 (N_6885,N_1139,N_4524);
and U6886 (N_6886,N_4918,N_1584);
or U6887 (N_6887,N_3366,N_3273);
and U6888 (N_6888,N_4551,N_3543);
and U6889 (N_6889,N_2950,N_4559);
or U6890 (N_6890,N_2264,N_3587);
nor U6891 (N_6891,N_1973,N_4010);
nor U6892 (N_6892,N_3521,N_4306);
xnor U6893 (N_6893,N_4718,N_3256);
xnor U6894 (N_6894,N_2778,N_3584);
or U6895 (N_6895,N_1636,N_4447);
or U6896 (N_6896,N_2941,N_689);
nand U6897 (N_6897,N_2312,N_159);
and U6898 (N_6898,N_4573,N_4911);
and U6899 (N_6899,N_2304,N_2902);
or U6900 (N_6900,N_4503,N_2467);
or U6901 (N_6901,N_2740,N_1169);
and U6902 (N_6902,N_970,N_1979);
xnor U6903 (N_6903,N_977,N_196);
and U6904 (N_6904,N_1111,N_1110);
and U6905 (N_6905,N_2274,N_4642);
nand U6906 (N_6906,N_821,N_1509);
and U6907 (N_6907,N_2184,N_2388);
and U6908 (N_6908,N_4581,N_3432);
nor U6909 (N_6909,N_4613,N_4761);
nor U6910 (N_6910,N_264,N_74);
xor U6911 (N_6911,N_2835,N_1129);
nor U6912 (N_6912,N_1798,N_442);
or U6913 (N_6913,N_1297,N_2524);
or U6914 (N_6914,N_375,N_2733);
and U6915 (N_6915,N_1761,N_917);
nor U6916 (N_6916,N_3567,N_200);
nand U6917 (N_6917,N_2317,N_3179);
nand U6918 (N_6918,N_4591,N_4040);
nand U6919 (N_6919,N_4749,N_1992);
nor U6920 (N_6920,N_3880,N_1325);
xor U6921 (N_6921,N_3788,N_3268);
nor U6922 (N_6922,N_1433,N_3895);
or U6923 (N_6923,N_3156,N_2713);
and U6924 (N_6924,N_2382,N_2670);
xor U6925 (N_6925,N_1,N_2671);
xor U6926 (N_6926,N_3760,N_51);
and U6927 (N_6927,N_2008,N_78);
nor U6928 (N_6928,N_2027,N_3631);
and U6929 (N_6929,N_3172,N_1314);
nor U6930 (N_6930,N_819,N_1022);
and U6931 (N_6931,N_320,N_547);
and U6932 (N_6932,N_4557,N_3988);
nor U6933 (N_6933,N_204,N_4086);
xnor U6934 (N_6934,N_4345,N_2656);
or U6935 (N_6935,N_3884,N_394);
nand U6936 (N_6936,N_3560,N_1821);
nor U6937 (N_6937,N_980,N_4411);
or U6938 (N_6938,N_4949,N_2013);
and U6939 (N_6939,N_3812,N_2297);
nor U6940 (N_6940,N_2090,N_2944);
and U6941 (N_6941,N_723,N_3472);
nor U6942 (N_6942,N_1172,N_4847);
or U6943 (N_6943,N_3894,N_177);
and U6944 (N_6944,N_3484,N_4263);
or U6945 (N_6945,N_1136,N_4615);
and U6946 (N_6946,N_3188,N_4542);
xnor U6947 (N_6947,N_4595,N_3096);
nor U6948 (N_6948,N_697,N_4060);
and U6949 (N_6949,N_185,N_3333);
nor U6950 (N_6950,N_80,N_1249);
nor U6951 (N_6951,N_3675,N_4404);
and U6952 (N_6952,N_1094,N_1998);
and U6953 (N_6953,N_521,N_647);
or U6954 (N_6954,N_1983,N_313);
and U6955 (N_6955,N_526,N_4580);
nand U6956 (N_6956,N_1086,N_4556);
nand U6957 (N_6957,N_3100,N_557);
xnor U6958 (N_6958,N_2260,N_4939);
nand U6959 (N_6959,N_379,N_4147);
nor U6960 (N_6960,N_3239,N_2286);
nand U6961 (N_6961,N_3310,N_2804);
nor U6962 (N_6962,N_3457,N_2261);
and U6963 (N_6963,N_4035,N_3353);
xor U6964 (N_6964,N_4282,N_218);
nor U6965 (N_6965,N_2774,N_4011);
nor U6966 (N_6966,N_3337,N_2803);
and U6967 (N_6967,N_3476,N_1597);
nand U6968 (N_6968,N_3332,N_4975);
or U6969 (N_6969,N_986,N_309);
nand U6970 (N_6970,N_3122,N_4484);
xnor U6971 (N_6971,N_1878,N_3570);
and U6972 (N_6972,N_2354,N_3742);
nor U6973 (N_6973,N_1556,N_4657);
or U6974 (N_6974,N_1805,N_4460);
or U6975 (N_6975,N_4143,N_3264);
and U6976 (N_6976,N_4527,N_2840);
nand U6977 (N_6977,N_2488,N_3665);
nand U6978 (N_6978,N_4222,N_237);
or U6979 (N_6979,N_3605,N_1336);
nor U6980 (N_6980,N_3980,N_91);
nor U6981 (N_6981,N_3555,N_745);
nand U6982 (N_6982,N_709,N_2881);
nand U6983 (N_6983,N_3058,N_242);
or U6984 (N_6984,N_4569,N_1774);
nor U6985 (N_6985,N_3921,N_3068);
nand U6986 (N_6986,N_3048,N_3166);
and U6987 (N_6987,N_1671,N_2628);
xor U6988 (N_6988,N_3699,N_1933);
nor U6989 (N_6989,N_1173,N_814);
and U6990 (N_6990,N_4583,N_1010);
or U6991 (N_6991,N_851,N_4707);
and U6992 (N_6992,N_3495,N_2817);
and U6993 (N_6993,N_3647,N_2805);
nand U6994 (N_6994,N_2505,N_4350);
nand U6995 (N_6995,N_593,N_462);
or U6996 (N_6996,N_4054,N_165);
nor U6997 (N_6997,N_346,N_848);
nand U6998 (N_6998,N_4094,N_1397);
nor U6999 (N_6999,N_4407,N_2878);
or U7000 (N_7000,N_3389,N_2814);
nand U7001 (N_7001,N_4200,N_3030);
xor U7002 (N_7002,N_947,N_3752);
nor U7003 (N_7003,N_2869,N_190);
xor U7004 (N_7004,N_1524,N_2167);
xnor U7005 (N_7005,N_511,N_3181);
xnor U7006 (N_7006,N_1467,N_4968);
nand U7007 (N_7007,N_525,N_3441);
nor U7008 (N_7008,N_3393,N_778);
or U7009 (N_7009,N_1984,N_2737);
or U7010 (N_7010,N_4536,N_1498);
nor U7011 (N_7011,N_4495,N_4601);
or U7012 (N_7012,N_3789,N_3566);
nand U7013 (N_7013,N_1746,N_226);
nor U7014 (N_7014,N_3444,N_1547);
nor U7015 (N_7015,N_3320,N_288);
nor U7016 (N_7016,N_2889,N_1786);
nand U7017 (N_7017,N_2230,N_541);
xnor U7018 (N_7018,N_4134,N_3622);
and U7019 (N_7019,N_2823,N_2641);
nand U7020 (N_7020,N_562,N_2085);
nand U7021 (N_7021,N_1715,N_4817);
or U7022 (N_7022,N_4240,N_1576);
xor U7023 (N_7023,N_4065,N_2610);
nand U7024 (N_7024,N_2440,N_3815);
and U7025 (N_7025,N_1797,N_2942);
xnor U7026 (N_7026,N_4217,N_2474);
xor U7027 (N_7027,N_2222,N_4927);
xor U7028 (N_7028,N_900,N_3260);
and U7029 (N_7029,N_3703,N_2492);
nor U7030 (N_7030,N_2988,N_2721);
and U7031 (N_7031,N_4399,N_1976);
xnor U7032 (N_7032,N_4137,N_3913);
nand U7033 (N_7033,N_2813,N_2548);
nand U7034 (N_7034,N_1617,N_4652);
nor U7035 (N_7035,N_1291,N_2538);
or U7036 (N_7036,N_2646,N_87);
and U7037 (N_7037,N_3545,N_2593);
and U7038 (N_7038,N_450,N_2851);
or U7039 (N_7039,N_75,N_3878);
or U7040 (N_7040,N_1293,N_1521);
nor U7041 (N_7041,N_895,N_830);
nor U7042 (N_7042,N_3551,N_3442);
and U7043 (N_7043,N_1748,N_483);
nand U7044 (N_7044,N_4245,N_4999);
and U7045 (N_7045,N_1868,N_4293);
xnor U7046 (N_7046,N_2614,N_4234);
nor U7047 (N_7047,N_2844,N_4603);
and U7048 (N_7048,N_1904,N_2163);
and U7049 (N_7049,N_2076,N_4579);
nand U7050 (N_7050,N_362,N_3685);
nor U7051 (N_7051,N_4574,N_1627);
and U7052 (N_7052,N_381,N_3049);
nor U7053 (N_7053,N_2137,N_2188);
nor U7054 (N_7054,N_4564,N_102);
xor U7055 (N_7055,N_577,N_2442);
xnor U7056 (N_7056,N_503,N_1252);
or U7057 (N_7057,N_68,N_56);
nor U7058 (N_7058,N_1073,N_952);
and U7059 (N_7059,N_2118,N_3314);
or U7060 (N_7060,N_2282,N_1882);
and U7061 (N_7061,N_2289,N_2480);
or U7062 (N_7062,N_2267,N_2042);
and U7063 (N_7063,N_3659,N_838);
nor U7064 (N_7064,N_1912,N_4988);
nand U7065 (N_7065,N_2157,N_3334);
xor U7066 (N_7066,N_1426,N_896);
and U7067 (N_7067,N_1168,N_189);
nor U7068 (N_7068,N_4755,N_2489);
nand U7069 (N_7069,N_686,N_861);
nor U7070 (N_7070,N_676,N_4746);
xnor U7071 (N_7071,N_2990,N_2410);
nor U7072 (N_7072,N_4441,N_1810);
or U7073 (N_7073,N_1236,N_1496);
xnor U7074 (N_7074,N_3912,N_958);
and U7075 (N_7075,N_2294,N_2624);
xor U7076 (N_7076,N_4387,N_4818);
or U7077 (N_7077,N_3824,N_4148);
xnor U7078 (N_7078,N_500,N_1374);
nor U7079 (N_7079,N_3571,N_62);
xnor U7080 (N_7080,N_4483,N_4361);
nand U7081 (N_7081,N_418,N_4798);
and U7082 (N_7082,N_3860,N_2861);
nor U7083 (N_7083,N_2971,N_3664);
nand U7084 (N_7084,N_1836,N_260);
nor U7085 (N_7085,N_1608,N_1840);
or U7086 (N_7086,N_225,N_2296);
xor U7087 (N_7087,N_3775,N_259);
and U7088 (N_7088,N_1994,N_1161);
nand U7089 (N_7089,N_4674,N_2559);
and U7090 (N_7090,N_862,N_2436);
nand U7091 (N_7091,N_2408,N_2370);
nand U7092 (N_7092,N_1403,N_3992);
or U7093 (N_7093,N_4577,N_2151);
or U7094 (N_7094,N_1981,N_1987);
nand U7095 (N_7095,N_664,N_4157);
nand U7096 (N_7096,N_3107,N_3599);
and U7097 (N_7097,N_4069,N_3501);
nor U7098 (N_7098,N_4515,N_426);
xnor U7099 (N_7099,N_4519,N_1845);
nor U7100 (N_7100,N_2218,N_656);
and U7101 (N_7101,N_2719,N_1736);
xor U7102 (N_7102,N_154,N_3074);
xnor U7103 (N_7103,N_3419,N_936);
nand U7104 (N_7104,N_2707,N_482);
xnor U7105 (N_7105,N_2590,N_3398);
or U7106 (N_7106,N_3086,N_2306);
and U7107 (N_7107,N_1570,N_3286);
xor U7108 (N_7108,N_4666,N_3981);
nand U7109 (N_7109,N_1791,N_3349);
nor U7110 (N_7110,N_1300,N_4284);
xnor U7111 (N_7111,N_60,N_4104);
nor U7112 (N_7112,N_4890,N_1744);
or U7113 (N_7113,N_2233,N_1434);
or U7114 (N_7114,N_4605,N_2075);
nor U7115 (N_7115,N_1326,N_1355);
xnor U7116 (N_7116,N_2661,N_4794);
nor U7117 (N_7117,N_1548,N_3467);
xnor U7118 (N_7118,N_1093,N_2831);
nand U7119 (N_7119,N_1497,N_3606);
or U7120 (N_7120,N_4259,N_4440);
nand U7121 (N_7121,N_1762,N_4472);
and U7122 (N_7122,N_2197,N_1694);
xnor U7123 (N_7123,N_4963,N_341);
xnor U7124 (N_7124,N_4619,N_1202);
or U7125 (N_7125,N_3705,N_1573);
nor U7126 (N_7126,N_3882,N_2745);
nand U7127 (N_7127,N_1261,N_3009);
xnor U7128 (N_7128,N_4986,N_3280);
and U7129 (N_7129,N_4555,N_370);
nor U7130 (N_7130,N_2221,N_2945);
nor U7131 (N_7131,N_2133,N_4064);
or U7132 (N_7132,N_351,N_2638);
nand U7133 (N_7133,N_1174,N_2515);
or U7134 (N_7134,N_3176,N_305);
and U7135 (N_7135,N_1600,N_3248);
nor U7136 (N_7136,N_1956,N_1049);
nand U7137 (N_7137,N_4552,N_3946);
xnor U7138 (N_7138,N_4187,N_1254);
nor U7139 (N_7139,N_4391,N_2227);
nand U7140 (N_7140,N_991,N_3447);
xor U7141 (N_7141,N_3582,N_4651);
nand U7142 (N_7142,N_4973,N_2571);
nor U7143 (N_7143,N_1120,N_3865);
xnor U7144 (N_7144,N_1795,N_3817);
or U7145 (N_7145,N_4486,N_4602);
nand U7146 (N_7146,N_2611,N_2330);
xnor U7147 (N_7147,N_4405,N_1009);
nand U7148 (N_7148,N_2673,N_3402);
xnor U7149 (N_7149,N_1028,N_3482);
nand U7150 (N_7150,N_4135,N_2812);
nand U7151 (N_7151,N_4656,N_3094);
nand U7152 (N_7152,N_1153,N_658);
xnor U7153 (N_7153,N_2441,N_2977);
nand U7154 (N_7154,N_2893,N_4782);
and U7155 (N_7155,N_4784,N_4594);
nor U7156 (N_7156,N_1942,N_187);
and U7157 (N_7157,N_1755,N_1665);
and U7158 (N_7158,N_3234,N_4905);
or U7159 (N_7159,N_1952,N_99);
nor U7160 (N_7160,N_1171,N_2963);
xnor U7161 (N_7161,N_3984,N_3906);
nor U7162 (N_7162,N_3028,N_1225);
or U7163 (N_7163,N_1476,N_3381);
and U7164 (N_7164,N_355,N_1683);
and U7165 (N_7165,N_3133,N_1209);
nor U7166 (N_7166,N_2466,N_378);
nor U7167 (N_7167,N_1644,N_4213);
and U7168 (N_7168,N_687,N_280);
nor U7169 (N_7169,N_1460,N_3229);
or U7170 (N_7170,N_3169,N_3035);
or U7171 (N_7171,N_587,N_182);
and U7172 (N_7172,N_2241,N_3886);
xnor U7173 (N_7173,N_4492,N_4744);
xor U7174 (N_7174,N_1277,N_468);
nor U7175 (N_7175,N_1157,N_3586);
nor U7176 (N_7176,N_4816,N_4298);
nand U7177 (N_7177,N_865,N_4386);
nor U7178 (N_7178,N_1007,N_4379);
nor U7179 (N_7179,N_1268,N_4166);
xor U7180 (N_7180,N_2456,N_1179);
or U7181 (N_7181,N_784,N_933);
and U7182 (N_7182,N_4161,N_1894);
and U7183 (N_7183,N_2123,N_1789);
xnor U7184 (N_7184,N_2346,N_404);
xor U7185 (N_7185,N_2243,N_4150);
nand U7186 (N_7186,N_3881,N_1907);
and U7187 (N_7187,N_1350,N_1084);
nor U7188 (N_7188,N_4081,N_2734);
or U7189 (N_7189,N_924,N_1159);
and U7190 (N_7190,N_2923,N_3124);
and U7191 (N_7191,N_3299,N_421);
nor U7192 (N_7192,N_4433,N_186);
or U7193 (N_7193,N_337,N_240);
xor U7194 (N_7194,N_3825,N_2322);
xnor U7195 (N_7195,N_141,N_1472);
and U7196 (N_7196,N_3377,N_433);
and U7197 (N_7197,N_876,N_2109);
or U7198 (N_7198,N_3835,N_2654);
nor U7199 (N_7199,N_444,N_4566);
nand U7200 (N_7200,N_3307,N_2210);
nor U7201 (N_7201,N_1489,N_4014);
or U7202 (N_7202,N_3295,N_1926);
nor U7203 (N_7203,N_1305,N_192);
nor U7204 (N_7204,N_128,N_4688);
xnor U7205 (N_7205,N_2381,N_2645);
or U7206 (N_7206,N_2213,N_2299);
or U7207 (N_7207,N_205,N_1112);
nand U7208 (N_7208,N_2735,N_2980);
and U7209 (N_7209,N_2580,N_545);
and U7210 (N_7210,N_575,N_1475);
and U7211 (N_7211,N_1226,N_553);
nor U7212 (N_7212,N_3493,N_903);
and U7213 (N_7213,N_3267,N_1727);
xnor U7214 (N_7214,N_465,N_2069);
or U7215 (N_7215,N_1319,N_233);
and U7216 (N_7216,N_2791,N_412);
or U7217 (N_7217,N_4458,N_3223);
nand U7218 (N_7218,N_4130,N_491);
or U7219 (N_7219,N_261,N_198);
nand U7220 (N_7220,N_451,N_23);
nor U7221 (N_7221,N_599,N_399);
nand U7222 (N_7222,N_4826,N_55);
nand U7223 (N_7223,N_4406,N_1365);
or U7224 (N_7224,N_4125,N_2226);
nand U7225 (N_7225,N_4106,N_3885);
xnor U7226 (N_7226,N_2199,N_2087);
nand U7227 (N_7227,N_3796,N_3135);
nand U7228 (N_7228,N_340,N_1899);
nand U7229 (N_7229,N_3388,N_1941);
nand U7230 (N_7230,N_4607,N_2217);
and U7231 (N_7231,N_2338,N_552);
and U7232 (N_7232,N_4336,N_3093);
nand U7233 (N_7233,N_152,N_3175);
xor U7234 (N_7234,N_453,N_2798);
nand U7235 (N_7235,N_2934,N_2839);
or U7236 (N_7236,N_114,N_1718);
or U7237 (N_7237,N_4047,N_3163);
or U7238 (N_7238,N_1441,N_631);
xor U7239 (N_7239,N_3019,N_4813);
nor U7240 (N_7240,N_1678,N_1215);
or U7241 (N_7241,N_3634,N_1822);
nor U7242 (N_7242,N_942,N_1639);
and U7243 (N_7243,N_517,N_1893);
or U7244 (N_7244,N_2937,N_1347);
or U7245 (N_7245,N_311,N_4236);
nor U7246 (N_7246,N_3127,N_4409);
nor U7247 (N_7247,N_649,N_3410);
and U7248 (N_7248,N_3938,N_4612);
nand U7249 (N_7249,N_363,N_3786);
nand U7250 (N_7250,N_274,N_4031);
nand U7251 (N_7251,N_1134,N_3707);
or U7252 (N_7252,N_95,N_300);
and U7253 (N_7253,N_2483,N_3771);
nor U7254 (N_7254,N_4751,N_1459);
nand U7255 (N_7255,N_1862,N_911);
or U7256 (N_7256,N_594,N_2391);
nand U7257 (N_7257,N_1302,N_2273);
and U7258 (N_7258,N_1723,N_661);
nand U7259 (N_7259,N_1771,N_1247);
xor U7260 (N_7260,N_67,N_2743);
nand U7261 (N_7261,N_4523,N_2016);
nand U7262 (N_7262,N_1880,N_262);
xor U7263 (N_7263,N_3165,N_2396);
xnor U7264 (N_7264,N_3232,N_2375);
nor U7265 (N_7265,N_2186,N_122);
nor U7266 (N_7266,N_1980,N_354);
xor U7267 (N_7267,N_847,N_1946);
and U7268 (N_7268,N_3759,N_584);
and U7269 (N_7269,N_2211,N_1380);
nand U7270 (N_7270,N_4728,N_2310);
nor U7271 (N_7271,N_1223,N_3064);
and U7272 (N_7272,N_1309,N_3741);
or U7273 (N_7273,N_4439,N_3655);
xor U7274 (N_7274,N_42,N_1849);
xor U7275 (N_7275,N_874,N_4255);
or U7276 (N_7276,N_624,N_1684);
or U7277 (N_7277,N_3205,N_1025);
nand U7278 (N_7278,N_2757,N_1488);
and U7279 (N_7279,N_863,N_825);
and U7280 (N_7280,N_1619,N_2770);
xnor U7281 (N_7281,N_3253,N_2680);
or U7282 (N_7282,N_4952,N_919);
xnor U7283 (N_7283,N_976,N_3838);
nand U7284 (N_7284,N_4211,N_2672);
and U7285 (N_7285,N_2060,N_840);
nand U7286 (N_7286,N_1844,N_4983);
nand U7287 (N_7287,N_476,N_4131);
xor U7288 (N_7288,N_4967,N_4254);
xnor U7289 (N_7289,N_118,N_1250);
and U7290 (N_7290,N_1219,N_2111);
or U7291 (N_7291,N_3070,N_2453);
nand U7292 (N_7292,N_397,N_4588);
xnor U7293 (N_7293,N_3195,N_1528);
and U7294 (N_7294,N_3216,N_600);
xor U7295 (N_7295,N_1724,N_948);
nor U7296 (N_7296,N_1424,N_4220);
nor U7297 (N_7297,N_2360,N_4670);
nor U7298 (N_7298,N_2539,N_3641);
nand U7299 (N_7299,N_4414,N_3115);
nand U7300 (N_7300,N_964,N_1649);
nand U7301 (N_7301,N_3950,N_2724);
nand U7302 (N_7302,N_371,N_249);
nor U7303 (N_7303,N_2983,N_1070);
xnor U7304 (N_7304,N_4090,N_3532);
nor U7305 (N_7305,N_2976,N_4855);
nor U7306 (N_7306,N_4175,N_389);
xnor U7307 (N_7307,N_2397,N_3050);
and U7308 (N_7308,N_2995,N_3598);
nor U7309 (N_7309,N_3283,N_4960);
and U7310 (N_7310,N_478,N_4832);
xnor U7311 (N_7311,N_2395,N_582);
nor U7312 (N_7312,N_4079,N_2458);
nand U7313 (N_7313,N_2690,N_927);
xnor U7314 (N_7314,N_2960,N_3780);
and U7315 (N_7315,N_57,N_1288);
xor U7316 (N_7316,N_855,N_88);
and U7317 (N_7317,N_1016,N_4793);
or U7318 (N_7318,N_3038,N_2355);
and U7319 (N_7319,N_4820,N_3971);
nand U7320 (N_7320,N_4956,N_3522);
nand U7321 (N_7321,N_5,N_3536);
xor U7322 (N_7322,N_4329,N_4155);
or U7323 (N_7323,N_3716,N_1881);
nor U7324 (N_7324,N_595,N_428);
nand U7325 (N_7325,N_2465,N_1131);
and U7326 (N_7326,N_2020,N_3418);
nand U7327 (N_7327,N_2597,N_4431);
nor U7328 (N_7328,N_598,N_4767);
nor U7329 (N_7329,N_2999,N_213);
nor U7330 (N_7330,N_4057,N_58);
nand U7331 (N_7331,N_1673,N_4128);
and U7332 (N_7332,N_2209,N_2836);
and U7333 (N_7333,N_1545,N_1705);
nand U7334 (N_7334,N_2648,N_4752);
and U7335 (N_7335,N_2473,N_4848);
or U7336 (N_7336,N_3480,N_3487);
nand U7337 (N_7337,N_484,N_3673);
nor U7338 (N_7338,N_1222,N_1538);
or U7339 (N_7339,N_1963,N_3033);
and U7340 (N_7340,N_3144,N_3591);
nor U7341 (N_7341,N_628,N_4589);
xnor U7342 (N_7342,N_2235,N_4096);
and U7343 (N_7343,N_718,N_1873);
and U7344 (N_7344,N_2125,N_4052);
and U7345 (N_7345,N_884,N_3428);
nor U7346 (N_7346,N_860,N_823);
xnor U7347 (N_7347,N_3010,N_2140);
nor U7348 (N_7348,N_850,N_1590);
nor U7349 (N_7349,N_72,N_3358);
or U7350 (N_7350,N_3425,N_1280);
nor U7351 (N_7351,N_839,N_4548);
xnor U7352 (N_7352,N_881,N_4824);
nand U7353 (N_7353,N_2392,N_1378);
or U7354 (N_7354,N_4498,N_3818);
nor U7355 (N_7355,N_657,N_932);
nor U7356 (N_7356,N_3473,N_4434);
nor U7357 (N_7357,N_4396,N_1533);
or U7358 (N_7358,N_2117,N_956);
nand U7359 (N_7359,N_90,N_3568);
xnor U7360 (N_7360,N_3511,N_4852);
xor U7361 (N_7361,N_3636,N_2400);
nand U7362 (N_7362,N_3542,N_2906);
or U7363 (N_7363,N_4420,N_2182);
nor U7364 (N_7364,N_4291,N_2728);
nand U7365 (N_7365,N_1167,N_3750);
xnor U7366 (N_7366,N_3831,N_232);
xnor U7367 (N_7367,N_515,N_1354);
xor U7368 (N_7368,N_4876,N_3963);
nand U7369 (N_7369,N_4265,N_2315);
or U7370 (N_7370,N_597,N_1431);
xnor U7371 (N_7371,N_722,N_1986);
and U7372 (N_7372,N_3749,N_1119);
or U7373 (N_7373,N_145,N_2155);
or U7374 (N_7374,N_2240,N_3530);
and U7375 (N_7375,N_905,N_4626);
or U7376 (N_7376,N_4232,N_606);
nor U7377 (N_7377,N_1611,N_4640);
and U7378 (N_7378,N_2810,N_324);
and U7379 (N_7379,N_2393,N_46);
nor U7380 (N_7380,N_518,N_4658);
xor U7381 (N_7381,N_270,N_1474);
nand U7382 (N_7382,N_40,N_2287);
xnor U7383 (N_7383,N_813,N_2452);
and U7384 (N_7384,N_4444,N_3051);
or U7385 (N_7385,N_3868,N_3386);
nand U7386 (N_7386,N_535,N_3845);
xor U7387 (N_7387,N_3821,N_2107);
and U7388 (N_7388,N_2341,N_1055);
xor U7389 (N_7389,N_37,N_2616);
and U7390 (N_7390,N_3269,N_2270);
nor U7391 (N_7391,N_907,N_4738);
or U7392 (N_7392,N_1801,N_3063);
or U7393 (N_7393,N_2863,N_1356);
nor U7394 (N_7394,N_1543,N_4452);
and U7395 (N_7395,N_1145,N_2371);
xor U7396 (N_7396,N_125,N_4308);
or U7397 (N_7397,N_3604,N_1057);
or U7398 (N_7398,N_1869,N_3723);
nand U7399 (N_7399,N_2936,N_3713);
and U7400 (N_7400,N_1971,N_4951);
nor U7401 (N_7401,N_2254,N_1599);
nor U7402 (N_7402,N_853,N_4554);
xor U7403 (N_7403,N_4671,N_3024);
nor U7404 (N_7404,N_2752,N_3525);
nor U7405 (N_7405,N_2097,N_1689);
nand U7406 (N_7406,N_2485,N_2108);
or U7407 (N_7407,N_4377,N_219);
nand U7408 (N_7408,N_776,N_831);
or U7409 (N_7409,N_558,N_3415);
nand U7410 (N_7410,N_3246,N_3121);
and U7411 (N_7411,N_2026,N_893);
xnor U7412 (N_7412,N_1091,N_1969);
nor U7413 (N_7413,N_151,N_4314);
nand U7414 (N_7414,N_1464,N_4323);
nor U7415 (N_7415,N_4283,N_3437);
nor U7416 (N_7416,N_3892,N_4430);
xor U7417 (N_7417,N_3157,N_2220);
xnor U7418 (N_7418,N_2954,N_1717);
or U7419 (N_7419,N_420,N_3795);
nor U7420 (N_7420,N_719,N_1088);
xor U7421 (N_7421,N_2577,N_2776);
or U7422 (N_7422,N_44,N_4083);
or U7423 (N_7423,N_818,N_3803);
nand U7424 (N_7424,N_820,N_4201);
or U7425 (N_7425,N_571,N_3721);
nor U7426 (N_7426,N_1271,N_2847);
nor U7427 (N_7427,N_2829,N_3110);
and U7428 (N_7428,N_2412,N_4721);
nand U7429 (N_7429,N_1218,N_2065);
and U7430 (N_7430,N_2793,N_3112);
nor U7431 (N_7431,N_4237,N_1970);
nor U7432 (N_7432,N_1368,N_1274);
xor U7433 (N_7433,N_4275,N_2348);
nor U7434 (N_7434,N_1231,N_2753);
nor U7435 (N_7435,N_3161,N_4445);
or U7436 (N_7436,N_209,N_3342);
and U7437 (N_7437,N_3652,N_4989);
nand U7438 (N_7438,N_3720,N_4132);
nand U7439 (N_7439,N_1752,N_302);
xnor U7440 (N_7440,N_3823,N_94);
nor U7441 (N_7441,N_1203,N_4678);
or U7442 (N_7442,N_1281,N_4972);
xnor U7443 (N_7443,N_3558,N_1753);
nor U7444 (N_7444,N_1150,N_611);
and U7445 (N_7445,N_1447,N_3203);
or U7446 (N_7446,N_1751,N_4931);
or U7447 (N_7447,N_1328,N_1914);
or U7448 (N_7448,N_1053,N_2558);
xnor U7449 (N_7449,N_4050,N_306);
and U7450 (N_7450,N_4372,N_3828);
nand U7451 (N_7451,N_4692,N_806);
xor U7452 (N_7452,N_796,N_2973);
or U7453 (N_7453,N_2247,N_760);
nand U7454 (N_7454,N_713,N_3781);
xnor U7455 (N_7455,N_2399,N_272);
or U7456 (N_7456,N_2970,N_3424);
nor U7457 (N_7457,N_1760,N_4225);
nand U7458 (N_7458,N_3959,N_4092);
xor U7459 (N_7459,N_913,N_2602);
xor U7460 (N_7460,N_2969,N_39);
nand U7461 (N_7461,N_3171,N_1697);
nand U7462 (N_7462,N_3270,N_4327);
or U7463 (N_7463,N_2068,N_3018);
nor U7464 (N_7464,N_2865,N_1081);
nand U7465 (N_7465,N_169,N_3814);
nor U7466 (N_7466,N_342,N_1949);
and U7467 (N_7467,N_2930,N_3574);
and U7468 (N_7468,N_3928,N_4270);
and U7469 (N_7469,N_566,N_191);
xnor U7470 (N_7470,N_4567,N_2154);
nor U7471 (N_7471,N_2809,N_2605);
xnor U7472 (N_7472,N_3186,N_3954);
and U7473 (N_7473,N_1177,N_1193);
nor U7474 (N_7474,N_3710,N_1102);
nor U7475 (N_7475,N_1232,N_1574);
nand U7476 (N_7476,N_4698,N_934);
and U7477 (N_7477,N_4266,N_642);
nand U7478 (N_7478,N_344,N_1950);
xnor U7479 (N_7479,N_730,N_1861);
nor U7480 (N_7480,N_4829,N_4087);
and U7481 (N_7481,N_4026,N_119);
and U7482 (N_7482,N_3520,N_4885);
xnor U7483 (N_7483,N_1149,N_3378);
or U7484 (N_7484,N_3029,N_3296);
and U7485 (N_7485,N_529,N_2773);
nor U7486 (N_7486,N_3977,N_2245);
xnor U7487 (N_7487,N_36,N_551);
nor U7488 (N_7488,N_2142,N_1298);
nand U7489 (N_7489,N_1641,N_3554);
nand U7490 (N_7490,N_3829,N_875);
nand U7491 (N_7491,N_2631,N_2113);
xnor U7492 (N_7492,N_1329,N_3201);
or U7493 (N_7493,N_372,N_3743);
and U7494 (N_7494,N_2553,N_3956);
xor U7495 (N_7495,N_2207,N_764);
nor U7496 (N_7496,N_1732,N_1935);
xor U7497 (N_7497,N_1335,N_1382);
nor U7498 (N_7498,N_2325,N_229);
nand U7499 (N_7499,N_4779,N_2694);
or U7500 (N_7500,N_1225,N_3856);
nor U7501 (N_7501,N_4092,N_3165);
xnor U7502 (N_7502,N_4326,N_3241);
xor U7503 (N_7503,N_3122,N_2108);
xnor U7504 (N_7504,N_1983,N_856);
nand U7505 (N_7505,N_1239,N_10);
nand U7506 (N_7506,N_4439,N_4414);
nand U7507 (N_7507,N_1527,N_3780);
or U7508 (N_7508,N_3059,N_1136);
nand U7509 (N_7509,N_4173,N_185);
xor U7510 (N_7510,N_1131,N_3461);
nand U7511 (N_7511,N_3703,N_2212);
nor U7512 (N_7512,N_1759,N_4951);
or U7513 (N_7513,N_3095,N_1293);
or U7514 (N_7514,N_3912,N_4055);
nand U7515 (N_7515,N_3206,N_1511);
xnor U7516 (N_7516,N_2779,N_274);
xor U7517 (N_7517,N_2798,N_3679);
nand U7518 (N_7518,N_4514,N_3720);
and U7519 (N_7519,N_2300,N_1532);
nand U7520 (N_7520,N_3595,N_1893);
nand U7521 (N_7521,N_3831,N_3993);
nand U7522 (N_7522,N_3878,N_4504);
xor U7523 (N_7523,N_1955,N_102);
xnor U7524 (N_7524,N_2151,N_270);
xor U7525 (N_7525,N_1394,N_2326);
nor U7526 (N_7526,N_3295,N_4194);
and U7527 (N_7527,N_978,N_1190);
and U7528 (N_7528,N_3576,N_2077);
xor U7529 (N_7529,N_186,N_1738);
xnor U7530 (N_7530,N_1241,N_4582);
and U7531 (N_7531,N_2962,N_3233);
nand U7532 (N_7532,N_2543,N_2699);
or U7533 (N_7533,N_3336,N_2363);
or U7534 (N_7534,N_284,N_4301);
and U7535 (N_7535,N_10,N_3531);
or U7536 (N_7536,N_4965,N_3256);
or U7537 (N_7537,N_1446,N_4448);
xor U7538 (N_7538,N_1836,N_1887);
xnor U7539 (N_7539,N_1916,N_1209);
or U7540 (N_7540,N_4305,N_210);
nand U7541 (N_7541,N_2808,N_553);
or U7542 (N_7542,N_838,N_3539);
nand U7543 (N_7543,N_3550,N_4473);
nor U7544 (N_7544,N_3184,N_4659);
and U7545 (N_7545,N_3965,N_4710);
or U7546 (N_7546,N_4103,N_3047);
nor U7547 (N_7547,N_1349,N_3264);
nand U7548 (N_7548,N_3469,N_1272);
and U7549 (N_7549,N_1678,N_3765);
nor U7550 (N_7550,N_3796,N_4476);
or U7551 (N_7551,N_2071,N_1506);
and U7552 (N_7552,N_397,N_4877);
nand U7553 (N_7553,N_2449,N_3905);
nand U7554 (N_7554,N_4343,N_3114);
or U7555 (N_7555,N_4745,N_4746);
and U7556 (N_7556,N_1524,N_4238);
or U7557 (N_7557,N_3941,N_1580);
xnor U7558 (N_7558,N_631,N_2478);
or U7559 (N_7559,N_4243,N_1673);
or U7560 (N_7560,N_232,N_3802);
and U7561 (N_7561,N_394,N_1273);
xor U7562 (N_7562,N_2525,N_1351);
xnor U7563 (N_7563,N_1179,N_806);
or U7564 (N_7564,N_4080,N_923);
or U7565 (N_7565,N_2332,N_1094);
nand U7566 (N_7566,N_978,N_3029);
and U7567 (N_7567,N_887,N_4267);
nand U7568 (N_7568,N_1435,N_571);
or U7569 (N_7569,N_3781,N_2525);
or U7570 (N_7570,N_1883,N_4888);
and U7571 (N_7571,N_2222,N_2744);
xor U7572 (N_7572,N_2213,N_4850);
nand U7573 (N_7573,N_3033,N_2914);
nand U7574 (N_7574,N_2490,N_2148);
nand U7575 (N_7575,N_4378,N_2822);
xor U7576 (N_7576,N_1346,N_700);
nand U7577 (N_7577,N_4955,N_3343);
nand U7578 (N_7578,N_2427,N_1947);
xnor U7579 (N_7579,N_3288,N_4017);
xnor U7580 (N_7580,N_356,N_2385);
or U7581 (N_7581,N_2134,N_1125);
or U7582 (N_7582,N_3420,N_4513);
xnor U7583 (N_7583,N_2024,N_1123);
or U7584 (N_7584,N_187,N_3982);
xnor U7585 (N_7585,N_3069,N_2783);
or U7586 (N_7586,N_4018,N_3492);
or U7587 (N_7587,N_3868,N_1042);
xor U7588 (N_7588,N_2029,N_1136);
xnor U7589 (N_7589,N_4500,N_1561);
nand U7590 (N_7590,N_984,N_3656);
xor U7591 (N_7591,N_4146,N_4514);
nor U7592 (N_7592,N_3266,N_4304);
nor U7593 (N_7593,N_3252,N_3395);
nand U7594 (N_7594,N_4248,N_1317);
or U7595 (N_7595,N_2850,N_722);
and U7596 (N_7596,N_304,N_3719);
nand U7597 (N_7597,N_4023,N_3285);
or U7598 (N_7598,N_3398,N_2238);
nor U7599 (N_7599,N_3021,N_2783);
xor U7600 (N_7600,N_4969,N_4023);
nand U7601 (N_7601,N_1945,N_3617);
or U7602 (N_7602,N_4750,N_2738);
and U7603 (N_7603,N_1454,N_428);
xor U7604 (N_7604,N_1224,N_715);
and U7605 (N_7605,N_2724,N_4699);
nor U7606 (N_7606,N_116,N_4809);
nor U7607 (N_7607,N_4428,N_2156);
and U7608 (N_7608,N_2459,N_4846);
or U7609 (N_7609,N_4864,N_2406);
nand U7610 (N_7610,N_974,N_3522);
nor U7611 (N_7611,N_955,N_2858);
or U7612 (N_7612,N_8,N_3687);
nand U7613 (N_7613,N_1385,N_4093);
or U7614 (N_7614,N_3291,N_2279);
nor U7615 (N_7615,N_4572,N_1679);
or U7616 (N_7616,N_1011,N_3220);
nor U7617 (N_7617,N_307,N_2094);
or U7618 (N_7618,N_137,N_1182);
xnor U7619 (N_7619,N_2982,N_1264);
and U7620 (N_7620,N_3143,N_4494);
nor U7621 (N_7621,N_1359,N_2202);
nand U7622 (N_7622,N_3866,N_1337);
nand U7623 (N_7623,N_2406,N_1875);
or U7624 (N_7624,N_2180,N_4025);
nand U7625 (N_7625,N_1285,N_4410);
nand U7626 (N_7626,N_4525,N_745);
or U7627 (N_7627,N_4293,N_1476);
xnor U7628 (N_7628,N_869,N_2856);
xor U7629 (N_7629,N_1239,N_1394);
and U7630 (N_7630,N_386,N_3818);
and U7631 (N_7631,N_1081,N_2630);
nor U7632 (N_7632,N_2543,N_35);
or U7633 (N_7633,N_492,N_2048);
nor U7634 (N_7634,N_2077,N_3743);
xnor U7635 (N_7635,N_4379,N_4143);
xor U7636 (N_7636,N_3561,N_1533);
nand U7637 (N_7637,N_4999,N_1245);
nand U7638 (N_7638,N_4185,N_340);
xnor U7639 (N_7639,N_3233,N_3075);
xor U7640 (N_7640,N_1680,N_2220);
nor U7641 (N_7641,N_4900,N_3760);
and U7642 (N_7642,N_36,N_53);
and U7643 (N_7643,N_4687,N_2787);
nand U7644 (N_7644,N_2046,N_2658);
nor U7645 (N_7645,N_3098,N_1342);
and U7646 (N_7646,N_2972,N_3197);
or U7647 (N_7647,N_1037,N_3528);
xnor U7648 (N_7648,N_3786,N_2306);
nand U7649 (N_7649,N_34,N_1906);
or U7650 (N_7650,N_602,N_2848);
xor U7651 (N_7651,N_374,N_2825);
nor U7652 (N_7652,N_2621,N_3624);
or U7653 (N_7653,N_3717,N_4608);
or U7654 (N_7654,N_3100,N_488);
xor U7655 (N_7655,N_3642,N_4581);
and U7656 (N_7656,N_1869,N_3354);
or U7657 (N_7657,N_40,N_3236);
xor U7658 (N_7658,N_4534,N_4899);
and U7659 (N_7659,N_1863,N_1209);
and U7660 (N_7660,N_1227,N_2227);
or U7661 (N_7661,N_4596,N_725);
nand U7662 (N_7662,N_1997,N_994);
nor U7663 (N_7663,N_608,N_4027);
nand U7664 (N_7664,N_1853,N_3087);
xor U7665 (N_7665,N_4935,N_4628);
and U7666 (N_7666,N_645,N_4879);
nor U7667 (N_7667,N_328,N_103);
nor U7668 (N_7668,N_1935,N_4354);
nand U7669 (N_7669,N_615,N_1173);
or U7670 (N_7670,N_3068,N_1963);
and U7671 (N_7671,N_465,N_1978);
nand U7672 (N_7672,N_431,N_654);
or U7673 (N_7673,N_3744,N_1940);
and U7674 (N_7674,N_2530,N_2572);
and U7675 (N_7675,N_3450,N_2121);
and U7676 (N_7676,N_368,N_3700);
nand U7677 (N_7677,N_1631,N_4599);
nor U7678 (N_7678,N_3460,N_1046);
nand U7679 (N_7679,N_1529,N_3256);
or U7680 (N_7680,N_2152,N_1591);
and U7681 (N_7681,N_303,N_1875);
or U7682 (N_7682,N_454,N_579);
and U7683 (N_7683,N_169,N_2631);
nor U7684 (N_7684,N_528,N_146);
xnor U7685 (N_7685,N_4480,N_952);
and U7686 (N_7686,N_4341,N_1588);
or U7687 (N_7687,N_2497,N_1466);
nor U7688 (N_7688,N_1060,N_4627);
or U7689 (N_7689,N_4993,N_3731);
nor U7690 (N_7690,N_2338,N_675);
and U7691 (N_7691,N_4516,N_1342);
or U7692 (N_7692,N_1939,N_3017);
and U7693 (N_7693,N_466,N_4227);
or U7694 (N_7694,N_980,N_2943);
and U7695 (N_7695,N_607,N_3622);
nor U7696 (N_7696,N_1175,N_2535);
nor U7697 (N_7697,N_4550,N_4652);
xor U7698 (N_7698,N_4687,N_3003);
nor U7699 (N_7699,N_385,N_1065);
and U7700 (N_7700,N_3484,N_3634);
xor U7701 (N_7701,N_1157,N_584);
nand U7702 (N_7702,N_776,N_398);
nand U7703 (N_7703,N_2733,N_629);
xnor U7704 (N_7704,N_3376,N_3690);
or U7705 (N_7705,N_758,N_3624);
xnor U7706 (N_7706,N_4948,N_3240);
and U7707 (N_7707,N_589,N_2663);
nor U7708 (N_7708,N_1887,N_3696);
nor U7709 (N_7709,N_4368,N_653);
and U7710 (N_7710,N_3020,N_3295);
nand U7711 (N_7711,N_2345,N_2458);
and U7712 (N_7712,N_1669,N_1608);
xnor U7713 (N_7713,N_2882,N_678);
xnor U7714 (N_7714,N_363,N_3943);
nand U7715 (N_7715,N_1995,N_2525);
nand U7716 (N_7716,N_1329,N_2272);
nor U7717 (N_7717,N_198,N_4958);
and U7718 (N_7718,N_4130,N_481);
and U7719 (N_7719,N_3545,N_2959);
nand U7720 (N_7720,N_162,N_4878);
nand U7721 (N_7721,N_345,N_1552);
or U7722 (N_7722,N_1157,N_723);
and U7723 (N_7723,N_1563,N_4487);
and U7724 (N_7724,N_2643,N_2652);
nor U7725 (N_7725,N_3925,N_1101);
and U7726 (N_7726,N_4773,N_389);
and U7727 (N_7727,N_1828,N_2912);
xor U7728 (N_7728,N_3470,N_3349);
nor U7729 (N_7729,N_2952,N_3246);
and U7730 (N_7730,N_4006,N_1095);
xor U7731 (N_7731,N_1259,N_2482);
and U7732 (N_7732,N_2230,N_20);
and U7733 (N_7733,N_3060,N_1700);
nand U7734 (N_7734,N_1835,N_87);
xor U7735 (N_7735,N_2981,N_1231);
and U7736 (N_7736,N_1343,N_3573);
xor U7737 (N_7737,N_1441,N_893);
nand U7738 (N_7738,N_2026,N_2391);
or U7739 (N_7739,N_3425,N_107);
xor U7740 (N_7740,N_881,N_2827);
xor U7741 (N_7741,N_357,N_1469);
and U7742 (N_7742,N_3867,N_4579);
xor U7743 (N_7743,N_112,N_744);
or U7744 (N_7744,N_4098,N_580);
nor U7745 (N_7745,N_1055,N_2808);
nand U7746 (N_7746,N_4975,N_3910);
or U7747 (N_7747,N_2847,N_1444);
or U7748 (N_7748,N_2824,N_3620);
and U7749 (N_7749,N_1743,N_1335);
and U7750 (N_7750,N_787,N_3853);
and U7751 (N_7751,N_398,N_1286);
or U7752 (N_7752,N_2356,N_3215);
and U7753 (N_7753,N_4875,N_3037);
xnor U7754 (N_7754,N_1975,N_1004);
nand U7755 (N_7755,N_550,N_3689);
nor U7756 (N_7756,N_97,N_1266);
and U7757 (N_7757,N_600,N_2229);
nor U7758 (N_7758,N_424,N_1340);
or U7759 (N_7759,N_167,N_2993);
xor U7760 (N_7760,N_1127,N_3924);
nand U7761 (N_7761,N_1424,N_4045);
xor U7762 (N_7762,N_2843,N_2542);
and U7763 (N_7763,N_4966,N_3468);
xnor U7764 (N_7764,N_3998,N_1002);
and U7765 (N_7765,N_3960,N_178);
nand U7766 (N_7766,N_901,N_482);
or U7767 (N_7767,N_3674,N_1314);
nor U7768 (N_7768,N_1158,N_3468);
or U7769 (N_7769,N_2080,N_2530);
nand U7770 (N_7770,N_1373,N_654);
xnor U7771 (N_7771,N_2034,N_2526);
nor U7772 (N_7772,N_2067,N_3859);
or U7773 (N_7773,N_3016,N_2842);
nor U7774 (N_7774,N_1616,N_1810);
or U7775 (N_7775,N_787,N_3052);
and U7776 (N_7776,N_2230,N_1261);
nand U7777 (N_7777,N_4095,N_179);
and U7778 (N_7778,N_2953,N_3094);
nor U7779 (N_7779,N_2119,N_1122);
nor U7780 (N_7780,N_1652,N_4446);
nor U7781 (N_7781,N_4512,N_1068);
nor U7782 (N_7782,N_2754,N_4583);
nand U7783 (N_7783,N_2990,N_905);
and U7784 (N_7784,N_3883,N_491);
nand U7785 (N_7785,N_2703,N_2855);
nor U7786 (N_7786,N_2465,N_811);
nor U7787 (N_7787,N_3474,N_1874);
or U7788 (N_7788,N_4189,N_2161);
or U7789 (N_7789,N_2118,N_1907);
xnor U7790 (N_7790,N_1246,N_389);
nand U7791 (N_7791,N_1096,N_3386);
or U7792 (N_7792,N_283,N_3564);
nand U7793 (N_7793,N_4667,N_4122);
and U7794 (N_7794,N_1929,N_1756);
xnor U7795 (N_7795,N_4452,N_1199);
and U7796 (N_7796,N_3645,N_3395);
xor U7797 (N_7797,N_4718,N_2379);
nor U7798 (N_7798,N_1548,N_989);
nand U7799 (N_7799,N_4518,N_2025);
nand U7800 (N_7800,N_3328,N_4669);
or U7801 (N_7801,N_3875,N_3844);
or U7802 (N_7802,N_4789,N_2488);
xnor U7803 (N_7803,N_430,N_2745);
nor U7804 (N_7804,N_2883,N_1513);
nand U7805 (N_7805,N_2471,N_3193);
nor U7806 (N_7806,N_3750,N_1019);
and U7807 (N_7807,N_378,N_4183);
nor U7808 (N_7808,N_2641,N_3580);
or U7809 (N_7809,N_2453,N_1500);
nor U7810 (N_7810,N_3163,N_3917);
nor U7811 (N_7811,N_1951,N_3859);
xor U7812 (N_7812,N_4464,N_3979);
nand U7813 (N_7813,N_779,N_4012);
and U7814 (N_7814,N_4811,N_198);
or U7815 (N_7815,N_4655,N_264);
nor U7816 (N_7816,N_3340,N_448);
xor U7817 (N_7817,N_3792,N_1996);
and U7818 (N_7818,N_2185,N_3441);
nor U7819 (N_7819,N_1352,N_1728);
or U7820 (N_7820,N_48,N_3318);
and U7821 (N_7821,N_188,N_4178);
nor U7822 (N_7822,N_4885,N_470);
nand U7823 (N_7823,N_2739,N_2858);
or U7824 (N_7824,N_1500,N_860);
and U7825 (N_7825,N_4300,N_4403);
or U7826 (N_7826,N_872,N_1389);
or U7827 (N_7827,N_399,N_1918);
nand U7828 (N_7828,N_1443,N_2654);
nor U7829 (N_7829,N_2848,N_2832);
nor U7830 (N_7830,N_504,N_1707);
nand U7831 (N_7831,N_3783,N_3152);
and U7832 (N_7832,N_1232,N_4906);
and U7833 (N_7833,N_2813,N_3324);
xnor U7834 (N_7834,N_2871,N_3731);
and U7835 (N_7835,N_4632,N_2324);
or U7836 (N_7836,N_2052,N_3632);
nor U7837 (N_7837,N_666,N_785);
or U7838 (N_7838,N_4273,N_103);
xor U7839 (N_7839,N_4952,N_2614);
nand U7840 (N_7840,N_2351,N_3082);
xnor U7841 (N_7841,N_216,N_1750);
xor U7842 (N_7842,N_4491,N_3094);
nand U7843 (N_7843,N_3577,N_2021);
nand U7844 (N_7844,N_1230,N_4270);
or U7845 (N_7845,N_4300,N_178);
nand U7846 (N_7846,N_653,N_4117);
or U7847 (N_7847,N_2672,N_358);
nor U7848 (N_7848,N_137,N_2965);
and U7849 (N_7849,N_2496,N_2797);
nand U7850 (N_7850,N_1193,N_4583);
xor U7851 (N_7851,N_2903,N_736);
and U7852 (N_7852,N_4009,N_1112);
and U7853 (N_7853,N_281,N_443);
and U7854 (N_7854,N_4883,N_605);
nand U7855 (N_7855,N_2618,N_4303);
nor U7856 (N_7856,N_2148,N_3139);
and U7857 (N_7857,N_4880,N_350);
and U7858 (N_7858,N_2532,N_602);
nor U7859 (N_7859,N_4811,N_105);
xnor U7860 (N_7860,N_1445,N_797);
nand U7861 (N_7861,N_111,N_4691);
xnor U7862 (N_7862,N_2558,N_2559);
or U7863 (N_7863,N_779,N_1823);
or U7864 (N_7864,N_2582,N_2173);
and U7865 (N_7865,N_2135,N_1462);
nor U7866 (N_7866,N_3385,N_2815);
and U7867 (N_7867,N_2128,N_1462);
nand U7868 (N_7868,N_3550,N_2628);
xnor U7869 (N_7869,N_280,N_1252);
or U7870 (N_7870,N_2876,N_3651);
and U7871 (N_7871,N_266,N_3406);
xnor U7872 (N_7872,N_1237,N_4512);
nand U7873 (N_7873,N_4966,N_3292);
or U7874 (N_7874,N_3783,N_3631);
and U7875 (N_7875,N_2166,N_4384);
xor U7876 (N_7876,N_2071,N_3518);
nor U7877 (N_7877,N_3230,N_4825);
and U7878 (N_7878,N_4011,N_657);
nand U7879 (N_7879,N_4328,N_4782);
and U7880 (N_7880,N_4467,N_4320);
or U7881 (N_7881,N_4413,N_940);
nand U7882 (N_7882,N_3550,N_125);
nor U7883 (N_7883,N_1559,N_2813);
and U7884 (N_7884,N_2143,N_230);
or U7885 (N_7885,N_3370,N_1947);
and U7886 (N_7886,N_2510,N_942);
or U7887 (N_7887,N_4348,N_347);
nand U7888 (N_7888,N_4341,N_4869);
nand U7889 (N_7889,N_647,N_2460);
or U7890 (N_7890,N_1552,N_2513);
xnor U7891 (N_7891,N_4668,N_1701);
or U7892 (N_7892,N_4060,N_4875);
nand U7893 (N_7893,N_3680,N_1912);
or U7894 (N_7894,N_2520,N_3331);
nor U7895 (N_7895,N_4077,N_4219);
and U7896 (N_7896,N_1049,N_2713);
xor U7897 (N_7897,N_753,N_1940);
xor U7898 (N_7898,N_1109,N_1175);
nor U7899 (N_7899,N_2665,N_4825);
nor U7900 (N_7900,N_2307,N_3379);
nand U7901 (N_7901,N_1138,N_1593);
and U7902 (N_7902,N_4737,N_3085);
or U7903 (N_7903,N_4121,N_3077);
and U7904 (N_7904,N_2458,N_1015);
xnor U7905 (N_7905,N_3123,N_1918);
nand U7906 (N_7906,N_2139,N_3954);
nor U7907 (N_7907,N_4369,N_1585);
nand U7908 (N_7908,N_1601,N_2170);
nand U7909 (N_7909,N_1038,N_3356);
nand U7910 (N_7910,N_40,N_2220);
nor U7911 (N_7911,N_2680,N_4730);
xnor U7912 (N_7912,N_4517,N_3085);
or U7913 (N_7913,N_3317,N_4618);
nand U7914 (N_7914,N_1183,N_3386);
nor U7915 (N_7915,N_4469,N_3609);
nand U7916 (N_7916,N_1104,N_3455);
or U7917 (N_7917,N_4959,N_3060);
nor U7918 (N_7918,N_2740,N_3400);
nor U7919 (N_7919,N_2983,N_4811);
nand U7920 (N_7920,N_684,N_4045);
nand U7921 (N_7921,N_2546,N_3834);
and U7922 (N_7922,N_2776,N_2092);
and U7923 (N_7923,N_2807,N_3862);
and U7924 (N_7924,N_2324,N_1834);
or U7925 (N_7925,N_3529,N_975);
and U7926 (N_7926,N_3490,N_3054);
nor U7927 (N_7927,N_2265,N_2517);
xor U7928 (N_7928,N_2210,N_83);
nand U7929 (N_7929,N_3133,N_1010);
nor U7930 (N_7930,N_490,N_3095);
xnor U7931 (N_7931,N_372,N_475);
nand U7932 (N_7932,N_4057,N_2677);
or U7933 (N_7933,N_2053,N_4673);
nor U7934 (N_7934,N_4321,N_3038);
or U7935 (N_7935,N_2944,N_4427);
and U7936 (N_7936,N_332,N_4463);
or U7937 (N_7937,N_3971,N_2576);
xnor U7938 (N_7938,N_1434,N_2381);
nand U7939 (N_7939,N_4583,N_1023);
and U7940 (N_7940,N_4042,N_3044);
nand U7941 (N_7941,N_2178,N_3081);
or U7942 (N_7942,N_967,N_154);
and U7943 (N_7943,N_4175,N_1697);
or U7944 (N_7944,N_2155,N_772);
or U7945 (N_7945,N_3406,N_2348);
nor U7946 (N_7946,N_3945,N_2895);
nand U7947 (N_7947,N_2573,N_3844);
nand U7948 (N_7948,N_4034,N_1141);
or U7949 (N_7949,N_3563,N_3361);
nor U7950 (N_7950,N_772,N_1631);
and U7951 (N_7951,N_3528,N_1674);
nand U7952 (N_7952,N_4180,N_4520);
nor U7953 (N_7953,N_4487,N_1939);
nor U7954 (N_7954,N_4202,N_4799);
xnor U7955 (N_7955,N_4599,N_1375);
or U7956 (N_7956,N_427,N_4042);
xnor U7957 (N_7957,N_3363,N_2613);
xor U7958 (N_7958,N_4126,N_1975);
nor U7959 (N_7959,N_2062,N_4599);
xnor U7960 (N_7960,N_1147,N_934);
and U7961 (N_7961,N_4326,N_3607);
nor U7962 (N_7962,N_4083,N_602);
and U7963 (N_7963,N_4163,N_4183);
or U7964 (N_7964,N_1851,N_1218);
and U7965 (N_7965,N_2314,N_4447);
and U7966 (N_7966,N_1626,N_4519);
and U7967 (N_7967,N_4090,N_247);
xor U7968 (N_7968,N_526,N_2562);
nand U7969 (N_7969,N_2761,N_812);
xor U7970 (N_7970,N_3506,N_3320);
nor U7971 (N_7971,N_4560,N_3601);
and U7972 (N_7972,N_606,N_1149);
nand U7973 (N_7973,N_1591,N_126);
and U7974 (N_7974,N_1977,N_3978);
and U7975 (N_7975,N_3623,N_1916);
and U7976 (N_7976,N_3314,N_700);
nand U7977 (N_7977,N_1695,N_2181);
nor U7978 (N_7978,N_4994,N_2682);
and U7979 (N_7979,N_1460,N_4041);
nand U7980 (N_7980,N_2822,N_4896);
nand U7981 (N_7981,N_29,N_1149);
nor U7982 (N_7982,N_2341,N_2469);
and U7983 (N_7983,N_1933,N_1084);
or U7984 (N_7984,N_2826,N_4941);
nand U7985 (N_7985,N_2544,N_2942);
nand U7986 (N_7986,N_3559,N_2719);
xnor U7987 (N_7987,N_1719,N_3083);
nor U7988 (N_7988,N_292,N_2906);
xnor U7989 (N_7989,N_4223,N_1745);
xnor U7990 (N_7990,N_1586,N_441);
nor U7991 (N_7991,N_4606,N_1456);
xnor U7992 (N_7992,N_514,N_613);
nand U7993 (N_7993,N_2520,N_2939);
xor U7994 (N_7994,N_4883,N_2789);
or U7995 (N_7995,N_257,N_127);
nor U7996 (N_7996,N_2944,N_4064);
or U7997 (N_7997,N_2366,N_1338);
nor U7998 (N_7998,N_3759,N_1377);
nor U7999 (N_7999,N_3852,N_3081);
nand U8000 (N_8000,N_967,N_606);
xnor U8001 (N_8001,N_4898,N_2553);
or U8002 (N_8002,N_2122,N_4506);
and U8003 (N_8003,N_1072,N_4430);
or U8004 (N_8004,N_3429,N_3663);
and U8005 (N_8005,N_3835,N_1267);
nand U8006 (N_8006,N_3826,N_1591);
or U8007 (N_8007,N_479,N_3491);
xor U8008 (N_8008,N_2031,N_2228);
or U8009 (N_8009,N_856,N_2910);
xor U8010 (N_8010,N_4600,N_4882);
and U8011 (N_8011,N_3213,N_1349);
nor U8012 (N_8012,N_2760,N_2685);
and U8013 (N_8013,N_3982,N_92);
xnor U8014 (N_8014,N_2659,N_553);
nand U8015 (N_8015,N_3482,N_425);
xor U8016 (N_8016,N_2289,N_1789);
nor U8017 (N_8017,N_330,N_275);
nor U8018 (N_8018,N_1039,N_1820);
nor U8019 (N_8019,N_3800,N_3130);
xor U8020 (N_8020,N_2722,N_3363);
nand U8021 (N_8021,N_3893,N_824);
xor U8022 (N_8022,N_477,N_547);
nand U8023 (N_8023,N_4665,N_1797);
and U8024 (N_8024,N_185,N_1275);
nor U8025 (N_8025,N_1007,N_4552);
and U8026 (N_8026,N_3740,N_4481);
nand U8027 (N_8027,N_4497,N_677);
nor U8028 (N_8028,N_3480,N_1288);
and U8029 (N_8029,N_4828,N_164);
and U8030 (N_8030,N_3537,N_3944);
nand U8031 (N_8031,N_2662,N_1272);
or U8032 (N_8032,N_3627,N_3985);
or U8033 (N_8033,N_3693,N_3576);
xnor U8034 (N_8034,N_3132,N_1856);
xnor U8035 (N_8035,N_4874,N_2604);
and U8036 (N_8036,N_4372,N_1435);
nand U8037 (N_8037,N_4189,N_891);
and U8038 (N_8038,N_2020,N_3298);
xor U8039 (N_8039,N_2428,N_4715);
and U8040 (N_8040,N_1688,N_1895);
nor U8041 (N_8041,N_2826,N_2259);
nor U8042 (N_8042,N_4201,N_2386);
and U8043 (N_8043,N_1197,N_338);
xor U8044 (N_8044,N_4051,N_311);
xnor U8045 (N_8045,N_4032,N_2324);
nor U8046 (N_8046,N_620,N_3406);
and U8047 (N_8047,N_2954,N_4391);
and U8048 (N_8048,N_2821,N_4886);
or U8049 (N_8049,N_1216,N_786);
nand U8050 (N_8050,N_2856,N_3231);
or U8051 (N_8051,N_1130,N_4631);
nor U8052 (N_8052,N_1860,N_3123);
nand U8053 (N_8053,N_230,N_24);
nor U8054 (N_8054,N_346,N_4331);
nand U8055 (N_8055,N_233,N_4117);
xnor U8056 (N_8056,N_1616,N_4210);
xnor U8057 (N_8057,N_1110,N_3823);
xor U8058 (N_8058,N_2243,N_1955);
xor U8059 (N_8059,N_4217,N_1116);
nand U8060 (N_8060,N_2864,N_1053);
and U8061 (N_8061,N_857,N_4009);
nor U8062 (N_8062,N_2311,N_3289);
nor U8063 (N_8063,N_3562,N_4825);
xnor U8064 (N_8064,N_4319,N_319);
nor U8065 (N_8065,N_539,N_2573);
xnor U8066 (N_8066,N_2078,N_653);
nor U8067 (N_8067,N_1121,N_4558);
or U8068 (N_8068,N_247,N_387);
xor U8069 (N_8069,N_3286,N_3467);
nand U8070 (N_8070,N_204,N_3332);
nor U8071 (N_8071,N_4439,N_1698);
xor U8072 (N_8072,N_2396,N_3499);
and U8073 (N_8073,N_4380,N_2426);
and U8074 (N_8074,N_2777,N_1593);
nor U8075 (N_8075,N_1411,N_1007);
or U8076 (N_8076,N_3071,N_4378);
or U8077 (N_8077,N_4881,N_3693);
or U8078 (N_8078,N_74,N_4297);
nand U8079 (N_8079,N_3999,N_4881);
xnor U8080 (N_8080,N_1548,N_3298);
xor U8081 (N_8081,N_3539,N_1682);
or U8082 (N_8082,N_1415,N_1563);
or U8083 (N_8083,N_2677,N_303);
nor U8084 (N_8084,N_134,N_257);
or U8085 (N_8085,N_4777,N_4885);
nor U8086 (N_8086,N_4517,N_1976);
nand U8087 (N_8087,N_1258,N_601);
nor U8088 (N_8088,N_1106,N_3060);
or U8089 (N_8089,N_2196,N_4897);
and U8090 (N_8090,N_666,N_1878);
xnor U8091 (N_8091,N_1407,N_177);
xor U8092 (N_8092,N_4631,N_4586);
nand U8093 (N_8093,N_2644,N_4839);
or U8094 (N_8094,N_4632,N_2788);
and U8095 (N_8095,N_3958,N_169);
nor U8096 (N_8096,N_291,N_303);
nor U8097 (N_8097,N_1142,N_959);
xor U8098 (N_8098,N_4150,N_1977);
and U8099 (N_8099,N_3937,N_1774);
and U8100 (N_8100,N_2875,N_170);
and U8101 (N_8101,N_4035,N_3539);
and U8102 (N_8102,N_970,N_4964);
xor U8103 (N_8103,N_377,N_179);
nand U8104 (N_8104,N_3946,N_4907);
nor U8105 (N_8105,N_1158,N_4270);
xnor U8106 (N_8106,N_2800,N_1833);
nor U8107 (N_8107,N_84,N_4072);
nor U8108 (N_8108,N_2450,N_3817);
xor U8109 (N_8109,N_2845,N_1592);
nor U8110 (N_8110,N_3135,N_4475);
and U8111 (N_8111,N_2193,N_1176);
nor U8112 (N_8112,N_1904,N_4776);
nor U8113 (N_8113,N_4791,N_4597);
xnor U8114 (N_8114,N_1463,N_220);
nand U8115 (N_8115,N_1050,N_2646);
nor U8116 (N_8116,N_4270,N_133);
nand U8117 (N_8117,N_2794,N_4050);
nor U8118 (N_8118,N_4763,N_4372);
and U8119 (N_8119,N_1324,N_3586);
xnor U8120 (N_8120,N_2332,N_2858);
nor U8121 (N_8121,N_1842,N_2774);
nor U8122 (N_8122,N_3387,N_1516);
nand U8123 (N_8123,N_4770,N_757);
nand U8124 (N_8124,N_1076,N_399);
and U8125 (N_8125,N_3485,N_2981);
xor U8126 (N_8126,N_4336,N_764);
xor U8127 (N_8127,N_4983,N_3681);
nor U8128 (N_8128,N_1021,N_3659);
nand U8129 (N_8129,N_2671,N_2900);
xnor U8130 (N_8130,N_405,N_2782);
nor U8131 (N_8131,N_4889,N_799);
and U8132 (N_8132,N_2899,N_2213);
nand U8133 (N_8133,N_1802,N_4865);
or U8134 (N_8134,N_2409,N_4791);
and U8135 (N_8135,N_1624,N_1737);
nand U8136 (N_8136,N_895,N_1930);
and U8137 (N_8137,N_960,N_2975);
nor U8138 (N_8138,N_4771,N_4395);
or U8139 (N_8139,N_3599,N_3855);
xor U8140 (N_8140,N_3776,N_2861);
nor U8141 (N_8141,N_1875,N_2521);
nor U8142 (N_8142,N_4440,N_1312);
and U8143 (N_8143,N_4504,N_3829);
and U8144 (N_8144,N_518,N_3734);
nand U8145 (N_8145,N_1073,N_1531);
and U8146 (N_8146,N_3502,N_4308);
xnor U8147 (N_8147,N_4272,N_3896);
nand U8148 (N_8148,N_4224,N_2112);
or U8149 (N_8149,N_2849,N_3800);
nand U8150 (N_8150,N_2566,N_3941);
and U8151 (N_8151,N_4415,N_3524);
and U8152 (N_8152,N_4743,N_2077);
and U8153 (N_8153,N_2634,N_4794);
nor U8154 (N_8154,N_1151,N_4712);
xnor U8155 (N_8155,N_2036,N_3200);
nor U8156 (N_8156,N_3826,N_1892);
xor U8157 (N_8157,N_1467,N_3445);
nand U8158 (N_8158,N_4750,N_3787);
nor U8159 (N_8159,N_3922,N_1292);
xor U8160 (N_8160,N_2969,N_4987);
or U8161 (N_8161,N_2986,N_2047);
and U8162 (N_8162,N_4937,N_3898);
nand U8163 (N_8163,N_1762,N_1953);
nor U8164 (N_8164,N_3747,N_2640);
nand U8165 (N_8165,N_2692,N_3001);
nor U8166 (N_8166,N_707,N_480);
or U8167 (N_8167,N_3184,N_4827);
xnor U8168 (N_8168,N_972,N_4044);
or U8169 (N_8169,N_2672,N_4852);
and U8170 (N_8170,N_905,N_1359);
nand U8171 (N_8171,N_3632,N_2247);
xnor U8172 (N_8172,N_4832,N_4582);
nor U8173 (N_8173,N_679,N_776);
xor U8174 (N_8174,N_2992,N_2116);
and U8175 (N_8175,N_951,N_2129);
xor U8176 (N_8176,N_4761,N_162);
nand U8177 (N_8177,N_3091,N_824);
or U8178 (N_8178,N_193,N_2179);
nor U8179 (N_8179,N_3103,N_4675);
and U8180 (N_8180,N_82,N_2503);
nand U8181 (N_8181,N_383,N_803);
xor U8182 (N_8182,N_747,N_4691);
xnor U8183 (N_8183,N_3588,N_3907);
nor U8184 (N_8184,N_4093,N_2090);
and U8185 (N_8185,N_904,N_117);
or U8186 (N_8186,N_4030,N_3493);
nor U8187 (N_8187,N_1312,N_3880);
nand U8188 (N_8188,N_3868,N_4736);
nand U8189 (N_8189,N_3966,N_212);
nor U8190 (N_8190,N_417,N_1890);
xor U8191 (N_8191,N_1529,N_4644);
and U8192 (N_8192,N_4671,N_2554);
or U8193 (N_8193,N_694,N_3463);
or U8194 (N_8194,N_3197,N_3160);
or U8195 (N_8195,N_2079,N_3529);
xnor U8196 (N_8196,N_4090,N_4350);
nand U8197 (N_8197,N_2905,N_2407);
or U8198 (N_8198,N_2452,N_2664);
nor U8199 (N_8199,N_1914,N_70);
nor U8200 (N_8200,N_1281,N_2099);
or U8201 (N_8201,N_1777,N_3478);
xor U8202 (N_8202,N_2722,N_4301);
nor U8203 (N_8203,N_2959,N_3027);
nand U8204 (N_8204,N_3158,N_2322);
nand U8205 (N_8205,N_97,N_257);
nand U8206 (N_8206,N_3103,N_2409);
xnor U8207 (N_8207,N_3242,N_2644);
and U8208 (N_8208,N_4,N_2562);
xnor U8209 (N_8209,N_4676,N_2670);
nor U8210 (N_8210,N_4611,N_3666);
or U8211 (N_8211,N_2968,N_1109);
nand U8212 (N_8212,N_1643,N_3507);
or U8213 (N_8213,N_2578,N_2697);
nand U8214 (N_8214,N_1346,N_1995);
nor U8215 (N_8215,N_1220,N_2496);
and U8216 (N_8216,N_3538,N_1967);
and U8217 (N_8217,N_2438,N_1082);
or U8218 (N_8218,N_2619,N_3515);
or U8219 (N_8219,N_1293,N_4344);
nor U8220 (N_8220,N_3877,N_285);
and U8221 (N_8221,N_104,N_3356);
or U8222 (N_8222,N_3248,N_2648);
and U8223 (N_8223,N_1496,N_4120);
and U8224 (N_8224,N_4686,N_1565);
or U8225 (N_8225,N_4658,N_3927);
nand U8226 (N_8226,N_4770,N_2057);
and U8227 (N_8227,N_595,N_773);
and U8228 (N_8228,N_3874,N_798);
nand U8229 (N_8229,N_200,N_4275);
nor U8230 (N_8230,N_4414,N_1282);
xnor U8231 (N_8231,N_870,N_1872);
and U8232 (N_8232,N_131,N_1119);
xor U8233 (N_8233,N_2842,N_1874);
xor U8234 (N_8234,N_3952,N_3681);
nor U8235 (N_8235,N_4788,N_4598);
and U8236 (N_8236,N_3730,N_4735);
nor U8237 (N_8237,N_1465,N_2223);
and U8238 (N_8238,N_90,N_4655);
nor U8239 (N_8239,N_1002,N_3154);
and U8240 (N_8240,N_3337,N_3584);
nand U8241 (N_8241,N_995,N_1875);
xnor U8242 (N_8242,N_1604,N_3494);
or U8243 (N_8243,N_335,N_3895);
nand U8244 (N_8244,N_1466,N_3590);
and U8245 (N_8245,N_3007,N_3902);
nor U8246 (N_8246,N_3921,N_3966);
or U8247 (N_8247,N_2068,N_2261);
xnor U8248 (N_8248,N_2531,N_3550);
nand U8249 (N_8249,N_4015,N_2365);
nor U8250 (N_8250,N_261,N_1305);
nor U8251 (N_8251,N_3783,N_1309);
xnor U8252 (N_8252,N_1014,N_1335);
and U8253 (N_8253,N_2673,N_1151);
nor U8254 (N_8254,N_3520,N_2147);
or U8255 (N_8255,N_2747,N_2226);
nand U8256 (N_8256,N_527,N_725);
nand U8257 (N_8257,N_1528,N_709);
and U8258 (N_8258,N_2050,N_3952);
nor U8259 (N_8259,N_2962,N_4118);
nand U8260 (N_8260,N_3667,N_1780);
nor U8261 (N_8261,N_4453,N_2253);
nand U8262 (N_8262,N_972,N_729);
and U8263 (N_8263,N_2223,N_74);
nor U8264 (N_8264,N_2377,N_4344);
and U8265 (N_8265,N_870,N_4287);
nand U8266 (N_8266,N_3709,N_2436);
and U8267 (N_8267,N_3774,N_573);
xnor U8268 (N_8268,N_1839,N_1904);
xor U8269 (N_8269,N_1289,N_3609);
nor U8270 (N_8270,N_244,N_1597);
xnor U8271 (N_8271,N_3306,N_4788);
xnor U8272 (N_8272,N_3481,N_63);
or U8273 (N_8273,N_2553,N_3111);
nand U8274 (N_8274,N_794,N_2438);
and U8275 (N_8275,N_984,N_1596);
or U8276 (N_8276,N_2512,N_552);
xnor U8277 (N_8277,N_1178,N_2711);
nand U8278 (N_8278,N_689,N_858);
xor U8279 (N_8279,N_4700,N_4605);
or U8280 (N_8280,N_2159,N_2470);
nor U8281 (N_8281,N_823,N_3883);
nand U8282 (N_8282,N_3657,N_1651);
xor U8283 (N_8283,N_823,N_600);
or U8284 (N_8284,N_4845,N_131);
nand U8285 (N_8285,N_1276,N_817);
xor U8286 (N_8286,N_1017,N_491);
and U8287 (N_8287,N_3786,N_2609);
or U8288 (N_8288,N_4883,N_41);
xnor U8289 (N_8289,N_876,N_1785);
or U8290 (N_8290,N_3761,N_1548);
and U8291 (N_8291,N_209,N_1642);
xor U8292 (N_8292,N_4435,N_4696);
nand U8293 (N_8293,N_898,N_401);
nor U8294 (N_8294,N_4491,N_3870);
nand U8295 (N_8295,N_3983,N_3127);
nor U8296 (N_8296,N_3729,N_2732);
nor U8297 (N_8297,N_1499,N_4625);
nor U8298 (N_8298,N_761,N_3540);
or U8299 (N_8299,N_912,N_2623);
xor U8300 (N_8300,N_1397,N_4875);
or U8301 (N_8301,N_4191,N_2100);
nor U8302 (N_8302,N_3305,N_4947);
or U8303 (N_8303,N_4614,N_3138);
nor U8304 (N_8304,N_1130,N_3471);
or U8305 (N_8305,N_1369,N_2286);
or U8306 (N_8306,N_4846,N_251);
xnor U8307 (N_8307,N_3102,N_1391);
nand U8308 (N_8308,N_3812,N_811);
xnor U8309 (N_8309,N_854,N_549);
nand U8310 (N_8310,N_2715,N_3587);
xnor U8311 (N_8311,N_2361,N_1934);
xor U8312 (N_8312,N_263,N_1742);
xor U8313 (N_8313,N_1417,N_3383);
and U8314 (N_8314,N_2480,N_459);
or U8315 (N_8315,N_246,N_4197);
nand U8316 (N_8316,N_3066,N_2229);
and U8317 (N_8317,N_3514,N_557);
and U8318 (N_8318,N_1072,N_2018);
and U8319 (N_8319,N_4982,N_3700);
or U8320 (N_8320,N_1261,N_1405);
and U8321 (N_8321,N_723,N_3092);
and U8322 (N_8322,N_2883,N_933);
and U8323 (N_8323,N_2547,N_2327);
nand U8324 (N_8324,N_88,N_753);
nor U8325 (N_8325,N_77,N_4046);
and U8326 (N_8326,N_2342,N_2485);
and U8327 (N_8327,N_3388,N_1881);
and U8328 (N_8328,N_854,N_1374);
nor U8329 (N_8329,N_1334,N_2511);
nand U8330 (N_8330,N_4083,N_3111);
nand U8331 (N_8331,N_3490,N_3815);
nand U8332 (N_8332,N_3355,N_65);
nand U8333 (N_8333,N_4737,N_217);
or U8334 (N_8334,N_1884,N_4997);
nor U8335 (N_8335,N_3188,N_773);
nand U8336 (N_8336,N_4418,N_1663);
nor U8337 (N_8337,N_439,N_4988);
xor U8338 (N_8338,N_2192,N_4855);
nor U8339 (N_8339,N_441,N_1115);
and U8340 (N_8340,N_936,N_1994);
nor U8341 (N_8341,N_4427,N_3360);
nand U8342 (N_8342,N_1223,N_2088);
or U8343 (N_8343,N_244,N_4864);
xor U8344 (N_8344,N_2750,N_1503);
or U8345 (N_8345,N_3138,N_1646);
or U8346 (N_8346,N_3940,N_1502);
nor U8347 (N_8347,N_29,N_4033);
xor U8348 (N_8348,N_1599,N_2222);
nand U8349 (N_8349,N_2148,N_3777);
xor U8350 (N_8350,N_383,N_2300);
nand U8351 (N_8351,N_3470,N_3266);
or U8352 (N_8352,N_4682,N_3468);
nand U8353 (N_8353,N_941,N_1501);
nand U8354 (N_8354,N_2565,N_1614);
and U8355 (N_8355,N_3182,N_3482);
and U8356 (N_8356,N_496,N_1249);
nand U8357 (N_8357,N_3360,N_2455);
or U8358 (N_8358,N_2627,N_3813);
xor U8359 (N_8359,N_3816,N_2252);
nor U8360 (N_8360,N_3510,N_2745);
nor U8361 (N_8361,N_3197,N_2987);
nor U8362 (N_8362,N_2461,N_2808);
and U8363 (N_8363,N_1335,N_2607);
and U8364 (N_8364,N_1211,N_1080);
nand U8365 (N_8365,N_3124,N_4726);
and U8366 (N_8366,N_64,N_2617);
nor U8367 (N_8367,N_3010,N_2783);
xnor U8368 (N_8368,N_3501,N_846);
nand U8369 (N_8369,N_2372,N_3798);
nor U8370 (N_8370,N_3403,N_3800);
xor U8371 (N_8371,N_3489,N_4628);
or U8372 (N_8372,N_2465,N_1768);
and U8373 (N_8373,N_2285,N_4547);
or U8374 (N_8374,N_4303,N_4275);
nand U8375 (N_8375,N_2614,N_3694);
nand U8376 (N_8376,N_3967,N_4064);
or U8377 (N_8377,N_2527,N_2220);
xor U8378 (N_8378,N_114,N_4791);
xnor U8379 (N_8379,N_1293,N_4408);
or U8380 (N_8380,N_714,N_642);
nor U8381 (N_8381,N_1123,N_4406);
or U8382 (N_8382,N_2661,N_4009);
and U8383 (N_8383,N_1582,N_201);
or U8384 (N_8384,N_4336,N_2925);
nor U8385 (N_8385,N_4071,N_1619);
or U8386 (N_8386,N_972,N_2185);
and U8387 (N_8387,N_354,N_4219);
xor U8388 (N_8388,N_3811,N_1271);
or U8389 (N_8389,N_4463,N_2470);
nor U8390 (N_8390,N_813,N_2686);
nand U8391 (N_8391,N_860,N_2333);
or U8392 (N_8392,N_2432,N_4624);
nor U8393 (N_8393,N_633,N_4488);
or U8394 (N_8394,N_2922,N_4430);
nor U8395 (N_8395,N_1824,N_64);
xnor U8396 (N_8396,N_908,N_323);
nor U8397 (N_8397,N_492,N_18);
xnor U8398 (N_8398,N_428,N_4988);
xor U8399 (N_8399,N_2153,N_1330);
or U8400 (N_8400,N_1911,N_1535);
and U8401 (N_8401,N_3729,N_4569);
nor U8402 (N_8402,N_2174,N_1786);
nand U8403 (N_8403,N_3132,N_4252);
nor U8404 (N_8404,N_3482,N_1282);
nor U8405 (N_8405,N_2985,N_3395);
and U8406 (N_8406,N_2511,N_1095);
and U8407 (N_8407,N_1287,N_4866);
and U8408 (N_8408,N_1482,N_2574);
nor U8409 (N_8409,N_2299,N_1422);
nor U8410 (N_8410,N_1616,N_1266);
xor U8411 (N_8411,N_4274,N_4968);
and U8412 (N_8412,N_3864,N_3424);
and U8413 (N_8413,N_2445,N_3540);
nor U8414 (N_8414,N_1415,N_2437);
xnor U8415 (N_8415,N_994,N_1273);
and U8416 (N_8416,N_2769,N_2130);
and U8417 (N_8417,N_569,N_1587);
and U8418 (N_8418,N_1967,N_785);
and U8419 (N_8419,N_2522,N_1349);
and U8420 (N_8420,N_4298,N_1040);
and U8421 (N_8421,N_2635,N_4436);
xnor U8422 (N_8422,N_2591,N_2687);
xor U8423 (N_8423,N_1668,N_3816);
or U8424 (N_8424,N_3027,N_4526);
xor U8425 (N_8425,N_2909,N_1872);
xor U8426 (N_8426,N_4133,N_1536);
nand U8427 (N_8427,N_4786,N_1426);
and U8428 (N_8428,N_444,N_3533);
or U8429 (N_8429,N_2787,N_1043);
or U8430 (N_8430,N_4077,N_100);
or U8431 (N_8431,N_2295,N_399);
nand U8432 (N_8432,N_1783,N_1302);
nand U8433 (N_8433,N_1442,N_1767);
nand U8434 (N_8434,N_3231,N_2361);
xor U8435 (N_8435,N_786,N_1769);
or U8436 (N_8436,N_2228,N_1693);
xor U8437 (N_8437,N_769,N_270);
nor U8438 (N_8438,N_3248,N_1390);
xnor U8439 (N_8439,N_605,N_2665);
nand U8440 (N_8440,N_2026,N_3787);
or U8441 (N_8441,N_4926,N_1859);
and U8442 (N_8442,N_1229,N_1238);
xor U8443 (N_8443,N_4000,N_4680);
or U8444 (N_8444,N_2348,N_571);
nor U8445 (N_8445,N_3066,N_4109);
or U8446 (N_8446,N_4146,N_1793);
nand U8447 (N_8447,N_1597,N_4312);
nand U8448 (N_8448,N_2240,N_1207);
and U8449 (N_8449,N_4493,N_3995);
nor U8450 (N_8450,N_4218,N_3731);
xnor U8451 (N_8451,N_2058,N_3929);
xor U8452 (N_8452,N_1951,N_3911);
nor U8453 (N_8453,N_3258,N_1703);
or U8454 (N_8454,N_4580,N_4338);
nor U8455 (N_8455,N_3033,N_4283);
xor U8456 (N_8456,N_3872,N_63);
and U8457 (N_8457,N_3970,N_2984);
nor U8458 (N_8458,N_522,N_2630);
nand U8459 (N_8459,N_4909,N_2290);
nor U8460 (N_8460,N_4674,N_3729);
nor U8461 (N_8461,N_2066,N_3678);
nor U8462 (N_8462,N_428,N_4761);
and U8463 (N_8463,N_1196,N_3650);
or U8464 (N_8464,N_1605,N_1599);
or U8465 (N_8465,N_877,N_4901);
or U8466 (N_8466,N_1852,N_2297);
and U8467 (N_8467,N_4993,N_153);
and U8468 (N_8468,N_247,N_4179);
nor U8469 (N_8469,N_205,N_4581);
xor U8470 (N_8470,N_2362,N_556);
or U8471 (N_8471,N_1099,N_848);
nand U8472 (N_8472,N_3989,N_1926);
or U8473 (N_8473,N_1316,N_2295);
and U8474 (N_8474,N_1934,N_3748);
or U8475 (N_8475,N_390,N_4690);
nor U8476 (N_8476,N_2795,N_1308);
and U8477 (N_8477,N_4467,N_1560);
nor U8478 (N_8478,N_1485,N_2277);
nor U8479 (N_8479,N_3327,N_2262);
xnor U8480 (N_8480,N_1097,N_3397);
or U8481 (N_8481,N_3263,N_4467);
or U8482 (N_8482,N_3819,N_922);
xnor U8483 (N_8483,N_1343,N_1788);
and U8484 (N_8484,N_1232,N_246);
nor U8485 (N_8485,N_2093,N_3535);
nor U8486 (N_8486,N_4469,N_4710);
xor U8487 (N_8487,N_1740,N_2065);
xnor U8488 (N_8488,N_1322,N_2666);
xor U8489 (N_8489,N_1663,N_2803);
and U8490 (N_8490,N_1337,N_3588);
or U8491 (N_8491,N_1761,N_1931);
xor U8492 (N_8492,N_2572,N_3181);
and U8493 (N_8493,N_4453,N_2004);
or U8494 (N_8494,N_23,N_1270);
nand U8495 (N_8495,N_4405,N_278);
nor U8496 (N_8496,N_832,N_3956);
nand U8497 (N_8497,N_2966,N_4418);
nor U8498 (N_8498,N_3292,N_474);
xnor U8499 (N_8499,N_1502,N_2699);
nand U8500 (N_8500,N_2973,N_3668);
and U8501 (N_8501,N_2533,N_669);
nand U8502 (N_8502,N_81,N_1087);
or U8503 (N_8503,N_751,N_929);
nand U8504 (N_8504,N_492,N_1260);
nor U8505 (N_8505,N_323,N_1875);
or U8506 (N_8506,N_4783,N_1552);
nor U8507 (N_8507,N_1369,N_257);
nand U8508 (N_8508,N_956,N_3606);
and U8509 (N_8509,N_42,N_2867);
xor U8510 (N_8510,N_3217,N_4396);
or U8511 (N_8511,N_4807,N_2256);
nor U8512 (N_8512,N_2296,N_4968);
or U8513 (N_8513,N_2633,N_4854);
xnor U8514 (N_8514,N_937,N_1377);
or U8515 (N_8515,N_1794,N_2018);
and U8516 (N_8516,N_1514,N_3281);
nand U8517 (N_8517,N_3540,N_2370);
nand U8518 (N_8518,N_2754,N_4145);
and U8519 (N_8519,N_2750,N_4408);
xor U8520 (N_8520,N_1920,N_1024);
nand U8521 (N_8521,N_1266,N_3295);
nor U8522 (N_8522,N_2150,N_3433);
nor U8523 (N_8523,N_4573,N_3642);
nand U8524 (N_8524,N_71,N_2120);
and U8525 (N_8525,N_1611,N_770);
and U8526 (N_8526,N_1935,N_2938);
or U8527 (N_8527,N_4243,N_213);
and U8528 (N_8528,N_2694,N_3682);
xor U8529 (N_8529,N_4491,N_4635);
and U8530 (N_8530,N_1371,N_1596);
or U8531 (N_8531,N_4027,N_2909);
nand U8532 (N_8532,N_1851,N_3354);
or U8533 (N_8533,N_2411,N_2413);
nand U8534 (N_8534,N_1115,N_3916);
xor U8535 (N_8535,N_1430,N_3505);
and U8536 (N_8536,N_1264,N_1985);
and U8537 (N_8537,N_2836,N_142);
and U8538 (N_8538,N_3202,N_3820);
and U8539 (N_8539,N_1559,N_628);
nand U8540 (N_8540,N_3862,N_4194);
xnor U8541 (N_8541,N_578,N_2740);
nand U8542 (N_8542,N_524,N_1858);
nand U8543 (N_8543,N_4759,N_4344);
nand U8544 (N_8544,N_2436,N_2140);
and U8545 (N_8545,N_525,N_2747);
xor U8546 (N_8546,N_4251,N_2216);
nor U8547 (N_8547,N_2221,N_1762);
xnor U8548 (N_8548,N_868,N_1677);
nor U8549 (N_8549,N_4144,N_1057);
nand U8550 (N_8550,N_4674,N_1991);
nand U8551 (N_8551,N_712,N_4826);
and U8552 (N_8552,N_4181,N_2733);
nand U8553 (N_8553,N_2686,N_1394);
and U8554 (N_8554,N_1216,N_4410);
nor U8555 (N_8555,N_2179,N_4801);
xnor U8556 (N_8556,N_2932,N_2443);
or U8557 (N_8557,N_2303,N_3446);
nor U8558 (N_8558,N_153,N_2027);
xnor U8559 (N_8559,N_1104,N_1919);
nand U8560 (N_8560,N_4789,N_1265);
or U8561 (N_8561,N_4532,N_1625);
and U8562 (N_8562,N_1986,N_1059);
or U8563 (N_8563,N_580,N_1028);
or U8564 (N_8564,N_4661,N_2330);
nor U8565 (N_8565,N_3450,N_4936);
xor U8566 (N_8566,N_4417,N_373);
and U8567 (N_8567,N_492,N_2698);
nor U8568 (N_8568,N_1904,N_1851);
and U8569 (N_8569,N_4023,N_2104);
xor U8570 (N_8570,N_2251,N_826);
nand U8571 (N_8571,N_1198,N_736);
nor U8572 (N_8572,N_44,N_1782);
xnor U8573 (N_8573,N_3487,N_121);
and U8574 (N_8574,N_169,N_640);
and U8575 (N_8575,N_1188,N_1275);
nor U8576 (N_8576,N_3390,N_4977);
nand U8577 (N_8577,N_1826,N_1401);
nand U8578 (N_8578,N_1796,N_103);
or U8579 (N_8579,N_1883,N_4245);
xor U8580 (N_8580,N_26,N_2764);
nand U8581 (N_8581,N_317,N_4582);
nor U8582 (N_8582,N_4484,N_2942);
and U8583 (N_8583,N_4891,N_428);
and U8584 (N_8584,N_4190,N_2704);
xnor U8585 (N_8585,N_2815,N_1353);
and U8586 (N_8586,N_3323,N_3037);
nand U8587 (N_8587,N_1207,N_376);
or U8588 (N_8588,N_1254,N_2277);
or U8589 (N_8589,N_1250,N_3277);
xor U8590 (N_8590,N_332,N_2912);
nand U8591 (N_8591,N_2841,N_2121);
or U8592 (N_8592,N_4628,N_2400);
nor U8593 (N_8593,N_1368,N_4570);
or U8594 (N_8594,N_3247,N_533);
and U8595 (N_8595,N_636,N_3593);
and U8596 (N_8596,N_3244,N_3702);
and U8597 (N_8597,N_3008,N_3427);
and U8598 (N_8598,N_338,N_3393);
xnor U8599 (N_8599,N_1231,N_3208);
or U8600 (N_8600,N_3234,N_893);
xor U8601 (N_8601,N_886,N_3469);
xnor U8602 (N_8602,N_4365,N_4686);
nand U8603 (N_8603,N_3931,N_3054);
nand U8604 (N_8604,N_3712,N_3003);
nand U8605 (N_8605,N_4920,N_3670);
xnor U8606 (N_8606,N_3765,N_887);
nand U8607 (N_8607,N_4668,N_2096);
nor U8608 (N_8608,N_4835,N_3693);
nand U8609 (N_8609,N_797,N_1024);
or U8610 (N_8610,N_844,N_336);
xnor U8611 (N_8611,N_4740,N_1257);
and U8612 (N_8612,N_362,N_4287);
nor U8613 (N_8613,N_2346,N_2306);
nand U8614 (N_8614,N_101,N_1876);
xor U8615 (N_8615,N_4550,N_596);
xor U8616 (N_8616,N_1492,N_4666);
or U8617 (N_8617,N_4488,N_4287);
or U8618 (N_8618,N_520,N_2229);
and U8619 (N_8619,N_2689,N_505);
xnor U8620 (N_8620,N_4283,N_4499);
nor U8621 (N_8621,N_677,N_818);
nor U8622 (N_8622,N_3772,N_3135);
xnor U8623 (N_8623,N_3903,N_1700);
nor U8624 (N_8624,N_4755,N_1310);
or U8625 (N_8625,N_4763,N_3224);
xnor U8626 (N_8626,N_552,N_2346);
nand U8627 (N_8627,N_4527,N_2954);
nand U8628 (N_8628,N_2503,N_1812);
or U8629 (N_8629,N_1063,N_3747);
and U8630 (N_8630,N_2450,N_4091);
or U8631 (N_8631,N_4334,N_4520);
nand U8632 (N_8632,N_3807,N_1395);
xor U8633 (N_8633,N_2018,N_1408);
nor U8634 (N_8634,N_4184,N_2638);
nor U8635 (N_8635,N_1955,N_2072);
or U8636 (N_8636,N_4065,N_3991);
and U8637 (N_8637,N_970,N_4716);
and U8638 (N_8638,N_1780,N_738);
xor U8639 (N_8639,N_438,N_1195);
or U8640 (N_8640,N_611,N_2557);
xnor U8641 (N_8641,N_208,N_4999);
xnor U8642 (N_8642,N_3325,N_1239);
xor U8643 (N_8643,N_1178,N_4269);
and U8644 (N_8644,N_3268,N_2679);
xor U8645 (N_8645,N_535,N_2228);
nor U8646 (N_8646,N_3255,N_2083);
xor U8647 (N_8647,N_4005,N_943);
or U8648 (N_8648,N_729,N_3380);
nand U8649 (N_8649,N_621,N_1223);
xnor U8650 (N_8650,N_308,N_4507);
and U8651 (N_8651,N_3388,N_3552);
nor U8652 (N_8652,N_2985,N_3748);
and U8653 (N_8653,N_3684,N_3871);
nor U8654 (N_8654,N_2703,N_2531);
xor U8655 (N_8655,N_855,N_2474);
nor U8656 (N_8656,N_600,N_261);
nor U8657 (N_8657,N_3040,N_459);
xor U8658 (N_8658,N_3317,N_3798);
nand U8659 (N_8659,N_3960,N_4125);
or U8660 (N_8660,N_4099,N_4044);
nand U8661 (N_8661,N_3857,N_3496);
nand U8662 (N_8662,N_452,N_1786);
xnor U8663 (N_8663,N_22,N_786);
nand U8664 (N_8664,N_313,N_2620);
or U8665 (N_8665,N_2659,N_1654);
and U8666 (N_8666,N_2797,N_691);
nand U8667 (N_8667,N_2572,N_1034);
nor U8668 (N_8668,N_4884,N_106);
nand U8669 (N_8669,N_1399,N_3405);
xnor U8670 (N_8670,N_853,N_2055);
and U8671 (N_8671,N_676,N_1600);
or U8672 (N_8672,N_1145,N_211);
or U8673 (N_8673,N_1215,N_1702);
and U8674 (N_8674,N_245,N_3302);
and U8675 (N_8675,N_4040,N_3713);
nor U8676 (N_8676,N_4355,N_1135);
nor U8677 (N_8677,N_3601,N_2883);
nand U8678 (N_8678,N_1784,N_1256);
and U8679 (N_8679,N_281,N_420);
nand U8680 (N_8680,N_4403,N_2126);
nand U8681 (N_8681,N_82,N_2436);
nand U8682 (N_8682,N_3677,N_998);
xnor U8683 (N_8683,N_1333,N_3630);
nand U8684 (N_8684,N_3616,N_743);
nor U8685 (N_8685,N_3804,N_931);
xnor U8686 (N_8686,N_3735,N_2648);
nor U8687 (N_8687,N_3543,N_1920);
xor U8688 (N_8688,N_4562,N_2061);
and U8689 (N_8689,N_1005,N_4875);
or U8690 (N_8690,N_738,N_25);
nor U8691 (N_8691,N_3214,N_2062);
and U8692 (N_8692,N_4079,N_1194);
and U8693 (N_8693,N_4754,N_3805);
nor U8694 (N_8694,N_4123,N_1082);
nand U8695 (N_8695,N_1489,N_4485);
and U8696 (N_8696,N_2216,N_3593);
nor U8697 (N_8697,N_2858,N_2821);
xor U8698 (N_8698,N_1054,N_1575);
and U8699 (N_8699,N_2690,N_2287);
xor U8700 (N_8700,N_966,N_2109);
and U8701 (N_8701,N_723,N_1704);
nand U8702 (N_8702,N_1210,N_128);
nand U8703 (N_8703,N_3112,N_251);
nor U8704 (N_8704,N_113,N_2094);
nor U8705 (N_8705,N_709,N_3825);
nand U8706 (N_8706,N_4121,N_2714);
nor U8707 (N_8707,N_1160,N_3141);
nand U8708 (N_8708,N_3366,N_1150);
and U8709 (N_8709,N_2439,N_3294);
xor U8710 (N_8710,N_1610,N_686);
nor U8711 (N_8711,N_3955,N_1048);
nor U8712 (N_8712,N_4228,N_2023);
nand U8713 (N_8713,N_3521,N_3274);
or U8714 (N_8714,N_4102,N_356);
or U8715 (N_8715,N_2767,N_3958);
nand U8716 (N_8716,N_3581,N_1701);
nor U8717 (N_8717,N_3348,N_3129);
nor U8718 (N_8718,N_4256,N_2929);
or U8719 (N_8719,N_1753,N_2471);
nand U8720 (N_8720,N_1343,N_4915);
xor U8721 (N_8721,N_2059,N_1302);
or U8722 (N_8722,N_1705,N_1250);
xnor U8723 (N_8723,N_1176,N_4489);
or U8724 (N_8724,N_3077,N_2125);
and U8725 (N_8725,N_1188,N_628);
nor U8726 (N_8726,N_4576,N_977);
nand U8727 (N_8727,N_4476,N_4786);
or U8728 (N_8728,N_3972,N_2595);
nand U8729 (N_8729,N_4041,N_2339);
nand U8730 (N_8730,N_4601,N_3808);
or U8731 (N_8731,N_4525,N_4349);
nor U8732 (N_8732,N_2800,N_654);
and U8733 (N_8733,N_421,N_4442);
or U8734 (N_8734,N_2167,N_2983);
xor U8735 (N_8735,N_2070,N_4342);
or U8736 (N_8736,N_3667,N_1664);
nand U8737 (N_8737,N_1687,N_1605);
nor U8738 (N_8738,N_3280,N_1714);
or U8739 (N_8739,N_1838,N_3052);
and U8740 (N_8740,N_929,N_1433);
nor U8741 (N_8741,N_4531,N_1899);
or U8742 (N_8742,N_4754,N_1769);
and U8743 (N_8743,N_1619,N_1730);
xor U8744 (N_8744,N_1142,N_2240);
or U8745 (N_8745,N_1038,N_1084);
xnor U8746 (N_8746,N_3700,N_3434);
nand U8747 (N_8747,N_399,N_26);
and U8748 (N_8748,N_3716,N_3565);
nand U8749 (N_8749,N_2739,N_2067);
and U8750 (N_8750,N_1978,N_3957);
nand U8751 (N_8751,N_463,N_762);
xnor U8752 (N_8752,N_2701,N_3830);
nand U8753 (N_8753,N_907,N_2195);
or U8754 (N_8754,N_4994,N_339);
nand U8755 (N_8755,N_3529,N_2962);
nand U8756 (N_8756,N_4557,N_1563);
xnor U8757 (N_8757,N_1876,N_710);
nor U8758 (N_8758,N_4245,N_4457);
nor U8759 (N_8759,N_3987,N_3796);
and U8760 (N_8760,N_1041,N_2043);
and U8761 (N_8761,N_1158,N_4226);
nand U8762 (N_8762,N_4023,N_3556);
xor U8763 (N_8763,N_1226,N_3245);
or U8764 (N_8764,N_4232,N_2614);
or U8765 (N_8765,N_246,N_463);
or U8766 (N_8766,N_1595,N_4222);
xnor U8767 (N_8767,N_3900,N_259);
xnor U8768 (N_8768,N_1507,N_1983);
or U8769 (N_8769,N_2078,N_690);
xor U8770 (N_8770,N_3708,N_3182);
xnor U8771 (N_8771,N_3660,N_4379);
nor U8772 (N_8772,N_3467,N_2260);
nor U8773 (N_8773,N_792,N_3862);
nor U8774 (N_8774,N_3485,N_862);
xnor U8775 (N_8775,N_3481,N_1916);
nor U8776 (N_8776,N_4034,N_3629);
or U8777 (N_8777,N_2045,N_4119);
or U8778 (N_8778,N_2028,N_1685);
xnor U8779 (N_8779,N_3674,N_1805);
and U8780 (N_8780,N_1160,N_338);
nand U8781 (N_8781,N_3215,N_1295);
and U8782 (N_8782,N_973,N_636);
and U8783 (N_8783,N_3738,N_4724);
and U8784 (N_8784,N_1823,N_2044);
xnor U8785 (N_8785,N_716,N_3944);
or U8786 (N_8786,N_1357,N_1673);
and U8787 (N_8787,N_2206,N_622);
xnor U8788 (N_8788,N_718,N_2101);
or U8789 (N_8789,N_1517,N_4473);
or U8790 (N_8790,N_3813,N_2164);
nand U8791 (N_8791,N_623,N_3159);
nand U8792 (N_8792,N_2998,N_2104);
xor U8793 (N_8793,N_1715,N_4615);
or U8794 (N_8794,N_1949,N_928);
and U8795 (N_8795,N_632,N_764);
and U8796 (N_8796,N_2205,N_4147);
or U8797 (N_8797,N_3250,N_3670);
or U8798 (N_8798,N_2924,N_3312);
nand U8799 (N_8799,N_1905,N_3355);
or U8800 (N_8800,N_3291,N_3276);
nor U8801 (N_8801,N_4184,N_4965);
and U8802 (N_8802,N_4580,N_3615);
xor U8803 (N_8803,N_1236,N_11);
or U8804 (N_8804,N_731,N_4991);
nor U8805 (N_8805,N_4262,N_1533);
and U8806 (N_8806,N_2938,N_177);
nand U8807 (N_8807,N_13,N_3);
nor U8808 (N_8808,N_499,N_3694);
and U8809 (N_8809,N_2344,N_4701);
nand U8810 (N_8810,N_94,N_257);
xor U8811 (N_8811,N_3854,N_3194);
and U8812 (N_8812,N_2480,N_3056);
nand U8813 (N_8813,N_4018,N_4752);
nor U8814 (N_8814,N_1861,N_3123);
and U8815 (N_8815,N_3965,N_2627);
nand U8816 (N_8816,N_3611,N_1612);
xnor U8817 (N_8817,N_2303,N_4253);
xnor U8818 (N_8818,N_2004,N_2979);
nor U8819 (N_8819,N_4605,N_2327);
or U8820 (N_8820,N_1844,N_4411);
and U8821 (N_8821,N_228,N_1477);
or U8822 (N_8822,N_2706,N_1360);
xor U8823 (N_8823,N_1296,N_652);
and U8824 (N_8824,N_872,N_344);
and U8825 (N_8825,N_3636,N_3526);
xnor U8826 (N_8826,N_1518,N_1580);
nor U8827 (N_8827,N_4396,N_2207);
nor U8828 (N_8828,N_3667,N_1386);
nand U8829 (N_8829,N_1576,N_987);
nand U8830 (N_8830,N_112,N_241);
nand U8831 (N_8831,N_4451,N_4188);
xnor U8832 (N_8832,N_1246,N_3888);
and U8833 (N_8833,N_4398,N_3427);
nand U8834 (N_8834,N_1881,N_886);
and U8835 (N_8835,N_2410,N_910);
xor U8836 (N_8836,N_4983,N_4220);
or U8837 (N_8837,N_1511,N_1138);
nor U8838 (N_8838,N_800,N_2468);
or U8839 (N_8839,N_2452,N_2534);
xor U8840 (N_8840,N_2995,N_2556);
nor U8841 (N_8841,N_885,N_362);
or U8842 (N_8842,N_4663,N_532);
and U8843 (N_8843,N_4308,N_1890);
and U8844 (N_8844,N_829,N_1956);
xnor U8845 (N_8845,N_4508,N_3963);
xor U8846 (N_8846,N_2551,N_2625);
or U8847 (N_8847,N_2830,N_2597);
and U8848 (N_8848,N_1142,N_2793);
and U8849 (N_8849,N_3245,N_49);
and U8850 (N_8850,N_4658,N_1606);
nor U8851 (N_8851,N_4674,N_831);
and U8852 (N_8852,N_1360,N_4024);
and U8853 (N_8853,N_3294,N_4029);
nand U8854 (N_8854,N_4681,N_656);
xnor U8855 (N_8855,N_40,N_4618);
or U8856 (N_8856,N_126,N_3576);
xor U8857 (N_8857,N_912,N_2935);
nand U8858 (N_8858,N_2032,N_2984);
or U8859 (N_8859,N_4289,N_365);
xor U8860 (N_8860,N_849,N_2210);
nor U8861 (N_8861,N_2120,N_2709);
nor U8862 (N_8862,N_1765,N_2046);
nor U8863 (N_8863,N_3075,N_3539);
and U8864 (N_8864,N_1978,N_3352);
or U8865 (N_8865,N_2537,N_1179);
and U8866 (N_8866,N_3308,N_2841);
and U8867 (N_8867,N_1794,N_4953);
nand U8868 (N_8868,N_1380,N_260);
nand U8869 (N_8869,N_2124,N_3567);
or U8870 (N_8870,N_3115,N_3740);
nor U8871 (N_8871,N_3528,N_2622);
nor U8872 (N_8872,N_1855,N_2537);
and U8873 (N_8873,N_1360,N_501);
and U8874 (N_8874,N_1459,N_3278);
nor U8875 (N_8875,N_3695,N_2236);
nand U8876 (N_8876,N_4475,N_2280);
xnor U8877 (N_8877,N_33,N_3061);
or U8878 (N_8878,N_2164,N_3267);
nand U8879 (N_8879,N_3342,N_3651);
nor U8880 (N_8880,N_4401,N_938);
nand U8881 (N_8881,N_4463,N_4538);
xnor U8882 (N_8882,N_392,N_3703);
and U8883 (N_8883,N_1333,N_4587);
and U8884 (N_8884,N_2092,N_4744);
nor U8885 (N_8885,N_4137,N_4695);
nand U8886 (N_8886,N_173,N_3682);
and U8887 (N_8887,N_1970,N_795);
nor U8888 (N_8888,N_1697,N_2927);
and U8889 (N_8889,N_3204,N_3709);
nor U8890 (N_8890,N_102,N_299);
and U8891 (N_8891,N_3390,N_411);
xnor U8892 (N_8892,N_207,N_4260);
or U8893 (N_8893,N_3301,N_2798);
nor U8894 (N_8894,N_1419,N_2700);
xor U8895 (N_8895,N_4213,N_3158);
nor U8896 (N_8896,N_4030,N_4923);
nand U8897 (N_8897,N_3880,N_4107);
nand U8898 (N_8898,N_1374,N_2460);
nor U8899 (N_8899,N_849,N_4730);
xor U8900 (N_8900,N_4413,N_1010);
nand U8901 (N_8901,N_2498,N_64);
or U8902 (N_8902,N_580,N_2049);
or U8903 (N_8903,N_3287,N_4687);
xnor U8904 (N_8904,N_3335,N_1915);
or U8905 (N_8905,N_3638,N_3319);
and U8906 (N_8906,N_4875,N_533);
nand U8907 (N_8907,N_3596,N_267);
xor U8908 (N_8908,N_35,N_359);
nor U8909 (N_8909,N_1957,N_3798);
or U8910 (N_8910,N_1168,N_2090);
and U8911 (N_8911,N_4633,N_3834);
nor U8912 (N_8912,N_4026,N_177);
xor U8913 (N_8913,N_4642,N_3362);
xnor U8914 (N_8914,N_3556,N_4287);
nand U8915 (N_8915,N_876,N_1036);
or U8916 (N_8916,N_1318,N_1402);
or U8917 (N_8917,N_3465,N_2852);
nand U8918 (N_8918,N_4528,N_4131);
nor U8919 (N_8919,N_2515,N_2541);
and U8920 (N_8920,N_1737,N_1107);
xnor U8921 (N_8921,N_3960,N_4607);
or U8922 (N_8922,N_4590,N_4220);
and U8923 (N_8923,N_4846,N_2497);
nor U8924 (N_8924,N_24,N_4626);
nor U8925 (N_8925,N_959,N_840);
nand U8926 (N_8926,N_2476,N_3844);
and U8927 (N_8927,N_3809,N_1808);
nand U8928 (N_8928,N_535,N_2177);
nand U8929 (N_8929,N_248,N_3391);
nor U8930 (N_8930,N_679,N_3309);
or U8931 (N_8931,N_2685,N_1021);
nor U8932 (N_8932,N_2932,N_2439);
or U8933 (N_8933,N_1432,N_4088);
and U8934 (N_8934,N_3632,N_4321);
nand U8935 (N_8935,N_2888,N_1627);
and U8936 (N_8936,N_3106,N_3231);
nor U8937 (N_8937,N_3006,N_1035);
or U8938 (N_8938,N_766,N_3291);
and U8939 (N_8939,N_3067,N_3598);
nand U8940 (N_8940,N_976,N_2957);
nor U8941 (N_8941,N_937,N_1993);
or U8942 (N_8942,N_866,N_4878);
nor U8943 (N_8943,N_802,N_278);
and U8944 (N_8944,N_4790,N_4025);
and U8945 (N_8945,N_4283,N_2918);
xnor U8946 (N_8946,N_325,N_2102);
nand U8947 (N_8947,N_4880,N_1767);
and U8948 (N_8948,N_1351,N_3431);
xnor U8949 (N_8949,N_1366,N_4023);
xor U8950 (N_8950,N_1692,N_529);
or U8951 (N_8951,N_740,N_3417);
nor U8952 (N_8952,N_1097,N_221);
and U8953 (N_8953,N_1121,N_1504);
xnor U8954 (N_8954,N_1448,N_3747);
nand U8955 (N_8955,N_4207,N_3386);
and U8956 (N_8956,N_3773,N_2931);
or U8957 (N_8957,N_3741,N_1598);
nand U8958 (N_8958,N_2478,N_109);
and U8959 (N_8959,N_1163,N_2317);
or U8960 (N_8960,N_2720,N_3291);
nand U8961 (N_8961,N_4664,N_2717);
and U8962 (N_8962,N_1962,N_2380);
and U8963 (N_8963,N_2892,N_2879);
nand U8964 (N_8964,N_2299,N_4977);
and U8965 (N_8965,N_1799,N_900);
or U8966 (N_8966,N_210,N_2829);
and U8967 (N_8967,N_4310,N_2299);
and U8968 (N_8968,N_327,N_674);
nor U8969 (N_8969,N_3334,N_541);
nand U8970 (N_8970,N_128,N_1816);
xnor U8971 (N_8971,N_1178,N_410);
or U8972 (N_8972,N_730,N_1599);
xor U8973 (N_8973,N_4802,N_3894);
xor U8974 (N_8974,N_2737,N_1361);
nand U8975 (N_8975,N_4283,N_4192);
nor U8976 (N_8976,N_923,N_1159);
nor U8977 (N_8977,N_3981,N_2234);
and U8978 (N_8978,N_2927,N_2829);
nor U8979 (N_8979,N_3396,N_4605);
nand U8980 (N_8980,N_2458,N_1081);
or U8981 (N_8981,N_1717,N_3459);
nor U8982 (N_8982,N_221,N_4825);
and U8983 (N_8983,N_1762,N_1853);
or U8984 (N_8984,N_1481,N_4255);
xnor U8985 (N_8985,N_591,N_523);
nor U8986 (N_8986,N_2827,N_3599);
xnor U8987 (N_8987,N_1333,N_1893);
or U8988 (N_8988,N_4148,N_4748);
or U8989 (N_8989,N_3550,N_2376);
xnor U8990 (N_8990,N_2331,N_1853);
nand U8991 (N_8991,N_2767,N_1185);
xnor U8992 (N_8992,N_973,N_4473);
and U8993 (N_8993,N_2392,N_172);
or U8994 (N_8994,N_3731,N_1707);
xnor U8995 (N_8995,N_2465,N_4874);
xor U8996 (N_8996,N_480,N_2493);
xor U8997 (N_8997,N_814,N_351);
xnor U8998 (N_8998,N_3126,N_2779);
nor U8999 (N_8999,N_3058,N_3960);
nand U9000 (N_9000,N_1371,N_2134);
nand U9001 (N_9001,N_2929,N_4162);
and U9002 (N_9002,N_941,N_4216);
and U9003 (N_9003,N_2345,N_3408);
xor U9004 (N_9004,N_2381,N_4852);
and U9005 (N_9005,N_90,N_3824);
and U9006 (N_9006,N_579,N_4472);
nand U9007 (N_9007,N_2938,N_3924);
nor U9008 (N_9008,N_2685,N_2269);
xor U9009 (N_9009,N_3190,N_459);
nand U9010 (N_9010,N_964,N_51);
xnor U9011 (N_9011,N_2870,N_2974);
nand U9012 (N_9012,N_1593,N_1813);
or U9013 (N_9013,N_1213,N_328);
nor U9014 (N_9014,N_2945,N_4470);
xor U9015 (N_9015,N_3815,N_3672);
nor U9016 (N_9016,N_4834,N_377);
and U9017 (N_9017,N_2367,N_4593);
xor U9018 (N_9018,N_4576,N_1576);
nor U9019 (N_9019,N_1016,N_2704);
and U9020 (N_9020,N_2992,N_1274);
xnor U9021 (N_9021,N_668,N_1608);
nand U9022 (N_9022,N_1188,N_374);
and U9023 (N_9023,N_3363,N_4097);
or U9024 (N_9024,N_4750,N_4351);
nand U9025 (N_9025,N_785,N_450);
nor U9026 (N_9026,N_4496,N_4230);
xnor U9027 (N_9027,N_2424,N_2368);
nand U9028 (N_9028,N_4710,N_251);
and U9029 (N_9029,N_1672,N_3597);
or U9030 (N_9030,N_4198,N_2866);
or U9031 (N_9031,N_2767,N_2909);
or U9032 (N_9032,N_125,N_417);
nand U9033 (N_9033,N_3152,N_2761);
nand U9034 (N_9034,N_3993,N_2225);
xnor U9035 (N_9035,N_314,N_4308);
xnor U9036 (N_9036,N_1899,N_2687);
nor U9037 (N_9037,N_4231,N_857);
or U9038 (N_9038,N_1045,N_4883);
and U9039 (N_9039,N_2872,N_3231);
nand U9040 (N_9040,N_2941,N_2879);
or U9041 (N_9041,N_3635,N_4796);
xnor U9042 (N_9042,N_2476,N_1468);
and U9043 (N_9043,N_2344,N_3659);
and U9044 (N_9044,N_1848,N_308);
nand U9045 (N_9045,N_3972,N_2625);
or U9046 (N_9046,N_292,N_4878);
nand U9047 (N_9047,N_3197,N_906);
nand U9048 (N_9048,N_3903,N_259);
xnor U9049 (N_9049,N_4815,N_1521);
and U9050 (N_9050,N_2102,N_1870);
nand U9051 (N_9051,N_1776,N_3835);
and U9052 (N_9052,N_1481,N_711);
xor U9053 (N_9053,N_3213,N_2528);
nand U9054 (N_9054,N_1978,N_518);
or U9055 (N_9055,N_1601,N_35);
or U9056 (N_9056,N_2188,N_1179);
or U9057 (N_9057,N_4187,N_303);
nor U9058 (N_9058,N_711,N_544);
xnor U9059 (N_9059,N_4576,N_566);
xnor U9060 (N_9060,N_3167,N_9);
and U9061 (N_9061,N_1454,N_2417);
and U9062 (N_9062,N_4579,N_525);
or U9063 (N_9063,N_4408,N_2471);
and U9064 (N_9064,N_2751,N_2454);
nor U9065 (N_9065,N_4235,N_1018);
and U9066 (N_9066,N_2317,N_2947);
xnor U9067 (N_9067,N_655,N_3122);
and U9068 (N_9068,N_3195,N_4239);
xor U9069 (N_9069,N_3281,N_1501);
nand U9070 (N_9070,N_3556,N_2581);
nor U9071 (N_9071,N_1084,N_1257);
nand U9072 (N_9072,N_2094,N_1658);
nor U9073 (N_9073,N_32,N_4317);
nand U9074 (N_9074,N_366,N_1122);
nor U9075 (N_9075,N_2177,N_923);
nor U9076 (N_9076,N_4731,N_382);
or U9077 (N_9077,N_1543,N_3591);
nand U9078 (N_9078,N_2448,N_687);
xnor U9079 (N_9079,N_4760,N_4756);
or U9080 (N_9080,N_3509,N_159);
nand U9081 (N_9081,N_3264,N_1718);
xor U9082 (N_9082,N_3930,N_2395);
xor U9083 (N_9083,N_3667,N_457);
xnor U9084 (N_9084,N_1932,N_4520);
nand U9085 (N_9085,N_3907,N_3057);
or U9086 (N_9086,N_869,N_625);
and U9087 (N_9087,N_3803,N_4247);
and U9088 (N_9088,N_4180,N_2682);
nor U9089 (N_9089,N_1358,N_3979);
and U9090 (N_9090,N_785,N_3234);
nand U9091 (N_9091,N_4579,N_4678);
or U9092 (N_9092,N_945,N_3130);
nor U9093 (N_9093,N_2155,N_4763);
or U9094 (N_9094,N_2005,N_4317);
xnor U9095 (N_9095,N_350,N_139);
or U9096 (N_9096,N_3090,N_4041);
nor U9097 (N_9097,N_2403,N_889);
and U9098 (N_9098,N_4931,N_659);
and U9099 (N_9099,N_2761,N_4279);
xnor U9100 (N_9100,N_2895,N_1975);
nor U9101 (N_9101,N_824,N_1730);
and U9102 (N_9102,N_436,N_4502);
or U9103 (N_9103,N_2190,N_4361);
or U9104 (N_9104,N_3967,N_4868);
nand U9105 (N_9105,N_3737,N_2874);
nand U9106 (N_9106,N_3415,N_1624);
nand U9107 (N_9107,N_4556,N_4894);
nor U9108 (N_9108,N_584,N_976);
nor U9109 (N_9109,N_2194,N_537);
or U9110 (N_9110,N_4561,N_1964);
nor U9111 (N_9111,N_85,N_1602);
nand U9112 (N_9112,N_4711,N_4248);
nor U9113 (N_9113,N_4766,N_4692);
and U9114 (N_9114,N_3403,N_4486);
nand U9115 (N_9115,N_4458,N_2343);
nand U9116 (N_9116,N_3156,N_4987);
nand U9117 (N_9117,N_2335,N_4651);
or U9118 (N_9118,N_22,N_2387);
nand U9119 (N_9119,N_3016,N_3556);
xor U9120 (N_9120,N_2037,N_3622);
or U9121 (N_9121,N_3059,N_953);
nor U9122 (N_9122,N_3818,N_1050);
nor U9123 (N_9123,N_2780,N_655);
and U9124 (N_9124,N_2773,N_1261);
nand U9125 (N_9125,N_3938,N_2124);
nand U9126 (N_9126,N_3186,N_4013);
nor U9127 (N_9127,N_4379,N_1863);
and U9128 (N_9128,N_4397,N_2300);
and U9129 (N_9129,N_4816,N_4706);
nor U9130 (N_9130,N_1399,N_938);
and U9131 (N_9131,N_4135,N_414);
nand U9132 (N_9132,N_2006,N_4314);
nor U9133 (N_9133,N_793,N_235);
or U9134 (N_9134,N_2432,N_4717);
nor U9135 (N_9135,N_2732,N_739);
nand U9136 (N_9136,N_746,N_1559);
nor U9137 (N_9137,N_2325,N_4948);
xor U9138 (N_9138,N_3831,N_4558);
nor U9139 (N_9139,N_2315,N_3175);
nand U9140 (N_9140,N_2143,N_4110);
xnor U9141 (N_9141,N_2306,N_572);
nand U9142 (N_9142,N_3894,N_2501);
nor U9143 (N_9143,N_4059,N_4733);
nand U9144 (N_9144,N_3110,N_2188);
nor U9145 (N_9145,N_3467,N_2981);
nor U9146 (N_9146,N_895,N_1182);
nor U9147 (N_9147,N_2542,N_261);
nand U9148 (N_9148,N_1217,N_4475);
nor U9149 (N_9149,N_3984,N_3209);
xor U9150 (N_9150,N_1273,N_2418);
or U9151 (N_9151,N_4457,N_2762);
xor U9152 (N_9152,N_1700,N_120);
nand U9153 (N_9153,N_2943,N_3662);
or U9154 (N_9154,N_2085,N_3696);
nand U9155 (N_9155,N_2985,N_3169);
nor U9156 (N_9156,N_3967,N_4760);
nand U9157 (N_9157,N_1467,N_4558);
nand U9158 (N_9158,N_2228,N_4006);
or U9159 (N_9159,N_277,N_4379);
or U9160 (N_9160,N_4581,N_2487);
or U9161 (N_9161,N_4120,N_1296);
xnor U9162 (N_9162,N_4458,N_323);
xnor U9163 (N_9163,N_283,N_822);
xnor U9164 (N_9164,N_4624,N_1421);
nand U9165 (N_9165,N_3161,N_607);
nor U9166 (N_9166,N_1280,N_4817);
nor U9167 (N_9167,N_2867,N_2974);
xnor U9168 (N_9168,N_3655,N_387);
or U9169 (N_9169,N_4411,N_1965);
and U9170 (N_9170,N_838,N_2313);
nand U9171 (N_9171,N_1221,N_2604);
xor U9172 (N_9172,N_745,N_99);
xor U9173 (N_9173,N_43,N_8);
or U9174 (N_9174,N_4968,N_2440);
or U9175 (N_9175,N_4831,N_4286);
and U9176 (N_9176,N_4938,N_1222);
or U9177 (N_9177,N_3781,N_966);
and U9178 (N_9178,N_2825,N_1397);
nand U9179 (N_9179,N_580,N_2127);
xor U9180 (N_9180,N_2545,N_4477);
nor U9181 (N_9181,N_3077,N_88);
xor U9182 (N_9182,N_1407,N_141);
nand U9183 (N_9183,N_830,N_3751);
nand U9184 (N_9184,N_1587,N_728);
or U9185 (N_9185,N_803,N_1869);
xnor U9186 (N_9186,N_2412,N_3742);
xor U9187 (N_9187,N_31,N_2337);
nor U9188 (N_9188,N_792,N_2559);
or U9189 (N_9189,N_2416,N_2900);
nand U9190 (N_9190,N_173,N_1343);
or U9191 (N_9191,N_255,N_1388);
and U9192 (N_9192,N_4277,N_2112);
xor U9193 (N_9193,N_1278,N_449);
and U9194 (N_9194,N_4962,N_1943);
nand U9195 (N_9195,N_3235,N_448);
or U9196 (N_9196,N_1346,N_3384);
nor U9197 (N_9197,N_4219,N_4590);
or U9198 (N_9198,N_1139,N_2739);
or U9199 (N_9199,N_515,N_3016);
xnor U9200 (N_9200,N_4162,N_3112);
and U9201 (N_9201,N_1181,N_2384);
nand U9202 (N_9202,N_4800,N_3537);
nand U9203 (N_9203,N_3929,N_4765);
nand U9204 (N_9204,N_184,N_2871);
nor U9205 (N_9205,N_2010,N_3722);
and U9206 (N_9206,N_2700,N_3376);
nand U9207 (N_9207,N_2351,N_332);
nor U9208 (N_9208,N_4558,N_1668);
and U9209 (N_9209,N_2436,N_3408);
nand U9210 (N_9210,N_1091,N_462);
nor U9211 (N_9211,N_3702,N_2902);
nand U9212 (N_9212,N_3528,N_70);
nor U9213 (N_9213,N_4716,N_864);
nor U9214 (N_9214,N_3613,N_3694);
xor U9215 (N_9215,N_151,N_1554);
or U9216 (N_9216,N_104,N_639);
nand U9217 (N_9217,N_496,N_1792);
xor U9218 (N_9218,N_4793,N_4913);
and U9219 (N_9219,N_4725,N_3749);
nor U9220 (N_9220,N_1967,N_4221);
and U9221 (N_9221,N_4806,N_2812);
nor U9222 (N_9222,N_3440,N_4951);
xor U9223 (N_9223,N_106,N_1456);
xor U9224 (N_9224,N_1850,N_1493);
nor U9225 (N_9225,N_2666,N_2307);
or U9226 (N_9226,N_1628,N_755);
and U9227 (N_9227,N_287,N_1422);
or U9228 (N_9228,N_4734,N_4689);
and U9229 (N_9229,N_1371,N_930);
xnor U9230 (N_9230,N_4803,N_4789);
or U9231 (N_9231,N_2573,N_3693);
nor U9232 (N_9232,N_2822,N_3842);
nand U9233 (N_9233,N_2912,N_256);
nor U9234 (N_9234,N_1499,N_751);
and U9235 (N_9235,N_2532,N_2713);
or U9236 (N_9236,N_3173,N_952);
nor U9237 (N_9237,N_2928,N_4945);
nand U9238 (N_9238,N_2223,N_4450);
and U9239 (N_9239,N_4177,N_949);
nand U9240 (N_9240,N_540,N_2131);
xor U9241 (N_9241,N_4344,N_2000);
or U9242 (N_9242,N_1058,N_1470);
nor U9243 (N_9243,N_718,N_274);
xor U9244 (N_9244,N_3228,N_3104);
nor U9245 (N_9245,N_3918,N_350);
nand U9246 (N_9246,N_2448,N_1747);
and U9247 (N_9247,N_1515,N_3425);
nand U9248 (N_9248,N_1620,N_431);
nand U9249 (N_9249,N_3899,N_815);
nor U9250 (N_9250,N_1718,N_2629);
nor U9251 (N_9251,N_793,N_3832);
and U9252 (N_9252,N_3679,N_176);
nand U9253 (N_9253,N_2809,N_4982);
xor U9254 (N_9254,N_2701,N_1480);
or U9255 (N_9255,N_2171,N_1954);
and U9256 (N_9256,N_3921,N_3479);
and U9257 (N_9257,N_3309,N_4415);
nand U9258 (N_9258,N_2031,N_594);
xor U9259 (N_9259,N_729,N_726);
xor U9260 (N_9260,N_2409,N_3980);
nand U9261 (N_9261,N_816,N_4991);
nor U9262 (N_9262,N_2202,N_3806);
and U9263 (N_9263,N_100,N_3733);
nand U9264 (N_9264,N_3770,N_2772);
or U9265 (N_9265,N_1681,N_101);
nand U9266 (N_9266,N_3219,N_2754);
nand U9267 (N_9267,N_3542,N_4914);
nor U9268 (N_9268,N_496,N_504);
or U9269 (N_9269,N_1587,N_3227);
nand U9270 (N_9270,N_3475,N_20);
and U9271 (N_9271,N_3237,N_1462);
or U9272 (N_9272,N_3889,N_1009);
nand U9273 (N_9273,N_4731,N_2649);
or U9274 (N_9274,N_2180,N_4198);
xor U9275 (N_9275,N_4549,N_3480);
and U9276 (N_9276,N_3850,N_3490);
nand U9277 (N_9277,N_859,N_48);
xnor U9278 (N_9278,N_1726,N_137);
or U9279 (N_9279,N_4095,N_2073);
and U9280 (N_9280,N_1443,N_3812);
and U9281 (N_9281,N_143,N_844);
and U9282 (N_9282,N_4531,N_2444);
nor U9283 (N_9283,N_7,N_4352);
and U9284 (N_9284,N_4173,N_4142);
nor U9285 (N_9285,N_3401,N_3218);
or U9286 (N_9286,N_4091,N_1347);
xnor U9287 (N_9287,N_357,N_290);
nand U9288 (N_9288,N_3228,N_3467);
or U9289 (N_9289,N_2388,N_2327);
and U9290 (N_9290,N_457,N_2142);
nor U9291 (N_9291,N_3869,N_2341);
nand U9292 (N_9292,N_748,N_2625);
or U9293 (N_9293,N_3230,N_3355);
xnor U9294 (N_9294,N_3450,N_3764);
or U9295 (N_9295,N_4020,N_3480);
or U9296 (N_9296,N_2378,N_2698);
or U9297 (N_9297,N_300,N_2312);
xnor U9298 (N_9298,N_2564,N_2478);
xor U9299 (N_9299,N_607,N_4971);
xor U9300 (N_9300,N_3806,N_587);
xor U9301 (N_9301,N_326,N_3372);
nor U9302 (N_9302,N_609,N_3349);
xor U9303 (N_9303,N_3078,N_3403);
and U9304 (N_9304,N_1081,N_3151);
xnor U9305 (N_9305,N_2939,N_1923);
nor U9306 (N_9306,N_181,N_2908);
and U9307 (N_9307,N_817,N_464);
xnor U9308 (N_9308,N_479,N_4171);
nand U9309 (N_9309,N_4029,N_2882);
or U9310 (N_9310,N_4409,N_2693);
nand U9311 (N_9311,N_3886,N_3566);
and U9312 (N_9312,N_260,N_4605);
or U9313 (N_9313,N_686,N_688);
or U9314 (N_9314,N_3052,N_4946);
and U9315 (N_9315,N_2633,N_993);
nor U9316 (N_9316,N_1083,N_2607);
and U9317 (N_9317,N_4074,N_816);
xnor U9318 (N_9318,N_1012,N_1729);
xor U9319 (N_9319,N_3881,N_720);
or U9320 (N_9320,N_1098,N_1069);
xor U9321 (N_9321,N_1200,N_1897);
or U9322 (N_9322,N_758,N_1454);
nand U9323 (N_9323,N_4276,N_2352);
xnor U9324 (N_9324,N_3366,N_1965);
and U9325 (N_9325,N_1847,N_1352);
nor U9326 (N_9326,N_1975,N_377);
nand U9327 (N_9327,N_4711,N_635);
xor U9328 (N_9328,N_424,N_3272);
nor U9329 (N_9329,N_139,N_4028);
nand U9330 (N_9330,N_1540,N_1311);
or U9331 (N_9331,N_1042,N_3417);
and U9332 (N_9332,N_152,N_2659);
or U9333 (N_9333,N_2418,N_3691);
nor U9334 (N_9334,N_3159,N_1294);
nor U9335 (N_9335,N_777,N_2967);
xnor U9336 (N_9336,N_825,N_2207);
nand U9337 (N_9337,N_177,N_311);
and U9338 (N_9338,N_1340,N_1289);
nand U9339 (N_9339,N_3986,N_4808);
or U9340 (N_9340,N_221,N_4654);
or U9341 (N_9341,N_901,N_4606);
nor U9342 (N_9342,N_1211,N_1108);
xnor U9343 (N_9343,N_3962,N_3698);
xnor U9344 (N_9344,N_1501,N_1458);
xor U9345 (N_9345,N_4817,N_3888);
xor U9346 (N_9346,N_1653,N_3911);
nor U9347 (N_9347,N_3591,N_2719);
or U9348 (N_9348,N_4738,N_2928);
nor U9349 (N_9349,N_2858,N_1512);
or U9350 (N_9350,N_1912,N_2043);
nor U9351 (N_9351,N_4219,N_4462);
nand U9352 (N_9352,N_4676,N_1787);
or U9353 (N_9353,N_1731,N_1380);
nand U9354 (N_9354,N_1811,N_4650);
nor U9355 (N_9355,N_543,N_1679);
or U9356 (N_9356,N_4723,N_1466);
and U9357 (N_9357,N_34,N_584);
xor U9358 (N_9358,N_2655,N_2668);
xnor U9359 (N_9359,N_1562,N_660);
nor U9360 (N_9360,N_16,N_4589);
xor U9361 (N_9361,N_2818,N_1875);
nand U9362 (N_9362,N_3902,N_3473);
and U9363 (N_9363,N_966,N_1845);
nor U9364 (N_9364,N_4039,N_473);
nor U9365 (N_9365,N_2860,N_4647);
nor U9366 (N_9366,N_1464,N_4210);
or U9367 (N_9367,N_4893,N_2957);
and U9368 (N_9368,N_4117,N_1340);
nor U9369 (N_9369,N_4455,N_3430);
nand U9370 (N_9370,N_795,N_501);
xor U9371 (N_9371,N_2504,N_2690);
xnor U9372 (N_9372,N_1935,N_2628);
xor U9373 (N_9373,N_760,N_1698);
nor U9374 (N_9374,N_3023,N_592);
and U9375 (N_9375,N_3210,N_229);
xnor U9376 (N_9376,N_3437,N_1562);
and U9377 (N_9377,N_3272,N_2782);
nor U9378 (N_9378,N_517,N_2019);
or U9379 (N_9379,N_1569,N_1336);
nand U9380 (N_9380,N_1542,N_4795);
nor U9381 (N_9381,N_2016,N_1308);
nand U9382 (N_9382,N_4164,N_2246);
xor U9383 (N_9383,N_1006,N_1980);
xnor U9384 (N_9384,N_4683,N_3008);
nand U9385 (N_9385,N_3911,N_4240);
and U9386 (N_9386,N_3339,N_2859);
nand U9387 (N_9387,N_31,N_1855);
nand U9388 (N_9388,N_1269,N_2686);
xor U9389 (N_9389,N_3591,N_575);
or U9390 (N_9390,N_4207,N_1321);
xor U9391 (N_9391,N_2426,N_1279);
nor U9392 (N_9392,N_565,N_324);
xor U9393 (N_9393,N_1441,N_4587);
nand U9394 (N_9394,N_3337,N_1179);
and U9395 (N_9395,N_4497,N_454);
and U9396 (N_9396,N_772,N_2651);
or U9397 (N_9397,N_4453,N_1662);
xor U9398 (N_9398,N_4497,N_3874);
nor U9399 (N_9399,N_2971,N_2735);
xor U9400 (N_9400,N_4640,N_4150);
and U9401 (N_9401,N_3189,N_4850);
nor U9402 (N_9402,N_901,N_3006);
nor U9403 (N_9403,N_1519,N_4769);
nand U9404 (N_9404,N_1358,N_4529);
and U9405 (N_9405,N_609,N_4736);
and U9406 (N_9406,N_3364,N_1579);
nand U9407 (N_9407,N_3089,N_4224);
xor U9408 (N_9408,N_1084,N_2484);
and U9409 (N_9409,N_4600,N_1407);
and U9410 (N_9410,N_2696,N_1739);
nor U9411 (N_9411,N_3114,N_4852);
nor U9412 (N_9412,N_4259,N_3952);
nor U9413 (N_9413,N_1113,N_395);
and U9414 (N_9414,N_1044,N_3993);
and U9415 (N_9415,N_2378,N_2331);
xnor U9416 (N_9416,N_3606,N_1224);
nor U9417 (N_9417,N_2533,N_4817);
nand U9418 (N_9418,N_4625,N_2771);
xnor U9419 (N_9419,N_1768,N_3639);
xor U9420 (N_9420,N_2158,N_3399);
and U9421 (N_9421,N_2322,N_4543);
xnor U9422 (N_9422,N_3512,N_1333);
or U9423 (N_9423,N_3752,N_1367);
nand U9424 (N_9424,N_2577,N_4031);
and U9425 (N_9425,N_1552,N_463);
and U9426 (N_9426,N_136,N_920);
or U9427 (N_9427,N_3235,N_3382);
nor U9428 (N_9428,N_3102,N_3060);
or U9429 (N_9429,N_3590,N_4115);
nand U9430 (N_9430,N_1098,N_4441);
nor U9431 (N_9431,N_686,N_4906);
or U9432 (N_9432,N_1042,N_3042);
and U9433 (N_9433,N_1647,N_3242);
or U9434 (N_9434,N_1076,N_3374);
or U9435 (N_9435,N_925,N_1563);
xor U9436 (N_9436,N_1208,N_911);
nor U9437 (N_9437,N_754,N_3165);
xnor U9438 (N_9438,N_4965,N_1014);
nand U9439 (N_9439,N_487,N_3944);
xnor U9440 (N_9440,N_4085,N_259);
or U9441 (N_9441,N_2075,N_646);
xor U9442 (N_9442,N_579,N_3595);
and U9443 (N_9443,N_4075,N_207);
or U9444 (N_9444,N_1357,N_631);
xnor U9445 (N_9445,N_945,N_390);
xor U9446 (N_9446,N_2206,N_716);
nor U9447 (N_9447,N_1176,N_2863);
nand U9448 (N_9448,N_2806,N_2626);
nor U9449 (N_9449,N_2297,N_4043);
xnor U9450 (N_9450,N_844,N_4004);
nand U9451 (N_9451,N_1382,N_3067);
xor U9452 (N_9452,N_4865,N_787);
nand U9453 (N_9453,N_1878,N_2034);
nor U9454 (N_9454,N_3892,N_259);
nand U9455 (N_9455,N_3799,N_4933);
or U9456 (N_9456,N_794,N_1561);
nor U9457 (N_9457,N_2537,N_3887);
nand U9458 (N_9458,N_4251,N_1758);
nor U9459 (N_9459,N_504,N_4916);
nor U9460 (N_9460,N_4388,N_156);
nor U9461 (N_9461,N_2617,N_1265);
nand U9462 (N_9462,N_3145,N_3547);
nand U9463 (N_9463,N_4138,N_3033);
nand U9464 (N_9464,N_311,N_1783);
and U9465 (N_9465,N_3319,N_2967);
or U9466 (N_9466,N_4600,N_3790);
or U9467 (N_9467,N_4003,N_1497);
or U9468 (N_9468,N_2593,N_1810);
and U9469 (N_9469,N_3149,N_1827);
nand U9470 (N_9470,N_469,N_4501);
and U9471 (N_9471,N_1307,N_2451);
xor U9472 (N_9472,N_1972,N_4760);
xor U9473 (N_9473,N_2034,N_3883);
nand U9474 (N_9474,N_2653,N_3617);
nand U9475 (N_9475,N_3671,N_1624);
and U9476 (N_9476,N_938,N_593);
or U9477 (N_9477,N_2106,N_4630);
xnor U9478 (N_9478,N_570,N_1835);
or U9479 (N_9479,N_299,N_4396);
and U9480 (N_9480,N_3046,N_4982);
nor U9481 (N_9481,N_1981,N_1033);
or U9482 (N_9482,N_1100,N_2963);
nand U9483 (N_9483,N_3250,N_2578);
or U9484 (N_9484,N_1231,N_3967);
nor U9485 (N_9485,N_2954,N_2617);
or U9486 (N_9486,N_1482,N_4193);
nand U9487 (N_9487,N_3624,N_4978);
xor U9488 (N_9488,N_651,N_4939);
nor U9489 (N_9489,N_3106,N_624);
nor U9490 (N_9490,N_1266,N_2467);
and U9491 (N_9491,N_412,N_4913);
nor U9492 (N_9492,N_2817,N_1801);
nor U9493 (N_9493,N_94,N_1772);
nor U9494 (N_9494,N_2697,N_36);
xor U9495 (N_9495,N_2930,N_2355);
nor U9496 (N_9496,N_1193,N_2263);
or U9497 (N_9497,N_3793,N_3512);
or U9498 (N_9498,N_3964,N_2869);
nand U9499 (N_9499,N_684,N_4831);
xnor U9500 (N_9500,N_3542,N_3888);
nand U9501 (N_9501,N_1595,N_858);
xor U9502 (N_9502,N_1528,N_1862);
nand U9503 (N_9503,N_2046,N_3520);
or U9504 (N_9504,N_1997,N_931);
xnor U9505 (N_9505,N_4469,N_3317);
and U9506 (N_9506,N_782,N_1227);
nor U9507 (N_9507,N_2763,N_2403);
nand U9508 (N_9508,N_3842,N_3251);
nand U9509 (N_9509,N_2490,N_100);
or U9510 (N_9510,N_170,N_612);
nor U9511 (N_9511,N_3221,N_2191);
or U9512 (N_9512,N_922,N_2797);
and U9513 (N_9513,N_319,N_3157);
nor U9514 (N_9514,N_4127,N_2285);
or U9515 (N_9515,N_4483,N_2331);
nand U9516 (N_9516,N_4967,N_4120);
nor U9517 (N_9517,N_4817,N_758);
nand U9518 (N_9518,N_3395,N_1566);
and U9519 (N_9519,N_2947,N_4328);
xnor U9520 (N_9520,N_665,N_2187);
and U9521 (N_9521,N_2751,N_799);
or U9522 (N_9522,N_3297,N_4840);
xnor U9523 (N_9523,N_1937,N_854);
nand U9524 (N_9524,N_12,N_2299);
xor U9525 (N_9525,N_2814,N_1482);
or U9526 (N_9526,N_3643,N_1780);
and U9527 (N_9527,N_1327,N_1683);
nand U9528 (N_9528,N_61,N_4785);
nor U9529 (N_9529,N_4029,N_3885);
nor U9530 (N_9530,N_4735,N_4454);
or U9531 (N_9531,N_4901,N_4764);
or U9532 (N_9532,N_857,N_3666);
xor U9533 (N_9533,N_162,N_2929);
or U9534 (N_9534,N_2710,N_4985);
or U9535 (N_9535,N_3512,N_3451);
nor U9536 (N_9536,N_3229,N_4787);
or U9537 (N_9537,N_4873,N_1131);
or U9538 (N_9538,N_2899,N_1831);
xnor U9539 (N_9539,N_3391,N_1182);
nand U9540 (N_9540,N_3820,N_1211);
and U9541 (N_9541,N_4826,N_567);
nor U9542 (N_9542,N_4109,N_1637);
or U9543 (N_9543,N_1932,N_3511);
nor U9544 (N_9544,N_4504,N_593);
or U9545 (N_9545,N_3598,N_3353);
xor U9546 (N_9546,N_3456,N_4882);
and U9547 (N_9547,N_460,N_91);
nand U9548 (N_9548,N_3511,N_667);
nor U9549 (N_9549,N_2704,N_305);
or U9550 (N_9550,N_3198,N_3709);
or U9551 (N_9551,N_1636,N_4792);
nand U9552 (N_9552,N_3297,N_2991);
nand U9553 (N_9553,N_265,N_3890);
nor U9554 (N_9554,N_3406,N_1384);
and U9555 (N_9555,N_4378,N_3845);
or U9556 (N_9556,N_66,N_4694);
xor U9557 (N_9557,N_3691,N_3647);
nor U9558 (N_9558,N_3889,N_2040);
nor U9559 (N_9559,N_2164,N_3482);
nand U9560 (N_9560,N_2502,N_1148);
or U9561 (N_9561,N_4826,N_1496);
and U9562 (N_9562,N_768,N_3380);
xor U9563 (N_9563,N_2924,N_612);
nand U9564 (N_9564,N_124,N_4426);
and U9565 (N_9565,N_2217,N_769);
or U9566 (N_9566,N_549,N_415);
or U9567 (N_9567,N_4771,N_1142);
or U9568 (N_9568,N_1285,N_2126);
nor U9569 (N_9569,N_2286,N_1111);
xnor U9570 (N_9570,N_3849,N_865);
or U9571 (N_9571,N_1549,N_937);
xor U9572 (N_9572,N_2578,N_3280);
and U9573 (N_9573,N_3610,N_4563);
and U9574 (N_9574,N_1650,N_1155);
and U9575 (N_9575,N_2522,N_3378);
and U9576 (N_9576,N_175,N_451);
or U9577 (N_9577,N_1581,N_1017);
nor U9578 (N_9578,N_2858,N_4807);
nand U9579 (N_9579,N_1477,N_458);
nor U9580 (N_9580,N_1664,N_2158);
nand U9581 (N_9581,N_1019,N_4228);
or U9582 (N_9582,N_925,N_3949);
and U9583 (N_9583,N_559,N_2847);
nor U9584 (N_9584,N_3854,N_4834);
nand U9585 (N_9585,N_4536,N_3388);
and U9586 (N_9586,N_312,N_89);
or U9587 (N_9587,N_1769,N_4951);
xnor U9588 (N_9588,N_3922,N_716);
or U9589 (N_9589,N_443,N_1446);
nand U9590 (N_9590,N_3445,N_2813);
or U9591 (N_9591,N_2434,N_4298);
xor U9592 (N_9592,N_3529,N_4871);
nor U9593 (N_9593,N_2886,N_3067);
xnor U9594 (N_9594,N_158,N_590);
and U9595 (N_9595,N_1821,N_215);
xnor U9596 (N_9596,N_78,N_4762);
nor U9597 (N_9597,N_2350,N_2825);
nor U9598 (N_9598,N_424,N_2398);
xnor U9599 (N_9599,N_4379,N_4635);
or U9600 (N_9600,N_1609,N_2345);
nor U9601 (N_9601,N_3368,N_4868);
nand U9602 (N_9602,N_2513,N_4988);
or U9603 (N_9603,N_1476,N_3317);
and U9604 (N_9604,N_4411,N_2622);
xnor U9605 (N_9605,N_257,N_4067);
nor U9606 (N_9606,N_2982,N_1631);
and U9607 (N_9607,N_538,N_3477);
xnor U9608 (N_9608,N_3830,N_3986);
or U9609 (N_9609,N_656,N_4182);
or U9610 (N_9610,N_415,N_710);
or U9611 (N_9611,N_3601,N_3044);
xnor U9612 (N_9612,N_1159,N_309);
xnor U9613 (N_9613,N_3558,N_312);
or U9614 (N_9614,N_3124,N_4847);
xnor U9615 (N_9615,N_3089,N_2890);
or U9616 (N_9616,N_3532,N_4764);
nand U9617 (N_9617,N_466,N_2966);
xor U9618 (N_9618,N_1573,N_2774);
nor U9619 (N_9619,N_1794,N_1254);
or U9620 (N_9620,N_3720,N_2182);
and U9621 (N_9621,N_1622,N_38);
or U9622 (N_9622,N_4269,N_727);
or U9623 (N_9623,N_679,N_1124);
or U9624 (N_9624,N_4654,N_4029);
or U9625 (N_9625,N_538,N_2752);
nor U9626 (N_9626,N_2531,N_2408);
xnor U9627 (N_9627,N_4882,N_287);
nor U9628 (N_9628,N_3213,N_3401);
and U9629 (N_9629,N_3070,N_2956);
or U9630 (N_9630,N_1827,N_3733);
and U9631 (N_9631,N_3135,N_916);
and U9632 (N_9632,N_2121,N_508);
or U9633 (N_9633,N_2069,N_4551);
xnor U9634 (N_9634,N_3871,N_437);
nor U9635 (N_9635,N_2244,N_3530);
and U9636 (N_9636,N_474,N_4807);
nor U9637 (N_9637,N_1155,N_4058);
and U9638 (N_9638,N_4380,N_803);
and U9639 (N_9639,N_4293,N_4302);
or U9640 (N_9640,N_4299,N_3906);
and U9641 (N_9641,N_2496,N_1952);
and U9642 (N_9642,N_4605,N_1012);
and U9643 (N_9643,N_4625,N_2651);
xor U9644 (N_9644,N_709,N_456);
or U9645 (N_9645,N_1438,N_898);
nand U9646 (N_9646,N_578,N_4156);
nor U9647 (N_9647,N_429,N_1531);
nor U9648 (N_9648,N_3225,N_2457);
nand U9649 (N_9649,N_3482,N_2173);
xor U9650 (N_9650,N_3479,N_4406);
or U9651 (N_9651,N_4439,N_1316);
and U9652 (N_9652,N_214,N_3645);
nand U9653 (N_9653,N_3073,N_1494);
xor U9654 (N_9654,N_4559,N_242);
or U9655 (N_9655,N_2220,N_2359);
nor U9656 (N_9656,N_3864,N_1002);
xnor U9657 (N_9657,N_2312,N_2631);
nor U9658 (N_9658,N_3007,N_1113);
nor U9659 (N_9659,N_1412,N_4156);
nor U9660 (N_9660,N_4124,N_1830);
nor U9661 (N_9661,N_2320,N_2615);
or U9662 (N_9662,N_4863,N_1467);
nand U9663 (N_9663,N_233,N_1838);
xor U9664 (N_9664,N_1995,N_1285);
and U9665 (N_9665,N_1268,N_4471);
xnor U9666 (N_9666,N_336,N_2514);
xnor U9667 (N_9667,N_2815,N_441);
and U9668 (N_9668,N_1909,N_4230);
xor U9669 (N_9669,N_1809,N_2992);
and U9670 (N_9670,N_4830,N_730);
and U9671 (N_9671,N_1861,N_4928);
nor U9672 (N_9672,N_1881,N_3469);
or U9673 (N_9673,N_2334,N_1315);
nor U9674 (N_9674,N_2495,N_4867);
xor U9675 (N_9675,N_2013,N_816);
nand U9676 (N_9676,N_1978,N_1204);
xnor U9677 (N_9677,N_2909,N_3538);
nand U9678 (N_9678,N_299,N_1123);
or U9679 (N_9679,N_737,N_3342);
and U9680 (N_9680,N_2999,N_4518);
and U9681 (N_9681,N_692,N_887);
nand U9682 (N_9682,N_63,N_533);
or U9683 (N_9683,N_1988,N_1146);
xor U9684 (N_9684,N_4341,N_780);
and U9685 (N_9685,N_2110,N_4550);
nand U9686 (N_9686,N_232,N_4513);
nor U9687 (N_9687,N_1010,N_449);
nand U9688 (N_9688,N_348,N_3500);
nor U9689 (N_9689,N_4310,N_895);
nand U9690 (N_9690,N_1675,N_290);
nand U9691 (N_9691,N_4925,N_589);
xor U9692 (N_9692,N_3716,N_1096);
nand U9693 (N_9693,N_1598,N_3298);
nor U9694 (N_9694,N_541,N_2741);
xnor U9695 (N_9695,N_950,N_493);
nand U9696 (N_9696,N_1704,N_4996);
nand U9697 (N_9697,N_1641,N_3814);
or U9698 (N_9698,N_4254,N_854);
xor U9699 (N_9699,N_957,N_3188);
and U9700 (N_9700,N_3643,N_2655);
and U9701 (N_9701,N_68,N_2812);
nand U9702 (N_9702,N_748,N_2386);
nor U9703 (N_9703,N_4854,N_2280);
or U9704 (N_9704,N_518,N_3808);
xnor U9705 (N_9705,N_2865,N_2482);
nand U9706 (N_9706,N_3998,N_4873);
and U9707 (N_9707,N_649,N_4670);
nand U9708 (N_9708,N_2181,N_3310);
or U9709 (N_9709,N_1841,N_825);
nor U9710 (N_9710,N_3047,N_788);
nor U9711 (N_9711,N_4775,N_3536);
xor U9712 (N_9712,N_1909,N_475);
nand U9713 (N_9713,N_3170,N_845);
and U9714 (N_9714,N_3813,N_2234);
and U9715 (N_9715,N_3205,N_4153);
nand U9716 (N_9716,N_3395,N_1023);
nand U9717 (N_9717,N_1755,N_3915);
or U9718 (N_9718,N_1070,N_1841);
or U9719 (N_9719,N_1907,N_4161);
nand U9720 (N_9720,N_2304,N_389);
xor U9721 (N_9721,N_1963,N_2142);
or U9722 (N_9722,N_3959,N_2413);
xor U9723 (N_9723,N_2147,N_4362);
or U9724 (N_9724,N_2676,N_914);
xor U9725 (N_9725,N_413,N_1180);
nand U9726 (N_9726,N_191,N_224);
xor U9727 (N_9727,N_4525,N_4198);
or U9728 (N_9728,N_3903,N_513);
xor U9729 (N_9729,N_4175,N_1972);
and U9730 (N_9730,N_869,N_4216);
nand U9731 (N_9731,N_1447,N_2603);
nor U9732 (N_9732,N_4564,N_2799);
nor U9733 (N_9733,N_75,N_4671);
and U9734 (N_9734,N_2852,N_1373);
xor U9735 (N_9735,N_869,N_2233);
and U9736 (N_9736,N_3014,N_899);
and U9737 (N_9737,N_3974,N_770);
nand U9738 (N_9738,N_909,N_4002);
nor U9739 (N_9739,N_2783,N_4866);
nor U9740 (N_9740,N_3257,N_341);
and U9741 (N_9741,N_3244,N_486);
nor U9742 (N_9742,N_3899,N_1807);
nand U9743 (N_9743,N_363,N_1431);
and U9744 (N_9744,N_4038,N_4584);
nor U9745 (N_9745,N_1307,N_4008);
xor U9746 (N_9746,N_2136,N_1767);
and U9747 (N_9747,N_3122,N_2869);
and U9748 (N_9748,N_2855,N_2960);
xor U9749 (N_9749,N_215,N_51);
nand U9750 (N_9750,N_832,N_1263);
xnor U9751 (N_9751,N_4721,N_1887);
or U9752 (N_9752,N_4358,N_1920);
and U9753 (N_9753,N_1003,N_601);
nor U9754 (N_9754,N_2431,N_2690);
or U9755 (N_9755,N_3718,N_2115);
and U9756 (N_9756,N_4690,N_1728);
nor U9757 (N_9757,N_2603,N_1325);
nor U9758 (N_9758,N_1318,N_738);
and U9759 (N_9759,N_3954,N_3450);
or U9760 (N_9760,N_3237,N_2811);
or U9761 (N_9761,N_4873,N_3548);
or U9762 (N_9762,N_4747,N_1093);
nand U9763 (N_9763,N_3088,N_4219);
or U9764 (N_9764,N_1154,N_2526);
nand U9765 (N_9765,N_2638,N_725);
and U9766 (N_9766,N_3643,N_4919);
xor U9767 (N_9767,N_4719,N_623);
or U9768 (N_9768,N_1536,N_3382);
nand U9769 (N_9769,N_574,N_1930);
xnor U9770 (N_9770,N_3844,N_4787);
nand U9771 (N_9771,N_2399,N_2531);
xor U9772 (N_9772,N_3710,N_2605);
nand U9773 (N_9773,N_1475,N_1455);
xor U9774 (N_9774,N_813,N_4054);
xor U9775 (N_9775,N_1778,N_3752);
or U9776 (N_9776,N_3898,N_1835);
nand U9777 (N_9777,N_1518,N_201);
xor U9778 (N_9778,N_558,N_705);
nor U9779 (N_9779,N_1614,N_1955);
nor U9780 (N_9780,N_3287,N_2713);
xor U9781 (N_9781,N_4641,N_2663);
and U9782 (N_9782,N_724,N_1809);
xnor U9783 (N_9783,N_2754,N_3431);
nor U9784 (N_9784,N_4009,N_418);
or U9785 (N_9785,N_1606,N_794);
nand U9786 (N_9786,N_4493,N_4544);
and U9787 (N_9787,N_1979,N_2445);
or U9788 (N_9788,N_305,N_3618);
nor U9789 (N_9789,N_4889,N_2684);
xnor U9790 (N_9790,N_2584,N_549);
and U9791 (N_9791,N_3091,N_567);
nand U9792 (N_9792,N_389,N_4078);
nor U9793 (N_9793,N_814,N_225);
nand U9794 (N_9794,N_717,N_570);
nor U9795 (N_9795,N_3883,N_4029);
xnor U9796 (N_9796,N_3198,N_559);
nand U9797 (N_9797,N_218,N_4660);
nor U9798 (N_9798,N_532,N_4633);
and U9799 (N_9799,N_830,N_2815);
or U9800 (N_9800,N_3211,N_2879);
xnor U9801 (N_9801,N_3801,N_4571);
xor U9802 (N_9802,N_2874,N_1410);
or U9803 (N_9803,N_1959,N_1053);
or U9804 (N_9804,N_1738,N_729);
xor U9805 (N_9805,N_343,N_3308);
xor U9806 (N_9806,N_236,N_4523);
nor U9807 (N_9807,N_733,N_367);
nand U9808 (N_9808,N_2780,N_3147);
nor U9809 (N_9809,N_607,N_3169);
and U9810 (N_9810,N_4646,N_99);
nand U9811 (N_9811,N_2146,N_3826);
and U9812 (N_9812,N_3046,N_4960);
and U9813 (N_9813,N_827,N_4290);
or U9814 (N_9814,N_4585,N_4846);
nor U9815 (N_9815,N_3233,N_4551);
nand U9816 (N_9816,N_3077,N_421);
nor U9817 (N_9817,N_3810,N_2179);
nand U9818 (N_9818,N_3276,N_899);
nor U9819 (N_9819,N_2119,N_2610);
nor U9820 (N_9820,N_1262,N_4449);
nand U9821 (N_9821,N_2151,N_3784);
nor U9822 (N_9822,N_3662,N_3609);
nand U9823 (N_9823,N_2181,N_1905);
xor U9824 (N_9824,N_2255,N_2997);
nor U9825 (N_9825,N_3853,N_4496);
nand U9826 (N_9826,N_3812,N_960);
nor U9827 (N_9827,N_2029,N_3891);
or U9828 (N_9828,N_831,N_2127);
nand U9829 (N_9829,N_140,N_751);
nor U9830 (N_9830,N_2113,N_4362);
or U9831 (N_9831,N_4482,N_3965);
or U9832 (N_9832,N_4977,N_964);
or U9833 (N_9833,N_408,N_1672);
and U9834 (N_9834,N_4330,N_2144);
nand U9835 (N_9835,N_2993,N_2618);
and U9836 (N_9836,N_2359,N_4699);
xnor U9837 (N_9837,N_2038,N_4080);
nor U9838 (N_9838,N_3220,N_2859);
and U9839 (N_9839,N_2476,N_1178);
nand U9840 (N_9840,N_1086,N_1544);
xnor U9841 (N_9841,N_569,N_1313);
or U9842 (N_9842,N_2334,N_4893);
nor U9843 (N_9843,N_392,N_3608);
xor U9844 (N_9844,N_643,N_3949);
and U9845 (N_9845,N_2494,N_3121);
nor U9846 (N_9846,N_1419,N_2321);
xnor U9847 (N_9847,N_4298,N_1949);
and U9848 (N_9848,N_659,N_2317);
nand U9849 (N_9849,N_4251,N_696);
nor U9850 (N_9850,N_1671,N_1098);
and U9851 (N_9851,N_2174,N_4239);
nand U9852 (N_9852,N_4597,N_4037);
nand U9853 (N_9853,N_4536,N_1695);
xnor U9854 (N_9854,N_4578,N_928);
xnor U9855 (N_9855,N_4535,N_650);
nor U9856 (N_9856,N_2299,N_2067);
or U9857 (N_9857,N_1785,N_4214);
nor U9858 (N_9858,N_161,N_140);
and U9859 (N_9859,N_3977,N_1480);
xor U9860 (N_9860,N_1949,N_4473);
or U9861 (N_9861,N_2787,N_4824);
or U9862 (N_9862,N_3218,N_3051);
and U9863 (N_9863,N_384,N_4908);
and U9864 (N_9864,N_4413,N_4173);
nor U9865 (N_9865,N_2486,N_1427);
or U9866 (N_9866,N_2868,N_3955);
nor U9867 (N_9867,N_515,N_767);
xnor U9868 (N_9868,N_1556,N_410);
xor U9869 (N_9869,N_2844,N_287);
and U9870 (N_9870,N_3462,N_2119);
nor U9871 (N_9871,N_3318,N_812);
and U9872 (N_9872,N_3800,N_886);
or U9873 (N_9873,N_4837,N_1872);
and U9874 (N_9874,N_3141,N_1967);
nor U9875 (N_9875,N_3382,N_3055);
and U9876 (N_9876,N_339,N_2741);
xor U9877 (N_9877,N_3838,N_4962);
and U9878 (N_9878,N_2557,N_4240);
and U9879 (N_9879,N_2228,N_4229);
nand U9880 (N_9880,N_2916,N_2778);
xor U9881 (N_9881,N_548,N_1216);
and U9882 (N_9882,N_2456,N_1167);
and U9883 (N_9883,N_1297,N_537);
and U9884 (N_9884,N_1801,N_3916);
nand U9885 (N_9885,N_1932,N_1903);
xor U9886 (N_9886,N_2720,N_520);
xnor U9887 (N_9887,N_2534,N_4452);
and U9888 (N_9888,N_2866,N_37);
nand U9889 (N_9889,N_2393,N_4084);
nor U9890 (N_9890,N_1181,N_1384);
nor U9891 (N_9891,N_3075,N_989);
nand U9892 (N_9892,N_4202,N_3881);
xor U9893 (N_9893,N_1573,N_3353);
and U9894 (N_9894,N_3312,N_1344);
xnor U9895 (N_9895,N_3703,N_145);
nor U9896 (N_9896,N_2014,N_3542);
and U9897 (N_9897,N_4742,N_3549);
or U9898 (N_9898,N_2050,N_699);
xnor U9899 (N_9899,N_110,N_2926);
or U9900 (N_9900,N_2977,N_3190);
nand U9901 (N_9901,N_2258,N_990);
nand U9902 (N_9902,N_4589,N_3202);
xnor U9903 (N_9903,N_233,N_2718);
xnor U9904 (N_9904,N_612,N_4327);
or U9905 (N_9905,N_1488,N_841);
nor U9906 (N_9906,N_3435,N_1899);
or U9907 (N_9907,N_1654,N_2846);
or U9908 (N_9908,N_3637,N_3376);
nand U9909 (N_9909,N_851,N_637);
and U9910 (N_9910,N_2947,N_1782);
nor U9911 (N_9911,N_602,N_2109);
and U9912 (N_9912,N_3031,N_4549);
nand U9913 (N_9913,N_4307,N_1401);
xnor U9914 (N_9914,N_2232,N_1169);
xnor U9915 (N_9915,N_660,N_2054);
or U9916 (N_9916,N_158,N_3193);
nor U9917 (N_9917,N_2801,N_4730);
or U9918 (N_9918,N_2376,N_655);
nor U9919 (N_9919,N_322,N_2264);
and U9920 (N_9920,N_2498,N_1056);
nand U9921 (N_9921,N_3588,N_2144);
xor U9922 (N_9922,N_1022,N_694);
nand U9923 (N_9923,N_2778,N_4101);
and U9924 (N_9924,N_4870,N_257);
or U9925 (N_9925,N_1310,N_4317);
and U9926 (N_9926,N_4268,N_3846);
nand U9927 (N_9927,N_4282,N_740);
nor U9928 (N_9928,N_1820,N_4093);
nand U9929 (N_9929,N_4742,N_1826);
or U9930 (N_9930,N_3782,N_3810);
or U9931 (N_9931,N_1720,N_4376);
and U9932 (N_9932,N_3372,N_4);
nand U9933 (N_9933,N_4555,N_1050);
or U9934 (N_9934,N_2618,N_2619);
nand U9935 (N_9935,N_359,N_1335);
and U9936 (N_9936,N_1614,N_4942);
xnor U9937 (N_9937,N_1808,N_1822);
nand U9938 (N_9938,N_567,N_2274);
xor U9939 (N_9939,N_3008,N_3432);
nand U9940 (N_9940,N_2518,N_1725);
xnor U9941 (N_9941,N_3015,N_4318);
or U9942 (N_9942,N_2573,N_3429);
or U9943 (N_9943,N_3890,N_816);
or U9944 (N_9944,N_3248,N_439);
and U9945 (N_9945,N_4729,N_1343);
or U9946 (N_9946,N_2159,N_4900);
nand U9947 (N_9947,N_2850,N_509);
or U9948 (N_9948,N_2930,N_1341);
xnor U9949 (N_9949,N_2298,N_2978);
nor U9950 (N_9950,N_4380,N_2450);
and U9951 (N_9951,N_4889,N_1574);
xor U9952 (N_9952,N_2271,N_235);
or U9953 (N_9953,N_4406,N_406);
xnor U9954 (N_9954,N_2835,N_4032);
nor U9955 (N_9955,N_2653,N_1497);
or U9956 (N_9956,N_4590,N_683);
and U9957 (N_9957,N_4452,N_2347);
and U9958 (N_9958,N_4352,N_302);
nand U9959 (N_9959,N_3332,N_3360);
or U9960 (N_9960,N_4151,N_2737);
nor U9961 (N_9961,N_976,N_2793);
or U9962 (N_9962,N_4043,N_4605);
nand U9963 (N_9963,N_4863,N_4339);
xor U9964 (N_9964,N_3960,N_3727);
nor U9965 (N_9965,N_2500,N_1417);
nor U9966 (N_9966,N_971,N_2815);
xnor U9967 (N_9967,N_513,N_4961);
and U9968 (N_9968,N_647,N_2619);
xor U9969 (N_9969,N_1056,N_3401);
xnor U9970 (N_9970,N_4572,N_877);
xnor U9971 (N_9971,N_674,N_1111);
or U9972 (N_9972,N_3629,N_611);
or U9973 (N_9973,N_2652,N_3933);
xor U9974 (N_9974,N_1325,N_3658);
nor U9975 (N_9975,N_137,N_1629);
xor U9976 (N_9976,N_4622,N_914);
nand U9977 (N_9977,N_4755,N_3088);
nor U9978 (N_9978,N_1744,N_1943);
nand U9979 (N_9979,N_3749,N_169);
and U9980 (N_9980,N_3052,N_4443);
nand U9981 (N_9981,N_2857,N_4878);
nand U9982 (N_9982,N_4415,N_1810);
nor U9983 (N_9983,N_4699,N_3533);
or U9984 (N_9984,N_2406,N_2714);
nand U9985 (N_9985,N_2827,N_2342);
and U9986 (N_9986,N_234,N_4095);
or U9987 (N_9987,N_4572,N_853);
xnor U9988 (N_9988,N_4484,N_2444);
nor U9989 (N_9989,N_3545,N_3302);
nand U9990 (N_9990,N_4309,N_4258);
nand U9991 (N_9991,N_1642,N_4625);
nand U9992 (N_9992,N_3134,N_2500);
xor U9993 (N_9993,N_2399,N_2294);
nand U9994 (N_9994,N_3652,N_1071);
and U9995 (N_9995,N_4684,N_875);
or U9996 (N_9996,N_4485,N_3913);
xor U9997 (N_9997,N_4049,N_1120);
xnor U9998 (N_9998,N_664,N_2277);
and U9999 (N_9999,N_274,N_1746);
nand U10000 (N_10000,N_6101,N_9190);
nand U10001 (N_10001,N_8614,N_5065);
or U10002 (N_10002,N_6662,N_6854);
nand U10003 (N_10003,N_8883,N_6750);
nor U10004 (N_10004,N_6269,N_8469);
nor U10005 (N_10005,N_6680,N_7949);
nor U10006 (N_10006,N_7676,N_9552);
and U10007 (N_10007,N_5384,N_9254);
and U10008 (N_10008,N_7614,N_5140);
and U10009 (N_10009,N_6597,N_7522);
xor U10010 (N_10010,N_5704,N_7042);
nand U10011 (N_10011,N_8783,N_8298);
nor U10012 (N_10012,N_9954,N_9029);
nand U10013 (N_10013,N_5499,N_8775);
or U10014 (N_10014,N_9713,N_7056);
xnor U10015 (N_10015,N_8326,N_5356);
xor U10016 (N_10016,N_6963,N_8677);
and U10017 (N_10017,N_5759,N_5978);
nand U10018 (N_10018,N_7916,N_5173);
nand U10019 (N_10019,N_9590,N_9622);
xor U10020 (N_10020,N_6618,N_7343);
xor U10021 (N_10021,N_9785,N_8649);
nor U10022 (N_10022,N_7662,N_6641);
and U10023 (N_10023,N_5123,N_6142);
nor U10024 (N_10024,N_6874,N_6021);
xor U10025 (N_10025,N_6199,N_6716);
xnor U10026 (N_10026,N_7431,N_6454);
nor U10027 (N_10027,N_6962,N_9940);
nand U10028 (N_10028,N_8537,N_8514);
and U10029 (N_10029,N_6350,N_9361);
nand U10030 (N_10030,N_9213,N_7736);
and U10031 (N_10031,N_5203,N_5376);
or U10032 (N_10032,N_9161,N_7051);
nand U10033 (N_10033,N_6032,N_9673);
and U10034 (N_10034,N_9446,N_6188);
nand U10035 (N_10035,N_7638,N_7724);
nand U10036 (N_10036,N_7110,N_5523);
nor U10037 (N_10037,N_6494,N_6445);
nand U10038 (N_10038,N_5280,N_9686);
nand U10039 (N_10039,N_9155,N_7000);
xnor U10040 (N_10040,N_7053,N_6325);
xor U10041 (N_10041,N_8927,N_9826);
or U10042 (N_10042,N_6908,N_9019);
or U10043 (N_10043,N_9242,N_7268);
or U10044 (N_10044,N_6234,N_6848);
or U10045 (N_10045,N_8860,N_5038);
nand U10046 (N_10046,N_6590,N_6010);
nand U10047 (N_10047,N_9601,N_6150);
or U10048 (N_10048,N_5176,N_6310);
xor U10049 (N_10049,N_6564,N_9442);
nor U10050 (N_10050,N_5373,N_9831);
and U10051 (N_10051,N_6363,N_8088);
xnor U10052 (N_10052,N_9145,N_9219);
or U10053 (N_10053,N_7377,N_6258);
nand U10054 (N_10054,N_6600,N_6852);
nand U10055 (N_10055,N_7549,N_6755);
nor U10056 (N_10056,N_8542,N_9605);
xnor U10057 (N_10057,N_5104,N_7931);
xnor U10058 (N_10058,N_5096,N_5840);
xnor U10059 (N_10059,N_9803,N_8386);
xnor U10060 (N_10060,N_8475,N_5421);
nor U10061 (N_10061,N_8809,N_6155);
nand U10062 (N_10062,N_6922,N_9726);
nand U10063 (N_10063,N_6099,N_7791);
xor U10064 (N_10064,N_8167,N_5702);
xnor U10065 (N_10065,N_6460,N_8874);
xor U10066 (N_10066,N_9285,N_9259);
xnor U10067 (N_10067,N_6499,N_5733);
nand U10068 (N_10068,N_6529,N_5342);
xor U10069 (N_10069,N_7561,N_6562);
nor U10070 (N_10070,N_7565,N_6131);
and U10071 (N_10071,N_8376,N_5858);
and U10072 (N_10072,N_6047,N_6067);
nor U10073 (N_10073,N_5133,N_8072);
xor U10074 (N_10074,N_5456,N_6975);
xnor U10075 (N_10075,N_8019,N_7180);
nor U10076 (N_10076,N_8596,N_6532);
nand U10077 (N_10077,N_5198,N_6723);
nand U10078 (N_10078,N_8574,N_8193);
xor U10079 (N_10079,N_7124,N_8132);
nand U10080 (N_10080,N_9563,N_5420);
xor U10081 (N_10081,N_8262,N_8000);
and U10082 (N_10082,N_9407,N_7658);
and U10083 (N_10083,N_7450,N_7536);
nand U10084 (N_10084,N_6498,N_6385);
nand U10085 (N_10085,N_6735,N_6113);
xor U10086 (N_10086,N_5713,N_7941);
nor U10087 (N_10087,N_7818,N_5069);
nand U10088 (N_10088,N_8374,N_9595);
or U10089 (N_10089,N_6262,N_5363);
xnor U10090 (N_10090,N_5929,N_8719);
xnor U10091 (N_10091,N_5541,N_5721);
xnor U10092 (N_10092,N_5475,N_7102);
xnor U10093 (N_10093,N_7652,N_5352);
nand U10094 (N_10094,N_5579,N_7860);
nor U10095 (N_10095,N_7111,N_9090);
and U10096 (N_10096,N_7965,N_6221);
nor U10097 (N_10097,N_6598,N_7260);
nor U10098 (N_10098,N_5077,N_9972);
or U10099 (N_10099,N_7103,N_9174);
xnor U10100 (N_10100,N_5874,N_8936);
xor U10101 (N_10101,N_7326,N_5872);
xnor U10102 (N_10102,N_6521,N_6901);
or U10103 (N_10103,N_7654,N_6629);
xnor U10104 (N_10104,N_7025,N_6283);
xnor U10105 (N_10105,N_7933,N_6765);
or U10106 (N_10106,N_8538,N_5417);
nor U10107 (N_10107,N_7415,N_5243);
and U10108 (N_10108,N_9750,N_6913);
and U10109 (N_10109,N_6278,N_8906);
xnor U10110 (N_10110,N_7578,N_9465);
and U10111 (N_10111,N_6126,N_5265);
xnor U10112 (N_10112,N_7361,N_5349);
or U10113 (N_10113,N_7360,N_8738);
nor U10114 (N_10114,N_5418,N_8996);
nor U10115 (N_10115,N_6941,N_5740);
xnor U10116 (N_10116,N_8482,N_7412);
and U10117 (N_10117,N_8236,N_6009);
and U10118 (N_10118,N_5508,N_8346);
nand U10119 (N_10119,N_5620,N_7568);
nor U10120 (N_10120,N_7976,N_6374);
or U10121 (N_10121,N_7250,N_7942);
and U10122 (N_10122,N_8016,N_9941);
nand U10123 (N_10123,N_5246,N_7191);
and U10124 (N_10124,N_5518,N_9844);
or U10125 (N_10125,N_7126,N_7641);
or U10126 (N_10126,N_5783,N_8759);
nor U10127 (N_10127,N_6610,N_9433);
nand U10128 (N_10128,N_9882,N_8309);
xnor U10129 (N_10129,N_7834,N_5327);
nor U10130 (N_10130,N_9360,N_8826);
or U10131 (N_10131,N_8395,N_5683);
or U10132 (N_10132,N_8354,N_8337);
nand U10133 (N_10133,N_5980,N_6703);
nor U10134 (N_10134,N_7492,N_8120);
and U10135 (N_10135,N_6452,N_6907);
nand U10136 (N_10136,N_6068,N_8934);
xor U10137 (N_10137,N_5837,N_9818);
nor U10138 (N_10138,N_6117,N_7176);
and U10139 (N_10139,N_5430,N_9500);
or U10140 (N_10140,N_9860,N_5478);
nand U10141 (N_10141,N_9887,N_5900);
and U10142 (N_10142,N_9576,N_9345);
xor U10143 (N_10143,N_6541,N_7593);
and U10144 (N_10144,N_6468,N_5023);
xnor U10145 (N_10145,N_8917,N_6835);
nor U10146 (N_10146,N_8561,N_5146);
nor U10147 (N_10147,N_9405,N_7314);
nand U10148 (N_10148,N_9146,N_9722);
nand U10149 (N_10149,N_7152,N_8666);
and U10150 (N_10150,N_8413,N_9062);
nand U10151 (N_10151,N_9497,N_9933);
nor U10152 (N_10152,N_8185,N_7732);
xor U10153 (N_10153,N_5865,N_5528);
nand U10154 (N_10154,N_6060,N_8636);
and U10155 (N_10155,N_7021,N_8368);
xor U10156 (N_10156,N_7455,N_7763);
nand U10157 (N_10157,N_5234,N_5167);
nor U10158 (N_10158,N_5545,N_8822);
and U10159 (N_10159,N_7304,N_7609);
or U10160 (N_10160,N_5469,N_5256);
nand U10161 (N_10161,N_8334,N_7703);
nand U10162 (N_10162,N_7892,N_9706);
nand U10163 (N_10163,N_6065,N_7777);
nor U10164 (N_10164,N_9178,N_5798);
and U10165 (N_10165,N_6991,N_7439);
or U10166 (N_10166,N_8194,N_5304);
nor U10167 (N_10167,N_9978,N_6790);
nand U10168 (N_10168,N_5306,N_9228);
xnor U10169 (N_10169,N_6326,N_5583);
or U10170 (N_10170,N_7929,N_7657);
and U10171 (N_10171,N_8231,N_6253);
and U10172 (N_10172,N_9124,N_6108);
nor U10173 (N_10173,N_7575,N_6298);
xnor U10174 (N_10174,N_6145,N_9930);
nor U10175 (N_10175,N_6589,N_7795);
xor U10176 (N_10176,N_5088,N_9028);
or U10177 (N_10177,N_7095,N_8720);
nand U10178 (N_10178,N_7643,N_5685);
nand U10179 (N_10179,N_7969,N_6969);
nand U10180 (N_10180,N_9589,N_9164);
or U10181 (N_10181,N_8498,N_9277);
xor U10182 (N_10182,N_7307,N_7623);
and U10183 (N_10183,N_6574,N_8074);
nor U10184 (N_10184,N_7980,N_6467);
or U10185 (N_10185,N_8307,N_8530);
or U10186 (N_10186,N_7369,N_7295);
and U10187 (N_10187,N_7153,N_7348);
nand U10188 (N_10188,N_5419,N_7092);
or U10189 (N_10189,N_8083,N_9044);
nand U10190 (N_10190,N_9583,N_6547);
xnor U10191 (N_10191,N_5789,N_8659);
nor U10192 (N_10192,N_5742,N_5559);
xnor U10193 (N_10193,N_8572,N_6213);
nand U10194 (N_10194,N_8246,N_9975);
nand U10195 (N_10195,N_5182,N_7039);
or U10196 (N_10196,N_7443,N_7221);
and U10197 (N_10197,N_9293,N_5926);
and U10198 (N_10198,N_7693,N_6202);
or U10199 (N_10199,N_5242,N_8004);
xnor U10200 (N_10200,N_5490,N_7647);
or U10201 (N_10201,N_6895,N_5054);
or U10202 (N_10202,N_9709,N_7774);
and U10203 (N_10203,N_8159,N_5962);
nand U10204 (N_10204,N_9689,N_9435);
nand U10205 (N_10205,N_7273,N_6870);
or U10206 (N_10206,N_6224,N_9564);
or U10207 (N_10207,N_7616,N_6942);
nand U10208 (N_10208,N_5932,N_7127);
and U10209 (N_10209,N_5017,N_8364);
or U10210 (N_10210,N_5928,N_8634);
nand U10211 (N_10211,N_8076,N_8771);
and U10212 (N_10212,N_9685,N_9241);
xnor U10213 (N_10213,N_9936,N_6539);
nor U10214 (N_10214,N_7441,N_7872);
nand U10215 (N_10215,N_7203,N_7007);
xor U10216 (N_10216,N_6190,N_7179);
nor U10217 (N_10217,N_7634,N_6809);
xor U10218 (N_10218,N_6658,N_7481);
and U10219 (N_10219,N_8734,N_6837);
nor U10220 (N_10220,N_9490,N_8360);
or U10221 (N_10221,N_6053,N_7253);
or U10222 (N_10222,N_8685,N_9392);
and U10223 (N_10223,N_6492,N_7138);
and U10224 (N_10224,N_8547,N_6265);
or U10225 (N_10225,N_7383,N_6977);
nor U10226 (N_10226,N_9870,N_9665);
xor U10227 (N_10227,N_5340,N_5682);
and U10228 (N_10228,N_6796,N_8317);
nor U10229 (N_10229,N_9886,N_7507);
nor U10230 (N_10230,N_5606,N_6125);
xor U10231 (N_10231,N_9784,N_5771);
nor U10232 (N_10232,N_8782,N_8447);
nor U10233 (N_10233,N_6517,N_5209);
nand U10234 (N_10234,N_5882,N_9206);
xor U10235 (N_10235,N_5515,N_5911);
nor U10236 (N_10236,N_6197,N_8095);
nand U10237 (N_10237,N_8950,N_8411);
nor U10238 (N_10238,N_9896,N_9512);
and U10239 (N_10239,N_6305,N_7466);
nor U10240 (N_10240,N_7216,N_9848);
and U10241 (N_10241,N_6888,N_8825);
or U10242 (N_10242,N_5153,N_5194);
nor U10243 (N_10243,N_9305,N_8150);
nor U10244 (N_10244,N_5630,N_7223);
xnor U10245 (N_10245,N_7644,N_8141);
xor U10246 (N_10246,N_6250,N_9515);
nor U10247 (N_10247,N_5205,N_6863);
nand U10248 (N_10248,N_7434,N_6294);
and U10249 (N_10249,N_9953,N_5655);
or U10250 (N_10250,N_7925,N_7493);
xor U10251 (N_10251,N_5122,N_6583);
nor U10252 (N_10252,N_8885,N_6228);
xnor U10253 (N_10253,N_8931,N_5378);
and U10254 (N_10254,N_8516,N_5633);
and U10255 (N_10255,N_6840,N_8375);
xor U10256 (N_10256,N_9203,N_7318);
or U10257 (N_10257,N_8505,N_8899);
nor U10258 (N_10258,N_8568,N_8701);
and U10259 (N_10259,N_7656,N_9885);
nor U10260 (N_10260,N_9710,N_7453);
xor U10261 (N_10261,N_6334,N_6940);
and U10262 (N_10262,N_9976,N_9063);
or U10263 (N_10263,N_8222,N_5641);
nand U10264 (N_10264,N_9276,N_6075);
nand U10265 (N_10265,N_5611,N_7875);
nor U10266 (N_10266,N_7890,N_7028);
nand U10267 (N_10267,N_7972,N_6005);
and U10268 (N_10268,N_8502,N_5811);
or U10269 (N_10269,N_7635,N_9175);
nor U10270 (N_10270,N_9142,N_5557);
or U10271 (N_10271,N_5647,N_5817);
nor U10272 (N_10272,N_8446,N_8722);
nand U10273 (N_10273,N_6024,N_5897);
or U10274 (N_10274,N_8357,N_9874);
and U10275 (N_10275,N_9973,N_6842);
and U10276 (N_10276,N_6509,N_5695);
nand U10277 (N_10277,N_6572,N_7444);
xor U10278 (N_10278,N_8064,N_6910);
and U10279 (N_10279,N_8247,N_9728);
xnor U10280 (N_10280,N_7442,N_7893);
or U10281 (N_10281,N_5072,N_6898);
nor U10282 (N_10282,N_7040,N_6011);
and U10283 (N_10283,N_8316,N_8990);
and U10284 (N_10284,N_9900,N_8291);
nor U10285 (N_10285,N_5890,N_5286);
xnor U10286 (N_10286,N_8163,N_5283);
nand U10287 (N_10287,N_7899,N_7086);
and U10288 (N_10288,N_9569,N_9895);
and U10289 (N_10289,N_7143,N_9267);
xnor U10290 (N_10290,N_7934,N_9861);
nand U10291 (N_10291,N_5662,N_8654);
xnor U10292 (N_10292,N_7224,N_6348);
and U10293 (N_10293,N_8292,N_6072);
or U10294 (N_10294,N_8420,N_5440);
nor U10295 (N_10295,N_5341,N_6535);
and U10296 (N_10296,N_7024,N_7142);
or U10297 (N_10297,N_6001,N_6554);
nor U10298 (N_10298,N_7731,N_8708);
nor U10299 (N_10299,N_7470,N_5521);
and U10300 (N_10300,N_8331,N_5687);
and U10301 (N_10301,N_5324,N_5555);
nand U10302 (N_10302,N_6829,N_8158);
nand U10303 (N_10303,N_9881,N_7873);
nand U10304 (N_10304,N_9399,N_8339);
xor U10305 (N_10305,N_6954,N_9769);
nor U10306 (N_10306,N_5019,N_8044);
nand U10307 (N_10307,N_6420,N_7744);
and U10308 (N_10308,N_5480,N_9693);
xnor U10309 (N_10309,N_5152,N_5726);
nor U10310 (N_10310,N_9107,N_8245);
nor U10311 (N_10311,N_7107,N_5329);
nand U10312 (N_10312,N_9716,N_8059);
nand U10313 (N_10313,N_9475,N_7263);
nor U10314 (N_10314,N_8126,N_7397);
nor U10315 (N_10315,N_7772,N_6791);
and U10316 (N_10316,N_9245,N_7150);
and U10317 (N_10317,N_6316,N_8090);
nor U10318 (N_10318,N_9695,N_6130);
or U10319 (N_10319,N_5032,N_7780);
xnor U10320 (N_10320,N_8746,N_7637);
nand U10321 (N_10321,N_6916,N_5714);
nor U10322 (N_10322,N_5427,N_5930);
and U10323 (N_10323,N_7759,N_8940);
and U10324 (N_10324,N_7388,N_5041);
nor U10325 (N_10325,N_6869,N_8871);
nor U10326 (N_10326,N_9408,N_6380);
nor U10327 (N_10327,N_9658,N_6612);
or U10328 (N_10328,N_7692,N_9151);
nand U10329 (N_10329,N_8554,N_8875);
nor U10330 (N_10330,N_8641,N_7132);
and U10331 (N_10331,N_9329,N_5253);
nand U10332 (N_10332,N_6948,N_8788);
nor U10333 (N_10333,N_8170,N_7541);
nand U10334 (N_10334,N_9113,N_6616);
xnor U10335 (N_10335,N_5411,N_5796);
and U10336 (N_10336,N_7236,N_9890);
nor U10337 (N_10337,N_7089,N_5048);
nand U10338 (N_10338,N_8551,N_8526);
and U10339 (N_10339,N_9415,N_5264);
xor U10340 (N_10340,N_7543,N_7300);
xnor U10341 (N_10341,N_5689,N_7427);
and U10342 (N_10342,N_5944,N_9369);
xnor U10343 (N_10343,N_7581,N_7385);
and U10344 (N_10344,N_5806,N_9342);
nand U10345 (N_10345,N_6872,N_8600);
and U10346 (N_10346,N_5103,N_8663);
and U10347 (N_10347,N_5617,N_6439);
and U10348 (N_10348,N_7174,N_9121);
xnor U10349 (N_10349,N_7367,N_8790);
xor U10350 (N_10350,N_7712,N_6759);
nor U10351 (N_10351,N_6409,N_6432);
or U10352 (N_10352,N_6438,N_9115);
or U10353 (N_10353,N_8112,N_5139);
and U10354 (N_10354,N_6244,N_8961);
nand U10355 (N_10355,N_6064,N_7014);
nor U10356 (N_10356,N_9303,N_9341);
and U10357 (N_10357,N_5595,N_7472);
nor U10358 (N_10358,N_8145,N_8872);
nor U10359 (N_10359,N_9042,N_9205);
nor U10360 (N_10360,N_7707,N_5912);
and U10361 (N_10361,N_6904,N_5948);
xor U10362 (N_10362,N_9774,N_8787);
xnor U10363 (N_10363,N_7109,N_8947);
and U10364 (N_10364,N_8035,N_7436);
and U10365 (N_10365,N_8082,N_9776);
nor U10366 (N_10366,N_9440,N_6285);
xor U10367 (N_10367,N_9328,N_9287);
nor U10368 (N_10368,N_5206,N_6366);
xnor U10369 (N_10369,N_7420,N_6792);
and U10370 (N_10370,N_8517,N_9035);
or U10371 (N_10371,N_6403,N_6646);
xor U10372 (N_10372,N_9112,N_6045);
and U10373 (N_10373,N_6605,N_5999);
nand U10374 (N_10374,N_7357,N_7363);
and U10375 (N_10375,N_6700,N_6328);
or U10376 (N_10376,N_7672,N_9625);
nand U10377 (N_10377,N_7359,N_8509);
nor U10378 (N_10378,N_6448,N_9809);
and U10379 (N_10379,N_9662,N_9983);
nand U10380 (N_10380,N_7349,N_8661);
and U10381 (N_10381,N_8199,N_7294);
and U10382 (N_10382,N_6808,N_8887);
nand U10383 (N_10383,N_9729,N_7022);
and U10384 (N_10384,N_9770,N_8816);
and U10385 (N_10385,N_8370,N_5387);
xnor U10386 (N_10386,N_6714,N_9891);
xnor U10387 (N_10387,N_9236,N_5942);
xor U10388 (N_10388,N_7468,N_7544);
nor U10389 (N_10389,N_9553,N_6665);
or U10390 (N_10390,N_7789,N_8018);
xnor U10391 (N_10391,N_9478,N_5879);
or U10392 (N_10392,N_7854,N_5201);
nor U10393 (N_10393,N_6480,N_9901);
nand U10394 (N_10394,N_8340,N_8136);
nor U10395 (N_10395,N_7379,N_9179);
nand U10396 (N_10396,N_8266,N_7782);
xnor U10397 (N_10397,N_9911,N_8415);
nand U10398 (N_10398,N_7998,N_5675);
and U10399 (N_10399,N_5805,N_9459);
nor U10400 (N_10400,N_5863,N_9763);
and U10401 (N_10401,N_9951,N_8905);
or U10402 (N_10402,N_6995,N_8534);
and U10403 (N_10403,N_6543,N_6429);
nand U10404 (N_10404,N_8117,N_9920);
or U10405 (N_10405,N_5601,N_9340);
nor U10406 (N_10406,N_5985,N_6819);
or U10407 (N_10407,N_7508,N_5414);
xor U10408 (N_10408,N_7469,N_7401);
nor U10409 (N_10409,N_6857,N_6151);
and U10410 (N_10410,N_6764,N_8249);
nor U10411 (N_10411,N_5287,N_7937);
xor U10412 (N_10412,N_7446,N_7560);
xnor U10413 (N_10413,N_6946,N_7999);
nand U10414 (N_10414,N_5272,N_7766);
or U10415 (N_10415,N_5836,N_6820);
nor U10416 (N_10416,N_6877,N_9637);
or U10417 (N_10417,N_5628,N_9410);
nor U10418 (N_10418,N_5336,N_6961);
xor U10419 (N_10419,N_9962,N_7210);
nor U10420 (N_10420,N_6324,N_5215);
nand U10421 (N_10421,N_9756,N_6440);
xnor U10422 (N_10422,N_8926,N_5268);
xor U10423 (N_10423,N_8098,N_5960);
nor U10424 (N_10424,N_8909,N_6177);
nand U10425 (N_10425,N_7402,N_6553);
xor U10426 (N_10426,N_6035,N_6036);
nor U10427 (N_10427,N_9130,N_8671);
or U10428 (N_10428,N_8847,N_7938);
xnor U10429 (N_10429,N_5860,N_7001);
and U10430 (N_10430,N_9078,N_8977);
and U10431 (N_10431,N_9788,N_5361);
or U10432 (N_10432,N_8692,N_9334);
and U10433 (N_10433,N_6319,N_8870);
nor U10434 (N_10434,N_7905,N_6172);
and U10435 (N_10435,N_8118,N_8405);
nand U10436 (N_10436,N_5642,N_9908);
and U10437 (N_10437,N_6091,N_8821);
nor U10438 (N_10438,N_7131,N_7205);
xor U10439 (N_10439,N_8608,N_8984);
or U10440 (N_10440,N_9066,N_5998);
nor U10441 (N_10441,N_6805,N_9696);
nor U10442 (N_10442,N_5185,N_8876);
nor U10443 (N_10443,N_7997,N_9129);
and U10444 (N_10444,N_5639,N_7832);
or U10445 (N_10445,N_7633,N_8862);
and U10446 (N_10446,N_9862,N_5461);
nand U10447 (N_10447,N_6653,N_6622);
and U10448 (N_10448,N_9220,N_5851);
or U10449 (N_10449,N_5121,N_9131);
xnor U10450 (N_10450,N_7606,N_5807);
or U10451 (N_10451,N_9742,N_5619);
nand U10452 (N_10452,N_7417,N_7192);
and U10453 (N_10453,N_9672,N_9543);
or U10454 (N_10454,N_7355,N_6892);
or U10455 (N_10455,N_6210,N_7322);
nand U10456 (N_10456,N_6463,N_6523);
and U10457 (N_10457,N_7002,N_7320);
nand U10458 (N_10458,N_6027,N_9389);
nand U10459 (N_10459,N_6191,N_6070);
or U10460 (N_10460,N_6431,N_5666);
or U10461 (N_10461,N_6849,N_9148);
and U10462 (N_10462,N_6165,N_9509);
nor U10463 (N_10463,N_5869,N_6433);
or U10464 (N_10464,N_5696,N_8010);
xnor U10465 (N_10465,N_6747,N_6660);
and U10466 (N_10466,N_9501,N_5514);
nor U10467 (N_10467,N_7052,N_8038);
and U10468 (N_10468,N_8699,N_5976);
nor U10469 (N_10469,N_9064,N_7806);
or U10470 (N_10470,N_8800,N_6745);
or U10471 (N_10471,N_5544,N_5204);
and U10472 (N_10472,N_6472,N_7297);
xnor U10473 (N_10473,N_6497,N_7995);
xor U10474 (N_10474,N_5765,N_8873);
nand U10475 (N_10475,N_5907,N_8901);
or U10476 (N_10476,N_7225,N_9336);
nor U10477 (N_10477,N_9181,N_7975);
or U10478 (N_10478,N_7050,N_5612);
or U10479 (N_10479,N_8029,N_5993);
or U10480 (N_10480,N_9652,N_7958);
nand U10481 (N_10481,N_7113,N_5729);
nand U10482 (N_10482,N_7309,N_9667);
nor U10483 (N_10483,N_7121,N_6772);
or U10484 (N_10484,N_8173,N_6314);
nor U10485 (N_10485,N_6181,N_9540);
xnor U10486 (N_10486,N_8588,N_8327);
and U10487 (N_10487,N_6783,N_9068);
or U10488 (N_10488,N_5901,N_5084);
nor U10489 (N_10489,N_8229,N_6821);
xnor U10490 (N_10490,N_9597,N_5070);
or U10491 (N_10491,N_6955,N_5006);
or U10492 (N_10492,N_8287,N_9486);
nor U10493 (N_10493,N_5558,N_7093);
or U10494 (N_10494,N_9257,N_9613);
xnor U10495 (N_10495,N_6540,N_9432);
and U10496 (N_10496,N_7666,N_6778);
nand U10497 (N_10497,N_5366,N_5569);
nor U10498 (N_10498,N_5149,N_8854);
or U10499 (N_10499,N_9524,N_9401);
or U10500 (N_10500,N_6087,N_8243);
or U10501 (N_10501,N_7213,N_5160);
xor U10502 (N_10502,N_8866,N_9153);
xnor U10503 (N_10503,N_6376,N_8465);
nor U10504 (N_10504,N_9720,N_6466);
and U10505 (N_10505,N_5142,N_8487);
xor U10506 (N_10506,N_7953,N_5660);
or U10507 (N_10507,N_7168,N_9663);
nor U10508 (N_10508,N_5255,N_6186);
nand U10509 (N_10509,N_9030,N_9079);
and U10510 (N_10510,N_5525,N_8383);
and U10511 (N_10511,N_6341,N_8426);
and U10512 (N_10512,N_7691,N_8938);
xnor U10513 (N_10513,N_5130,N_8494);
and U10514 (N_10514,N_9226,N_5476);
or U10515 (N_10515,N_9183,N_5575);
and U10516 (N_10516,N_6650,N_5720);
or U10517 (N_10517,N_6028,N_9103);
nor U10518 (N_10518,N_8815,N_8282);
nor U10519 (N_10519,N_9905,N_5574);
and U10520 (N_10520,N_5883,N_5290);
nor U10521 (N_10521,N_5030,N_8717);
or U10522 (N_10522,N_7188,N_6671);
xnor U10523 (N_10523,N_9436,N_7499);
or U10524 (N_10524,N_7811,N_7342);
or U10525 (N_10525,N_8645,N_9996);
nand U10526 (N_10526,N_8226,N_7917);
and U10527 (N_10527,N_5227,N_7135);
nor U10528 (N_10528,N_7869,N_7010);
nor U10529 (N_10529,N_8599,N_5994);
and U10530 (N_10530,N_9768,N_7098);
and U10531 (N_10531,N_7084,N_5034);
nand U10532 (N_10532,N_5403,N_5891);
and U10533 (N_10533,N_8148,N_7407);
or U10534 (N_10534,N_9570,N_8884);
nand U10535 (N_10535,N_6359,N_6798);
and U10536 (N_10536,N_6824,N_5086);
xnor U10537 (N_10537,N_7796,N_5320);
nand U10538 (N_10538,N_5552,N_9222);
nand U10539 (N_10539,N_6971,N_8868);
xor U10540 (N_10540,N_8253,N_6885);
xor U10541 (N_10541,N_7101,N_9707);
and U10542 (N_10542,N_5024,N_7206);
nand U10543 (N_10543,N_7483,N_6549);
nor U10544 (N_10544,N_5331,N_8479);
and U10545 (N_10545,N_6174,N_7923);
or U10546 (N_10546,N_6766,N_8020);
nand U10547 (N_10547,N_9347,N_6882);
nor U10548 (N_10548,N_6012,N_7595);
or U10549 (N_10549,N_6303,N_8916);
or U10550 (N_10550,N_7038,N_8976);
xnor U10551 (N_10551,N_8155,N_6457);
or U10552 (N_10552,N_7408,N_9926);
nand U10553 (N_10553,N_5230,N_6382);
nand U10554 (N_10554,N_5681,N_6743);
nand U10555 (N_10555,N_6508,N_8613);
or U10556 (N_10556,N_6370,N_6301);
nor U10557 (N_10557,N_8466,N_9320);
and U10558 (N_10558,N_7484,N_8971);
or U10559 (N_10559,N_8280,N_5593);
and U10560 (N_10560,N_9959,N_5522);
nor U10561 (N_10561,N_6566,N_8552);
nor U10562 (N_10562,N_9538,N_6287);
xnor U10563 (N_10563,N_9152,N_7338);
nand U10564 (N_10564,N_5279,N_9758);
xnor U10565 (N_10565,N_8433,N_5066);
or U10566 (N_10566,N_8784,N_9839);
and U10567 (N_10567,N_6683,N_9521);
or U10568 (N_10568,N_5766,N_9099);
nor U10569 (N_10569,N_6833,N_5652);
xnor U10570 (N_10570,N_6694,N_5827);
nand U10571 (N_10571,N_8056,N_8628);
nor U10572 (N_10572,N_8994,N_6693);
and U10573 (N_10573,N_5531,N_7345);
nand U10574 (N_10574,N_5894,N_9310);
nand U10575 (N_10575,N_8937,N_6020);
or U10576 (N_10576,N_9780,N_7296);
xnor U10577 (N_10577,N_6899,N_7773);
or U10578 (N_10578,N_7520,N_8259);
xnor U10579 (N_10579,N_5275,N_9123);
and U10580 (N_10580,N_9733,N_5902);
and U10581 (N_10581,N_7846,N_5546);
nand U10582 (N_10582,N_8171,N_5097);
xnor U10583 (N_10583,N_7029,N_6416);
or U10584 (N_10584,N_7758,N_6295);
nor U10585 (N_10585,N_8102,N_6736);
nand U10586 (N_10586,N_9302,N_7735);
or U10587 (N_10587,N_6640,N_6691);
xor U10588 (N_10588,N_9708,N_8028);
and U10589 (N_10589,N_8914,N_6596);
or U10590 (N_10590,N_9761,N_7686);
nand U10591 (N_10591,N_8414,N_9469);
nor U10592 (N_10592,N_9558,N_5512);
xnor U10593 (N_10593,N_9906,N_5550);
or U10594 (N_10594,N_5310,N_6677);
nand U10595 (N_10595,N_5899,N_9476);
xnor U10596 (N_10596,N_7974,N_5884);
nand U10597 (N_10597,N_7747,N_7639);
and U10598 (N_10598,N_6569,N_8615);
and U10599 (N_10599,N_7670,N_5752);
nand U10600 (N_10600,N_9738,N_8642);
nor U10601 (N_10601,N_5779,N_5450);
xor U10602 (N_10602,N_6231,N_9843);
or U10603 (N_10603,N_8443,N_7347);
nor U10604 (N_10604,N_9391,N_7971);
and U10605 (N_10605,N_5012,N_5964);
xnor U10606 (N_10606,N_9909,N_9913);
and U10607 (N_10607,N_6644,N_5375);
nand U10608 (N_10608,N_5300,N_5118);
xnor U10609 (N_10609,N_6827,N_5707);
or U10610 (N_10610,N_7506,N_9918);
xnor U10611 (N_10611,N_5382,N_7171);
xor U10612 (N_10612,N_6744,N_5257);
or U10613 (N_10613,N_8086,N_7587);
or U10614 (N_10614,N_6752,N_8449);
nor U10615 (N_10615,N_8138,N_7381);
xnor U10616 (N_10616,N_6169,N_5953);
and U10617 (N_10617,N_6237,N_8186);
and U10618 (N_10618,N_5814,N_6964);
xor U10619 (N_10619,N_7898,N_9775);
and U10620 (N_10620,N_6927,N_7805);
and U10621 (N_10621,N_5409,N_9439);
and U10622 (N_10622,N_9621,N_9114);
xor U10623 (N_10623,N_8892,N_5395);
nand U10624 (N_10624,N_5358,N_5802);
nand U10625 (N_10625,N_9872,N_6158);
xor U10626 (N_10626,N_9473,N_5232);
and U10627 (N_10627,N_5760,N_7495);
xor U10628 (N_10628,N_8045,N_7677);
and U10629 (N_10629,N_7497,N_5432);
nor U10630 (N_10630,N_5429,N_5433);
and U10631 (N_10631,N_7428,N_7572);
nor U10632 (N_10632,N_5249,N_9634);
nand U10633 (N_10633,N_8216,N_8353);
nor U10634 (N_10634,N_5679,N_7880);
xor U10635 (N_10635,N_7727,N_5369);
nor U10636 (N_10636,N_6911,N_8993);
or U10637 (N_10637,N_8725,N_5015);
xor U10638 (N_10638,N_5248,N_6050);
xnor U10639 (N_10639,N_8198,N_6601);
xnor U10640 (N_10640,N_7720,N_8714);
xnor U10641 (N_10641,N_8891,N_8202);
nand U10642 (N_10642,N_9585,N_5841);
nand U10643 (N_10643,N_9883,N_7234);
nor U10644 (N_10644,N_5171,N_7500);
or U10645 (N_10645,N_6249,N_9841);
xnor U10646 (N_10646,N_5917,N_7668);
and U10647 (N_10647,N_5889,N_5921);
and U10648 (N_10648,N_8470,N_6980);
or U10649 (N_10649,N_6085,N_5954);
nor U10650 (N_10650,N_9105,N_9795);
xnor U10651 (N_10651,N_9249,N_8939);
nor U10652 (N_10652,N_7855,N_9868);
xor U10653 (N_10653,N_6461,N_5795);
and U10654 (N_10654,N_7229,N_9636);
or U10655 (N_10655,N_9474,N_5968);
or U10656 (N_10656,N_7829,N_9483);
nand U10657 (N_10657,N_7714,N_5002);
xor U10658 (N_10658,N_8078,N_6176);
or U10659 (N_10659,N_6281,N_5370);
nor U10660 (N_10660,N_5925,N_8753);
nor U10661 (N_10661,N_8380,N_6845);
or U10662 (N_10662,N_6161,N_9168);
and U10663 (N_10663,N_9496,N_6648);
xor U10664 (N_10664,N_5830,N_9830);
nand U10665 (N_10665,N_6659,N_5676);
nor U10666 (N_10666,N_8674,N_7475);
nand U10667 (N_10667,N_9154,N_6318);
or U10668 (N_10668,N_8995,N_9966);
and U10669 (N_10669,N_8427,N_7618);
or U10670 (N_10670,N_5645,N_5129);
and U10671 (N_10671,N_9529,N_7785);
xor U10672 (N_10672,N_9288,N_7650);
and U10673 (N_10673,N_7087,N_5905);
or U10674 (N_10674,N_8007,N_9527);
xnor U10675 (N_10675,N_5670,N_9849);
xor U10676 (N_10676,N_6464,N_8592);
or U10677 (N_10677,N_8341,N_6217);
and U10678 (N_10678,N_6692,N_5799);
nor U10679 (N_10679,N_9485,N_7708);
nand U10680 (N_10680,N_8265,N_8768);
xnor U10681 (N_10681,N_6266,N_9426);
nand U10682 (N_10682,N_8273,N_9037);
and U10683 (N_10683,N_9947,N_9845);
or U10684 (N_10684,N_6211,N_7745);
nor U10685 (N_10685,N_9825,N_5183);
and U10686 (N_10686,N_6696,N_5092);
xnor U10687 (N_10687,N_6102,N_6943);
or U10688 (N_10688,N_7505,N_9182);
and U10689 (N_10689,N_6652,N_8290);
xor U10690 (N_10690,N_7946,N_6733);
and U10691 (N_10691,N_9318,N_8336);
and U10692 (N_10692,N_8382,N_9295);
xor U10693 (N_10693,N_5080,N_7259);
nand U10694 (N_10694,N_7013,N_5138);
nor U10695 (N_10695,N_5856,N_7374);
nor U10696 (N_10696,N_5757,N_6611);
and U10697 (N_10697,N_7871,N_6414);
or U10698 (N_10698,N_7678,N_5308);
nor U10699 (N_10699,N_7755,N_8576);
nor U10700 (N_10700,N_8718,N_9586);
or U10701 (N_10701,N_9314,N_8619);
and U10702 (N_10702,N_5388,N_8450);
xor U10703 (N_10703,N_9059,N_9492);
nor U10704 (N_10704,N_8711,N_8693);
nand U10705 (N_10705,N_8472,N_7943);
xor U10706 (N_10706,N_5235,N_7312);
or U10707 (N_10707,N_9544,N_9869);
or U10708 (N_10708,N_5365,N_5425);
and U10709 (N_10709,N_9299,N_5705);
nor U10710 (N_10710,N_7681,N_6484);
xnor U10711 (N_10711,N_7725,N_5282);
xor U10712 (N_10712,N_9565,N_7112);
xor U10713 (N_10713,N_5397,N_9917);
nor U10714 (N_10714,N_7684,N_6932);
nand U10715 (N_10715,N_9366,N_7046);
nand U10716 (N_10716,N_9949,N_9413);
nand U10717 (N_10717,N_6639,N_5244);
nand U10718 (N_10718,N_8070,N_9017);
and U10719 (N_10719,N_6565,N_5175);
or U10720 (N_10720,N_7166,N_5453);
xor U10721 (N_10721,N_9128,N_9127);
or U10722 (N_10722,N_5824,N_6116);
nand U10723 (N_10723,N_9960,N_8952);
and U10724 (N_10724,N_6844,N_6227);
xnor U10725 (N_10725,N_9945,N_8763);
nand U10726 (N_10726,N_5990,N_6801);
or U10727 (N_10727,N_6581,N_6793);
nor U10728 (N_10728,N_6811,N_5941);
or U10729 (N_10729,N_6933,N_6399);
and U10730 (N_10730,N_8841,N_6000);
nand U10731 (N_10731,N_6602,N_8461);
xor U10732 (N_10732,N_5786,N_6542);
nor U10733 (N_10733,N_9322,N_8349);
nand U10734 (N_10734,N_9614,N_8408);
xor U10735 (N_10735,N_8780,N_8284);
and U10736 (N_10736,N_9863,N_6682);
nor U10737 (N_10737,N_5770,N_6264);
nand U10738 (N_10738,N_5314,N_5058);
nor U10739 (N_10739,N_8625,N_8313);
or U10740 (N_10740,N_8754,N_5504);
nor U10741 (N_10741,N_6889,N_5636);
nand U10742 (N_10742,N_6118,N_6245);
or U10743 (N_10743,N_6993,N_9324);
or U10744 (N_10744,N_9921,N_6056);
nand U10745 (N_10745,N_7246,N_6832);
nor U10746 (N_10746,N_6704,N_9548);
or U10747 (N_10747,N_7733,N_6476);
and U10748 (N_10748,N_5095,N_8463);
xnor U10749 (N_10749,N_9542,N_7532);
xor U10750 (N_10750,N_8587,N_5044);
or U10751 (N_10751,N_5471,N_8422);
or U10752 (N_10752,N_7966,N_9743);
nor U10753 (N_10753,N_9498,N_9383);
xor U10754 (N_10754,N_8635,N_9537);
and U10755 (N_10755,N_9040,N_8301);
or U10756 (N_10756,N_7926,N_7884);
and U10757 (N_10757,N_9790,N_6311);
or U10758 (N_10758,N_7422,N_6897);
and U10759 (N_10759,N_9902,N_8921);
and U10760 (N_10760,N_9608,N_8491);
xnor U10761 (N_10761,N_9022,N_6437);
or U10762 (N_10762,N_5483,N_8988);
or U10763 (N_10763,N_7243,N_9778);
nor U10764 (N_10764,N_9039,N_7209);
nand U10765 (N_10765,N_9670,N_8579);
nand U10766 (N_10766,N_9980,N_6477);
and U10767 (N_10767,N_8524,N_6415);
nor U10768 (N_10768,N_6133,N_5446);
xnor U10769 (N_10769,N_8240,N_7944);
or U10770 (N_10770,N_8101,N_8288);
or U10771 (N_10771,N_8673,N_7594);
and U10772 (N_10772,N_5423,N_7850);
and U10773 (N_10773,N_8540,N_6841);
nand U10774 (N_10774,N_7425,N_7181);
and U10775 (N_10775,N_8859,N_5748);
nand U10776 (N_10776,N_6526,N_7280);
xnor U10777 (N_10777,N_8781,N_8306);
nand U10778 (N_10778,N_6656,N_8830);
or U10779 (N_10779,N_8221,N_5000);
nand U10780 (N_10780,N_7891,N_6054);
xor U10781 (N_10781,N_6339,N_6626);
xor U10782 (N_10782,N_5460,N_8513);
and U10783 (N_10783,N_8071,N_9612);
or U10784 (N_10784,N_7395,N_5697);
nor U10785 (N_10785,N_6926,N_7511);
nand U10786 (N_10786,N_9256,N_5131);
nand U10787 (N_10787,N_7489,N_9525);
or U10788 (N_10788,N_6673,N_6689);
nand U10789 (N_10789,N_6215,N_7145);
nor U10790 (N_10790,N_7903,N_7419);
and U10791 (N_10791,N_9997,N_8694);
or U10792 (N_10792,N_9916,N_8626);
xnor U10793 (N_10793,N_5750,N_9173);
or U10794 (N_10794,N_7396,N_6088);
or U10795 (N_10795,N_7090,N_7608);
and U10796 (N_10796,N_6313,N_6705);
nor U10797 (N_10797,N_5986,N_8580);
nand U10798 (N_10798,N_7649,N_7619);
and U10799 (N_10799,N_6929,N_5746);
nor U10800 (N_10800,N_7833,N_7003);
or U10801 (N_10801,N_9086,N_6725);
or U10802 (N_10802,N_6937,N_6029);
or U10803 (N_10803,N_7457,N_6090);
or U10804 (N_10804,N_6651,N_6746);
or U10805 (N_10805,N_9700,N_8833);
nand U10806 (N_10806,N_5916,N_6092);
or U10807 (N_10807,N_6315,N_9604);
nand U10808 (N_10808,N_9104,N_9157);
nor U10809 (N_10809,N_7394,N_6579);
nand U10810 (N_10810,N_8715,N_9227);
nor U10811 (N_10811,N_9223,N_7125);
and U10812 (N_10812,N_6205,N_6110);
and U10813 (N_10813,N_6768,N_6069);
and U10814 (N_10814,N_8431,N_9332);
and U10815 (N_10815,N_7841,N_9671);
or U10816 (N_10816,N_7576,N_5218);
or U10817 (N_10817,N_9888,N_9629);
xnor U10818 (N_10818,N_6972,N_9201);
and U10819 (N_10819,N_8888,N_9854);
nor U10820 (N_10820,N_8137,N_8161);
nand U10821 (N_10821,N_8772,N_8766);
nor U10822 (N_10822,N_8621,N_9246);
and U10823 (N_10823,N_8541,N_7680);
or U10824 (N_10824,N_5371,N_5669);
or U10825 (N_10825,N_8904,N_9745);
or U10826 (N_10826,N_7554,N_8704);
or U10827 (N_10827,N_6400,N_5042);
and U10828 (N_10828,N_7058,N_8658);
nor U10829 (N_10829,N_9970,N_6847);
and U10830 (N_10830,N_7586,N_7403);
nor U10831 (N_10831,N_7908,N_8054);
or U10832 (N_10832,N_7272,N_5588);
and U10833 (N_10833,N_5346,N_7238);
xor U10834 (N_10834,N_9573,N_5847);
nand U10835 (N_10835,N_5589,N_8435);
nand U10836 (N_10836,N_8951,N_5680);
nand U10837 (N_10837,N_5335,N_9603);
nand U10838 (N_10838,N_7982,N_5793);
or U10839 (N_10839,N_5043,N_8527);
nor U10840 (N_10840,N_6055,N_7464);
and U10841 (N_10841,N_7826,N_6327);
nor U10842 (N_10842,N_8756,N_6781);
or U10843 (N_10843,N_7227,N_5486);
nand U10844 (N_10844,N_7199,N_6930);
and U10845 (N_10845,N_9735,N_7275);
or U10846 (N_10846,N_8945,N_8667);
or U10847 (N_10847,N_5491,N_8319);
and U10848 (N_10848,N_9986,N_9014);
nor U10849 (N_10849,N_8767,N_6635);
nand U10850 (N_10850,N_6173,N_8147);
nor U10851 (N_10851,N_6753,N_7251);
or U10852 (N_10852,N_5267,N_5318);
or U10853 (N_10853,N_9823,N_5724);
nor U10854 (N_10854,N_7219,N_9265);
nor U10855 (N_10855,N_5500,N_7148);
nand U10856 (N_10856,N_7055,N_8304);
or U10857 (N_10857,N_5114,N_8960);
or U10858 (N_10858,N_6357,N_8321);
nand U10859 (N_10859,N_8594,N_7099);
and U10860 (N_10860,N_5156,N_7141);
xnor U10861 (N_10861,N_6621,N_5288);
xnor U10862 (N_10862,N_9674,N_7067);
and U10863 (N_10863,N_7339,N_6119);
nand U10864 (N_10864,N_5277,N_8662);
or U10865 (N_10865,N_7366,N_5758);
nor U10866 (N_10866,N_6140,N_5584);
and U10867 (N_10867,N_5741,N_9749);
nand U10868 (N_10868,N_9704,N_5321);
xnor U10869 (N_10869,N_7237,N_9381);
nor U10870 (N_10870,N_5803,N_6861);
xnor U10871 (N_10871,N_6994,N_5113);
xnor U10872 (N_10872,N_9834,N_6757);
or U10873 (N_10873,N_9160,N_7144);
nand U10874 (N_10874,N_6663,N_7274);
nor U10875 (N_10875,N_7977,N_5715);
xnor U10876 (N_10876,N_9169,N_8980);
xnor U10877 (N_10877,N_9789,N_6442);
or U10878 (N_10878,N_8843,N_8103);
nand U10879 (N_10879,N_7332,N_9297);
and U10880 (N_10880,N_9307,N_8910);
and U10881 (N_10881,N_7648,N_7449);
xor U10882 (N_10882,N_9132,N_8553);
or U10883 (N_10883,N_8755,N_8428);
or U10884 (N_10884,N_8985,N_8957);
or U10885 (N_10885,N_9194,N_7947);
nor U10886 (N_10886,N_5116,N_7054);
or U10887 (N_10887,N_6519,N_8080);
or U10888 (N_10888,N_6267,N_8590);
nand U10889 (N_10889,N_5829,N_5983);
and U10890 (N_10890,N_8133,N_9499);
and U10891 (N_10891,N_8002,N_5516);
and U10892 (N_10892,N_8972,N_6506);
or U10893 (N_10893,N_5864,N_8244);
or U10894 (N_10894,N_9734,N_6711);
or U10895 (N_10895,N_9176,N_7118);
or U10896 (N_10896,N_8577,N_9136);
or U10897 (N_10897,N_7045,N_9400);
xor U10898 (N_10898,N_8219,N_8365);
or U10899 (N_10899,N_8536,N_6123);
xor U10900 (N_10900,N_5238,N_7671);
or U10901 (N_10901,N_9262,N_9056);
nand U10902 (N_10902,N_9533,N_8801);
nor U10903 (N_10903,N_8128,N_8091);
and U10904 (N_10904,N_9551,N_6352);
nand U10905 (N_10905,N_7986,N_9046);
nor U10906 (N_10906,N_8591,N_5506);
nor U10907 (N_10907,N_5867,N_5591);
or U10908 (N_10908,N_9717,N_9339);
xor U10909 (N_10909,N_9319,N_8531);
xor U10910 (N_10910,N_5602,N_9325);
xor U10911 (N_10911,N_8686,N_9836);
xnor U10912 (N_10912,N_6240,N_9073);
and U10913 (N_10913,N_8499,N_9260);
nand U10914 (N_10914,N_7557,N_9101);
nand U10915 (N_10915,N_9859,N_7409);
nand U10916 (N_10916,N_5245,N_7911);
nor U10917 (N_10917,N_9231,N_6485);
nand U10918 (N_10918,N_6320,N_8242);
nand U10919 (N_10919,N_6571,N_6545);
xnor U10920 (N_10920,N_6081,N_6873);
xor U10921 (N_10921,N_5437,N_8190);
and U10922 (N_10922,N_5903,N_9427);
nor U10923 (N_10923,N_7525,N_8157);
xor U10924 (N_10924,N_5207,N_5457);
and U10925 (N_10925,N_6960,N_5162);
xor U10926 (N_10926,N_9372,N_6722);
nand U10927 (N_10927,N_5184,N_5228);
nand U10928 (N_10928,N_9599,N_7134);
nor U10929 (N_10929,N_9067,N_5538);
xor U10930 (N_10930,N_6931,N_9495);
or U10931 (N_10931,N_8933,N_7912);
and U10932 (N_10932,N_8507,N_7673);
or U10933 (N_10933,N_9852,N_5488);
nor U10934 (N_10934,N_6360,N_9939);
xor U10935 (N_10935,N_8882,N_6006);
nand U10936 (N_10936,N_8834,N_8168);
and U10937 (N_10937,N_8911,N_7517);
xor U10938 (N_10938,N_9727,N_5489);
nand U10939 (N_10939,N_8890,N_5339);
nor U10940 (N_10940,N_9653,N_6741);
or U10941 (N_10941,N_5319,N_8665);
nand U10942 (N_10942,N_5157,N_8311);
xnor U10943 (N_10943,N_8338,N_9139);
xnor U10944 (N_10944,N_6138,N_7719);
and U10945 (N_10945,N_9592,N_5568);
or U10946 (N_10946,N_6046,N_5507);
nand U10947 (N_10947,N_6201,N_8400);
and U10948 (N_10948,N_5927,N_9787);
nand U10949 (N_10949,N_7083,N_6351);
nand U10950 (N_10950,N_6906,N_5561);
and U10951 (N_10951,N_9416,N_5819);
nand U10952 (N_10952,N_7380,N_8481);
nor U10953 (N_10953,N_7849,N_6346);
nand U10954 (N_10954,N_9358,N_5394);
and U10955 (N_10955,N_6361,N_7994);
nand U10956 (N_10956,N_5992,N_5274);
or U10957 (N_10957,N_8060,N_6077);
and U10958 (N_10958,N_9087,N_6193);
nand U10959 (N_10959,N_7252,N_8254);
nor U10960 (N_10960,N_8774,N_6670);
xnor U10961 (N_10961,N_8657,N_7154);
nand U10962 (N_10962,N_5711,N_9215);
and U10963 (N_10963,N_7330,N_5237);
xnor U10964 (N_10964,N_9922,N_5284);
or U10965 (N_10965,N_6979,N_9150);
or U10966 (N_10966,N_8630,N_5571);
and U10967 (N_10967,N_8691,N_7551);
nand U10968 (N_10968,N_9134,N_9919);
and U10969 (N_10969,N_7451,N_6720);
nor U10970 (N_10970,N_5839,N_8857);
xnor U10971 (N_10971,N_5835,N_8377);
nor U10972 (N_10972,N_8955,N_6568);
xor U10973 (N_10973,N_8624,N_6063);
and U10974 (N_10974,N_9365,N_5607);
or U10975 (N_10975,N_7257,N_6275);
xor U10976 (N_10976,N_9929,N_5465);
nor U10977 (N_10977,N_9214,N_9458);
nor U10978 (N_10978,N_5402,N_7993);
xor U10979 (N_10979,N_5451,N_8728);
and U10980 (N_10980,N_6608,N_7071);
nor U10981 (N_10981,N_6719,N_7808);
xnor U10982 (N_10982,N_7172,N_8256);
nand U10983 (N_10983,N_5970,N_5778);
or U10984 (N_10984,N_6162,N_6496);
xor U10985 (N_10985,N_9777,N_6799);
nand U10986 (N_10986,N_7807,N_6358);
xnor U10987 (N_10987,N_7044,N_7352);
nand U10988 (N_10988,N_5570,N_6623);
or U10989 (N_10989,N_5578,N_9216);
and U10990 (N_10990,N_6578,N_9363);
or U10991 (N_10991,N_6007,N_5374);
nand U10992 (N_10992,N_8281,N_9757);
or U10993 (N_10993,N_6216,N_9532);
nor U10994 (N_10994,N_6776,N_5511);
nor U10995 (N_10995,N_5452,N_6627);
xnor U10996 (N_10996,N_6002,N_9343);
nor U10997 (N_10997,N_5412,N_5126);
and U10998 (N_10998,N_7738,N_5045);
nor U10999 (N_10999,N_7163,N_9632);
and U11000 (N_11000,N_7386,N_8631);
or U11001 (N_11001,N_7410,N_9093);
nor U11002 (N_11002,N_6309,N_7498);
nand U11003 (N_11003,N_9623,N_8858);
nand U11004 (N_11004,N_7717,N_5503);
xnor U11005 (N_11005,N_5624,N_7245);
nor U11006 (N_11006,N_6153,N_7710);
nor U11007 (N_11007,N_7922,N_6712);
nor U11008 (N_11008,N_8312,N_8879);
nor U11009 (N_11009,N_9606,N_5061);
nand U11010 (N_11010,N_5347,N_8308);
nand U11011 (N_11011,N_9403,N_7302);
nand U11012 (N_11012,N_6534,N_9025);
xor U11013 (N_11013,N_7548,N_9163);
nand U11014 (N_11014,N_7902,N_8026);
nand U11015 (N_11015,N_6427,N_7526);
nor U11016 (N_11016,N_8959,N_7504);
nand U11017 (N_11017,N_9526,N_9977);
xnor U11018 (N_11018,N_7376,N_5147);
nand U11019 (N_11019,N_6560,N_6383);
nand U11020 (N_11020,N_5047,N_7020);
and U11021 (N_11021,N_6546,N_5868);
nor U11022 (N_11022,N_9418,N_6074);
and U11023 (N_11023,N_9417,N_5031);
xor U11024 (N_11024,N_5299,N_6364);
xor U11025 (N_11025,N_5716,N_8181);
nand U11026 (N_11026,N_9278,N_5734);
or U11027 (N_11027,N_6797,N_9865);
nand U11028 (N_11028,N_5845,N_8818);
and U11029 (N_11029,N_9052,N_9813);
nand U11030 (N_11030,N_7432,N_6241);
or U11031 (N_11031,N_7861,N_6170);
xor U11032 (N_11032,N_9751,N_5351);
nand U11033 (N_11033,N_7512,N_5439);
or U11034 (N_11034,N_9192,N_8999);
nor U11035 (N_11035,N_7948,N_8997);
nor U11036 (N_11036,N_8681,N_8039);
or U11037 (N_11037,N_9348,N_7185);
and U11038 (N_11038,N_6040,N_5494);
or U11039 (N_11039,N_7137,N_8131);
or U11040 (N_11040,N_6812,N_9760);
xnor U11041 (N_11041,N_9335,N_9971);
and U11042 (N_11042,N_9074,N_8706);
xor U11043 (N_11043,N_8578,N_8385);
and U11044 (N_11044,N_6742,N_5192);
nor U11045 (N_11045,N_5014,N_5605);
nand U11046 (N_11046,N_9344,N_6335);
or U11047 (N_11047,N_6229,N_5399);
xnor U11048 (N_11048,N_6502,N_8741);
or U11049 (N_11049,N_6588,N_8467);
or U11050 (N_11050,N_8647,N_6834);
nor U11051 (N_11051,N_7723,N_6458);
xnor U11052 (N_11052,N_8515,N_7375);
xnor U11053 (N_11053,N_5885,N_6107);
or U11054 (N_11054,N_8895,N_9600);
or U11055 (N_11055,N_6879,N_5648);
nor U11056 (N_11056,N_7856,N_5709);
or U11057 (N_11057,N_9648,N_8670);
and U11058 (N_11058,N_5161,N_9012);
xnor U11059 (N_11059,N_8723,N_5573);
xor U11060 (N_11060,N_9875,N_5774);
xor U11061 (N_11061,N_5051,N_5474);
nand U11062 (N_11062,N_9268,N_9506);
and U11063 (N_11063,N_5208,N_8584);
and U11064 (N_11064,N_9261,N_7413);
nor U11065 (N_11065,N_7306,N_7640);
xor U11066 (N_11066,N_5415,N_9024);
xnor U11067 (N_11067,N_6031,N_5266);
and U11068 (N_11068,N_7836,N_5876);
xor U11069 (N_11069,N_6410,N_7155);
nand U11070 (N_11070,N_6853,N_5316);
xnor U11071 (N_11071,N_8687,N_6424);
and U11072 (N_11072,N_5010,N_6858);
and U11073 (N_11073,N_5136,N_5018);
nand U11074 (N_11074,N_6392,N_9005);
xor U11075 (N_11075,N_5492,N_6959);
and U11076 (N_11076,N_6538,N_9555);
nor U11077 (N_11077,N_5210,N_5634);
or U11078 (N_11078,N_6788,N_9258);
xor U11079 (N_11079,N_7291,N_7091);
nand U11080 (N_11080,N_7405,N_9824);
nand U11081 (N_11081,N_9422,N_5477);
nand U11082 (N_11082,N_6634,N_8250);
or U11083 (N_11083,N_5197,N_7779);
nand U11084 (N_11084,N_6871,N_6058);
nor U11085 (N_11085,N_5124,N_6935);
nand U11086 (N_11086,N_6968,N_9306);
and U11087 (N_11087,N_6418,N_8838);
and U11088 (N_11088,N_9076,N_7981);
and U11089 (N_11089,N_7585,N_9669);
or U11090 (N_11090,N_7685,N_6343);
or U11091 (N_11091,N_8632,N_9447);
and U11092 (N_11092,N_8769,N_9508);
or U11093 (N_11093,N_7351,N_8478);
or U11094 (N_11094,N_5247,N_5191);
nand U11095 (N_11095,N_9645,N_7627);
or U11096 (N_11096,N_6342,N_7909);
or U11097 (N_11097,N_7271,N_9805);
or U11098 (N_11098,N_6769,N_5200);
xor U11099 (N_11099,N_6300,N_8212);
xnor U11100 (N_11100,N_9656,N_9833);
or U11101 (N_11101,N_9266,N_9864);
and U11102 (N_11102,N_8575,N_5269);
nand U11103 (N_11103,N_7078,N_9428);
and U11104 (N_11104,N_7461,N_5853);
nand U11105 (N_11105,N_7590,N_6482);
or U11106 (N_11106,N_7228,N_8271);
or U11107 (N_11107,N_5344,N_8749);
nand U11108 (N_11108,N_9368,N_5360);
nor U11109 (N_11109,N_8352,N_5600);
nand U11110 (N_11110,N_7265,N_7008);
xnor U11111 (N_11111,N_9185,N_6026);
nor U11112 (N_11112,N_8424,N_7041);
nand U11113 (N_11113,N_7104,N_6604);
nor U11114 (N_11114,N_9948,N_9133);
nor U11115 (N_11115,N_8855,N_9057);
and U11116 (N_11116,N_8085,N_5664);
nor U11117 (N_11117,N_5638,N_6921);
xnor U11118 (N_11118,N_7839,N_6062);
nor U11119 (N_11119,N_5408,N_9296);
xor U11120 (N_11120,N_9943,N_8521);
and U11121 (N_11121,N_9092,N_7831);
nor U11122 (N_11122,N_5958,N_5001);
nand U11123 (N_11123,N_7233,N_7604);
or U11124 (N_11124,N_9584,N_9251);
nand U11125 (N_11125,N_6232,N_9556);
nand U11126 (N_11126,N_5343,N_8067);
nand U11127 (N_11127,N_7823,N_5691);
nand U11128 (N_11128,N_5924,N_6945);
nand U11129 (N_11129,N_9294,N_8778);
nor U11130 (N_11130,N_9196,N_7202);
and U11131 (N_11131,N_5276,N_9932);
xor U11132 (N_11132,N_6726,N_6676);
and U11133 (N_11133,N_9250,N_7406);
or U11134 (N_11134,N_6890,N_5271);
nand U11135 (N_11135,N_9376,N_7803);
nor U11136 (N_11136,N_7932,N_5226);
or U11137 (N_11137,N_5762,N_5005);
nor U11138 (N_11138,N_6014,N_6548);
and U11139 (N_11139,N_6291,N_7389);
or U11140 (N_11140,N_5463,N_9858);
or U11141 (N_11141,N_9677,N_8656);
nand U11142 (N_11142,N_6992,N_7992);
xnor U11143 (N_11143,N_8208,N_9587);
and U11144 (N_11144,N_8929,N_9903);
nor U11145 (N_11145,N_8274,N_5049);
xnor U11146 (N_11146,N_9687,N_9545);
nor U11147 (N_11147,N_8005,N_9159);
nor U11148 (N_11148,N_7528,N_9688);
or U11149 (N_11149,N_7061,N_8107);
nand U11150 (N_11150,N_7515,N_8930);
xnor U11151 (N_11151,N_7438,N_9739);
nand U11152 (N_11152,N_6976,N_9315);
nor U11153 (N_11153,N_9607,N_8146);
xor U11154 (N_11154,N_5656,N_5513);
nor U11155 (N_11155,N_5211,N_8548);
and U11156 (N_11156,N_6740,N_7927);
nand U11157 (N_11157,N_7283,N_6329);
nor U11158 (N_11158,N_9484,N_6146);
nor U11159 (N_11159,N_6257,N_6949);
or U11160 (N_11160,N_8844,N_9006);
and U11161 (N_11161,N_8065,N_6638);
xor U11162 (N_11162,N_7675,N_9773);
and U11163 (N_11163,N_8777,N_5164);
nand U11164 (N_11164,N_9853,N_8438);
xor U11165 (N_11165,N_5540,N_9702);
and U11166 (N_11166,N_7742,N_9117);
nor U11167 (N_11167,N_8432,N_5046);
nor U11168 (N_11168,N_7817,N_5567);
and U11169 (N_11169,N_7535,N_7182);
xnor U11170 (N_11170,N_7445,N_8629);
xor U11171 (N_11171,N_7208,N_7600);
xor U11172 (N_11172,N_8452,N_9616);
and U11173 (N_11173,N_5100,N_6550);
or U11174 (N_11174,N_8925,N_8747);
xor U11175 (N_11175,N_9061,N_6378);
nand U11176 (N_11176,N_8609,N_6171);
or U11177 (N_11177,N_7715,N_7488);
and U11178 (N_11178,N_9138,N_7480);
and U11179 (N_11179,N_6207,N_6732);
nand U11180 (N_11180,N_5466,N_8602);
or U11181 (N_11181,N_6767,N_8850);
and U11182 (N_11182,N_7799,N_8314);
nor U11183 (N_11183,N_8998,N_9471);
and U11184 (N_11184,N_6701,N_6471);
nand U11185 (N_11185,N_5108,N_9627);
nor U11186 (N_11186,N_9598,N_6446);
and U11187 (N_11187,N_8840,N_7285);
or U11188 (N_11188,N_7760,N_9211);
xor U11189 (N_11189,N_9631,N_6179);
or U11190 (N_11190,N_5362,N_7603);
or U11191 (N_11191,N_7157,N_9450);
and U11192 (N_11192,N_5763,N_8023);
nand U11193 (N_11193,N_7204,N_6180);
xnor U11194 (N_11194,N_7494,N_9406);
or U11195 (N_11195,N_6198,N_9810);
xnor U11196 (N_11196,N_9594,N_6134);
and U11197 (N_11197,N_5193,N_7429);
nand U11198 (N_11198,N_9676,N_6256);
nor U11199 (N_11199,N_9937,N_5761);
nand U11200 (N_11200,N_8106,N_7156);
and U11201 (N_11201,N_8861,N_5576);
and U11202 (N_11202,N_7496,N_7527);
xor U11203 (N_11203,N_8986,N_8224);
or U11204 (N_11204,N_6436,N_7646);
nor U11205 (N_11205,N_7697,N_7750);
xor U11206 (N_11206,N_5844,N_6938);
xor U11207 (N_11207,N_8528,N_7319);
and U11208 (N_11208,N_9070,N_7797);
xor U11209 (N_11209,N_5079,N_9666);
xor U11210 (N_11210,N_5972,N_9423);
nor U11211 (N_11211,N_6637,N_9679);
nor U11212 (N_11212,N_7292,N_9582);
and U11213 (N_11213,N_9050,N_8978);
and U11214 (N_11214,N_9619,N_8831);
and U11215 (N_11215,N_8345,N_5127);
nand U11216 (N_11216,N_8616,N_6802);
xnor U11217 (N_11217,N_7165,N_8409);
xnor U11218 (N_11218,N_8690,N_9367);
xor U11219 (N_11219,N_5445,N_8073);
or U11220 (N_11220,N_7959,N_5454);
nor U11221 (N_11221,N_8484,N_5270);
and U11222 (N_11222,N_8569,N_7258);
and U11223 (N_11223,N_5661,N_5564);
nor U11224 (N_11224,N_8050,N_5777);
and U11225 (N_11225,N_5029,N_7810);
and U11226 (N_11226,N_5982,N_7062);
nand U11227 (N_11227,N_9641,N_8519);
nor U11228 (N_11228,N_9723,N_8165);
nand U11229 (N_11229,N_7301,N_9047);
nor U11230 (N_11230,N_5337,N_5674);
nand U11231 (N_11231,N_8079,N_6120);
or U11232 (N_11232,N_8490,N_7398);
or U11233 (N_11233,N_5221,N_7631);
nor U11234 (N_11234,N_5392,N_7956);
or U11235 (N_11235,N_7542,N_8886);
and U11236 (N_11236,N_5952,N_7085);
nor U11237 (N_11237,N_9481,N_6563);
xnor U11238 (N_11238,N_6272,N_7852);
or U11239 (N_11239,N_7962,N_5801);
nand U11240 (N_11240,N_5229,N_7421);
and U11241 (N_11241,N_5289,N_5170);
nand U11242 (N_11242,N_8143,N_9993);
or U11243 (N_11243,N_6104,N_9857);
or U11244 (N_11244,N_5254,N_7070);
nor U11245 (N_11245,N_5083,N_5794);
nor U11246 (N_11246,N_6293,N_5273);
nand U11247 (N_11247,N_7068,N_7973);
xnor U11248 (N_11248,N_6738,N_8182);
nand U11249 (N_11249,N_9737,N_6559);
nor U11250 (N_11250,N_6044,N_7373);
xnor U11251 (N_11251,N_6504,N_6254);
or U11252 (N_11252,N_6973,N_8974);
and U11253 (N_11253,N_7244,N_9284);
xnor U11254 (N_11254,N_8464,N_9725);
and U11255 (N_11255,N_9197,N_5174);
or U11256 (N_11256,N_5385,N_8573);
nor U11257 (N_11257,N_9541,N_9374);
nor U11258 (N_11258,N_7626,N_9111);
nor U11259 (N_11259,N_7739,N_9472);
and U11260 (N_11260,N_5974,N_7411);
xor U11261 (N_11261,N_7756,N_7060);
nand U11262 (N_11262,N_9985,N_5878);
and U11263 (N_11263,N_7814,N_6421);
nor U11264 (N_11264,N_5587,N_7983);
nand U11265 (N_11265,N_6277,N_6956);
nand U11266 (N_11266,N_5725,N_8444);
and U11267 (N_11267,N_5866,N_9007);
or U11268 (N_11268,N_7088,N_6368);
nor U11269 (N_11269,N_9771,N_7315);
xor U11270 (N_11270,N_7970,N_9907);
or U11271 (N_11271,N_7705,N_5775);
nor U11272 (N_11272,N_9732,N_5062);
or U11273 (N_11273,N_7116,N_9782);
and U11274 (N_11274,N_8021,N_5718);
or U11275 (N_11275,N_7564,N_9815);
or U11276 (N_11276,N_8660,N_8611);
or U11277 (N_11277,N_8794,N_8742);
xor U11278 (N_11278,N_8501,N_7169);
xnor U11279 (N_11279,N_9796,N_9539);
nand U11280 (N_11280,N_8726,N_5977);
and U11281 (N_11281,N_6669,N_9089);
xnor U11282 (N_11282,N_6615,N_6394);
nor U11283 (N_11283,N_9456,N_5111);
nor U11284 (N_11284,N_8503,N_7632);
and U11285 (N_11285,N_7919,N_6132);
nand U11286 (N_11286,N_7335,N_7888);
and U11287 (N_11287,N_9682,N_9800);
nor U11288 (N_11288,N_9802,N_8418);
nor U11289 (N_11289,N_6505,N_6270);
nand U11290 (N_11290,N_5653,N_5132);
nand U11291 (N_11291,N_9311,N_8607);
nor U11292 (N_11292,N_7881,N_9938);
or U11293 (N_11293,N_7991,N_5497);
nor U11294 (N_11294,N_9191,N_9331);
and U11295 (N_11295,N_7768,N_8518);
nand U11296 (N_11296,N_6970,N_7945);
xnor U11297 (N_11297,N_9102,N_7674);
and U11298 (N_11298,N_6771,N_9031);
xor U11299 (N_11299,N_7207,N_9255);
and U11300 (N_11300,N_8122,N_8539);
nand U11301 (N_11301,N_7877,N_8344);
or U11302 (N_11302,N_7160,N_9455);
and U11303 (N_11303,N_5614,N_5303);
and U11304 (N_11304,N_5223,N_6167);
or U11305 (N_11305,N_9522,N_9766);
nor U11306 (N_11306,N_8451,N_9814);
xnor U11307 (N_11307,N_8401,N_5509);
nor U11308 (N_11308,N_5259,N_6387);
xor U11309 (N_11309,N_7299,N_7195);
nor U11310 (N_11310,N_6248,N_7365);
or U11311 (N_11311,N_8358,N_5233);
or U11312 (N_11312,N_5678,N_9321);
nor U11313 (N_11313,N_5212,N_8166);
nand U11314 (N_11314,N_5117,N_7748);
xor U11315 (N_11315,N_5333,N_8727);
nand U11316 (N_11316,N_5442,N_7313);
or U11317 (N_11317,N_5893,N_7629);
and U11318 (N_11318,N_5181,N_8920);
xor U11319 (N_11319,N_7241,N_8812);
nand U11320 (N_11320,N_8679,N_8398);
nand U11321 (N_11321,N_9195,N_9468);
or U11322 (N_11322,N_7540,N_6143);
nor U11323 (N_11323,N_8762,N_8622);
and U11324 (N_11324,N_5553,N_5703);
nand U11325 (N_11325,N_6331,N_5776);
xnor U11326 (N_11326,N_7645,N_7073);
or U11327 (N_11327,N_5749,N_6280);
or U11328 (N_11328,N_9835,N_9354);
and U11329 (N_11329,N_8912,N_8154);
xnor U11330 (N_11330,N_9741,N_9482);
nor U11331 (N_11331,N_9397,N_5971);
and U11332 (N_11332,N_8052,N_9248);
nor U11333 (N_11333,N_9866,N_7018);
xnor U11334 (N_11334,N_8795,N_6178);
nor U11335 (N_11335,N_6606,N_8179);
or U11336 (N_11336,N_7689,N_8713);
or U11337 (N_11337,N_8732,N_8589);
xor U11338 (N_11338,N_7329,N_7262);
nand U11339 (N_11339,N_7987,N_7478);
nand U11340 (N_11340,N_6721,N_7545);
nand U11341 (N_11341,N_9333,N_6567);
nand U11342 (N_11342,N_7218,N_5285);
nand U11343 (N_11343,N_5172,N_7122);
nand U11344 (N_11344,N_9988,N_6607);
nor U11345 (N_11345,N_7057,N_8956);
nand U11346 (N_11346,N_7651,N_5886);
nor U11347 (N_11347,N_6080,N_9141);
xnor U11348 (N_11348,N_9373,N_6795);
xor U11349 (N_11349,N_8305,N_5537);
nor U11350 (N_11350,N_7978,N_8556);
or U11351 (N_11351,N_6023,N_8235);
and U11352 (N_11352,N_9821,N_7390);
and U11353 (N_11353,N_8550,N_9523);
nand U11354 (N_11354,N_9994,N_5618);
nand U11355 (N_11355,N_7458,N_7939);
xor U11356 (N_11356,N_9503,N_5293);
or U11357 (N_11357,N_7364,N_7761);
xnor U11358 (N_11358,N_5580,N_9298);
or U11359 (N_11359,N_6226,N_7334);
or U11360 (N_11360,N_6411,N_6187);
xor U11361 (N_11361,N_7011,N_7889);
nor U11362 (N_11362,N_8436,N_5791);
or U11363 (N_11363,N_7751,N_7699);
and U11364 (N_11364,N_5751,N_5906);
and U11365 (N_11365,N_9967,N_6184);
xnor U11366 (N_11366,N_7918,N_5717);
xnor U11367 (N_11367,N_8151,N_8798);
or U11368 (N_11368,N_7311,N_8416);
nand U11369 (N_11369,N_6456,N_9892);
nor U11370 (N_11370,N_6632,N_8839);
and U11371 (N_11371,N_7935,N_7990);
xor U11372 (N_11372,N_6390,N_5565);
and U11373 (N_11373,N_7487,N_9678);
nor U11374 (N_11374,N_5727,N_7894);
and U11375 (N_11375,N_5644,N_8342);
or U11376 (N_11376,N_5554,N_7848);
nand U11377 (N_11377,N_9602,N_7082);
xnor U11378 (N_11378,N_7988,N_8394);
nand U11379 (N_11379,N_8739,N_7006);
or U11380 (N_11380,N_8211,N_5599);
xor U11381 (N_11381,N_6957,N_6365);
or U11382 (N_11382,N_7081,N_5572);
nor U11383 (N_11383,N_8897,N_7602);
or U11384 (N_11384,N_8402,N_7711);
or U11385 (N_11385,N_6924,N_5093);
and U11386 (N_11386,N_8680,N_8637);
nand U11387 (N_11387,N_6985,N_8017);
nand U11388 (N_11388,N_8651,N_5800);
nand U11389 (N_11389,N_7337,N_9177);
and U11390 (N_11390,N_7802,N_6379);
nand U11391 (N_11391,N_5631,N_8125);
and U11392 (N_11392,N_9120,N_7702);
nand U11393 (N_11393,N_7023,N_8543);
xor U11394 (N_11394,N_8743,N_9715);
or U11395 (N_11395,N_6843,N_9817);
xor U11396 (N_11396,N_5949,N_6628);
and U11397 (N_11397,N_6643,N_7323);
nor U11398 (N_11398,N_5719,N_9764);
xnor U11399 (N_11399,N_8042,N_7928);
xor U11400 (N_11400,N_5997,N_9240);
nor U11401 (N_11401,N_8560,N_6575);
xnor U11402 (N_11402,N_9491,N_6292);
and U11403 (N_11403,N_8032,N_5918);
xor U11404 (N_11404,N_8948,N_5764);
or U11405 (N_11405,N_8672,N_8810);
nand U11406 (N_11406,N_5037,N_9928);
nand U11407 (N_11407,N_6947,N_5542);
and U11408 (N_11408,N_5188,N_5616);
and U11409 (N_11409,N_6891,N_8084);
xnor U11410 (N_11410,N_8878,N_8160);
or U11411 (N_11411,N_8523,N_7286);
or U11412 (N_11412,N_8003,N_6222);
nand U11413 (N_11413,N_6576,N_8178);
nor U11414 (N_11414,N_9894,N_8967);
nor U11415 (N_11415,N_7589,N_9356);
or U11416 (N_11416,N_8049,N_8964);
or U11417 (N_11417,N_8258,N_6388);
xor U11418 (N_11418,N_8119,N_7235);
or U11419 (N_11419,N_9032,N_9229);
nand U11420 (N_11420,N_5040,N_7105);
xnor U11421 (N_11421,N_6989,N_5772);
or U11422 (N_11422,N_7968,N_7336);
and U11423 (N_11423,N_7173,N_8012);
nor U11424 (N_11424,N_5566,N_6412);
and U11425 (N_11425,N_5535,N_9877);
xnor U11426 (N_11426,N_5615,N_7630);
and U11427 (N_11427,N_8006,N_5216);
nor U11428 (N_11428,N_6859,N_7698);
or U11429 (N_11429,N_6990,N_8267);
nand U11430 (N_11430,N_9867,N_5597);
and U11431 (N_11431,N_6157,N_6094);
and U11432 (N_11432,N_6988,N_5737);
and U11433 (N_11433,N_5963,N_7305);
nor U11434 (N_11434,N_7266,N_5422);
nand U11435 (N_11435,N_9189,N_5913);
or U11436 (N_11436,N_9463,N_8162);
or U11437 (N_11437,N_9914,N_5424);
or U11438 (N_11438,N_8397,N_5213);
nor U11439 (N_11439,N_8207,N_8724);
or U11440 (N_11440,N_9239,N_8135);
nand U11441 (N_11441,N_5158,N_6592);
or U11442 (N_11442,N_7454,N_8559);
xnor U11443 (N_11443,N_8856,N_5085);
and U11444 (N_11444,N_7108,N_6304);
nand U11445 (N_11445,N_9001,N_5464);
or U11446 (N_11446,N_9300,N_8707);
or U11447 (N_11447,N_5231,N_9430);
xor U11448 (N_11448,N_5473,N_8217);
or U11449 (N_11449,N_6749,N_9873);
nor U11450 (N_11450,N_9510,N_7539);
nor U11451 (N_11451,N_9304,N_6585);
xor U11452 (N_11452,N_6299,N_8175);
or U11453 (N_11453,N_9806,N_9822);
nand U11454 (N_11454,N_5060,N_7749);
and U11455 (N_11455,N_7624,N_9000);
nor U11456 (N_11456,N_7217,N_6071);
nor U11457 (N_11457,N_5936,N_6684);
or U11458 (N_11458,N_5768,N_9698);
or U11459 (N_11459,N_5101,N_7096);
and U11460 (N_11460,N_5328,N_6758);
and U11461 (N_11461,N_9684,N_6552);
or U11462 (N_11462,N_7059,N_9045);
and U11463 (N_11463,N_6323,N_9253);
or U11464 (N_11464,N_5873,N_8220);
nand U11465 (N_11465,N_7035,N_8350);
and U11466 (N_11466,N_5834,N_8034);
xnor U11467 (N_11467,N_7015,N_7844);
nor U11468 (N_11468,N_9470,N_7184);
nand U11469 (N_11469,N_5064,N_8566);
nand U11470 (N_11470,N_7321,N_6981);
or U11471 (N_11471,N_9349,N_6447);
or U11472 (N_11472,N_7317,N_8652);
or U11473 (N_11473,N_8495,N_8263);
or U11474 (N_11474,N_5627,N_6428);
nand U11475 (N_11475,N_7764,N_9946);
xnor U11476 (N_11476,N_5447,N_9898);
nor U11477 (N_11477,N_6122,N_8824);
nand U11478 (N_11478,N_7809,N_6867);
nand U11479 (N_11479,N_6902,N_6594);
nor U11480 (N_11480,N_8832,N_7886);
nor U11481 (N_11481,N_8919,N_8129);
xor U11482 (N_11482,N_5313,N_5519);
and U11483 (N_11483,N_6884,N_7864);
nor U11484 (N_11484,N_6242,N_7716);
and U11485 (N_11485,N_8881,N_8324);
nand U11486 (N_11486,N_5693,N_8700);
or U11487 (N_11487,N_9359,N_5581);
xnor U11488 (N_11488,N_9644,N_6803);
and U11489 (N_11489,N_6435,N_5106);
xnor U11490 (N_11490,N_7047,N_8644);
and U11491 (N_11491,N_8793,N_9308);
nor U11492 (N_11492,N_8440,N_8532);
or U11493 (N_11493,N_8123,N_5563);
nand U11494 (N_11494,N_9827,N_9384);
nor U11495 (N_11495,N_9660,N_5938);
xor U11496 (N_11496,N_9200,N_7622);
and U11497 (N_11497,N_7440,N_6290);
nand U11498 (N_11498,N_8041,N_6685);
or U11499 (N_11499,N_8089,N_8241);
nand U11500 (N_11500,N_6111,N_8702);
and U11501 (N_11501,N_8214,N_9212);
or U11502 (N_11502,N_7825,N_7897);
nand U11503 (N_11503,N_8867,N_5428);
xnor U11504 (N_11504,N_8329,N_9692);
xor U11505 (N_11505,N_6260,N_9379);
and U11506 (N_11506,N_7862,N_7757);
xor U11507 (N_11507,N_8303,N_6958);
nor U11508 (N_11508,N_5377,N_5348);
nand U11509 (N_11509,N_7694,N_5915);
xor U11510 (N_11510,N_7879,N_9596);
nand U11511 (N_11511,N_6273,N_7955);
and U11512 (N_11512,N_6330,N_9398);
nand U11513 (N_11513,N_8379,N_5773);
xnor U11514 (N_11514,N_7746,N_9944);
and U11515 (N_11515,N_8520,N_5608);
or U11516 (N_11516,N_8913,N_8740);
nand U11517 (N_11517,N_9668,N_6373);
nor U11518 (N_11518,N_5898,N_9283);
nor U11519 (N_11519,N_8633,N_9577);
or U11520 (N_11520,N_8823,N_7344);
xnor U11521 (N_11521,N_7232,N_5444);
nor U11522 (N_11522,N_5613,N_6084);
and U11523 (N_11523,N_8508,N_7577);
nor U11524 (N_11524,N_5846,N_7574);
or U11525 (N_11525,N_6831,N_5120);
nor U11526 (N_11526,N_8598,N_8846);
xnor U11527 (N_11527,N_6189,N_7793);
or U11528 (N_11528,N_9982,N_5389);
and U11529 (N_11529,N_9166,N_8437);
xor U11530 (N_11530,N_9643,N_7706);
xnor U11531 (N_11531,N_5168,N_7794);
and U11532 (N_11532,N_8124,N_9462);
nor U11533 (N_11533,N_7985,N_9628);
nor U11534 (N_11534,N_5698,N_5931);
nand U11535 (N_11535,N_6883,N_7289);
and U11536 (N_11536,N_7835,N_7264);
nor U11537 (N_11537,N_8563,N_5236);
or U11538 (N_11538,N_8389,N_6814);
nand U11539 (N_11539,N_9961,N_9380);
nand U11540 (N_11540,N_7851,N_9832);
xnor U11541 (N_11541,N_8675,N_9346);
or U11542 (N_11542,N_8105,N_9020);
and U11543 (N_11543,N_7017,N_7076);
nand U11544 (N_11544,N_6706,N_8836);
nor U11545 (N_11545,N_7859,N_5785);
or U11546 (N_11546,N_8942,N_7787);
or U11547 (N_11547,N_8111,N_9143);
xor U11548 (N_11548,N_7178,N_8941);
nor U11549 (N_11549,N_9593,N_7226);
nor U11550 (N_11550,N_6115,N_5241);
and U11551 (N_11551,N_7546,N_5322);
xnor U11552 (N_11552,N_9106,N_5090);
nor U11553 (N_11553,N_9630,N_7695);
xnor U11554 (N_11554,N_8646,N_9021);
nor U11555 (N_11555,N_7700,N_8387);
xor U11556 (N_11556,N_6880,N_6404);
nand U11557 (N_11557,N_5663,N_5007);
and U11558 (N_11558,N_9762,N_9992);
or U11559 (N_11559,N_8077,N_8014);
nand U11560 (N_11560,N_5496,N_9317);
nor U11561 (N_11561,N_6731,N_8737);
xor U11562 (N_11562,N_5119,N_9578);
or U11563 (N_11563,N_6034,N_5712);
or U11564 (N_11564,N_6043,N_8898);
or U11565 (N_11565,N_7066,N_7074);
xor U11566 (N_11566,N_7462,N_6465);
or U11567 (N_11567,N_8093,N_9846);
xor U11568 (N_11568,N_9807,N_8758);
and U11569 (N_11569,N_6423,N_8116);
or U11570 (N_11570,N_7596,N_9083);
or U11571 (N_11571,N_9487,N_8367);
nand U11572 (N_11572,N_5050,N_7910);
nor U11573 (N_11573,N_6106,N_7713);
nor U11574 (N_11574,N_6846,N_5880);
xor U11575 (N_11575,N_8347,N_9033);
nand U11576 (N_11576,N_6586,N_7655);
nor U11577 (N_11577,N_8225,N_5436);
or U11578 (N_11578,N_8299,N_7529);
or U11579 (N_11579,N_7820,N_6223);
xnor U11580 (N_11580,N_7308,N_8195);
nor U11581 (N_11581,N_5723,N_5441);
nand U11582 (N_11582,N_8837,N_9210);
and U11583 (N_11583,N_6515,N_9071);
or U11584 (N_11584,N_8351,N_7812);
or U11585 (N_11585,N_6434,N_5220);
or U11586 (N_11586,N_6004,N_6558);
nor U11587 (N_11587,N_9535,N_9023);
or U11588 (N_11588,N_6398,N_5781);
xor U11589 (N_11589,N_6076,N_8140);
nor U11590 (N_11590,N_5769,N_8545);
and U11591 (N_11591,N_7778,N_6220);
nor U11592 (N_11592,N_6698,N_9193);
xor U11593 (N_11593,N_8200,N_5134);
and U11594 (N_11594,N_5448,N_9323);
or U11595 (N_11595,N_8903,N_5407);
nand U11596 (N_11596,N_7447,N_9871);
and U11597 (N_11597,N_6308,N_7679);
xnor U11598 (N_11598,N_5143,N_7615);
and U11599 (N_11599,N_6998,N_6061);
or U11600 (N_11600,N_8595,N_9118);
or U11601 (N_11601,N_7065,N_5109);
xnor U11602 (N_11602,N_8448,N_5850);
or U11603 (N_11603,N_6967,N_7391);
nand U11604 (N_11604,N_8230,N_6322);
or U11605 (N_11605,N_5832,N_7097);
or U11606 (N_11606,N_6520,N_5150);
xor U11607 (N_11607,N_7866,N_6344);
nor U11608 (N_11608,N_8407,N_5529);
nand U11609 (N_11609,N_6333,N_6763);
and U11610 (N_11610,N_5524,N_9879);
nor U11611 (N_11611,N_7984,N_8525);
xor U11612 (N_11612,N_9122,N_5485);
or U11613 (N_11613,N_9419,N_6751);
nand U11614 (N_11614,N_6909,N_8828);
nand U11615 (N_11615,N_5610,N_5843);
and U11616 (N_11616,N_6263,N_8468);
or U11617 (N_11617,N_8366,N_8805);
nand U11618 (N_11618,N_5861,N_9316);
and U11619 (N_11619,N_6192,N_9080);
nor U11620 (N_11620,N_8802,N_6479);
nor U11621 (N_11621,N_8001,N_8570);
nand U11622 (N_11622,N_6103,N_5623);
or U11623 (N_11623,N_5144,N_6235);
nor U11624 (N_11624,N_8544,N_6664);
and U11625 (N_11625,N_9225,N_6317);
xor U11626 (N_11626,N_6530,N_6095);
or U11627 (N_11627,N_5141,N_9520);
xor U11628 (N_11628,N_5292,N_9438);
nand U11629 (N_11629,N_7569,N_6739);
and U11630 (N_11630,N_7269,N_9184);
nor U11631 (N_11631,N_8008,N_6406);
nand U11632 (N_11632,N_9013,N_6225);
nand U11633 (N_11633,N_8359,N_8493);
xnor U11634 (N_11634,N_9350,N_8522);
or U11635 (N_11635,N_6978,N_5792);
xor U11636 (N_11636,N_9048,N_6881);
nor U11637 (N_11637,N_5590,N_7530);
nor U11638 (N_11638,N_6666,N_8204);
xnor U11639 (N_11639,N_8183,N_8617);
xor U11640 (N_11640,N_9856,N_8712);
xor U11641 (N_11641,N_7729,N_8664);
or U11642 (N_11642,N_6756,N_5239);
xor U11643 (N_11643,N_6018,N_9493);
and U11644 (N_11644,N_6015,N_6236);
nor U11645 (N_11645,N_5462,N_6203);
nor U11646 (N_11646,N_8423,N_6524);
nor U11647 (N_11647,N_8460,N_8033);
or U11648 (N_11648,N_9910,N_5739);
nand U11649 (N_11649,N_5431,N_7960);
xnor U11650 (N_11650,N_5562,N_8172);
xor U11651 (N_11651,N_9414,N_8817);
nand U11652 (N_11652,N_9424,N_7669);
and U11653 (N_11653,N_5087,N_6944);
nor U11654 (N_11654,N_6728,N_9518);
xor U11655 (N_11655,N_6462,N_9162);
or U11656 (N_11656,N_6093,N_6667);
nor U11657 (N_11657,N_7740,N_9452);
and U11658 (N_11658,N_9338,N_5812);
or U11659 (N_11659,N_6730,N_8412);
nor U11660 (N_11660,N_9724,N_9235);
or U11661 (N_11661,N_5530,N_8922);
nor U11662 (N_11662,N_9791,N_6580);
nor U11663 (N_11663,N_9269,N_9588);
nor U11664 (N_11664,N_8239,N_9094);
xor U11665 (N_11665,N_8820,N_7293);
and U11666 (N_11666,N_6939,N_6503);
or U11667 (N_11667,N_8924,N_8075);
and U11668 (N_11668,N_9792,N_5743);
xor U11669 (N_11669,N_5877,N_6156);
or U11670 (N_11670,N_6297,N_5278);
xnor U11671 (N_11671,N_7537,N_5604);
and U11672 (N_11672,N_9058,N_5252);
nor U11673 (N_11673,N_7821,N_8954);
nand U11674 (N_11674,N_8968,N_8745);
and U11675 (N_11675,N_8969,N_8485);
nand U11676 (N_11676,N_7924,N_6013);
nor U11677 (N_11677,N_6082,N_8979);
xnor U11678 (N_11678,N_7792,N_7753);
xnor U11679 (N_11679,N_7819,N_9850);
and U11680 (N_11680,N_9395,N_7356);
or U11681 (N_11681,N_6699,N_7214);
xor U11682 (N_11682,N_8811,N_5326);
nor U11683 (N_11683,N_9394,N_8943);
nand U11684 (N_11684,N_7430,N_8094);
nor U11685 (N_11685,N_9448,N_7904);
nand U11686 (N_11686,N_5151,N_7324);
nand U11687 (N_11687,N_6233,N_8923);
or U11688 (N_11688,N_6518,N_9591);
and U11689 (N_11689,N_9554,N_8381);
or U11690 (N_11690,N_5307,N_5438);
nor U11691 (N_11691,N_8114,N_5443);
and U11692 (N_11692,N_6332,N_7547);
xnor U11693 (N_11693,N_8962,N_9026);
and U11694 (N_11694,N_8982,N_7372);
or U11695 (N_11695,N_8459,N_9301);
and U11696 (N_11696,N_7690,N_5075);
or U11697 (N_11697,N_6354,N_9444);
and U11698 (N_11698,N_5556,N_8302);
xnor U11699 (N_11699,N_5989,N_5073);
and U11700 (N_11700,N_5534,N_6051);
nand U11701 (N_11701,N_7830,N_9572);
or U11702 (N_11702,N_8252,N_6500);
or U11703 (N_11703,N_7617,N_6356);
and U11704 (N_11704,N_9077,N_8104);
nor U11705 (N_11705,N_9387,N_6782);
nor U11706 (N_11706,N_8852,N_9263);
xor U11707 (N_11707,N_5033,N_5987);
xor U11708 (N_11708,N_7114,N_7562);
or U11709 (N_11709,N_8555,N_6183);
xnor U11710 (N_11710,N_9633,N_9984);
and U11711 (N_11711,N_6813,N_6405);
or U11712 (N_11712,N_6230,N_7378);
nand U11713 (N_11713,N_6491,N_5353);
nor U11714 (N_11714,N_7119,N_9581);
xor U11715 (N_11715,N_6923,N_6614);
or U11716 (N_11716,N_9649,N_6817);
nor U11717 (N_11717,N_5393,N_6396);
xnor U11718 (N_11718,N_5036,N_7194);
or U11719 (N_11719,N_5594,N_9272);
nor U11720 (N_11720,N_6876,N_8261);
and U11721 (N_11721,N_7278,N_6166);
nor U11722 (N_11722,N_9897,N_5383);
and U11723 (N_11723,N_5659,N_7816);
and U11724 (N_11724,N_6038,N_7913);
nor U11725 (N_11725,N_8785,N_6397);
xnor U11726 (N_11726,N_5291,N_5063);
and U11727 (N_11727,N_7509,N_5818);
or U11728 (N_11728,N_7043,N_6800);
and U11729 (N_11729,N_7502,N_5325);
nor U11730 (N_11730,N_8748,N_8097);
nor U11731 (N_11731,N_9647,N_7721);
nand U11732 (N_11732,N_9445,N_6599);
or U11733 (N_11733,N_5609,N_7437);
or U11734 (N_11734,N_9638,N_6717);
nor U11735 (N_11735,N_8643,N_7328);
or U11736 (N_11736,N_6984,N_5920);
nor U11737 (N_11737,N_7531,N_5626);
or U11738 (N_11738,N_7967,N_8773);
and U11739 (N_11739,N_7754,N_6996);
and U11740 (N_11740,N_5493,N_5966);
or U11741 (N_11741,N_6048,N_6381);
and U11742 (N_11742,N_5939,N_9075);
and U11743 (N_11743,N_9746,N_8294);
and U11744 (N_11744,N_6950,N_7770);
or U11745 (N_11745,N_8676,N_9731);
or U11746 (N_11746,N_9516,N_8048);
nor U11747 (N_11747,N_5180,N_5808);
and U11748 (N_11748,N_9072,N_5165);
and U11749 (N_11749,N_9199,N_5217);
and U11750 (N_11750,N_8233,N_6914);
or U11751 (N_11751,N_8209,N_7771);
nor U11752 (N_11752,N_5039,N_5317);
nand U11753 (N_11753,N_8057,N_8206);
xor U11754 (N_11754,N_7704,N_5547);
xnor U11755 (N_11755,N_5416,N_7077);
xor U11756 (N_11756,N_5875,N_8682);
nand U11757 (N_11757,N_9377,N_9390);
xor U11758 (N_11758,N_6204,N_7660);
nor U11759 (N_11759,N_5991,N_9207);
and U11760 (N_11760,N_8695,N_7026);
or U11761 (N_11761,N_5357,N_5004);
nor U11762 (N_11762,N_8215,N_6780);
or U11763 (N_11763,N_9158,N_9309);
nand U11764 (N_11764,N_8442,N_9165);
xor U11765 (N_11765,N_6912,N_9964);
and U11766 (N_11766,N_5410,N_8372);
and U11767 (N_11767,N_8144,N_5099);
and U11768 (N_11768,N_7800,N_9880);
nor U11769 (N_11769,N_7491,N_7486);
xnor U11770 (N_11770,N_8223,N_8765);
or U11771 (N_11771,N_9204,N_6864);
xor U11772 (N_11772,N_5078,N_8108);
and U11773 (N_11773,N_5667,N_8257);
and U11774 (N_11774,N_5914,N_9955);
nand U11775 (N_11775,N_6587,N_7247);
and U11776 (N_11776,N_7563,N_8184);
and U11777 (N_11777,N_6200,N_8915);
and U11778 (N_11778,N_6896,N_9016);
xor U11779 (N_11779,N_5148,N_6105);
xor U11780 (N_11780,N_7393,N_5677);
nor U11781 (N_11781,N_8480,N_5825);
xor U11782 (N_11782,N_7870,N_7592);
nand U11783 (N_11783,N_5323,N_8419);
and U11784 (N_11784,N_8149,N_6894);
and U11785 (N_11785,N_7790,N_7907);
or U11786 (N_11786,N_6773,N_7270);
or U11787 (N_11787,N_8620,N_8689);
xor U11788 (N_11788,N_9187,N_6017);
and U11789 (N_11789,N_9579,N_5658);
or U11790 (N_11790,N_5020,N_9889);
and U11791 (N_11791,N_6862,N_5187);
nand U11792 (N_11792,N_6395,N_6707);
and U11793 (N_11793,N_9280,N_5459);
or U11794 (N_11794,N_6148,N_6489);
nand U11795 (N_11795,N_6196,N_6830);
xnor U11796 (N_11796,N_8234,N_5258);
xor U11797 (N_11797,N_9274,N_6645);
xnor U11798 (N_11798,N_7664,N_5981);
and U11799 (N_11799,N_7979,N_8473);
nor U11800 (N_11800,N_5996,N_8760);
and U11801 (N_11801,N_5826,N_7954);
or U11802 (N_11802,N_5517,N_7822);
nor U11803 (N_11803,N_9925,N_5533);
xnor U11804 (N_11804,N_6185,N_8610);
nor U11805 (N_11805,N_8434,N_5426);
or U11806 (N_11806,N_9519,N_7211);
xor U11807 (N_11807,N_9289,N_7485);
xor U11808 (N_11808,N_5301,N_7636);
and U11809 (N_11809,N_7853,N_8283);
xor U11810 (N_11810,N_7824,N_8655);
xor U11811 (N_11811,N_5596,N_6109);
or U11812 (N_11812,N_7249,N_9969);
nand U11813 (N_11813,N_9779,N_6083);
and U11814 (N_11814,N_9828,N_6807);
nand U11815 (N_11815,N_7063,N_9188);
nor U11816 (N_11816,N_9530,N_5842);
nand U11817 (N_11817,N_5738,N_7414);
and U11818 (N_11818,N_6525,N_9517);
nor U11819 (N_11819,N_7123,N_8100);
or U11820 (N_11820,N_6279,N_5068);
and U11821 (N_11821,N_7242,N_6393);
nand U11822 (N_11822,N_6507,N_5635);
or U11823 (N_11823,N_6078,N_8439);
or U11824 (N_11824,N_7482,N_9243);
or U11825 (N_11825,N_5699,N_6868);
and U11826 (N_11826,N_8404,N_6986);
xnor U11827 (N_11827,N_9755,N_8177);
xor U11828 (N_11828,N_5107,N_9549);
xor U11829 (N_11829,N_9477,N_5334);
nand U11830 (N_11830,N_9797,N_8218);
nor U11831 (N_11831,N_6709,N_8286);
nor U11832 (N_11832,N_5688,N_8391);
xnor U11833 (N_11833,N_5155,N_6246);
and U11834 (N_11834,N_8457,N_6059);
and U11835 (N_11835,N_7611,N_8348);
and U11836 (N_11836,N_6823,N_7256);
nor U11837 (N_11837,N_8474,N_6049);
or U11838 (N_11838,N_6983,N_9987);
nand U11839 (N_11839,N_9837,N_6407);
xnor U11840 (N_11840,N_8966,N_9829);
nand U11841 (N_11841,N_8880,N_7248);
nand U11842 (N_11842,N_6856,N_8188);
or U11843 (N_11843,N_5359,N_5145);
xor U11844 (N_11844,N_6997,N_7741);
xnor U11845 (N_11845,N_6557,N_7783);
and U11846 (N_11846,N_8361,N_5943);
and U11847 (N_11847,N_5401,N_7303);
xor U11848 (N_11848,N_8797,N_6296);
nor U11849 (N_11849,N_7158,N_6137);
and U11850 (N_11850,N_8483,N_7327);
and U11851 (N_11851,N_6469,N_9878);
and U11852 (N_11852,N_5178,N_8011);
nor U11853 (N_11853,N_9053,N_5646);
xor U11854 (N_11854,N_5640,N_6470);
nor U11855 (N_11855,N_7418,N_9651);
and U11856 (N_11856,N_9429,N_5708);
and U11857 (N_11857,N_7193,N_8729);
or U11858 (N_11858,N_9699,N_5747);
or U11859 (N_11859,N_6371,N_5057);
nand U11860 (N_11860,N_9069,N_7868);
nand U11861 (N_11861,N_6401,N_8055);
nand U11862 (N_11862,N_6449,N_8430);
or U11863 (N_11863,N_8180,N_7162);
or U11864 (N_11864,N_9935,N_6338);
xnor U11865 (N_11865,N_7222,N_9753);
xor U11866 (N_11866,N_5934,N_8260);
nand U11867 (N_11867,N_5028,N_9794);
nand U11868 (N_11868,N_8496,N_5672);
or U11869 (N_11869,N_5790,N_5115);
nor U11870 (N_11870,N_6455,N_7197);
or U11871 (N_11871,N_8251,N_7620);
and U11872 (N_11872,N_9559,N_7368);
nand U11873 (N_11873,N_6362,N_6377);
or U11874 (N_11874,N_7610,N_7187);
nor U11875 (N_11875,N_8343,N_8908);
and U11876 (N_11876,N_8462,N_5753);
and U11877 (N_11877,N_8991,N_8761);
nor U11878 (N_11878,N_9847,N_6748);
xor U11879 (N_11879,N_5154,N_6079);
xnor U11880 (N_11880,N_8981,N_5577);
xnor U11881 (N_11881,N_9355,N_8210);
or U11882 (N_11882,N_5950,N_5881);
xnor U11883 (N_11883,N_5298,N_6678);
nand U11884 (N_11884,N_7788,N_6661);
xor U11885 (N_11885,N_6718,N_8653);
nor U11886 (N_11886,N_8593,N_6052);
xor U11887 (N_11887,N_6478,N_8896);
or U11888 (N_11888,N_9617,N_8066);
xnor U11889 (N_11889,N_6754,N_8022);
nand U11890 (N_11890,N_6239,N_9421);
nor U11891 (N_11891,N_8445,N_8458);
nand U11892 (N_11892,N_8639,N_5919);
nand U11893 (N_11893,N_5003,N_9546);
nor U11894 (N_11894,N_7325,N_8500);
or U11895 (N_11895,N_5922,N_8835);
or U11896 (N_11896,N_5400,N_9958);
xor U11897 (N_11897,N_9467,N_8792);
nor U11898 (N_11898,N_8396,N_8721);
nand U11899 (N_11899,N_9004,N_9091);
nor U11900 (N_11900,N_7784,N_8272);
nor U11901 (N_11901,N_6965,N_7696);
xor U11902 (N_11902,N_6620,N_9409);
nor U11903 (N_11903,N_9149,N_6657);
xor U11904 (N_11904,N_5975,N_6511);
or U11905 (N_11905,N_9237,N_7287);
and U11906 (N_11906,N_9218,N_8092);
nand U11907 (N_11907,N_5262,N_5091);
nand U11908 (N_11908,N_7254,N_7914);
or U11909 (N_11909,N_5910,N_6570);
xor U11910 (N_11910,N_6384,N_9116);
nand U11911 (N_11911,N_9561,N_6114);
xnor U11912 (N_11912,N_9327,N_6128);
nor U11913 (N_11913,N_8813,N_5892);
nor U11914 (N_11914,N_6851,N_5390);
nand U11915 (N_11915,N_8156,N_8696);
xnor U11916 (N_11916,N_9140,N_6514);
or U11917 (N_11917,N_8030,N_9362);
nor U11918 (N_11918,N_9271,N_6925);
or U11919 (N_11919,N_8949,N_6674);
nor U11920 (N_11920,N_5021,N_9095);
nand U11921 (N_11921,N_5888,N_6345);
xnor U11922 (N_11922,N_6702,N_5745);
nor U11923 (N_11923,N_7288,N_5305);
nor U11924 (N_11924,N_6822,N_6261);
nor U11925 (N_11925,N_5787,N_7687);
nor U11926 (N_11926,N_9041,N_9981);
and U11927 (N_11927,N_5951,N_9661);
nor U11928 (N_11928,N_6160,N_9657);
nor U11929 (N_11929,N_8963,N_5125);
and U11930 (N_11930,N_7170,N_9292);
xor U11931 (N_11931,N_7467,N_9534);
nand U11932 (N_11932,N_8684,N_5945);
and U11933 (N_11933,N_7183,N_9055);
or U11934 (N_11934,N_9353,N_8603);
and U11935 (N_11935,N_8355,N_6353);
nand U11936 (N_11936,N_9851,N_8333);
and U11937 (N_11937,N_7598,N_8907);
nand U11938 (N_11938,N_9618,N_6591);
nand U11939 (N_11939,N_5008,N_5472);
xnor U11940 (N_11940,N_9536,N_5449);
nor U11941 (N_11941,N_7663,N_6625);
nand U11942 (N_11942,N_8735,N_6483);
and U11943 (N_11943,N_9352,N_9611);
or U11944 (N_11944,N_7628,N_8269);
or U11945 (N_11945,N_7424,N_9388);
nor U11946 (N_11946,N_5833,N_5671);
nand U11947 (N_11947,N_6475,N_5498);
nor U11948 (N_11948,N_9655,N_7878);
nand U11949 (N_11949,N_5854,N_8604);
and U11950 (N_11950,N_8944,N_9640);
nand U11951 (N_11951,N_8134,N_6613);
nor U11952 (N_11952,N_8378,N_8187);
or U11953 (N_11953,N_5055,N_6855);
or U11954 (N_11954,N_5756,N_9167);
nor U11955 (N_11955,N_9126,N_6238);
nor U11956 (N_11956,N_7231,N_7190);
xor U11957 (N_11957,N_6459,N_6920);
nand U11958 (N_11958,N_6152,N_7133);
nor U11959 (N_11959,N_8043,N_9927);
xor U11960 (N_11960,N_8893,N_9125);
xnor U11961 (N_11961,N_6775,N_8601);
nand U11962 (N_11962,N_8698,N_5059);
or U11963 (N_11963,N_7516,N_8323);
xnor U11964 (N_11964,N_6019,N_8068);
nor U11965 (N_11965,N_7392,N_8803);
or U11966 (N_11966,N_7743,N_9098);
nand U11967 (N_11967,N_9488,N_9730);
nand U11968 (N_11968,N_9437,N_8789);
nor U11969 (N_11969,N_8770,N_8356);
and U11970 (N_11970,N_7580,N_9008);
and U11971 (N_11971,N_6647,N_5332);
and U11972 (N_11972,N_6402,N_7290);
nand U11973 (N_11973,N_5526,N_6584);
nor U11974 (N_11974,N_7032,N_5965);
or U11975 (N_11975,N_5532,N_7597);
nand U11976 (N_11976,N_7737,N_6642);
or U11977 (N_11977,N_6042,N_5700);
xor U11978 (N_11978,N_9694,N_5199);
nand U11979 (N_11979,N_9290,N_8492);
nand U11980 (N_11980,N_9100,N_9703);
nor U11981 (N_11981,N_9286,N_8864);
nand U11982 (N_11982,N_8388,N_8557);
nand U11983 (N_11983,N_8849,N_9281);
or U11984 (N_11984,N_7963,N_8549);
xor U11985 (N_11985,N_5586,N_7200);
xnor U11986 (N_11986,N_9956,N_8845);
and U11987 (N_11987,N_7460,N_6826);
nor U11988 (N_11988,N_9838,N_7161);
nor U11989 (N_11989,N_8650,N_7828);
xor U11990 (N_11990,N_5434,N_8318);
or U11991 (N_11991,N_6025,N_9466);
or U11992 (N_11992,N_5435,N_6850);
nor U11993 (N_11993,N_8970,N_6513);
nand U11994 (N_11994,N_5548,N_7667);
and U11995 (N_11995,N_9420,N_9393);
xnor U11996 (N_11996,N_7882,N_5089);
and U11997 (N_11997,N_8293,N_6919);
xor U11998 (N_11998,N_5816,N_9765);
or U11999 (N_11999,N_7147,N_7471);
xor U12000 (N_12000,N_5782,N_8332);
nand U12001 (N_12001,N_8456,N_6619);
xor U12002 (N_12002,N_7534,N_6144);
xor U12003 (N_12003,N_8535,N_8709);
and U12004 (N_12004,N_9893,N_8384);
xnor U12005 (N_12005,N_9505,N_5338);
nor U12006 (N_12006,N_8829,N_7120);
nand U12007 (N_12007,N_7284,N_8730);
nand U12008 (N_12008,N_6804,N_5935);
nor U12009 (N_12009,N_8983,N_9567);
or U12010 (N_12010,N_7607,N_9279);
or U12011 (N_12011,N_9404,N_6168);
nor U12012 (N_12012,N_9675,N_7362);
and U12013 (N_12013,N_6147,N_8113);
xnor U12014 (N_12014,N_7901,N_9480);
xnor U12015 (N_12015,N_6163,N_5643);
or U12016 (N_12016,N_8110,N_9884);
nor U12017 (N_12017,N_6451,N_5056);
and U12018 (N_12018,N_9974,N_8417);
nand U12019 (N_12019,N_8330,N_7769);
xnor U12020 (N_12020,N_7843,N_9721);
nor U12021 (N_12021,N_9170,N_8069);
xnor U12022 (N_12022,N_8047,N_6195);
xnor U12023 (N_12023,N_7140,N_7382);
nor U12024 (N_12024,N_8533,N_9224);
nor U12025 (N_12025,N_6762,N_7665);
xor U12026 (N_12026,N_5484,N_7100);
nand U12027 (N_12027,N_5973,N_9547);
nand U12028 (N_12028,N_6016,N_5297);
xor U12029 (N_12029,N_7012,N_7883);
or U12030 (N_12030,N_9088,N_8441);
nor U12031 (N_12031,N_5598,N_9842);
and U12032 (N_12032,N_6734,N_9566);
nand U12033 (N_12033,N_7559,N_5946);
nor U12034 (N_12034,N_7298,N_7718);
or U12035 (N_12035,N_7387,N_9979);
and U12036 (N_12036,N_5686,N_6208);
nand U12037 (N_12037,N_7613,N_9109);
or U12038 (N_12038,N_5169,N_9411);
nor U12039 (N_12039,N_8703,N_5053);
and U12040 (N_12040,N_5694,N_7255);
nor U12041 (N_12041,N_9425,N_8062);
nand U12042 (N_12042,N_9264,N_9876);
or U12043 (N_12043,N_8203,N_7477);
xor U12044 (N_12044,N_8808,N_6784);
xor U12045 (N_12045,N_7538,N_7175);
nand U12046 (N_12046,N_6654,N_7239);
and U12047 (N_12047,N_9639,N_8953);
nand U12048 (N_12048,N_6030,N_7583);
xor U12049 (N_12049,N_6488,N_6633);
nor U12050 (N_12050,N_9441,N_8285);
nand U12051 (N_12051,N_7033,N_7556);
nor U12052 (N_12052,N_5458,N_8421);
or U12053 (N_12053,N_7801,N_8335);
or U12054 (N_12054,N_9575,N_9147);
or U12055 (N_12055,N_7463,N_5961);
or U12056 (N_12056,N_6900,N_8581);
or U12057 (N_12057,N_6724,N_9275);
xnor U12058 (N_12058,N_9654,N_6551);
nor U12059 (N_12059,N_8248,N_9574);
or U12060 (N_12060,N_6593,N_9659);
xnor U12061 (N_12061,N_9957,N_6336);
nand U12062 (N_12062,N_6838,N_7064);
nand U12063 (N_12063,N_6450,N_6251);
or U12064 (N_12064,N_9952,N_9230);
and U12065 (N_12065,N_5788,N_9963);
nand U12066 (N_12066,N_9273,N_7031);
and U12067 (N_12067,N_6098,N_9208);
or U12068 (N_12068,N_8842,N_8814);
nor U12069 (N_12069,N_5186,N_9550);
or U12070 (N_12070,N_5520,N_6284);
and U12071 (N_12071,N_6887,N_5821);
and U12072 (N_12072,N_5665,N_6690);
nand U12073 (N_12073,N_8678,N_6182);
or U12074 (N_12074,N_7350,N_6124);
nor U12075 (N_12075,N_5673,N_5988);
nor U12076 (N_12076,N_6934,N_8973);
xnor U12077 (N_12077,N_5067,N_6729);
or U12078 (N_12078,N_8562,N_8932);
nor U12079 (N_12079,N_6636,N_5940);
and U12080 (N_12080,N_7876,N_7080);
or U12081 (N_12081,N_7030,N_6555);
nor U12082 (N_12082,N_9011,N_6255);
and U12083 (N_12083,N_5368,N_8848);
or U12084 (N_12084,N_8851,N_5979);
or U12085 (N_12085,N_5871,N_5350);
or U12086 (N_12086,N_6495,N_8328);
nand U12087 (N_12087,N_7865,N_9082);
nand U12088 (N_12088,N_6306,N_5372);
nand U12089 (N_12089,N_6918,N_9767);
nor U12090 (N_12090,N_7333,N_8013);
nor U12091 (N_12091,N_9198,N_6999);
and U12092 (N_12092,N_9454,N_5651);
and U12093 (N_12093,N_9504,N_8277);
and U12094 (N_12094,N_8264,N_6243);
or U12095 (N_12095,N_8894,N_7139);
and U12096 (N_12096,N_5413,N_6761);
xnor U12097 (N_12097,N_7212,N_7473);
or U12098 (N_12098,N_9364,N_8139);
or U12099 (N_12099,N_7371,N_8363);
nor U12100 (N_12100,N_8454,N_6206);
or U12101 (N_12101,N_6695,N_7989);
and U12102 (N_12102,N_7456,N_8369);
nand U12103 (N_12103,N_5189,N_7433);
and U12104 (N_12104,N_5052,N_5909);
nand U12105 (N_12105,N_8564,N_5632);
nor U12106 (N_12106,N_5582,N_6391);
nand U12107 (N_12107,N_8205,N_9137);
xor U12108 (N_12108,N_7435,N_6473);
nor U12109 (N_12109,N_6194,N_8025);
nand U12110 (N_12110,N_5098,N_7957);
and U12111 (N_12111,N_5701,N_6917);
xor U12112 (N_12112,N_7804,N_6259);
xnor U12113 (N_12113,N_5797,N_5294);
nand U12114 (N_12114,N_8799,N_9119);
and U12115 (N_12115,N_6556,N_5190);
nand U12116 (N_12116,N_9820,N_9233);
and U12117 (N_12117,N_8476,N_8087);
and U12118 (N_12118,N_8425,N_5684);
or U12119 (N_12119,N_8232,N_6100);
nor U12120 (N_12120,N_5355,N_7276);
nor U12121 (N_12121,N_7164,N_5855);
or U12122 (N_12122,N_7776,N_6774);
or U12123 (N_12123,N_6066,N_6760);
nor U12124 (N_12124,N_9396,N_6218);
nor U12125 (N_12125,N_7004,N_6022);
xor U12126 (N_12126,N_6214,N_5380);
or U12127 (N_12127,N_7709,N_9650);
xnor U12128 (N_12128,N_8197,N_5657);
and U12129 (N_12129,N_6951,N_5809);
or U12130 (N_12130,N_9009,N_7921);
nor U12131 (N_12131,N_9995,N_8061);
nand U12132 (N_12132,N_7136,N_9252);
or U12133 (N_12133,N_8053,N_6686);
nand U12134 (N_12134,N_5549,N_6715);
nand U12135 (N_12135,N_7503,N_7423);
xor U12136 (N_12136,N_5011,N_8121);
xnor U12137 (N_12137,N_6490,N_6679);
or U12138 (N_12138,N_9135,N_6630);
or U12139 (N_12139,N_5933,N_8744);
or U12140 (N_12140,N_5102,N_6866);
nand U12141 (N_12141,N_7588,N_6141);
and U12142 (N_12142,N_5852,N_8176);
nand U12143 (N_12143,N_8279,N_9690);
nor U12144 (N_12144,N_9513,N_5482);
or U12145 (N_12145,N_7915,N_7518);
xor U12146 (N_12146,N_6302,N_9385);
and U12147 (N_12147,N_8565,N_8511);
xor U12148 (N_12148,N_8779,N_9412);
or U12149 (N_12149,N_6516,N_9772);
or U12150 (N_12150,N_5923,N_7688);
nand U12151 (N_12151,N_5468,N_9580);
xnor U12152 (N_12152,N_9999,N_6681);
nand U12153 (N_12153,N_7767,N_9624);
nor U12154 (N_12154,N_9326,N_7075);
nand U12155 (N_12155,N_5025,N_7519);
nand U12156 (N_12156,N_5166,N_7930);
xnor U12157 (N_12157,N_7895,N_8989);
or U12158 (N_12158,N_6905,N_6039);
and U12159 (N_12159,N_7282,N_9626);
and U12160 (N_12160,N_7358,N_8504);
xnor U12161 (N_12161,N_9232,N_5367);
xnor U12162 (N_12162,N_9615,N_8099);
or U12163 (N_12163,N_5625,N_9934);
nor U12164 (N_12164,N_5094,N_8046);
and U12165 (N_12165,N_7465,N_9489);
or U12166 (N_12166,N_6089,N_9747);
xnor U12167 (N_12167,N_8393,N_7177);
nand U12168 (N_12168,N_9054,N_8804);
and U12169 (N_12169,N_6127,N_5379);
or U12170 (N_12170,N_6785,N_5240);
nand U12171 (N_12171,N_8390,N_5202);
nand U12172 (N_12172,N_8295,N_8115);
xnor U12173 (N_12173,N_8051,N_5022);
and U12174 (N_12174,N_7521,N_5543);
nand U12175 (N_12175,N_7920,N_5904);
nor U12176 (N_12176,N_7316,N_9610);
or U12177 (N_12177,N_6878,N_5251);
nor U12178 (N_12178,N_5732,N_9015);
nor U12179 (N_12179,N_7752,N_5481);
nor U12180 (N_12180,N_6307,N_6097);
nor U12181 (N_12181,N_5296,N_7838);
nand U12182 (N_12182,N_6789,N_7331);
nor U12183 (N_12183,N_5654,N_9479);
xor U12184 (N_12184,N_9609,N_7281);
and U12185 (N_12185,N_6573,N_9511);
xor U12186 (N_12186,N_6312,N_7567);
nor U12187 (N_12187,N_6386,N_8371);
or U12188 (N_12188,N_7896,N_8510);
and U12189 (N_12189,N_5074,N_6609);
or U12190 (N_12190,N_5177,N_8486);
nand U12191 (N_12191,N_7146,N_8406);
xor U12192 (N_12192,N_9457,N_5479);
nand U12193 (N_12193,N_7346,N_9312);
nand U12194 (N_12194,N_8688,N_8024);
or U12195 (N_12195,N_8786,N_8638);
and U12196 (N_12196,N_7661,N_9084);
or U12197 (N_12197,N_9531,N_7653);
and U12198 (N_12198,N_8668,N_5071);
and U12199 (N_12199,N_6003,N_9855);
nand U12200 (N_12200,N_5345,N_6688);
or U12201 (N_12201,N_9156,N_5009);
nand U12202 (N_12202,N_5585,N_6839);
and U12203 (N_12203,N_9034,N_6865);
nand U12204 (N_12204,N_5250,N_5822);
nor U12205 (N_12205,N_8127,N_9002);
nand U12206 (N_12206,N_6149,N_7550);
and U12207 (N_12207,N_7584,N_9812);
xnor U12208 (N_12208,N_5957,N_6408);
nand U12209 (N_12209,N_6349,N_9085);
nor U12210 (N_12210,N_7612,N_7579);
xor U12211 (N_12211,N_7555,N_6369);
xnor U12212 (N_12212,N_7072,N_5838);
xnor U12213 (N_12213,N_5731,N_6493);
and U12214 (N_12214,N_7186,N_5225);
and U12215 (N_12215,N_8213,N_6915);
nor U12216 (N_12216,N_7936,N_7426);
nor U12217 (N_12217,N_7566,N_8196);
and U12218 (N_12218,N_6164,N_8697);
xnor U12219 (N_12219,N_9965,N_6875);
xor U12220 (N_12220,N_6247,N_5895);
or U12221 (N_12221,N_8403,N_8627);
nand U12222 (N_12222,N_6787,N_5813);
xnor U12223 (N_12223,N_6825,N_7553);
nand U12224 (N_12224,N_9646,N_8865);
or U12225 (N_12225,N_8586,N_9942);
xor U12226 (N_12226,N_8900,N_8237);
nand U12227 (N_12227,N_6544,N_6595);
nand U12228 (N_12228,N_6710,N_7149);
nand U12229 (N_12229,N_8238,N_6419);
or U12230 (N_12230,N_6582,N_8710);
xnor U12231 (N_12231,N_9434,N_8152);
nand U12232 (N_12232,N_5527,N_6347);
nand U12233 (N_12233,N_8455,N_7501);
nand U12234 (N_12234,N_5312,N_5754);
nand U12235 (N_12235,N_5728,N_8669);
and U12236 (N_12236,N_8322,N_6340);
or U12237 (N_12237,N_8683,N_6271);
or U12238 (N_12238,N_8488,N_7198);
and U12239 (N_12239,N_5135,N_8315);
nor U12240 (N_12240,N_8191,N_9754);
and U12241 (N_12241,N_5260,N_7151);
nand U12242 (N_12242,N_7106,N_7514);
or U12243 (N_12243,N_7961,N_7857);
or U12244 (N_12244,N_6008,N_7683);
or U12245 (N_12245,N_8853,N_7570);
xor U12246 (N_12246,N_9337,N_8889);
xor U12247 (N_12247,N_6041,N_6209);
nor U12248 (N_12248,N_9386,N_7340);
or U12249 (N_12249,N_8752,N_8918);
nor U12250 (N_12250,N_9270,N_5495);
nor U12251 (N_12251,N_5969,N_9036);
xnor U12252 (N_12252,N_8189,N_5467);
nor U12253 (N_12253,N_7016,N_8169);
or U12254 (N_12254,N_7621,N_9382);
nor U12255 (N_12255,N_6375,N_7037);
nand U12256 (N_12256,N_8546,N_9375);
or U12257 (N_12257,N_6836,N_6675);
and U12258 (N_12258,N_9003,N_7726);
nand U12259 (N_12259,N_7642,N_8807);
and U12260 (N_12260,N_6033,N_9180);
xor U12261 (N_12261,N_6444,N_5560);
and U12262 (N_12262,N_9313,N_5820);
xnor U12263 (N_12263,N_7840,N_7582);
xor U12264 (N_12264,N_7354,N_6474);
and U12265 (N_12265,N_5722,N_6413);
xnor U12266 (N_12266,N_7847,N_9697);
xor U12267 (N_12267,N_5179,N_6537);
xnor U12268 (N_12268,N_7599,N_7005);
nor U12269 (N_12269,N_9816,N_9899);
xor U12270 (N_12270,N_9620,N_5354);
nor U12271 (N_12271,N_5849,N_5405);
nor U12272 (N_12272,N_5487,N_5311);
and U12273 (N_12273,N_6786,N_8776);
or U12274 (N_12274,N_7996,N_8585);
nand U12275 (N_12275,N_7196,N_8877);
and U12276 (N_12276,N_8946,N_5736);
nor U12277 (N_12277,N_7267,N_8827);
and U12278 (N_12278,N_6810,N_9096);
nand U12279 (N_12279,N_5027,N_9171);
and U12280 (N_12280,N_9528,N_5302);
nand U12281 (N_12281,N_8109,N_7404);
and U12282 (N_12282,N_9370,N_7069);
nor U12283 (N_12283,N_9571,N_7510);
nor U12284 (N_12284,N_9748,N_5637);
nor U12285 (N_12285,N_5391,N_6818);
and U12286 (N_12286,N_7950,N_5309);
nand U12287 (N_12287,N_8300,N_5650);
xor U12288 (N_12288,N_9804,N_7940);
and U12289 (N_12289,N_8806,N_8027);
nor U12290 (N_12290,N_7952,N_6129);
xnor U12291 (N_12291,N_7845,N_8965);
nor U12292 (N_12292,N_8750,N_6481);
nand U12293 (N_12293,N_7900,N_7277);
nand U12294 (N_12294,N_9209,N_7906);
or U12295 (N_12295,N_8289,N_6086);
or U12296 (N_12296,N_6453,N_7240);
xnor U12297 (N_12297,N_7786,N_5692);
nor U12298 (N_12298,N_8296,N_8497);
xor U12299 (N_12299,N_7399,N_6708);
or U12300 (N_12300,N_7858,N_5295);
and U12301 (N_12301,N_9801,N_5195);
xor U12302 (N_12302,N_9244,N_9904);
or U12303 (N_12303,N_6816,N_6531);
or U12304 (N_12304,N_5281,N_7230);
nor U12305 (N_12305,N_8791,N_5128);
nand U12306 (N_12306,N_9282,N_9744);
nand U12307 (N_12307,N_9451,N_8164);
xnor U12308 (N_12308,N_9781,N_9950);
or U12309 (N_12309,N_7523,N_5896);
nand U12310 (N_12310,N_8512,N_6159);
xnor U12311 (N_12311,N_8278,N_7034);
xor U12312 (N_12312,N_9453,N_8153);
nor U12313 (N_12313,N_9460,N_8268);
nand U12314 (N_12314,N_8320,N_6486);
nor U12315 (N_12315,N_6337,N_9238);
or U12316 (N_12316,N_5603,N_7159);
and U12317 (N_12317,N_7887,N_5629);
nor U12318 (N_12318,N_5501,N_9108);
and U12319 (N_12319,N_5735,N_6510);
xor U12320 (N_12320,N_7964,N_7027);
xor U12321 (N_12321,N_6527,N_6268);
nand U12322 (N_12322,N_8270,N_6096);
and U12323 (N_12323,N_9991,N_5196);
nor U12324 (N_12324,N_5404,N_6536);
or U12325 (N_12325,N_8255,N_8583);
and U12326 (N_12326,N_5536,N_8731);
xor U12327 (N_12327,N_7762,N_5455);
xor U12328 (N_12328,N_9642,N_8040);
xor U12329 (N_12329,N_9043,N_7459);
nor U12330 (N_12330,N_7079,N_8228);
nor U12331 (N_12331,N_9989,N_5621);
nand U12332 (N_12332,N_8130,N_6425);
or U12333 (N_12333,N_9714,N_7813);
or U12334 (N_12334,N_9968,N_8764);
or U12335 (N_12335,N_7128,N_9736);
or U12336 (N_12336,N_5815,N_8192);
nor U12337 (N_12337,N_7730,N_7130);
xor U12338 (N_12338,N_8096,N_6443);
nor U12339 (N_12339,N_8640,N_6617);
nor U12340 (N_12340,N_9915,N_6779);
nor U12341 (N_12341,N_9923,N_6828);
and U12342 (N_12342,N_8529,N_7722);
nand U12343 (N_12343,N_7036,N_6974);
and U12344 (N_12344,N_5848,N_5219);
nor U12345 (N_12345,N_5755,N_7261);
nand U12346 (N_12346,N_5381,N_9683);
xor U12347 (N_12347,N_7827,N_6952);
xor U12348 (N_12348,N_5690,N_7476);
and U12349 (N_12349,N_9051,N_7310);
nor U12350 (N_12350,N_8863,N_5956);
and U12351 (N_12351,N_8605,N_9038);
and U12352 (N_12352,N_9217,N_9705);
nor U12353 (N_12353,N_6441,N_7448);
xor U12354 (N_12354,N_6139,N_9110);
and U12355 (N_12355,N_6806,N_9924);
xnor U12356 (N_12356,N_7353,N_7591);
and U12357 (N_12357,N_6136,N_9759);
or U12358 (N_12358,N_7094,N_6073);
or U12359 (N_12359,N_6487,N_5396);
or U12360 (N_12360,N_5937,N_9378);
or U12361 (N_12361,N_7571,N_8310);
xnor U12362 (N_12362,N_6135,N_5710);
nor U12363 (N_12363,N_8276,N_8174);
nor U12364 (N_12364,N_5470,N_8716);
or U12365 (N_12365,N_6512,N_9560);
and U12366 (N_12366,N_8992,N_5984);
and U12367 (N_12367,N_6522,N_5947);
xnor U12368 (N_12368,N_7167,N_5539);
and U12369 (N_12369,N_6777,N_5214);
nand U12370 (N_12370,N_5668,N_8567);
nor U12371 (N_12371,N_9144,N_6121);
nor U12372 (N_12372,N_7215,N_9330);
nor U12373 (N_12373,N_8036,N_8736);
nand U12374 (N_12374,N_8582,N_9719);
xor U12375 (N_12375,N_6274,N_5767);
or U12376 (N_12376,N_7798,N_7558);
and U12377 (N_12377,N_7400,N_9502);
nor U12378 (N_12378,N_5551,N_5163);
xnor U12379 (N_12379,N_9010,N_8037);
or U12380 (N_12380,N_6953,N_8597);
or U12381 (N_12381,N_8373,N_6966);
or U12382 (N_12382,N_6276,N_5823);
xnor U12383 (N_12383,N_9065,N_8571);
nand U12384 (N_12384,N_7781,N_6624);
nand U12385 (N_12385,N_9912,N_6903);
nand U12386 (N_12386,N_9247,N_9202);
xnor U12387 (N_12387,N_8275,N_9718);
xnor U12388 (N_12388,N_9783,N_9712);
nor U12389 (N_12389,N_7815,N_6367);
nor U12390 (N_12390,N_8975,N_5859);
and U12391 (N_12391,N_8606,N_7490);
nand U12392 (N_12392,N_6501,N_7842);
nand U12393 (N_12393,N_8325,N_9808);
nor U12394 (N_12394,N_5112,N_8958);
nor U12395 (N_12395,N_5081,N_6321);
or U12396 (N_12396,N_5592,N_7513);
and U12397 (N_12397,N_6668,N_6252);
nand U12398 (N_12398,N_9461,N_8471);
nor U12399 (N_12399,N_6687,N_9291);
xnor U12400 (N_12400,N_8648,N_5035);
or U12401 (N_12401,N_6987,N_8015);
nor U12402 (N_12402,N_8935,N_5222);
xnor U12403 (N_12403,N_9431,N_9464);
and U12404 (N_12404,N_8558,N_7189);
and U12405 (N_12405,N_5137,N_8399);
or U12406 (N_12406,N_9691,N_6417);
xnor U12407 (N_12407,N_5406,N_7117);
nor U12408 (N_12408,N_6697,N_9635);
nand U12409 (N_12409,N_8058,N_9840);
nand U12410 (N_12410,N_6286,N_8297);
xnor U12411 (N_12411,N_9402,N_7775);
or U12412 (N_12412,N_9664,N_9740);
xnor U12413 (N_12413,N_8869,N_8618);
and U12414 (N_12414,N_5887,N_7728);
and U12415 (N_12415,N_5649,N_9798);
nand U12416 (N_12416,N_6288,N_8410);
nor U12417 (N_12417,N_9081,N_9681);
xor U12418 (N_12418,N_7019,N_5398);
nand U12419 (N_12419,N_7048,N_9494);
nor U12420 (N_12420,N_9514,N_6528);
nor U12421 (N_12421,N_5744,N_7479);
xor U12422 (N_12422,N_8796,N_8705);
nand U12423 (N_12423,N_9819,N_8612);
or U12424 (N_12424,N_5263,N_7129);
or U12425 (N_12425,N_5810,N_7863);
and U12426 (N_12426,N_6893,N_6355);
xnor U12427 (N_12427,N_9172,N_5105);
xnor U12428 (N_12428,N_5315,N_8031);
nor U12429 (N_12429,N_5505,N_8392);
and U12430 (N_12430,N_8477,N_9711);
and U12431 (N_12431,N_5502,N_5780);
nor U12432 (N_12432,N_6737,N_6154);
and U12433 (N_12433,N_5622,N_9234);
xor U12434 (N_12434,N_9060,N_5967);
and U12435 (N_12435,N_7765,N_7867);
xor U12436 (N_12436,N_6577,N_7279);
and U12437 (N_12437,N_7341,N_9752);
nand U12438 (N_12438,N_5831,N_8362);
nor U12439 (N_12439,N_5784,N_9799);
xor U12440 (N_12440,N_5870,N_5959);
and U12441 (N_12441,N_6057,N_7701);
nand U12442 (N_12442,N_7220,N_6815);
and U12443 (N_12443,N_6727,N_7370);
and U12444 (N_12444,N_8081,N_6770);
xnor U12445 (N_12445,N_6794,N_7009);
xnor U12446 (N_12446,N_6649,N_9097);
xor U12447 (N_12447,N_6422,N_8453);
nor U12448 (N_12448,N_8063,N_9793);
nor U12449 (N_12449,N_8819,N_5026);
and U12450 (N_12450,N_6603,N_5110);
xnor U12451 (N_12451,N_9811,N_8733);
xnor U12452 (N_12452,N_9186,N_6928);
nand U12453 (N_12453,N_5908,N_7601);
or U12454 (N_12454,N_9371,N_8142);
xnor U12455 (N_12455,N_7605,N_7533);
xnor U12456 (N_12456,N_5082,N_7384);
and U12457 (N_12457,N_6282,N_5955);
xnor U12458 (N_12458,N_8506,N_9562);
xor U12459 (N_12459,N_6886,N_5330);
nand U12460 (N_12460,N_7524,N_7115);
xnor U12461 (N_12461,N_7049,N_6655);
and U12462 (N_12462,N_8987,N_9931);
nor U12463 (N_12463,N_7625,N_8757);
and U12464 (N_12464,N_6426,N_7416);
nor U12465 (N_12465,N_6982,N_5510);
and U12466 (N_12466,N_7659,N_5159);
and U12467 (N_12467,N_7552,N_9443);
nand U12468 (N_12468,N_5261,N_9357);
and U12469 (N_12469,N_9990,N_7573);
and U12470 (N_12470,N_5013,N_7452);
nand U12471 (N_12471,N_7885,N_7837);
and U12472 (N_12472,N_9568,N_9786);
nor U12473 (N_12473,N_9027,N_5386);
or U12474 (N_12474,N_5364,N_7682);
nor U12475 (N_12475,N_9049,N_6212);
xnor U12476 (N_12476,N_9557,N_8009);
xnor U12477 (N_12477,N_6631,N_8623);
or U12478 (N_12478,N_8489,N_7734);
and U12479 (N_12479,N_6936,N_6430);
and U12480 (N_12480,N_6713,N_5706);
nand U12481 (N_12481,N_6672,N_6037);
nor U12482 (N_12482,N_6112,N_8751);
or U12483 (N_12483,N_9221,N_7874);
nor U12484 (N_12484,N_9449,N_5804);
nand U12485 (N_12485,N_5862,N_9701);
xnor U12486 (N_12486,N_6175,N_8227);
and U12487 (N_12487,N_5224,N_9680);
xor U12488 (N_12488,N_9507,N_6860);
xor U12489 (N_12489,N_7201,N_5076);
nand U12490 (N_12490,N_5730,N_6561);
nand U12491 (N_12491,N_6533,N_6372);
and U12492 (N_12492,N_5857,N_5995);
and U12493 (N_12493,N_6289,N_7474);
and U12494 (N_12494,N_9351,N_6389);
nor U12495 (N_12495,N_5828,N_8429);
xnor U12496 (N_12496,N_5016,N_7951);
nand U12497 (N_12497,N_9998,N_9018);
and U12498 (N_12498,N_8902,N_6219);
nor U12499 (N_12499,N_8928,N_8201);
nand U12500 (N_12500,N_9564,N_6322);
or U12501 (N_12501,N_6809,N_5173);
nor U12502 (N_12502,N_8207,N_8768);
nor U12503 (N_12503,N_6010,N_6114);
nand U12504 (N_12504,N_6298,N_7466);
nor U12505 (N_12505,N_9112,N_8572);
and U12506 (N_12506,N_7138,N_7426);
or U12507 (N_12507,N_7714,N_5249);
nor U12508 (N_12508,N_5179,N_8584);
nand U12509 (N_12509,N_9310,N_8920);
xor U12510 (N_12510,N_7795,N_5833);
xor U12511 (N_12511,N_8856,N_8450);
xor U12512 (N_12512,N_9871,N_5215);
and U12513 (N_12513,N_6761,N_6781);
nand U12514 (N_12514,N_6681,N_9094);
nand U12515 (N_12515,N_9321,N_8774);
nand U12516 (N_12516,N_5206,N_7347);
nand U12517 (N_12517,N_6651,N_5370);
xor U12518 (N_12518,N_6038,N_7317);
xnor U12519 (N_12519,N_8946,N_7769);
xor U12520 (N_12520,N_5784,N_5462);
and U12521 (N_12521,N_9191,N_5890);
nor U12522 (N_12522,N_7348,N_7180);
nand U12523 (N_12523,N_9477,N_6945);
xnor U12524 (N_12524,N_5524,N_7436);
nand U12525 (N_12525,N_9278,N_9321);
xor U12526 (N_12526,N_7288,N_5721);
xor U12527 (N_12527,N_7879,N_6914);
nor U12528 (N_12528,N_6656,N_8719);
nand U12529 (N_12529,N_5391,N_7786);
nand U12530 (N_12530,N_8762,N_6911);
or U12531 (N_12531,N_7439,N_7650);
or U12532 (N_12532,N_9359,N_5531);
and U12533 (N_12533,N_9994,N_5929);
xnor U12534 (N_12534,N_5712,N_6806);
nand U12535 (N_12535,N_5475,N_6668);
nor U12536 (N_12536,N_5589,N_9746);
xnor U12537 (N_12537,N_8240,N_5554);
nor U12538 (N_12538,N_7124,N_7426);
nor U12539 (N_12539,N_7587,N_6924);
xnor U12540 (N_12540,N_6758,N_8277);
or U12541 (N_12541,N_8433,N_7552);
or U12542 (N_12542,N_5447,N_7744);
or U12543 (N_12543,N_9248,N_5856);
xnor U12544 (N_12544,N_6459,N_7883);
and U12545 (N_12545,N_7421,N_7914);
or U12546 (N_12546,N_5032,N_8047);
and U12547 (N_12547,N_7008,N_5481);
xor U12548 (N_12548,N_5300,N_8167);
nand U12549 (N_12549,N_6254,N_6613);
and U12550 (N_12550,N_9257,N_7478);
xnor U12551 (N_12551,N_5496,N_8607);
and U12552 (N_12552,N_7751,N_7598);
nand U12553 (N_12553,N_7392,N_6586);
xor U12554 (N_12554,N_5790,N_8345);
nand U12555 (N_12555,N_8341,N_6497);
nor U12556 (N_12556,N_9591,N_5365);
nand U12557 (N_12557,N_8511,N_8987);
or U12558 (N_12558,N_9477,N_9737);
xor U12559 (N_12559,N_6667,N_8584);
or U12560 (N_12560,N_9145,N_5786);
nor U12561 (N_12561,N_8143,N_5289);
or U12562 (N_12562,N_7676,N_6378);
nand U12563 (N_12563,N_6500,N_9962);
nand U12564 (N_12564,N_9002,N_8758);
nor U12565 (N_12565,N_6478,N_8521);
xor U12566 (N_12566,N_9921,N_8719);
or U12567 (N_12567,N_7682,N_8763);
xnor U12568 (N_12568,N_7617,N_7920);
xnor U12569 (N_12569,N_7010,N_8084);
and U12570 (N_12570,N_8421,N_7630);
or U12571 (N_12571,N_9442,N_7379);
or U12572 (N_12572,N_6313,N_8324);
or U12573 (N_12573,N_7440,N_5451);
nand U12574 (N_12574,N_6484,N_5924);
xor U12575 (N_12575,N_7734,N_8082);
and U12576 (N_12576,N_7477,N_7106);
and U12577 (N_12577,N_5265,N_7290);
nor U12578 (N_12578,N_7842,N_9479);
or U12579 (N_12579,N_9031,N_7446);
and U12580 (N_12580,N_9473,N_6430);
nor U12581 (N_12581,N_9968,N_8654);
xor U12582 (N_12582,N_9675,N_7321);
xor U12583 (N_12583,N_7093,N_5096);
or U12584 (N_12584,N_8937,N_6417);
nand U12585 (N_12585,N_7773,N_7996);
nor U12586 (N_12586,N_9274,N_8358);
xor U12587 (N_12587,N_6688,N_6289);
nor U12588 (N_12588,N_5228,N_9006);
nand U12589 (N_12589,N_9423,N_9850);
nor U12590 (N_12590,N_9784,N_6884);
and U12591 (N_12591,N_9617,N_7657);
nand U12592 (N_12592,N_9166,N_9753);
or U12593 (N_12593,N_7936,N_7243);
or U12594 (N_12594,N_7166,N_5033);
nor U12595 (N_12595,N_7115,N_6294);
and U12596 (N_12596,N_9684,N_7405);
or U12597 (N_12597,N_5257,N_9781);
and U12598 (N_12598,N_5261,N_7744);
and U12599 (N_12599,N_5284,N_8049);
nor U12600 (N_12600,N_7285,N_6757);
or U12601 (N_12601,N_8429,N_8408);
xnor U12602 (N_12602,N_8103,N_7472);
or U12603 (N_12603,N_9763,N_9912);
and U12604 (N_12604,N_5035,N_5404);
nand U12605 (N_12605,N_7678,N_9994);
nor U12606 (N_12606,N_7334,N_6701);
and U12607 (N_12607,N_7873,N_8995);
nand U12608 (N_12608,N_9964,N_7886);
and U12609 (N_12609,N_7152,N_5541);
and U12610 (N_12610,N_9849,N_8802);
or U12611 (N_12611,N_6696,N_8503);
nand U12612 (N_12612,N_8738,N_5172);
xor U12613 (N_12613,N_8159,N_5978);
xnor U12614 (N_12614,N_5189,N_7115);
or U12615 (N_12615,N_5175,N_8191);
and U12616 (N_12616,N_9503,N_6014);
and U12617 (N_12617,N_8645,N_6450);
nor U12618 (N_12618,N_7048,N_5463);
xnor U12619 (N_12619,N_7025,N_6802);
nor U12620 (N_12620,N_7728,N_8970);
xnor U12621 (N_12621,N_5046,N_7216);
and U12622 (N_12622,N_5666,N_7914);
nand U12623 (N_12623,N_5197,N_9611);
nand U12624 (N_12624,N_7983,N_9549);
xor U12625 (N_12625,N_8138,N_7422);
xor U12626 (N_12626,N_6947,N_6212);
and U12627 (N_12627,N_7226,N_7006);
and U12628 (N_12628,N_5593,N_8477);
and U12629 (N_12629,N_6169,N_7344);
nand U12630 (N_12630,N_8317,N_9532);
and U12631 (N_12631,N_9737,N_8729);
and U12632 (N_12632,N_5865,N_8305);
nor U12633 (N_12633,N_8424,N_9033);
and U12634 (N_12634,N_8612,N_9454);
nor U12635 (N_12635,N_9581,N_5610);
xnor U12636 (N_12636,N_5079,N_5920);
or U12637 (N_12637,N_6248,N_7630);
nand U12638 (N_12638,N_5571,N_5419);
and U12639 (N_12639,N_8753,N_8124);
or U12640 (N_12640,N_8431,N_6674);
nand U12641 (N_12641,N_5486,N_5591);
nor U12642 (N_12642,N_7561,N_6526);
and U12643 (N_12643,N_5707,N_6254);
nand U12644 (N_12644,N_8886,N_6177);
or U12645 (N_12645,N_7943,N_7789);
or U12646 (N_12646,N_6623,N_8078);
or U12647 (N_12647,N_7758,N_7272);
and U12648 (N_12648,N_6441,N_6058);
xnor U12649 (N_12649,N_7872,N_9880);
and U12650 (N_12650,N_5378,N_6358);
or U12651 (N_12651,N_8613,N_6924);
nor U12652 (N_12652,N_9708,N_9749);
xnor U12653 (N_12653,N_7766,N_7523);
or U12654 (N_12654,N_5827,N_8355);
or U12655 (N_12655,N_9149,N_6186);
and U12656 (N_12656,N_7695,N_5786);
nor U12657 (N_12657,N_5590,N_5054);
and U12658 (N_12658,N_5236,N_5654);
nor U12659 (N_12659,N_8055,N_6941);
and U12660 (N_12660,N_6711,N_8409);
or U12661 (N_12661,N_8265,N_7433);
or U12662 (N_12662,N_8247,N_6246);
and U12663 (N_12663,N_7299,N_5183);
or U12664 (N_12664,N_5447,N_7030);
xor U12665 (N_12665,N_8686,N_6041);
or U12666 (N_12666,N_5457,N_5641);
or U12667 (N_12667,N_6274,N_7294);
xnor U12668 (N_12668,N_7238,N_7557);
nand U12669 (N_12669,N_5201,N_6301);
and U12670 (N_12670,N_8027,N_9867);
nor U12671 (N_12671,N_9453,N_6631);
nor U12672 (N_12672,N_5540,N_9174);
xnor U12673 (N_12673,N_7090,N_5813);
xnor U12674 (N_12674,N_6502,N_5438);
and U12675 (N_12675,N_5527,N_8291);
nor U12676 (N_12676,N_5243,N_7965);
nor U12677 (N_12677,N_5381,N_8291);
or U12678 (N_12678,N_6472,N_9307);
and U12679 (N_12679,N_7870,N_5198);
or U12680 (N_12680,N_8404,N_7246);
nor U12681 (N_12681,N_6958,N_7921);
xnor U12682 (N_12682,N_9252,N_9858);
and U12683 (N_12683,N_9473,N_5819);
or U12684 (N_12684,N_6604,N_8227);
nor U12685 (N_12685,N_9095,N_5955);
or U12686 (N_12686,N_7754,N_7752);
and U12687 (N_12687,N_7001,N_8646);
nor U12688 (N_12688,N_6794,N_8105);
nand U12689 (N_12689,N_7901,N_7802);
xor U12690 (N_12690,N_9436,N_9657);
or U12691 (N_12691,N_6951,N_9101);
nand U12692 (N_12692,N_6485,N_7837);
xor U12693 (N_12693,N_9486,N_9995);
xnor U12694 (N_12694,N_8481,N_9287);
nand U12695 (N_12695,N_7360,N_9322);
nor U12696 (N_12696,N_6415,N_8201);
nor U12697 (N_12697,N_7575,N_8681);
and U12698 (N_12698,N_5643,N_7152);
and U12699 (N_12699,N_8740,N_6625);
xor U12700 (N_12700,N_8523,N_5384);
nor U12701 (N_12701,N_8692,N_8507);
nor U12702 (N_12702,N_7710,N_6724);
and U12703 (N_12703,N_8437,N_7577);
nor U12704 (N_12704,N_7653,N_6984);
and U12705 (N_12705,N_5899,N_6175);
nor U12706 (N_12706,N_9302,N_7821);
xor U12707 (N_12707,N_7024,N_7087);
nand U12708 (N_12708,N_8515,N_9409);
and U12709 (N_12709,N_9716,N_5922);
nor U12710 (N_12710,N_6262,N_5433);
and U12711 (N_12711,N_9461,N_6654);
and U12712 (N_12712,N_7233,N_6721);
nor U12713 (N_12713,N_8896,N_5906);
nor U12714 (N_12714,N_8299,N_5585);
nor U12715 (N_12715,N_6327,N_7104);
and U12716 (N_12716,N_9979,N_5991);
and U12717 (N_12717,N_8869,N_7822);
nor U12718 (N_12718,N_5843,N_6721);
xnor U12719 (N_12719,N_5920,N_8807);
xnor U12720 (N_12720,N_8245,N_8531);
nor U12721 (N_12721,N_8835,N_6287);
nand U12722 (N_12722,N_8731,N_9453);
and U12723 (N_12723,N_5068,N_8423);
nand U12724 (N_12724,N_9245,N_5017);
nand U12725 (N_12725,N_5130,N_8345);
and U12726 (N_12726,N_7159,N_6229);
xor U12727 (N_12727,N_5775,N_8096);
xor U12728 (N_12728,N_6001,N_5028);
and U12729 (N_12729,N_6329,N_5203);
nor U12730 (N_12730,N_8099,N_8960);
xnor U12731 (N_12731,N_9858,N_8347);
nor U12732 (N_12732,N_5064,N_8652);
xor U12733 (N_12733,N_7162,N_8406);
or U12734 (N_12734,N_7369,N_7638);
or U12735 (N_12735,N_9111,N_6061);
and U12736 (N_12736,N_7126,N_8111);
and U12737 (N_12737,N_6350,N_7871);
nand U12738 (N_12738,N_6920,N_5549);
and U12739 (N_12739,N_8556,N_6624);
and U12740 (N_12740,N_5068,N_5978);
xnor U12741 (N_12741,N_9010,N_6293);
nand U12742 (N_12742,N_5468,N_9479);
nand U12743 (N_12743,N_7149,N_9921);
or U12744 (N_12744,N_6742,N_8416);
or U12745 (N_12745,N_7974,N_8973);
xor U12746 (N_12746,N_7535,N_6007);
and U12747 (N_12747,N_8633,N_8586);
or U12748 (N_12748,N_5197,N_9670);
nor U12749 (N_12749,N_7090,N_8891);
or U12750 (N_12750,N_7395,N_5454);
xnor U12751 (N_12751,N_8580,N_7543);
or U12752 (N_12752,N_9101,N_9269);
or U12753 (N_12753,N_5769,N_6925);
xnor U12754 (N_12754,N_9800,N_5228);
xnor U12755 (N_12755,N_9225,N_5708);
or U12756 (N_12756,N_6498,N_5706);
or U12757 (N_12757,N_9947,N_9719);
or U12758 (N_12758,N_7779,N_8157);
nor U12759 (N_12759,N_7262,N_7564);
or U12760 (N_12760,N_9026,N_7714);
or U12761 (N_12761,N_9727,N_8019);
nor U12762 (N_12762,N_7327,N_8128);
and U12763 (N_12763,N_9345,N_7891);
xnor U12764 (N_12764,N_6760,N_6979);
xnor U12765 (N_12765,N_5906,N_9679);
and U12766 (N_12766,N_9183,N_5433);
nand U12767 (N_12767,N_6877,N_6726);
nor U12768 (N_12768,N_8137,N_5795);
nor U12769 (N_12769,N_7132,N_5090);
nor U12770 (N_12770,N_8365,N_6012);
xnor U12771 (N_12771,N_6629,N_9417);
or U12772 (N_12772,N_8416,N_7187);
nor U12773 (N_12773,N_5874,N_6669);
and U12774 (N_12774,N_8065,N_5256);
and U12775 (N_12775,N_6823,N_8762);
nand U12776 (N_12776,N_7435,N_9401);
and U12777 (N_12777,N_5240,N_5278);
and U12778 (N_12778,N_8320,N_9642);
and U12779 (N_12779,N_9706,N_9991);
or U12780 (N_12780,N_6125,N_5988);
and U12781 (N_12781,N_7444,N_6342);
and U12782 (N_12782,N_9647,N_5083);
and U12783 (N_12783,N_5273,N_5256);
nand U12784 (N_12784,N_7124,N_6186);
or U12785 (N_12785,N_9413,N_6787);
and U12786 (N_12786,N_9235,N_5535);
and U12787 (N_12787,N_7401,N_6546);
xnor U12788 (N_12788,N_7073,N_9419);
nor U12789 (N_12789,N_9469,N_9129);
nor U12790 (N_12790,N_8238,N_5903);
or U12791 (N_12791,N_8900,N_7218);
nor U12792 (N_12792,N_6360,N_7536);
nor U12793 (N_12793,N_7510,N_8702);
nor U12794 (N_12794,N_9057,N_8360);
nor U12795 (N_12795,N_9380,N_9182);
xnor U12796 (N_12796,N_5804,N_9494);
nor U12797 (N_12797,N_9690,N_6488);
nand U12798 (N_12798,N_9677,N_6608);
and U12799 (N_12799,N_6659,N_8656);
and U12800 (N_12800,N_5666,N_8550);
and U12801 (N_12801,N_5983,N_6513);
and U12802 (N_12802,N_7429,N_9027);
nor U12803 (N_12803,N_7639,N_8612);
nor U12804 (N_12804,N_9581,N_9666);
or U12805 (N_12805,N_8128,N_8626);
nand U12806 (N_12806,N_8545,N_5024);
nor U12807 (N_12807,N_6359,N_7549);
nor U12808 (N_12808,N_7638,N_9382);
nand U12809 (N_12809,N_8376,N_8681);
xor U12810 (N_12810,N_9776,N_9778);
and U12811 (N_12811,N_8881,N_8691);
or U12812 (N_12812,N_9411,N_6294);
nor U12813 (N_12813,N_7568,N_8743);
or U12814 (N_12814,N_7102,N_9687);
xor U12815 (N_12815,N_5325,N_8512);
xor U12816 (N_12816,N_8371,N_5115);
nand U12817 (N_12817,N_6589,N_7647);
or U12818 (N_12818,N_9699,N_8301);
xor U12819 (N_12819,N_8206,N_8897);
xor U12820 (N_12820,N_5639,N_9266);
or U12821 (N_12821,N_9990,N_8357);
nand U12822 (N_12822,N_7934,N_6285);
nand U12823 (N_12823,N_9754,N_8956);
xnor U12824 (N_12824,N_5298,N_5195);
and U12825 (N_12825,N_6030,N_8561);
and U12826 (N_12826,N_9720,N_9946);
and U12827 (N_12827,N_5067,N_7600);
nand U12828 (N_12828,N_7083,N_5839);
or U12829 (N_12829,N_7578,N_5959);
nand U12830 (N_12830,N_9605,N_7428);
and U12831 (N_12831,N_6372,N_8748);
xor U12832 (N_12832,N_9222,N_6228);
and U12833 (N_12833,N_8520,N_5794);
and U12834 (N_12834,N_8683,N_9754);
and U12835 (N_12835,N_7895,N_7463);
xnor U12836 (N_12836,N_5583,N_7553);
xor U12837 (N_12837,N_5033,N_7234);
xnor U12838 (N_12838,N_7252,N_9175);
and U12839 (N_12839,N_9730,N_6616);
or U12840 (N_12840,N_9445,N_8537);
nand U12841 (N_12841,N_8204,N_8632);
xor U12842 (N_12842,N_9972,N_5270);
xor U12843 (N_12843,N_5105,N_6459);
or U12844 (N_12844,N_7459,N_7437);
nand U12845 (N_12845,N_5859,N_6548);
xor U12846 (N_12846,N_7424,N_9812);
or U12847 (N_12847,N_6771,N_8735);
and U12848 (N_12848,N_8386,N_8949);
or U12849 (N_12849,N_9038,N_6838);
or U12850 (N_12850,N_8787,N_8060);
nor U12851 (N_12851,N_6883,N_9261);
xnor U12852 (N_12852,N_7562,N_8515);
and U12853 (N_12853,N_9007,N_5935);
and U12854 (N_12854,N_5803,N_5504);
xnor U12855 (N_12855,N_7540,N_6851);
or U12856 (N_12856,N_9254,N_8383);
and U12857 (N_12857,N_6668,N_6776);
nand U12858 (N_12858,N_5391,N_8868);
nand U12859 (N_12859,N_9829,N_6873);
and U12860 (N_12860,N_8326,N_6155);
xnor U12861 (N_12861,N_8851,N_9345);
or U12862 (N_12862,N_5539,N_5472);
or U12863 (N_12863,N_9845,N_5121);
and U12864 (N_12864,N_6948,N_7703);
xor U12865 (N_12865,N_8364,N_7450);
or U12866 (N_12866,N_9728,N_6828);
nand U12867 (N_12867,N_7976,N_6637);
nor U12868 (N_12868,N_7441,N_9965);
nand U12869 (N_12869,N_8591,N_5999);
xnor U12870 (N_12870,N_6492,N_7549);
nor U12871 (N_12871,N_9175,N_7972);
and U12872 (N_12872,N_6696,N_9337);
xor U12873 (N_12873,N_8908,N_5903);
nand U12874 (N_12874,N_9174,N_8313);
nor U12875 (N_12875,N_6058,N_7508);
xnor U12876 (N_12876,N_9803,N_6067);
or U12877 (N_12877,N_8123,N_8696);
or U12878 (N_12878,N_8341,N_8459);
xor U12879 (N_12879,N_5666,N_9319);
or U12880 (N_12880,N_6149,N_6558);
xnor U12881 (N_12881,N_6878,N_8043);
or U12882 (N_12882,N_9836,N_5054);
nor U12883 (N_12883,N_5153,N_5510);
nor U12884 (N_12884,N_9712,N_8948);
and U12885 (N_12885,N_5923,N_8960);
nand U12886 (N_12886,N_6535,N_9799);
xor U12887 (N_12887,N_6059,N_7361);
xnor U12888 (N_12888,N_9938,N_6716);
and U12889 (N_12889,N_8539,N_8591);
or U12890 (N_12890,N_9403,N_5610);
nand U12891 (N_12891,N_6620,N_7606);
nor U12892 (N_12892,N_9064,N_7591);
xor U12893 (N_12893,N_5697,N_7591);
nor U12894 (N_12894,N_5373,N_6789);
and U12895 (N_12895,N_5557,N_9342);
nor U12896 (N_12896,N_7583,N_7600);
nor U12897 (N_12897,N_7174,N_6246);
nand U12898 (N_12898,N_8408,N_5087);
xor U12899 (N_12899,N_8012,N_9477);
and U12900 (N_12900,N_6042,N_6812);
nor U12901 (N_12901,N_7084,N_8318);
or U12902 (N_12902,N_5719,N_6031);
nor U12903 (N_12903,N_9182,N_6009);
nand U12904 (N_12904,N_8400,N_9779);
nor U12905 (N_12905,N_6752,N_7587);
nor U12906 (N_12906,N_8497,N_8275);
nor U12907 (N_12907,N_5430,N_6046);
or U12908 (N_12908,N_9186,N_7312);
and U12909 (N_12909,N_6684,N_6249);
nand U12910 (N_12910,N_9104,N_8279);
nor U12911 (N_12911,N_5269,N_7291);
and U12912 (N_12912,N_8696,N_8012);
and U12913 (N_12913,N_8775,N_9396);
or U12914 (N_12914,N_8127,N_6934);
xor U12915 (N_12915,N_5722,N_6254);
or U12916 (N_12916,N_8920,N_7821);
nand U12917 (N_12917,N_5136,N_5376);
or U12918 (N_12918,N_9600,N_7102);
or U12919 (N_12919,N_5342,N_5823);
or U12920 (N_12920,N_9033,N_8400);
and U12921 (N_12921,N_9296,N_8491);
and U12922 (N_12922,N_6129,N_8532);
or U12923 (N_12923,N_5355,N_6185);
or U12924 (N_12924,N_5964,N_7559);
nor U12925 (N_12925,N_7477,N_6437);
nor U12926 (N_12926,N_6972,N_8738);
nand U12927 (N_12927,N_5863,N_8857);
or U12928 (N_12928,N_6300,N_7073);
nand U12929 (N_12929,N_9324,N_8736);
nand U12930 (N_12930,N_9237,N_8221);
or U12931 (N_12931,N_9549,N_6984);
and U12932 (N_12932,N_7555,N_5991);
and U12933 (N_12933,N_5095,N_6199);
or U12934 (N_12934,N_7918,N_6305);
nand U12935 (N_12935,N_6198,N_7862);
nor U12936 (N_12936,N_6306,N_6779);
nand U12937 (N_12937,N_7779,N_6740);
xnor U12938 (N_12938,N_9368,N_8954);
xnor U12939 (N_12939,N_7510,N_6024);
nor U12940 (N_12940,N_9296,N_6099);
nor U12941 (N_12941,N_9370,N_5624);
and U12942 (N_12942,N_6410,N_9449);
or U12943 (N_12943,N_6876,N_9057);
and U12944 (N_12944,N_6525,N_6976);
nor U12945 (N_12945,N_6708,N_5076);
nor U12946 (N_12946,N_8247,N_7869);
nor U12947 (N_12947,N_5220,N_7033);
or U12948 (N_12948,N_5571,N_7509);
xor U12949 (N_12949,N_7136,N_7727);
nor U12950 (N_12950,N_5263,N_6793);
xor U12951 (N_12951,N_8817,N_6471);
xnor U12952 (N_12952,N_5905,N_7397);
nor U12953 (N_12953,N_8182,N_9089);
xor U12954 (N_12954,N_5094,N_9230);
nor U12955 (N_12955,N_7000,N_8434);
nor U12956 (N_12956,N_6330,N_6694);
xor U12957 (N_12957,N_8247,N_6652);
xnor U12958 (N_12958,N_6561,N_7941);
nand U12959 (N_12959,N_8860,N_7043);
xnor U12960 (N_12960,N_9523,N_7191);
or U12961 (N_12961,N_6203,N_8725);
nand U12962 (N_12962,N_6786,N_6273);
nor U12963 (N_12963,N_5014,N_8897);
nor U12964 (N_12964,N_5667,N_5879);
and U12965 (N_12965,N_7461,N_8285);
nor U12966 (N_12966,N_6868,N_5882);
and U12967 (N_12967,N_7873,N_5361);
or U12968 (N_12968,N_5547,N_7748);
nor U12969 (N_12969,N_5156,N_5913);
and U12970 (N_12970,N_7320,N_7893);
and U12971 (N_12971,N_7134,N_9790);
or U12972 (N_12972,N_9263,N_9740);
nor U12973 (N_12973,N_8657,N_5843);
or U12974 (N_12974,N_5129,N_7539);
or U12975 (N_12975,N_7414,N_8705);
nand U12976 (N_12976,N_9891,N_9350);
nor U12977 (N_12977,N_6757,N_8176);
nand U12978 (N_12978,N_7558,N_9646);
nor U12979 (N_12979,N_8893,N_8419);
xor U12980 (N_12980,N_7088,N_6041);
nand U12981 (N_12981,N_6645,N_5695);
and U12982 (N_12982,N_7970,N_9162);
nand U12983 (N_12983,N_6133,N_9449);
nor U12984 (N_12984,N_6605,N_9228);
or U12985 (N_12985,N_9571,N_7766);
nor U12986 (N_12986,N_6990,N_6981);
xor U12987 (N_12987,N_5379,N_9672);
nor U12988 (N_12988,N_6590,N_7951);
nand U12989 (N_12989,N_6812,N_5539);
and U12990 (N_12990,N_5543,N_5731);
nor U12991 (N_12991,N_6348,N_7669);
nor U12992 (N_12992,N_6239,N_8410);
nand U12993 (N_12993,N_9740,N_9891);
nand U12994 (N_12994,N_5883,N_5056);
and U12995 (N_12995,N_7215,N_5936);
or U12996 (N_12996,N_6187,N_7880);
and U12997 (N_12997,N_6532,N_9507);
xor U12998 (N_12998,N_7328,N_7295);
and U12999 (N_12999,N_6507,N_9312);
nand U13000 (N_13000,N_6138,N_7096);
and U13001 (N_13001,N_9708,N_5975);
nand U13002 (N_13002,N_5535,N_8376);
or U13003 (N_13003,N_7446,N_7078);
or U13004 (N_13004,N_6930,N_7665);
and U13005 (N_13005,N_6541,N_6581);
and U13006 (N_13006,N_8071,N_6697);
nand U13007 (N_13007,N_8794,N_6995);
nor U13008 (N_13008,N_5675,N_6182);
xor U13009 (N_13009,N_8340,N_5591);
xor U13010 (N_13010,N_8386,N_9348);
xor U13011 (N_13011,N_6374,N_6018);
nand U13012 (N_13012,N_6805,N_9677);
nand U13013 (N_13013,N_8142,N_5328);
xnor U13014 (N_13014,N_7656,N_8227);
and U13015 (N_13015,N_8396,N_7850);
nor U13016 (N_13016,N_7513,N_8153);
or U13017 (N_13017,N_6676,N_6589);
xnor U13018 (N_13018,N_9619,N_9120);
or U13019 (N_13019,N_6820,N_6626);
xor U13020 (N_13020,N_6834,N_8074);
or U13021 (N_13021,N_9776,N_9481);
and U13022 (N_13022,N_7809,N_7850);
nor U13023 (N_13023,N_6439,N_5053);
and U13024 (N_13024,N_7593,N_8403);
nand U13025 (N_13025,N_9465,N_7615);
nor U13026 (N_13026,N_6866,N_5040);
nor U13027 (N_13027,N_7336,N_6717);
nor U13028 (N_13028,N_5205,N_9563);
xnor U13029 (N_13029,N_8227,N_7255);
nor U13030 (N_13030,N_8529,N_8567);
nor U13031 (N_13031,N_7501,N_7672);
nand U13032 (N_13032,N_7588,N_6958);
xnor U13033 (N_13033,N_6671,N_9318);
nor U13034 (N_13034,N_7006,N_7967);
nor U13035 (N_13035,N_5181,N_9197);
nor U13036 (N_13036,N_9113,N_7646);
nand U13037 (N_13037,N_7376,N_5939);
or U13038 (N_13038,N_6313,N_7619);
xor U13039 (N_13039,N_7268,N_9054);
xor U13040 (N_13040,N_8618,N_8804);
and U13041 (N_13041,N_9507,N_6329);
and U13042 (N_13042,N_5227,N_8390);
and U13043 (N_13043,N_6114,N_6796);
nor U13044 (N_13044,N_5785,N_8524);
or U13045 (N_13045,N_8617,N_5061);
xor U13046 (N_13046,N_7906,N_8099);
nor U13047 (N_13047,N_9448,N_7557);
xnor U13048 (N_13048,N_7426,N_5096);
nand U13049 (N_13049,N_6560,N_9831);
and U13050 (N_13050,N_5275,N_6572);
or U13051 (N_13051,N_9935,N_6524);
xor U13052 (N_13052,N_7214,N_6544);
or U13053 (N_13053,N_5749,N_7684);
and U13054 (N_13054,N_9280,N_8388);
nor U13055 (N_13055,N_9118,N_7385);
nand U13056 (N_13056,N_6614,N_7126);
or U13057 (N_13057,N_9279,N_8093);
or U13058 (N_13058,N_9593,N_9337);
nor U13059 (N_13059,N_7771,N_6412);
nor U13060 (N_13060,N_6795,N_7397);
xor U13061 (N_13061,N_7145,N_7210);
nor U13062 (N_13062,N_5551,N_7794);
or U13063 (N_13063,N_7127,N_6114);
xor U13064 (N_13064,N_5985,N_9078);
nor U13065 (N_13065,N_5326,N_9592);
or U13066 (N_13066,N_8051,N_7932);
and U13067 (N_13067,N_8927,N_8876);
xor U13068 (N_13068,N_9964,N_9106);
xnor U13069 (N_13069,N_7376,N_5506);
and U13070 (N_13070,N_8170,N_8088);
and U13071 (N_13071,N_7124,N_9214);
nor U13072 (N_13072,N_8719,N_9379);
xnor U13073 (N_13073,N_9574,N_8602);
xnor U13074 (N_13074,N_7263,N_6178);
xor U13075 (N_13075,N_5430,N_6479);
or U13076 (N_13076,N_9531,N_5599);
nor U13077 (N_13077,N_8671,N_8286);
and U13078 (N_13078,N_8869,N_5295);
nand U13079 (N_13079,N_7435,N_6262);
nand U13080 (N_13080,N_5535,N_5310);
and U13081 (N_13081,N_8068,N_8169);
or U13082 (N_13082,N_9394,N_8542);
or U13083 (N_13083,N_7682,N_6023);
nand U13084 (N_13084,N_9668,N_5052);
xnor U13085 (N_13085,N_5890,N_7703);
and U13086 (N_13086,N_6765,N_5780);
or U13087 (N_13087,N_6323,N_9273);
nand U13088 (N_13088,N_8256,N_6742);
xor U13089 (N_13089,N_9296,N_6413);
nand U13090 (N_13090,N_9335,N_6694);
and U13091 (N_13091,N_9961,N_6165);
xor U13092 (N_13092,N_9304,N_6112);
and U13093 (N_13093,N_7140,N_5910);
xor U13094 (N_13094,N_8308,N_9031);
nor U13095 (N_13095,N_7630,N_8557);
xnor U13096 (N_13096,N_5689,N_5704);
and U13097 (N_13097,N_8992,N_5760);
or U13098 (N_13098,N_9018,N_9259);
and U13099 (N_13099,N_9183,N_8802);
nor U13100 (N_13100,N_6894,N_8301);
nand U13101 (N_13101,N_9638,N_9162);
and U13102 (N_13102,N_9313,N_9564);
and U13103 (N_13103,N_5108,N_6021);
and U13104 (N_13104,N_7921,N_7149);
nand U13105 (N_13105,N_5677,N_5058);
nand U13106 (N_13106,N_7994,N_9488);
or U13107 (N_13107,N_7071,N_6782);
nor U13108 (N_13108,N_8121,N_6933);
or U13109 (N_13109,N_9252,N_8797);
and U13110 (N_13110,N_8473,N_8748);
or U13111 (N_13111,N_6528,N_7476);
xnor U13112 (N_13112,N_9413,N_8687);
xnor U13113 (N_13113,N_5414,N_7310);
nand U13114 (N_13114,N_7060,N_8751);
nand U13115 (N_13115,N_9372,N_9865);
and U13116 (N_13116,N_5087,N_5357);
nor U13117 (N_13117,N_5579,N_5691);
xnor U13118 (N_13118,N_6104,N_7134);
xor U13119 (N_13119,N_8209,N_9763);
and U13120 (N_13120,N_8884,N_9404);
or U13121 (N_13121,N_6814,N_6227);
and U13122 (N_13122,N_5575,N_9071);
or U13123 (N_13123,N_9085,N_9614);
and U13124 (N_13124,N_5750,N_9466);
xnor U13125 (N_13125,N_8168,N_7933);
nand U13126 (N_13126,N_9630,N_7550);
and U13127 (N_13127,N_6599,N_6907);
or U13128 (N_13128,N_7667,N_6571);
xnor U13129 (N_13129,N_5249,N_8491);
xnor U13130 (N_13130,N_8803,N_7730);
xor U13131 (N_13131,N_8472,N_9817);
nor U13132 (N_13132,N_6516,N_6416);
nand U13133 (N_13133,N_5687,N_9903);
xnor U13134 (N_13134,N_5153,N_6269);
nor U13135 (N_13135,N_9706,N_9426);
or U13136 (N_13136,N_9625,N_5360);
nand U13137 (N_13137,N_9160,N_8413);
and U13138 (N_13138,N_7479,N_8608);
and U13139 (N_13139,N_9230,N_5702);
nand U13140 (N_13140,N_6036,N_7389);
nor U13141 (N_13141,N_6005,N_6370);
nor U13142 (N_13142,N_8855,N_6748);
and U13143 (N_13143,N_5726,N_8342);
nand U13144 (N_13144,N_8697,N_6424);
xnor U13145 (N_13145,N_7149,N_5784);
nor U13146 (N_13146,N_5704,N_5220);
nor U13147 (N_13147,N_6863,N_5916);
nor U13148 (N_13148,N_7769,N_7969);
xor U13149 (N_13149,N_7255,N_9382);
and U13150 (N_13150,N_8276,N_5047);
nand U13151 (N_13151,N_8713,N_8619);
or U13152 (N_13152,N_8521,N_8663);
xor U13153 (N_13153,N_5116,N_6582);
or U13154 (N_13154,N_6038,N_7989);
xnor U13155 (N_13155,N_8973,N_6781);
and U13156 (N_13156,N_5692,N_5946);
and U13157 (N_13157,N_9982,N_8321);
nor U13158 (N_13158,N_9657,N_6926);
and U13159 (N_13159,N_6761,N_9573);
xnor U13160 (N_13160,N_9189,N_8639);
nor U13161 (N_13161,N_7205,N_7541);
nand U13162 (N_13162,N_8452,N_6532);
and U13163 (N_13163,N_9138,N_9477);
nor U13164 (N_13164,N_8208,N_9758);
or U13165 (N_13165,N_5195,N_8117);
and U13166 (N_13166,N_6495,N_5469);
or U13167 (N_13167,N_5863,N_7302);
or U13168 (N_13168,N_5515,N_6209);
nor U13169 (N_13169,N_8735,N_8845);
nor U13170 (N_13170,N_6231,N_9781);
xnor U13171 (N_13171,N_8834,N_7980);
and U13172 (N_13172,N_5496,N_8340);
and U13173 (N_13173,N_9979,N_8829);
or U13174 (N_13174,N_6751,N_8549);
nand U13175 (N_13175,N_9655,N_8625);
xor U13176 (N_13176,N_7309,N_7767);
or U13177 (N_13177,N_6459,N_9128);
or U13178 (N_13178,N_5613,N_9478);
or U13179 (N_13179,N_7124,N_9400);
and U13180 (N_13180,N_9186,N_5040);
nor U13181 (N_13181,N_8068,N_8686);
nand U13182 (N_13182,N_5510,N_7713);
nor U13183 (N_13183,N_7390,N_5278);
or U13184 (N_13184,N_9408,N_9188);
xor U13185 (N_13185,N_8756,N_5237);
nand U13186 (N_13186,N_5696,N_8669);
or U13187 (N_13187,N_9896,N_7873);
xor U13188 (N_13188,N_9055,N_6348);
or U13189 (N_13189,N_7655,N_7035);
xor U13190 (N_13190,N_6613,N_6991);
and U13191 (N_13191,N_8433,N_6163);
xnor U13192 (N_13192,N_8582,N_5087);
or U13193 (N_13193,N_7445,N_6538);
xnor U13194 (N_13194,N_8895,N_9393);
or U13195 (N_13195,N_9763,N_7849);
or U13196 (N_13196,N_9355,N_7673);
or U13197 (N_13197,N_7450,N_6113);
nor U13198 (N_13198,N_8081,N_7734);
nor U13199 (N_13199,N_6330,N_7907);
or U13200 (N_13200,N_9823,N_5945);
xor U13201 (N_13201,N_8400,N_9394);
and U13202 (N_13202,N_7409,N_5315);
xor U13203 (N_13203,N_5646,N_7348);
or U13204 (N_13204,N_8161,N_7398);
or U13205 (N_13205,N_8675,N_9262);
nor U13206 (N_13206,N_8979,N_5664);
nand U13207 (N_13207,N_5688,N_5004);
or U13208 (N_13208,N_9762,N_8719);
xnor U13209 (N_13209,N_6409,N_9797);
nand U13210 (N_13210,N_5614,N_7420);
nor U13211 (N_13211,N_6533,N_6994);
xor U13212 (N_13212,N_9783,N_9790);
xnor U13213 (N_13213,N_5541,N_6362);
nand U13214 (N_13214,N_6067,N_5914);
xor U13215 (N_13215,N_7277,N_8471);
xnor U13216 (N_13216,N_7677,N_8933);
or U13217 (N_13217,N_8722,N_9212);
nor U13218 (N_13218,N_7472,N_7970);
nand U13219 (N_13219,N_7703,N_8181);
nand U13220 (N_13220,N_5193,N_5450);
and U13221 (N_13221,N_6684,N_5566);
nand U13222 (N_13222,N_5075,N_8752);
nor U13223 (N_13223,N_8923,N_9267);
and U13224 (N_13224,N_7544,N_9256);
and U13225 (N_13225,N_7868,N_6341);
nor U13226 (N_13226,N_9756,N_6702);
nor U13227 (N_13227,N_6342,N_5044);
xor U13228 (N_13228,N_5574,N_7583);
nand U13229 (N_13229,N_5890,N_5437);
and U13230 (N_13230,N_7040,N_7524);
nor U13231 (N_13231,N_9086,N_6108);
and U13232 (N_13232,N_5841,N_5886);
nor U13233 (N_13233,N_7336,N_5115);
or U13234 (N_13234,N_5165,N_6836);
and U13235 (N_13235,N_7068,N_9505);
or U13236 (N_13236,N_9282,N_7943);
nor U13237 (N_13237,N_9015,N_8494);
or U13238 (N_13238,N_6819,N_9790);
or U13239 (N_13239,N_9223,N_8803);
nand U13240 (N_13240,N_9645,N_8882);
nor U13241 (N_13241,N_6647,N_6731);
nor U13242 (N_13242,N_9212,N_5187);
nor U13243 (N_13243,N_8573,N_9483);
and U13244 (N_13244,N_7633,N_7670);
nand U13245 (N_13245,N_5387,N_9292);
xnor U13246 (N_13246,N_9913,N_8920);
or U13247 (N_13247,N_6871,N_8985);
or U13248 (N_13248,N_6666,N_5789);
nand U13249 (N_13249,N_6338,N_7812);
and U13250 (N_13250,N_8362,N_9245);
nor U13251 (N_13251,N_7672,N_6646);
or U13252 (N_13252,N_9823,N_6173);
xor U13253 (N_13253,N_8544,N_9027);
nand U13254 (N_13254,N_9462,N_9271);
nor U13255 (N_13255,N_6052,N_9395);
nor U13256 (N_13256,N_5698,N_8010);
nand U13257 (N_13257,N_8916,N_7000);
or U13258 (N_13258,N_6743,N_8212);
xor U13259 (N_13259,N_5679,N_7650);
xor U13260 (N_13260,N_6443,N_8652);
nand U13261 (N_13261,N_5898,N_6241);
nand U13262 (N_13262,N_5675,N_7383);
or U13263 (N_13263,N_6582,N_8330);
xnor U13264 (N_13264,N_9874,N_5046);
nand U13265 (N_13265,N_5452,N_8452);
or U13266 (N_13266,N_6829,N_8009);
or U13267 (N_13267,N_5411,N_9155);
or U13268 (N_13268,N_7930,N_8510);
and U13269 (N_13269,N_8338,N_6932);
or U13270 (N_13270,N_8721,N_9625);
and U13271 (N_13271,N_6801,N_8771);
nand U13272 (N_13272,N_8669,N_9930);
xor U13273 (N_13273,N_6331,N_9591);
xor U13274 (N_13274,N_7074,N_8280);
nand U13275 (N_13275,N_8415,N_7769);
nand U13276 (N_13276,N_6608,N_5364);
and U13277 (N_13277,N_8861,N_8213);
or U13278 (N_13278,N_7277,N_5858);
xor U13279 (N_13279,N_8494,N_7346);
and U13280 (N_13280,N_9585,N_6183);
or U13281 (N_13281,N_7435,N_7813);
nor U13282 (N_13282,N_9254,N_9534);
and U13283 (N_13283,N_5782,N_7055);
and U13284 (N_13284,N_7145,N_8917);
xnor U13285 (N_13285,N_6941,N_6158);
and U13286 (N_13286,N_9636,N_5375);
nor U13287 (N_13287,N_8799,N_8852);
xor U13288 (N_13288,N_5156,N_8552);
nand U13289 (N_13289,N_9122,N_5449);
and U13290 (N_13290,N_7292,N_6658);
or U13291 (N_13291,N_8256,N_9303);
or U13292 (N_13292,N_9209,N_7473);
nor U13293 (N_13293,N_9214,N_6610);
nor U13294 (N_13294,N_5588,N_8500);
or U13295 (N_13295,N_9192,N_9553);
or U13296 (N_13296,N_9643,N_8125);
or U13297 (N_13297,N_9849,N_9986);
nand U13298 (N_13298,N_8145,N_9219);
xor U13299 (N_13299,N_8789,N_7303);
nor U13300 (N_13300,N_6758,N_7132);
or U13301 (N_13301,N_7766,N_9333);
nor U13302 (N_13302,N_6681,N_5186);
and U13303 (N_13303,N_6011,N_9845);
nand U13304 (N_13304,N_8940,N_8543);
or U13305 (N_13305,N_5806,N_6618);
or U13306 (N_13306,N_6017,N_7216);
nor U13307 (N_13307,N_8351,N_9731);
or U13308 (N_13308,N_6528,N_8356);
nand U13309 (N_13309,N_8756,N_7385);
nand U13310 (N_13310,N_5134,N_9916);
or U13311 (N_13311,N_8645,N_6837);
xnor U13312 (N_13312,N_9475,N_9376);
or U13313 (N_13313,N_6533,N_8704);
nor U13314 (N_13314,N_8430,N_9866);
or U13315 (N_13315,N_8057,N_9379);
nor U13316 (N_13316,N_5710,N_7948);
nand U13317 (N_13317,N_5914,N_6346);
nor U13318 (N_13318,N_9770,N_6876);
or U13319 (N_13319,N_7463,N_9071);
xor U13320 (N_13320,N_8415,N_8525);
nand U13321 (N_13321,N_7626,N_6026);
xnor U13322 (N_13322,N_8364,N_6527);
xnor U13323 (N_13323,N_8779,N_5602);
nand U13324 (N_13324,N_9812,N_7812);
nor U13325 (N_13325,N_5152,N_5097);
or U13326 (N_13326,N_9130,N_9508);
or U13327 (N_13327,N_5496,N_7010);
and U13328 (N_13328,N_5157,N_7493);
xor U13329 (N_13329,N_5106,N_9597);
and U13330 (N_13330,N_9164,N_6933);
xor U13331 (N_13331,N_8179,N_7618);
or U13332 (N_13332,N_8634,N_8722);
nor U13333 (N_13333,N_5576,N_5641);
and U13334 (N_13334,N_5018,N_8874);
nand U13335 (N_13335,N_5244,N_8850);
and U13336 (N_13336,N_9233,N_5497);
xor U13337 (N_13337,N_8799,N_7738);
and U13338 (N_13338,N_8559,N_7047);
xnor U13339 (N_13339,N_6127,N_7379);
and U13340 (N_13340,N_5131,N_7070);
nor U13341 (N_13341,N_8814,N_7690);
xor U13342 (N_13342,N_8675,N_8749);
nand U13343 (N_13343,N_5642,N_5645);
and U13344 (N_13344,N_6834,N_6969);
xnor U13345 (N_13345,N_5868,N_5990);
and U13346 (N_13346,N_5842,N_7681);
and U13347 (N_13347,N_6059,N_9204);
or U13348 (N_13348,N_6974,N_7770);
xor U13349 (N_13349,N_5925,N_6838);
xor U13350 (N_13350,N_7100,N_5568);
nor U13351 (N_13351,N_8375,N_5934);
xor U13352 (N_13352,N_6013,N_9927);
nand U13353 (N_13353,N_7382,N_9179);
and U13354 (N_13354,N_6513,N_9153);
or U13355 (N_13355,N_7608,N_7471);
xnor U13356 (N_13356,N_8418,N_6347);
nand U13357 (N_13357,N_7632,N_9253);
and U13358 (N_13358,N_6604,N_6894);
and U13359 (N_13359,N_8020,N_7302);
nand U13360 (N_13360,N_6690,N_5955);
and U13361 (N_13361,N_9139,N_7316);
nand U13362 (N_13362,N_6248,N_7998);
and U13363 (N_13363,N_9497,N_8814);
xnor U13364 (N_13364,N_8949,N_7475);
or U13365 (N_13365,N_8409,N_5789);
xnor U13366 (N_13366,N_5094,N_5547);
xor U13367 (N_13367,N_8138,N_6279);
xor U13368 (N_13368,N_8476,N_7217);
xor U13369 (N_13369,N_5285,N_5021);
and U13370 (N_13370,N_7217,N_8625);
or U13371 (N_13371,N_6222,N_7878);
xor U13372 (N_13372,N_6148,N_6430);
or U13373 (N_13373,N_8100,N_5166);
nand U13374 (N_13374,N_9136,N_7851);
nand U13375 (N_13375,N_8908,N_9344);
xnor U13376 (N_13376,N_8618,N_9837);
nand U13377 (N_13377,N_7665,N_7529);
nor U13378 (N_13378,N_7354,N_5482);
nand U13379 (N_13379,N_5272,N_9399);
xor U13380 (N_13380,N_6129,N_5154);
and U13381 (N_13381,N_7581,N_7338);
xnor U13382 (N_13382,N_7292,N_7946);
and U13383 (N_13383,N_8275,N_5536);
nand U13384 (N_13384,N_8778,N_5999);
nand U13385 (N_13385,N_8971,N_7830);
xor U13386 (N_13386,N_6010,N_6502);
or U13387 (N_13387,N_5573,N_6348);
nand U13388 (N_13388,N_6832,N_9991);
and U13389 (N_13389,N_8776,N_9120);
xor U13390 (N_13390,N_7322,N_5533);
or U13391 (N_13391,N_7610,N_5382);
nor U13392 (N_13392,N_6200,N_9888);
nor U13393 (N_13393,N_5571,N_9909);
nor U13394 (N_13394,N_9907,N_9441);
nand U13395 (N_13395,N_5714,N_6962);
and U13396 (N_13396,N_8140,N_9720);
or U13397 (N_13397,N_6679,N_7392);
xnor U13398 (N_13398,N_8126,N_8613);
and U13399 (N_13399,N_9004,N_6059);
nor U13400 (N_13400,N_6136,N_6672);
or U13401 (N_13401,N_7092,N_5222);
nand U13402 (N_13402,N_7425,N_5954);
xnor U13403 (N_13403,N_5026,N_7080);
nand U13404 (N_13404,N_7255,N_8848);
or U13405 (N_13405,N_5257,N_6686);
nor U13406 (N_13406,N_7099,N_5744);
nand U13407 (N_13407,N_7241,N_7719);
and U13408 (N_13408,N_7264,N_8903);
or U13409 (N_13409,N_9532,N_7463);
nor U13410 (N_13410,N_5654,N_7793);
xor U13411 (N_13411,N_8838,N_6074);
and U13412 (N_13412,N_7071,N_6054);
or U13413 (N_13413,N_8915,N_8963);
xor U13414 (N_13414,N_9189,N_7785);
nor U13415 (N_13415,N_8515,N_8155);
xor U13416 (N_13416,N_8218,N_6844);
or U13417 (N_13417,N_7062,N_8267);
xor U13418 (N_13418,N_5166,N_8076);
nor U13419 (N_13419,N_5060,N_5102);
and U13420 (N_13420,N_9977,N_7270);
and U13421 (N_13421,N_9766,N_9059);
nand U13422 (N_13422,N_5392,N_8047);
and U13423 (N_13423,N_6177,N_8146);
xnor U13424 (N_13424,N_6846,N_5200);
and U13425 (N_13425,N_7427,N_9973);
nor U13426 (N_13426,N_5445,N_5920);
and U13427 (N_13427,N_5949,N_7651);
xnor U13428 (N_13428,N_8185,N_6230);
xor U13429 (N_13429,N_9497,N_7027);
xnor U13430 (N_13430,N_5967,N_9853);
nor U13431 (N_13431,N_6001,N_5681);
xor U13432 (N_13432,N_9579,N_6278);
and U13433 (N_13433,N_5177,N_8716);
nand U13434 (N_13434,N_9120,N_5689);
nor U13435 (N_13435,N_8669,N_8140);
and U13436 (N_13436,N_6458,N_9261);
or U13437 (N_13437,N_8764,N_9670);
nand U13438 (N_13438,N_8892,N_8570);
nand U13439 (N_13439,N_5964,N_5663);
or U13440 (N_13440,N_8945,N_7320);
xor U13441 (N_13441,N_8015,N_7353);
and U13442 (N_13442,N_6000,N_7791);
and U13443 (N_13443,N_8627,N_6516);
xnor U13444 (N_13444,N_6762,N_7650);
nor U13445 (N_13445,N_5186,N_6092);
or U13446 (N_13446,N_5639,N_6638);
nand U13447 (N_13447,N_5230,N_7237);
nor U13448 (N_13448,N_8787,N_9516);
nor U13449 (N_13449,N_5866,N_7607);
nor U13450 (N_13450,N_9680,N_8443);
nor U13451 (N_13451,N_9506,N_9845);
nand U13452 (N_13452,N_9253,N_7466);
nand U13453 (N_13453,N_6357,N_6405);
nor U13454 (N_13454,N_7330,N_7873);
or U13455 (N_13455,N_5879,N_6837);
and U13456 (N_13456,N_7903,N_6201);
nand U13457 (N_13457,N_7749,N_8658);
nor U13458 (N_13458,N_6925,N_9741);
and U13459 (N_13459,N_6820,N_7306);
or U13460 (N_13460,N_5891,N_9321);
nor U13461 (N_13461,N_5613,N_6095);
nor U13462 (N_13462,N_6306,N_9227);
xnor U13463 (N_13463,N_9926,N_5905);
nor U13464 (N_13464,N_8688,N_5505);
and U13465 (N_13465,N_5863,N_8995);
nand U13466 (N_13466,N_8411,N_8229);
and U13467 (N_13467,N_6621,N_7544);
and U13468 (N_13468,N_8943,N_9662);
xor U13469 (N_13469,N_8223,N_8624);
and U13470 (N_13470,N_9045,N_6091);
nand U13471 (N_13471,N_7777,N_7797);
nand U13472 (N_13472,N_5980,N_7443);
xnor U13473 (N_13473,N_8598,N_5302);
and U13474 (N_13474,N_8424,N_8877);
and U13475 (N_13475,N_7353,N_8951);
or U13476 (N_13476,N_6513,N_7518);
xor U13477 (N_13477,N_9712,N_9615);
and U13478 (N_13478,N_8936,N_8356);
and U13479 (N_13479,N_7123,N_8701);
and U13480 (N_13480,N_6355,N_8102);
nor U13481 (N_13481,N_6396,N_7277);
nand U13482 (N_13482,N_7039,N_5487);
nor U13483 (N_13483,N_5064,N_8203);
and U13484 (N_13484,N_9020,N_7117);
xor U13485 (N_13485,N_5992,N_8080);
or U13486 (N_13486,N_9824,N_5481);
xnor U13487 (N_13487,N_7852,N_8852);
xor U13488 (N_13488,N_6020,N_8096);
nor U13489 (N_13489,N_8892,N_5448);
nand U13490 (N_13490,N_7370,N_8761);
and U13491 (N_13491,N_9854,N_5279);
nor U13492 (N_13492,N_8122,N_9824);
nand U13493 (N_13493,N_7550,N_6580);
and U13494 (N_13494,N_9216,N_9411);
nand U13495 (N_13495,N_5931,N_6603);
and U13496 (N_13496,N_8778,N_5782);
or U13497 (N_13497,N_7492,N_9301);
or U13498 (N_13498,N_9416,N_7488);
nor U13499 (N_13499,N_5472,N_9290);
or U13500 (N_13500,N_8678,N_9039);
nor U13501 (N_13501,N_8528,N_7124);
nor U13502 (N_13502,N_7077,N_8006);
or U13503 (N_13503,N_5814,N_8960);
xor U13504 (N_13504,N_8908,N_8521);
nand U13505 (N_13505,N_8874,N_8902);
xor U13506 (N_13506,N_5560,N_7470);
xor U13507 (N_13507,N_6740,N_8956);
or U13508 (N_13508,N_5698,N_6976);
or U13509 (N_13509,N_7304,N_6601);
and U13510 (N_13510,N_5184,N_7322);
xor U13511 (N_13511,N_8775,N_9967);
nor U13512 (N_13512,N_9117,N_6803);
xnor U13513 (N_13513,N_7451,N_7174);
nand U13514 (N_13514,N_6878,N_7978);
and U13515 (N_13515,N_9068,N_9404);
and U13516 (N_13516,N_6236,N_6823);
nand U13517 (N_13517,N_5775,N_7423);
xor U13518 (N_13518,N_9169,N_9574);
nor U13519 (N_13519,N_7400,N_7900);
xnor U13520 (N_13520,N_7058,N_5130);
and U13521 (N_13521,N_6908,N_5278);
and U13522 (N_13522,N_6251,N_7546);
and U13523 (N_13523,N_5662,N_6873);
and U13524 (N_13524,N_5444,N_5760);
nand U13525 (N_13525,N_6034,N_8898);
nor U13526 (N_13526,N_8777,N_6792);
nand U13527 (N_13527,N_6022,N_7626);
and U13528 (N_13528,N_6492,N_7710);
and U13529 (N_13529,N_9270,N_8955);
or U13530 (N_13530,N_7272,N_9565);
nand U13531 (N_13531,N_5884,N_8209);
nor U13532 (N_13532,N_6031,N_6042);
and U13533 (N_13533,N_7378,N_5938);
or U13534 (N_13534,N_6173,N_7812);
nor U13535 (N_13535,N_9355,N_7819);
and U13536 (N_13536,N_6093,N_9851);
and U13537 (N_13537,N_5823,N_8403);
nor U13538 (N_13538,N_9381,N_7422);
nor U13539 (N_13539,N_8500,N_6698);
or U13540 (N_13540,N_6291,N_6056);
xnor U13541 (N_13541,N_7960,N_9453);
xor U13542 (N_13542,N_9050,N_5637);
or U13543 (N_13543,N_9034,N_9411);
and U13544 (N_13544,N_9170,N_9902);
nand U13545 (N_13545,N_6614,N_9490);
nand U13546 (N_13546,N_9694,N_5251);
or U13547 (N_13547,N_9788,N_6836);
xnor U13548 (N_13548,N_5343,N_8607);
and U13549 (N_13549,N_7055,N_6829);
nor U13550 (N_13550,N_8107,N_6331);
or U13551 (N_13551,N_9033,N_6994);
and U13552 (N_13552,N_9506,N_9404);
and U13553 (N_13553,N_9048,N_7601);
and U13554 (N_13554,N_5992,N_7767);
and U13555 (N_13555,N_5073,N_8618);
and U13556 (N_13556,N_6249,N_5197);
or U13557 (N_13557,N_6846,N_7846);
and U13558 (N_13558,N_9786,N_6378);
xnor U13559 (N_13559,N_6402,N_8530);
nor U13560 (N_13560,N_8473,N_8784);
and U13561 (N_13561,N_8155,N_8694);
xor U13562 (N_13562,N_5994,N_5453);
or U13563 (N_13563,N_8267,N_6895);
or U13564 (N_13564,N_6014,N_6653);
xor U13565 (N_13565,N_5078,N_9887);
xnor U13566 (N_13566,N_5372,N_9631);
nand U13567 (N_13567,N_7420,N_9347);
and U13568 (N_13568,N_8415,N_9349);
or U13569 (N_13569,N_7432,N_9540);
or U13570 (N_13570,N_6925,N_8572);
xnor U13571 (N_13571,N_7303,N_5778);
nor U13572 (N_13572,N_7968,N_5539);
xor U13573 (N_13573,N_8586,N_9910);
or U13574 (N_13574,N_9047,N_5479);
nand U13575 (N_13575,N_5443,N_8945);
nor U13576 (N_13576,N_7853,N_9557);
and U13577 (N_13577,N_5908,N_7271);
xor U13578 (N_13578,N_6556,N_7607);
nor U13579 (N_13579,N_6284,N_7361);
xor U13580 (N_13580,N_6318,N_5663);
nand U13581 (N_13581,N_5806,N_5332);
nand U13582 (N_13582,N_8916,N_6821);
and U13583 (N_13583,N_6442,N_5296);
nand U13584 (N_13584,N_5815,N_8836);
nor U13585 (N_13585,N_9888,N_9158);
nand U13586 (N_13586,N_5935,N_9647);
nor U13587 (N_13587,N_8551,N_9822);
xnor U13588 (N_13588,N_7234,N_9097);
or U13589 (N_13589,N_9915,N_9112);
or U13590 (N_13590,N_7124,N_9361);
nand U13591 (N_13591,N_5345,N_9249);
nor U13592 (N_13592,N_8315,N_7569);
nor U13593 (N_13593,N_7250,N_6544);
xor U13594 (N_13594,N_5351,N_5609);
xor U13595 (N_13595,N_8773,N_7672);
nor U13596 (N_13596,N_6237,N_5536);
or U13597 (N_13597,N_8413,N_8391);
or U13598 (N_13598,N_5208,N_7931);
xor U13599 (N_13599,N_6684,N_9545);
and U13600 (N_13600,N_7352,N_6038);
or U13601 (N_13601,N_5886,N_6916);
xnor U13602 (N_13602,N_8936,N_5114);
and U13603 (N_13603,N_6618,N_7969);
and U13604 (N_13604,N_6104,N_9782);
nand U13605 (N_13605,N_8363,N_6632);
or U13606 (N_13606,N_8282,N_6109);
xor U13607 (N_13607,N_5661,N_6379);
and U13608 (N_13608,N_7581,N_6404);
nor U13609 (N_13609,N_8725,N_5245);
or U13610 (N_13610,N_5746,N_8750);
xnor U13611 (N_13611,N_6136,N_6558);
nor U13612 (N_13612,N_7091,N_6554);
and U13613 (N_13613,N_8246,N_9782);
nor U13614 (N_13614,N_9327,N_9103);
or U13615 (N_13615,N_8773,N_5099);
and U13616 (N_13616,N_8082,N_9172);
xor U13617 (N_13617,N_7793,N_8200);
or U13618 (N_13618,N_8414,N_8245);
nand U13619 (N_13619,N_9216,N_5770);
nor U13620 (N_13620,N_9641,N_7454);
or U13621 (N_13621,N_6282,N_9145);
nand U13622 (N_13622,N_7463,N_7379);
nor U13623 (N_13623,N_9517,N_7026);
nor U13624 (N_13624,N_7798,N_9950);
nand U13625 (N_13625,N_8820,N_8685);
xnor U13626 (N_13626,N_5213,N_8834);
xnor U13627 (N_13627,N_5482,N_5171);
nand U13628 (N_13628,N_9899,N_9117);
nor U13629 (N_13629,N_7914,N_9132);
nand U13630 (N_13630,N_9946,N_7125);
nor U13631 (N_13631,N_5198,N_7939);
or U13632 (N_13632,N_7601,N_5690);
nor U13633 (N_13633,N_7816,N_9714);
xnor U13634 (N_13634,N_5582,N_5016);
and U13635 (N_13635,N_8826,N_7293);
and U13636 (N_13636,N_8899,N_7757);
nor U13637 (N_13637,N_6409,N_7605);
nand U13638 (N_13638,N_5787,N_7417);
xnor U13639 (N_13639,N_6565,N_6391);
nand U13640 (N_13640,N_7860,N_9681);
or U13641 (N_13641,N_5769,N_6705);
nand U13642 (N_13642,N_6749,N_8543);
or U13643 (N_13643,N_6552,N_8135);
nor U13644 (N_13644,N_7655,N_6485);
nand U13645 (N_13645,N_9226,N_6282);
nand U13646 (N_13646,N_7498,N_8667);
xor U13647 (N_13647,N_7241,N_9020);
nor U13648 (N_13648,N_9557,N_5393);
nand U13649 (N_13649,N_7846,N_5251);
xnor U13650 (N_13650,N_8981,N_8205);
xnor U13651 (N_13651,N_6719,N_9200);
nor U13652 (N_13652,N_9451,N_6688);
xnor U13653 (N_13653,N_8446,N_7024);
and U13654 (N_13654,N_6965,N_6655);
nor U13655 (N_13655,N_8035,N_6337);
nand U13656 (N_13656,N_7383,N_9047);
nor U13657 (N_13657,N_5272,N_8872);
nor U13658 (N_13658,N_7536,N_7210);
xnor U13659 (N_13659,N_8432,N_7251);
nor U13660 (N_13660,N_5865,N_5499);
nand U13661 (N_13661,N_7005,N_7647);
xnor U13662 (N_13662,N_6386,N_7687);
and U13663 (N_13663,N_6885,N_6411);
nor U13664 (N_13664,N_6400,N_6378);
nor U13665 (N_13665,N_7828,N_6709);
and U13666 (N_13666,N_9582,N_9398);
nor U13667 (N_13667,N_7809,N_5933);
nand U13668 (N_13668,N_7842,N_5107);
nand U13669 (N_13669,N_9915,N_8589);
nor U13670 (N_13670,N_9339,N_5499);
and U13671 (N_13671,N_8639,N_6844);
nor U13672 (N_13672,N_6180,N_6280);
nor U13673 (N_13673,N_5441,N_7578);
xnor U13674 (N_13674,N_7109,N_5933);
nor U13675 (N_13675,N_5574,N_5626);
nor U13676 (N_13676,N_8479,N_6719);
xnor U13677 (N_13677,N_8456,N_9836);
nor U13678 (N_13678,N_5635,N_6241);
nand U13679 (N_13679,N_5602,N_9989);
and U13680 (N_13680,N_8358,N_7035);
nor U13681 (N_13681,N_6909,N_8318);
nand U13682 (N_13682,N_7320,N_8050);
or U13683 (N_13683,N_5630,N_5516);
xor U13684 (N_13684,N_7753,N_9754);
nor U13685 (N_13685,N_5537,N_7043);
and U13686 (N_13686,N_9594,N_7844);
or U13687 (N_13687,N_6682,N_7984);
or U13688 (N_13688,N_8813,N_9365);
or U13689 (N_13689,N_5159,N_9770);
xor U13690 (N_13690,N_7669,N_7198);
nor U13691 (N_13691,N_9992,N_6553);
or U13692 (N_13692,N_5829,N_7383);
or U13693 (N_13693,N_9790,N_9660);
nor U13694 (N_13694,N_5181,N_8337);
xor U13695 (N_13695,N_5374,N_8148);
nor U13696 (N_13696,N_5205,N_5284);
and U13697 (N_13697,N_8092,N_6151);
or U13698 (N_13698,N_8085,N_6073);
xnor U13699 (N_13699,N_5907,N_5692);
or U13700 (N_13700,N_7603,N_8209);
xnor U13701 (N_13701,N_9157,N_5048);
xnor U13702 (N_13702,N_8486,N_7437);
and U13703 (N_13703,N_6642,N_9957);
nor U13704 (N_13704,N_5979,N_9353);
xor U13705 (N_13705,N_8463,N_6064);
and U13706 (N_13706,N_5145,N_7714);
or U13707 (N_13707,N_7092,N_6285);
or U13708 (N_13708,N_9432,N_7690);
nand U13709 (N_13709,N_9278,N_7509);
xor U13710 (N_13710,N_8064,N_7657);
nor U13711 (N_13711,N_8494,N_9633);
or U13712 (N_13712,N_7385,N_9808);
nand U13713 (N_13713,N_8627,N_5707);
and U13714 (N_13714,N_8299,N_6765);
or U13715 (N_13715,N_7101,N_7106);
xnor U13716 (N_13716,N_6622,N_5554);
xor U13717 (N_13717,N_8405,N_7315);
nand U13718 (N_13718,N_8388,N_8335);
nand U13719 (N_13719,N_7999,N_8712);
nor U13720 (N_13720,N_8188,N_5466);
nand U13721 (N_13721,N_7949,N_6883);
nand U13722 (N_13722,N_8353,N_7023);
nor U13723 (N_13723,N_5522,N_9414);
and U13724 (N_13724,N_5993,N_7890);
or U13725 (N_13725,N_9023,N_5735);
nor U13726 (N_13726,N_7222,N_5113);
xor U13727 (N_13727,N_6374,N_7599);
or U13728 (N_13728,N_5247,N_7043);
nor U13729 (N_13729,N_9510,N_5531);
and U13730 (N_13730,N_6915,N_7899);
nand U13731 (N_13731,N_9183,N_7211);
nand U13732 (N_13732,N_8558,N_6484);
or U13733 (N_13733,N_9014,N_9883);
nor U13734 (N_13734,N_8336,N_6889);
nor U13735 (N_13735,N_7402,N_8221);
xnor U13736 (N_13736,N_7866,N_7717);
or U13737 (N_13737,N_5967,N_9619);
or U13738 (N_13738,N_6746,N_6621);
xor U13739 (N_13739,N_5287,N_6683);
nand U13740 (N_13740,N_5943,N_7772);
and U13741 (N_13741,N_6602,N_9016);
or U13742 (N_13742,N_9887,N_5315);
and U13743 (N_13743,N_5900,N_7605);
and U13744 (N_13744,N_6247,N_7922);
nor U13745 (N_13745,N_8972,N_9310);
nand U13746 (N_13746,N_9082,N_5309);
xor U13747 (N_13747,N_8519,N_8336);
and U13748 (N_13748,N_8103,N_8744);
or U13749 (N_13749,N_7476,N_9686);
xnor U13750 (N_13750,N_9341,N_8791);
nand U13751 (N_13751,N_8118,N_8177);
and U13752 (N_13752,N_7960,N_5910);
and U13753 (N_13753,N_6214,N_7333);
xor U13754 (N_13754,N_8607,N_5202);
nor U13755 (N_13755,N_9544,N_9780);
and U13756 (N_13756,N_6936,N_8580);
or U13757 (N_13757,N_6571,N_9601);
and U13758 (N_13758,N_7186,N_5137);
and U13759 (N_13759,N_7053,N_5874);
nor U13760 (N_13760,N_6427,N_7060);
nor U13761 (N_13761,N_8501,N_7630);
and U13762 (N_13762,N_5236,N_6188);
nand U13763 (N_13763,N_6944,N_7669);
and U13764 (N_13764,N_8996,N_6405);
and U13765 (N_13765,N_8803,N_6251);
nor U13766 (N_13766,N_5805,N_7321);
xnor U13767 (N_13767,N_5693,N_5975);
or U13768 (N_13768,N_7063,N_7458);
nand U13769 (N_13769,N_7896,N_6781);
xnor U13770 (N_13770,N_8639,N_7305);
nor U13771 (N_13771,N_6018,N_8504);
nand U13772 (N_13772,N_6462,N_9795);
or U13773 (N_13773,N_7789,N_6841);
xnor U13774 (N_13774,N_8165,N_7467);
nand U13775 (N_13775,N_5908,N_5096);
nand U13776 (N_13776,N_5024,N_8991);
nor U13777 (N_13777,N_8978,N_5160);
nand U13778 (N_13778,N_5818,N_7311);
or U13779 (N_13779,N_7514,N_8665);
xnor U13780 (N_13780,N_8695,N_8766);
nand U13781 (N_13781,N_7881,N_9116);
xnor U13782 (N_13782,N_9391,N_8929);
nor U13783 (N_13783,N_6013,N_7372);
nand U13784 (N_13784,N_8181,N_5107);
nor U13785 (N_13785,N_7341,N_5176);
nand U13786 (N_13786,N_7217,N_8484);
or U13787 (N_13787,N_6030,N_9980);
or U13788 (N_13788,N_7120,N_6634);
nand U13789 (N_13789,N_8976,N_6425);
nor U13790 (N_13790,N_9608,N_8769);
or U13791 (N_13791,N_9417,N_6476);
nand U13792 (N_13792,N_6964,N_8823);
and U13793 (N_13793,N_5840,N_7265);
xor U13794 (N_13794,N_8311,N_8746);
xor U13795 (N_13795,N_6190,N_6806);
nand U13796 (N_13796,N_8146,N_7750);
and U13797 (N_13797,N_6168,N_7703);
xor U13798 (N_13798,N_8235,N_7594);
and U13799 (N_13799,N_7784,N_8090);
nand U13800 (N_13800,N_5519,N_8661);
xor U13801 (N_13801,N_9251,N_6984);
and U13802 (N_13802,N_5835,N_5745);
and U13803 (N_13803,N_5800,N_7067);
or U13804 (N_13804,N_7487,N_7141);
xor U13805 (N_13805,N_5404,N_8851);
and U13806 (N_13806,N_8957,N_7282);
nor U13807 (N_13807,N_8446,N_5928);
xnor U13808 (N_13808,N_7257,N_7653);
nand U13809 (N_13809,N_8723,N_6799);
and U13810 (N_13810,N_9982,N_5915);
nand U13811 (N_13811,N_5147,N_9226);
nand U13812 (N_13812,N_9377,N_5421);
nand U13813 (N_13813,N_7854,N_5833);
nand U13814 (N_13814,N_8347,N_9215);
xnor U13815 (N_13815,N_7257,N_5568);
or U13816 (N_13816,N_6876,N_9513);
or U13817 (N_13817,N_6565,N_5105);
xnor U13818 (N_13818,N_8089,N_8061);
nor U13819 (N_13819,N_6990,N_7435);
nor U13820 (N_13820,N_8593,N_5693);
and U13821 (N_13821,N_5307,N_7405);
nor U13822 (N_13822,N_8610,N_6017);
nand U13823 (N_13823,N_8657,N_7969);
and U13824 (N_13824,N_8350,N_9533);
or U13825 (N_13825,N_9716,N_7408);
or U13826 (N_13826,N_6245,N_5774);
xor U13827 (N_13827,N_9318,N_8833);
xnor U13828 (N_13828,N_6302,N_6106);
nor U13829 (N_13829,N_7887,N_8175);
xor U13830 (N_13830,N_9034,N_7252);
or U13831 (N_13831,N_7148,N_7330);
nor U13832 (N_13832,N_9580,N_6993);
xnor U13833 (N_13833,N_5032,N_9678);
or U13834 (N_13834,N_7790,N_5308);
xor U13835 (N_13835,N_9449,N_9985);
nand U13836 (N_13836,N_9043,N_5107);
and U13837 (N_13837,N_5118,N_8123);
or U13838 (N_13838,N_9326,N_6543);
xnor U13839 (N_13839,N_5410,N_7806);
or U13840 (N_13840,N_9773,N_9902);
xor U13841 (N_13841,N_9481,N_6717);
xor U13842 (N_13842,N_7615,N_7909);
or U13843 (N_13843,N_5246,N_5875);
and U13844 (N_13844,N_8901,N_5732);
xor U13845 (N_13845,N_5233,N_7658);
nor U13846 (N_13846,N_7064,N_8464);
xnor U13847 (N_13847,N_9236,N_6858);
nand U13848 (N_13848,N_9665,N_9240);
nand U13849 (N_13849,N_9655,N_7701);
nand U13850 (N_13850,N_9353,N_9892);
nor U13851 (N_13851,N_9964,N_8495);
nand U13852 (N_13852,N_5985,N_5986);
xnor U13853 (N_13853,N_7134,N_9475);
or U13854 (N_13854,N_5990,N_8102);
nor U13855 (N_13855,N_5754,N_5425);
xnor U13856 (N_13856,N_9390,N_7399);
nand U13857 (N_13857,N_5159,N_8653);
nor U13858 (N_13858,N_6379,N_7155);
and U13859 (N_13859,N_6964,N_6290);
or U13860 (N_13860,N_9275,N_7600);
or U13861 (N_13861,N_5553,N_6706);
and U13862 (N_13862,N_7197,N_5939);
or U13863 (N_13863,N_8364,N_5318);
nand U13864 (N_13864,N_8996,N_7597);
nand U13865 (N_13865,N_9166,N_6302);
and U13866 (N_13866,N_6667,N_5554);
or U13867 (N_13867,N_5279,N_7112);
nand U13868 (N_13868,N_6048,N_9830);
or U13869 (N_13869,N_7970,N_6061);
or U13870 (N_13870,N_6366,N_9360);
nand U13871 (N_13871,N_7082,N_9875);
xor U13872 (N_13872,N_9882,N_7635);
xor U13873 (N_13873,N_5617,N_6701);
or U13874 (N_13874,N_8953,N_8172);
nor U13875 (N_13875,N_6351,N_7440);
xor U13876 (N_13876,N_7512,N_6376);
and U13877 (N_13877,N_5801,N_8313);
nand U13878 (N_13878,N_7219,N_8043);
nor U13879 (N_13879,N_8158,N_5228);
and U13880 (N_13880,N_8071,N_7800);
nand U13881 (N_13881,N_7688,N_5297);
or U13882 (N_13882,N_9428,N_9061);
nand U13883 (N_13883,N_8222,N_9529);
nor U13884 (N_13884,N_5480,N_5215);
xnor U13885 (N_13885,N_9792,N_5636);
or U13886 (N_13886,N_9388,N_7640);
or U13887 (N_13887,N_8590,N_9843);
nand U13888 (N_13888,N_9976,N_9522);
xor U13889 (N_13889,N_8359,N_7917);
nor U13890 (N_13890,N_6194,N_9206);
and U13891 (N_13891,N_8640,N_9479);
and U13892 (N_13892,N_9725,N_9360);
nor U13893 (N_13893,N_5210,N_6833);
xnor U13894 (N_13894,N_5632,N_7672);
xor U13895 (N_13895,N_6456,N_9879);
and U13896 (N_13896,N_7023,N_9742);
nand U13897 (N_13897,N_9449,N_8493);
or U13898 (N_13898,N_6026,N_7244);
and U13899 (N_13899,N_7815,N_9597);
or U13900 (N_13900,N_6673,N_6240);
and U13901 (N_13901,N_5410,N_5674);
or U13902 (N_13902,N_9084,N_5912);
nand U13903 (N_13903,N_7510,N_6669);
or U13904 (N_13904,N_7212,N_9074);
xor U13905 (N_13905,N_6658,N_8721);
and U13906 (N_13906,N_7057,N_9506);
nand U13907 (N_13907,N_9545,N_7004);
nor U13908 (N_13908,N_8966,N_7504);
nand U13909 (N_13909,N_7986,N_8384);
nand U13910 (N_13910,N_7502,N_8328);
nor U13911 (N_13911,N_8676,N_6266);
nand U13912 (N_13912,N_7093,N_8538);
nor U13913 (N_13913,N_5631,N_8870);
xor U13914 (N_13914,N_5184,N_7153);
and U13915 (N_13915,N_6728,N_7541);
nor U13916 (N_13916,N_5781,N_5946);
nor U13917 (N_13917,N_5328,N_5830);
xnor U13918 (N_13918,N_6648,N_6103);
nor U13919 (N_13919,N_6203,N_9419);
or U13920 (N_13920,N_5646,N_9991);
nor U13921 (N_13921,N_5077,N_8285);
nand U13922 (N_13922,N_6765,N_7530);
xnor U13923 (N_13923,N_5626,N_5829);
nor U13924 (N_13924,N_8465,N_8261);
nor U13925 (N_13925,N_5651,N_6718);
nand U13926 (N_13926,N_6758,N_9441);
and U13927 (N_13927,N_6645,N_9513);
and U13928 (N_13928,N_8657,N_6204);
nor U13929 (N_13929,N_8837,N_6453);
nor U13930 (N_13930,N_9857,N_9400);
nor U13931 (N_13931,N_5314,N_9435);
and U13932 (N_13932,N_8637,N_5216);
and U13933 (N_13933,N_5864,N_6985);
nand U13934 (N_13934,N_5293,N_5278);
or U13935 (N_13935,N_8063,N_6563);
or U13936 (N_13936,N_8228,N_7584);
xor U13937 (N_13937,N_5367,N_9334);
xnor U13938 (N_13938,N_7156,N_8975);
xor U13939 (N_13939,N_6085,N_6227);
nor U13940 (N_13940,N_7588,N_6914);
nand U13941 (N_13941,N_7739,N_6107);
xnor U13942 (N_13942,N_5142,N_5567);
xor U13943 (N_13943,N_9482,N_7395);
nor U13944 (N_13944,N_9833,N_8645);
and U13945 (N_13945,N_6793,N_6586);
xnor U13946 (N_13946,N_9026,N_6665);
xnor U13947 (N_13947,N_9645,N_8767);
nand U13948 (N_13948,N_5928,N_7972);
xor U13949 (N_13949,N_9286,N_6764);
nor U13950 (N_13950,N_9319,N_9028);
nand U13951 (N_13951,N_6978,N_6252);
nand U13952 (N_13952,N_9197,N_7425);
or U13953 (N_13953,N_8271,N_7443);
and U13954 (N_13954,N_6166,N_6950);
nor U13955 (N_13955,N_9389,N_6392);
nor U13956 (N_13956,N_7620,N_5038);
xor U13957 (N_13957,N_8336,N_7814);
xor U13958 (N_13958,N_6330,N_7160);
and U13959 (N_13959,N_9345,N_8261);
or U13960 (N_13960,N_6223,N_7429);
xnor U13961 (N_13961,N_9011,N_8472);
and U13962 (N_13962,N_9060,N_9550);
and U13963 (N_13963,N_5399,N_9734);
and U13964 (N_13964,N_9103,N_5158);
nand U13965 (N_13965,N_5660,N_7359);
xnor U13966 (N_13966,N_5231,N_9536);
or U13967 (N_13967,N_6483,N_8145);
and U13968 (N_13968,N_9623,N_5284);
nor U13969 (N_13969,N_5971,N_6035);
nand U13970 (N_13970,N_9625,N_9300);
nor U13971 (N_13971,N_5395,N_9615);
xor U13972 (N_13972,N_6141,N_8518);
xnor U13973 (N_13973,N_6434,N_8766);
and U13974 (N_13974,N_9102,N_9518);
nor U13975 (N_13975,N_5627,N_5113);
nor U13976 (N_13976,N_5157,N_5963);
nand U13977 (N_13977,N_8809,N_7833);
xnor U13978 (N_13978,N_5750,N_7427);
nand U13979 (N_13979,N_6079,N_7554);
or U13980 (N_13980,N_9793,N_9957);
and U13981 (N_13981,N_6272,N_6630);
xor U13982 (N_13982,N_7235,N_5213);
and U13983 (N_13983,N_8156,N_7947);
nor U13984 (N_13984,N_9383,N_9615);
nand U13985 (N_13985,N_5042,N_5090);
or U13986 (N_13986,N_5690,N_8929);
and U13987 (N_13987,N_8826,N_6060);
nor U13988 (N_13988,N_8778,N_6163);
nor U13989 (N_13989,N_8480,N_6753);
or U13990 (N_13990,N_8807,N_5595);
nand U13991 (N_13991,N_6240,N_5786);
xnor U13992 (N_13992,N_7887,N_6458);
xnor U13993 (N_13993,N_5242,N_5180);
nand U13994 (N_13994,N_5090,N_8034);
and U13995 (N_13995,N_7711,N_9909);
and U13996 (N_13996,N_8613,N_7354);
nor U13997 (N_13997,N_6184,N_7991);
or U13998 (N_13998,N_5150,N_8216);
and U13999 (N_13999,N_9699,N_8891);
or U14000 (N_14000,N_9211,N_9728);
nor U14001 (N_14001,N_7609,N_9370);
or U14002 (N_14002,N_6996,N_9049);
and U14003 (N_14003,N_9897,N_5630);
and U14004 (N_14004,N_8785,N_7059);
xor U14005 (N_14005,N_8329,N_5228);
nand U14006 (N_14006,N_9087,N_7072);
or U14007 (N_14007,N_7257,N_9205);
or U14008 (N_14008,N_9111,N_9903);
and U14009 (N_14009,N_7633,N_7986);
nor U14010 (N_14010,N_8595,N_9329);
nand U14011 (N_14011,N_6147,N_5381);
or U14012 (N_14012,N_8841,N_5321);
nand U14013 (N_14013,N_8573,N_9808);
nor U14014 (N_14014,N_6500,N_7937);
nand U14015 (N_14015,N_5954,N_7509);
or U14016 (N_14016,N_8366,N_7936);
xnor U14017 (N_14017,N_7307,N_8122);
and U14018 (N_14018,N_5771,N_5276);
nor U14019 (N_14019,N_5099,N_8406);
nor U14020 (N_14020,N_9915,N_9626);
xor U14021 (N_14021,N_7013,N_5177);
nor U14022 (N_14022,N_5712,N_6978);
nand U14023 (N_14023,N_8956,N_9434);
nand U14024 (N_14024,N_7372,N_5018);
nand U14025 (N_14025,N_8375,N_7538);
or U14026 (N_14026,N_5945,N_5676);
nand U14027 (N_14027,N_7673,N_6842);
xnor U14028 (N_14028,N_8146,N_7420);
and U14029 (N_14029,N_8619,N_5834);
or U14030 (N_14030,N_5144,N_8646);
xnor U14031 (N_14031,N_6963,N_7569);
xor U14032 (N_14032,N_8133,N_9606);
and U14033 (N_14033,N_8629,N_5743);
and U14034 (N_14034,N_6552,N_7170);
nand U14035 (N_14035,N_5151,N_5782);
nand U14036 (N_14036,N_7248,N_7835);
and U14037 (N_14037,N_9188,N_5220);
nor U14038 (N_14038,N_9384,N_5570);
or U14039 (N_14039,N_7735,N_8999);
nor U14040 (N_14040,N_6954,N_5984);
nor U14041 (N_14041,N_5579,N_6944);
or U14042 (N_14042,N_5567,N_9531);
or U14043 (N_14043,N_6769,N_8316);
and U14044 (N_14044,N_5218,N_6795);
and U14045 (N_14045,N_9264,N_9738);
nand U14046 (N_14046,N_7267,N_7735);
xor U14047 (N_14047,N_5513,N_7781);
nand U14048 (N_14048,N_9607,N_8889);
nand U14049 (N_14049,N_8791,N_6953);
nor U14050 (N_14050,N_9812,N_8892);
or U14051 (N_14051,N_8359,N_6208);
xnor U14052 (N_14052,N_9484,N_5086);
and U14053 (N_14053,N_6798,N_7773);
or U14054 (N_14054,N_7261,N_9248);
or U14055 (N_14055,N_5103,N_9709);
or U14056 (N_14056,N_8616,N_7236);
nand U14057 (N_14057,N_7503,N_6962);
or U14058 (N_14058,N_8471,N_5471);
nor U14059 (N_14059,N_6420,N_8881);
xnor U14060 (N_14060,N_5576,N_7683);
nand U14061 (N_14061,N_7121,N_7579);
nand U14062 (N_14062,N_9310,N_7787);
or U14063 (N_14063,N_8861,N_7828);
xor U14064 (N_14064,N_7793,N_7021);
and U14065 (N_14065,N_5034,N_6497);
and U14066 (N_14066,N_5030,N_8313);
or U14067 (N_14067,N_7953,N_5837);
or U14068 (N_14068,N_6983,N_7825);
nand U14069 (N_14069,N_8272,N_6058);
nor U14070 (N_14070,N_7349,N_8241);
nor U14071 (N_14071,N_5807,N_9919);
nor U14072 (N_14072,N_7314,N_9280);
nor U14073 (N_14073,N_9263,N_6780);
xnor U14074 (N_14074,N_7849,N_9027);
or U14075 (N_14075,N_7077,N_6633);
xor U14076 (N_14076,N_7270,N_6097);
nor U14077 (N_14077,N_8370,N_6803);
xor U14078 (N_14078,N_7750,N_8367);
nor U14079 (N_14079,N_5397,N_8731);
and U14080 (N_14080,N_9049,N_8969);
and U14081 (N_14081,N_6485,N_7028);
xnor U14082 (N_14082,N_9628,N_7408);
and U14083 (N_14083,N_5132,N_7514);
xor U14084 (N_14084,N_7951,N_6546);
or U14085 (N_14085,N_7827,N_5969);
and U14086 (N_14086,N_7602,N_7830);
xor U14087 (N_14087,N_7725,N_8255);
nand U14088 (N_14088,N_6224,N_6386);
or U14089 (N_14089,N_7564,N_8989);
and U14090 (N_14090,N_7079,N_5659);
nand U14091 (N_14091,N_6080,N_9558);
nor U14092 (N_14092,N_8273,N_9465);
xor U14093 (N_14093,N_5373,N_8305);
or U14094 (N_14094,N_5695,N_5441);
nand U14095 (N_14095,N_7322,N_7578);
nor U14096 (N_14096,N_5380,N_7227);
and U14097 (N_14097,N_5650,N_6897);
and U14098 (N_14098,N_7642,N_6841);
and U14099 (N_14099,N_5785,N_7438);
nor U14100 (N_14100,N_7040,N_6142);
nor U14101 (N_14101,N_5509,N_5659);
or U14102 (N_14102,N_7075,N_8184);
xor U14103 (N_14103,N_7732,N_6253);
xnor U14104 (N_14104,N_5228,N_7053);
and U14105 (N_14105,N_9869,N_6646);
xnor U14106 (N_14106,N_6116,N_7945);
nor U14107 (N_14107,N_8113,N_5544);
or U14108 (N_14108,N_6832,N_9650);
nand U14109 (N_14109,N_7509,N_6032);
and U14110 (N_14110,N_6607,N_5623);
nand U14111 (N_14111,N_7419,N_7076);
or U14112 (N_14112,N_5538,N_6886);
and U14113 (N_14113,N_5623,N_6422);
nand U14114 (N_14114,N_8542,N_9714);
nand U14115 (N_14115,N_8983,N_9901);
xor U14116 (N_14116,N_6969,N_6193);
nand U14117 (N_14117,N_5529,N_8223);
and U14118 (N_14118,N_9677,N_9166);
or U14119 (N_14119,N_8013,N_5099);
nor U14120 (N_14120,N_5077,N_6849);
nand U14121 (N_14121,N_7153,N_6366);
xor U14122 (N_14122,N_9983,N_7122);
and U14123 (N_14123,N_6044,N_7506);
nand U14124 (N_14124,N_7747,N_8741);
and U14125 (N_14125,N_7951,N_9237);
and U14126 (N_14126,N_6707,N_8792);
or U14127 (N_14127,N_7761,N_9558);
nor U14128 (N_14128,N_6987,N_8854);
or U14129 (N_14129,N_9481,N_5420);
and U14130 (N_14130,N_9236,N_9900);
nand U14131 (N_14131,N_7085,N_6213);
nor U14132 (N_14132,N_5134,N_9521);
or U14133 (N_14133,N_9485,N_5455);
xor U14134 (N_14134,N_8109,N_6343);
xor U14135 (N_14135,N_5599,N_6777);
xnor U14136 (N_14136,N_6406,N_5090);
xnor U14137 (N_14137,N_5874,N_8370);
and U14138 (N_14138,N_8140,N_6028);
or U14139 (N_14139,N_5387,N_7817);
and U14140 (N_14140,N_6068,N_5743);
and U14141 (N_14141,N_8369,N_9060);
and U14142 (N_14142,N_8476,N_6397);
nand U14143 (N_14143,N_7840,N_5065);
nor U14144 (N_14144,N_5540,N_7372);
nand U14145 (N_14145,N_6269,N_8307);
or U14146 (N_14146,N_6146,N_8978);
xnor U14147 (N_14147,N_6528,N_8745);
and U14148 (N_14148,N_5058,N_7036);
xor U14149 (N_14149,N_7769,N_6375);
nor U14150 (N_14150,N_9061,N_6342);
nand U14151 (N_14151,N_7152,N_8988);
nand U14152 (N_14152,N_6499,N_7047);
nor U14153 (N_14153,N_5404,N_5579);
and U14154 (N_14154,N_7213,N_9957);
or U14155 (N_14155,N_7051,N_6419);
nand U14156 (N_14156,N_5539,N_8217);
and U14157 (N_14157,N_6814,N_6111);
and U14158 (N_14158,N_6045,N_9094);
nor U14159 (N_14159,N_6908,N_8300);
nor U14160 (N_14160,N_6551,N_5726);
xor U14161 (N_14161,N_6780,N_6726);
and U14162 (N_14162,N_7888,N_6102);
nor U14163 (N_14163,N_6351,N_7466);
nor U14164 (N_14164,N_7078,N_6506);
or U14165 (N_14165,N_9251,N_5964);
and U14166 (N_14166,N_9030,N_8298);
nor U14167 (N_14167,N_6327,N_8404);
nand U14168 (N_14168,N_6638,N_7979);
nand U14169 (N_14169,N_5415,N_5859);
nor U14170 (N_14170,N_5743,N_8361);
nand U14171 (N_14171,N_6369,N_6233);
xnor U14172 (N_14172,N_5997,N_9020);
or U14173 (N_14173,N_9498,N_7673);
and U14174 (N_14174,N_5282,N_6282);
xor U14175 (N_14175,N_8842,N_5131);
xnor U14176 (N_14176,N_5273,N_7442);
nand U14177 (N_14177,N_6039,N_7226);
xor U14178 (N_14178,N_9984,N_7003);
xnor U14179 (N_14179,N_5381,N_7479);
nor U14180 (N_14180,N_5129,N_5894);
and U14181 (N_14181,N_9228,N_6541);
nand U14182 (N_14182,N_5606,N_7736);
or U14183 (N_14183,N_9368,N_5779);
xnor U14184 (N_14184,N_8438,N_9110);
or U14185 (N_14185,N_7577,N_5000);
nor U14186 (N_14186,N_7076,N_9167);
nor U14187 (N_14187,N_5811,N_9904);
xor U14188 (N_14188,N_8068,N_5827);
nand U14189 (N_14189,N_7747,N_9164);
xnor U14190 (N_14190,N_7926,N_9516);
nand U14191 (N_14191,N_8729,N_5387);
xor U14192 (N_14192,N_8134,N_9280);
and U14193 (N_14193,N_5399,N_6058);
and U14194 (N_14194,N_6250,N_6472);
xor U14195 (N_14195,N_7094,N_5594);
and U14196 (N_14196,N_7528,N_8451);
nand U14197 (N_14197,N_7726,N_9316);
and U14198 (N_14198,N_6907,N_6556);
nand U14199 (N_14199,N_5197,N_5798);
and U14200 (N_14200,N_7497,N_9045);
xnor U14201 (N_14201,N_5167,N_8321);
nand U14202 (N_14202,N_8136,N_8052);
nand U14203 (N_14203,N_7563,N_8268);
xor U14204 (N_14204,N_9906,N_6305);
nor U14205 (N_14205,N_5168,N_5332);
and U14206 (N_14206,N_8337,N_8073);
or U14207 (N_14207,N_9066,N_7222);
nand U14208 (N_14208,N_7072,N_6199);
nand U14209 (N_14209,N_5736,N_8124);
and U14210 (N_14210,N_5276,N_5899);
nand U14211 (N_14211,N_7648,N_8632);
xor U14212 (N_14212,N_6907,N_8078);
nor U14213 (N_14213,N_8110,N_9061);
xor U14214 (N_14214,N_9017,N_6973);
and U14215 (N_14215,N_8267,N_5866);
and U14216 (N_14216,N_7746,N_8222);
nand U14217 (N_14217,N_7912,N_6924);
and U14218 (N_14218,N_5095,N_9014);
and U14219 (N_14219,N_9474,N_7585);
xor U14220 (N_14220,N_7300,N_5699);
xor U14221 (N_14221,N_5668,N_9684);
nor U14222 (N_14222,N_8641,N_6632);
nand U14223 (N_14223,N_7908,N_6180);
and U14224 (N_14224,N_6115,N_9655);
xnor U14225 (N_14225,N_7338,N_7992);
and U14226 (N_14226,N_8088,N_7798);
nand U14227 (N_14227,N_9992,N_8432);
nor U14228 (N_14228,N_8576,N_7207);
and U14229 (N_14229,N_5198,N_6450);
or U14230 (N_14230,N_9918,N_9196);
nand U14231 (N_14231,N_7129,N_9640);
and U14232 (N_14232,N_8009,N_5835);
nor U14233 (N_14233,N_7214,N_9122);
xnor U14234 (N_14234,N_5032,N_5661);
and U14235 (N_14235,N_9928,N_7896);
or U14236 (N_14236,N_6420,N_6806);
nor U14237 (N_14237,N_7950,N_9365);
nand U14238 (N_14238,N_6075,N_7154);
and U14239 (N_14239,N_7378,N_7924);
and U14240 (N_14240,N_7529,N_8921);
nor U14241 (N_14241,N_5500,N_8724);
nor U14242 (N_14242,N_6222,N_7824);
xnor U14243 (N_14243,N_6831,N_6867);
or U14244 (N_14244,N_6453,N_8156);
xor U14245 (N_14245,N_9823,N_9581);
xnor U14246 (N_14246,N_5965,N_8614);
or U14247 (N_14247,N_6207,N_6090);
nand U14248 (N_14248,N_7583,N_7790);
or U14249 (N_14249,N_6732,N_6948);
nand U14250 (N_14250,N_6635,N_6491);
nand U14251 (N_14251,N_9863,N_7160);
xnor U14252 (N_14252,N_5036,N_8841);
and U14253 (N_14253,N_5500,N_6576);
xnor U14254 (N_14254,N_7155,N_9604);
and U14255 (N_14255,N_7408,N_5184);
nor U14256 (N_14256,N_5671,N_6689);
nor U14257 (N_14257,N_5313,N_7257);
or U14258 (N_14258,N_7456,N_6906);
nor U14259 (N_14259,N_6372,N_6388);
nand U14260 (N_14260,N_9735,N_8100);
nand U14261 (N_14261,N_5800,N_9946);
nor U14262 (N_14262,N_5573,N_5613);
or U14263 (N_14263,N_8208,N_8835);
nand U14264 (N_14264,N_7667,N_5113);
or U14265 (N_14265,N_5278,N_8620);
nand U14266 (N_14266,N_5060,N_8848);
xnor U14267 (N_14267,N_5720,N_6040);
nand U14268 (N_14268,N_5013,N_8130);
xnor U14269 (N_14269,N_7550,N_8233);
nor U14270 (N_14270,N_5308,N_9821);
or U14271 (N_14271,N_6902,N_6465);
or U14272 (N_14272,N_9482,N_8163);
nor U14273 (N_14273,N_7855,N_7913);
nor U14274 (N_14274,N_7595,N_5995);
and U14275 (N_14275,N_6170,N_7404);
and U14276 (N_14276,N_7239,N_7391);
and U14277 (N_14277,N_7200,N_5450);
nor U14278 (N_14278,N_5603,N_7536);
nand U14279 (N_14279,N_7833,N_5611);
xnor U14280 (N_14280,N_6635,N_5865);
or U14281 (N_14281,N_6016,N_9215);
and U14282 (N_14282,N_8226,N_8077);
nand U14283 (N_14283,N_8143,N_9673);
nand U14284 (N_14284,N_7042,N_5813);
or U14285 (N_14285,N_8321,N_5341);
nor U14286 (N_14286,N_8886,N_5107);
nor U14287 (N_14287,N_9911,N_8497);
nand U14288 (N_14288,N_8881,N_7516);
or U14289 (N_14289,N_9462,N_9698);
and U14290 (N_14290,N_7935,N_5301);
or U14291 (N_14291,N_9079,N_9346);
nand U14292 (N_14292,N_5508,N_8151);
or U14293 (N_14293,N_7389,N_6058);
nor U14294 (N_14294,N_9146,N_8925);
nand U14295 (N_14295,N_5466,N_8591);
and U14296 (N_14296,N_9508,N_7338);
and U14297 (N_14297,N_5267,N_9291);
nand U14298 (N_14298,N_6609,N_9531);
and U14299 (N_14299,N_9011,N_6089);
nor U14300 (N_14300,N_7469,N_7921);
nor U14301 (N_14301,N_7477,N_5233);
nor U14302 (N_14302,N_8738,N_9183);
xnor U14303 (N_14303,N_8744,N_9317);
or U14304 (N_14304,N_6344,N_6449);
nand U14305 (N_14305,N_9393,N_7136);
nor U14306 (N_14306,N_8621,N_9677);
and U14307 (N_14307,N_7797,N_9527);
and U14308 (N_14308,N_9111,N_8328);
and U14309 (N_14309,N_7034,N_9161);
nor U14310 (N_14310,N_9123,N_6746);
and U14311 (N_14311,N_8562,N_5088);
nor U14312 (N_14312,N_5539,N_9382);
and U14313 (N_14313,N_8862,N_5538);
or U14314 (N_14314,N_6091,N_5533);
or U14315 (N_14315,N_6435,N_8606);
and U14316 (N_14316,N_7881,N_6683);
nor U14317 (N_14317,N_5307,N_5825);
nand U14318 (N_14318,N_8312,N_5937);
nand U14319 (N_14319,N_5231,N_6529);
xor U14320 (N_14320,N_8224,N_8558);
and U14321 (N_14321,N_6459,N_8418);
and U14322 (N_14322,N_6533,N_6468);
or U14323 (N_14323,N_8457,N_7330);
or U14324 (N_14324,N_6286,N_7647);
nor U14325 (N_14325,N_7564,N_8238);
nand U14326 (N_14326,N_9261,N_5988);
xnor U14327 (N_14327,N_7247,N_6857);
nand U14328 (N_14328,N_9628,N_7506);
or U14329 (N_14329,N_7567,N_6743);
nand U14330 (N_14330,N_5998,N_5355);
and U14331 (N_14331,N_7250,N_6576);
nor U14332 (N_14332,N_9584,N_5888);
nand U14333 (N_14333,N_9774,N_9452);
or U14334 (N_14334,N_8961,N_8200);
nand U14335 (N_14335,N_7648,N_9561);
and U14336 (N_14336,N_6981,N_7448);
and U14337 (N_14337,N_7314,N_7303);
and U14338 (N_14338,N_7848,N_8900);
nand U14339 (N_14339,N_9667,N_8431);
xor U14340 (N_14340,N_7280,N_5525);
xnor U14341 (N_14341,N_6944,N_5692);
and U14342 (N_14342,N_9055,N_6127);
nand U14343 (N_14343,N_9406,N_7120);
xnor U14344 (N_14344,N_7094,N_5699);
nor U14345 (N_14345,N_7370,N_6860);
nor U14346 (N_14346,N_8836,N_8983);
nand U14347 (N_14347,N_8497,N_8723);
nand U14348 (N_14348,N_8680,N_7973);
or U14349 (N_14349,N_5046,N_6543);
nand U14350 (N_14350,N_8312,N_5722);
nor U14351 (N_14351,N_6393,N_6097);
nor U14352 (N_14352,N_5664,N_8396);
or U14353 (N_14353,N_9550,N_6327);
xnor U14354 (N_14354,N_7282,N_5288);
or U14355 (N_14355,N_7304,N_5943);
nor U14356 (N_14356,N_8258,N_5646);
nor U14357 (N_14357,N_8609,N_9594);
and U14358 (N_14358,N_5913,N_5573);
nand U14359 (N_14359,N_8329,N_6573);
nor U14360 (N_14360,N_7101,N_9232);
xnor U14361 (N_14361,N_6120,N_7715);
nor U14362 (N_14362,N_5010,N_7080);
xor U14363 (N_14363,N_6848,N_6914);
and U14364 (N_14364,N_6033,N_6077);
xnor U14365 (N_14365,N_6057,N_6159);
nor U14366 (N_14366,N_5978,N_5953);
xnor U14367 (N_14367,N_5250,N_5790);
nor U14368 (N_14368,N_7471,N_7596);
nand U14369 (N_14369,N_8146,N_6515);
and U14370 (N_14370,N_6258,N_5099);
nor U14371 (N_14371,N_9232,N_6951);
nand U14372 (N_14372,N_6502,N_8003);
nand U14373 (N_14373,N_8660,N_7489);
nor U14374 (N_14374,N_6763,N_9728);
xor U14375 (N_14375,N_7735,N_7378);
or U14376 (N_14376,N_7477,N_5235);
or U14377 (N_14377,N_7947,N_6769);
and U14378 (N_14378,N_7117,N_9859);
nor U14379 (N_14379,N_6574,N_8148);
nor U14380 (N_14380,N_5005,N_9859);
nand U14381 (N_14381,N_7097,N_7492);
and U14382 (N_14382,N_7454,N_5904);
and U14383 (N_14383,N_5414,N_7285);
and U14384 (N_14384,N_6566,N_9233);
xor U14385 (N_14385,N_5491,N_7878);
xnor U14386 (N_14386,N_6334,N_6904);
nor U14387 (N_14387,N_8746,N_9779);
or U14388 (N_14388,N_6066,N_9910);
xnor U14389 (N_14389,N_5976,N_5265);
or U14390 (N_14390,N_9021,N_9339);
nand U14391 (N_14391,N_8813,N_7382);
and U14392 (N_14392,N_9258,N_6853);
and U14393 (N_14393,N_6129,N_5986);
or U14394 (N_14394,N_9583,N_8850);
nor U14395 (N_14395,N_5663,N_6699);
nand U14396 (N_14396,N_9601,N_8767);
nor U14397 (N_14397,N_9943,N_8247);
nand U14398 (N_14398,N_5896,N_8468);
nand U14399 (N_14399,N_9776,N_5312);
nand U14400 (N_14400,N_6372,N_7809);
xnor U14401 (N_14401,N_8378,N_9526);
and U14402 (N_14402,N_7842,N_6881);
nand U14403 (N_14403,N_8558,N_7848);
or U14404 (N_14404,N_9144,N_6230);
and U14405 (N_14405,N_5895,N_7514);
or U14406 (N_14406,N_9749,N_7963);
xor U14407 (N_14407,N_5380,N_9036);
xor U14408 (N_14408,N_6587,N_9278);
and U14409 (N_14409,N_6746,N_5462);
nand U14410 (N_14410,N_9775,N_8583);
and U14411 (N_14411,N_5565,N_9745);
xnor U14412 (N_14412,N_9511,N_6940);
xor U14413 (N_14413,N_9560,N_5500);
and U14414 (N_14414,N_9872,N_6570);
xnor U14415 (N_14415,N_5340,N_5401);
xor U14416 (N_14416,N_7739,N_6558);
nand U14417 (N_14417,N_6174,N_6134);
nand U14418 (N_14418,N_6181,N_7153);
or U14419 (N_14419,N_6298,N_7875);
xnor U14420 (N_14420,N_6563,N_9362);
and U14421 (N_14421,N_5604,N_7215);
xor U14422 (N_14422,N_7163,N_6704);
xor U14423 (N_14423,N_9669,N_6404);
and U14424 (N_14424,N_5309,N_6350);
or U14425 (N_14425,N_6759,N_6059);
xnor U14426 (N_14426,N_5333,N_7190);
nand U14427 (N_14427,N_8349,N_5751);
nor U14428 (N_14428,N_7457,N_5641);
nor U14429 (N_14429,N_6629,N_5724);
nand U14430 (N_14430,N_7096,N_9268);
nor U14431 (N_14431,N_5044,N_7950);
or U14432 (N_14432,N_6507,N_9689);
and U14433 (N_14433,N_8744,N_5630);
nand U14434 (N_14434,N_6602,N_7872);
nor U14435 (N_14435,N_8018,N_5400);
nand U14436 (N_14436,N_7852,N_6751);
nor U14437 (N_14437,N_8386,N_5054);
nor U14438 (N_14438,N_5783,N_6162);
xnor U14439 (N_14439,N_7008,N_5560);
nand U14440 (N_14440,N_9088,N_5971);
or U14441 (N_14441,N_5354,N_8631);
nor U14442 (N_14442,N_6793,N_8377);
nor U14443 (N_14443,N_7654,N_7481);
nand U14444 (N_14444,N_5062,N_5437);
or U14445 (N_14445,N_7998,N_9158);
nand U14446 (N_14446,N_6835,N_9206);
and U14447 (N_14447,N_5232,N_8942);
xnor U14448 (N_14448,N_9544,N_6210);
nor U14449 (N_14449,N_9156,N_5361);
xnor U14450 (N_14450,N_5710,N_9296);
nor U14451 (N_14451,N_5520,N_5020);
nor U14452 (N_14452,N_8835,N_6441);
nor U14453 (N_14453,N_7232,N_7053);
or U14454 (N_14454,N_7490,N_8491);
or U14455 (N_14455,N_8419,N_6102);
or U14456 (N_14456,N_9572,N_5079);
nand U14457 (N_14457,N_9222,N_5028);
nor U14458 (N_14458,N_8899,N_6982);
or U14459 (N_14459,N_8967,N_9928);
xnor U14460 (N_14460,N_7294,N_9131);
and U14461 (N_14461,N_9932,N_8223);
or U14462 (N_14462,N_8640,N_5259);
or U14463 (N_14463,N_9326,N_6432);
and U14464 (N_14464,N_6420,N_7478);
xor U14465 (N_14465,N_5149,N_9980);
nor U14466 (N_14466,N_8843,N_9774);
or U14467 (N_14467,N_9737,N_5427);
nor U14468 (N_14468,N_7352,N_8326);
nand U14469 (N_14469,N_6511,N_7374);
nor U14470 (N_14470,N_6826,N_7674);
nand U14471 (N_14471,N_5321,N_5309);
nand U14472 (N_14472,N_7736,N_7275);
xor U14473 (N_14473,N_9623,N_7115);
or U14474 (N_14474,N_6805,N_7040);
and U14475 (N_14475,N_5290,N_7652);
nor U14476 (N_14476,N_6960,N_7686);
xnor U14477 (N_14477,N_6424,N_8736);
xnor U14478 (N_14478,N_8594,N_5196);
nand U14479 (N_14479,N_8716,N_6504);
nor U14480 (N_14480,N_6664,N_8204);
xnor U14481 (N_14481,N_7356,N_7871);
and U14482 (N_14482,N_5766,N_9186);
nor U14483 (N_14483,N_7218,N_5601);
xnor U14484 (N_14484,N_9790,N_5942);
and U14485 (N_14485,N_8070,N_8275);
nor U14486 (N_14486,N_7543,N_5045);
xor U14487 (N_14487,N_6811,N_8352);
nor U14488 (N_14488,N_7835,N_7236);
nor U14489 (N_14489,N_7255,N_5404);
or U14490 (N_14490,N_6733,N_7106);
or U14491 (N_14491,N_8598,N_6302);
nor U14492 (N_14492,N_6331,N_6148);
or U14493 (N_14493,N_8917,N_5260);
and U14494 (N_14494,N_9936,N_9526);
nand U14495 (N_14495,N_9733,N_7790);
xnor U14496 (N_14496,N_5296,N_9508);
xor U14497 (N_14497,N_7583,N_7565);
nand U14498 (N_14498,N_8238,N_5733);
and U14499 (N_14499,N_9707,N_8732);
nand U14500 (N_14500,N_7758,N_5088);
nand U14501 (N_14501,N_9072,N_5757);
nand U14502 (N_14502,N_8516,N_7422);
or U14503 (N_14503,N_5957,N_8063);
or U14504 (N_14504,N_9550,N_7585);
or U14505 (N_14505,N_5984,N_9888);
xnor U14506 (N_14506,N_8594,N_7204);
or U14507 (N_14507,N_8122,N_5436);
nand U14508 (N_14508,N_8783,N_5249);
nand U14509 (N_14509,N_8257,N_6460);
nor U14510 (N_14510,N_6367,N_6980);
or U14511 (N_14511,N_9661,N_8915);
and U14512 (N_14512,N_9405,N_7930);
nor U14513 (N_14513,N_5837,N_9536);
and U14514 (N_14514,N_7842,N_8257);
or U14515 (N_14515,N_6681,N_6804);
nor U14516 (N_14516,N_5270,N_7474);
nand U14517 (N_14517,N_9902,N_5612);
nand U14518 (N_14518,N_5706,N_8445);
and U14519 (N_14519,N_7698,N_6640);
nor U14520 (N_14520,N_7367,N_9204);
nor U14521 (N_14521,N_7946,N_8283);
and U14522 (N_14522,N_6631,N_9381);
or U14523 (N_14523,N_5437,N_6294);
nor U14524 (N_14524,N_7503,N_8580);
nor U14525 (N_14525,N_7638,N_9495);
and U14526 (N_14526,N_8686,N_6329);
or U14527 (N_14527,N_8722,N_9554);
xnor U14528 (N_14528,N_8109,N_5115);
and U14529 (N_14529,N_8692,N_9788);
and U14530 (N_14530,N_5011,N_7349);
and U14531 (N_14531,N_9780,N_5985);
or U14532 (N_14532,N_7854,N_6314);
and U14533 (N_14533,N_6195,N_7979);
xnor U14534 (N_14534,N_5043,N_5233);
nor U14535 (N_14535,N_5791,N_5359);
xor U14536 (N_14536,N_5920,N_8943);
or U14537 (N_14537,N_5929,N_9571);
and U14538 (N_14538,N_5573,N_8596);
nor U14539 (N_14539,N_5403,N_8917);
xnor U14540 (N_14540,N_8859,N_5010);
or U14541 (N_14541,N_7456,N_5894);
and U14542 (N_14542,N_8593,N_6501);
and U14543 (N_14543,N_7394,N_6946);
xor U14544 (N_14544,N_5147,N_9568);
nor U14545 (N_14545,N_8603,N_8044);
or U14546 (N_14546,N_8368,N_9490);
nor U14547 (N_14547,N_6045,N_6572);
or U14548 (N_14548,N_9268,N_8613);
xnor U14549 (N_14549,N_5698,N_8762);
xor U14550 (N_14550,N_8709,N_6247);
and U14551 (N_14551,N_9424,N_8358);
nand U14552 (N_14552,N_6736,N_5490);
and U14553 (N_14553,N_8794,N_8791);
and U14554 (N_14554,N_6856,N_7642);
nand U14555 (N_14555,N_8351,N_8792);
xor U14556 (N_14556,N_8671,N_8222);
xor U14557 (N_14557,N_6109,N_7175);
nand U14558 (N_14558,N_8988,N_5384);
or U14559 (N_14559,N_7801,N_7268);
and U14560 (N_14560,N_5644,N_7948);
xor U14561 (N_14561,N_5004,N_7664);
or U14562 (N_14562,N_7601,N_7065);
nor U14563 (N_14563,N_9789,N_6622);
and U14564 (N_14564,N_5470,N_5102);
nand U14565 (N_14565,N_7104,N_9285);
nand U14566 (N_14566,N_6469,N_8272);
xor U14567 (N_14567,N_5422,N_9680);
xnor U14568 (N_14568,N_8807,N_7377);
nand U14569 (N_14569,N_5040,N_6864);
and U14570 (N_14570,N_7876,N_9998);
or U14571 (N_14571,N_8246,N_5108);
nand U14572 (N_14572,N_5655,N_5672);
or U14573 (N_14573,N_6922,N_8406);
nor U14574 (N_14574,N_8922,N_7348);
or U14575 (N_14575,N_5029,N_6220);
nand U14576 (N_14576,N_6843,N_7831);
and U14577 (N_14577,N_6546,N_8998);
and U14578 (N_14578,N_9708,N_5589);
and U14579 (N_14579,N_9686,N_6350);
nand U14580 (N_14580,N_8741,N_9326);
xor U14581 (N_14581,N_6568,N_8048);
nand U14582 (N_14582,N_6580,N_8912);
or U14583 (N_14583,N_7096,N_8087);
nor U14584 (N_14584,N_6690,N_6568);
nand U14585 (N_14585,N_9708,N_7891);
nand U14586 (N_14586,N_5491,N_5216);
xor U14587 (N_14587,N_7097,N_7246);
nand U14588 (N_14588,N_6817,N_5796);
and U14589 (N_14589,N_8662,N_5472);
nand U14590 (N_14590,N_9224,N_7294);
xor U14591 (N_14591,N_8023,N_7887);
nand U14592 (N_14592,N_9120,N_6960);
xnor U14593 (N_14593,N_9258,N_5457);
xor U14594 (N_14594,N_9436,N_6727);
or U14595 (N_14595,N_5560,N_9955);
xor U14596 (N_14596,N_8595,N_5885);
and U14597 (N_14597,N_6105,N_6470);
xor U14598 (N_14598,N_9813,N_6080);
nand U14599 (N_14599,N_7452,N_6918);
or U14600 (N_14600,N_8354,N_6057);
nand U14601 (N_14601,N_8924,N_8366);
xor U14602 (N_14602,N_7021,N_7499);
nor U14603 (N_14603,N_9219,N_8553);
nand U14604 (N_14604,N_8401,N_7869);
or U14605 (N_14605,N_6226,N_5912);
and U14606 (N_14606,N_7258,N_8191);
nand U14607 (N_14607,N_6923,N_6305);
xor U14608 (N_14608,N_9109,N_8195);
and U14609 (N_14609,N_9891,N_8914);
nor U14610 (N_14610,N_5066,N_8944);
and U14611 (N_14611,N_9341,N_6492);
xnor U14612 (N_14612,N_9015,N_7683);
nor U14613 (N_14613,N_7180,N_6307);
and U14614 (N_14614,N_8210,N_9991);
or U14615 (N_14615,N_6119,N_6986);
nand U14616 (N_14616,N_5778,N_9314);
and U14617 (N_14617,N_7686,N_7337);
xnor U14618 (N_14618,N_5060,N_7244);
or U14619 (N_14619,N_8828,N_9489);
nand U14620 (N_14620,N_9986,N_6064);
nor U14621 (N_14621,N_8498,N_6056);
nand U14622 (N_14622,N_9811,N_7508);
or U14623 (N_14623,N_6492,N_8942);
nand U14624 (N_14624,N_7206,N_5273);
nand U14625 (N_14625,N_6796,N_7917);
or U14626 (N_14626,N_6515,N_6615);
or U14627 (N_14627,N_9112,N_9990);
nand U14628 (N_14628,N_7524,N_5103);
xor U14629 (N_14629,N_9715,N_6226);
xor U14630 (N_14630,N_5648,N_9619);
nand U14631 (N_14631,N_6042,N_6120);
and U14632 (N_14632,N_8451,N_7495);
nor U14633 (N_14633,N_6897,N_9082);
nor U14634 (N_14634,N_6503,N_6565);
nand U14635 (N_14635,N_6805,N_5089);
or U14636 (N_14636,N_8275,N_5442);
or U14637 (N_14637,N_5196,N_9095);
nor U14638 (N_14638,N_9952,N_6053);
or U14639 (N_14639,N_7074,N_8347);
xnor U14640 (N_14640,N_7205,N_6132);
nor U14641 (N_14641,N_7329,N_8443);
nand U14642 (N_14642,N_9156,N_7609);
and U14643 (N_14643,N_5630,N_9228);
and U14644 (N_14644,N_7483,N_9222);
or U14645 (N_14645,N_9953,N_9364);
nor U14646 (N_14646,N_5341,N_8894);
and U14647 (N_14647,N_8237,N_8083);
nor U14648 (N_14648,N_7493,N_8727);
nor U14649 (N_14649,N_6068,N_9696);
nor U14650 (N_14650,N_9925,N_6285);
nand U14651 (N_14651,N_9978,N_7862);
xnor U14652 (N_14652,N_6359,N_6005);
nor U14653 (N_14653,N_7308,N_7977);
or U14654 (N_14654,N_6172,N_7222);
nor U14655 (N_14655,N_7345,N_6660);
nand U14656 (N_14656,N_6193,N_5516);
or U14657 (N_14657,N_7098,N_6142);
and U14658 (N_14658,N_8524,N_7362);
or U14659 (N_14659,N_8121,N_8698);
nand U14660 (N_14660,N_9368,N_7940);
nor U14661 (N_14661,N_9599,N_5110);
and U14662 (N_14662,N_6000,N_8500);
or U14663 (N_14663,N_5628,N_7386);
nand U14664 (N_14664,N_8919,N_8365);
nand U14665 (N_14665,N_6883,N_5005);
or U14666 (N_14666,N_6204,N_7850);
and U14667 (N_14667,N_8995,N_7159);
nand U14668 (N_14668,N_8946,N_9056);
and U14669 (N_14669,N_7884,N_9853);
and U14670 (N_14670,N_5626,N_8491);
and U14671 (N_14671,N_5822,N_7182);
nor U14672 (N_14672,N_9870,N_7394);
and U14673 (N_14673,N_5541,N_7110);
nor U14674 (N_14674,N_8159,N_8073);
xor U14675 (N_14675,N_7345,N_5164);
and U14676 (N_14676,N_5502,N_6895);
nand U14677 (N_14677,N_8945,N_7135);
nor U14678 (N_14678,N_9596,N_5351);
and U14679 (N_14679,N_8179,N_7225);
and U14680 (N_14680,N_9572,N_7835);
nand U14681 (N_14681,N_6025,N_6122);
and U14682 (N_14682,N_9913,N_7888);
and U14683 (N_14683,N_8359,N_8392);
nor U14684 (N_14684,N_5513,N_8111);
and U14685 (N_14685,N_5551,N_5130);
and U14686 (N_14686,N_7454,N_7131);
or U14687 (N_14687,N_5477,N_7550);
or U14688 (N_14688,N_9748,N_9727);
nor U14689 (N_14689,N_5304,N_5683);
and U14690 (N_14690,N_5723,N_8790);
or U14691 (N_14691,N_9423,N_9501);
xnor U14692 (N_14692,N_9916,N_8985);
nand U14693 (N_14693,N_7945,N_8655);
or U14694 (N_14694,N_8099,N_6358);
or U14695 (N_14695,N_5235,N_9926);
nand U14696 (N_14696,N_8391,N_5012);
or U14697 (N_14697,N_5900,N_5495);
nand U14698 (N_14698,N_8122,N_7053);
nor U14699 (N_14699,N_7752,N_5039);
nor U14700 (N_14700,N_9178,N_8272);
xnor U14701 (N_14701,N_6143,N_5298);
xnor U14702 (N_14702,N_9764,N_8185);
nand U14703 (N_14703,N_9987,N_6082);
xnor U14704 (N_14704,N_7328,N_7301);
nor U14705 (N_14705,N_9850,N_5391);
or U14706 (N_14706,N_8610,N_7789);
nand U14707 (N_14707,N_9902,N_6536);
nand U14708 (N_14708,N_9739,N_8765);
nand U14709 (N_14709,N_7712,N_5888);
and U14710 (N_14710,N_9290,N_8950);
nor U14711 (N_14711,N_7821,N_9052);
or U14712 (N_14712,N_6293,N_7315);
nand U14713 (N_14713,N_9432,N_6979);
nand U14714 (N_14714,N_6217,N_8352);
nand U14715 (N_14715,N_9540,N_8002);
nand U14716 (N_14716,N_8895,N_5738);
nor U14717 (N_14717,N_6805,N_7748);
nand U14718 (N_14718,N_6103,N_5628);
xnor U14719 (N_14719,N_8679,N_6273);
and U14720 (N_14720,N_5005,N_9782);
xnor U14721 (N_14721,N_5524,N_9546);
or U14722 (N_14722,N_8920,N_5821);
and U14723 (N_14723,N_9554,N_9191);
xor U14724 (N_14724,N_6388,N_7091);
xnor U14725 (N_14725,N_8331,N_7279);
or U14726 (N_14726,N_8374,N_7393);
and U14727 (N_14727,N_5459,N_8620);
and U14728 (N_14728,N_8129,N_5293);
nor U14729 (N_14729,N_6102,N_9690);
nor U14730 (N_14730,N_5962,N_5663);
or U14731 (N_14731,N_5537,N_9428);
and U14732 (N_14732,N_9097,N_5589);
nor U14733 (N_14733,N_9163,N_6044);
and U14734 (N_14734,N_9939,N_6153);
nor U14735 (N_14735,N_6826,N_9356);
nor U14736 (N_14736,N_6087,N_6871);
nor U14737 (N_14737,N_8188,N_6470);
xnor U14738 (N_14738,N_5175,N_7700);
nor U14739 (N_14739,N_9966,N_6173);
or U14740 (N_14740,N_9790,N_8511);
and U14741 (N_14741,N_5842,N_5599);
and U14742 (N_14742,N_6783,N_5635);
and U14743 (N_14743,N_9115,N_9801);
or U14744 (N_14744,N_9904,N_5694);
nor U14745 (N_14745,N_7592,N_8696);
nand U14746 (N_14746,N_7878,N_8821);
xnor U14747 (N_14747,N_6590,N_5928);
and U14748 (N_14748,N_5299,N_5507);
and U14749 (N_14749,N_8095,N_6646);
nor U14750 (N_14750,N_7611,N_7317);
xnor U14751 (N_14751,N_7309,N_8342);
nand U14752 (N_14752,N_7114,N_6517);
and U14753 (N_14753,N_8043,N_5122);
nor U14754 (N_14754,N_7304,N_7231);
or U14755 (N_14755,N_6965,N_7559);
nand U14756 (N_14756,N_5168,N_5890);
or U14757 (N_14757,N_7472,N_8369);
and U14758 (N_14758,N_9944,N_7920);
nand U14759 (N_14759,N_5113,N_6673);
nand U14760 (N_14760,N_7678,N_7260);
and U14761 (N_14761,N_8083,N_8974);
or U14762 (N_14762,N_7242,N_9673);
or U14763 (N_14763,N_6535,N_7643);
xor U14764 (N_14764,N_8911,N_9211);
xor U14765 (N_14765,N_9589,N_8755);
and U14766 (N_14766,N_5004,N_9446);
xnor U14767 (N_14767,N_9994,N_6682);
or U14768 (N_14768,N_7472,N_7537);
nand U14769 (N_14769,N_7143,N_8618);
nand U14770 (N_14770,N_6645,N_7844);
nor U14771 (N_14771,N_8284,N_5504);
xnor U14772 (N_14772,N_9676,N_8156);
xor U14773 (N_14773,N_6714,N_8812);
or U14774 (N_14774,N_8162,N_8772);
nor U14775 (N_14775,N_8016,N_9276);
nand U14776 (N_14776,N_9101,N_9198);
nand U14777 (N_14777,N_5272,N_6184);
or U14778 (N_14778,N_7881,N_7563);
nand U14779 (N_14779,N_7576,N_9982);
xnor U14780 (N_14780,N_5248,N_8971);
nor U14781 (N_14781,N_8370,N_6314);
nand U14782 (N_14782,N_7899,N_9159);
or U14783 (N_14783,N_9331,N_8761);
or U14784 (N_14784,N_6239,N_5607);
nand U14785 (N_14785,N_9769,N_9973);
nor U14786 (N_14786,N_8925,N_9547);
and U14787 (N_14787,N_6851,N_5046);
nand U14788 (N_14788,N_9661,N_8762);
and U14789 (N_14789,N_9554,N_7196);
nor U14790 (N_14790,N_6562,N_9391);
and U14791 (N_14791,N_8798,N_8299);
or U14792 (N_14792,N_9353,N_8635);
nor U14793 (N_14793,N_8740,N_7771);
or U14794 (N_14794,N_6389,N_5234);
xnor U14795 (N_14795,N_9409,N_9009);
and U14796 (N_14796,N_7623,N_6295);
nor U14797 (N_14797,N_7630,N_8542);
or U14798 (N_14798,N_7302,N_7315);
or U14799 (N_14799,N_6926,N_6538);
xor U14800 (N_14800,N_6191,N_9936);
nand U14801 (N_14801,N_9844,N_8172);
nand U14802 (N_14802,N_5161,N_8161);
nand U14803 (N_14803,N_5790,N_9456);
and U14804 (N_14804,N_8174,N_6258);
xor U14805 (N_14805,N_7417,N_5574);
nor U14806 (N_14806,N_6842,N_6796);
xor U14807 (N_14807,N_7579,N_5014);
and U14808 (N_14808,N_6402,N_7890);
xor U14809 (N_14809,N_7081,N_9536);
xor U14810 (N_14810,N_9806,N_8780);
nor U14811 (N_14811,N_8493,N_8149);
nand U14812 (N_14812,N_7238,N_9728);
nor U14813 (N_14813,N_6457,N_5493);
and U14814 (N_14814,N_7870,N_7061);
xnor U14815 (N_14815,N_6450,N_8332);
nor U14816 (N_14816,N_8025,N_6148);
or U14817 (N_14817,N_5494,N_5991);
or U14818 (N_14818,N_9770,N_6572);
xnor U14819 (N_14819,N_5703,N_7592);
or U14820 (N_14820,N_5807,N_6814);
xor U14821 (N_14821,N_8576,N_9805);
or U14822 (N_14822,N_5155,N_7532);
nand U14823 (N_14823,N_7201,N_9514);
and U14824 (N_14824,N_7028,N_9223);
nand U14825 (N_14825,N_6713,N_5791);
nand U14826 (N_14826,N_8073,N_5703);
nand U14827 (N_14827,N_9129,N_6493);
nor U14828 (N_14828,N_8056,N_9886);
nor U14829 (N_14829,N_8615,N_9754);
or U14830 (N_14830,N_7330,N_5529);
xnor U14831 (N_14831,N_7937,N_9393);
xnor U14832 (N_14832,N_9756,N_5964);
nor U14833 (N_14833,N_5776,N_8078);
xnor U14834 (N_14834,N_5898,N_5626);
nand U14835 (N_14835,N_9191,N_6244);
or U14836 (N_14836,N_7363,N_8478);
nor U14837 (N_14837,N_9070,N_9220);
nor U14838 (N_14838,N_7130,N_8107);
xnor U14839 (N_14839,N_7983,N_8768);
and U14840 (N_14840,N_6213,N_8677);
or U14841 (N_14841,N_8519,N_9509);
nor U14842 (N_14842,N_5829,N_8133);
and U14843 (N_14843,N_6051,N_7989);
xor U14844 (N_14844,N_9722,N_7445);
nor U14845 (N_14845,N_8354,N_5902);
xor U14846 (N_14846,N_8850,N_6092);
or U14847 (N_14847,N_7671,N_5883);
xnor U14848 (N_14848,N_7552,N_8358);
nand U14849 (N_14849,N_5248,N_7587);
nand U14850 (N_14850,N_9131,N_9442);
xor U14851 (N_14851,N_6809,N_7670);
and U14852 (N_14852,N_8989,N_5304);
nand U14853 (N_14853,N_6292,N_9273);
nor U14854 (N_14854,N_7566,N_7396);
xnor U14855 (N_14855,N_8751,N_5949);
nand U14856 (N_14856,N_7284,N_9187);
nand U14857 (N_14857,N_5571,N_5207);
and U14858 (N_14858,N_9325,N_6171);
xnor U14859 (N_14859,N_6332,N_9668);
nand U14860 (N_14860,N_5646,N_6721);
nand U14861 (N_14861,N_6791,N_7538);
and U14862 (N_14862,N_7989,N_6540);
xor U14863 (N_14863,N_7971,N_8133);
xor U14864 (N_14864,N_7943,N_9603);
and U14865 (N_14865,N_9850,N_6556);
or U14866 (N_14866,N_6067,N_5084);
and U14867 (N_14867,N_8979,N_7188);
nor U14868 (N_14868,N_8986,N_5229);
nor U14869 (N_14869,N_6603,N_7493);
nand U14870 (N_14870,N_8897,N_8235);
or U14871 (N_14871,N_9894,N_6579);
nand U14872 (N_14872,N_5647,N_8848);
nor U14873 (N_14873,N_5194,N_7545);
xnor U14874 (N_14874,N_9116,N_8378);
or U14875 (N_14875,N_9711,N_6481);
xor U14876 (N_14876,N_5147,N_7529);
nand U14877 (N_14877,N_5125,N_8619);
nor U14878 (N_14878,N_6388,N_9603);
or U14879 (N_14879,N_5968,N_8678);
nand U14880 (N_14880,N_7940,N_6898);
xnor U14881 (N_14881,N_9839,N_8445);
nor U14882 (N_14882,N_5099,N_9379);
nor U14883 (N_14883,N_8828,N_9478);
or U14884 (N_14884,N_5321,N_6716);
xor U14885 (N_14885,N_8500,N_9168);
nand U14886 (N_14886,N_8160,N_6985);
nand U14887 (N_14887,N_6632,N_8515);
and U14888 (N_14888,N_9281,N_8749);
and U14889 (N_14889,N_6933,N_7476);
xnor U14890 (N_14890,N_5655,N_8715);
or U14891 (N_14891,N_5036,N_5094);
and U14892 (N_14892,N_9880,N_9817);
xnor U14893 (N_14893,N_7908,N_6800);
and U14894 (N_14894,N_7280,N_9946);
xor U14895 (N_14895,N_5462,N_7412);
xnor U14896 (N_14896,N_8204,N_7920);
and U14897 (N_14897,N_7250,N_5442);
nor U14898 (N_14898,N_5943,N_9826);
and U14899 (N_14899,N_6576,N_7924);
xor U14900 (N_14900,N_6905,N_6117);
xnor U14901 (N_14901,N_6288,N_5178);
nor U14902 (N_14902,N_6558,N_6121);
or U14903 (N_14903,N_7791,N_7751);
xor U14904 (N_14904,N_7002,N_5823);
xnor U14905 (N_14905,N_9958,N_6626);
or U14906 (N_14906,N_7366,N_5727);
nor U14907 (N_14907,N_5969,N_6971);
nor U14908 (N_14908,N_9185,N_8062);
nor U14909 (N_14909,N_8231,N_5805);
and U14910 (N_14910,N_6015,N_5433);
xor U14911 (N_14911,N_6183,N_6280);
nor U14912 (N_14912,N_9548,N_7111);
nor U14913 (N_14913,N_9163,N_8561);
and U14914 (N_14914,N_7719,N_9738);
or U14915 (N_14915,N_6935,N_6274);
xnor U14916 (N_14916,N_8596,N_7388);
xor U14917 (N_14917,N_8433,N_7535);
nand U14918 (N_14918,N_5177,N_8394);
nor U14919 (N_14919,N_6413,N_6725);
nand U14920 (N_14920,N_8534,N_5132);
xnor U14921 (N_14921,N_9249,N_5008);
xor U14922 (N_14922,N_5430,N_7479);
nand U14923 (N_14923,N_9041,N_8310);
nor U14924 (N_14924,N_8883,N_7985);
and U14925 (N_14925,N_8033,N_9498);
xor U14926 (N_14926,N_7312,N_8772);
and U14927 (N_14927,N_8223,N_7770);
xor U14928 (N_14928,N_6281,N_8143);
nor U14929 (N_14929,N_8845,N_7163);
nor U14930 (N_14930,N_6158,N_8643);
nand U14931 (N_14931,N_8229,N_5048);
nor U14932 (N_14932,N_5382,N_7756);
or U14933 (N_14933,N_5313,N_8628);
xnor U14934 (N_14934,N_5506,N_9268);
and U14935 (N_14935,N_9868,N_9062);
or U14936 (N_14936,N_9857,N_9927);
or U14937 (N_14937,N_9342,N_7240);
and U14938 (N_14938,N_7083,N_8922);
xnor U14939 (N_14939,N_7600,N_6439);
xnor U14940 (N_14940,N_7524,N_6365);
or U14941 (N_14941,N_8653,N_9577);
xor U14942 (N_14942,N_8503,N_9728);
and U14943 (N_14943,N_9121,N_9180);
nor U14944 (N_14944,N_5720,N_5264);
nand U14945 (N_14945,N_5636,N_8572);
nand U14946 (N_14946,N_6452,N_7893);
or U14947 (N_14947,N_7576,N_7405);
nor U14948 (N_14948,N_9678,N_6412);
nand U14949 (N_14949,N_7207,N_7832);
nand U14950 (N_14950,N_8944,N_9794);
and U14951 (N_14951,N_9814,N_7806);
xnor U14952 (N_14952,N_8441,N_8446);
and U14953 (N_14953,N_9669,N_6974);
or U14954 (N_14954,N_9546,N_6717);
or U14955 (N_14955,N_8345,N_8989);
nor U14956 (N_14956,N_8713,N_8074);
or U14957 (N_14957,N_5318,N_6433);
or U14958 (N_14958,N_6917,N_9707);
xnor U14959 (N_14959,N_5667,N_6440);
and U14960 (N_14960,N_5594,N_8758);
nand U14961 (N_14961,N_8084,N_8199);
nand U14962 (N_14962,N_6481,N_6269);
xnor U14963 (N_14963,N_7049,N_5740);
and U14964 (N_14964,N_5384,N_5863);
and U14965 (N_14965,N_8835,N_6491);
or U14966 (N_14966,N_9297,N_7737);
nand U14967 (N_14967,N_5365,N_8299);
nor U14968 (N_14968,N_5195,N_9018);
and U14969 (N_14969,N_9552,N_9065);
and U14970 (N_14970,N_6530,N_9275);
xor U14971 (N_14971,N_9013,N_6311);
nand U14972 (N_14972,N_8472,N_6079);
and U14973 (N_14973,N_7354,N_7140);
and U14974 (N_14974,N_8567,N_6598);
nor U14975 (N_14975,N_6589,N_8227);
nand U14976 (N_14976,N_7782,N_6532);
and U14977 (N_14977,N_8677,N_5586);
nand U14978 (N_14978,N_7924,N_9471);
nor U14979 (N_14979,N_7042,N_5049);
and U14980 (N_14980,N_5695,N_5828);
nor U14981 (N_14981,N_9093,N_5499);
or U14982 (N_14982,N_9474,N_5802);
and U14983 (N_14983,N_9054,N_8330);
nand U14984 (N_14984,N_5169,N_7012);
xnor U14985 (N_14985,N_9174,N_8919);
or U14986 (N_14986,N_7571,N_7314);
xnor U14987 (N_14987,N_9505,N_6556);
nor U14988 (N_14988,N_7993,N_9930);
nor U14989 (N_14989,N_7504,N_6362);
nand U14990 (N_14990,N_6161,N_5984);
nand U14991 (N_14991,N_5007,N_6176);
xor U14992 (N_14992,N_6579,N_9458);
nand U14993 (N_14993,N_6048,N_7620);
nor U14994 (N_14994,N_7876,N_7936);
nor U14995 (N_14995,N_5994,N_6201);
nand U14996 (N_14996,N_5896,N_5949);
or U14997 (N_14997,N_9908,N_7868);
nand U14998 (N_14998,N_9733,N_9568);
nand U14999 (N_14999,N_7776,N_5132);
nor UO_0 (O_0,N_12964,N_11295);
and UO_1 (O_1,N_12070,N_12535);
xor UO_2 (O_2,N_13408,N_12954);
nand UO_3 (O_3,N_12199,N_13655);
and UO_4 (O_4,N_11500,N_12947);
and UO_5 (O_5,N_12529,N_13502);
nor UO_6 (O_6,N_14127,N_10804);
and UO_7 (O_7,N_13596,N_13218);
or UO_8 (O_8,N_13770,N_11967);
and UO_9 (O_9,N_12416,N_11702);
xnor UO_10 (O_10,N_10806,N_14339);
nor UO_11 (O_11,N_11568,N_11431);
and UO_12 (O_12,N_14940,N_14797);
nor UO_13 (O_13,N_12846,N_10367);
nand UO_14 (O_14,N_13099,N_14451);
and UO_15 (O_15,N_12566,N_13925);
and UO_16 (O_16,N_13063,N_14118);
nand UO_17 (O_17,N_12014,N_13721);
xnor UO_18 (O_18,N_14543,N_12662);
or UO_19 (O_19,N_14427,N_10583);
or UO_20 (O_20,N_13455,N_12700);
nor UO_21 (O_21,N_13600,N_12955);
nor UO_22 (O_22,N_11784,N_12029);
or UO_23 (O_23,N_13298,N_13639);
nand UO_24 (O_24,N_14328,N_13584);
xnor UO_25 (O_25,N_10356,N_12851);
xor UO_26 (O_26,N_12977,N_10377);
or UO_27 (O_27,N_12429,N_12194);
nor UO_28 (O_28,N_11403,N_10411);
or UO_29 (O_29,N_10038,N_14743);
nor UO_30 (O_30,N_14863,N_13301);
nor UO_31 (O_31,N_13884,N_10584);
or UO_32 (O_32,N_12334,N_12757);
nor UO_33 (O_33,N_12033,N_10253);
xnor UO_34 (O_34,N_14463,N_11007);
and UO_35 (O_35,N_13253,N_10887);
or UO_36 (O_36,N_13848,N_14270);
xnor UO_37 (O_37,N_11055,N_14216);
nand UO_38 (O_38,N_12316,N_14417);
nand UO_39 (O_39,N_12492,N_13146);
xor UO_40 (O_40,N_10258,N_14034);
nand UO_41 (O_41,N_11277,N_14258);
nor UO_42 (O_42,N_12143,N_10589);
nor UO_43 (O_43,N_11175,N_10421);
and UO_44 (O_44,N_12067,N_14063);
xnor UO_45 (O_45,N_12807,N_10381);
or UO_46 (O_46,N_13534,N_13254);
xnor UO_47 (O_47,N_10579,N_12369);
and UO_48 (O_48,N_10051,N_13193);
nand UO_49 (O_49,N_12078,N_10448);
xor UO_50 (O_50,N_14828,N_10594);
nand UO_51 (O_51,N_12630,N_13391);
xor UO_52 (O_52,N_14899,N_12465);
nand UO_53 (O_53,N_11700,N_12975);
nor UO_54 (O_54,N_13958,N_11670);
or UO_55 (O_55,N_13693,N_12017);
or UO_56 (O_56,N_13134,N_12799);
nand UO_57 (O_57,N_10209,N_14713);
nor UO_58 (O_58,N_13729,N_12277);
or UO_59 (O_59,N_12036,N_13519);
and UO_60 (O_60,N_11559,N_12288);
nand UO_61 (O_61,N_12755,N_13797);
and UO_62 (O_62,N_14016,N_11337);
or UO_63 (O_63,N_10453,N_10774);
and UO_64 (O_64,N_13978,N_13646);
or UO_65 (O_65,N_14554,N_14210);
and UO_66 (O_66,N_12681,N_11617);
nor UO_67 (O_67,N_13690,N_11313);
and UO_68 (O_68,N_13834,N_10093);
nand UO_69 (O_69,N_11254,N_10597);
nor UO_70 (O_70,N_10437,N_14742);
xor UO_71 (O_71,N_12372,N_13389);
xor UO_72 (O_72,N_14702,N_13730);
nand UO_73 (O_73,N_12306,N_12667);
and UO_74 (O_74,N_13742,N_12497);
nor UO_75 (O_75,N_10728,N_10376);
and UO_76 (O_76,N_10251,N_13713);
nand UO_77 (O_77,N_11163,N_14213);
xor UO_78 (O_78,N_12158,N_14791);
and UO_79 (O_79,N_10245,N_14286);
or UO_80 (O_80,N_14668,N_10516);
nor UO_81 (O_81,N_14059,N_11872);
nand UO_82 (O_82,N_14294,N_14586);
nand UO_83 (O_83,N_13987,N_11888);
nand UO_84 (O_84,N_11467,N_11488);
nand UO_85 (O_85,N_14235,N_13572);
nor UO_86 (O_86,N_11933,N_13044);
nand UO_87 (O_87,N_10927,N_12902);
nor UO_88 (O_88,N_13479,N_14255);
xnor UO_89 (O_89,N_12875,N_12574);
nor UO_90 (O_90,N_11035,N_14137);
xor UO_91 (O_91,N_13334,N_12329);
and UO_92 (O_92,N_14612,N_12778);
or UO_93 (O_93,N_11239,N_10212);
and UO_94 (O_94,N_14849,N_10297);
nand UO_95 (O_95,N_10656,N_12003);
xor UO_96 (O_96,N_11356,N_12819);
or UO_97 (O_97,N_11961,N_10125);
xor UO_98 (O_98,N_10240,N_12233);
xor UO_99 (O_99,N_12570,N_12146);
and UO_100 (O_100,N_11144,N_12990);
and UO_101 (O_101,N_10676,N_10724);
nor UO_102 (O_102,N_10200,N_12622);
or UO_103 (O_103,N_14448,N_10529);
or UO_104 (O_104,N_10341,N_11381);
xnor UO_105 (O_105,N_10807,N_11126);
nor UO_106 (O_106,N_11739,N_13811);
nand UO_107 (O_107,N_10073,N_11331);
or UO_108 (O_108,N_11519,N_11034);
nor UO_109 (O_109,N_11200,N_14266);
xnor UO_110 (O_110,N_12792,N_12589);
or UO_111 (O_111,N_14480,N_10213);
or UO_112 (O_112,N_11466,N_13297);
xnor UO_113 (O_113,N_14009,N_10990);
and UO_114 (O_114,N_12770,N_11544);
and UO_115 (O_115,N_10497,N_12654);
xnor UO_116 (O_116,N_11038,N_10737);
and UO_117 (O_117,N_14139,N_10829);
or UO_118 (O_118,N_11651,N_11526);
xnor UO_119 (O_119,N_11733,N_13920);
or UO_120 (O_120,N_11927,N_11300);
and UO_121 (O_121,N_14169,N_14674);
nand UO_122 (O_122,N_11432,N_14380);
or UO_123 (O_123,N_13355,N_13205);
nor UO_124 (O_124,N_13016,N_14881);
nor UO_125 (O_125,N_14880,N_10417);
or UO_126 (O_126,N_10171,N_11706);
xor UO_127 (O_127,N_12820,N_14798);
or UO_128 (O_128,N_12668,N_11977);
xnor UO_129 (O_129,N_10653,N_14116);
or UO_130 (O_130,N_12400,N_11713);
nand UO_131 (O_131,N_10886,N_12279);
or UO_132 (O_132,N_11899,N_12883);
or UO_133 (O_133,N_12172,N_10031);
nor UO_134 (O_134,N_14305,N_14188);
or UO_135 (O_135,N_14581,N_11222);
and UO_136 (O_136,N_10474,N_14708);
or UO_137 (O_137,N_10866,N_14144);
xnor UO_138 (O_138,N_11496,N_13335);
and UO_139 (O_139,N_14683,N_11723);
nand UO_140 (O_140,N_12319,N_12395);
or UO_141 (O_141,N_11025,N_12650);
and UO_142 (O_142,N_11252,N_13842);
xor UO_143 (O_143,N_11475,N_10204);
nor UO_144 (O_144,N_14942,N_11352);
and UO_145 (O_145,N_12076,N_14322);
or UO_146 (O_146,N_10285,N_10298);
nand UO_147 (O_147,N_12506,N_12950);
and UO_148 (O_148,N_10135,N_10063);
and UO_149 (O_149,N_14620,N_12080);
and UO_150 (O_150,N_12691,N_12679);
or UO_151 (O_151,N_12601,N_14453);
or UO_152 (O_152,N_11399,N_10416);
xnor UO_153 (O_153,N_10199,N_11894);
and UO_154 (O_154,N_12835,N_12243);
and UO_155 (O_155,N_13381,N_10752);
and UO_156 (O_156,N_10470,N_13496);
nand UO_157 (O_157,N_12494,N_12043);
nor UO_158 (O_158,N_10483,N_12002);
or UO_159 (O_159,N_14747,N_12422);
xnor UO_160 (O_160,N_13701,N_13943);
or UO_161 (O_161,N_11465,N_11584);
or UO_162 (O_162,N_11452,N_14660);
or UO_163 (O_163,N_12921,N_11645);
and UO_164 (O_164,N_12396,N_14512);
or UO_165 (O_165,N_13450,N_10596);
nand UO_166 (O_166,N_11718,N_12719);
nand UO_167 (O_167,N_13598,N_14547);
or UO_168 (O_168,N_13086,N_12849);
or UO_169 (O_169,N_14385,N_10352);
or UO_170 (O_170,N_10748,N_10238);
nand UO_171 (O_171,N_11778,N_10864);
nor UO_172 (O_172,N_14055,N_12345);
nand UO_173 (O_173,N_13832,N_14419);
nor UO_174 (O_174,N_11990,N_14654);
xnor UO_175 (O_175,N_10154,N_11549);
nor UO_176 (O_176,N_10754,N_13021);
and UO_177 (O_177,N_11834,N_13163);
nand UO_178 (O_178,N_10023,N_10469);
nor UO_179 (O_179,N_12845,N_11176);
nand UO_180 (O_180,N_12683,N_11677);
nor UO_181 (O_181,N_12123,N_10492);
nand UO_182 (O_182,N_14414,N_14723);
nor UO_183 (O_183,N_14399,N_10787);
nand UO_184 (O_184,N_13268,N_14580);
xnor UO_185 (O_185,N_11386,N_11540);
or UO_186 (O_186,N_10142,N_13169);
xor UO_187 (O_187,N_10185,N_12932);
nor UO_188 (O_188,N_12793,N_12058);
nor UO_189 (O_189,N_12042,N_14051);
xnor UO_190 (O_190,N_13932,N_14875);
or UO_191 (O_191,N_10932,N_13759);
xnor UO_192 (O_192,N_14376,N_13156);
xor UO_193 (O_193,N_11151,N_11181);
nor UO_194 (O_194,N_12737,N_10180);
nor UO_195 (O_195,N_12624,N_12263);
or UO_196 (O_196,N_11269,N_14653);
and UO_197 (O_197,N_13185,N_13845);
and UO_198 (O_198,N_13039,N_13919);
or UO_199 (O_199,N_10822,N_11213);
or UO_200 (O_200,N_10090,N_10161);
or UO_201 (O_201,N_12546,N_12915);
and UO_202 (O_202,N_12407,N_11976);
and UO_203 (O_203,N_12335,N_10471);
or UO_204 (O_204,N_12040,N_10153);
nor UO_205 (O_205,N_12717,N_13672);
and UO_206 (O_206,N_10973,N_10010);
and UO_207 (O_207,N_12696,N_13878);
or UO_208 (O_208,N_10928,N_13855);
nand UO_209 (O_209,N_12397,N_12694);
nor UO_210 (O_210,N_13524,N_11287);
and UO_211 (O_211,N_12145,N_11656);
and UO_212 (O_212,N_10184,N_13535);
xnor UO_213 (O_213,N_12004,N_10109);
nor UO_214 (O_214,N_10770,N_11384);
nor UO_215 (O_215,N_13509,N_13140);
or UO_216 (O_216,N_11204,N_12094);
xnor UO_217 (O_217,N_14768,N_12560);
nor UO_218 (O_218,N_11059,N_12294);
nand UO_219 (O_219,N_14181,N_12262);
xnor UO_220 (O_220,N_12897,N_14811);
nand UO_221 (O_221,N_11944,N_10160);
nor UO_222 (O_222,N_14582,N_10699);
nor UO_223 (O_223,N_13810,N_10466);
nor UO_224 (O_224,N_10922,N_11813);
or UO_225 (O_225,N_13242,N_14390);
xor UO_226 (O_226,N_13123,N_10612);
xor UO_227 (O_227,N_13325,N_14311);
nor UO_228 (O_228,N_11604,N_12657);
xnor UO_229 (O_229,N_10564,N_14633);
and UO_230 (O_230,N_13059,N_14796);
xor UO_231 (O_231,N_14238,N_10134);
nand UO_232 (O_232,N_14388,N_13684);
and UO_233 (O_233,N_14436,N_13981);
or UO_234 (O_234,N_10027,N_11971);
and UO_235 (O_235,N_13788,N_14622);
nand UO_236 (O_236,N_14966,N_11903);
or UO_237 (O_237,N_13424,N_14087);
nor UO_238 (O_238,N_14319,N_10781);
and UO_239 (O_239,N_12027,N_14550);
xor UO_240 (O_240,N_12871,N_14386);
and UO_241 (O_241,N_13631,N_13037);
and UO_242 (O_242,N_14918,N_10461);
nand UO_243 (O_243,N_10802,N_13966);
xnor UO_244 (O_244,N_12842,N_14840);
nand UO_245 (O_245,N_12870,N_13265);
nand UO_246 (O_246,N_13340,N_14284);
nand UO_247 (O_247,N_12477,N_11861);
nand UO_248 (O_248,N_12826,N_12249);
and UO_249 (O_249,N_12658,N_10302);
nor UO_250 (O_250,N_14870,N_10982);
or UO_251 (O_251,N_10828,N_11516);
nor UO_252 (O_252,N_12858,N_12399);
and UO_253 (O_253,N_13635,N_11491);
nor UO_254 (O_254,N_10116,N_12805);
xnor UO_255 (O_255,N_14326,N_13210);
nand UO_256 (O_256,N_12804,N_14409);
xor UO_257 (O_257,N_10995,N_13793);
and UO_258 (O_258,N_11004,N_10476);
or UO_259 (O_259,N_10370,N_14128);
xor UO_260 (O_260,N_14561,N_11566);
xor UO_261 (O_261,N_13963,N_11486);
nor UO_262 (O_262,N_13776,N_12054);
nand UO_263 (O_263,N_10966,N_12287);
and UO_264 (O_264,N_11551,N_13652);
xor UO_265 (O_265,N_14891,N_14135);
nand UO_266 (O_266,N_13587,N_11987);
xor UO_267 (O_267,N_12364,N_14021);
xor UO_268 (O_268,N_11804,N_14335);
nor UO_269 (O_269,N_13533,N_12255);
nor UO_270 (O_270,N_13187,N_14952);
xor UO_271 (O_271,N_14267,N_13720);
nor UO_272 (O_272,N_13907,N_10276);
and UO_273 (O_273,N_13594,N_11309);
or UO_274 (O_274,N_10835,N_10955);
xor UO_275 (O_275,N_11202,N_11818);
or UO_276 (O_276,N_10003,N_13518);
or UO_277 (O_277,N_12984,N_13816);
nor UO_278 (O_278,N_14770,N_10337);
nand UO_279 (O_279,N_11797,N_10956);
and UO_280 (O_280,N_10576,N_13277);
nor UO_281 (O_281,N_11093,N_14243);
and UO_282 (O_282,N_11740,N_10799);
and UO_283 (O_283,N_14005,N_14013);
nand UO_284 (O_284,N_13260,N_11595);
or UO_285 (O_285,N_12527,N_14161);
and UO_286 (O_286,N_11564,N_12142);
or UO_287 (O_287,N_13317,N_14902);
and UO_288 (O_288,N_10042,N_10017);
or UO_289 (O_289,N_13013,N_14956);
nand UO_290 (O_290,N_14734,N_13179);
nor UO_291 (O_291,N_14854,N_11900);
nor UO_292 (O_292,N_10499,N_12237);
or UO_293 (O_293,N_11117,N_10145);
nand UO_294 (O_294,N_14502,N_10801);
and UO_295 (O_295,N_11019,N_12026);
or UO_296 (O_296,N_13200,N_13227);
xnor UO_297 (O_297,N_14040,N_10895);
or UO_298 (O_298,N_13459,N_12159);
nor UO_299 (O_299,N_13551,N_12413);
xor UO_300 (O_300,N_11455,N_14520);
nand UO_301 (O_301,N_10338,N_13444);
or UO_302 (O_302,N_12852,N_10057);
nand UO_303 (O_303,N_10299,N_12920);
xor UO_304 (O_304,N_13611,N_13570);
nand UO_305 (O_305,N_13195,N_11964);
and UO_306 (O_306,N_13500,N_14108);
and UO_307 (O_307,N_12959,N_14705);
or UO_308 (O_308,N_13700,N_10128);
nand UO_309 (O_309,N_10293,N_14571);
and UO_310 (O_310,N_11327,N_14221);
xnor UO_311 (O_311,N_14605,N_14408);
or UO_312 (O_312,N_11103,N_11314);
and UO_313 (O_313,N_14469,N_14279);
or UO_314 (O_314,N_10190,N_13423);
and UO_315 (O_315,N_10143,N_14995);
xnor UO_316 (O_316,N_10552,N_11116);
xor UO_317 (O_317,N_10254,N_10625);
xnor UO_318 (O_318,N_11115,N_10713);
xor UO_319 (O_319,N_12165,N_11916);
and UO_320 (O_320,N_12854,N_10132);
and UO_321 (O_321,N_10919,N_13120);
and UO_322 (O_322,N_14292,N_14497);
nor UO_323 (O_323,N_13688,N_12953);
nor UO_324 (O_324,N_12367,N_13457);
and UO_325 (O_325,N_14324,N_14236);
nor UO_326 (O_326,N_14194,N_12878);
and UO_327 (O_327,N_12522,N_14814);
or UO_328 (O_328,N_14232,N_10503);
nand UO_329 (O_329,N_14538,N_13249);
or UO_330 (O_330,N_10182,N_14862);
xnor UO_331 (O_331,N_13817,N_14533);
xor UO_332 (O_332,N_10741,N_14984);
or UO_333 (O_333,N_10778,N_14084);
nor UO_334 (O_334,N_12602,N_12960);
nor UO_335 (O_335,N_11541,N_10062);
and UO_336 (O_336,N_13328,N_13419);
and UO_337 (O_337,N_13549,N_13209);
nor UO_338 (O_338,N_14699,N_13972);
nand UO_339 (O_339,N_10407,N_14320);
nor UO_340 (O_340,N_13960,N_10179);
and UO_341 (O_341,N_13141,N_14688);
and UO_342 (O_342,N_10217,N_13349);
or UO_343 (O_343,N_10599,N_14123);
nor UO_344 (O_344,N_12134,N_12130);
or UO_345 (O_345,N_13090,N_12711);
or UO_346 (O_346,N_10506,N_10414);
and UO_347 (O_347,N_12742,N_11279);
and UO_348 (O_348,N_13917,N_14015);
nor UO_349 (O_349,N_13677,N_14733);
and UO_350 (O_350,N_12347,N_13442);
xnor UO_351 (O_351,N_11823,N_10273);
or UO_352 (O_352,N_12115,N_11765);
nand UO_353 (O_353,N_10723,N_10015);
xor UO_354 (O_354,N_13875,N_11957);
or UO_355 (O_355,N_12350,N_10224);
or UO_356 (O_356,N_14962,N_11368);
nand UO_357 (O_357,N_11511,N_12796);
xnor UO_358 (O_358,N_10330,N_13213);
xnor UO_359 (O_359,N_12016,N_10991);
nand UO_360 (O_360,N_10423,N_12060);
or UO_361 (O_361,N_12880,N_12154);
nand UO_362 (O_362,N_14931,N_14429);
xor UO_363 (O_363,N_13903,N_13626);
and UO_364 (O_364,N_11935,N_12712);
xnor UO_365 (O_365,N_12768,N_10084);
xnor UO_366 (O_366,N_11679,N_11535);
nand UO_367 (O_367,N_12714,N_10277);
and UO_368 (O_368,N_10907,N_13112);
xor UO_369 (O_369,N_13220,N_14331);
or UO_370 (O_370,N_10156,N_14314);
nand UO_371 (O_371,N_14532,N_12197);
or UO_372 (O_372,N_10521,N_12850);
xnor UO_373 (O_373,N_13080,N_10127);
xor UO_374 (O_374,N_12252,N_12776);
xnor UO_375 (O_375,N_13353,N_14576);
xor UO_376 (O_376,N_13130,N_14100);
or UO_377 (O_377,N_13024,N_13826);
xor UO_378 (O_378,N_13405,N_11472);
xnor UO_379 (O_379,N_10112,N_13303);
nor UO_380 (O_380,N_14053,N_10518);
xnor UO_381 (O_381,N_14499,N_11746);
and UO_382 (O_382,N_13870,N_12232);
xor UO_383 (O_383,N_11842,N_14707);
and UO_384 (O_384,N_10219,N_13077);
or UO_385 (O_385,N_11460,N_12122);
or UO_386 (O_386,N_12353,N_13038);
xor UO_387 (O_387,N_12663,N_11264);
nand UO_388 (O_388,N_12087,N_12967);
nor UO_389 (O_389,N_12392,N_12615);
and UO_390 (O_390,N_11777,N_10721);
and UO_391 (O_391,N_11908,N_13497);
or UO_392 (O_392,N_10236,N_12519);
nand UO_393 (O_393,N_11658,N_10571);
xnor UO_394 (O_394,N_14035,N_13168);
or UO_395 (O_395,N_10261,N_14075);
nand UO_396 (O_396,N_14514,N_11879);
and UO_397 (O_397,N_14275,N_13930);
nor UO_398 (O_398,N_13223,N_10379);
nor UO_399 (O_399,N_14295,N_13098);
xor UO_400 (O_400,N_14046,N_12110);
and UO_401 (O_401,N_12983,N_10290);
nor UO_402 (O_402,N_12769,N_12376);
and UO_403 (O_403,N_13886,N_12448);
and UO_404 (O_404,N_12857,N_10681);
nand UO_405 (O_405,N_14458,N_13245);
nand UO_406 (O_406,N_12718,N_12750);
and UO_407 (O_407,N_14313,N_14352);
or UO_408 (O_408,N_14640,N_10440);
nand UO_409 (O_409,N_10647,N_13791);
and UO_410 (O_410,N_14510,N_11463);
and UO_411 (O_411,N_13913,N_12951);
xor UO_412 (O_412,N_10908,N_10567);
and UO_413 (O_413,N_12030,N_13618);
and UO_414 (O_414,N_13426,N_13456);
or UO_415 (O_415,N_10152,N_14321);
or UO_416 (O_416,N_10308,N_14407);
nand UO_417 (O_417,N_11958,N_10074);
nor UO_418 (O_418,N_13427,N_10332);
and UO_419 (O_419,N_10147,N_13786);
nor UO_420 (O_420,N_10668,N_12720);
nor UO_421 (O_421,N_12149,N_11644);
nor UO_422 (O_422,N_10641,N_13372);
nor UO_423 (O_423,N_12569,N_14093);
nand UO_424 (O_424,N_11965,N_13507);
nand UO_425 (O_425,N_11856,N_14047);
or UO_426 (O_426,N_11847,N_14579);
nand UO_427 (O_427,N_10747,N_14527);
nand UO_428 (O_428,N_10896,N_11322);
or UO_429 (O_429,N_13188,N_10030);
xnor UO_430 (O_430,N_12409,N_13715);
nor UO_431 (O_431,N_11930,N_12470);
or UO_432 (O_432,N_10755,N_14193);
and UO_433 (O_433,N_13243,N_10333);
and UO_434 (O_434,N_11884,N_12640);
xnor UO_435 (O_435,N_12341,N_13591);
nand UO_436 (O_436,N_12735,N_14518);
or UO_437 (O_437,N_14949,N_13679);
xor UO_438 (O_438,N_11245,N_13799);
xnor UO_439 (O_439,N_10222,N_13540);
nand UO_440 (O_440,N_13458,N_14774);
and UO_441 (O_441,N_13199,N_13064);
or UO_442 (O_442,N_13809,N_11119);
and UO_443 (O_443,N_14416,N_14631);
nand UO_444 (O_444,N_10201,N_14360);
xnor UO_445 (O_445,N_13109,N_10616);
nor UO_446 (O_446,N_11569,N_11415);
xor UO_447 (O_447,N_10316,N_10148);
nand UO_448 (O_448,N_14757,N_14245);
xor UO_449 (O_449,N_13663,N_13320);
nand UO_450 (O_450,N_13544,N_10005);
xor UO_451 (O_451,N_14070,N_12173);
nor UO_452 (O_452,N_10661,N_13009);
nand UO_453 (O_453,N_10060,N_10591);
nand UO_454 (O_454,N_10227,N_12840);
nand UO_455 (O_455,N_10208,N_13796);
or UO_456 (O_456,N_12082,N_14648);
xor UO_457 (O_457,N_12208,N_12664);
nor UO_458 (O_458,N_14739,N_14993);
or UO_459 (O_459,N_10763,N_11555);
xnor UO_460 (O_460,N_12862,N_11143);
nand UO_461 (O_461,N_10071,N_10646);
and UO_462 (O_462,N_10615,N_11859);
nor UO_463 (O_463,N_14603,N_11229);
or UO_464 (O_464,N_14761,N_13728);
or UO_465 (O_465,N_12402,N_11328);
nand UO_466 (O_466,N_10243,N_10834);
xor UO_467 (O_467,N_10702,N_13812);
xnor UO_468 (O_468,N_12317,N_10794);
xnor UO_469 (O_469,N_10412,N_13373);
or UO_470 (O_470,N_10020,N_12178);
nand UO_471 (O_471,N_12096,N_13154);
xor UO_472 (O_472,N_12424,N_12176);
and UO_473 (O_473,N_12503,N_12022);
xor UO_474 (O_474,N_13025,N_11835);
and UO_475 (O_475,N_11639,N_14866);
or UO_476 (O_476,N_10342,N_14342);
nor UO_477 (O_477,N_14056,N_12486);
and UO_478 (O_478,N_13856,N_14687);
or UO_479 (O_479,N_14735,N_11233);
xnor UO_480 (O_480,N_14293,N_13530);
and UO_481 (O_481,N_10235,N_13698);
and UO_482 (O_482,N_12642,N_13051);
nor UO_483 (O_483,N_14837,N_13173);
nor UO_484 (O_484,N_12726,N_10335);
xor UO_485 (O_485,N_11985,N_11866);
nor UO_486 (O_486,N_13703,N_14208);
xnor UO_487 (O_487,N_13725,N_10904);
and UO_488 (O_488,N_14104,N_11819);
nand UO_489 (O_489,N_13089,N_13377);
nor UO_490 (O_490,N_13621,N_13395);
nand UO_491 (O_491,N_14864,N_12135);
or UO_492 (O_492,N_14485,N_12710);
xor UO_493 (O_493,N_14254,N_12435);
nand UO_494 (O_494,N_13827,N_13364);
nand UO_495 (O_495,N_12291,N_12573);
and UO_496 (O_496,N_13062,N_12698);
or UO_497 (O_497,N_11572,N_11203);
nand UO_498 (O_498,N_13036,N_12517);
xnor UO_499 (O_499,N_14555,N_11024);
and UO_500 (O_500,N_13678,N_10013);
nor UO_501 (O_501,N_10124,N_11710);
and UO_502 (O_502,N_11824,N_10534);
nor UO_503 (O_503,N_14172,N_12659);
or UO_504 (O_504,N_14452,N_13017);
and UO_505 (O_505,N_10856,N_12905);
and UO_506 (O_506,N_11137,N_13144);
and UO_507 (O_507,N_13516,N_14782);
nor UO_508 (O_508,N_12542,N_12469);
and UO_509 (O_509,N_14099,N_10674);
and UO_510 (O_510,N_11928,N_11748);
or UO_511 (O_511,N_13740,N_10272);
nand UO_512 (O_512,N_12764,N_10710);
and UO_513 (O_513,N_13022,N_12481);
and UO_514 (O_514,N_14264,N_14560);
or UO_515 (O_515,N_11089,N_11148);
and UO_516 (O_516,N_13503,N_14378);
nand UO_517 (O_517,N_12295,N_10631);
nor UO_518 (O_518,N_10099,N_11557);
nor UO_519 (O_519,N_13177,N_10434);
nor UO_520 (O_520,N_10322,N_11329);
nand UO_521 (O_521,N_12919,N_14804);
and UO_522 (O_522,N_11422,N_14248);
nor UO_523 (O_523,N_13766,N_11406);
xor UO_524 (O_524,N_12012,N_14646);
and UO_525 (O_525,N_12612,N_11454);
nor UO_526 (O_526,N_11456,N_14164);
xnor UO_527 (O_527,N_10853,N_14886);
nand UO_528 (O_528,N_13401,N_13346);
nand UO_529 (O_529,N_12161,N_13939);
nor UO_530 (O_530,N_13476,N_12886);
xnor UO_531 (O_531,N_13654,N_10375);
and UO_532 (O_532,N_10089,N_10515);
or UO_533 (O_533,N_13211,N_12818);
nor UO_534 (O_534,N_10292,N_14979);
and UO_535 (O_535,N_11211,N_14600);
nand UO_536 (O_536,N_14111,N_13250);
or UO_537 (O_537,N_12013,N_10540);
or UO_538 (O_538,N_13440,N_13924);
nand UO_539 (O_539,N_11489,N_12625);
or UO_540 (O_540,N_13110,N_13961);
and UO_541 (O_541,N_10050,N_10851);
nand UO_542 (O_542,N_14746,N_14106);
nand UO_543 (O_543,N_14022,N_14839);
nor UO_544 (O_544,N_11377,N_11954);
nor UO_545 (O_545,N_11937,N_14685);
or UO_546 (O_546,N_11573,N_13904);
nand UO_547 (O_547,N_11194,N_13829);
nor UO_548 (O_548,N_11407,N_10274);
nand UO_549 (O_549,N_13840,N_14988);
xor UO_550 (O_550,N_13935,N_13998);
nor UO_551 (O_551,N_10178,N_11123);
nor UO_552 (O_552,N_10790,N_14630);
nand UO_553 (O_553,N_10939,N_13851);
and UO_554 (O_554,N_10961,N_11696);
or UO_555 (O_555,N_14191,N_10789);
nand UO_556 (O_556,N_12911,N_12695);
or UO_557 (O_557,N_11947,N_10924);
nand UO_558 (O_558,N_11110,N_11798);
nor UO_559 (O_559,N_11864,N_14537);
xnor UO_560 (O_560,N_12235,N_12245);
nor UO_561 (O_561,N_11762,N_12586);
nor UO_562 (O_562,N_14549,N_11811);
or UO_563 (O_563,N_12355,N_13993);
nor UO_564 (O_564,N_14365,N_12075);
xnor UO_565 (O_565,N_10662,N_14392);
nand UO_566 (O_566,N_13367,N_14044);
and UO_567 (O_567,N_12261,N_10347);
xnor UO_568 (O_568,N_11354,N_13893);
nor UO_569 (O_569,N_12998,N_10810);
nor UO_570 (O_570,N_14397,N_14917);
xor UO_571 (O_571,N_12128,N_13314);
and UO_572 (O_572,N_10749,N_14825);
nor UO_573 (O_573,N_14626,N_12461);
and UO_574 (O_574,N_11707,N_12937);
or UO_575 (O_575,N_10523,N_14615);
and UO_576 (O_576,N_11450,N_13955);
or UO_577 (O_577,N_13042,N_12285);
or UO_578 (O_578,N_13485,N_12127);
and UO_579 (O_579,N_11652,N_14426);
or UO_580 (O_580,N_11298,N_11855);
nor UO_581 (O_581,N_14991,N_10210);
xor UO_582 (O_582,N_14278,N_12073);
and UO_583 (O_583,N_13398,N_11830);
nand UO_584 (O_584,N_11493,N_11131);
xnor UO_585 (O_585,N_10507,N_14986);
and UO_586 (O_586,N_11111,N_13096);
nor UO_587 (O_587,N_13833,N_13581);
and UO_588 (O_588,N_11766,N_11220);
and UO_589 (O_589,N_10351,N_12203);
and UO_590 (O_590,N_11974,N_12485);
xnor UO_591 (O_591,N_10603,N_13436);
or UO_592 (O_592,N_11728,N_13716);
xnor UO_593 (O_593,N_12311,N_11552);
and UO_594 (O_594,N_10400,N_14004);
or UO_595 (O_595,N_10280,N_10729);
or UO_596 (O_596,N_10771,N_12383);
or UO_597 (O_597,N_10783,N_12147);
or UO_598 (O_598,N_11036,N_11484);
xor UO_599 (O_599,N_13289,N_12798);
or UO_600 (O_600,N_11880,N_10938);
and UO_601 (O_601,N_14091,N_11938);
and UO_602 (O_602,N_14969,N_12510);
and UO_603 (O_603,N_13839,N_13131);
and UO_604 (O_604,N_14186,N_12848);
nand UO_605 (O_605,N_11416,N_14412);
nor UO_606 (O_606,N_13049,N_11217);
or UO_607 (O_607,N_12860,N_11387);
nor UO_608 (O_608,N_13157,N_14487);
nand UO_609 (O_609,N_13074,N_14948);
xor UO_610 (O_610,N_13874,N_14277);
nor UO_611 (O_611,N_11192,N_14291);
nand UO_612 (O_612,N_11359,N_11168);
or UO_613 (O_613,N_13915,N_10353);
xnor UO_614 (O_614,N_13814,N_11380);
nand UO_615 (O_615,N_10248,N_11438);
or UO_616 (O_616,N_14629,N_12767);
and UO_617 (O_617,N_10942,N_13569);
and UO_618 (O_618,N_12466,N_10092);
and UO_619 (O_619,N_14251,N_13309);
and UO_620 (O_620,N_10988,N_12653);
nor UO_621 (O_621,N_12031,N_10220);
nand UO_622 (O_622,N_14649,N_10891);
or UO_623 (O_623,N_14884,N_10879);
nand UO_624 (O_624,N_13916,N_13868);
nor UO_625 (O_625,N_11737,N_11694);
nor UO_626 (O_626,N_12066,N_14489);
or UO_627 (O_627,N_10241,N_11468);
xor UO_628 (O_628,N_12867,N_14425);
nand UO_629 (O_629,N_10767,N_12783);
and UO_630 (O_630,N_10820,N_13333);
or UO_631 (O_631,N_14239,N_10174);
xor UO_632 (O_632,N_12912,N_10700);
nor UO_633 (O_633,N_14588,N_11097);
and UO_634 (O_634,N_12270,N_10717);
or UO_635 (O_635,N_11771,N_13033);
or UO_636 (O_636,N_10573,N_12206);
or UO_637 (O_637,N_11242,N_12336);
nor UO_638 (O_638,N_10989,N_12274);
xor UO_639 (O_639,N_14204,N_13722);
nor UO_640 (O_640,N_13241,N_11120);
nand UO_641 (O_641,N_13318,N_10494);
nor UO_642 (O_642,N_11166,N_14060);
nor UO_643 (O_643,N_12427,N_14975);
and UO_644 (O_644,N_13836,N_14006);
nand UO_645 (O_645,N_13505,N_10812);
xnor UO_646 (O_646,N_12062,N_10336);
nor UO_647 (O_647,N_10486,N_11371);
nand UO_648 (O_648,N_14066,N_11079);
xor UO_649 (O_649,N_13757,N_13975);
nor UO_650 (O_650,N_14889,N_10561);
nand UO_651 (O_651,N_14477,N_11132);
and UO_652 (O_652,N_10346,N_12202);
and UO_653 (O_653,N_10855,N_11324);
xnor UO_654 (O_654,N_10727,N_10905);
xor UO_655 (O_655,N_11689,N_13433);
nand UO_656 (O_656,N_14350,N_10357);
nand UO_657 (O_657,N_14460,N_10309);
xnor UO_658 (O_658,N_12739,N_13206);
or UO_659 (O_659,N_11446,N_14464);
and UO_660 (O_660,N_10159,N_13711);
and UO_661 (O_661,N_12224,N_12215);
xnor UO_662 (O_662,N_12312,N_10659);
and UO_663 (O_663,N_12479,N_13030);
and UO_664 (O_664,N_10649,N_13630);
nand UO_665 (O_665,N_14544,N_12432);
nand UO_666 (O_666,N_10041,N_13452);
nor UO_667 (O_667,N_12447,N_13180);
nand UO_668 (O_668,N_10488,N_11571);
xnor UO_669 (O_669,N_12117,N_10570);
nor UO_670 (O_670,N_11430,N_11505);
and UO_671 (O_671,N_11726,N_14001);
xnor UO_672 (O_672,N_10860,N_11357);
nand UO_673 (O_673,N_10260,N_10172);
or UO_674 (O_674,N_10198,N_12637);
or UO_675 (O_675,N_11753,N_13599);
or UO_676 (O_676,N_11518,N_13539);
or UO_677 (O_677,N_14769,N_11634);
or UO_678 (O_678,N_14298,N_13097);
or UO_679 (O_679,N_14945,N_10595);
or UO_680 (O_680,N_12756,N_12868);
or UO_681 (O_681,N_14574,N_10635);
or UO_682 (O_682,N_12204,N_11921);
and UO_683 (O_683,N_13813,N_14026);
or UO_684 (O_684,N_11863,N_10165);
or UO_685 (O_685,N_11917,N_13480);
and UO_686 (O_686,N_11072,N_11436);
and UO_687 (O_687,N_13750,N_12238);
and UO_688 (O_688,N_13495,N_12974);
and UO_689 (O_689,N_13523,N_10326);
xnor UO_690 (O_690,N_11993,N_11624);
nor UO_691 (O_691,N_11822,N_11304);
xor UO_692 (O_692,N_14632,N_10923);
or UO_693 (O_693,N_14736,N_11752);
and UO_694 (O_694,N_13947,N_10279);
nor UO_695 (O_695,N_14812,N_13733);
and UO_696 (O_696,N_12041,N_11315);
xnor UO_697 (O_697,N_13807,N_13625);
nor UO_698 (O_698,N_13506,N_14228);
nand UO_699 (O_699,N_10738,N_12419);
nor UO_700 (O_700,N_12386,N_11712);
nor UO_701 (O_701,N_12061,N_12425);
nor UO_702 (O_702,N_14050,N_11228);
or UO_703 (O_703,N_13737,N_10575);
or UO_704 (O_704,N_10740,N_12313);
or UO_705 (O_705,N_13215,N_14096);
nor UO_706 (O_706,N_10898,N_14503);
nor UO_707 (O_707,N_14637,N_14928);
and UO_708 (O_708,N_14765,N_11758);
xnor UO_709 (O_709,N_10123,N_11469);
nor UO_710 (O_710,N_10824,N_11683);
or UO_711 (O_711,N_14618,N_13453);
nor UO_712 (O_712,N_10175,N_10313);
nand UO_713 (O_713,N_12039,N_10839);
nand UO_714 (O_714,N_13831,N_13667);
or UO_715 (O_715,N_10994,N_13449);
nand UO_716 (O_716,N_11716,N_11068);
nand UO_717 (O_717,N_12266,N_10536);
or UO_718 (O_718,N_14616,N_10053);
xnor UO_719 (O_719,N_13018,N_11391);
nor UO_720 (O_720,N_11597,N_13057);
nor UO_721 (O_721,N_10630,N_13984);
or UO_722 (O_722,N_11109,N_13137);
nand UO_723 (O_723,N_12610,N_14391);
or UO_724 (O_724,N_11409,N_10232);
nand UO_725 (O_725,N_10399,N_11626);
xor UO_726 (O_726,N_10882,N_11458);
or UO_727 (O_727,N_11182,N_14474);
or UO_728 (O_728,N_11630,N_14696);
or UO_729 (O_729,N_10832,N_11730);
and UO_730 (O_730,N_11543,N_13352);
or UO_731 (O_731,N_10121,N_11895);
xnor UO_732 (O_732,N_13956,N_12889);
xnor UO_733 (O_733,N_14517,N_10859);
nor UO_734 (O_734,N_10444,N_10024);
nand UO_735 (O_735,N_10054,N_12946);
and UO_736 (O_736,N_13985,N_12504);
or UO_737 (O_737,N_12009,N_14909);
xor UO_738 (O_738,N_11461,N_12354);
nor UO_739 (O_739,N_14359,N_14115);
nand UO_740 (O_740,N_11026,N_11305);
and UO_741 (O_741,N_13803,N_10374);
and UO_742 (O_742,N_13538,N_10691);
or UO_743 (O_743,N_12103,N_12189);
or UO_744 (O_744,N_14418,N_12548);
and UO_745 (O_745,N_12749,N_14751);
xnor UO_746 (O_746,N_13000,N_13411);
and UO_747 (O_747,N_14383,N_10872);
and UO_748 (O_748,N_14714,N_12704);
or UO_749 (O_749,N_10598,N_12728);
and UO_750 (O_750,N_10590,N_11299);
or UO_751 (O_751,N_12556,N_10250);
or UO_752 (O_752,N_14658,N_10113);
and UO_753 (O_753,N_14865,N_11383);
nor UO_754 (O_754,N_10294,N_10618);
and UO_755 (O_755,N_12938,N_12956);
nor UO_756 (O_756,N_11638,N_14572);
nor UO_757 (O_757,N_12549,N_11705);
nor UO_758 (O_758,N_13577,N_14887);
and UO_759 (O_759,N_13446,N_11339);
and UO_760 (O_760,N_13365,N_10795);
nand UO_761 (O_761,N_10344,N_12001);
and UO_762 (O_762,N_12644,N_11561);
or UO_763 (O_763,N_12543,N_10965);
xnor UO_764 (O_764,N_10163,N_14915);
nand UO_765 (O_765,N_12411,N_11016);
nand UO_766 (O_766,N_10544,N_12195);
nor UO_767 (O_767,N_14130,N_11814);
nor UO_768 (O_768,N_12550,N_14645);
nor UO_769 (O_769,N_11043,N_14895);
and UO_770 (O_770,N_14030,N_10070);
xnor UO_771 (O_771,N_13121,N_10753);
xnor UO_772 (O_772,N_10672,N_12822);
nand UO_773 (O_773,N_13094,N_14478);
nand UO_774 (O_774,N_13777,N_11069);
nand UO_775 (O_775,N_14069,N_11852);
xnor UO_776 (O_776,N_11527,N_10869);
or UO_777 (O_777,N_10650,N_10100);
and UO_778 (O_778,N_13148,N_13670);
or UO_779 (O_779,N_13158,N_11171);
and UO_780 (O_780,N_12148,N_12370);
or UO_781 (O_781,N_10601,N_11514);
and UO_782 (O_782,N_11581,N_13704);
and UO_783 (O_783,N_14530,N_10894);
nor UO_784 (O_784,N_10917,N_10348);
nand UO_785 (O_785,N_12157,N_14604);
nand UO_786 (O_786,N_12280,N_10751);
nand UO_787 (O_787,N_14848,N_12217);
xnor UO_788 (O_788,N_12049,N_14597);
or UO_789 (O_789,N_11187,N_11362);
nor UO_790 (O_790,N_13264,N_11769);
nor UO_791 (O_791,N_14844,N_13633);
xnor UO_792 (O_792,N_13448,N_14608);
and UO_793 (O_793,N_14719,N_13393);
or UO_794 (O_794,N_12356,N_11152);
or UO_795 (O_795,N_13251,N_14017);
nor UO_796 (O_796,N_10509,N_11952);
and UO_797 (O_797,N_13366,N_11760);
nor UO_798 (O_798,N_14166,N_13143);
xnor UO_799 (O_799,N_14934,N_11084);
or UO_800 (O_800,N_13020,N_13432);
xor UO_801 (O_801,N_13270,N_14725);
or UO_802 (O_802,N_13321,N_10757);
nand UO_803 (O_803,N_11174,N_11922);
and UO_804 (O_804,N_10983,N_10874);
or UO_805 (O_805,N_12426,N_13830);
xor UO_806 (O_806,N_12365,N_14421);
xnor UO_807 (O_807,N_12192,N_10122);
and UO_808 (O_808,N_11998,N_13537);
xnor UO_809 (O_809,N_14566,N_13034);
and UO_810 (O_810,N_10743,N_14290);
xnor UO_811 (O_811,N_10047,N_13370);
or UO_812 (O_812,N_12784,N_10837);
xor UO_813 (O_813,N_14958,N_13382);
or UO_814 (O_814,N_11201,N_12387);
or UO_815 (O_815,N_10664,N_14472);
and UO_816 (O_816,N_10340,N_10543);
xnor UO_817 (O_817,N_10501,N_13542);
nor UO_818 (O_818,N_14795,N_14444);
or UO_819 (O_819,N_11153,N_12884);
xnor UO_820 (O_820,N_11991,N_11234);
xor UO_821 (O_821,N_11881,N_13047);
nand UO_822 (O_822,N_10909,N_13779);
or UO_823 (O_823,N_11378,N_12816);
xnor UO_824 (O_824,N_12682,N_12655);
xor UO_825 (O_825,N_11161,N_13573);
or UO_826 (O_826,N_11812,N_11749);
nor UO_827 (O_827,N_10697,N_10442);
nor UO_828 (O_828,N_11601,N_13441);
xnor UO_829 (O_829,N_10186,N_14819);
and UO_830 (O_830,N_13403,N_10526);
nand UO_831 (O_831,N_11846,N_10884);
and UO_832 (O_832,N_10401,N_12772);
nor UO_833 (O_833,N_14307,N_13853);
nor UO_834 (O_834,N_14901,N_12824);
nand UO_835 (O_835,N_13601,N_10247);
and UO_836 (O_836,N_14095,N_12450);
or UO_837 (O_837,N_11057,N_13100);
and UO_838 (O_838,N_11833,N_10857);
nor UO_839 (O_839,N_13843,N_11911);
and UO_840 (O_840,N_14872,N_13237);
nor UO_841 (O_841,N_13061,N_13460);
and UO_842 (O_842,N_12209,N_13085);
and UO_843 (O_843,N_12524,N_11787);
nor UO_844 (O_844,N_14994,N_12460);
xnor UO_845 (O_845,N_13876,N_10780);
and UO_846 (O_846,N_14253,N_12371);
xor UO_847 (O_847,N_13790,N_13986);
and UO_848 (O_848,N_10900,N_12308);
xnor UO_849 (O_849,N_10666,N_10314);
xor UO_850 (O_850,N_13015,N_12724);
or UO_851 (O_851,N_11311,N_12310);
nor UO_852 (O_852,N_10520,N_13221);
nor UO_853 (O_853,N_12170,N_11936);
or UO_854 (O_854,N_10962,N_13881);
nor UO_855 (O_855,N_11653,N_10363);
xor UO_856 (O_856,N_10067,N_12636);
nand UO_857 (O_857,N_11524,N_12180);
and UO_858 (O_858,N_13012,N_14920);
or UO_859 (O_859,N_14000,N_13617);
xor UO_860 (O_860,N_12575,N_11897);
nand UO_861 (O_861,N_14415,N_13478);
nand UO_862 (O_862,N_12412,N_14752);
and UO_863 (O_863,N_14717,N_12333);
xor UO_864 (O_864,N_13230,N_10513);
nand UO_865 (O_865,N_14085,N_14783);
nor UO_866 (O_866,N_12989,N_13789);
or UO_867 (O_867,N_14595,N_13233);
and UO_868 (O_868,N_13326,N_10768);
and UO_869 (O_869,N_14155,N_11816);
xnor UO_870 (O_870,N_14771,N_12090);
nor UO_871 (O_871,N_12939,N_12686);
and UO_872 (O_872,N_11780,N_11404);
xnor UO_873 (O_873,N_11681,N_14850);
nand UO_874 (O_874,N_10383,N_11792);
nor UO_875 (O_875,N_11248,N_14082);
nor UO_876 (O_876,N_10282,N_13226);
and UO_877 (O_877,N_12190,N_11104);
nand UO_878 (O_878,N_14202,N_12689);
xnor UO_879 (O_879,N_14457,N_10141);
or UO_880 (O_880,N_13708,N_12496);
xnor UO_881 (O_881,N_14806,N_14967);
xnor UO_882 (O_882,N_14471,N_12604);
nor UO_883 (O_883,N_10675,N_11860);
nor UO_884 (O_884,N_14535,N_12366);
nand UO_885 (O_885,N_12018,N_14265);
xnor UO_886 (O_886,N_12008,N_14856);
and UO_887 (O_887,N_14233,N_14430);
nor UO_888 (O_888,N_10081,N_12785);
nor UO_889 (O_889,N_13681,N_10192);
nand UO_890 (O_890,N_11266,N_12286);
nand UO_891 (O_891,N_13648,N_14465);
nor UO_892 (O_892,N_11218,N_11487);
nand UO_893 (O_893,N_11809,N_11688);
and UO_894 (O_894,N_11926,N_13905);
and UO_895 (O_895,N_11189,N_11969);
nand UO_896 (O_896,N_12813,N_12808);
nand UO_897 (O_897,N_10360,N_14585);
and UO_898 (O_898,N_10007,N_14109);
xor UO_899 (O_899,N_11241,N_12817);
nand UO_900 (O_900,N_14634,N_11732);
or UO_901 (O_901,N_13609,N_10438);
xor UO_902 (O_902,N_14627,N_14996);
xnor UO_903 (O_903,N_11291,N_12388);
nor UO_904 (O_904,N_12513,N_11960);
and UO_905 (O_905,N_10478,N_11546);
nand UO_906 (O_906,N_11857,N_14110);
nand UO_907 (O_907,N_12229,N_11946);
and UO_908 (O_908,N_12774,N_13723);
and UO_909 (O_909,N_13970,N_13582);
and UO_910 (O_910,N_11224,N_13272);
and UO_911 (O_911,N_14759,N_10968);
nand UO_912 (O_912,N_14377,N_11310);
nor UO_913 (O_913,N_13239,N_10663);
nand UO_914 (O_914,N_11006,N_11212);
nand UO_915 (O_915,N_12374,N_14141);
nand UO_916 (O_916,N_11389,N_10016);
nand UO_917 (O_917,N_13406,N_10237);
xor UO_918 (O_918,N_14014,N_10511);
nor UO_919 (O_919,N_12417,N_11457);
and UO_920 (O_920,N_10422,N_11350);
and UO_921 (O_921,N_13499,N_10604);
and UO_922 (O_922,N_14932,N_13971);
and UO_923 (O_923,N_14296,N_13528);
and UO_924 (O_924,N_12071,N_14479);
nand UO_925 (O_925,N_11288,N_11610);
xor UO_926 (O_926,N_14215,N_10731);
nand UO_927 (O_927,N_10532,N_12458);
nand UO_928 (O_928,N_14755,N_11263);
nor UO_929 (O_929,N_12271,N_11196);
nand UO_930 (O_930,N_12538,N_12568);
or UO_931 (O_931,N_10088,N_12023);
and UO_932 (O_932,N_14067,N_11210);
nand UO_933 (O_933,N_14564,N_11756);
and UO_934 (O_934,N_11776,N_10979);
nor UO_935 (O_935,N_10648,N_11542);
nand UO_936 (O_936,N_10960,N_10069);
nand UO_937 (O_937,N_11968,N_12941);
or UO_938 (O_938,N_13999,N_11221);
nor UO_939 (O_939,N_10993,N_14212);
or UO_940 (O_940,N_14484,N_10189);
nand UO_941 (O_941,N_14033,N_12678);
nor UO_942 (O_942,N_11708,N_13280);
nor UO_943 (O_943,N_12995,N_12649);
nor UO_944 (O_944,N_13197,N_12899);
xor UO_945 (O_945,N_13712,N_10371);
nor UO_946 (O_946,N_11138,N_11061);
nand UO_947 (O_947,N_14504,N_14261);
nand UO_948 (O_948,N_12182,N_10937);
nand UO_949 (O_949,N_14841,N_14832);
nand UO_950 (O_950,N_13647,N_13060);
nand UO_951 (O_951,N_12948,N_14794);
nor UO_952 (O_952,N_10164,N_13011);
xnor UO_953 (O_953,N_11494,N_14972);
or UO_954 (O_954,N_14269,N_12120);
xor UO_955 (O_955,N_14488,N_10542);
nor UO_956 (O_956,N_10975,N_14018);
xnor UO_957 (O_957,N_13738,N_14963);
xnor UO_958 (O_958,N_13238,N_14861);
nor UO_959 (O_959,N_10918,N_11147);
nand UO_960 (O_960,N_13741,N_10068);
or UO_961 (O_961,N_12131,N_14635);
nor UO_962 (O_962,N_10695,N_12021);
xnor UO_963 (O_963,N_13936,N_11827);
nand UO_964 (O_964,N_12766,N_14432);
nand UO_965 (O_965,N_11445,N_11021);
and UO_966 (O_966,N_10193,N_12254);
and UO_967 (O_967,N_13668,N_12155);
nand UO_968 (O_968,N_12439,N_11825);
or UO_969 (O_969,N_11433,N_11464);
or UO_970 (O_970,N_12379,N_11578);
and UO_971 (O_971,N_14358,N_12588);
nor UO_972 (O_972,N_13472,N_11000);
nor UO_973 (O_973,N_12898,N_12102);
or UO_974 (O_974,N_12598,N_10772);
xor UO_975 (O_975,N_14450,N_13486);
nor UO_976 (O_976,N_12708,N_14048);
or UO_977 (O_977,N_14237,N_14925);
nor UO_978 (O_978,N_10581,N_12906);
nor UO_979 (O_979,N_11408,N_14760);
nand UO_980 (O_980,N_12732,N_14944);
nand UO_981 (O_981,N_12153,N_14423);
nor UO_982 (O_982,N_13858,N_11376);
nand UO_983 (O_983,N_14929,N_11125);
xor UO_984 (O_984,N_10096,N_14156);
nor UO_985 (O_985,N_11301,N_12765);
xnor UO_986 (O_986,N_12759,N_11280);
nor UO_987 (O_987,N_11041,N_10528);
nand UO_988 (O_988,N_13043,N_10462);
xnor UO_989 (O_989,N_13965,N_14189);
and UO_990 (O_990,N_14766,N_11142);
nand UO_991 (O_991,N_14730,N_11956);
xor UO_992 (O_992,N_14521,N_10670);
or UO_993 (O_993,N_13494,N_10380);
or UO_994 (O_994,N_10097,N_13604);
or UO_995 (O_995,N_14131,N_14602);
xor UO_996 (O_996,N_11858,N_14971);
or UO_997 (O_997,N_12876,N_11247);
and UO_998 (O_998,N_12580,N_13135);
or UO_999 (O_999,N_11091,N_11849);
or UO_1000 (O_1000,N_12997,N_13806);
nor UO_1001 (O_1001,N_10914,N_12323);
xor UO_1002 (O_1002,N_12843,N_12741);
nor UO_1003 (O_1003,N_10562,N_11039);
nor UO_1004 (O_1004,N_11790,N_14955);
nor UO_1005 (O_1005,N_12385,N_14662);
nor UO_1006 (O_1006,N_14244,N_12595);
xor UO_1007 (O_1007,N_10249,N_14793);
nand UO_1008 (O_1008,N_11731,N_13360);
nand UO_1009 (O_1009,N_11530,N_13412);
xor UO_1010 (O_1010,N_10390,N_11801);
xor UO_1011 (O_1011,N_11599,N_13052);
or UO_1012 (O_1012,N_13232,N_14938);
nand UO_1013 (O_1013,N_10064,N_13988);
nor UO_1014 (O_1014,N_14973,N_13410);
nor UO_1015 (O_1015,N_14534,N_10759);
nor UO_1016 (O_1016,N_11483,N_11070);
and UO_1017 (O_1017,N_12895,N_11741);
xor UO_1018 (O_1018,N_12256,N_10101);
and UO_1019 (O_1019,N_14025,N_12687);
xnor UO_1020 (O_1020,N_11358,N_13661);
and UO_1021 (O_1021,N_11501,N_14097);
nand UO_1022 (O_1022,N_11556,N_12377);
xnor UO_1023 (O_1023,N_12452,N_14394);
and UO_1024 (O_1024,N_12674,N_14900);
nand UO_1025 (O_1025,N_14336,N_14710);
xor UO_1026 (O_1026,N_11660,N_14071);
nor UO_1027 (O_1027,N_14641,N_13212);
xor UO_1028 (O_1028,N_11770,N_14316);
xor UO_1029 (O_1029,N_10539,N_13383);
xnor UO_1030 (O_1030,N_13808,N_13161);
or UO_1031 (O_1031,N_12476,N_13040);
nor UO_1032 (O_1032,N_13536,N_11523);
nor UO_1033 (O_1033,N_10009,N_14644);
nand UO_1034 (O_1034,N_14598,N_11851);
nor UO_1035 (O_1035,N_11478,N_12339);
and UO_1036 (O_1036,N_10610,N_12923);
and UO_1037 (O_1037,N_12827,N_12320);
xor UO_1038 (O_1038,N_12576,N_11918);
and UO_1039 (O_1039,N_12791,N_10733);
or UO_1040 (O_1040,N_13997,N_13322);
nor UO_1041 (O_1041,N_13784,N_14345);
and UO_1042 (O_1042,N_14762,N_14138);
nand UO_1043 (O_1043,N_10014,N_12278);
nor UO_1044 (O_1044,N_14947,N_11796);
nand UO_1045 (O_1045,N_14306,N_14160);
nand UO_1046 (O_1046,N_14800,N_12487);
xor UO_1047 (O_1047,N_14851,N_13323);
nor UO_1048 (O_1048,N_10018,N_13643);
nand UO_1049 (O_1049,N_10557,N_11703);
or UO_1050 (O_1050,N_13153,N_11763);
or UO_1051 (O_1051,N_10456,N_14187);
xor UO_1052 (O_1052,N_14732,N_13804);
nand UO_1053 (O_1053,N_11934,N_10639);
and UO_1054 (O_1054,N_10485,N_11293);
xnor UO_1055 (O_1055,N_14673,N_10495);
and UO_1056 (O_1056,N_10847,N_12301);
and UO_1057 (O_1057,N_13775,N_12037);
nor UO_1058 (O_1058,N_10425,N_12318);
nand UO_1059 (O_1059,N_14843,N_14801);
nand UO_1060 (O_1060,N_14036,N_14098);
or UO_1061 (O_1061,N_11669,N_13104);
and UO_1062 (O_1062,N_14885,N_13136);
or UO_1063 (O_1063,N_14803,N_13707);
and UO_1064 (O_1064,N_10651,N_14404);
xor UO_1065 (O_1065,N_12651,N_12258);
nand UO_1066 (O_1066,N_13204,N_14957);
xnor UO_1067 (O_1067,N_12982,N_11018);
or UO_1068 (O_1068,N_14625,N_11845);
or UO_1069 (O_1069,N_10711,N_13562);
or UO_1070 (O_1070,N_14498,N_12092);
xor UO_1071 (O_1071,N_12281,N_10435);
or UO_1072 (O_1072,N_14455,N_13019);
or UO_1073 (O_1073,N_11725,N_10537);
xnor UO_1074 (O_1074,N_14821,N_12474);
nand UO_1075 (O_1075,N_13773,N_12495);
nor UO_1076 (O_1076,N_12338,N_14368);
xor UO_1077 (O_1077,N_12085,N_12561);
and UO_1078 (O_1078,N_11939,N_13548);
nor UO_1079 (O_1079,N_12596,N_10324);
nor UO_1080 (O_1080,N_11128,N_12641);
nand UO_1081 (O_1081,N_10021,N_10368);
or UO_1082 (O_1082,N_11915,N_10756);
nand UO_1083 (O_1083,N_12415,N_11611);
and UO_1084 (O_1084,N_10077,N_10555);
or UO_1085 (O_1085,N_14344,N_10373);
xor UO_1086 (O_1086,N_11914,N_10138);
and UO_1087 (O_1087,N_14587,N_14077);
xor UO_1088 (O_1088,N_13937,N_11788);
nor UO_1089 (O_1089,N_14496,N_14206);
nand UO_1090 (O_1090,N_10387,N_14838);
or UO_1091 (O_1091,N_10867,N_13361);
nand UO_1092 (O_1092,N_11548,N_11064);
or UO_1093 (O_1093,N_12944,N_11251);
or UO_1094 (O_1094,N_12554,N_11657);
or UO_1095 (O_1095,N_12661,N_14671);
xnor UO_1096 (O_1096,N_12518,N_14859);
and UO_1097 (O_1097,N_10343,N_13835);
nor UO_1098 (O_1098,N_12324,N_14575);
and UO_1099 (O_1099,N_13081,N_10176);
and UO_1100 (O_1100,N_12292,N_10079);
or UO_1101 (O_1101,N_10976,N_14570);
xor UO_1102 (O_1102,N_12855,N_11037);
or UO_1103 (O_1103,N_13922,N_12375);
nor UO_1104 (O_1104,N_10930,N_13088);
xnor UO_1105 (O_1105,N_14195,N_14285);
and UO_1106 (O_1106,N_11612,N_13614);
xor UO_1107 (O_1107,N_12966,N_14440);
or UO_1108 (O_1108,N_10196,N_13149);
and UO_1109 (O_1109,N_12251,N_14643);
nor UO_1110 (O_1110,N_13844,N_10677);
or UO_1111 (O_1111,N_10111,N_12931);
or UO_1112 (O_1112,N_13256,N_14964);
or UO_1113 (O_1113,N_13954,N_12760);
nand UO_1114 (O_1114,N_14287,N_12887);
nand UO_1115 (O_1115,N_14167,N_14756);
or UO_1116 (O_1116,N_11342,N_11547);
nand UO_1117 (O_1117,N_14052,N_11253);
xor UO_1118 (O_1118,N_14834,N_11983);
or UO_1119 (O_1119,N_12952,N_14476);
or UO_1120 (O_1120,N_14402,N_10981);
or UO_1121 (O_1121,N_10846,N_14650);
and UO_1122 (O_1122,N_10609,N_12024);
nor UO_1123 (O_1123,N_12825,N_10295);
nand UO_1124 (O_1124,N_13934,N_12337);
nor UO_1125 (O_1125,N_13687,N_10468);
nor UO_1126 (O_1126,N_12083,N_10311);
and UO_1127 (O_1127,N_13468,N_14628);
xor UO_1128 (O_1128,N_13852,N_13356);
xor UO_1129 (O_1129,N_12357,N_13114);
nor UO_1130 (O_1130,N_11402,N_12779);
xor UO_1131 (O_1131,N_14722,N_10687);
xor UO_1132 (O_1132,N_12198,N_12702);
or UO_1133 (O_1133,N_13866,N_12685);
and UO_1134 (O_1134,N_12248,N_10065);
and UO_1135 (O_1135,N_12652,N_14525);
nand UO_1136 (O_1136,N_13894,N_13525);
nor UO_1137 (O_1137,N_11032,N_12684);
nand UO_1138 (O_1138,N_11374,N_12482);
and UO_1139 (O_1139,N_14214,N_11179);
xor UO_1140 (O_1140,N_12098,N_11088);
nor UO_1141 (O_1141,N_11121,N_13510);
and UO_1142 (O_1142,N_11485,N_14374);
and UO_1143 (O_1143,N_10242,N_13683);
or UO_1144 (O_1144,N_12930,N_14513);
and UO_1145 (O_1145,N_10963,N_14669);
nor UO_1146 (O_1146,N_13491,N_14367);
nand UO_1147 (O_1147,N_11874,N_14105);
xor UO_1148 (O_1148,N_12446,N_12406);
or UO_1149 (O_1149,N_11410,N_13379);
and UO_1150 (O_1150,N_13122,N_13921);
and UO_1151 (O_1151,N_13557,N_13101);
nor UO_1152 (O_1152,N_10722,N_10818);
nand UO_1153 (O_1153,N_14524,N_14129);
and UO_1154 (O_1154,N_10758,N_12327);
and UO_1155 (O_1155,N_13498,N_12421);
nor UO_1156 (O_1156,N_13908,N_11366);
nand UO_1157 (O_1157,N_14983,N_12234);
nor UO_1158 (O_1158,N_13764,N_13801);
and UO_1159 (O_1159,N_12926,N_11896);
and UO_1160 (O_1160,N_11806,N_12483);
xnor UO_1161 (O_1161,N_10283,N_10082);
and UO_1162 (O_1162,N_12521,N_10739);
and UO_1163 (O_1163,N_12536,N_11648);
nor UO_1164 (O_1164,N_10890,N_14197);
and UO_1165 (O_1165,N_13392,N_12343);
nand UO_1166 (O_1166,N_12250,N_14492);
and UO_1167 (O_1167,N_10429,N_10139);
nand UO_1168 (O_1168,N_14327,N_10764);
and UO_1169 (O_1169,N_13224,N_11426);
and UO_1170 (O_1170,N_11363,N_10044);
and UO_1171 (O_1171,N_14434,N_11047);
nor UO_1172 (O_1172,N_11332,N_11022);
or UO_1173 (O_1173,N_13607,N_12267);
xnor UO_1174 (O_1174,N_13304,N_12803);
nor UO_1175 (O_1175,N_12428,N_11843);
or UO_1176 (O_1176,N_10246,N_13362);
nand UO_1177 (O_1177,N_13483,N_10278);
and UO_1178 (O_1178,N_11462,N_10964);
nor UO_1179 (O_1179,N_12782,N_13056);
and UO_1180 (O_1180,N_11099,N_13731);
xor UO_1181 (O_1181,N_14700,N_13589);
xor UO_1182 (O_1182,N_10393,N_10943);
or UO_1183 (O_1183,N_10858,N_14354);
nor UO_1184 (O_1184,N_10025,N_11294);
xor UO_1185 (O_1185,N_11704,N_14371);
or UO_1186 (O_1186,N_13475,N_13045);
xnor UO_1187 (O_1187,N_11885,N_11102);
xnor UO_1188 (O_1188,N_10593,N_10307);
or UO_1189 (O_1189,N_11420,N_10372);
nor UO_1190 (O_1190,N_11274,N_14283);
nand UO_1191 (O_1191,N_12314,N_10777);
and UO_1192 (O_1192,N_13912,N_10305);
and UO_1193 (O_1193,N_14028,N_13166);
nor UO_1194 (O_1194,N_14332,N_11130);
and UO_1195 (O_1195,N_13944,N_11992);
or UO_1196 (O_1196,N_13103,N_10266);
nor UO_1197 (O_1197,N_14090,N_13559);
or UO_1198 (O_1198,N_11640,N_13306);
nand UO_1199 (O_1199,N_13692,N_11275);
xnor UO_1200 (O_1200,N_13860,N_10239);
or UO_1201 (O_1201,N_13923,N_11347);
xor UO_1202 (O_1202,N_14882,N_12839);
or UO_1203 (O_1203,N_14508,N_12055);
and UO_1204 (O_1204,N_11870,N_11060);
or UO_1205 (O_1205,N_12063,N_13709);
and UO_1206 (O_1206,N_14406,N_13555);
xor UO_1207 (O_1207,N_13332,N_14807);
or UO_1208 (O_1208,N_10482,N_10133);
nand UO_1209 (O_1209,N_10323,N_10409);
xnor UO_1210 (O_1210,N_12979,N_12991);
nor UO_1211 (O_1211,N_11320,N_14974);
nor UO_1212 (O_1212,N_11439,N_10967);
or UO_1213 (O_1213,N_11642,N_10978);
nor UO_1214 (O_1214,N_13429,N_14744);
nor UO_1215 (O_1215,N_14970,N_12740);
xnor UO_1216 (O_1216,N_11209,N_14809);
and UO_1217 (O_1217,N_13190,N_13106);
and UO_1218 (O_1218,N_12112,N_13357);
and UO_1219 (O_1219,N_11943,N_11667);
or UO_1220 (O_1220,N_13138,N_12214);
nor UO_1221 (O_1221,N_14437,N_11165);
or UO_1222 (O_1222,N_11715,N_13841);
xor UO_1223 (O_1223,N_14062,N_12059);
or UO_1224 (O_1224,N_10833,N_10549);
nor UO_1225 (O_1225,N_12116,N_13567);
xor UO_1226 (O_1226,N_10958,N_12993);
or UO_1227 (O_1227,N_14968,N_11932);
xnor UO_1228 (O_1228,N_11051,N_13117);
nor UO_1229 (O_1229,N_12268,N_13588);
or UO_1230 (O_1230,N_11945,N_10572);
nand UO_1231 (O_1231,N_13070,N_10607);
nand UO_1232 (O_1232,N_12559,N_10527);
or UO_1233 (O_1233,N_11257,N_13324);
nand UO_1234 (O_1234,N_10765,N_12531);
and UO_1235 (O_1235,N_13949,N_10726);
and UO_1236 (O_1236,N_14246,N_11272);
or UO_1237 (O_1237,N_12330,N_12821);
or UO_1238 (O_1238,N_14552,N_13959);
nand UO_1239 (O_1239,N_13568,N_11563);
xnor UO_1240 (O_1240,N_13225,N_12885);
nor UO_1241 (O_1241,N_13780,N_12048);
nand UO_1242 (O_1242,N_12656,N_12414);
xnor UO_1243 (O_1243,N_10959,N_11244);
xor UO_1244 (O_1244,N_11775,N_11318);
xor UO_1245 (O_1245,N_12298,N_13164);
xnor UO_1246 (O_1246,N_14431,N_10032);
xnor UO_1247 (O_1247,N_11574,N_14847);
nand UO_1248 (O_1248,N_11498,N_14256);
or UO_1249 (O_1249,N_13753,N_12187);
xor UO_1250 (O_1250,N_13470,N_13443);
xnor UO_1251 (O_1251,N_13718,N_12787);
nor UO_1252 (O_1252,N_13911,N_11418);
or UO_1253 (O_1253,N_12220,N_14728);
and UO_1254 (O_1254,N_12913,N_11185);
xnor UO_1255 (O_1255,N_10947,N_11081);
and UO_1256 (O_1256,N_10850,N_13702);
or UO_1257 (O_1257,N_13992,N_13492);
and UO_1258 (O_1258,N_14589,N_10508);
nand UO_1259 (O_1259,N_10957,N_12015);
nand UO_1260 (O_1260,N_12551,N_11989);
nand UO_1261 (O_1261,N_14976,N_14401);
nand UO_1262 (O_1262,N_10550,N_12302);
nor UO_1263 (O_1263,N_10852,N_14698);
nor UO_1264 (O_1264,N_14505,N_13462);
nand UO_1265 (O_1265,N_14023,N_13007);
nor UO_1266 (O_1266,N_12581,N_14655);
and UO_1267 (O_1267,N_11902,N_13151);
nand UO_1268 (O_1268,N_13348,N_13805);
or UO_1269 (O_1269,N_14613,N_11193);
and UO_1270 (O_1270,N_12591,N_14177);
or UO_1271 (O_1271,N_11191,N_13758);
xor UO_1272 (O_1272,N_14081,N_14031);
and UO_1273 (O_1273,N_11575,N_14042);
xnor UO_1274 (O_1274,N_14817,N_10619);
xor UO_1275 (O_1275,N_13940,N_14540);
nor UO_1276 (O_1276,N_12404,N_11312);
xor UO_1277 (O_1277,N_14303,N_10998);
nand UO_1278 (O_1278,N_14583,N_10496);
or UO_1279 (O_1279,N_10854,N_10892);
nand UO_1280 (O_1280,N_12480,N_12627);
or UO_1281 (O_1281,N_13967,N_13128);
and UO_1282 (O_1282,N_12359,N_11424);
xor UO_1283 (O_1283,N_10873,N_12914);
or UO_1284 (O_1284,N_14370,N_13258);
nor UO_1285 (O_1285,N_11261,N_14482);
nand UO_1286 (O_1286,N_10705,N_13719);
nand UO_1287 (O_1287,N_11565,N_10150);
or UO_1288 (O_1288,N_11396,N_10329);
and UO_1289 (O_1289,N_11447,N_14682);
nand UO_1290 (O_1290,N_10463,N_13615);
xnor UO_1291 (O_1291,N_12828,N_14666);
or UO_1292 (O_1292,N_11742,N_14853);
and UO_1293 (O_1293,N_12006,N_13657);
xnor UO_1294 (O_1294,N_14200,N_14231);
nor UO_1295 (O_1295,N_11745,N_10136);
nand UO_1296 (O_1296,N_11105,N_10431);
and UO_1297 (O_1297,N_11227,N_14568);
or UO_1298 (O_1298,N_12869,N_11249);
nand UO_1299 (O_1299,N_10848,N_12265);
and UO_1300 (O_1300,N_14263,N_14490);
and UO_1301 (O_1301,N_14831,N_11836);
nand UO_1302 (O_1302,N_14545,N_11095);
nand UO_1303 (O_1303,N_12368,N_14086);
nand UO_1304 (O_1304,N_13263,N_10841);
and UO_1305 (O_1305,N_13186,N_12701);
nor UO_1306 (O_1306,N_13299,N_10578);
xnor UO_1307 (O_1307,N_13850,N_10952);
and UO_1308 (O_1308,N_12490,N_13724);
and UO_1309 (O_1309,N_14852,N_14729);
nor UO_1310 (O_1310,N_11628,N_14315);
nand UO_1311 (O_1311,N_11913,N_12978);
or UO_1312 (O_1312,N_13865,N_14609);
and UO_1313 (O_1313,N_11986,N_10933);
nor UO_1314 (O_1314,N_12669,N_11141);
xor UO_1315 (O_1315,N_11395,N_11664);
nand UO_1316 (O_1316,N_11577,N_10634);
and UO_1317 (O_1317,N_13115,N_13420);
xor UO_1318 (O_1318,N_12815,N_13347);
xnor UO_1319 (O_1319,N_11623,N_13522);
nor UO_1320 (O_1320,N_14462,N_12806);
nor UO_1321 (O_1321,N_13977,N_10586);
xnor UO_1322 (O_1322,N_12384,N_10689);
xnor UO_1323 (O_1323,N_10761,N_14822);
or UO_1324 (O_1324,N_10577,N_14773);
nand UO_1325 (O_1325,N_14509,N_13246);
or UO_1326 (O_1326,N_10257,N_12780);
nor UO_1327 (O_1327,N_12207,N_13028);
or UO_1328 (O_1328,N_12114,N_13583);
or UO_1329 (O_1329,N_11178,N_12363);
or UO_1330 (O_1330,N_14606,N_11782);
nor UO_1331 (O_1331,N_13649,N_13994);
nor UO_1332 (O_1332,N_10563,N_13563);
or UO_1333 (O_1333,N_10115,N_11815);
or UO_1334 (O_1334,N_10712,N_14262);
nand UO_1335 (O_1335,N_11255,N_12467);
xor UO_1336 (O_1336,N_11853,N_14684);
and UO_1337 (O_1337,N_11073,N_13255);
nand UO_1338 (O_1338,N_12936,N_13578);
nand UO_1339 (O_1339,N_10334,N_13973);
nor UO_1340 (O_1340,N_12462,N_14136);
and UO_1341 (O_1341,N_14002,N_12430);
or UO_1342 (O_1342,N_13545,N_10086);
nor UO_1343 (O_1343,N_14539,N_14679);
xnor UO_1344 (O_1344,N_10194,N_13527);
nand UO_1345 (O_1345,N_13402,N_13899);
and UO_1346 (O_1346,N_13732,N_13107);
and UO_1347 (O_1347,N_14145,N_12028);
or UO_1348 (O_1348,N_11910,N_11636);
or UO_1349 (O_1349,N_12325,N_13409);
or UO_1350 (O_1350,N_14923,N_12240);
or UO_1351 (O_1351,N_13300,N_13734);
xor UO_1352 (O_1352,N_13274,N_11226);
or UO_1353 (O_1353,N_12908,N_11616);
nand UO_1354 (O_1354,N_10654,N_10912);
or UO_1355 (O_1355,N_12156,N_12838);
xor UO_1356 (O_1356,N_14916,N_11286);
or UO_1357 (O_1357,N_11405,N_14012);
or UO_1358 (O_1358,N_13396,N_14346);
nand UO_1359 (O_1359,N_14758,N_12558);
nor UO_1360 (O_1360,N_14175,N_12631);
and UO_1361 (O_1361,N_14827,N_11686);
xnor UO_1362 (O_1362,N_14159,N_14716);
nand UO_1363 (O_1363,N_14907,N_11831);
xnor UO_1364 (O_1364,N_11643,N_13517);
nor UO_1365 (O_1365,N_12859,N_12599);
nor UO_1366 (O_1366,N_13417,N_13896);
xor UO_1367 (O_1367,N_10559,N_12592);
nor UO_1368 (O_1368,N_11772,N_10870);
nor UO_1369 (O_1369,N_12917,N_14170);
xnor UO_1370 (O_1370,N_11154,N_13909);
nor UO_1371 (O_1371,N_10658,N_12007);
or UO_1372 (O_1372,N_14780,N_14997);
nand UO_1373 (O_1373,N_11054,N_13862);
nand UO_1374 (O_1374,N_10312,N_11027);
xnor UO_1375 (O_1375,N_13035,N_14032);
nand UO_1376 (O_1376,N_11184,N_10107);
or UO_1377 (O_1377,N_10813,N_13454);
nand UO_1378 (O_1378,N_14721,N_11474);
and UO_1379 (O_1379,N_11805,N_12800);
nor UO_1380 (O_1380,N_11877,N_14435);
nor UO_1381 (O_1381,N_13302,N_10325);
nand UO_1382 (O_1382,N_13787,N_14312);
nand UO_1383 (O_1383,N_14011,N_13783);
and UO_1384 (O_1384,N_13504,N_14405);
nand UO_1385 (O_1385,N_10114,N_11307);
and UO_1386 (O_1386,N_14792,N_11663);
nand UO_1387 (O_1387,N_11440,N_10517);
nand UO_1388 (O_1388,N_11023,N_10315);
nor UO_1389 (O_1389,N_11177,N_12326);
nor UO_1390 (O_1390,N_14389,N_11898);
nand UO_1391 (O_1391,N_10637,N_10788);
xnor UO_1392 (O_1392,N_10636,N_14785);
nor UO_1393 (O_1393,N_12746,N_11052);
and UO_1394 (O_1394,N_13312,N_12847);
or UO_1395 (O_1395,N_10106,N_12949);
nand UO_1396 (O_1396,N_14102,N_14777);
nand UO_1397 (O_1397,N_13342,N_12594);
and UO_1398 (O_1398,N_10028,N_13050);
nor UO_1399 (O_1399,N_14438,N_11160);
xnor UO_1400 (O_1400,N_14877,N_13095);
nand UO_1401 (O_1401,N_14205,N_10033);
and UO_1402 (O_1402,N_13428,N_11015);
and UO_1403 (O_1403,N_10744,N_14664);
or UO_1404 (O_1404,N_11419,N_11216);
xnor UO_1405 (O_1405,N_14441,N_10195);
nor UO_1406 (O_1406,N_11080,N_12454);
nand UO_1407 (O_1407,N_14424,N_12688);
nor UO_1408 (O_1408,N_14855,N_12734);
nand UO_1409 (O_1409,N_14443,N_14536);
and UO_1410 (O_1410,N_10270,N_11582);
nor UO_1411 (O_1411,N_10187,N_11781);
xnor UO_1412 (O_1412,N_13178,N_13473);
nand UO_1413 (O_1413,N_12582,N_10701);
nor UO_1414 (O_1414,N_10715,N_12101);
or UO_1415 (O_1415,N_14663,N_12716);
nor UO_1416 (O_1416,N_12405,N_10541);
xnor UO_1417 (O_1417,N_10693,N_13287);
or UO_1418 (O_1418,N_13641,N_14922);
or UO_1419 (O_1419,N_11134,N_14092);
xnor UO_1420 (O_1420,N_11297,N_13906);
nand UO_1421 (O_1421,N_11236,N_10655);
xor UO_1422 (O_1422,N_11868,N_13198);
xnor UO_1423 (O_1423,N_10766,N_12525);
xor UO_1424 (O_1424,N_11495,N_11981);
xnor UO_1425 (O_1425,N_10883,N_12730);
or UO_1426 (O_1426,N_12633,N_10502);
xnor UO_1427 (O_1427,N_11509,N_12853);
or UO_1428 (O_1428,N_12537,N_10083);
xor UO_1429 (O_1429,N_12167,N_13755);
nor UO_1430 (O_1430,N_12441,N_11321);
or UO_1431 (O_1431,N_12236,N_14329);
nand UO_1432 (O_1432,N_14506,N_10776);
xor UO_1433 (O_1433,N_10587,N_12675);
xor UO_1434 (O_1434,N_14816,N_14447);
xnor UO_1435 (O_1435,N_14833,N_14985);
nor UO_1436 (O_1436,N_14546,N_10971);
and UO_1437 (O_1437,N_13653,N_11924);
and UO_1438 (O_1438,N_12464,N_14523);
or UO_1439 (O_1439,N_12099,N_10358);
nor UO_1440 (O_1440,N_10035,N_14158);
nor UO_1441 (O_1441,N_13752,N_10481);
nor UO_1442 (O_1442,N_12342,N_14893);
nand UO_1443 (O_1443,N_11106,N_12986);
nand UO_1444 (O_1444,N_13951,N_11912);
or UO_1445 (O_1445,N_14511,N_10420);
xnor UO_1446 (O_1446,N_11714,N_14121);
xnor UO_1447 (O_1447,N_12555,N_11214);
xnor UO_1448 (O_1448,N_11206,N_14379);
or UO_1449 (O_1449,N_11393,N_11159);
and UO_1450 (O_1450,N_12177,N_12218);
and UO_1451 (O_1451,N_11379,N_13369);
nor UO_1452 (O_1452,N_11720,N_14357);
nor UO_1453 (O_1453,N_12297,N_13315);
xnor UO_1454 (O_1454,N_10395,N_14507);
nor UO_1455 (O_1455,N_11385,N_11030);
nor UO_1456 (O_1456,N_11397,N_11923);
and UO_1457 (O_1457,N_13229,N_11865);
xor UO_1458 (O_1458,N_13664,N_14289);
nand UO_1459 (O_1459,N_12617,N_13818);
nand UO_1460 (O_1460,N_10548,N_11199);
or UO_1461 (O_1461,N_10264,N_11083);
and UO_1462 (O_1462,N_14953,N_13425);
nand UO_1463 (O_1463,N_11149,N_14260);
nand UO_1464 (O_1464,N_13214,N_14987);
nor UO_1465 (O_1465,N_13942,N_14281);
nand UO_1466 (O_1466,N_11886,N_11560);
and UO_1467 (O_1467,N_10926,N_11951);
nor UO_1468 (O_1468,N_13368,N_10779);
nand UO_1469 (O_1469,N_14252,N_10745);
or UO_1470 (O_1470,N_11755,N_12672);
and UO_1471 (O_1471,N_11662,N_14165);
nor UO_1472 (O_1472,N_12801,N_14173);
nor UO_1473 (O_1473,N_12150,N_11632);
nand UO_1474 (O_1474,N_14395,N_11980);
nor UO_1475 (O_1475,N_13515,N_12185);
nor UO_1476 (O_1476,N_13400,N_13933);
nor UO_1477 (O_1477,N_12705,N_10265);
nand UO_1478 (O_1478,N_11062,N_14182);
or UO_1479 (O_1479,N_12958,N_13467);
nor UO_1480 (O_1480,N_12745,N_14317);
and UO_1481 (O_1481,N_14493,N_10120);
nand UO_1482 (O_1482,N_12105,N_11303);
xor UO_1483 (O_1483,N_11999,N_12068);
xnor UO_1484 (O_1484,N_14951,N_11931);
xor UO_1485 (O_1485,N_11173,N_10617);
xnor UO_1486 (O_1486,N_11335,N_14930);
and UO_1487 (O_1487,N_11090,N_10464);
and UO_1488 (O_1488,N_13802,N_13883);
nor UO_1489 (O_1489,N_10384,N_12584);
xor UO_1490 (O_1490,N_12670,N_13068);
xor UO_1491 (O_1491,N_12754,N_10987);
nand UO_1492 (O_1492,N_10730,N_10946);
nor UO_1493 (O_1493,N_11588,N_11365);
xnor UO_1494 (O_1494,N_13082,N_12331);
nor UO_1495 (O_1495,N_12812,N_13471);
or UO_1496 (O_1496,N_11590,N_13438);
nor UO_1497 (O_1497,N_14201,N_11620);
xnor UO_1498 (O_1498,N_10614,N_13512);
xnor UO_1499 (O_1499,N_13132,N_14652);
nand UO_1500 (O_1500,N_11124,N_13285);
xor UO_1501 (O_1501,N_13815,N_10934);
and UO_1502 (O_1502,N_14913,N_14325);
and UO_1503 (O_1503,N_13290,N_12403);
or UO_1504 (O_1504,N_10303,N_11341);
or UO_1505 (O_1505,N_14413,N_13463);
or UO_1506 (O_1506,N_14207,N_14943);
nor UO_1507 (O_1507,N_14142,N_13231);
nor UO_1508 (O_1508,N_12613,N_14748);
and UO_1509 (O_1509,N_13343,N_14361);
xor UO_1510 (O_1510,N_13682,N_14961);
nor UO_1511 (O_1511,N_13622,N_12035);
nor UO_1512 (O_1512,N_13820,N_13464);
or UO_1513 (O_1513,N_13477,N_14247);
or UO_1514 (O_1514,N_11558,N_10545);
nand UO_1515 (O_1515,N_10707,N_11970);
nand UO_1516 (O_1516,N_13928,N_11512);
and UO_1517 (O_1517,N_11876,N_12163);
nor UO_1518 (O_1518,N_10183,N_11966);
and UO_1519 (O_1519,N_13608,N_11602);
nor UO_1520 (O_1520,N_14693,N_11223);
and UO_1521 (O_1521,N_10039,N_13296);
xor UO_1522 (O_1522,N_14027,N_13824);
or UO_1523 (O_1523,N_11699,N_13613);
and UO_1524 (O_1524,N_13345,N_13785);
nand UO_1525 (O_1525,N_13341,N_13658);
or UO_1526 (O_1526,N_13167,N_13651);
xnor UO_1527 (O_1527,N_11854,N_13508);
nand UO_1528 (O_1528,N_10671,N_11906);
nor UO_1529 (O_1529,N_12152,N_10382);
nor UO_1530 (O_1530,N_10229,N_10811);
or UO_1531 (O_1531,N_13872,N_11893);
or UO_1532 (O_1532,N_12879,N_13031);
or UO_1533 (O_1533,N_13261,N_12046);
or UO_1534 (O_1534,N_13248,N_14921);
xor UO_1535 (O_1535,N_11074,N_14183);
or UO_1536 (O_1536,N_10585,N_13976);
or UO_1537 (O_1537,N_14601,N_13948);
nand UO_1538 (O_1538,N_10361,N_14154);
nor UO_1539 (O_1539,N_11118,N_14553);
nand UO_1540 (O_1540,N_11268,N_12475);
and UO_1541 (O_1541,N_10628,N_10969);
nor UO_1542 (O_1542,N_10645,N_11698);
and UO_1543 (O_1543,N_10708,N_12442);
xnor UO_1544 (O_1544,N_13165,N_11270);
nor UO_1545 (O_1545,N_11330,N_14939);
nand UO_1546 (O_1546,N_13058,N_11690);
xor UO_1547 (O_1547,N_12269,N_14835);
and UO_1548 (O_1548,N_13338,N_12423);
nor UO_1549 (O_1549,N_11449,N_12509);
nand UO_1550 (O_1550,N_14879,N_14308);
nand UO_1551 (O_1551,N_13941,N_13996);
xnor UO_1552 (O_1552,N_11348,N_12969);
nand UO_1553 (O_1553,N_14351,N_14323);
nand UO_1554 (O_1554,N_12283,N_13385);
xnor UO_1555 (O_1555,N_12676,N_13952);
nor UO_1556 (O_1556,N_13794,N_10796);
xor UO_1557 (O_1557,N_11443,N_10760);
nand UO_1558 (O_1558,N_14147,N_11108);
nand UO_1559 (O_1559,N_12019,N_12488);
and UO_1560 (O_1560,N_10880,N_13863);
and UO_1561 (O_1561,N_12541,N_12864);
xnor UO_1562 (O_1562,N_12247,N_14846);
nand UO_1563 (O_1563,N_10306,N_12567);
nor UO_1564 (O_1564,N_11878,N_14898);
nor UO_1565 (O_1565,N_10118,N_11112);
nor UO_1566 (O_1566,N_10040,N_12205);
nand UO_1567 (O_1567,N_12713,N_12715);
nor UO_1568 (O_1568,N_12410,N_13026);
nand UO_1569 (O_1569,N_11697,N_14890);
or UO_1570 (O_1570,N_12445,N_11791);
and UO_1571 (O_1571,N_13066,N_12091);
or UO_1572 (O_1572,N_13394,N_10827);
xnor UO_1573 (O_1573,N_13418,N_11534);
nand UO_1574 (O_1574,N_10984,N_11208);
and UO_1575 (O_1575,N_13637,N_12221);
xor UO_1576 (O_1576,N_14456,N_10475);
and UO_1577 (O_1577,N_11668,N_14494);
or UO_1578 (O_1578,N_12349,N_11325);
nor UO_1579 (O_1579,N_10268,N_10473);
and UO_1580 (O_1580,N_13628,N_10389);
nand UO_1581 (O_1581,N_11973,N_13778);
xor UO_1582 (O_1582,N_14242,N_10447);
or UO_1583 (O_1583,N_13399,N_13606);
xor UO_1584 (O_1584,N_14180,N_12985);
nand UO_1585 (O_1585,N_13208,N_11984);
and UO_1586 (O_1586,N_13795,N_14366);
nand UO_1587 (O_1587,N_12246,N_10684);
nor UO_1588 (O_1588,N_11596,N_13520);
or UO_1589 (O_1589,N_11504,N_13575);
nand UO_1590 (O_1590,N_12832,N_12775);
nand UO_1591 (O_1591,N_14711,N_10087);
xnor UO_1592 (O_1592,N_13754,N_13240);
and UO_1593 (O_1593,N_12647,N_12398);
nor UO_1594 (O_1594,N_13610,N_12380);
xnor UO_1595 (O_1595,N_12736,N_10094);
and UO_1596 (O_1596,N_11622,N_14057);
xnor UO_1597 (O_1597,N_10011,N_14268);
xnor UO_1598 (O_1598,N_12196,N_13390);
and UO_1599 (O_1599,N_13259,N_14403);
xor UO_1600 (O_1600,N_12089,N_13727);
nand UO_1601 (O_1601,N_14459,N_11273);
or UO_1602 (O_1602,N_13236,N_11675);
xor UO_1603 (O_1603,N_13561,N_11398);
nand UO_1604 (O_1604,N_12874,N_13267);
xnor UO_1605 (O_1605,N_14338,N_13735);
nor UO_1606 (O_1606,N_10103,N_14883);
nand UO_1607 (O_1607,N_10657,N_14667);
or UO_1608 (O_1608,N_13969,N_14387);
nor UO_1609 (O_1609,N_12523,N_10632);
and UO_1610 (O_1610,N_11136,N_13363);
xor UO_1611 (O_1611,N_10627,N_11050);
and UO_1612 (O_1612,N_11625,N_11757);
xor UO_1613 (O_1613,N_10951,N_12600);
xor UO_1614 (O_1614,N_10889,N_14692);
nand UO_1615 (O_1615,N_10206,N_11164);
and UO_1616 (O_1616,N_14878,N_13586);
nor UO_1617 (O_1617,N_11793,N_14369);
or UO_1618 (O_1618,N_13111,N_10823);
or UO_1619 (O_1619,N_14072,N_12533);
or UO_1620 (O_1620,N_11078,N_14657);
xor UO_1621 (O_1621,N_11633,N_13546);
nor UO_1622 (O_1622,N_10443,N_14767);
or UO_1623 (O_1623,N_13897,N_14250);
nand UO_1624 (O_1624,N_13819,N_12643);
nor UO_1625 (O_1625,N_10862,N_11437);
or UO_1626 (O_1626,N_14954,N_12809);
and UO_1627 (O_1627,N_14694,N_10267);
or UO_1628 (O_1628,N_11444,N_10432);
nand UO_1629 (O_1629,N_12833,N_10001);
nor UO_1630 (O_1630,N_12861,N_10868);
xor UO_1631 (O_1631,N_10491,N_14500);
xor UO_1632 (O_1632,N_11441,N_11655);
nand UO_1633 (O_1633,N_10620,N_13991);
xnor UO_1634 (O_1634,N_10718,N_12160);
xnor UO_1635 (O_1635,N_11157,N_13374);
xor UO_1636 (O_1636,N_12378,N_12299);
nand UO_1637 (O_1637,N_11676,N_13023);
nand UO_1638 (O_1638,N_13465,N_12034);
nand UO_1639 (O_1639,N_14519,N_12665);
nor UO_1640 (O_1640,N_10775,N_14788);
nor UO_1641 (O_1641,N_10652,N_12169);
xnor UO_1642 (O_1642,N_10046,N_11613);
or UO_1643 (O_1643,N_10750,N_10792);
nor UO_1644 (O_1644,N_12965,N_14592);
and UO_1645 (O_1645,N_10734,N_14209);
nand UO_1646 (O_1646,N_10075,N_13275);
or UO_1647 (O_1647,N_14467,N_14830);
or UO_1648 (O_1648,N_11336,N_13782);
xnor UO_1649 (O_1649,N_14998,N_10830);
or UO_1650 (O_1650,N_10131,N_13822);
nor UO_1651 (O_1651,N_12010,N_10455);
xnor UO_1652 (O_1652,N_13129,N_14978);
nand UO_1653 (O_1653,N_11994,N_11326);
xnor UO_1654 (O_1654,N_14157,N_12309);
or UO_1655 (O_1655,N_13656,N_14965);
and UO_1656 (O_1656,N_10091,N_13747);
and UO_1657 (O_1657,N_10026,N_14678);
or UO_1658 (O_1658,N_13145,N_11592);
nor UO_1659 (O_1659,N_10439,N_10327);
nor UO_1660 (O_1660,N_12107,N_10538);
nor UO_1661 (O_1661,N_12361,N_13093);
and UO_1662 (O_1662,N_12093,N_12962);
and UO_1663 (O_1663,N_11779,N_10913);
nand UO_1664 (O_1664,N_12391,N_13490);
and UO_1665 (O_1665,N_12394,N_12045);
xor UO_1666 (O_1666,N_11014,N_14054);
or UO_1667 (O_1667,N_13541,N_12332);
nor UO_1668 (O_1668,N_13946,N_12500);
nand UO_1669 (O_1669,N_13482,N_13118);
nor UO_1670 (O_1670,N_12863,N_12881);
and UO_1671 (O_1671,N_11502,N_12390);
nand UO_1672 (O_1672,N_11761,N_10623);
xor UO_1673 (O_1673,N_12171,N_12289);
xnor UO_1674 (O_1674,N_11344,N_13055);
xor UO_1675 (O_1675,N_11997,N_10519);
and UO_1676 (O_1676,N_11807,N_11240);
and UO_1677 (O_1677,N_11646,N_11265);
xor UO_1678 (O_1678,N_10977,N_12577);
nand UO_1679 (O_1679,N_14061,N_10673);
nor UO_1680 (O_1680,N_14223,N_11388);
or UO_1681 (O_1681,N_14065,N_14125);
nor UO_1682 (O_1682,N_12463,N_14935);
nand UO_1683 (O_1683,N_14008,N_14340);
xor UO_1684 (O_1684,N_12401,N_12242);
nand UO_1685 (O_1685,N_11162,N_11871);
or UO_1686 (O_1686,N_13593,N_10080);
xor UO_1687 (O_1687,N_10678,N_12440);
and UO_1688 (O_1688,N_14912,N_13889);
and UO_1689 (O_1689,N_14114,N_10066);
and UO_1690 (O_1690,N_14080,N_12212);
or UO_1691 (O_1691,N_14304,N_13001);
nor UO_1692 (O_1692,N_13387,N_10002);
nor UO_1693 (O_1693,N_14754,N_11481);
or UO_1694 (O_1694,N_10397,N_12725);
nor UO_1695 (O_1695,N_12837,N_10925);
nor UO_1696 (O_1696,N_12508,N_10600);
or UO_1697 (O_1697,N_11840,N_14680);
nor UO_1698 (O_1698,N_13762,N_12971);
and UO_1699 (O_1699,N_12032,N_14989);
or UO_1700 (O_1700,N_14163,N_12578);
and UO_1701 (O_1701,N_10049,N_13384);
nor UO_1702 (O_1702,N_13847,N_14908);
nand UO_1703 (O_1703,N_14936,N_13439);
nor UO_1704 (O_1704,N_14910,N_13571);
and UO_1705 (O_1705,N_12565,N_13914);
nand UO_1706 (O_1706,N_11820,N_12904);
nand UO_1707 (O_1707,N_14078,N_11183);
xor UO_1708 (O_1708,N_13176,N_12175);
and UO_1709 (O_1709,N_12620,N_11197);
and UO_1710 (O_1710,N_13744,N_13926);
nor UO_1711 (O_1711,N_13798,N_12137);
nor UO_1712 (O_1712,N_10644,N_13378);
nor UO_1713 (O_1713,N_14842,N_12916);
or UO_1714 (O_1714,N_12455,N_12968);
nand UO_1715 (O_1715,N_14422,N_12179);
and UO_1716 (O_1716,N_14446,N_13680);
and UO_1717 (O_1717,N_14273,N_11665);
or UO_1718 (O_1718,N_14120,N_12942);
nor UO_1719 (O_1719,N_11158,N_10275);
and UO_1720 (O_1720,N_11671,N_11750);
nor UO_1721 (O_1721,N_14038,N_10467);
xor UO_1722 (O_1722,N_14584,N_12296);
or UO_1723 (O_1723,N_13172,N_14867);
and UO_1724 (O_1724,N_11522,N_10535);
nor UO_1725 (O_1725,N_11580,N_10378);
or UO_1726 (O_1726,N_10479,N_13743);
xnor UO_1727 (O_1727,N_10863,N_13756);
or UO_1728 (O_1728,N_11576,N_12731);
and UO_1729 (O_1729,N_13902,N_11594);
and UO_1730 (O_1730,N_12943,N_14926);
xnor UO_1731 (O_1731,N_10949,N_10410);
xor UO_1732 (O_1732,N_13898,N_14076);
nor UO_1733 (O_1733,N_12489,N_14874);
nand UO_1734 (O_1734,N_11979,N_14541);
and UO_1735 (O_1735,N_14903,N_10665);
xor UO_1736 (O_1736,N_11476,N_11429);
nor UO_1737 (O_1737,N_11583,N_13244);
or UO_1738 (O_1738,N_14483,N_12191);
or UO_1739 (O_1739,N_13931,N_10679);
nor UO_1740 (O_1740,N_10694,N_10181);
nand UO_1741 (O_1741,N_14738,N_14558);
or UO_1742 (O_1742,N_13484,N_11423);
nor UO_1743 (O_1743,N_14486,N_10019);
xnor UO_1744 (O_1744,N_13170,N_13828);
nand UO_1745 (O_1745,N_10512,N_13466);
xor UO_1746 (O_1746,N_12389,N_13087);
and UO_1747 (O_1747,N_13980,N_11427);
xor UO_1748 (O_1748,N_11012,N_10493);
nand UO_1749 (O_1749,N_10076,N_10061);
nand UO_1750 (O_1750,N_11520,N_13072);
nor UO_1751 (O_1751,N_10805,N_10166);
and UO_1752 (O_1752,N_12632,N_10716);
or UO_1753 (O_1753,N_12970,N_12706);
nor UO_1754 (O_1754,N_10899,N_10878);
nor UO_1755 (O_1755,N_12590,N_11256);
xor UO_1756 (O_1756,N_13008,N_14860);
nor UO_1757 (O_1757,N_14396,N_11919);
or UO_1758 (O_1758,N_13386,N_11046);
nor UO_1759 (O_1759,N_14590,N_13048);
nand UO_1760 (O_1760,N_13375,N_14309);
nor UO_1761 (O_1761,N_11754,N_12144);
xor UO_1762 (O_1762,N_10791,N_11647);
or UO_1763 (O_1763,N_10997,N_14297);
nor UO_1764 (O_1764,N_14565,N_11615);
nor UO_1765 (O_1765,N_13619,N_12722);
nand UO_1766 (O_1766,N_10911,N_11086);
and UO_1767 (O_1767,N_10207,N_14249);
nand UO_1768 (O_1768,N_11821,N_11607);
and UO_1769 (O_1769,N_14271,N_13623);
and UO_1770 (O_1770,N_13673,N_11372);
and UO_1771 (O_1771,N_14808,N_12909);
nor UO_1772 (O_1772,N_13662,N_10319);
and UO_1773 (O_1773,N_13746,N_13108);
or UO_1774 (O_1774,N_14990,N_11810);
and UO_1775 (O_1775,N_13685,N_10167);
and UO_1776 (O_1776,N_13771,N_14171);
nor UO_1777 (O_1777,N_10935,N_12834);
and UO_1778 (O_1778,N_14272,N_11049);
and UO_1779 (O_1779,N_13767,N_10558);
and UO_1780 (O_1780,N_13189,N_11005);
and UO_1781 (O_1781,N_10669,N_12903);
nor UO_1782 (O_1782,N_10626,N_11031);
or UO_1783 (O_1783,N_12910,N_11098);
nand UO_1784 (O_1784,N_13196,N_12692);
nand UO_1785 (O_1785,N_11850,N_11631);
nor UO_1786 (O_1786,N_12038,N_10052);
and UO_1787 (O_1787,N_12125,N_14010);
nor UO_1788 (O_1788,N_10547,N_13344);
xor UO_1789 (O_1789,N_10624,N_13376);
nand UO_1790 (O_1790,N_12393,N_13983);
or UO_1791 (O_1791,N_13488,N_10177);
or UO_1792 (O_1792,N_11188,N_10105);
or UO_1793 (O_1793,N_14599,N_12922);
or UO_1794 (O_1794,N_11513,N_10885);
xnor UO_1795 (O_1795,N_11401,N_12933);
nor UO_1796 (O_1796,N_12053,N_10514);
or UO_1797 (O_1797,N_11621,N_13029);
nand UO_1798 (O_1798,N_10108,N_12276);
nor UO_1799 (O_1799,N_14445,N_11150);
and UO_1800 (O_1800,N_11873,N_10793);
and UO_1801 (O_1801,N_10888,N_11250);
nor UO_1802 (O_1802,N_11122,N_10354);
xnor UO_1803 (O_1803,N_14981,N_13461);
xnor UO_1804 (O_1804,N_13469,N_11219);
or UO_1805 (O_1805,N_12227,N_11695);
xor UO_1806 (O_1806,N_12126,N_12225);
nor UO_1807 (O_1807,N_11056,N_12811);
and UO_1808 (O_1808,N_11586,N_11799);
and UO_1809 (O_1809,N_11167,N_10459);
and UO_1810 (O_1810,N_11094,N_13671);
xor UO_1811 (O_1811,N_13612,N_11901);
or UO_1812 (O_1812,N_13105,N_11492);
or UO_1813 (O_1813,N_12639,N_11909);
nand UO_1814 (O_1814,N_10244,N_13638);
xor UO_1815 (O_1815,N_14107,N_14400);
and UO_1816 (O_1816,N_11267,N_12124);
nand UO_1817 (O_1817,N_12638,N_14563);
nor UO_1818 (O_1818,N_11490,N_11243);
or UO_1819 (O_1819,N_14333,N_10875);
nor UO_1820 (O_1820,N_13474,N_14122);
nand UO_1821 (O_1821,N_12162,N_13437);
or UO_1822 (O_1822,N_14168,N_11346);
nand UO_1823 (O_1823,N_14927,N_12925);
and UO_1824 (O_1824,N_11666,N_13119);
nand UO_1825 (O_1825,N_12434,N_13413);
nand UO_1826 (O_1826,N_11562,N_13768);
nand UO_1827 (O_1827,N_13950,N_10954);
and UO_1828 (O_1828,N_11231,N_11306);
or UO_1829 (O_1829,N_12473,N_12360);
xor UO_1830 (O_1830,N_10012,N_10331);
nor UO_1831 (O_1831,N_11837,N_11451);
or UO_1832 (O_1832,N_11259,N_14356);
xnor UO_1833 (O_1833,N_11276,N_10844);
and UO_1834 (O_1834,N_12752,N_13974);
and UO_1835 (O_1835,N_11618,N_12797);
xor UO_1836 (O_1836,N_10188,N_11156);
nand UO_1837 (O_1837,N_13336,N_13005);
nand UO_1838 (O_1838,N_14611,N_10629);
or UO_1839 (O_1839,N_11230,N_11435);
nand UO_1840 (O_1840,N_11800,N_14594);
xor UO_1841 (O_1841,N_14301,N_13282);
nand UO_1842 (O_1842,N_14410,N_11735);
and UO_1843 (O_1843,N_12011,N_11693);
nor UO_1844 (O_1844,N_14787,N_12315);
nor UO_1845 (O_1845,N_14153,N_13281);
or UO_1846 (O_1846,N_12451,N_11789);
and UO_1847 (O_1847,N_12553,N_13566);
nor UO_1848 (O_1848,N_14198,N_13710);
nand UO_1849 (O_1849,N_13632,N_10231);
nand UO_1850 (O_1850,N_10059,N_13726);
nor UO_1851 (O_1851,N_10769,N_13837);
nor UO_1852 (O_1852,N_12940,N_12113);
nor UO_1853 (O_1853,N_13091,N_13002);
nand UO_1854 (O_1854,N_10098,N_14043);
nor UO_1855 (O_1855,N_11673,N_11205);
xor UO_1856 (O_1856,N_12408,N_12228);
and UO_1857 (O_1857,N_13595,N_11421);
or UO_1858 (O_1858,N_13882,N_10714);
or UO_1859 (O_1859,N_10450,N_12539);
or UO_1860 (O_1860,N_13084,N_12673);
nand UO_1861 (O_1861,N_13514,N_14337);
xor UO_1862 (O_1862,N_10746,N_10104);
or UO_1863 (O_1863,N_12980,N_10391);
xnor UO_1864 (O_1864,N_11650,N_13216);
and UO_1865 (O_1865,N_11767,N_10843);
or UO_1866 (O_1866,N_13397,N_13276);
and UO_1867 (O_1867,N_10055,N_10808);
nand UO_1868 (O_1868,N_13329,N_13371);
nand UO_1869 (O_1869,N_13351,N_13160);
or UO_1870 (O_1870,N_11905,N_11925);
xnor UO_1871 (O_1871,N_13447,N_12000);
and UO_1872 (O_1872,N_13686,N_12564);
xnor UO_1873 (O_1873,N_10130,N_14029);
nor UO_1874 (O_1874,N_14058,N_12456);
nand UO_1875 (O_1875,N_10259,N_14162);
nand UO_1876 (O_1876,N_10255,N_13763);
and UO_1877 (O_1877,N_10897,N_12660);
or UO_1878 (O_1878,N_14676,N_10505);
or UO_1879 (O_1879,N_13574,N_12583);
and UO_1880 (O_1880,N_14763,N_10489);
xnor UO_1881 (O_1881,N_11503,N_14148);
and UO_1882 (O_1882,N_10415,N_10413);
xor UO_1883 (O_1883,N_14776,N_12418);
and UO_1884 (O_1884,N_14019,N_14911);
nand UO_1885 (O_1885,N_11361,N_12987);
nand UO_1886 (O_1886,N_14897,N_13407);
nand UO_1887 (O_1887,N_11009,N_12823);
nor UO_1888 (O_1888,N_12471,N_11453);
nand UO_1889 (O_1889,N_14007,N_13191);
and UO_1890 (O_1890,N_11832,N_12507);
xnor UO_1891 (O_1891,N_14892,N_12097);
and UO_1892 (O_1892,N_12253,N_10110);
nor UO_1893 (O_1893,N_11308,N_11722);
nor UO_1894 (O_1894,N_10162,N_11962);
nor UO_1895 (O_1895,N_10972,N_11764);
and UO_1896 (O_1896,N_13659,N_11521);
nand UO_1897 (O_1897,N_10205,N_14190);
xor UO_1898 (O_1898,N_11390,N_13305);
nor UO_1899 (O_1899,N_12478,N_10366);
nor UO_1900 (O_1900,N_13945,N_14636);
xnor UO_1901 (O_1901,N_13990,N_11982);
or UO_1902 (O_1902,N_11198,N_10840);
or UO_1903 (O_1903,N_14873,N_11232);
nor UO_1904 (O_1904,N_11482,N_10703);
nand UO_1905 (O_1905,N_12272,N_12981);
and UO_1906 (O_1906,N_11040,N_14150);
nand UO_1907 (O_1907,N_10985,N_13800);
nor UO_1908 (O_1908,N_11785,N_12443);
nor UO_1909 (O_1909,N_11528,N_12697);
or UO_1910 (O_1910,N_11538,N_14381);
xnor UO_1911 (O_1911,N_11869,N_10394);
or UO_1912 (O_1912,N_10056,N_12300);
or UO_1913 (O_1913,N_14845,N_11282);
nand UO_1914 (O_1914,N_12119,N_12545);
xor UO_1915 (O_1915,N_13069,N_11360);
or UO_1916 (O_1916,N_13202,N_10735);
or UO_1917 (O_1917,N_14617,N_10140);
or UO_1918 (O_1918,N_13739,N_12890);
nand UO_1919 (O_1919,N_14896,N_12381);
or UO_1920 (O_1920,N_14176,N_13481);
nor UO_1921 (O_1921,N_14184,N_10000);
nor UO_1922 (O_1922,N_14230,N_13521);
and UO_1923 (O_1923,N_14695,N_11988);
xor UO_1924 (O_1924,N_10119,N_14531);
nor UO_1925 (O_1925,N_14623,N_11593);
or UO_1926 (O_1926,N_10472,N_12888);
nand UO_1927 (O_1927,N_14373,N_10642);
nor UO_1928 (O_1928,N_11479,N_10078);
or UO_1929 (O_1929,N_10286,N_11907);
nor UO_1930 (O_1930,N_10271,N_12065);
or UO_1931 (O_1931,N_10117,N_10043);
xnor UO_1932 (O_1932,N_14037,N_11394);
nand UO_1933 (O_1933,N_12544,N_11011);
and UO_1934 (O_1934,N_14750,N_10498);
nor UO_1935 (O_1935,N_13501,N_14134);
xnor UO_1936 (O_1936,N_11682,N_12239);
nand UO_1937 (O_1937,N_11719,N_10838);
or UO_1938 (O_1938,N_13938,N_11101);
and UO_1939 (O_1939,N_11100,N_11691);
and UO_1940 (O_1940,N_12520,N_13543);
or UO_1941 (O_1941,N_11351,N_10436);
and UO_1942 (O_1942,N_14960,N_11972);
or UO_1943 (O_1943,N_10608,N_13674);
nand UO_1944 (O_1944,N_10611,N_13854);
xor UO_1945 (O_1945,N_14152,N_10008);
nand UO_1946 (O_1946,N_12810,N_13511);
nor UO_1947 (O_1947,N_12623,N_12109);
and UO_1948 (O_1948,N_12282,N_11649);
nand UO_1949 (O_1949,N_12290,N_11302);
nand UO_1950 (O_1950,N_10686,N_10408);
or UO_1951 (O_1951,N_13445,N_14619);
nand UO_1952 (O_1952,N_11507,N_14178);
xor UO_1953 (O_1953,N_10784,N_10709);
nor UO_1954 (O_1954,N_14805,N_10643);
nor UO_1955 (O_1955,N_13116,N_14119);
xor UO_1956 (O_1956,N_14741,N_14257);
nor UO_1957 (O_1957,N_14726,N_14133);
nand UO_1958 (O_1958,N_13644,N_13645);
and UO_1959 (O_1959,N_11428,N_14041);
xor UO_1960 (O_1960,N_14241,N_10441);
and UO_1961 (O_1961,N_13014,N_14302);
and UO_1962 (O_1962,N_13532,N_12358);
nor UO_1963 (O_1963,N_11950,N_10287);
or UO_1964 (O_1964,N_10252,N_13388);
xor UO_1965 (O_1965,N_13597,N_13887);
nor UO_1966 (O_1966,N_11803,N_13288);
nor UO_1967 (O_1967,N_10449,N_10034);
or UO_1968 (O_1968,N_11338,N_14639);
xnor UO_1969 (O_1969,N_14094,N_10477);
or UO_1970 (O_1970,N_10950,N_14775);
and UO_1971 (O_1971,N_13650,N_11743);
nor UO_1972 (O_1972,N_12918,N_14225);
or UO_1973 (O_1973,N_14179,N_14784);
xor UO_1974 (O_1974,N_12244,N_10910);
xnor UO_1975 (O_1975,N_13918,N_10445);
and UO_1976 (O_1976,N_10364,N_14569);
nand UO_1977 (O_1977,N_11515,N_10974);
or UO_1978 (O_1978,N_11550,N_11685);
nor UO_1979 (O_1979,N_13354,N_11082);
and UO_1980 (O_1980,N_10706,N_11606);
nor UO_1981 (O_1981,N_12491,N_13487);
and UO_1982 (O_1982,N_12841,N_13192);
nor UO_1983 (O_1983,N_12540,N_12307);
nor UO_1984 (O_1984,N_13194,N_12174);
and UO_1985 (O_1985,N_10226,N_12129);
nor UO_1986 (O_1986,N_11672,N_11848);
xor UO_1987 (O_1987,N_13553,N_13665);
nor UO_1988 (O_1988,N_11382,N_10876);
nand UO_1989 (O_1989,N_11892,N_12721);
and UO_1990 (O_1990,N_10405,N_11459);
or UO_1991 (O_1991,N_13885,N_14372);
nand UO_1992 (O_1992,N_11875,N_13666);
nor UO_1993 (O_1993,N_12164,N_12264);
nor UO_1994 (O_1994,N_11862,N_13624);
nand UO_1995 (O_1995,N_12005,N_10903);
xnor UO_1996 (O_1996,N_12025,N_12707);
or UO_1997 (O_1997,N_14941,N_13203);
xor UO_1998 (O_1998,N_14439,N_11107);
xnor UO_1999 (O_1999,N_11585,N_13979);
endmodule