module basic_750_5000_1000_50_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_502,In_595);
and U1 (N_1,In_169,In_191);
nor U2 (N_2,In_636,In_547);
and U3 (N_3,In_190,In_469);
nand U4 (N_4,In_685,In_440);
or U5 (N_5,In_149,In_375);
nor U6 (N_6,In_543,In_50);
and U7 (N_7,In_429,In_171);
nor U8 (N_8,In_549,In_418);
or U9 (N_9,In_309,In_145);
and U10 (N_10,In_527,In_43);
nand U11 (N_11,In_295,In_715);
and U12 (N_12,In_210,In_37);
nor U13 (N_13,In_555,In_660);
nand U14 (N_14,In_187,In_120);
nor U15 (N_15,In_218,In_328);
xor U16 (N_16,In_28,In_673);
or U17 (N_17,In_147,In_220);
and U18 (N_18,In_578,In_136);
and U19 (N_19,In_367,In_53);
nand U20 (N_20,In_742,In_679);
or U21 (N_21,In_677,In_522);
nand U22 (N_22,In_513,In_669);
nand U23 (N_23,In_695,In_124);
nand U24 (N_24,In_117,In_161);
xor U25 (N_25,In_610,In_58);
and U26 (N_26,In_496,In_322);
nor U27 (N_27,In_40,In_510);
and U28 (N_28,In_457,In_259);
or U29 (N_29,In_617,In_27);
xnor U30 (N_30,In_122,In_616);
and U31 (N_31,In_420,In_545);
or U32 (N_32,In_443,In_654);
nor U33 (N_33,In_729,In_411);
or U34 (N_34,In_503,In_258);
xor U35 (N_35,In_123,In_84);
or U36 (N_36,In_376,In_554);
and U37 (N_37,In_747,In_6);
nand U38 (N_38,In_726,In_703);
and U39 (N_39,In_22,In_693);
nand U40 (N_40,In_463,In_339);
nand U41 (N_41,In_432,In_236);
nand U42 (N_42,In_38,In_459);
nand U43 (N_43,In_458,In_581);
and U44 (N_44,In_51,In_366);
or U45 (N_45,In_431,In_242);
and U46 (N_46,In_604,In_582);
and U47 (N_47,In_114,In_219);
nand U48 (N_48,In_134,In_425);
and U49 (N_49,In_738,In_714);
and U50 (N_50,In_204,In_54);
nand U51 (N_51,In_273,In_100);
or U52 (N_52,In_18,In_326);
or U53 (N_53,In_241,In_415);
nand U54 (N_54,In_629,In_72);
nand U55 (N_55,In_137,In_683);
nor U56 (N_56,In_427,In_47);
or U57 (N_57,In_202,In_437);
and U58 (N_58,In_436,In_515);
nand U59 (N_59,In_368,In_630);
or U60 (N_60,In_489,In_705);
xnor U61 (N_61,In_529,In_154);
and U62 (N_62,In_310,In_419);
and U63 (N_63,In_716,In_19);
nor U64 (N_64,In_221,In_294);
or U65 (N_65,In_324,In_166);
or U66 (N_66,In_168,In_587);
or U67 (N_67,In_377,In_181);
nor U68 (N_68,In_130,In_44);
nand U69 (N_69,In_88,In_243);
nand U70 (N_70,In_179,In_397);
nand U71 (N_71,In_645,In_113);
nor U72 (N_72,In_697,In_68);
xor U73 (N_73,In_129,In_434);
xor U74 (N_74,In_281,In_460);
nand U75 (N_75,In_721,In_495);
nor U76 (N_76,In_699,In_234);
or U77 (N_77,In_369,In_409);
or U78 (N_78,In_125,In_265);
and U79 (N_79,In_280,In_652);
or U80 (N_80,In_135,In_674);
or U81 (N_81,In_602,In_702);
or U82 (N_82,In_183,In_186);
nand U83 (N_83,In_539,In_570);
nor U84 (N_84,In_665,In_141);
nor U85 (N_85,In_173,In_524);
nor U86 (N_86,In_533,In_170);
or U87 (N_87,In_650,In_453);
xnor U88 (N_88,In_467,In_269);
and U89 (N_89,In_25,In_379);
and U90 (N_90,In_151,In_678);
nor U91 (N_91,In_52,In_518);
xor U92 (N_92,In_658,In_385);
xor U93 (N_93,In_10,In_526);
nand U94 (N_94,In_207,In_481);
xor U95 (N_95,In_593,In_416);
nor U96 (N_96,In_253,In_138);
nand U97 (N_97,In_468,In_689);
and U98 (N_98,In_709,In_198);
and U99 (N_99,In_567,In_89);
nor U100 (N_100,In_492,In_724);
nand U101 (N_101,In_192,N_80);
and U102 (N_102,In_732,In_164);
xor U103 (N_103,In_748,In_316);
and U104 (N_104,N_7,In_337);
or U105 (N_105,In_395,In_390);
nand U106 (N_106,In_277,In_291);
and U107 (N_107,In_189,In_574);
or U108 (N_108,In_249,In_107);
nand U109 (N_109,In_426,In_354);
and U110 (N_110,In_162,In_256);
nand U111 (N_111,N_58,In_470);
and U112 (N_112,In_165,In_392);
nand U113 (N_113,N_8,In_178);
and U114 (N_114,In_696,In_384);
nor U115 (N_115,N_23,In_306);
nor U116 (N_116,In_564,In_201);
xor U117 (N_117,In_386,In_356);
and U118 (N_118,In_410,In_150);
xor U119 (N_119,In_508,In_235);
nor U120 (N_120,In_180,In_13);
nor U121 (N_121,In_304,In_723);
and U122 (N_122,N_22,In_225);
nor U123 (N_123,In_512,In_506);
and U124 (N_124,N_94,In_176);
or U125 (N_125,In_586,In_535);
or U126 (N_126,N_10,In_692);
xor U127 (N_127,In_653,In_23);
xnor U128 (N_128,N_3,In_623);
nor U129 (N_129,In_655,In_589);
and U130 (N_130,In_139,In_101);
and U131 (N_131,In_625,In_77);
nor U132 (N_132,In_483,In_327);
nand U133 (N_133,In_528,In_577);
nor U134 (N_134,In_296,In_501);
or U135 (N_135,In_142,In_228);
or U136 (N_136,N_51,N_72);
nor U137 (N_137,N_12,In_601);
or U138 (N_138,In_321,In_93);
or U139 (N_139,In_303,In_659);
xnor U140 (N_140,In_98,In_559);
nand U141 (N_141,In_30,In_494);
and U142 (N_142,In_487,In_507);
nor U143 (N_143,In_81,In_194);
nand U144 (N_144,N_62,In_741);
xnor U145 (N_145,In_305,In_214);
xor U146 (N_146,N_38,In_223);
or U147 (N_147,In_509,In_371);
nand U148 (N_148,In_360,In_278);
or U149 (N_149,In_355,In_465);
nand U150 (N_150,In_378,In_598);
nand U151 (N_151,In_284,In_103);
nand U152 (N_152,In_229,N_69);
and U153 (N_153,In_745,In_553);
and U154 (N_154,In_102,In_605);
nor U155 (N_155,N_4,In_21);
xor U156 (N_156,In_346,N_30);
and U157 (N_157,N_87,In_631);
nand U158 (N_158,In_690,In_76);
or U159 (N_159,In_153,In_11);
and U160 (N_160,In_148,In_591);
nor U161 (N_161,In_711,In_222);
or U162 (N_162,In_710,In_232);
nand U163 (N_163,In_448,In_664);
and U164 (N_164,N_55,N_28);
or U165 (N_165,In_661,N_26);
and U166 (N_166,N_5,N_19);
nor U167 (N_167,In_621,In_740);
nor U168 (N_168,In_473,In_29);
or U169 (N_169,In_330,In_572);
or U170 (N_170,In_466,In_600);
or U171 (N_171,In_66,In_16);
nand U172 (N_172,In_442,In_302);
and U173 (N_173,In_521,In_195);
nor U174 (N_174,N_2,In_238);
and U175 (N_175,N_43,In_87);
nand U176 (N_176,In_637,In_594);
nor U177 (N_177,In_612,In_708);
nor U178 (N_178,N_97,In_211);
and U179 (N_179,In_405,In_676);
or U180 (N_180,In_647,In_184);
nand U181 (N_181,In_86,In_199);
and U182 (N_182,In_333,In_718);
xor U183 (N_183,In_701,In_35);
nand U184 (N_184,In_694,In_618);
nor U185 (N_185,In_566,In_633);
nand U186 (N_186,In_65,In_110);
nand U187 (N_187,In_585,In_413);
nor U188 (N_188,In_583,In_290);
or U189 (N_189,In_670,N_16);
nor U190 (N_190,In_41,In_562);
and U191 (N_191,In_71,In_287);
or U192 (N_192,In_728,In_331);
xnor U193 (N_193,N_50,In_688);
and U194 (N_194,In_450,In_456);
nand U195 (N_195,In_224,In_441);
or U196 (N_196,In_364,In_83);
nand U197 (N_197,In_200,In_212);
and U198 (N_198,In_462,N_46);
nand U199 (N_199,N_82,N_91);
and U200 (N_200,In_540,In_252);
nand U201 (N_201,In_109,In_254);
nand U202 (N_202,N_9,In_606);
nand U203 (N_203,In_641,In_428);
nor U204 (N_204,N_192,In_584);
or U205 (N_205,In_511,In_447);
or U206 (N_206,N_96,In_603);
nor U207 (N_207,N_78,In_336);
nand U208 (N_208,In_451,N_57);
nor U209 (N_209,In_56,N_182);
nand U210 (N_210,In_244,N_140);
nor U211 (N_211,N_66,In_749);
and U212 (N_212,In_283,In_126);
or U213 (N_213,In_311,In_250);
or U214 (N_214,In_412,N_110);
nand U215 (N_215,In_597,In_92);
xor U216 (N_216,In_663,In_62);
or U217 (N_217,N_135,N_104);
and U218 (N_218,In_569,N_111);
and U219 (N_219,N_103,In_155);
nand U220 (N_220,In_96,N_166);
nand U221 (N_221,N_165,In_45);
nand U222 (N_222,N_125,In_651);
nor U223 (N_223,In_362,N_47);
nand U224 (N_224,N_159,In_445);
nor U225 (N_225,N_186,In_4);
and U226 (N_226,N_199,In_128);
nor U227 (N_227,In_550,In_299);
nand U228 (N_228,N_34,In_505);
and U229 (N_229,In_479,N_171);
or U230 (N_230,N_180,In_163);
and U231 (N_231,In_285,N_76);
or U232 (N_232,N_120,In_203);
and U233 (N_233,In_42,In_237);
nor U234 (N_234,In_735,In_140);
and U235 (N_235,In_516,In_157);
nand U236 (N_236,In_691,N_146);
and U237 (N_237,In_575,In_490);
nand U238 (N_238,N_68,In_8);
or U239 (N_239,N_116,In_497);
and U240 (N_240,In_675,In_247);
nor U241 (N_241,In_382,In_268);
nand U242 (N_242,In_596,In_143);
nor U243 (N_243,In_733,N_131);
nand U244 (N_244,In_609,In_391);
nor U245 (N_245,N_191,In_438);
nor U246 (N_246,N_147,N_25);
nor U247 (N_247,In_94,In_626);
or U248 (N_248,N_20,In_292);
nor U249 (N_249,In_14,In_720);
and U250 (N_250,N_158,N_73);
or U251 (N_251,In_614,In_484);
and U252 (N_252,In_576,N_188);
and U253 (N_253,In_565,In_422);
and U254 (N_254,In_667,In_657);
nor U255 (N_255,N_44,In_643);
or U256 (N_256,In_91,N_33);
and U257 (N_257,In_197,In_69);
xor U258 (N_258,N_175,N_59);
or U259 (N_259,In_408,In_119);
nor U260 (N_260,In_682,In_286);
nor U261 (N_261,N_100,In_739);
nand U262 (N_262,In_613,In_70);
nand U263 (N_263,N_27,In_396);
or U264 (N_264,In_312,N_194);
xor U265 (N_265,N_13,In_132);
or U266 (N_266,In_55,N_148);
and U267 (N_267,In_344,In_725);
or U268 (N_268,N_144,N_31);
xnor U269 (N_269,In_607,In_624);
nor U270 (N_270,In_105,In_345);
nand U271 (N_271,In_31,In_538);
or U272 (N_272,In_80,N_106);
nor U273 (N_273,In_534,N_113);
or U274 (N_274,In_639,In_288);
or U275 (N_275,In_209,In_736);
nor U276 (N_276,In_628,N_6);
or U277 (N_277,In_731,In_317);
and U278 (N_278,In_627,N_161);
and U279 (N_279,N_70,In_656);
xor U280 (N_280,In_323,In_320);
nand U281 (N_281,In_79,In_340);
nand U282 (N_282,In_568,In_571);
nor U283 (N_283,In_34,In_158);
or U284 (N_284,In_619,N_195);
nor U285 (N_285,In_403,In_372);
nand U286 (N_286,N_193,N_168);
nor U287 (N_287,N_75,In_167);
and U288 (N_288,In_213,In_106);
xor U289 (N_289,In_421,In_293);
xnor U290 (N_290,N_124,N_81);
xnor U291 (N_291,N_52,N_101);
and U292 (N_292,N_130,In_46);
nor U293 (N_293,In_423,N_150);
or U294 (N_294,N_185,In_439);
nand U295 (N_295,In_592,N_86);
nand U296 (N_296,N_123,In_231);
and U297 (N_297,In_17,In_363);
nor U298 (N_298,In_267,N_89);
nand U299 (N_299,In_251,In_358);
nor U300 (N_300,N_259,N_289);
nor U301 (N_301,In_245,N_42);
xnor U302 (N_302,In_260,In_49);
nand U303 (N_303,N_154,N_18);
nor U304 (N_304,N_234,N_261);
nand U305 (N_305,In_446,N_255);
nor U306 (N_306,In_504,N_142);
or U307 (N_307,In_215,In_712);
or U308 (N_308,N_37,In_406);
nor U309 (N_309,In_620,In_75);
and U310 (N_310,In_590,N_201);
or U311 (N_311,N_24,In_638);
and U312 (N_312,In_615,In_348);
and U313 (N_313,In_552,N_200);
xnor U314 (N_314,N_215,In_357);
or U315 (N_315,N_272,In_144);
or U316 (N_316,N_243,N_267);
nand U317 (N_317,In_2,In_520);
nor U318 (N_318,In_246,In_546);
nor U319 (N_319,N_160,In_64);
nor U320 (N_320,In_700,In_3);
and U321 (N_321,In_523,In_205);
nor U322 (N_322,N_143,In_112);
nor U323 (N_323,In_118,In_744);
nand U324 (N_324,In_681,In_159);
nor U325 (N_325,N_88,N_241);
nor U326 (N_326,N_293,In_370);
and U327 (N_327,In_580,N_238);
nand U328 (N_328,In_279,N_246);
nor U329 (N_329,In_573,In_282);
nand U330 (N_330,N_253,In_532);
and U331 (N_331,In_717,N_213);
nand U332 (N_332,In_414,In_99);
or U333 (N_333,N_162,In_671);
or U334 (N_334,N_77,N_269);
nor U335 (N_335,In_579,In_61);
nand U336 (N_336,In_248,In_57);
and U337 (N_337,In_477,In_684);
and U338 (N_338,In_338,In_261);
nand U339 (N_339,N_211,N_63);
nor U340 (N_340,N_134,N_139);
or U341 (N_341,In_297,N_184);
nand U342 (N_342,N_71,In_435);
nor U343 (N_343,In_476,N_83);
or U344 (N_344,N_11,N_177);
nand U345 (N_345,N_126,In_97);
nor U346 (N_346,In_387,In_672);
xor U347 (N_347,In_632,N_245);
nor U348 (N_348,N_270,In_454);
nor U349 (N_349,In_257,In_217);
and U350 (N_350,N_90,N_108);
nor U351 (N_351,In_264,N_299);
nor U352 (N_352,In_687,In_734);
or U353 (N_353,In_152,In_393);
nor U354 (N_354,N_216,N_105);
and U355 (N_355,In_325,In_233);
and U356 (N_356,In_108,In_704);
nand U357 (N_357,In_7,In_500);
nor U358 (N_358,In_263,In_353);
or U359 (N_359,N_54,N_95);
and U360 (N_360,N_117,N_264);
nor U361 (N_361,N_223,In_719);
or U362 (N_362,N_15,N_1);
xor U363 (N_363,N_210,N_256);
nand U364 (N_364,N_179,N_254);
nand U365 (N_365,N_277,In_381);
or U366 (N_366,In_746,N_262);
nor U367 (N_367,In_271,In_424);
nor U368 (N_368,In_334,In_646);
and U369 (N_369,In_115,In_649);
nor U370 (N_370,In_270,In_541);
and U371 (N_371,In_0,N_132);
and U372 (N_372,In_26,In_73);
nor U373 (N_373,N_298,In_266);
and U374 (N_374,N_85,In_12);
and U375 (N_375,N_294,N_292);
nor U376 (N_376,In_662,In_563);
nor U377 (N_377,In_491,In_635);
and U378 (N_378,In_640,N_221);
nand U379 (N_379,In_478,N_244);
or U380 (N_380,N_172,N_115);
nor U381 (N_381,N_174,N_240);
or U382 (N_382,N_279,In_116);
nand U383 (N_383,In_560,In_74);
and U384 (N_384,N_35,N_297);
or U385 (N_385,In_226,In_359);
or U386 (N_386,N_258,In_707);
and U387 (N_387,N_141,In_525);
or U388 (N_388,N_217,N_64);
nor U389 (N_389,N_45,In_20);
or U390 (N_390,N_263,In_329);
nand U391 (N_391,In_350,N_296);
and U392 (N_392,In_536,In_308);
and U393 (N_393,In_680,N_65);
xor U394 (N_394,In_111,In_146);
and U395 (N_395,In_373,N_84);
nand U396 (N_396,N_251,In_33);
xor U397 (N_397,N_291,In_433);
nand U398 (N_398,N_260,N_230);
or U399 (N_399,In_318,In_361);
or U400 (N_400,N_281,In_648);
nand U401 (N_401,N_137,In_274);
nand U402 (N_402,In_208,N_338);
and U403 (N_403,N_344,N_359);
nor U404 (N_404,N_310,In_85);
nand U405 (N_405,N_396,In_558);
nand U406 (N_406,In_193,N_242);
nor U407 (N_407,In_319,N_271);
nor U408 (N_408,In_666,N_372);
nand U409 (N_409,N_214,In_722);
nor U410 (N_410,N_17,In_698);
or U411 (N_411,In_307,In_133);
and U412 (N_412,N_278,N_363);
nand U413 (N_413,N_324,N_364);
xor U414 (N_414,N_301,N_219);
and U415 (N_415,In_275,N_226);
nor U416 (N_416,N_358,N_74);
nand U417 (N_417,In_298,N_320);
or U418 (N_418,In_59,In_498);
xnor U419 (N_419,N_170,N_335);
or U420 (N_420,In_255,N_250);
nor U421 (N_421,In_127,N_21);
nand U422 (N_422,N_119,In_175);
or U423 (N_423,N_304,N_339);
nand U424 (N_424,In_499,In_343);
or U425 (N_425,In_517,N_373);
nor U426 (N_426,In_160,In_402);
nand U427 (N_427,N_391,N_375);
or U428 (N_428,In_404,In_341);
nand U429 (N_429,N_365,In_67);
or U430 (N_430,N_206,N_118);
nor U431 (N_431,N_196,In_36);
and U432 (N_432,N_284,N_381);
nor U433 (N_433,N_398,N_208);
xnor U434 (N_434,N_239,In_60);
or U435 (N_435,In_188,N_114);
or U436 (N_436,N_282,In_417);
nor U437 (N_437,N_376,In_300);
nor U438 (N_438,N_222,In_556);
nor U439 (N_439,N_212,N_312);
nor U440 (N_440,In_82,In_352);
nand U441 (N_441,N_341,N_163);
xnor U442 (N_442,In_104,N_93);
nand U443 (N_443,In_449,N_56);
or U444 (N_444,In_727,N_181);
and U445 (N_445,N_249,In_349);
nand U446 (N_446,N_280,N_315);
nor U447 (N_447,In_388,In_475);
and U448 (N_448,In_713,N_32);
nor U449 (N_449,In_174,N_39);
and U450 (N_450,N_287,N_390);
and U451 (N_451,In_474,In_544);
nand U452 (N_452,N_388,N_225);
or U453 (N_453,N_190,N_79);
nor U454 (N_454,N_368,N_155);
xnor U455 (N_455,N_343,N_169);
and U456 (N_456,In_471,N_205);
nand U457 (N_457,N_197,N_367);
nand U458 (N_458,N_99,In_486);
nor U459 (N_459,N_317,In_530);
and U460 (N_460,N_207,N_286);
nor U461 (N_461,N_360,N_347);
and U462 (N_462,N_354,N_257);
xor U463 (N_463,In_313,N_151);
and U464 (N_464,N_227,In_9);
nand U465 (N_465,N_112,In_131);
nand U466 (N_466,In_39,N_353);
and U467 (N_467,In_347,N_275);
nor U468 (N_468,N_349,In_380);
or U469 (N_469,N_164,In_216);
xor U470 (N_470,In_542,N_389);
or U471 (N_471,In_599,N_136);
or U472 (N_472,In_493,N_302);
and U473 (N_473,In_455,In_686);
nor U474 (N_474,N_129,N_247);
xor U475 (N_475,In_240,N_319);
or U476 (N_476,N_268,N_322);
nand U477 (N_477,N_321,In_239);
or U478 (N_478,In_374,In_706);
nor U479 (N_479,In_548,N_187);
or U480 (N_480,In_644,N_229);
and U481 (N_481,N_14,N_307);
and U482 (N_482,In_24,In_63);
and U483 (N_483,N_236,N_305);
nor U484 (N_484,In_461,N_366);
or U485 (N_485,In_401,N_128);
nand U486 (N_486,In_185,In_383);
nor U487 (N_487,In_557,N_386);
nor U488 (N_488,N_313,In_15);
nand U489 (N_489,N_274,In_389);
and U490 (N_490,In_444,In_398);
nand U491 (N_491,N_167,N_393);
nor U492 (N_492,In_230,N_232);
and U493 (N_493,In_332,N_345);
nand U494 (N_494,N_121,N_326);
and U495 (N_495,N_316,In_289);
nand U496 (N_496,N_102,In_90);
or U497 (N_497,N_276,N_380);
or U498 (N_498,In_485,N_290);
nand U499 (N_499,In_743,In_156);
xnor U500 (N_500,N_67,In_622);
nor U501 (N_501,N_189,N_336);
and U502 (N_502,N_401,N_416);
nand U503 (N_503,N_288,N_252);
nand U504 (N_504,N_369,N_228);
nand U505 (N_505,N_414,N_122);
and U506 (N_506,N_433,N_387);
or U507 (N_507,N_308,N_486);
nor U508 (N_508,N_340,N_443);
or U509 (N_509,N_404,N_346);
nor U510 (N_510,N_472,N_496);
or U511 (N_511,N_248,N_295);
nand U512 (N_512,N_394,N_487);
and U513 (N_513,N_464,In_276);
nand U514 (N_514,N_337,N_478);
or U515 (N_515,N_447,In_737);
and U516 (N_516,N_403,N_374);
or U517 (N_517,N_455,In_537);
or U518 (N_518,N_49,N_453);
and U519 (N_519,N_352,N_325);
nand U520 (N_520,N_451,N_456);
and U521 (N_521,N_98,N_471);
nor U522 (N_522,In_262,N_328);
xor U523 (N_523,N_427,N_384);
or U524 (N_524,N_371,N_311);
and U525 (N_525,In_1,N_418);
nor U526 (N_526,N_490,In_472);
nor U527 (N_527,In_588,N_484);
xnor U528 (N_528,N_458,N_399);
nor U529 (N_529,N_480,N_497);
nand U530 (N_530,N_475,N_421);
or U531 (N_531,N_385,N_273);
and U532 (N_532,N_430,N_468);
nand U533 (N_533,N_483,N_465);
and U534 (N_534,In_452,N_149);
nand U535 (N_535,N_309,In_315);
or U536 (N_536,N_356,N_449);
nand U537 (N_537,N_265,N_406);
or U538 (N_538,N_209,N_429);
xor U539 (N_539,N_362,In_272);
xnor U540 (N_540,N_314,N_29);
and U541 (N_541,N_419,N_0);
and U542 (N_542,In_342,In_172);
nand U543 (N_543,N_342,N_145);
xor U544 (N_544,N_470,N_329);
and U545 (N_545,N_400,In_608);
xnor U546 (N_546,N_378,In_611);
or U547 (N_547,N_395,N_474);
or U548 (N_548,N_424,In_430);
and U549 (N_549,N_382,N_351);
or U550 (N_550,N_204,In_400);
nor U551 (N_551,N_485,In_32);
nor U552 (N_552,N_40,N_495);
nand U553 (N_553,N_48,N_202);
nor U554 (N_554,In_480,N_420);
nand U555 (N_555,N_203,N_482);
nor U556 (N_556,N_231,N_409);
nand U557 (N_557,N_379,N_488);
nand U558 (N_558,In_335,N_334);
nand U559 (N_559,N_462,N_333);
xor U560 (N_560,N_370,In_301);
nand U561 (N_561,N_415,N_178);
or U562 (N_562,In_196,N_410);
nand U563 (N_563,N_361,N_153);
nor U564 (N_564,N_233,N_463);
and U565 (N_565,N_383,N_454);
nand U566 (N_566,N_457,N_36);
nand U567 (N_567,N_425,N_355);
nor U568 (N_568,In_642,N_411);
or U569 (N_569,N_436,N_498);
nand U570 (N_570,In_182,N_441);
xor U571 (N_571,N_392,N_138);
nand U572 (N_572,N_109,N_440);
nor U573 (N_573,N_467,N_331);
nand U574 (N_574,In_551,In_514);
nand U575 (N_575,N_422,N_432);
or U576 (N_576,N_450,In_730);
or U577 (N_577,In_464,N_53);
or U578 (N_578,N_489,In_177);
xnor U579 (N_579,N_459,N_152);
xor U580 (N_580,In_206,N_444);
or U581 (N_581,N_435,N_41);
and U582 (N_582,In_314,N_417);
and U583 (N_583,N_466,N_491);
and U584 (N_584,In_48,N_357);
or U585 (N_585,N_285,In_488);
nor U586 (N_586,N_224,N_442);
xnor U587 (N_587,N_266,N_439);
and U588 (N_588,In_634,N_348);
and U589 (N_589,N_452,N_460);
or U590 (N_590,In_407,N_446);
nor U591 (N_591,N_492,N_438);
nand U592 (N_592,N_183,In_365);
xor U593 (N_593,N_461,N_448);
or U594 (N_594,N_237,In_394);
nor U595 (N_595,N_173,N_494);
and U596 (N_596,N_350,N_235);
or U597 (N_597,In_227,N_493);
or U598 (N_598,N_377,In_561);
or U599 (N_599,N_477,In_482);
or U600 (N_600,N_557,N_531);
or U601 (N_601,N_511,N_575);
nand U602 (N_602,N_512,N_529);
and U603 (N_603,N_327,N_549);
nand U604 (N_604,N_514,N_407);
nand U605 (N_605,N_501,N_510);
nor U606 (N_606,N_587,N_551);
xor U607 (N_607,N_517,N_555);
nand U608 (N_608,N_506,N_537);
xor U609 (N_609,N_518,N_476);
nor U610 (N_610,N_573,N_569);
and U611 (N_611,N_220,N_445);
nor U612 (N_612,In_121,N_426);
nand U613 (N_613,N_554,N_198);
or U614 (N_614,N_543,In_95);
and U615 (N_615,N_568,N_541);
nand U616 (N_616,N_571,N_330);
nor U617 (N_617,N_520,N_157);
nor U618 (N_618,N_579,N_437);
and U619 (N_619,N_594,N_563);
nand U620 (N_620,N_597,N_559);
nand U621 (N_621,N_508,N_61);
nand U622 (N_622,N_397,N_522);
nor U623 (N_623,N_513,N_431);
nor U624 (N_624,N_576,N_499);
and U625 (N_625,N_519,N_332);
or U626 (N_626,N_552,N_402);
nor U627 (N_627,In_668,N_585);
and U628 (N_628,N_566,N_283);
or U629 (N_629,N_408,N_500);
xor U630 (N_630,N_534,N_524);
and U631 (N_631,N_581,N_525);
or U632 (N_632,N_300,N_323);
nor U633 (N_633,N_572,N_533);
nor U634 (N_634,N_405,N_218);
or U635 (N_635,N_509,N_538);
nor U636 (N_636,N_176,N_530);
or U637 (N_637,N_156,N_532);
nor U638 (N_638,N_526,In_399);
nor U639 (N_639,N_528,N_580);
nand U640 (N_640,N_596,N_428);
xnor U641 (N_641,N_521,N_107);
xor U642 (N_642,N_306,N_584);
xnor U643 (N_643,In_351,N_527);
nand U644 (N_644,N_413,N_507);
xor U645 (N_645,N_481,N_469);
nor U646 (N_646,N_505,N_598);
or U647 (N_647,N_565,N_590);
nand U648 (N_648,N_545,N_553);
and U649 (N_649,N_515,N_504);
and U650 (N_650,N_547,N_570);
nand U651 (N_651,N_578,N_539);
xor U652 (N_652,In_531,N_60);
and U653 (N_653,N_591,N_564);
or U654 (N_654,N_133,N_479);
or U655 (N_655,In_78,N_556);
or U656 (N_656,N_574,N_558);
or U657 (N_657,N_546,N_127);
or U658 (N_658,In_5,N_318);
or U659 (N_659,N_583,N_586);
xor U660 (N_660,N_550,N_599);
or U661 (N_661,N_562,N_542);
xor U662 (N_662,N_536,N_582);
and U663 (N_663,N_535,N_303);
or U664 (N_664,N_434,N_540);
and U665 (N_665,N_502,N_503);
or U666 (N_666,N_412,N_561);
and U667 (N_667,N_595,N_523);
and U668 (N_668,N_592,N_588);
xor U669 (N_669,N_516,N_589);
nand U670 (N_670,N_548,N_92);
or U671 (N_671,N_577,N_560);
or U672 (N_672,N_593,N_567);
nand U673 (N_673,N_544,N_473);
nor U674 (N_674,N_423,In_519);
and U675 (N_675,N_523,N_573);
and U676 (N_676,N_541,N_323);
nor U677 (N_677,N_569,N_428);
or U678 (N_678,In_668,N_589);
and U679 (N_679,N_306,In_519);
or U680 (N_680,N_585,N_303);
nor U681 (N_681,N_330,N_476);
nor U682 (N_682,N_596,N_593);
nor U683 (N_683,N_574,N_548);
xnor U684 (N_684,N_156,N_220);
nor U685 (N_685,N_517,N_542);
xor U686 (N_686,N_550,N_539);
or U687 (N_687,N_306,N_473);
nand U688 (N_688,N_547,N_157);
nor U689 (N_689,N_500,N_595);
xor U690 (N_690,N_590,N_542);
and U691 (N_691,N_547,N_553);
nand U692 (N_692,N_590,N_552);
and U693 (N_693,N_518,N_330);
nor U694 (N_694,N_586,N_332);
and U695 (N_695,N_598,N_589);
or U696 (N_696,N_540,N_593);
or U697 (N_697,N_426,N_573);
nand U698 (N_698,N_597,N_569);
or U699 (N_699,N_220,N_473);
or U700 (N_700,N_698,N_668);
nor U701 (N_701,N_680,N_623);
nor U702 (N_702,N_621,N_627);
or U703 (N_703,N_638,N_637);
nand U704 (N_704,N_641,N_662);
nor U705 (N_705,N_619,N_610);
or U706 (N_706,N_665,N_652);
or U707 (N_707,N_697,N_676);
and U708 (N_708,N_602,N_691);
nand U709 (N_709,N_689,N_673);
and U710 (N_710,N_626,N_695);
nand U711 (N_711,N_645,N_692);
or U712 (N_712,N_616,N_677);
and U713 (N_713,N_674,N_628);
nand U714 (N_714,N_622,N_669);
and U715 (N_715,N_681,N_661);
and U716 (N_716,N_694,N_603);
nand U717 (N_717,N_649,N_632);
nand U718 (N_718,N_671,N_686);
nand U719 (N_719,N_642,N_634);
nor U720 (N_720,N_651,N_685);
and U721 (N_721,N_664,N_653);
nor U722 (N_722,N_687,N_672);
and U723 (N_723,N_690,N_625);
and U724 (N_724,N_640,N_604);
and U725 (N_725,N_659,N_663);
or U726 (N_726,N_655,N_679);
or U727 (N_727,N_630,N_696);
and U728 (N_728,N_607,N_624);
and U729 (N_729,N_670,N_683);
nand U730 (N_730,N_629,N_639);
xnor U731 (N_731,N_678,N_620);
nand U732 (N_732,N_600,N_611);
and U733 (N_733,N_688,N_633);
xnor U734 (N_734,N_648,N_650);
nand U735 (N_735,N_654,N_618);
or U736 (N_736,N_646,N_615);
or U737 (N_737,N_660,N_656);
or U738 (N_738,N_635,N_601);
nand U739 (N_739,N_667,N_699);
or U740 (N_740,N_644,N_613);
xnor U741 (N_741,N_612,N_617);
nor U742 (N_742,N_631,N_675);
xor U743 (N_743,N_682,N_609);
or U744 (N_744,N_666,N_647);
and U745 (N_745,N_606,N_657);
nor U746 (N_746,N_605,N_643);
nor U747 (N_747,N_636,N_684);
nand U748 (N_748,N_614,N_608);
or U749 (N_749,N_658,N_693);
xnor U750 (N_750,N_630,N_622);
nand U751 (N_751,N_685,N_627);
nand U752 (N_752,N_657,N_615);
and U753 (N_753,N_688,N_670);
and U754 (N_754,N_662,N_604);
or U755 (N_755,N_663,N_615);
and U756 (N_756,N_602,N_600);
and U757 (N_757,N_640,N_689);
xor U758 (N_758,N_681,N_625);
nor U759 (N_759,N_678,N_666);
nand U760 (N_760,N_627,N_602);
nand U761 (N_761,N_659,N_680);
or U762 (N_762,N_681,N_616);
nor U763 (N_763,N_639,N_699);
nand U764 (N_764,N_688,N_655);
and U765 (N_765,N_688,N_663);
nor U766 (N_766,N_613,N_629);
or U767 (N_767,N_617,N_683);
and U768 (N_768,N_618,N_613);
and U769 (N_769,N_669,N_655);
nand U770 (N_770,N_659,N_621);
or U771 (N_771,N_656,N_624);
nor U772 (N_772,N_665,N_626);
nand U773 (N_773,N_694,N_689);
nand U774 (N_774,N_631,N_621);
and U775 (N_775,N_633,N_669);
and U776 (N_776,N_653,N_639);
nand U777 (N_777,N_643,N_636);
nor U778 (N_778,N_683,N_656);
and U779 (N_779,N_692,N_618);
or U780 (N_780,N_677,N_623);
xor U781 (N_781,N_673,N_610);
nand U782 (N_782,N_655,N_649);
nand U783 (N_783,N_686,N_667);
nand U784 (N_784,N_600,N_608);
xnor U785 (N_785,N_609,N_626);
or U786 (N_786,N_682,N_631);
and U787 (N_787,N_630,N_661);
nand U788 (N_788,N_617,N_607);
nand U789 (N_789,N_635,N_659);
nor U790 (N_790,N_672,N_618);
or U791 (N_791,N_664,N_666);
and U792 (N_792,N_632,N_653);
nand U793 (N_793,N_611,N_652);
or U794 (N_794,N_629,N_672);
or U795 (N_795,N_694,N_649);
xnor U796 (N_796,N_626,N_693);
xor U797 (N_797,N_663,N_674);
nand U798 (N_798,N_643,N_627);
nor U799 (N_799,N_697,N_616);
nand U800 (N_800,N_782,N_739);
and U801 (N_801,N_727,N_799);
or U802 (N_802,N_776,N_766);
or U803 (N_803,N_700,N_774);
xnor U804 (N_804,N_731,N_771);
xnor U805 (N_805,N_742,N_757);
nor U806 (N_806,N_747,N_710);
nand U807 (N_807,N_712,N_704);
nand U808 (N_808,N_795,N_706);
or U809 (N_809,N_773,N_767);
and U810 (N_810,N_755,N_707);
nand U811 (N_811,N_775,N_796);
and U812 (N_812,N_785,N_702);
or U813 (N_813,N_737,N_725);
nor U814 (N_814,N_728,N_736);
and U815 (N_815,N_759,N_703);
and U816 (N_816,N_715,N_792);
nor U817 (N_817,N_789,N_735);
or U818 (N_818,N_780,N_758);
nand U819 (N_819,N_754,N_717);
nand U820 (N_820,N_701,N_714);
and U821 (N_821,N_793,N_777);
and U822 (N_822,N_770,N_768);
xor U823 (N_823,N_720,N_779);
nand U824 (N_824,N_711,N_723);
and U825 (N_825,N_761,N_781);
nor U826 (N_826,N_778,N_751);
nand U827 (N_827,N_765,N_762);
and U828 (N_828,N_763,N_786);
xnor U829 (N_829,N_716,N_729);
and U830 (N_830,N_756,N_705);
and U831 (N_831,N_744,N_713);
and U832 (N_832,N_708,N_752);
or U833 (N_833,N_760,N_764);
nor U834 (N_834,N_722,N_790);
xnor U835 (N_835,N_746,N_797);
or U836 (N_836,N_718,N_769);
nand U837 (N_837,N_738,N_788);
and U838 (N_838,N_719,N_733);
nand U839 (N_839,N_753,N_787);
nor U840 (N_840,N_791,N_745);
xor U841 (N_841,N_741,N_794);
or U842 (N_842,N_721,N_709);
or U843 (N_843,N_783,N_730);
nor U844 (N_844,N_743,N_740);
nor U845 (N_845,N_784,N_724);
and U846 (N_846,N_749,N_772);
nor U847 (N_847,N_726,N_748);
nor U848 (N_848,N_734,N_750);
nand U849 (N_849,N_732,N_798);
or U850 (N_850,N_726,N_791);
and U851 (N_851,N_742,N_759);
xor U852 (N_852,N_779,N_714);
and U853 (N_853,N_794,N_739);
or U854 (N_854,N_744,N_778);
or U855 (N_855,N_721,N_775);
and U856 (N_856,N_764,N_743);
and U857 (N_857,N_771,N_770);
nand U858 (N_858,N_717,N_729);
or U859 (N_859,N_747,N_791);
nor U860 (N_860,N_795,N_709);
nand U861 (N_861,N_784,N_718);
and U862 (N_862,N_754,N_715);
and U863 (N_863,N_724,N_730);
or U864 (N_864,N_723,N_716);
or U865 (N_865,N_726,N_779);
xor U866 (N_866,N_747,N_713);
and U867 (N_867,N_714,N_798);
nor U868 (N_868,N_744,N_724);
nor U869 (N_869,N_795,N_707);
or U870 (N_870,N_704,N_713);
xor U871 (N_871,N_703,N_701);
xor U872 (N_872,N_710,N_748);
xor U873 (N_873,N_772,N_722);
nand U874 (N_874,N_798,N_766);
nand U875 (N_875,N_772,N_740);
or U876 (N_876,N_796,N_707);
xnor U877 (N_877,N_731,N_730);
and U878 (N_878,N_706,N_759);
and U879 (N_879,N_741,N_781);
xor U880 (N_880,N_743,N_737);
or U881 (N_881,N_717,N_796);
nor U882 (N_882,N_700,N_771);
and U883 (N_883,N_730,N_758);
xor U884 (N_884,N_789,N_772);
and U885 (N_885,N_790,N_746);
and U886 (N_886,N_707,N_769);
nand U887 (N_887,N_771,N_751);
and U888 (N_888,N_770,N_777);
nor U889 (N_889,N_704,N_755);
nand U890 (N_890,N_715,N_786);
nand U891 (N_891,N_765,N_759);
or U892 (N_892,N_729,N_758);
or U893 (N_893,N_750,N_793);
or U894 (N_894,N_720,N_718);
or U895 (N_895,N_730,N_744);
nand U896 (N_896,N_708,N_780);
nand U897 (N_897,N_719,N_709);
nand U898 (N_898,N_753,N_741);
and U899 (N_899,N_796,N_779);
xnor U900 (N_900,N_874,N_853);
xor U901 (N_901,N_883,N_801);
or U902 (N_902,N_881,N_845);
nand U903 (N_903,N_810,N_821);
nand U904 (N_904,N_829,N_807);
and U905 (N_905,N_855,N_843);
xnor U906 (N_906,N_865,N_866);
or U907 (N_907,N_806,N_889);
nand U908 (N_908,N_847,N_896);
nor U909 (N_909,N_891,N_879);
nor U910 (N_910,N_875,N_838);
and U911 (N_911,N_839,N_840);
nand U912 (N_912,N_846,N_886);
xnor U913 (N_913,N_814,N_805);
nor U914 (N_914,N_868,N_817);
xor U915 (N_915,N_898,N_870);
nand U916 (N_916,N_833,N_852);
and U917 (N_917,N_832,N_802);
nand U918 (N_918,N_861,N_835);
nor U919 (N_919,N_848,N_827);
or U920 (N_920,N_858,N_819);
or U921 (N_921,N_818,N_823);
or U922 (N_922,N_876,N_844);
and U923 (N_923,N_884,N_871);
nand U924 (N_924,N_893,N_841);
or U925 (N_925,N_815,N_820);
nand U926 (N_926,N_842,N_872);
nor U927 (N_927,N_860,N_863);
or U928 (N_928,N_878,N_811);
nor U929 (N_929,N_894,N_831);
nand U930 (N_930,N_825,N_800);
or U931 (N_931,N_895,N_824);
and U932 (N_932,N_887,N_864);
nor U933 (N_933,N_849,N_828);
nand U934 (N_934,N_897,N_822);
and U935 (N_935,N_851,N_834);
xor U936 (N_936,N_882,N_857);
nor U937 (N_937,N_826,N_830);
and U938 (N_938,N_812,N_873);
and U939 (N_939,N_862,N_836);
nand U940 (N_940,N_877,N_892);
xor U941 (N_941,N_816,N_837);
or U942 (N_942,N_899,N_890);
nor U943 (N_943,N_850,N_854);
nand U944 (N_944,N_888,N_869);
or U945 (N_945,N_880,N_859);
nand U946 (N_946,N_813,N_803);
or U947 (N_947,N_804,N_856);
or U948 (N_948,N_867,N_809);
xor U949 (N_949,N_808,N_885);
or U950 (N_950,N_834,N_861);
nor U951 (N_951,N_866,N_875);
xor U952 (N_952,N_802,N_833);
or U953 (N_953,N_820,N_842);
or U954 (N_954,N_899,N_896);
and U955 (N_955,N_822,N_877);
and U956 (N_956,N_879,N_876);
nor U957 (N_957,N_897,N_846);
or U958 (N_958,N_845,N_818);
nand U959 (N_959,N_883,N_848);
and U960 (N_960,N_825,N_841);
nand U961 (N_961,N_893,N_810);
nand U962 (N_962,N_890,N_837);
nand U963 (N_963,N_894,N_827);
xor U964 (N_964,N_868,N_848);
nor U965 (N_965,N_850,N_881);
nor U966 (N_966,N_875,N_830);
and U967 (N_967,N_821,N_897);
or U968 (N_968,N_851,N_871);
nor U969 (N_969,N_899,N_885);
nand U970 (N_970,N_861,N_862);
nor U971 (N_971,N_888,N_855);
xnor U972 (N_972,N_819,N_800);
and U973 (N_973,N_864,N_875);
nand U974 (N_974,N_849,N_872);
nor U975 (N_975,N_826,N_821);
and U976 (N_976,N_891,N_825);
nor U977 (N_977,N_839,N_883);
nor U978 (N_978,N_808,N_876);
xor U979 (N_979,N_851,N_892);
nor U980 (N_980,N_842,N_828);
or U981 (N_981,N_810,N_867);
or U982 (N_982,N_830,N_831);
or U983 (N_983,N_800,N_828);
xnor U984 (N_984,N_899,N_879);
xor U985 (N_985,N_821,N_869);
or U986 (N_986,N_855,N_853);
nand U987 (N_987,N_850,N_859);
nand U988 (N_988,N_865,N_826);
and U989 (N_989,N_801,N_821);
nor U990 (N_990,N_828,N_815);
and U991 (N_991,N_883,N_802);
and U992 (N_992,N_846,N_864);
or U993 (N_993,N_878,N_889);
nand U994 (N_994,N_825,N_867);
or U995 (N_995,N_832,N_880);
and U996 (N_996,N_823,N_816);
xor U997 (N_997,N_884,N_846);
nor U998 (N_998,N_866,N_858);
and U999 (N_999,N_898,N_897);
xor U1000 (N_1000,N_973,N_948);
and U1001 (N_1001,N_931,N_992);
or U1002 (N_1002,N_953,N_943);
xor U1003 (N_1003,N_926,N_945);
nor U1004 (N_1004,N_937,N_905);
nand U1005 (N_1005,N_923,N_969);
nor U1006 (N_1006,N_985,N_910);
or U1007 (N_1007,N_947,N_990);
nand U1008 (N_1008,N_934,N_986);
and U1009 (N_1009,N_959,N_968);
or U1010 (N_1010,N_979,N_960);
nor U1011 (N_1011,N_976,N_994);
or U1012 (N_1012,N_942,N_932);
nor U1013 (N_1013,N_956,N_927);
nor U1014 (N_1014,N_950,N_970);
nor U1015 (N_1015,N_925,N_929);
nand U1016 (N_1016,N_966,N_964);
nand U1017 (N_1017,N_919,N_902);
and U1018 (N_1018,N_961,N_982);
or U1019 (N_1019,N_944,N_922);
and U1020 (N_1020,N_998,N_967);
nor U1021 (N_1021,N_921,N_984);
or U1022 (N_1022,N_916,N_997);
nor U1023 (N_1023,N_935,N_940);
and U1024 (N_1024,N_955,N_981);
nand U1025 (N_1025,N_908,N_988);
nand U1026 (N_1026,N_999,N_924);
and U1027 (N_1027,N_907,N_954);
and U1028 (N_1028,N_977,N_901);
or U1029 (N_1029,N_978,N_989);
or U1030 (N_1030,N_951,N_996);
nor U1031 (N_1031,N_941,N_906);
nand U1032 (N_1032,N_938,N_913);
nand U1033 (N_1033,N_920,N_958);
or U1034 (N_1034,N_930,N_914);
xnor U1035 (N_1035,N_900,N_946);
nand U1036 (N_1036,N_991,N_962);
and U1037 (N_1037,N_971,N_912);
and U1038 (N_1038,N_918,N_975);
or U1039 (N_1039,N_995,N_933);
and U1040 (N_1040,N_957,N_917);
or U1041 (N_1041,N_972,N_909);
and U1042 (N_1042,N_911,N_949);
nor U1043 (N_1043,N_903,N_980);
nand U1044 (N_1044,N_952,N_993);
nor U1045 (N_1045,N_983,N_939);
nor U1046 (N_1046,N_974,N_936);
or U1047 (N_1047,N_965,N_963);
nand U1048 (N_1048,N_904,N_987);
nor U1049 (N_1049,N_928,N_915);
xor U1050 (N_1050,N_975,N_923);
nand U1051 (N_1051,N_996,N_981);
and U1052 (N_1052,N_958,N_971);
nor U1053 (N_1053,N_926,N_967);
nand U1054 (N_1054,N_900,N_904);
and U1055 (N_1055,N_924,N_971);
or U1056 (N_1056,N_988,N_957);
or U1057 (N_1057,N_942,N_930);
or U1058 (N_1058,N_959,N_955);
xor U1059 (N_1059,N_969,N_978);
xnor U1060 (N_1060,N_973,N_901);
or U1061 (N_1061,N_966,N_949);
nand U1062 (N_1062,N_953,N_937);
and U1063 (N_1063,N_938,N_949);
xor U1064 (N_1064,N_972,N_966);
and U1065 (N_1065,N_935,N_915);
or U1066 (N_1066,N_977,N_974);
or U1067 (N_1067,N_924,N_976);
nor U1068 (N_1068,N_979,N_906);
or U1069 (N_1069,N_920,N_962);
xor U1070 (N_1070,N_975,N_920);
and U1071 (N_1071,N_999,N_903);
nor U1072 (N_1072,N_930,N_923);
and U1073 (N_1073,N_906,N_996);
xor U1074 (N_1074,N_917,N_932);
nand U1075 (N_1075,N_970,N_939);
and U1076 (N_1076,N_924,N_981);
nor U1077 (N_1077,N_906,N_911);
or U1078 (N_1078,N_919,N_964);
nand U1079 (N_1079,N_901,N_966);
nor U1080 (N_1080,N_958,N_981);
nand U1081 (N_1081,N_989,N_975);
and U1082 (N_1082,N_981,N_922);
or U1083 (N_1083,N_902,N_905);
or U1084 (N_1084,N_971,N_902);
or U1085 (N_1085,N_946,N_983);
or U1086 (N_1086,N_992,N_974);
or U1087 (N_1087,N_935,N_967);
nor U1088 (N_1088,N_989,N_966);
nand U1089 (N_1089,N_916,N_949);
or U1090 (N_1090,N_958,N_964);
or U1091 (N_1091,N_960,N_990);
nand U1092 (N_1092,N_925,N_933);
and U1093 (N_1093,N_953,N_923);
and U1094 (N_1094,N_924,N_933);
nor U1095 (N_1095,N_966,N_959);
nor U1096 (N_1096,N_914,N_907);
nor U1097 (N_1097,N_918,N_916);
and U1098 (N_1098,N_998,N_909);
or U1099 (N_1099,N_928,N_939);
nor U1100 (N_1100,N_1077,N_1098);
nand U1101 (N_1101,N_1049,N_1018);
or U1102 (N_1102,N_1030,N_1053);
nand U1103 (N_1103,N_1013,N_1086);
and U1104 (N_1104,N_1055,N_1029);
nor U1105 (N_1105,N_1062,N_1044);
xnor U1106 (N_1106,N_1069,N_1000);
nor U1107 (N_1107,N_1009,N_1073);
or U1108 (N_1108,N_1076,N_1089);
and U1109 (N_1109,N_1008,N_1001);
or U1110 (N_1110,N_1088,N_1033);
xor U1111 (N_1111,N_1046,N_1068);
nor U1112 (N_1112,N_1094,N_1003);
nand U1113 (N_1113,N_1012,N_1056);
nand U1114 (N_1114,N_1064,N_1063);
nor U1115 (N_1115,N_1005,N_1083);
or U1116 (N_1116,N_1092,N_1078);
and U1117 (N_1117,N_1075,N_1011);
nand U1118 (N_1118,N_1043,N_1097);
or U1119 (N_1119,N_1093,N_1079);
nor U1120 (N_1120,N_1084,N_1010);
nor U1121 (N_1121,N_1061,N_1042);
and U1122 (N_1122,N_1047,N_1025);
and U1123 (N_1123,N_1067,N_1020);
nor U1124 (N_1124,N_1090,N_1087);
or U1125 (N_1125,N_1037,N_1080);
or U1126 (N_1126,N_1026,N_1032);
nor U1127 (N_1127,N_1028,N_1041);
xor U1128 (N_1128,N_1006,N_1021);
xor U1129 (N_1129,N_1082,N_1022);
and U1130 (N_1130,N_1052,N_1081);
xnor U1131 (N_1131,N_1024,N_1015);
nor U1132 (N_1132,N_1027,N_1002);
xnor U1133 (N_1133,N_1031,N_1036);
and U1134 (N_1134,N_1059,N_1014);
or U1135 (N_1135,N_1071,N_1016);
nor U1136 (N_1136,N_1054,N_1038);
nand U1137 (N_1137,N_1096,N_1039);
nor U1138 (N_1138,N_1070,N_1099);
and U1139 (N_1139,N_1060,N_1004);
nor U1140 (N_1140,N_1035,N_1034);
nor U1141 (N_1141,N_1095,N_1085);
or U1142 (N_1142,N_1065,N_1058);
or U1143 (N_1143,N_1048,N_1050);
or U1144 (N_1144,N_1045,N_1023);
or U1145 (N_1145,N_1019,N_1051);
nand U1146 (N_1146,N_1017,N_1072);
and U1147 (N_1147,N_1066,N_1074);
xor U1148 (N_1148,N_1091,N_1007);
nor U1149 (N_1149,N_1040,N_1057);
nor U1150 (N_1150,N_1010,N_1011);
or U1151 (N_1151,N_1075,N_1038);
or U1152 (N_1152,N_1029,N_1067);
or U1153 (N_1153,N_1093,N_1073);
or U1154 (N_1154,N_1008,N_1069);
or U1155 (N_1155,N_1031,N_1011);
nor U1156 (N_1156,N_1082,N_1087);
and U1157 (N_1157,N_1064,N_1023);
and U1158 (N_1158,N_1080,N_1073);
or U1159 (N_1159,N_1094,N_1045);
nand U1160 (N_1160,N_1028,N_1034);
nand U1161 (N_1161,N_1077,N_1073);
xnor U1162 (N_1162,N_1038,N_1030);
nand U1163 (N_1163,N_1051,N_1009);
nor U1164 (N_1164,N_1008,N_1006);
nand U1165 (N_1165,N_1012,N_1044);
or U1166 (N_1166,N_1053,N_1005);
nand U1167 (N_1167,N_1013,N_1076);
and U1168 (N_1168,N_1008,N_1039);
nand U1169 (N_1169,N_1079,N_1075);
xnor U1170 (N_1170,N_1057,N_1096);
nand U1171 (N_1171,N_1063,N_1040);
and U1172 (N_1172,N_1063,N_1046);
or U1173 (N_1173,N_1004,N_1064);
nand U1174 (N_1174,N_1068,N_1037);
nand U1175 (N_1175,N_1098,N_1002);
or U1176 (N_1176,N_1080,N_1065);
or U1177 (N_1177,N_1076,N_1001);
xor U1178 (N_1178,N_1025,N_1019);
or U1179 (N_1179,N_1049,N_1092);
nand U1180 (N_1180,N_1078,N_1090);
nor U1181 (N_1181,N_1055,N_1070);
or U1182 (N_1182,N_1042,N_1083);
and U1183 (N_1183,N_1079,N_1077);
or U1184 (N_1184,N_1014,N_1043);
or U1185 (N_1185,N_1095,N_1064);
nand U1186 (N_1186,N_1095,N_1065);
nor U1187 (N_1187,N_1096,N_1087);
nor U1188 (N_1188,N_1022,N_1064);
or U1189 (N_1189,N_1039,N_1061);
and U1190 (N_1190,N_1075,N_1058);
or U1191 (N_1191,N_1006,N_1003);
and U1192 (N_1192,N_1005,N_1004);
and U1193 (N_1193,N_1046,N_1009);
nor U1194 (N_1194,N_1051,N_1024);
or U1195 (N_1195,N_1077,N_1016);
or U1196 (N_1196,N_1088,N_1000);
or U1197 (N_1197,N_1072,N_1033);
and U1198 (N_1198,N_1090,N_1024);
xor U1199 (N_1199,N_1066,N_1024);
nor U1200 (N_1200,N_1162,N_1101);
nor U1201 (N_1201,N_1194,N_1135);
xnor U1202 (N_1202,N_1145,N_1105);
and U1203 (N_1203,N_1148,N_1147);
nand U1204 (N_1204,N_1130,N_1168);
or U1205 (N_1205,N_1138,N_1131);
nor U1206 (N_1206,N_1142,N_1174);
nand U1207 (N_1207,N_1104,N_1160);
and U1208 (N_1208,N_1173,N_1134);
or U1209 (N_1209,N_1163,N_1136);
or U1210 (N_1210,N_1182,N_1124);
nand U1211 (N_1211,N_1180,N_1156);
nor U1212 (N_1212,N_1157,N_1115);
and U1213 (N_1213,N_1140,N_1141);
or U1214 (N_1214,N_1166,N_1189);
and U1215 (N_1215,N_1170,N_1144);
or U1216 (N_1216,N_1190,N_1165);
nand U1217 (N_1217,N_1196,N_1195);
xnor U1218 (N_1218,N_1127,N_1113);
xor U1219 (N_1219,N_1126,N_1133);
or U1220 (N_1220,N_1129,N_1164);
nand U1221 (N_1221,N_1161,N_1178);
or U1222 (N_1222,N_1171,N_1150);
nand U1223 (N_1223,N_1146,N_1177);
and U1224 (N_1224,N_1151,N_1192);
or U1225 (N_1225,N_1188,N_1159);
or U1226 (N_1226,N_1181,N_1110);
nand U1227 (N_1227,N_1155,N_1118);
or U1228 (N_1228,N_1186,N_1154);
or U1229 (N_1229,N_1100,N_1187);
xnor U1230 (N_1230,N_1132,N_1122);
and U1231 (N_1231,N_1102,N_1193);
nor U1232 (N_1232,N_1108,N_1114);
nand U1233 (N_1233,N_1125,N_1152);
or U1234 (N_1234,N_1153,N_1175);
and U1235 (N_1235,N_1112,N_1169);
nand U1236 (N_1236,N_1103,N_1167);
and U1237 (N_1237,N_1185,N_1143);
and U1238 (N_1238,N_1107,N_1121);
or U1239 (N_1239,N_1117,N_1128);
nand U1240 (N_1240,N_1109,N_1199);
or U1241 (N_1241,N_1119,N_1176);
and U1242 (N_1242,N_1179,N_1137);
nand U1243 (N_1243,N_1158,N_1139);
nor U1244 (N_1244,N_1149,N_1120);
nor U1245 (N_1245,N_1184,N_1198);
or U1246 (N_1246,N_1183,N_1172);
nand U1247 (N_1247,N_1123,N_1197);
nand U1248 (N_1248,N_1191,N_1116);
nand U1249 (N_1249,N_1111,N_1106);
and U1250 (N_1250,N_1186,N_1196);
nor U1251 (N_1251,N_1177,N_1105);
nor U1252 (N_1252,N_1101,N_1158);
or U1253 (N_1253,N_1143,N_1184);
nand U1254 (N_1254,N_1119,N_1138);
nand U1255 (N_1255,N_1139,N_1181);
nand U1256 (N_1256,N_1121,N_1120);
xnor U1257 (N_1257,N_1147,N_1197);
xnor U1258 (N_1258,N_1190,N_1157);
or U1259 (N_1259,N_1104,N_1165);
or U1260 (N_1260,N_1109,N_1182);
or U1261 (N_1261,N_1185,N_1157);
or U1262 (N_1262,N_1107,N_1132);
and U1263 (N_1263,N_1114,N_1160);
nor U1264 (N_1264,N_1161,N_1173);
nand U1265 (N_1265,N_1151,N_1186);
nor U1266 (N_1266,N_1196,N_1183);
and U1267 (N_1267,N_1181,N_1104);
nand U1268 (N_1268,N_1168,N_1186);
or U1269 (N_1269,N_1193,N_1140);
xnor U1270 (N_1270,N_1154,N_1103);
or U1271 (N_1271,N_1158,N_1121);
and U1272 (N_1272,N_1144,N_1125);
nor U1273 (N_1273,N_1105,N_1191);
and U1274 (N_1274,N_1112,N_1103);
or U1275 (N_1275,N_1181,N_1191);
or U1276 (N_1276,N_1196,N_1110);
xnor U1277 (N_1277,N_1125,N_1122);
and U1278 (N_1278,N_1199,N_1122);
xnor U1279 (N_1279,N_1187,N_1177);
or U1280 (N_1280,N_1159,N_1168);
nand U1281 (N_1281,N_1118,N_1177);
nor U1282 (N_1282,N_1109,N_1131);
nand U1283 (N_1283,N_1191,N_1174);
and U1284 (N_1284,N_1181,N_1165);
and U1285 (N_1285,N_1195,N_1108);
xor U1286 (N_1286,N_1141,N_1100);
nor U1287 (N_1287,N_1194,N_1158);
nor U1288 (N_1288,N_1190,N_1100);
or U1289 (N_1289,N_1173,N_1103);
nand U1290 (N_1290,N_1112,N_1153);
nand U1291 (N_1291,N_1177,N_1195);
nor U1292 (N_1292,N_1109,N_1105);
nand U1293 (N_1293,N_1101,N_1116);
nor U1294 (N_1294,N_1160,N_1152);
and U1295 (N_1295,N_1193,N_1105);
nand U1296 (N_1296,N_1154,N_1177);
and U1297 (N_1297,N_1197,N_1102);
nor U1298 (N_1298,N_1139,N_1178);
or U1299 (N_1299,N_1137,N_1174);
nand U1300 (N_1300,N_1247,N_1279);
and U1301 (N_1301,N_1270,N_1232);
nor U1302 (N_1302,N_1215,N_1269);
nand U1303 (N_1303,N_1231,N_1242);
nand U1304 (N_1304,N_1237,N_1236);
or U1305 (N_1305,N_1210,N_1213);
or U1306 (N_1306,N_1244,N_1264);
nand U1307 (N_1307,N_1201,N_1278);
and U1308 (N_1308,N_1297,N_1295);
nand U1309 (N_1309,N_1274,N_1263);
or U1310 (N_1310,N_1235,N_1257);
nand U1311 (N_1311,N_1207,N_1285);
and U1312 (N_1312,N_1256,N_1293);
nand U1313 (N_1313,N_1220,N_1251);
xor U1314 (N_1314,N_1248,N_1240);
and U1315 (N_1315,N_1281,N_1292);
nand U1316 (N_1316,N_1202,N_1284);
nor U1317 (N_1317,N_1252,N_1280);
xor U1318 (N_1318,N_1294,N_1260);
nand U1319 (N_1319,N_1226,N_1277);
xor U1320 (N_1320,N_1271,N_1209);
or U1321 (N_1321,N_1298,N_1299);
or U1322 (N_1322,N_1223,N_1286);
and U1323 (N_1323,N_1203,N_1262);
nand U1324 (N_1324,N_1204,N_1261);
nand U1325 (N_1325,N_1239,N_1214);
and U1326 (N_1326,N_1249,N_1216);
nor U1327 (N_1327,N_1291,N_1208);
or U1328 (N_1328,N_1206,N_1217);
nand U1329 (N_1329,N_1221,N_1289);
nand U1330 (N_1330,N_1265,N_1224);
nor U1331 (N_1331,N_1282,N_1211);
nor U1332 (N_1332,N_1222,N_1266);
xor U1333 (N_1333,N_1267,N_1233);
nor U1334 (N_1334,N_1219,N_1246);
nor U1335 (N_1335,N_1200,N_1228);
nor U1336 (N_1336,N_1268,N_1283);
nand U1337 (N_1337,N_1245,N_1212);
and U1338 (N_1338,N_1288,N_1275);
nor U1339 (N_1339,N_1205,N_1276);
nand U1340 (N_1340,N_1287,N_1255);
nor U1341 (N_1341,N_1250,N_1259);
nor U1342 (N_1342,N_1241,N_1238);
or U1343 (N_1343,N_1227,N_1234);
nor U1344 (N_1344,N_1258,N_1225);
or U1345 (N_1345,N_1254,N_1230);
nor U1346 (N_1346,N_1218,N_1272);
or U1347 (N_1347,N_1253,N_1290);
nor U1348 (N_1348,N_1296,N_1243);
nor U1349 (N_1349,N_1229,N_1273);
nand U1350 (N_1350,N_1265,N_1292);
nand U1351 (N_1351,N_1271,N_1211);
xnor U1352 (N_1352,N_1258,N_1218);
nor U1353 (N_1353,N_1249,N_1264);
and U1354 (N_1354,N_1210,N_1231);
or U1355 (N_1355,N_1286,N_1248);
or U1356 (N_1356,N_1286,N_1219);
and U1357 (N_1357,N_1268,N_1223);
or U1358 (N_1358,N_1239,N_1275);
nor U1359 (N_1359,N_1202,N_1228);
nand U1360 (N_1360,N_1273,N_1212);
or U1361 (N_1361,N_1261,N_1242);
and U1362 (N_1362,N_1244,N_1272);
and U1363 (N_1363,N_1217,N_1248);
xnor U1364 (N_1364,N_1251,N_1244);
nor U1365 (N_1365,N_1290,N_1248);
or U1366 (N_1366,N_1260,N_1293);
nor U1367 (N_1367,N_1238,N_1293);
nand U1368 (N_1368,N_1272,N_1234);
and U1369 (N_1369,N_1274,N_1271);
or U1370 (N_1370,N_1249,N_1257);
nand U1371 (N_1371,N_1254,N_1286);
nor U1372 (N_1372,N_1260,N_1235);
and U1373 (N_1373,N_1241,N_1215);
and U1374 (N_1374,N_1259,N_1254);
or U1375 (N_1375,N_1298,N_1289);
nor U1376 (N_1376,N_1232,N_1227);
or U1377 (N_1377,N_1293,N_1244);
and U1378 (N_1378,N_1271,N_1281);
or U1379 (N_1379,N_1286,N_1289);
nand U1380 (N_1380,N_1252,N_1269);
nand U1381 (N_1381,N_1238,N_1236);
nand U1382 (N_1382,N_1251,N_1227);
nand U1383 (N_1383,N_1259,N_1275);
and U1384 (N_1384,N_1217,N_1241);
nand U1385 (N_1385,N_1208,N_1210);
nand U1386 (N_1386,N_1256,N_1286);
and U1387 (N_1387,N_1258,N_1290);
and U1388 (N_1388,N_1260,N_1273);
xnor U1389 (N_1389,N_1261,N_1200);
and U1390 (N_1390,N_1284,N_1238);
nor U1391 (N_1391,N_1204,N_1278);
and U1392 (N_1392,N_1231,N_1291);
nor U1393 (N_1393,N_1286,N_1236);
and U1394 (N_1394,N_1288,N_1277);
nor U1395 (N_1395,N_1268,N_1202);
nor U1396 (N_1396,N_1213,N_1293);
or U1397 (N_1397,N_1240,N_1275);
nor U1398 (N_1398,N_1287,N_1230);
nor U1399 (N_1399,N_1204,N_1263);
or U1400 (N_1400,N_1351,N_1399);
xor U1401 (N_1401,N_1395,N_1367);
nor U1402 (N_1402,N_1356,N_1326);
or U1403 (N_1403,N_1323,N_1378);
nor U1404 (N_1404,N_1305,N_1353);
and U1405 (N_1405,N_1372,N_1324);
xor U1406 (N_1406,N_1388,N_1334);
or U1407 (N_1407,N_1359,N_1315);
nor U1408 (N_1408,N_1343,N_1379);
and U1409 (N_1409,N_1374,N_1339);
xnor U1410 (N_1410,N_1308,N_1341);
xor U1411 (N_1411,N_1380,N_1390);
nor U1412 (N_1412,N_1376,N_1369);
or U1413 (N_1413,N_1358,N_1333);
and U1414 (N_1414,N_1396,N_1300);
and U1415 (N_1415,N_1342,N_1301);
and U1416 (N_1416,N_1383,N_1364);
nor U1417 (N_1417,N_1311,N_1318);
and U1418 (N_1418,N_1313,N_1349);
nor U1419 (N_1419,N_1352,N_1316);
and U1420 (N_1420,N_1354,N_1350);
and U1421 (N_1421,N_1363,N_1309);
and U1422 (N_1422,N_1303,N_1377);
xor U1423 (N_1423,N_1393,N_1307);
nor U1424 (N_1424,N_1332,N_1361);
or U1425 (N_1425,N_1346,N_1306);
nand U1426 (N_1426,N_1362,N_1373);
and U1427 (N_1427,N_1344,N_1389);
nor U1428 (N_1428,N_1391,N_1381);
nor U1429 (N_1429,N_1366,N_1328);
nand U1430 (N_1430,N_1304,N_1394);
and U1431 (N_1431,N_1321,N_1325);
and U1432 (N_1432,N_1330,N_1317);
or U1433 (N_1433,N_1302,N_1368);
or U1434 (N_1434,N_1331,N_1329);
xor U1435 (N_1435,N_1337,N_1370);
and U1436 (N_1436,N_1398,N_1320);
nor U1437 (N_1437,N_1347,N_1386);
nand U1438 (N_1438,N_1336,N_1348);
nand U1439 (N_1439,N_1371,N_1310);
or U1440 (N_1440,N_1314,N_1365);
nand U1441 (N_1441,N_1340,N_1355);
nor U1442 (N_1442,N_1382,N_1335);
or U1443 (N_1443,N_1360,N_1385);
and U1444 (N_1444,N_1357,N_1387);
xor U1445 (N_1445,N_1375,N_1384);
xnor U1446 (N_1446,N_1392,N_1327);
and U1447 (N_1447,N_1322,N_1319);
or U1448 (N_1448,N_1338,N_1345);
or U1449 (N_1449,N_1312,N_1397);
and U1450 (N_1450,N_1386,N_1373);
nor U1451 (N_1451,N_1335,N_1340);
nand U1452 (N_1452,N_1325,N_1389);
nand U1453 (N_1453,N_1309,N_1391);
or U1454 (N_1454,N_1379,N_1329);
or U1455 (N_1455,N_1387,N_1368);
nor U1456 (N_1456,N_1316,N_1347);
or U1457 (N_1457,N_1328,N_1324);
and U1458 (N_1458,N_1327,N_1319);
xnor U1459 (N_1459,N_1323,N_1329);
or U1460 (N_1460,N_1344,N_1354);
xnor U1461 (N_1461,N_1344,N_1321);
and U1462 (N_1462,N_1303,N_1327);
and U1463 (N_1463,N_1346,N_1319);
nand U1464 (N_1464,N_1316,N_1330);
and U1465 (N_1465,N_1329,N_1312);
nand U1466 (N_1466,N_1378,N_1341);
nor U1467 (N_1467,N_1349,N_1399);
or U1468 (N_1468,N_1304,N_1361);
nor U1469 (N_1469,N_1389,N_1303);
nor U1470 (N_1470,N_1344,N_1379);
and U1471 (N_1471,N_1301,N_1349);
xor U1472 (N_1472,N_1348,N_1309);
nor U1473 (N_1473,N_1320,N_1347);
or U1474 (N_1474,N_1304,N_1357);
or U1475 (N_1475,N_1372,N_1370);
nor U1476 (N_1476,N_1347,N_1356);
or U1477 (N_1477,N_1388,N_1393);
nor U1478 (N_1478,N_1313,N_1348);
or U1479 (N_1479,N_1369,N_1399);
and U1480 (N_1480,N_1372,N_1338);
and U1481 (N_1481,N_1362,N_1340);
or U1482 (N_1482,N_1399,N_1389);
or U1483 (N_1483,N_1379,N_1335);
or U1484 (N_1484,N_1364,N_1387);
and U1485 (N_1485,N_1382,N_1378);
nand U1486 (N_1486,N_1395,N_1387);
or U1487 (N_1487,N_1363,N_1393);
and U1488 (N_1488,N_1339,N_1372);
nand U1489 (N_1489,N_1366,N_1347);
xor U1490 (N_1490,N_1395,N_1307);
nor U1491 (N_1491,N_1319,N_1334);
nand U1492 (N_1492,N_1306,N_1387);
nor U1493 (N_1493,N_1364,N_1313);
or U1494 (N_1494,N_1396,N_1324);
and U1495 (N_1495,N_1358,N_1372);
or U1496 (N_1496,N_1332,N_1382);
xnor U1497 (N_1497,N_1313,N_1355);
nor U1498 (N_1498,N_1365,N_1312);
nor U1499 (N_1499,N_1321,N_1307);
and U1500 (N_1500,N_1465,N_1484);
or U1501 (N_1501,N_1488,N_1448);
nand U1502 (N_1502,N_1443,N_1441);
nand U1503 (N_1503,N_1473,N_1466);
nor U1504 (N_1504,N_1485,N_1474);
and U1505 (N_1505,N_1453,N_1478);
nand U1506 (N_1506,N_1475,N_1497);
or U1507 (N_1507,N_1444,N_1409);
nor U1508 (N_1508,N_1400,N_1463);
xnor U1509 (N_1509,N_1417,N_1467);
or U1510 (N_1510,N_1471,N_1487);
nand U1511 (N_1511,N_1480,N_1472);
and U1512 (N_1512,N_1437,N_1438);
nand U1513 (N_1513,N_1459,N_1406);
and U1514 (N_1514,N_1434,N_1495);
and U1515 (N_1515,N_1486,N_1412);
nand U1516 (N_1516,N_1482,N_1470);
nand U1517 (N_1517,N_1489,N_1425);
nor U1518 (N_1518,N_1429,N_1469);
nand U1519 (N_1519,N_1450,N_1419);
or U1520 (N_1520,N_1423,N_1454);
and U1521 (N_1521,N_1492,N_1447);
and U1522 (N_1522,N_1408,N_1462);
nor U1523 (N_1523,N_1430,N_1439);
or U1524 (N_1524,N_1479,N_1410);
and U1525 (N_1525,N_1494,N_1402);
or U1526 (N_1526,N_1498,N_1407);
nor U1527 (N_1527,N_1493,N_1420);
or U1528 (N_1528,N_1416,N_1458);
or U1529 (N_1529,N_1426,N_1477);
and U1530 (N_1530,N_1491,N_1413);
nand U1531 (N_1531,N_1440,N_1455);
nand U1532 (N_1532,N_1411,N_1405);
nor U1533 (N_1533,N_1457,N_1452);
nor U1534 (N_1534,N_1403,N_1435);
nand U1535 (N_1535,N_1456,N_1481);
or U1536 (N_1536,N_1421,N_1401);
or U1537 (N_1537,N_1424,N_1418);
xnor U1538 (N_1538,N_1464,N_1460);
and U1539 (N_1539,N_1422,N_1436);
or U1540 (N_1540,N_1449,N_1451);
nor U1541 (N_1541,N_1490,N_1404);
nand U1542 (N_1542,N_1483,N_1432);
nor U1543 (N_1543,N_1445,N_1415);
nor U1544 (N_1544,N_1442,N_1499);
nand U1545 (N_1545,N_1428,N_1414);
and U1546 (N_1546,N_1446,N_1433);
and U1547 (N_1547,N_1496,N_1427);
or U1548 (N_1548,N_1468,N_1476);
and U1549 (N_1549,N_1461,N_1431);
and U1550 (N_1550,N_1428,N_1487);
nor U1551 (N_1551,N_1419,N_1437);
or U1552 (N_1552,N_1447,N_1445);
and U1553 (N_1553,N_1458,N_1440);
and U1554 (N_1554,N_1413,N_1400);
and U1555 (N_1555,N_1492,N_1458);
or U1556 (N_1556,N_1458,N_1435);
and U1557 (N_1557,N_1454,N_1424);
xnor U1558 (N_1558,N_1440,N_1410);
xor U1559 (N_1559,N_1441,N_1400);
nand U1560 (N_1560,N_1439,N_1403);
nand U1561 (N_1561,N_1423,N_1474);
nand U1562 (N_1562,N_1422,N_1465);
or U1563 (N_1563,N_1423,N_1495);
nand U1564 (N_1564,N_1431,N_1420);
and U1565 (N_1565,N_1479,N_1432);
nor U1566 (N_1566,N_1462,N_1426);
nand U1567 (N_1567,N_1423,N_1401);
nand U1568 (N_1568,N_1491,N_1430);
and U1569 (N_1569,N_1457,N_1498);
nor U1570 (N_1570,N_1406,N_1402);
nor U1571 (N_1571,N_1494,N_1434);
or U1572 (N_1572,N_1431,N_1415);
nand U1573 (N_1573,N_1457,N_1494);
xor U1574 (N_1574,N_1444,N_1410);
nand U1575 (N_1575,N_1402,N_1487);
nor U1576 (N_1576,N_1460,N_1473);
nand U1577 (N_1577,N_1431,N_1401);
and U1578 (N_1578,N_1495,N_1402);
or U1579 (N_1579,N_1466,N_1482);
nor U1580 (N_1580,N_1461,N_1438);
nor U1581 (N_1581,N_1463,N_1439);
or U1582 (N_1582,N_1427,N_1439);
nand U1583 (N_1583,N_1489,N_1479);
and U1584 (N_1584,N_1463,N_1430);
nand U1585 (N_1585,N_1467,N_1485);
and U1586 (N_1586,N_1425,N_1480);
nor U1587 (N_1587,N_1464,N_1421);
or U1588 (N_1588,N_1433,N_1400);
or U1589 (N_1589,N_1434,N_1440);
xnor U1590 (N_1590,N_1412,N_1497);
nand U1591 (N_1591,N_1423,N_1419);
and U1592 (N_1592,N_1455,N_1402);
and U1593 (N_1593,N_1496,N_1473);
and U1594 (N_1594,N_1422,N_1430);
nor U1595 (N_1595,N_1486,N_1425);
nor U1596 (N_1596,N_1411,N_1444);
or U1597 (N_1597,N_1437,N_1456);
nor U1598 (N_1598,N_1432,N_1480);
nand U1599 (N_1599,N_1499,N_1413);
nand U1600 (N_1600,N_1544,N_1572);
nor U1601 (N_1601,N_1547,N_1570);
or U1602 (N_1602,N_1594,N_1582);
xor U1603 (N_1603,N_1527,N_1566);
or U1604 (N_1604,N_1502,N_1510);
nor U1605 (N_1605,N_1552,N_1596);
or U1606 (N_1606,N_1581,N_1592);
nor U1607 (N_1607,N_1577,N_1545);
and U1608 (N_1608,N_1576,N_1519);
and U1609 (N_1609,N_1537,N_1526);
or U1610 (N_1610,N_1589,N_1516);
and U1611 (N_1611,N_1571,N_1597);
nand U1612 (N_1612,N_1524,N_1551);
nand U1613 (N_1613,N_1557,N_1543);
and U1614 (N_1614,N_1532,N_1573);
nand U1615 (N_1615,N_1506,N_1522);
nand U1616 (N_1616,N_1501,N_1529);
or U1617 (N_1617,N_1559,N_1569);
and U1618 (N_1618,N_1538,N_1535);
nor U1619 (N_1619,N_1565,N_1525);
xnor U1620 (N_1620,N_1518,N_1588);
nand U1621 (N_1621,N_1536,N_1562);
nor U1622 (N_1622,N_1586,N_1598);
and U1623 (N_1623,N_1555,N_1504);
nand U1624 (N_1624,N_1534,N_1595);
nand U1625 (N_1625,N_1507,N_1512);
or U1626 (N_1626,N_1556,N_1542);
nor U1627 (N_1627,N_1591,N_1540);
nor U1628 (N_1628,N_1554,N_1517);
nand U1629 (N_1629,N_1503,N_1530);
or U1630 (N_1630,N_1511,N_1599);
nor U1631 (N_1631,N_1528,N_1587);
nor U1632 (N_1632,N_1500,N_1567);
nor U1633 (N_1633,N_1505,N_1550);
nand U1634 (N_1634,N_1539,N_1509);
nand U1635 (N_1635,N_1515,N_1533);
or U1636 (N_1636,N_1578,N_1560);
nor U1637 (N_1637,N_1553,N_1513);
and U1638 (N_1638,N_1585,N_1568);
nand U1639 (N_1639,N_1521,N_1520);
nand U1640 (N_1640,N_1584,N_1546);
and U1641 (N_1641,N_1541,N_1593);
and U1642 (N_1642,N_1590,N_1548);
and U1643 (N_1643,N_1564,N_1563);
or U1644 (N_1644,N_1583,N_1579);
xnor U1645 (N_1645,N_1561,N_1575);
and U1646 (N_1646,N_1508,N_1523);
nand U1647 (N_1647,N_1514,N_1580);
nand U1648 (N_1648,N_1531,N_1558);
and U1649 (N_1649,N_1549,N_1574);
nor U1650 (N_1650,N_1513,N_1529);
and U1651 (N_1651,N_1597,N_1523);
nor U1652 (N_1652,N_1594,N_1584);
nor U1653 (N_1653,N_1581,N_1588);
nand U1654 (N_1654,N_1569,N_1537);
and U1655 (N_1655,N_1524,N_1503);
and U1656 (N_1656,N_1582,N_1581);
and U1657 (N_1657,N_1536,N_1576);
xor U1658 (N_1658,N_1575,N_1560);
nand U1659 (N_1659,N_1554,N_1588);
or U1660 (N_1660,N_1584,N_1569);
xor U1661 (N_1661,N_1511,N_1547);
and U1662 (N_1662,N_1587,N_1524);
nand U1663 (N_1663,N_1594,N_1507);
nand U1664 (N_1664,N_1590,N_1506);
and U1665 (N_1665,N_1503,N_1527);
and U1666 (N_1666,N_1522,N_1573);
nand U1667 (N_1667,N_1528,N_1538);
and U1668 (N_1668,N_1535,N_1597);
nand U1669 (N_1669,N_1548,N_1525);
and U1670 (N_1670,N_1546,N_1515);
nand U1671 (N_1671,N_1583,N_1543);
nor U1672 (N_1672,N_1582,N_1565);
and U1673 (N_1673,N_1533,N_1505);
and U1674 (N_1674,N_1541,N_1517);
or U1675 (N_1675,N_1539,N_1521);
or U1676 (N_1676,N_1569,N_1565);
or U1677 (N_1677,N_1545,N_1565);
and U1678 (N_1678,N_1598,N_1501);
nand U1679 (N_1679,N_1570,N_1506);
nand U1680 (N_1680,N_1535,N_1588);
nor U1681 (N_1681,N_1564,N_1599);
xor U1682 (N_1682,N_1548,N_1536);
nor U1683 (N_1683,N_1537,N_1545);
nand U1684 (N_1684,N_1539,N_1527);
or U1685 (N_1685,N_1570,N_1582);
or U1686 (N_1686,N_1537,N_1535);
and U1687 (N_1687,N_1519,N_1582);
and U1688 (N_1688,N_1568,N_1535);
xnor U1689 (N_1689,N_1561,N_1523);
nor U1690 (N_1690,N_1542,N_1506);
nand U1691 (N_1691,N_1563,N_1513);
or U1692 (N_1692,N_1531,N_1528);
and U1693 (N_1693,N_1558,N_1534);
nor U1694 (N_1694,N_1520,N_1563);
xor U1695 (N_1695,N_1508,N_1551);
or U1696 (N_1696,N_1556,N_1514);
nor U1697 (N_1697,N_1591,N_1577);
nor U1698 (N_1698,N_1539,N_1515);
nand U1699 (N_1699,N_1587,N_1521);
and U1700 (N_1700,N_1634,N_1659);
nor U1701 (N_1701,N_1648,N_1646);
or U1702 (N_1702,N_1631,N_1666);
and U1703 (N_1703,N_1603,N_1682);
nor U1704 (N_1704,N_1692,N_1688);
nor U1705 (N_1705,N_1697,N_1694);
nand U1706 (N_1706,N_1686,N_1628);
nand U1707 (N_1707,N_1690,N_1643);
nand U1708 (N_1708,N_1622,N_1621);
or U1709 (N_1709,N_1614,N_1689);
nor U1710 (N_1710,N_1684,N_1651);
or U1711 (N_1711,N_1683,N_1606);
xor U1712 (N_1712,N_1620,N_1632);
nand U1713 (N_1713,N_1638,N_1644);
and U1714 (N_1714,N_1640,N_1696);
nor U1715 (N_1715,N_1662,N_1635);
xnor U1716 (N_1716,N_1641,N_1655);
nand U1717 (N_1717,N_1674,N_1676);
nand U1718 (N_1718,N_1691,N_1650);
nand U1719 (N_1719,N_1608,N_1613);
xnor U1720 (N_1720,N_1675,N_1681);
xor U1721 (N_1721,N_1605,N_1699);
or U1722 (N_1722,N_1670,N_1612);
nand U1723 (N_1723,N_1639,N_1673);
nand U1724 (N_1724,N_1668,N_1663);
and U1725 (N_1725,N_1654,N_1625);
nand U1726 (N_1726,N_1664,N_1629);
xnor U1727 (N_1727,N_1604,N_1633);
or U1728 (N_1728,N_1607,N_1658);
and U1729 (N_1729,N_1609,N_1669);
and U1730 (N_1730,N_1626,N_1678);
xnor U1731 (N_1731,N_1636,N_1610);
nor U1732 (N_1732,N_1616,N_1618);
or U1733 (N_1733,N_1695,N_1656);
or U1734 (N_1734,N_1619,N_1611);
or U1735 (N_1735,N_1601,N_1671);
nor U1736 (N_1736,N_1657,N_1680);
and U1737 (N_1737,N_1630,N_1623);
and U1738 (N_1738,N_1672,N_1667);
nor U1739 (N_1739,N_1687,N_1642);
nor U1740 (N_1740,N_1615,N_1600);
nand U1741 (N_1741,N_1661,N_1693);
and U1742 (N_1742,N_1685,N_1647);
nor U1743 (N_1743,N_1698,N_1679);
and U1744 (N_1744,N_1660,N_1649);
xnor U1745 (N_1745,N_1627,N_1677);
or U1746 (N_1746,N_1645,N_1617);
and U1747 (N_1747,N_1624,N_1637);
nor U1748 (N_1748,N_1665,N_1652);
nand U1749 (N_1749,N_1653,N_1602);
nor U1750 (N_1750,N_1620,N_1661);
and U1751 (N_1751,N_1673,N_1658);
and U1752 (N_1752,N_1608,N_1667);
nand U1753 (N_1753,N_1651,N_1698);
nor U1754 (N_1754,N_1678,N_1694);
nand U1755 (N_1755,N_1686,N_1678);
and U1756 (N_1756,N_1667,N_1678);
and U1757 (N_1757,N_1690,N_1657);
and U1758 (N_1758,N_1629,N_1600);
nand U1759 (N_1759,N_1654,N_1621);
nor U1760 (N_1760,N_1680,N_1612);
or U1761 (N_1761,N_1651,N_1648);
nor U1762 (N_1762,N_1637,N_1644);
or U1763 (N_1763,N_1637,N_1609);
or U1764 (N_1764,N_1609,N_1625);
nor U1765 (N_1765,N_1640,N_1678);
xor U1766 (N_1766,N_1604,N_1670);
nor U1767 (N_1767,N_1653,N_1678);
or U1768 (N_1768,N_1690,N_1666);
nand U1769 (N_1769,N_1677,N_1672);
and U1770 (N_1770,N_1636,N_1657);
and U1771 (N_1771,N_1632,N_1646);
nand U1772 (N_1772,N_1653,N_1615);
nor U1773 (N_1773,N_1691,N_1646);
nand U1774 (N_1774,N_1668,N_1621);
xnor U1775 (N_1775,N_1654,N_1684);
or U1776 (N_1776,N_1667,N_1617);
and U1777 (N_1777,N_1689,N_1639);
nand U1778 (N_1778,N_1668,N_1693);
and U1779 (N_1779,N_1603,N_1616);
and U1780 (N_1780,N_1634,N_1653);
xor U1781 (N_1781,N_1647,N_1699);
xor U1782 (N_1782,N_1664,N_1612);
nand U1783 (N_1783,N_1681,N_1671);
nor U1784 (N_1784,N_1620,N_1681);
nor U1785 (N_1785,N_1623,N_1658);
nand U1786 (N_1786,N_1690,N_1640);
or U1787 (N_1787,N_1672,N_1634);
and U1788 (N_1788,N_1680,N_1616);
nand U1789 (N_1789,N_1614,N_1637);
or U1790 (N_1790,N_1619,N_1658);
nor U1791 (N_1791,N_1618,N_1699);
and U1792 (N_1792,N_1676,N_1610);
nand U1793 (N_1793,N_1658,N_1698);
xnor U1794 (N_1794,N_1691,N_1638);
nor U1795 (N_1795,N_1608,N_1696);
and U1796 (N_1796,N_1657,N_1604);
nor U1797 (N_1797,N_1664,N_1613);
nor U1798 (N_1798,N_1678,N_1636);
or U1799 (N_1799,N_1654,N_1622);
xnor U1800 (N_1800,N_1702,N_1794);
or U1801 (N_1801,N_1796,N_1779);
nand U1802 (N_1802,N_1704,N_1795);
and U1803 (N_1803,N_1750,N_1769);
nor U1804 (N_1804,N_1771,N_1729);
or U1805 (N_1805,N_1737,N_1716);
nand U1806 (N_1806,N_1757,N_1777);
nor U1807 (N_1807,N_1713,N_1752);
or U1808 (N_1808,N_1765,N_1723);
nor U1809 (N_1809,N_1740,N_1754);
nand U1810 (N_1810,N_1708,N_1761);
xnor U1811 (N_1811,N_1741,N_1742);
or U1812 (N_1812,N_1780,N_1764);
or U1813 (N_1813,N_1774,N_1721);
xnor U1814 (N_1814,N_1743,N_1747);
nand U1815 (N_1815,N_1753,N_1772);
nand U1816 (N_1816,N_1759,N_1751);
or U1817 (N_1817,N_1785,N_1782);
or U1818 (N_1818,N_1730,N_1793);
or U1819 (N_1819,N_1781,N_1710);
nor U1820 (N_1820,N_1731,N_1727);
xor U1821 (N_1821,N_1715,N_1749);
xnor U1822 (N_1822,N_1786,N_1714);
or U1823 (N_1823,N_1768,N_1789);
xor U1824 (N_1824,N_1711,N_1790);
nor U1825 (N_1825,N_1773,N_1739);
and U1826 (N_1826,N_1755,N_1706);
nand U1827 (N_1827,N_1736,N_1788);
nor U1828 (N_1828,N_1798,N_1760);
nor U1829 (N_1829,N_1734,N_1756);
nand U1830 (N_1830,N_1775,N_1746);
and U1831 (N_1831,N_1717,N_1705);
and U1832 (N_1832,N_1725,N_1718);
and U1833 (N_1833,N_1762,N_1700);
nor U1834 (N_1834,N_1748,N_1784);
and U1835 (N_1835,N_1744,N_1720);
nor U1836 (N_1836,N_1797,N_1728);
nand U1837 (N_1837,N_1758,N_1709);
nor U1838 (N_1838,N_1763,N_1738);
or U1839 (N_1839,N_1712,N_1732);
xor U1840 (N_1840,N_1776,N_1783);
nor U1841 (N_1841,N_1767,N_1766);
nand U1842 (N_1842,N_1707,N_1770);
nor U1843 (N_1843,N_1733,N_1701);
or U1844 (N_1844,N_1778,N_1724);
nor U1845 (N_1845,N_1703,N_1735);
or U1846 (N_1846,N_1726,N_1719);
xnor U1847 (N_1847,N_1799,N_1791);
or U1848 (N_1848,N_1787,N_1745);
and U1849 (N_1849,N_1722,N_1792);
nand U1850 (N_1850,N_1722,N_1710);
nor U1851 (N_1851,N_1798,N_1747);
nand U1852 (N_1852,N_1784,N_1787);
nor U1853 (N_1853,N_1758,N_1768);
nor U1854 (N_1854,N_1779,N_1733);
nand U1855 (N_1855,N_1701,N_1736);
and U1856 (N_1856,N_1788,N_1778);
nand U1857 (N_1857,N_1764,N_1749);
or U1858 (N_1858,N_1725,N_1773);
xor U1859 (N_1859,N_1739,N_1797);
and U1860 (N_1860,N_1783,N_1720);
and U1861 (N_1861,N_1701,N_1715);
nand U1862 (N_1862,N_1724,N_1771);
or U1863 (N_1863,N_1788,N_1733);
nand U1864 (N_1864,N_1708,N_1741);
nand U1865 (N_1865,N_1779,N_1776);
nor U1866 (N_1866,N_1765,N_1735);
nand U1867 (N_1867,N_1744,N_1792);
or U1868 (N_1868,N_1767,N_1720);
nor U1869 (N_1869,N_1776,N_1716);
nor U1870 (N_1870,N_1733,N_1738);
nand U1871 (N_1871,N_1730,N_1775);
nand U1872 (N_1872,N_1752,N_1754);
nor U1873 (N_1873,N_1741,N_1730);
nand U1874 (N_1874,N_1798,N_1723);
nor U1875 (N_1875,N_1776,N_1761);
and U1876 (N_1876,N_1791,N_1767);
nand U1877 (N_1877,N_1713,N_1792);
nand U1878 (N_1878,N_1775,N_1764);
nand U1879 (N_1879,N_1708,N_1782);
and U1880 (N_1880,N_1728,N_1783);
and U1881 (N_1881,N_1795,N_1760);
nor U1882 (N_1882,N_1728,N_1704);
or U1883 (N_1883,N_1709,N_1787);
or U1884 (N_1884,N_1711,N_1718);
and U1885 (N_1885,N_1747,N_1774);
or U1886 (N_1886,N_1778,N_1749);
or U1887 (N_1887,N_1734,N_1780);
xnor U1888 (N_1888,N_1775,N_1780);
xor U1889 (N_1889,N_1777,N_1768);
and U1890 (N_1890,N_1795,N_1762);
nor U1891 (N_1891,N_1736,N_1718);
nor U1892 (N_1892,N_1730,N_1782);
nor U1893 (N_1893,N_1776,N_1765);
nand U1894 (N_1894,N_1721,N_1709);
nor U1895 (N_1895,N_1797,N_1762);
nor U1896 (N_1896,N_1751,N_1798);
and U1897 (N_1897,N_1707,N_1731);
and U1898 (N_1898,N_1799,N_1706);
or U1899 (N_1899,N_1753,N_1771);
nor U1900 (N_1900,N_1812,N_1870);
and U1901 (N_1901,N_1884,N_1810);
nand U1902 (N_1902,N_1821,N_1879);
nor U1903 (N_1903,N_1820,N_1829);
or U1904 (N_1904,N_1860,N_1858);
xnor U1905 (N_1905,N_1853,N_1877);
and U1906 (N_1906,N_1808,N_1866);
or U1907 (N_1907,N_1896,N_1873);
nor U1908 (N_1908,N_1830,N_1842);
nand U1909 (N_1909,N_1844,N_1836);
or U1910 (N_1910,N_1802,N_1882);
nand U1911 (N_1911,N_1826,N_1883);
xnor U1912 (N_1912,N_1869,N_1876);
nor U1913 (N_1913,N_1813,N_1854);
or U1914 (N_1914,N_1804,N_1875);
xnor U1915 (N_1915,N_1837,N_1849);
xor U1916 (N_1916,N_1818,N_1806);
and U1917 (N_1917,N_1828,N_1861);
nand U1918 (N_1918,N_1827,N_1893);
nor U1919 (N_1919,N_1809,N_1817);
or U1920 (N_1920,N_1859,N_1864);
nor U1921 (N_1921,N_1811,N_1863);
and U1922 (N_1922,N_1855,N_1825);
nand U1923 (N_1923,N_1898,N_1839);
and U1924 (N_1924,N_1840,N_1851);
xnor U1925 (N_1925,N_1815,N_1889);
nand U1926 (N_1926,N_1897,N_1823);
and U1927 (N_1927,N_1899,N_1880);
xor U1928 (N_1928,N_1857,N_1868);
nand U1929 (N_1929,N_1814,N_1805);
nor U1930 (N_1930,N_1822,N_1832);
nand U1931 (N_1931,N_1848,N_1807);
nor U1932 (N_1932,N_1856,N_1865);
and U1933 (N_1933,N_1881,N_1872);
nand U1934 (N_1934,N_1894,N_1891);
and U1935 (N_1935,N_1824,N_1888);
or U1936 (N_1936,N_1816,N_1831);
or U1937 (N_1937,N_1841,N_1846);
nor U1938 (N_1938,N_1887,N_1838);
nand U1939 (N_1939,N_1890,N_1895);
and U1940 (N_1940,N_1800,N_1801);
and U1941 (N_1941,N_1867,N_1874);
or U1942 (N_1942,N_1834,N_1847);
nand U1943 (N_1943,N_1850,N_1803);
or U1944 (N_1944,N_1819,N_1892);
or U1945 (N_1945,N_1871,N_1833);
xnor U1946 (N_1946,N_1852,N_1885);
nor U1947 (N_1947,N_1886,N_1845);
nand U1948 (N_1948,N_1878,N_1843);
nor U1949 (N_1949,N_1862,N_1835);
nand U1950 (N_1950,N_1842,N_1879);
nand U1951 (N_1951,N_1867,N_1842);
nor U1952 (N_1952,N_1829,N_1836);
xor U1953 (N_1953,N_1860,N_1810);
and U1954 (N_1954,N_1812,N_1854);
nor U1955 (N_1955,N_1846,N_1899);
or U1956 (N_1956,N_1891,N_1806);
or U1957 (N_1957,N_1859,N_1869);
nand U1958 (N_1958,N_1883,N_1840);
nor U1959 (N_1959,N_1855,N_1886);
nor U1960 (N_1960,N_1858,N_1807);
nor U1961 (N_1961,N_1840,N_1836);
nand U1962 (N_1962,N_1865,N_1821);
nand U1963 (N_1963,N_1846,N_1868);
xnor U1964 (N_1964,N_1804,N_1838);
and U1965 (N_1965,N_1836,N_1873);
xor U1966 (N_1966,N_1838,N_1888);
and U1967 (N_1967,N_1887,N_1803);
nor U1968 (N_1968,N_1813,N_1851);
nor U1969 (N_1969,N_1837,N_1871);
and U1970 (N_1970,N_1807,N_1853);
or U1971 (N_1971,N_1854,N_1858);
or U1972 (N_1972,N_1822,N_1871);
nor U1973 (N_1973,N_1841,N_1864);
xor U1974 (N_1974,N_1834,N_1827);
nand U1975 (N_1975,N_1830,N_1872);
nor U1976 (N_1976,N_1809,N_1811);
or U1977 (N_1977,N_1889,N_1806);
nand U1978 (N_1978,N_1857,N_1873);
or U1979 (N_1979,N_1883,N_1880);
nor U1980 (N_1980,N_1862,N_1894);
nand U1981 (N_1981,N_1816,N_1887);
nor U1982 (N_1982,N_1824,N_1886);
nand U1983 (N_1983,N_1880,N_1823);
and U1984 (N_1984,N_1882,N_1880);
and U1985 (N_1985,N_1885,N_1840);
and U1986 (N_1986,N_1873,N_1817);
nor U1987 (N_1987,N_1812,N_1815);
and U1988 (N_1988,N_1802,N_1865);
or U1989 (N_1989,N_1856,N_1803);
xnor U1990 (N_1990,N_1817,N_1894);
nor U1991 (N_1991,N_1873,N_1861);
nand U1992 (N_1992,N_1822,N_1873);
nand U1993 (N_1993,N_1860,N_1891);
xor U1994 (N_1994,N_1844,N_1800);
and U1995 (N_1995,N_1896,N_1894);
or U1996 (N_1996,N_1892,N_1873);
xor U1997 (N_1997,N_1838,N_1807);
nor U1998 (N_1998,N_1815,N_1894);
nand U1999 (N_1999,N_1877,N_1896);
and U2000 (N_2000,N_1918,N_1914);
nor U2001 (N_2001,N_1920,N_1982);
or U2002 (N_2002,N_1967,N_1921);
and U2003 (N_2003,N_1922,N_1942);
nand U2004 (N_2004,N_1961,N_1976);
nor U2005 (N_2005,N_1904,N_1963);
or U2006 (N_2006,N_1974,N_1960);
nand U2007 (N_2007,N_1912,N_1955);
or U2008 (N_2008,N_1925,N_1903);
nand U2009 (N_2009,N_1924,N_1994);
and U2010 (N_2010,N_1995,N_1935);
or U2011 (N_2011,N_1954,N_1991);
and U2012 (N_2012,N_1964,N_1940);
and U2013 (N_2013,N_1928,N_1953);
nand U2014 (N_2014,N_1999,N_1962);
and U2015 (N_2015,N_1948,N_1958);
or U2016 (N_2016,N_1992,N_1900);
or U2017 (N_2017,N_1966,N_1996);
xnor U2018 (N_2018,N_1984,N_1977);
or U2019 (N_2019,N_1998,N_1926);
nand U2020 (N_2020,N_1979,N_1931);
and U2021 (N_2021,N_1944,N_1937);
and U2022 (N_2022,N_1941,N_1930);
nand U2023 (N_2023,N_1970,N_1983);
and U2024 (N_2024,N_1986,N_1956);
nor U2025 (N_2025,N_1978,N_1933);
nand U2026 (N_2026,N_1945,N_1913);
xor U2027 (N_2027,N_1910,N_1936);
nand U2028 (N_2028,N_1916,N_1943);
or U2029 (N_2029,N_1923,N_1909);
xnor U2030 (N_2030,N_1929,N_1949);
nor U2031 (N_2031,N_1939,N_1927);
or U2032 (N_2032,N_1950,N_1907);
nand U2033 (N_2033,N_1902,N_1990);
nand U2034 (N_2034,N_1972,N_1938);
and U2035 (N_2035,N_1957,N_1932);
xor U2036 (N_2036,N_1980,N_1917);
xor U2037 (N_2037,N_1968,N_1906);
or U2038 (N_2038,N_1981,N_1975);
and U2039 (N_2039,N_1952,N_1969);
nor U2040 (N_2040,N_1988,N_1915);
or U2041 (N_2041,N_1989,N_1973);
nand U2042 (N_2042,N_1965,N_1919);
xor U2043 (N_2043,N_1997,N_1959);
or U2044 (N_2044,N_1971,N_1947);
and U2045 (N_2045,N_1901,N_1905);
nand U2046 (N_2046,N_1951,N_1985);
nor U2047 (N_2047,N_1987,N_1934);
nand U2048 (N_2048,N_1946,N_1908);
nor U2049 (N_2049,N_1993,N_1911);
nand U2050 (N_2050,N_1911,N_1913);
and U2051 (N_2051,N_1975,N_1971);
xnor U2052 (N_2052,N_1950,N_1908);
xnor U2053 (N_2053,N_1981,N_1938);
and U2054 (N_2054,N_1965,N_1949);
nand U2055 (N_2055,N_1985,N_1901);
nand U2056 (N_2056,N_1974,N_1906);
or U2057 (N_2057,N_1908,N_1948);
and U2058 (N_2058,N_1910,N_1984);
or U2059 (N_2059,N_1941,N_1917);
nand U2060 (N_2060,N_1944,N_1931);
or U2061 (N_2061,N_1951,N_1929);
or U2062 (N_2062,N_1952,N_1958);
nand U2063 (N_2063,N_1904,N_1902);
xnor U2064 (N_2064,N_1967,N_1946);
nand U2065 (N_2065,N_1989,N_1948);
or U2066 (N_2066,N_1911,N_1953);
or U2067 (N_2067,N_1986,N_1914);
and U2068 (N_2068,N_1964,N_1952);
or U2069 (N_2069,N_1946,N_1922);
xnor U2070 (N_2070,N_1996,N_1931);
or U2071 (N_2071,N_1976,N_1996);
nand U2072 (N_2072,N_1952,N_1995);
nor U2073 (N_2073,N_1904,N_1998);
nor U2074 (N_2074,N_1956,N_1920);
nand U2075 (N_2075,N_1915,N_1908);
nor U2076 (N_2076,N_1922,N_1983);
xor U2077 (N_2077,N_1908,N_1981);
nand U2078 (N_2078,N_1900,N_1924);
nand U2079 (N_2079,N_1925,N_1988);
and U2080 (N_2080,N_1986,N_1930);
nor U2081 (N_2081,N_1998,N_1995);
nand U2082 (N_2082,N_1956,N_1959);
xor U2083 (N_2083,N_1919,N_1926);
nand U2084 (N_2084,N_1998,N_1909);
or U2085 (N_2085,N_1989,N_1926);
nor U2086 (N_2086,N_1988,N_1970);
xnor U2087 (N_2087,N_1942,N_1908);
and U2088 (N_2088,N_1934,N_1902);
nand U2089 (N_2089,N_1976,N_1939);
xnor U2090 (N_2090,N_1970,N_1949);
and U2091 (N_2091,N_1979,N_1921);
nor U2092 (N_2092,N_1990,N_1980);
nand U2093 (N_2093,N_1940,N_1958);
or U2094 (N_2094,N_1964,N_1951);
and U2095 (N_2095,N_1940,N_1931);
nand U2096 (N_2096,N_1982,N_1998);
xnor U2097 (N_2097,N_1933,N_1957);
and U2098 (N_2098,N_1953,N_1955);
xor U2099 (N_2099,N_1986,N_1926);
nand U2100 (N_2100,N_2075,N_2095);
nand U2101 (N_2101,N_2057,N_2044);
xnor U2102 (N_2102,N_2077,N_2005);
or U2103 (N_2103,N_2062,N_2051);
nand U2104 (N_2104,N_2058,N_2072);
nor U2105 (N_2105,N_2063,N_2034);
or U2106 (N_2106,N_2067,N_2061);
and U2107 (N_2107,N_2025,N_2010);
nor U2108 (N_2108,N_2023,N_2042);
nand U2109 (N_2109,N_2086,N_2045);
nor U2110 (N_2110,N_2032,N_2098);
xnor U2111 (N_2111,N_2066,N_2093);
and U2112 (N_2112,N_2085,N_2038);
nor U2113 (N_2113,N_2089,N_2090);
nor U2114 (N_2114,N_2009,N_2073);
or U2115 (N_2115,N_2004,N_2001);
nand U2116 (N_2116,N_2015,N_2046);
or U2117 (N_2117,N_2031,N_2097);
nor U2118 (N_2118,N_2028,N_2035);
nand U2119 (N_2119,N_2059,N_2091);
nor U2120 (N_2120,N_2081,N_2041);
nand U2121 (N_2121,N_2054,N_2083);
nor U2122 (N_2122,N_2017,N_2024);
and U2123 (N_2123,N_2027,N_2018);
nor U2124 (N_2124,N_2026,N_2039);
and U2125 (N_2125,N_2021,N_2088);
nor U2126 (N_2126,N_2019,N_2076);
and U2127 (N_2127,N_2074,N_2096);
and U2128 (N_2128,N_2050,N_2013);
or U2129 (N_2129,N_2071,N_2070);
nor U2130 (N_2130,N_2052,N_2002);
nor U2131 (N_2131,N_2030,N_2043);
nor U2132 (N_2132,N_2014,N_2040);
or U2133 (N_2133,N_2033,N_2049);
nand U2134 (N_2134,N_2008,N_2016);
and U2135 (N_2135,N_2080,N_2099);
and U2136 (N_2136,N_2036,N_2094);
nor U2137 (N_2137,N_2003,N_2065);
xor U2138 (N_2138,N_2037,N_2029);
and U2139 (N_2139,N_2000,N_2055);
and U2140 (N_2140,N_2012,N_2020);
nand U2141 (N_2141,N_2084,N_2053);
and U2142 (N_2142,N_2079,N_2022);
nand U2143 (N_2143,N_2060,N_2006);
or U2144 (N_2144,N_2078,N_2056);
and U2145 (N_2145,N_2048,N_2047);
or U2146 (N_2146,N_2082,N_2092);
or U2147 (N_2147,N_2068,N_2087);
nor U2148 (N_2148,N_2007,N_2064);
xor U2149 (N_2149,N_2011,N_2069);
and U2150 (N_2150,N_2080,N_2086);
and U2151 (N_2151,N_2094,N_2096);
nor U2152 (N_2152,N_2021,N_2083);
and U2153 (N_2153,N_2002,N_2019);
xnor U2154 (N_2154,N_2002,N_2083);
nand U2155 (N_2155,N_2055,N_2065);
and U2156 (N_2156,N_2054,N_2044);
nor U2157 (N_2157,N_2029,N_2059);
and U2158 (N_2158,N_2011,N_2061);
xor U2159 (N_2159,N_2025,N_2043);
and U2160 (N_2160,N_2046,N_2052);
nor U2161 (N_2161,N_2013,N_2032);
or U2162 (N_2162,N_2001,N_2018);
or U2163 (N_2163,N_2043,N_2018);
and U2164 (N_2164,N_2089,N_2017);
nand U2165 (N_2165,N_2080,N_2046);
and U2166 (N_2166,N_2041,N_2017);
or U2167 (N_2167,N_2008,N_2061);
nor U2168 (N_2168,N_2052,N_2090);
or U2169 (N_2169,N_2008,N_2004);
or U2170 (N_2170,N_2039,N_2070);
nor U2171 (N_2171,N_2023,N_2073);
nand U2172 (N_2172,N_2095,N_2053);
nor U2173 (N_2173,N_2075,N_2068);
nand U2174 (N_2174,N_2055,N_2031);
and U2175 (N_2175,N_2016,N_2052);
xnor U2176 (N_2176,N_2085,N_2048);
nand U2177 (N_2177,N_2095,N_2099);
or U2178 (N_2178,N_2045,N_2057);
nor U2179 (N_2179,N_2088,N_2079);
nor U2180 (N_2180,N_2063,N_2076);
nand U2181 (N_2181,N_2012,N_2070);
and U2182 (N_2182,N_2000,N_2005);
nor U2183 (N_2183,N_2088,N_2027);
and U2184 (N_2184,N_2058,N_2005);
or U2185 (N_2185,N_2053,N_2056);
and U2186 (N_2186,N_2073,N_2044);
nor U2187 (N_2187,N_2041,N_2062);
and U2188 (N_2188,N_2051,N_2071);
nand U2189 (N_2189,N_2021,N_2008);
nor U2190 (N_2190,N_2009,N_2012);
or U2191 (N_2191,N_2018,N_2057);
xnor U2192 (N_2192,N_2004,N_2076);
nor U2193 (N_2193,N_2095,N_2085);
nand U2194 (N_2194,N_2048,N_2092);
nor U2195 (N_2195,N_2081,N_2058);
or U2196 (N_2196,N_2060,N_2055);
nor U2197 (N_2197,N_2053,N_2071);
nor U2198 (N_2198,N_2085,N_2046);
or U2199 (N_2199,N_2074,N_2021);
or U2200 (N_2200,N_2172,N_2151);
nand U2201 (N_2201,N_2177,N_2147);
or U2202 (N_2202,N_2161,N_2150);
or U2203 (N_2203,N_2128,N_2164);
and U2204 (N_2204,N_2191,N_2142);
xor U2205 (N_2205,N_2122,N_2104);
and U2206 (N_2206,N_2145,N_2158);
nor U2207 (N_2207,N_2187,N_2196);
or U2208 (N_2208,N_2165,N_2107);
nand U2209 (N_2209,N_2162,N_2100);
or U2210 (N_2210,N_2146,N_2111);
nand U2211 (N_2211,N_2188,N_2135);
and U2212 (N_2212,N_2192,N_2112);
or U2213 (N_2213,N_2183,N_2171);
and U2214 (N_2214,N_2117,N_2173);
and U2215 (N_2215,N_2166,N_2105);
or U2216 (N_2216,N_2155,N_2102);
nor U2217 (N_2217,N_2109,N_2148);
and U2218 (N_2218,N_2130,N_2114);
and U2219 (N_2219,N_2182,N_2134);
or U2220 (N_2220,N_2195,N_2119);
xor U2221 (N_2221,N_2168,N_2149);
or U2222 (N_2222,N_2194,N_2139);
and U2223 (N_2223,N_2156,N_2108);
nor U2224 (N_2224,N_2133,N_2184);
nor U2225 (N_2225,N_2197,N_2125);
or U2226 (N_2226,N_2179,N_2115);
nor U2227 (N_2227,N_2136,N_2110);
and U2228 (N_2228,N_2138,N_2154);
nand U2229 (N_2229,N_2123,N_2116);
or U2230 (N_2230,N_2186,N_2190);
or U2231 (N_2231,N_2120,N_2176);
and U2232 (N_2232,N_2106,N_2101);
nand U2233 (N_2233,N_2132,N_2180);
or U2234 (N_2234,N_2152,N_2160);
nor U2235 (N_2235,N_2137,N_2189);
xor U2236 (N_2236,N_2199,N_2143);
nand U2237 (N_2237,N_2141,N_2129);
xnor U2238 (N_2238,N_2153,N_2169);
nor U2239 (N_2239,N_2103,N_2185);
nor U2240 (N_2240,N_2163,N_2159);
nor U2241 (N_2241,N_2118,N_2167);
and U2242 (N_2242,N_2127,N_2181);
and U2243 (N_2243,N_2113,N_2175);
nor U2244 (N_2244,N_2124,N_2157);
or U2245 (N_2245,N_2126,N_2193);
nand U2246 (N_2246,N_2121,N_2178);
and U2247 (N_2247,N_2198,N_2170);
nand U2248 (N_2248,N_2131,N_2140);
nor U2249 (N_2249,N_2174,N_2144);
nand U2250 (N_2250,N_2142,N_2148);
xnor U2251 (N_2251,N_2145,N_2138);
or U2252 (N_2252,N_2116,N_2178);
and U2253 (N_2253,N_2153,N_2128);
nand U2254 (N_2254,N_2116,N_2107);
or U2255 (N_2255,N_2177,N_2178);
nor U2256 (N_2256,N_2113,N_2134);
nand U2257 (N_2257,N_2197,N_2168);
or U2258 (N_2258,N_2191,N_2148);
or U2259 (N_2259,N_2116,N_2133);
nor U2260 (N_2260,N_2147,N_2102);
or U2261 (N_2261,N_2122,N_2103);
nor U2262 (N_2262,N_2159,N_2120);
nand U2263 (N_2263,N_2139,N_2151);
and U2264 (N_2264,N_2105,N_2143);
and U2265 (N_2265,N_2110,N_2143);
xor U2266 (N_2266,N_2136,N_2106);
or U2267 (N_2267,N_2155,N_2120);
nand U2268 (N_2268,N_2181,N_2176);
or U2269 (N_2269,N_2181,N_2109);
and U2270 (N_2270,N_2172,N_2150);
xnor U2271 (N_2271,N_2163,N_2188);
nand U2272 (N_2272,N_2128,N_2169);
and U2273 (N_2273,N_2197,N_2139);
or U2274 (N_2274,N_2178,N_2102);
and U2275 (N_2275,N_2113,N_2146);
nor U2276 (N_2276,N_2185,N_2142);
nor U2277 (N_2277,N_2119,N_2161);
xnor U2278 (N_2278,N_2189,N_2196);
or U2279 (N_2279,N_2147,N_2192);
nor U2280 (N_2280,N_2131,N_2103);
and U2281 (N_2281,N_2159,N_2153);
xnor U2282 (N_2282,N_2183,N_2177);
or U2283 (N_2283,N_2104,N_2178);
or U2284 (N_2284,N_2178,N_2194);
or U2285 (N_2285,N_2107,N_2119);
and U2286 (N_2286,N_2147,N_2190);
nor U2287 (N_2287,N_2146,N_2119);
nand U2288 (N_2288,N_2109,N_2192);
and U2289 (N_2289,N_2162,N_2131);
nand U2290 (N_2290,N_2141,N_2139);
nor U2291 (N_2291,N_2193,N_2117);
xor U2292 (N_2292,N_2102,N_2111);
and U2293 (N_2293,N_2152,N_2107);
xnor U2294 (N_2294,N_2180,N_2140);
nand U2295 (N_2295,N_2164,N_2110);
nor U2296 (N_2296,N_2127,N_2131);
nand U2297 (N_2297,N_2128,N_2152);
nand U2298 (N_2298,N_2199,N_2178);
and U2299 (N_2299,N_2158,N_2134);
nand U2300 (N_2300,N_2218,N_2221);
xnor U2301 (N_2301,N_2248,N_2282);
nand U2302 (N_2302,N_2245,N_2260);
nor U2303 (N_2303,N_2229,N_2284);
and U2304 (N_2304,N_2294,N_2212);
or U2305 (N_2305,N_2231,N_2226);
or U2306 (N_2306,N_2210,N_2213);
and U2307 (N_2307,N_2280,N_2269);
or U2308 (N_2308,N_2242,N_2239);
nand U2309 (N_2309,N_2270,N_2202);
or U2310 (N_2310,N_2253,N_2211);
nand U2311 (N_2311,N_2216,N_2276);
or U2312 (N_2312,N_2208,N_2214);
or U2313 (N_2313,N_2278,N_2258);
nor U2314 (N_2314,N_2289,N_2256);
nor U2315 (N_2315,N_2283,N_2287);
nand U2316 (N_2316,N_2259,N_2271);
or U2317 (N_2317,N_2267,N_2261);
or U2318 (N_2318,N_2262,N_2298);
xor U2319 (N_2319,N_2292,N_2291);
nand U2320 (N_2320,N_2274,N_2243);
nor U2321 (N_2321,N_2265,N_2251);
nand U2322 (N_2322,N_2286,N_2257);
or U2323 (N_2323,N_2230,N_2217);
and U2324 (N_2324,N_2264,N_2219);
nand U2325 (N_2325,N_2275,N_2234);
and U2326 (N_2326,N_2224,N_2273);
nor U2327 (N_2327,N_2236,N_2206);
nor U2328 (N_2328,N_2295,N_2222);
or U2329 (N_2329,N_2281,N_2201);
nor U2330 (N_2330,N_2290,N_2235);
and U2331 (N_2331,N_2272,N_2279);
and U2332 (N_2332,N_2263,N_2228);
and U2333 (N_2333,N_2296,N_2204);
nor U2334 (N_2334,N_2233,N_2268);
xnor U2335 (N_2335,N_2299,N_2246);
and U2336 (N_2336,N_2241,N_2200);
xor U2337 (N_2337,N_2203,N_2215);
or U2338 (N_2338,N_2249,N_2225);
xnor U2339 (N_2339,N_2247,N_2237);
nand U2340 (N_2340,N_2252,N_2227);
nand U2341 (N_2341,N_2238,N_2223);
and U2342 (N_2342,N_2266,N_2255);
and U2343 (N_2343,N_2277,N_2288);
nor U2344 (N_2344,N_2293,N_2209);
nor U2345 (N_2345,N_2254,N_2244);
nand U2346 (N_2346,N_2285,N_2205);
and U2347 (N_2347,N_2207,N_2297);
and U2348 (N_2348,N_2220,N_2250);
nor U2349 (N_2349,N_2232,N_2240);
or U2350 (N_2350,N_2291,N_2256);
or U2351 (N_2351,N_2277,N_2263);
nor U2352 (N_2352,N_2204,N_2232);
nand U2353 (N_2353,N_2211,N_2294);
nor U2354 (N_2354,N_2207,N_2287);
and U2355 (N_2355,N_2283,N_2236);
and U2356 (N_2356,N_2224,N_2267);
nand U2357 (N_2357,N_2272,N_2283);
and U2358 (N_2358,N_2206,N_2269);
nor U2359 (N_2359,N_2299,N_2292);
nor U2360 (N_2360,N_2281,N_2232);
nor U2361 (N_2361,N_2286,N_2229);
nand U2362 (N_2362,N_2213,N_2236);
nand U2363 (N_2363,N_2222,N_2202);
nor U2364 (N_2364,N_2208,N_2294);
xnor U2365 (N_2365,N_2233,N_2248);
nor U2366 (N_2366,N_2274,N_2284);
nor U2367 (N_2367,N_2249,N_2284);
nor U2368 (N_2368,N_2236,N_2243);
nand U2369 (N_2369,N_2213,N_2203);
nor U2370 (N_2370,N_2236,N_2279);
nand U2371 (N_2371,N_2226,N_2242);
or U2372 (N_2372,N_2275,N_2237);
nand U2373 (N_2373,N_2212,N_2226);
or U2374 (N_2374,N_2213,N_2260);
nor U2375 (N_2375,N_2261,N_2277);
and U2376 (N_2376,N_2223,N_2263);
and U2377 (N_2377,N_2270,N_2219);
and U2378 (N_2378,N_2250,N_2269);
nand U2379 (N_2379,N_2217,N_2294);
or U2380 (N_2380,N_2271,N_2227);
and U2381 (N_2381,N_2232,N_2229);
nand U2382 (N_2382,N_2250,N_2206);
nand U2383 (N_2383,N_2290,N_2259);
nor U2384 (N_2384,N_2262,N_2267);
nand U2385 (N_2385,N_2215,N_2284);
or U2386 (N_2386,N_2251,N_2244);
or U2387 (N_2387,N_2264,N_2237);
or U2388 (N_2388,N_2270,N_2277);
nor U2389 (N_2389,N_2239,N_2297);
xnor U2390 (N_2390,N_2231,N_2212);
nor U2391 (N_2391,N_2259,N_2221);
and U2392 (N_2392,N_2286,N_2239);
nand U2393 (N_2393,N_2202,N_2261);
and U2394 (N_2394,N_2299,N_2239);
nor U2395 (N_2395,N_2200,N_2206);
nor U2396 (N_2396,N_2221,N_2243);
or U2397 (N_2397,N_2237,N_2278);
or U2398 (N_2398,N_2254,N_2295);
nor U2399 (N_2399,N_2246,N_2253);
nor U2400 (N_2400,N_2333,N_2378);
nand U2401 (N_2401,N_2304,N_2356);
xor U2402 (N_2402,N_2391,N_2395);
nor U2403 (N_2403,N_2339,N_2375);
and U2404 (N_2404,N_2393,N_2377);
or U2405 (N_2405,N_2341,N_2387);
xnor U2406 (N_2406,N_2316,N_2397);
nand U2407 (N_2407,N_2343,N_2370);
nor U2408 (N_2408,N_2373,N_2398);
nor U2409 (N_2409,N_2388,N_2300);
or U2410 (N_2410,N_2322,N_2357);
nor U2411 (N_2411,N_2324,N_2392);
and U2412 (N_2412,N_2361,N_2347);
nand U2413 (N_2413,N_2321,N_2394);
or U2414 (N_2414,N_2379,N_2327);
and U2415 (N_2415,N_2381,N_2323);
and U2416 (N_2416,N_2372,N_2376);
nand U2417 (N_2417,N_2349,N_2328);
and U2418 (N_2418,N_2311,N_2334);
nor U2419 (N_2419,N_2362,N_2306);
nor U2420 (N_2420,N_2354,N_2371);
nor U2421 (N_2421,N_2364,N_2390);
or U2422 (N_2422,N_2345,N_2363);
nand U2423 (N_2423,N_2320,N_2380);
and U2424 (N_2424,N_2382,N_2338);
xor U2425 (N_2425,N_2318,N_2369);
or U2426 (N_2426,N_2342,N_2308);
xor U2427 (N_2427,N_2368,N_2355);
xor U2428 (N_2428,N_2374,N_2337);
nand U2429 (N_2429,N_2344,N_2325);
nor U2430 (N_2430,N_2331,N_2360);
nand U2431 (N_2431,N_2350,N_2326);
or U2432 (N_2432,N_2367,N_2307);
or U2433 (N_2433,N_2309,N_2352);
nand U2434 (N_2434,N_2396,N_2358);
or U2435 (N_2435,N_2385,N_2319);
nand U2436 (N_2436,N_2301,N_2353);
and U2437 (N_2437,N_2340,N_2330);
xor U2438 (N_2438,N_2365,N_2351);
or U2439 (N_2439,N_2389,N_2366);
nand U2440 (N_2440,N_2329,N_2312);
and U2441 (N_2441,N_2315,N_2305);
nand U2442 (N_2442,N_2332,N_2303);
nor U2443 (N_2443,N_2317,N_2348);
nor U2444 (N_2444,N_2310,N_2399);
nor U2445 (N_2445,N_2386,N_2314);
nand U2446 (N_2446,N_2313,N_2302);
nor U2447 (N_2447,N_2383,N_2346);
and U2448 (N_2448,N_2384,N_2336);
and U2449 (N_2449,N_2359,N_2335);
or U2450 (N_2450,N_2387,N_2338);
or U2451 (N_2451,N_2361,N_2351);
and U2452 (N_2452,N_2336,N_2399);
or U2453 (N_2453,N_2334,N_2327);
nand U2454 (N_2454,N_2391,N_2372);
nand U2455 (N_2455,N_2354,N_2334);
nand U2456 (N_2456,N_2340,N_2397);
or U2457 (N_2457,N_2330,N_2383);
nor U2458 (N_2458,N_2357,N_2347);
and U2459 (N_2459,N_2391,N_2384);
xor U2460 (N_2460,N_2376,N_2300);
nor U2461 (N_2461,N_2316,N_2301);
nor U2462 (N_2462,N_2369,N_2386);
or U2463 (N_2463,N_2398,N_2391);
and U2464 (N_2464,N_2399,N_2364);
and U2465 (N_2465,N_2390,N_2367);
xnor U2466 (N_2466,N_2394,N_2382);
and U2467 (N_2467,N_2366,N_2363);
or U2468 (N_2468,N_2318,N_2312);
xnor U2469 (N_2469,N_2308,N_2316);
or U2470 (N_2470,N_2324,N_2345);
nor U2471 (N_2471,N_2330,N_2333);
xnor U2472 (N_2472,N_2376,N_2329);
nand U2473 (N_2473,N_2382,N_2324);
and U2474 (N_2474,N_2372,N_2349);
nand U2475 (N_2475,N_2350,N_2320);
nand U2476 (N_2476,N_2306,N_2346);
and U2477 (N_2477,N_2375,N_2302);
nor U2478 (N_2478,N_2347,N_2344);
xor U2479 (N_2479,N_2340,N_2303);
xor U2480 (N_2480,N_2380,N_2304);
xnor U2481 (N_2481,N_2301,N_2342);
and U2482 (N_2482,N_2350,N_2359);
nand U2483 (N_2483,N_2371,N_2379);
xnor U2484 (N_2484,N_2327,N_2312);
nor U2485 (N_2485,N_2338,N_2340);
nand U2486 (N_2486,N_2302,N_2360);
nor U2487 (N_2487,N_2373,N_2328);
nor U2488 (N_2488,N_2312,N_2330);
nand U2489 (N_2489,N_2311,N_2360);
or U2490 (N_2490,N_2329,N_2373);
and U2491 (N_2491,N_2349,N_2347);
nand U2492 (N_2492,N_2362,N_2346);
xor U2493 (N_2493,N_2322,N_2335);
nand U2494 (N_2494,N_2396,N_2332);
nand U2495 (N_2495,N_2300,N_2351);
and U2496 (N_2496,N_2308,N_2384);
nor U2497 (N_2497,N_2352,N_2357);
nand U2498 (N_2498,N_2317,N_2322);
and U2499 (N_2499,N_2344,N_2332);
or U2500 (N_2500,N_2457,N_2479);
nor U2501 (N_2501,N_2441,N_2486);
or U2502 (N_2502,N_2433,N_2485);
nand U2503 (N_2503,N_2462,N_2472);
xnor U2504 (N_2504,N_2413,N_2448);
or U2505 (N_2505,N_2487,N_2447);
and U2506 (N_2506,N_2474,N_2429);
nor U2507 (N_2507,N_2498,N_2404);
nand U2508 (N_2508,N_2469,N_2480);
nor U2509 (N_2509,N_2478,N_2461);
and U2510 (N_2510,N_2491,N_2475);
or U2511 (N_2511,N_2430,N_2445);
nor U2512 (N_2512,N_2453,N_2434);
nand U2513 (N_2513,N_2476,N_2432);
nor U2514 (N_2514,N_2449,N_2499);
nor U2515 (N_2515,N_2415,N_2436);
nor U2516 (N_2516,N_2496,N_2428);
nand U2517 (N_2517,N_2455,N_2421);
nor U2518 (N_2518,N_2438,N_2419);
nand U2519 (N_2519,N_2488,N_2437);
nand U2520 (N_2520,N_2467,N_2458);
xor U2521 (N_2521,N_2425,N_2440);
xnor U2522 (N_2522,N_2477,N_2463);
xnor U2523 (N_2523,N_2435,N_2482);
and U2524 (N_2524,N_2490,N_2443);
nor U2525 (N_2525,N_2465,N_2405);
nand U2526 (N_2526,N_2422,N_2450);
nand U2527 (N_2527,N_2492,N_2427);
nand U2528 (N_2528,N_2473,N_2466);
nor U2529 (N_2529,N_2484,N_2402);
or U2530 (N_2530,N_2407,N_2451);
or U2531 (N_2531,N_2444,N_2431);
and U2532 (N_2532,N_2493,N_2410);
nor U2533 (N_2533,N_2412,N_2470);
nor U2534 (N_2534,N_2416,N_2452);
nand U2535 (N_2535,N_2414,N_2426);
or U2536 (N_2536,N_2481,N_2401);
or U2537 (N_2537,N_2400,N_2423);
nor U2538 (N_2538,N_2417,N_2418);
or U2539 (N_2539,N_2471,N_2424);
nand U2540 (N_2540,N_2408,N_2406);
nor U2541 (N_2541,N_2420,N_2495);
and U2542 (N_2542,N_2494,N_2454);
xor U2543 (N_2543,N_2464,N_2459);
nand U2544 (N_2544,N_2456,N_2403);
and U2545 (N_2545,N_2439,N_2483);
nand U2546 (N_2546,N_2446,N_2409);
nor U2547 (N_2547,N_2460,N_2497);
nand U2548 (N_2548,N_2468,N_2411);
and U2549 (N_2549,N_2489,N_2442);
nand U2550 (N_2550,N_2407,N_2481);
and U2551 (N_2551,N_2487,N_2445);
nand U2552 (N_2552,N_2467,N_2408);
or U2553 (N_2553,N_2486,N_2432);
or U2554 (N_2554,N_2461,N_2405);
nand U2555 (N_2555,N_2447,N_2418);
nor U2556 (N_2556,N_2459,N_2452);
nor U2557 (N_2557,N_2499,N_2460);
nor U2558 (N_2558,N_2416,N_2463);
or U2559 (N_2559,N_2494,N_2420);
or U2560 (N_2560,N_2401,N_2426);
nand U2561 (N_2561,N_2408,N_2481);
and U2562 (N_2562,N_2402,N_2497);
or U2563 (N_2563,N_2469,N_2406);
nand U2564 (N_2564,N_2473,N_2406);
nand U2565 (N_2565,N_2426,N_2487);
xor U2566 (N_2566,N_2485,N_2408);
nor U2567 (N_2567,N_2410,N_2473);
xnor U2568 (N_2568,N_2491,N_2494);
nand U2569 (N_2569,N_2438,N_2437);
or U2570 (N_2570,N_2450,N_2434);
nand U2571 (N_2571,N_2430,N_2463);
or U2572 (N_2572,N_2472,N_2413);
nor U2573 (N_2573,N_2467,N_2477);
and U2574 (N_2574,N_2490,N_2426);
and U2575 (N_2575,N_2443,N_2483);
nor U2576 (N_2576,N_2470,N_2413);
and U2577 (N_2577,N_2497,N_2473);
nor U2578 (N_2578,N_2455,N_2412);
or U2579 (N_2579,N_2417,N_2462);
and U2580 (N_2580,N_2408,N_2429);
and U2581 (N_2581,N_2457,N_2471);
nand U2582 (N_2582,N_2475,N_2458);
nor U2583 (N_2583,N_2450,N_2462);
and U2584 (N_2584,N_2446,N_2449);
and U2585 (N_2585,N_2474,N_2467);
xor U2586 (N_2586,N_2484,N_2446);
nor U2587 (N_2587,N_2416,N_2449);
xor U2588 (N_2588,N_2457,N_2435);
or U2589 (N_2589,N_2486,N_2411);
nor U2590 (N_2590,N_2488,N_2412);
and U2591 (N_2591,N_2420,N_2411);
and U2592 (N_2592,N_2479,N_2485);
nand U2593 (N_2593,N_2428,N_2481);
xnor U2594 (N_2594,N_2487,N_2472);
nand U2595 (N_2595,N_2493,N_2460);
and U2596 (N_2596,N_2437,N_2472);
nand U2597 (N_2597,N_2434,N_2475);
nand U2598 (N_2598,N_2470,N_2427);
or U2599 (N_2599,N_2402,N_2479);
nand U2600 (N_2600,N_2542,N_2587);
nor U2601 (N_2601,N_2547,N_2538);
or U2602 (N_2602,N_2573,N_2527);
nor U2603 (N_2603,N_2531,N_2530);
and U2604 (N_2604,N_2578,N_2565);
and U2605 (N_2605,N_2549,N_2525);
and U2606 (N_2606,N_2536,N_2580);
nor U2607 (N_2607,N_2556,N_2500);
xor U2608 (N_2608,N_2563,N_2513);
or U2609 (N_2609,N_2521,N_2540);
and U2610 (N_2610,N_2522,N_2506);
nor U2611 (N_2611,N_2539,N_2515);
nor U2612 (N_2612,N_2544,N_2553);
nand U2613 (N_2613,N_2516,N_2576);
nor U2614 (N_2614,N_2507,N_2564);
xnor U2615 (N_2615,N_2597,N_2550);
nor U2616 (N_2616,N_2528,N_2501);
xor U2617 (N_2617,N_2532,N_2590);
nand U2618 (N_2618,N_2599,N_2584);
or U2619 (N_2619,N_2593,N_2552);
nand U2620 (N_2620,N_2561,N_2577);
nand U2621 (N_2621,N_2524,N_2535);
or U2622 (N_2622,N_2509,N_2554);
and U2623 (N_2623,N_2546,N_2508);
and U2624 (N_2624,N_2555,N_2541);
and U2625 (N_2625,N_2596,N_2558);
and U2626 (N_2626,N_2579,N_2598);
nand U2627 (N_2627,N_2519,N_2592);
nand U2628 (N_2628,N_2585,N_2586);
nor U2629 (N_2629,N_2588,N_2594);
and U2630 (N_2630,N_2510,N_2523);
nand U2631 (N_2631,N_2572,N_2560);
nand U2632 (N_2632,N_2570,N_2504);
or U2633 (N_2633,N_2548,N_2582);
nor U2634 (N_2634,N_2574,N_2589);
and U2635 (N_2635,N_2514,N_2557);
or U2636 (N_2636,N_2551,N_2517);
nand U2637 (N_2637,N_2545,N_2562);
xor U2638 (N_2638,N_2505,N_2583);
and U2639 (N_2639,N_2595,N_2503);
nand U2640 (N_2640,N_2529,N_2559);
nand U2641 (N_2641,N_2591,N_2569);
nor U2642 (N_2642,N_2543,N_2526);
nor U2643 (N_2643,N_2567,N_2502);
and U2644 (N_2644,N_2571,N_2568);
nor U2645 (N_2645,N_2581,N_2537);
or U2646 (N_2646,N_2575,N_2566);
nor U2647 (N_2647,N_2512,N_2520);
nand U2648 (N_2648,N_2533,N_2518);
nand U2649 (N_2649,N_2534,N_2511);
and U2650 (N_2650,N_2556,N_2586);
or U2651 (N_2651,N_2509,N_2572);
and U2652 (N_2652,N_2557,N_2512);
nor U2653 (N_2653,N_2594,N_2571);
nand U2654 (N_2654,N_2567,N_2597);
nand U2655 (N_2655,N_2589,N_2502);
and U2656 (N_2656,N_2516,N_2574);
nand U2657 (N_2657,N_2560,N_2538);
and U2658 (N_2658,N_2520,N_2524);
or U2659 (N_2659,N_2594,N_2505);
or U2660 (N_2660,N_2515,N_2510);
nand U2661 (N_2661,N_2538,N_2518);
nor U2662 (N_2662,N_2549,N_2533);
and U2663 (N_2663,N_2519,N_2513);
nor U2664 (N_2664,N_2590,N_2549);
and U2665 (N_2665,N_2562,N_2578);
nor U2666 (N_2666,N_2512,N_2528);
and U2667 (N_2667,N_2505,N_2561);
nand U2668 (N_2668,N_2511,N_2542);
or U2669 (N_2669,N_2521,N_2538);
and U2670 (N_2670,N_2511,N_2508);
and U2671 (N_2671,N_2554,N_2567);
nor U2672 (N_2672,N_2523,N_2531);
nor U2673 (N_2673,N_2593,N_2585);
and U2674 (N_2674,N_2539,N_2520);
or U2675 (N_2675,N_2537,N_2539);
nor U2676 (N_2676,N_2584,N_2535);
and U2677 (N_2677,N_2507,N_2572);
or U2678 (N_2678,N_2538,N_2504);
nor U2679 (N_2679,N_2579,N_2593);
nand U2680 (N_2680,N_2525,N_2550);
or U2681 (N_2681,N_2557,N_2561);
or U2682 (N_2682,N_2560,N_2508);
nand U2683 (N_2683,N_2525,N_2531);
or U2684 (N_2684,N_2589,N_2560);
nand U2685 (N_2685,N_2504,N_2555);
or U2686 (N_2686,N_2553,N_2562);
nor U2687 (N_2687,N_2547,N_2548);
or U2688 (N_2688,N_2554,N_2573);
xnor U2689 (N_2689,N_2548,N_2532);
nand U2690 (N_2690,N_2546,N_2524);
nor U2691 (N_2691,N_2562,N_2590);
xnor U2692 (N_2692,N_2564,N_2569);
and U2693 (N_2693,N_2524,N_2525);
nand U2694 (N_2694,N_2513,N_2517);
nor U2695 (N_2695,N_2512,N_2542);
or U2696 (N_2696,N_2529,N_2508);
nand U2697 (N_2697,N_2561,N_2517);
or U2698 (N_2698,N_2582,N_2599);
xnor U2699 (N_2699,N_2529,N_2567);
or U2700 (N_2700,N_2610,N_2694);
or U2701 (N_2701,N_2634,N_2623);
or U2702 (N_2702,N_2680,N_2632);
nand U2703 (N_2703,N_2604,N_2665);
nor U2704 (N_2704,N_2687,N_2602);
or U2705 (N_2705,N_2636,N_2631);
nand U2706 (N_2706,N_2639,N_2600);
and U2707 (N_2707,N_2612,N_2635);
nand U2708 (N_2708,N_2677,N_2674);
nor U2709 (N_2709,N_2654,N_2671);
or U2710 (N_2710,N_2670,N_2637);
nand U2711 (N_2711,N_2653,N_2603);
or U2712 (N_2712,N_2679,N_2648);
and U2713 (N_2713,N_2656,N_2613);
xor U2714 (N_2714,N_2622,N_2690);
and U2715 (N_2715,N_2668,N_2649);
and U2716 (N_2716,N_2696,N_2660);
nand U2717 (N_2717,N_2667,N_2642);
or U2718 (N_2718,N_2630,N_2606);
and U2719 (N_2719,N_2614,N_2657);
nor U2720 (N_2720,N_2684,N_2618);
nor U2721 (N_2721,N_2681,N_2669);
or U2722 (N_2722,N_2699,N_2628);
and U2723 (N_2723,N_2647,N_2659);
and U2724 (N_2724,N_2605,N_2640);
nand U2725 (N_2725,N_2619,N_2688);
nor U2726 (N_2726,N_2609,N_2646);
xor U2727 (N_2727,N_2644,N_2629);
and U2728 (N_2728,N_2672,N_2601);
or U2729 (N_2729,N_2645,N_2678);
nor U2730 (N_2730,N_2655,N_2617);
and U2731 (N_2731,N_2676,N_2611);
and U2732 (N_2732,N_2658,N_2624);
nand U2733 (N_2733,N_2607,N_2643);
or U2734 (N_2734,N_2686,N_2615);
nor U2735 (N_2735,N_2698,N_2692);
or U2736 (N_2736,N_2693,N_2650);
nor U2737 (N_2737,N_2663,N_2626);
or U2738 (N_2738,N_2685,N_2662);
and U2739 (N_2739,N_2608,N_2652);
or U2740 (N_2740,N_2625,N_2697);
xnor U2741 (N_2741,N_2633,N_2620);
or U2742 (N_2742,N_2661,N_2641);
nor U2743 (N_2743,N_2666,N_2627);
nand U2744 (N_2744,N_2689,N_2675);
nand U2745 (N_2745,N_2651,N_2664);
and U2746 (N_2746,N_2621,N_2673);
xnor U2747 (N_2747,N_2683,N_2682);
and U2748 (N_2748,N_2691,N_2616);
nand U2749 (N_2749,N_2695,N_2638);
or U2750 (N_2750,N_2601,N_2640);
nor U2751 (N_2751,N_2679,N_2605);
and U2752 (N_2752,N_2651,N_2614);
nand U2753 (N_2753,N_2601,N_2662);
or U2754 (N_2754,N_2601,N_2616);
xor U2755 (N_2755,N_2628,N_2683);
or U2756 (N_2756,N_2691,N_2688);
or U2757 (N_2757,N_2687,N_2662);
or U2758 (N_2758,N_2677,N_2644);
nand U2759 (N_2759,N_2689,N_2647);
and U2760 (N_2760,N_2642,N_2657);
and U2761 (N_2761,N_2672,N_2635);
and U2762 (N_2762,N_2672,N_2692);
and U2763 (N_2763,N_2660,N_2631);
nor U2764 (N_2764,N_2649,N_2676);
nor U2765 (N_2765,N_2635,N_2683);
and U2766 (N_2766,N_2601,N_2668);
and U2767 (N_2767,N_2672,N_2661);
nor U2768 (N_2768,N_2645,N_2682);
nand U2769 (N_2769,N_2688,N_2614);
nand U2770 (N_2770,N_2644,N_2615);
xnor U2771 (N_2771,N_2636,N_2640);
or U2772 (N_2772,N_2651,N_2696);
or U2773 (N_2773,N_2677,N_2602);
xnor U2774 (N_2774,N_2686,N_2657);
and U2775 (N_2775,N_2683,N_2669);
nand U2776 (N_2776,N_2630,N_2650);
or U2777 (N_2777,N_2635,N_2625);
nor U2778 (N_2778,N_2620,N_2632);
or U2779 (N_2779,N_2661,N_2613);
or U2780 (N_2780,N_2669,N_2666);
or U2781 (N_2781,N_2628,N_2624);
and U2782 (N_2782,N_2618,N_2656);
or U2783 (N_2783,N_2641,N_2614);
xor U2784 (N_2784,N_2662,N_2650);
nand U2785 (N_2785,N_2623,N_2683);
nand U2786 (N_2786,N_2636,N_2623);
and U2787 (N_2787,N_2620,N_2684);
and U2788 (N_2788,N_2605,N_2617);
nor U2789 (N_2789,N_2697,N_2609);
and U2790 (N_2790,N_2673,N_2631);
or U2791 (N_2791,N_2692,N_2674);
and U2792 (N_2792,N_2676,N_2606);
or U2793 (N_2793,N_2610,N_2607);
nor U2794 (N_2794,N_2618,N_2687);
or U2795 (N_2795,N_2611,N_2624);
xor U2796 (N_2796,N_2651,N_2671);
or U2797 (N_2797,N_2620,N_2699);
nor U2798 (N_2798,N_2658,N_2629);
xnor U2799 (N_2799,N_2640,N_2671);
nand U2800 (N_2800,N_2742,N_2744);
nor U2801 (N_2801,N_2717,N_2768);
and U2802 (N_2802,N_2731,N_2709);
and U2803 (N_2803,N_2778,N_2780);
nand U2804 (N_2804,N_2725,N_2735);
and U2805 (N_2805,N_2798,N_2779);
xor U2806 (N_2806,N_2783,N_2701);
and U2807 (N_2807,N_2732,N_2782);
nor U2808 (N_2808,N_2700,N_2730);
nor U2809 (N_2809,N_2781,N_2747);
xor U2810 (N_2810,N_2718,N_2790);
nor U2811 (N_2811,N_2796,N_2795);
xor U2812 (N_2812,N_2743,N_2772);
xor U2813 (N_2813,N_2786,N_2762);
or U2814 (N_2814,N_2722,N_2711);
nor U2815 (N_2815,N_2749,N_2793);
nor U2816 (N_2816,N_2754,N_2787);
nor U2817 (N_2817,N_2771,N_2770);
and U2818 (N_2818,N_2785,N_2774);
xnor U2819 (N_2819,N_2767,N_2737);
nor U2820 (N_2820,N_2758,N_2757);
nand U2821 (N_2821,N_2753,N_2784);
xor U2822 (N_2822,N_2703,N_2763);
or U2823 (N_2823,N_2766,N_2704);
nand U2824 (N_2824,N_2705,N_2729);
or U2825 (N_2825,N_2775,N_2728);
nor U2826 (N_2826,N_2765,N_2777);
nor U2827 (N_2827,N_2724,N_2746);
nand U2828 (N_2828,N_2713,N_2756);
nand U2829 (N_2829,N_2764,N_2706);
nor U2830 (N_2830,N_2797,N_2734);
nor U2831 (N_2831,N_2750,N_2773);
nor U2832 (N_2832,N_2719,N_2745);
nand U2833 (N_2833,N_2712,N_2788);
or U2834 (N_2834,N_2791,N_2714);
nand U2835 (N_2835,N_2738,N_2789);
and U2836 (N_2836,N_2769,N_2792);
nand U2837 (N_2837,N_2733,N_2740);
nor U2838 (N_2838,N_2702,N_2710);
and U2839 (N_2839,N_2708,N_2759);
xor U2840 (N_2840,N_2723,N_2761);
nand U2841 (N_2841,N_2752,N_2720);
or U2842 (N_2842,N_2776,N_2739);
nand U2843 (N_2843,N_2751,N_2721);
and U2844 (N_2844,N_2715,N_2716);
and U2845 (N_2845,N_2794,N_2741);
and U2846 (N_2846,N_2799,N_2727);
and U2847 (N_2847,N_2755,N_2760);
or U2848 (N_2848,N_2707,N_2726);
and U2849 (N_2849,N_2748,N_2736);
nand U2850 (N_2850,N_2771,N_2722);
and U2851 (N_2851,N_2761,N_2717);
and U2852 (N_2852,N_2743,N_2771);
and U2853 (N_2853,N_2729,N_2764);
xnor U2854 (N_2854,N_2784,N_2740);
nor U2855 (N_2855,N_2728,N_2786);
nor U2856 (N_2856,N_2721,N_2789);
and U2857 (N_2857,N_2743,N_2701);
nor U2858 (N_2858,N_2709,N_2746);
nor U2859 (N_2859,N_2724,N_2772);
or U2860 (N_2860,N_2789,N_2783);
or U2861 (N_2861,N_2789,N_2741);
nor U2862 (N_2862,N_2786,N_2748);
or U2863 (N_2863,N_2782,N_2724);
xor U2864 (N_2864,N_2795,N_2700);
or U2865 (N_2865,N_2731,N_2708);
and U2866 (N_2866,N_2737,N_2775);
or U2867 (N_2867,N_2787,N_2776);
nor U2868 (N_2868,N_2738,N_2701);
nand U2869 (N_2869,N_2744,N_2731);
nand U2870 (N_2870,N_2795,N_2740);
or U2871 (N_2871,N_2761,N_2732);
and U2872 (N_2872,N_2729,N_2720);
nand U2873 (N_2873,N_2752,N_2741);
nor U2874 (N_2874,N_2774,N_2782);
xnor U2875 (N_2875,N_2784,N_2731);
and U2876 (N_2876,N_2793,N_2701);
nor U2877 (N_2877,N_2732,N_2788);
nand U2878 (N_2878,N_2799,N_2752);
nor U2879 (N_2879,N_2790,N_2729);
or U2880 (N_2880,N_2710,N_2731);
nand U2881 (N_2881,N_2704,N_2728);
nand U2882 (N_2882,N_2725,N_2742);
or U2883 (N_2883,N_2748,N_2744);
or U2884 (N_2884,N_2703,N_2776);
or U2885 (N_2885,N_2760,N_2730);
nand U2886 (N_2886,N_2714,N_2797);
nor U2887 (N_2887,N_2724,N_2722);
or U2888 (N_2888,N_2726,N_2733);
nand U2889 (N_2889,N_2778,N_2734);
and U2890 (N_2890,N_2740,N_2799);
nand U2891 (N_2891,N_2786,N_2706);
nor U2892 (N_2892,N_2769,N_2742);
and U2893 (N_2893,N_2780,N_2710);
nand U2894 (N_2894,N_2711,N_2749);
or U2895 (N_2895,N_2787,N_2789);
nand U2896 (N_2896,N_2717,N_2719);
nand U2897 (N_2897,N_2743,N_2746);
nor U2898 (N_2898,N_2750,N_2765);
nand U2899 (N_2899,N_2707,N_2709);
and U2900 (N_2900,N_2857,N_2844);
xor U2901 (N_2901,N_2896,N_2874);
and U2902 (N_2902,N_2813,N_2895);
or U2903 (N_2903,N_2855,N_2808);
nand U2904 (N_2904,N_2882,N_2837);
or U2905 (N_2905,N_2880,N_2864);
xnor U2906 (N_2906,N_2860,N_2873);
or U2907 (N_2907,N_2886,N_2858);
nor U2908 (N_2908,N_2819,N_2823);
nand U2909 (N_2909,N_2821,N_2850);
xnor U2910 (N_2910,N_2817,N_2894);
nor U2911 (N_2911,N_2822,N_2890);
nor U2912 (N_2912,N_2877,N_2828);
nor U2913 (N_2913,N_2851,N_2818);
nor U2914 (N_2914,N_2826,N_2809);
xor U2915 (N_2915,N_2861,N_2842);
nand U2916 (N_2916,N_2846,N_2832);
nor U2917 (N_2917,N_2820,N_2802);
or U2918 (N_2918,N_2854,N_2827);
xnor U2919 (N_2919,N_2806,N_2801);
nor U2920 (N_2920,N_2870,N_2897);
nor U2921 (N_2921,N_2872,N_2899);
or U2922 (N_2922,N_2878,N_2805);
nor U2923 (N_2923,N_2830,N_2881);
and U2924 (N_2924,N_2867,N_2825);
xor U2925 (N_2925,N_2835,N_2856);
nand U2926 (N_2926,N_2833,N_2824);
and U2927 (N_2927,N_2876,N_2814);
nor U2928 (N_2928,N_2865,N_2831);
or U2929 (N_2929,N_2812,N_2853);
and U2930 (N_2930,N_2898,N_2863);
and U2931 (N_2931,N_2843,N_2848);
or U2932 (N_2932,N_2841,N_2811);
and U2933 (N_2933,N_2887,N_2847);
nor U2934 (N_2934,N_2879,N_2829);
or U2935 (N_2935,N_2889,N_2869);
nor U2936 (N_2936,N_2804,N_2815);
and U2937 (N_2937,N_2871,N_2859);
nor U2938 (N_2938,N_2838,N_2885);
or U2939 (N_2939,N_2845,N_2810);
and U2940 (N_2940,N_2866,N_2849);
and U2941 (N_2941,N_2891,N_2888);
xnor U2942 (N_2942,N_2803,N_2862);
nand U2943 (N_2943,N_2868,N_2839);
or U2944 (N_2944,N_2893,N_2875);
and U2945 (N_2945,N_2816,N_2807);
nor U2946 (N_2946,N_2884,N_2883);
or U2947 (N_2947,N_2800,N_2834);
nand U2948 (N_2948,N_2840,N_2892);
nand U2949 (N_2949,N_2836,N_2852);
nor U2950 (N_2950,N_2888,N_2819);
nand U2951 (N_2951,N_2878,N_2826);
and U2952 (N_2952,N_2835,N_2883);
or U2953 (N_2953,N_2893,N_2821);
and U2954 (N_2954,N_2892,N_2842);
or U2955 (N_2955,N_2827,N_2853);
nor U2956 (N_2956,N_2874,N_2876);
nor U2957 (N_2957,N_2889,N_2864);
nor U2958 (N_2958,N_2866,N_2885);
xnor U2959 (N_2959,N_2883,N_2830);
and U2960 (N_2960,N_2818,N_2812);
or U2961 (N_2961,N_2805,N_2800);
and U2962 (N_2962,N_2827,N_2857);
xnor U2963 (N_2963,N_2824,N_2853);
or U2964 (N_2964,N_2821,N_2833);
nand U2965 (N_2965,N_2825,N_2874);
and U2966 (N_2966,N_2821,N_2834);
or U2967 (N_2967,N_2816,N_2867);
nand U2968 (N_2968,N_2821,N_2895);
nor U2969 (N_2969,N_2859,N_2820);
xnor U2970 (N_2970,N_2823,N_2810);
and U2971 (N_2971,N_2837,N_2810);
nand U2972 (N_2972,N_2870,N_2865);
and U2973 (N_2973,N_2804,N_2818);
or U2974 (N_2974,N_2859,N_2869);
nand U2975 (N_2975,N_2812,N_2895);
and U2976 (N_2976,N_2853,N_2870);
and U2977 (N_2977,N_2885,N_2831);
and U2978 (N_2978,N_2851,N_2831);
nor U2979 (N_2979,N_2806,N_2880);
nand U2980 (N_2980,N_2871,N_2883);
xnor U2981 (N_2981,N_2873,N_2898);
nand U2982 (N_2982,N_2810,N_2851);
xnor U2983 (N_2983,N_2844,N_2898);
and U2984 (N_2984,N_2816,N_2811);
and U2985 (N_2985,N_2837,N_2866);
xnor U2986 (N_2986,N_2846,N_2878);
and U2987 (N_2987,N_2888,N_2878);
nor U2988 (N_2988,N_2880,N_2856);
nand U2989 (N_2989,N_2851,N_2893);
nor U2990 (N_2990,N_2854,N_2843);
nor U2991 (N_2991,N_2893,N_2831);
xnor U2992 (N_2992,N_2837,N_2887);
and U2993 (N_2993,N_2808,N_2895);
nand U2994 (N_2994,N_2843,N_2840);
or U2995 (N_2995,N_2815,N_2849);
xor U2996 (N_2996,N_2800,N_2895);
and U2997 (N_2997,N_2878,N_2835);
nand U2998 (N_2998,N_2863,N_2804);
and U2999 (N_2999,N_2808,N_2846);
and U3000 (N_3000,N_2991,N_2920);
nand U3001 (N_3001,N_2921,N_2938);
nor U3002 (N_3002,N_2914,N_2981);
or U3003 (N_3003,N_2937,N_2932);
and U3004 (N_3004,N_2975,N_2901);
xor U3005 (N_3005,N_2979,N_2917);
nor U3006 (N_3006,N_2982,N_2987);
and U3007 (N_3007,N_2942,N_2905);
nor U3008 (N_3008,N_2954,N_2926);
and U3009 (N_3009,N_2971,N_2933);
or U3010 (N_3010,N_2919,N_2997);
nand U3011 (N_3011,N_2963,N_2962);
nor U3012 (N_3012,N_2939,N_2998);
nand U3013 (N_3013,N_2993,N_2951);
xnor U3014 (N_3014,N_2957,N_2949);
nor U3015 (N_3015,N_2911,N_2968);
nand U3016 (N_3016,N_2955,N_2980);
and U3017 (N_3017,N_2970,N_2906);
nor U3018 (N_3018,N_2902,N_2967);
or U3019 (N_3019,N_2913,N_2922);
or U3020 (N_3020,N_2923,N_2928);
xor U3021 (N_3021,N_2908,N_2918);
nand U3022 (N_3022,N_2994,N_2929);
and U3023 (N_3023,N_2960,N_2969);
or U3024 (N_3024,N_2974,N_2988);
nor U3025 (N_3025,N_2977,N_2953);
nand U3026 (N_3026,N_2945,N_2912);
or U3027 (N_3027,N_2989,N_2934);
or U3028 (N_3028,N_2965,N_2999);
or U3029 (N_3029,N_2976,N_2903);
and U3030 (N_3030,N_2940,N_2958);
and U3031 (N_3031,N_2978,N_2946);
nand U3032 (N_3032,N_2935,N_2950);
nand U3033 (N_3033,N_2995,N_2990);
nor U3034 (N_3034,N_2973,N_2956);
and U3035 (N_3035,N_2925,N_2964);
or U3036 (N_3036,N_2916,N_2924);
nand U3037 (N_3037,N_2948,N_2996);
nor U3038 (N_3038,N_2983,N_2947);
nor U3039 (N_3039,N_2936,N_2952);
xnor U3040 (N_3040,N_2909,N_2927);
nor U3041 (N_3041,N_2966,N_2930);
nor U3042 (N_3042,N_2907,N_2986);
and U3043 (N_3043,N_2944,N_2904);
or U3044 (N_3044,N_2972,N_2910);
or U3045 (N_3045,N_2931,N_2985);
nor U3046 (N_3046,N_2941,N_2992);
xnor U3047 (N_3047,N_2961,N_2984);
and U3048 (N_3048,N_2943,N_2959);
nor U3049 (N_3049,N_2915,N_2900);
or U3050 (N_3050,N_2968,N_2913);
nand U3051 (N_3051,N_2984,N_2979);
and U3052 (N_3052,N_2993,N_2912);
nand U3053 (N_3053,N_2902,N_2925);
or U3054 (N_3054,N_2981,N_2928);
xor U3055 (N_3055,N_2929,N_2971);
nand U3056 (N_3056,N_2959,N_2977);
nand U3057 (N_3057,N_2926,N_2956);
and U3058 (N_3058,N_2911,N_2942);
and U3059 (N_3059,N_2987,N_2934);
nand U3060 (N_3060,N_2944,N_2968);
nand U3061 (N_3061,N_2971,N_2901);
nor U3062 (N_3062,N_2919,N_2971);
nor U3063 (N_3063,N_2966,N_2975);
and U3064 (N_3064,N_2911,N_2997);
xnor U3065 (N_3065,N_2995,N_2913);
nor U3066 (N_3066,N_2906,N_2974);
nand U3067 (N_3067,N_2927,N_2989);
or U3068 (N_3068,N_2924,N_2963);
xor U3069 (N_3069,N_2924,N_2978);
nand U3070 (N_3070,N_2997,N_2961);
and U3071 (N_3071,N_2957,N_2994);
xor U3072 (N_3072,N_2906,N_2929);
nor U3073 (N_3073,N_2942,N_2917);
or U3074 (N_3074,N_2923,N_2905);
and U3075 (N_3075,N_2994,N_2956);
and U3076 (N_3076,N_2972,N_2921);
and U3077 (N_3077,N_2987,N_2993);
nor U3078 (N_3078,N_2931,N_2976);
and U3079 (N_3079,N_2924,N_2923);
xnor U3080 (N_3080,N_2969,N_2987);
or U3081 (N_3081,N_2934,N_2955);
and U3082 (N_3082,N_2939,N_2999);
xor U3083 (N_3083,N_2907,N_2927);
nor U3084 (N_3084,N_2995,N_2941);
nand U3085 (N_3085,N_2922,N_2940);
and U3086 (N_3086,N_2900,N_2931);
or U3087 (N_3087,N_2948,N_2969);
nor U3088 (N_3088,N_2952,N_2972);
nand U3089 (N_3089,N_2946,N_2935);
nand U3090 (N_3090,N_2976,N_2982);
and U3091 (N_3091,N_2939,N_2965);
nor U3092 (N_3092,N_2976,N_2983);
xor U3093 (N_3093,N_2962,N_2916);
nand U3094 (N_3094,N_2918,N_2993);
xor U3095 (N_3095,N_2900,N_2948);
nor U3096 (N_3096,N_2955,N_2940);
nor U3097 (N_3097,N_2943,N_2937);
or U3098 (N_3098,N_2947,N_2910);
and U3099 (N_3099,N_2929,N_2909);
nor U3100 (N_3100,N_3005,N_3071);
nand U3101 (N_3101,N_3083,N_3052);
or U3102 (N_3102,N_3028,N_3031);
xnor U3103 (N_3103,N_3084,N_3002);
nor U3104 (N_3104,N_3063,N_3073);
or U3105 (N_3105,N_3012,N_3017);
and U3106 (N_3106,N_3081,N_3075);
nand U3107 (N_3107,N_3007,N_3090);
nand U3108 (N_3108,N_3010,N_3056);
nand U3109 (N_3109,N_3086,N_3016);
nand U3110 (N_3110,N_3003,N_3041);
and U3111 (N_3111,N_3087,N_3000);
nand U3112 (N_3112,N_3051,N_3080);
xnor U3113 (N_3113,N_3036,N_3048);
nor U3114 (N_3114,N_3018,N_3009);
nand U3115 (N_3115,N_3019,N_3085);
and U3116 (N_3116,N_3093,N_3091);
nor U3117 (N_3117,N_3040,N_3059);
xor U3118 (N_3118,N_3029,N_3067);
nand U3119 (N_3119,N_3096,N_3047);
nand U3120 (N_3120,N_3054,N_3094);
or U3121 (N_3121,N_3092,N_3082);
xnor U3122 (N_3122,N_3057,N_3035);
or U3123 (N_3123,N_3070,N_3050);
nor U3124 (N_3124,N_3004,N_3033);
nor U3125 (N_3125,N_3039,N_3034);
or U3126 (N_3126,N_3088,N_3023);
and U3127 (N_3127,N_3065,N_3030);
xor U3128 (N_3128,N_3032,N_3058);
nor U3129 (N_3129,N_3072,N_3022);
nand U3130 (N_3130,N_3079,N_3025);
nand U3131 (N_3131,N_3024,N_3045);
nor U3132 (N_3132,N_3001,N_3069);
or U3133 (N_3133,N_3055,N_3068);
or U3134 (N_3134,N_3049,N_3013);
and U3135 (N_3135,N_3061,N_3021);
nor U3136 (N_3136,N_3060,N_3074);
and U3137 (N_3137,N_3089,N_3043);
nor U3138 (N_3138,N_3006,N_3044);
nand U3139 (N_3139,N_3042,N_3078);
and U3140 (N_3140,N_3064,N_3046);
nand U3141 (N_3141,N_3008,N_3027);
xor U3142 (N_3142,N_3014,N_3095);
and U3143 (N_3143,N_3098,N_3076);
or U3144 (N_3144,N_3020,N_3099);
and U3145 (N_3145,N_3011,N_3062);
nand U3146 (N_3146,N_3077,N_3026);
or U3147 (N_3147,N_3066,N_3037);
nand U3148 (N_3148,N_3038,N_3097);
nand U3149 (N_3149,N_3053,N_3015);
nand U3150 (N_3150,N_3058,N_3071);
nor U3151 (N_3151,N_3015,N_3060);
nand U3152 (N_3152,N_3008,N_3004);
nor U3153 (N_3153,N_3013,N_3088);
and U3154 (N_3154,N_3074,N_3021);
nand U3155 (N_3155,N_3010,N_3014);
nor U3156 (N_3156,N_3030,N_3026);
and U3157 (N_3157,N_3060,N_3076);
and U3158 (N_3158,N_3066,N_3042);
and U3159 (N_3159,N_3021,N_3085);
or U3160 (N_3160,N_3030,N_3066);
and U3161 (N_3161,N_3079,N_3064);
or U3162 (N_3162,N_3089,N_3003);
and U3163 (N_3163,N_3050,N_3028);
nand U3164 (N_3164,N_3055,N_3035);
nor U3165 (N_3165,N_3028,N_3026);
nor U3166 (N_3166,N_3081,N_3024);
and U3167 (N_3167,N_3097,N_3051);
and U3168 (N_3168,N_3017,N_3030);
nand U3169 (N_3169,N_3042,N_3098);
or U3170 (N_3170,N_3085,N_3020);
and U3171 (N_3171,N_3013,N_3045);
or U3172 (N_3172,N_3053,N_3081);
and U3173 (N_3173,N_3063,N_3018);
and U3174 (N_3174,N_3031,N_3047);
nor U3175 (N_3175,N_3054,N_3008);
nand U3176 (N_3176,N_3048,N_3073);
or U3177 (N_3177,N_3094,N_3059);
and U3178 (N_3178,N_3005,N_3033);
nand U3179 (N_3179,N_3067,N_3063);
nand U3180 (N_3180,N_3034,N_3083);
or U3181 (N_3181,N_3093,N_3098);
and U3182 (N_3182,N_3054,N_3095);
or U3183 (N_3183,N_3055,N_3007);
nand U3184 (N_3184,N_3008,N_3046);
xnor U3185 (N_3185,N_3064,N_3056);
nor U3186 (N_3186,N_3058,N_3099);
nor U3187 (N_3187,N_3005,N_3068);
nor U3188 (N_3188,N_3097,N_3087);
nor U3189 (N_3189,N_3065,N_3010);
or U3190 (N_3190,N_3028,N_3066);
nor U3191 (N_3191,N_3035,N_3091);
and U3192 (N_3192,N_3008,N_3096);
xnor U3193 (N_3193,N_3048,N_3080);
nor U3194 (N_3194,N_3004,N_3063);
nand U3195 (N_3195,N_3004,N_3020);
and U3196 (N_3196,N_3081,N_3015);
and U3197 (N_3197,N_3002,N_3060);
nand U3198 (N_3198,N_3046,N_3079);
nand U3199 (N_3199,N_3034,N_3068);
and U3200 (N_3200,N_3105,N_3176);
nor U3201 (N_3201,N_3151,N_3150);
or U3202 (N_3202,N_3101,N_3132);
nor U3203 (N_3203,N_3117,N_3186);
and U3204 (N_3204,N_3153,N_3193);
nor U3205 (N_3205,N_3164,N_3166);
nor U3206 (N_3206,N_3115,N_3160);
or U3207 (N_3207,N_3103,N_3171);
nand U3208 (N_3208,N_3125,N_3179);
or U3209 (N_3209,N_3192,N_3128);
and U3210 (N_3210,N_3118,N_3144);
and U3211 (N_3211,N_3162,N_3121);
xnor U3212 (N_3212,N_3134,N_3116);
nor U3213 (N_3213,N_3188,N_3114);
nand U3214 (N_3214,N_3163,N_3161);
nand U3215 (N_3215,N_3167,N_3122);
and U3216 (N_3216,N_3108,N_3185);
nand U3217 (N_3217,N_3159,N_3123);
and U3218 (N_3218,N_3145,N_3109);
nand U3219 (N_3219,N_3180,N_3170);
or U3220 (N_3220,N_3168,N_3199);
nor U3221 (N_3221,N_3102,N_3106);
nor U3222 (N_3222,N_3195,N_3182);
nand U3223 (N_3223,N_3107,N_3181);
nor U3224 (N_3224,N_3157,N_3198);
xor U3225 (N_3225,N_3183,N_3131);
and U3226 (N_3226,N_3177,N_3154);
nor U3227 (N_3227,N_3174,N_3104);
and U3228 (N_3228,N_3156,N_3135);
or U3229 (N_3229,N_3148,N_3137);
and U3230 (N_3230,N_3189,N_3158);
and U3231 (N_3231,N_3165,N_3112);
nor U3232 (N_3232,N_3173,N_3155);
nor U3233 (N_3233,N_3133,N_3130);
or U3234 (N_3234,N_3172,N_3147);
xor U3235 (N_3235,N_3152,N_3178);
nor U3236 (N_3236,N_3191,N_3169);
nand U3237 (N_3237,N_3197,N_3100);
and U3238 (N_3238,N_3126,N_3110);
or U3239 (N_3239,N_3194,N_3111);
nor U3240 (N_3240,N_3119,N_3127);
nand U3241 (N_3241,N_3190,N_3184);
or U3242 (N_3242,N_3140,N_3113);
nor U3243 (N_3243,N_3143,N_3142);
nand U3244 (N_3244,N_3124,N_3141);
nand U3245 (N_3245,N_3146,N_3187);
nand U3246 (N_3246,N_3136,N_3139);
and U3247 (N_3247,N_3196,N_3138);
nand U3248 (N_3248,N_3129,N_3175);
xnor U3249 (N_3249,N_3120,N_3149);
nand U3250 (N_3250,N_3111,N_3106);
nor U3251 (N_3251,N_3119,N_3173);
nor U3252 (N_3252,N_3111,N_3110);
nand U3253 (N_3253,N_3130,N_3184);
nand U3254 (N_3254,N_3163,N_3173);
nor U3255 (N_3255,N_3169,N_3133);
xor U3256 (N_3256,N_3120,N_3107);
and U3257 (N_3257,N_3127,N_3197);
nand U3258 (N_3258,N_3139,N_3162);
or U3259 (N_3259,N_3193,N_3166);
nor U3260 (N_3260,N_3128,N_3132);
and U3261 (N_3261,N_3143,N_3127);
or U3262 (N_3262,N_3125,N_3141);
nand U3263 (N_3263,N_3112,N_3102);
or U3264 (N_3264,N_3182,N_3162);
xor U3265 (N_3265,N_3195,N_3104);
and U3266 (N_3266,N_3102,N_3128);
nand U3267 (N_3267,N_3135,N_3107);
nor U3268 (N_3268,N_3178,N_3183);
xnor U3269 (N_3269,N_3113,N_3126);
and U3270 (N_3270,N_3127,N_3123);
or U3271 (N_3271,N_3113,N_3118);
and U3272 (N_3272,N_3130,N_3189);
nor U3273 (N_3273,N_3142,N_3146);
and U3274 (N_3274,N_3160,N_3196);
or U3275 (N_3275,N_3142,N_3101);
or U3276 (N_3276,N_3150,N_3115);
or U3277 (N_3277,N_3134,N_3153);
nor U3278 (N_3278,N_3131,N_3189);
and U3279 (N_3279,N_3104,N_3103);
nor U3280 (N_3280,N_3171,N_3175);
xor U3281 (N_3281,N_3158,N_3136);
nand U3282 (N_3282,N_3185,N_3191);
or U3283 (N_3283,N_3136,N_3120);
nor U3284 (N_3284,N_3165,N_3168);
xor U3285 (N_3285,N_3154,N_3199);
or U3286 (N_3286,N_3123,N_3177);
nand U3287 (N_3287,N_3154,N_3117);
nand U3288 (N_3288,N_3150,N_3103);
or U3289 (N_3289,N_3196,N_3159);
xor U3290 (N_3290,N_3190,N_3107);
or U3291 (N_3291,N_3186,N_3175);
nand U3292 (N_3292,N_3163,N_3113);
nor U3293 (N_3293,N_3184,N_3188);
or U3294 (N_3294,N_3139,N_3188);
or U3295 (N_3295,N_3101,N_3143);
or U3296 (N_3296,N_3147,N_3112);
nand U3297 (N_3297,N_3168,N_3104);
or U3298 (N_3298,N_3184,N_3107);
or U3299 (N_3299,N_3134,N_3136);
and U3300 (N_3300,N_3227,N_3285);
nand U3301 (N_3301,N_3218,N_3272);
nand U3302 (N_3302,N_3252,N_3271);
nor U3303 (N_3303,N_3261,N_3265);
xor U3304 (N_3304,N_3291,N_3266);
nand U3305 (N_3305,N_3247,N_3242);
or U3306 (N_3306,N_3290,N_3208);
or U3307 (N_3307,N_3287,N_3207);
and U3308 (N_3308,N_3296,N_3228);
nand U3309 (N_3309,N_3213,N_3256);
nand U3310 (N_3310,N_3230,N_3225);
nor U3311 (N_3311,N_3248,N_3257);
nand U3312 (N_3312,N_3221,N_3212);
nor U3313 (N_3313,N_3243,N_3286);
and U3314 (N_3314,N_3281,N_3202);
nand U3315 (N_3315,N_3299,N_3220);
or U3316 (N_3316,N_3206,N_3253);
nand U3317 (N_3317,N_3264,N_3293);
or U3318 (N_3318,N_3275,N_3283);
or U3319 (N_3319,N_3284,N_3236);
or U3320 (N_3320,N_3232,N_3269);
or U3321 (N_3321,N_3240,N_3260);
xnor U3322 (N_3322,N_3280,N_3274);
or U3323 (N_3323,N_3282,N_3262);
and U3324 (N_3324,N_3210,N_3238);
nand U3325 (N_3325,N_3263,N_3211);
or U3326 (N_3326,N_3209,N_3294);
and U3327 (N_3327,N_3259,N_3216);
nor U3328 (N_3328,N_3295,N_3203);
nor U3329 (N_3329,N_3251,N_3223);
nand U3330 (N_3330,N_3279,N_3222);
xor U3331 (N_3331,N_3241,N_3292);
or U3332 (N_3332,N_3219,N_3215);
or U3333 (N_3333,N_3201,N_3249);
or U3334 (N_3334,N_3204,N_3278);
or U3335 (N_3335,N_3245,N_3233);
or U3336 (N_3336,N_3200,N_3270);
xor U3337 (N_3337,N_3239,N_3255);
nand U3338 (N_3338,N_3217,N_3288);
nor U3339 (N_3339,N_3258,N_3229);
nand U3340 (N_3340,N_3250,N_3231);
and U3341 (N_3341,N_3205,N_3276);
or U3342 (N_3342,N_3298,N_3237);
nand U3343 (N_3343,N_3235,N_3224);
or U3344 (N_3344,N_3244,N_3268);
or U3345 (N_3345,N_3289,N_3234);
xnor U3346 (N_3346,N_3273,N_3267);
or U3347 (N_3347,N_3214,N_3297);
nand U3348 (N_3348,N_3254,N_3246);
nor U3349 (N_3349,N_3226,N_3277);
and U3350 (N_3350,N_3245,N_3246);
or U3351 (N_3351,N_3268,N_3281);
nor U3352 (N_3352,N_3285,N_3229);
and U3353 (N_3353,N_3260,N_3291);
nor U3354 (N_3354,N_3251,N_3219);
and U3355 (N_3355,N_3273,N_3271);
and U3356 (N_3356,N_3247,N_3285);
and U3357 (N_3357,N_3257,N_3267);
xnor U3358 (N_3358,N_3227,N_3273);
nand U3359 (N_3359,N_3251,N_3228);
nor U3360 (N_3360,N_3249,N_3292);
and U3361 (N_3361,N_3288,N_3253);
or U3362 (N_3362,N_3279,N_3235);
nor U3363 (N_3363,N_3239,N_3205);
nor U3364 (N_3364,N_3200,N_3218);
or U3365 (N_3365,N_3214,N_3254);
or U3366 (N_3366,N_3253,N_3274);
and U3367 (N_3367,N_3231,N_3208);
and U3368 (N_3368,N_3220,N_3233);
nor U3369 (N_3369,N_3208,N_3227);
or U3370 (N_3370,N_3229,N_3263);
or U3371 (N_3371,N_3211,N_3288);
xnor U3372 (N_3372,N_3236,N_3210);
nand U3373 (N_3373,N_3287,N_3260);
and U3374 (N_3374,N_3211,N_3213);
nor U3375 (N_3375,N_3257,N_3243);
or U3376 (N_3376,N_3276,N_3230);
nor U3377 (N_3377,N_3233,N_3264);
xor U3378 (N_3378,N_3269,N_3231);
nand U3379 (N_3379,N_3215,N_3229);
and U3380 (N_3380,N_3235,N_3230);
nor U3381 (N_3381,N_3240,N_3264);
and U3382 (N_3382,N_3234,N_3263);
nor U3383 (N_3383,N_3291,N_3200);
nor U3384 (N_3384,N_3261,N_3238);
nor U3385 (N_3385,N_3242,N_3283);
nand U3386 (N_3386,N_3295,N_3299);
nor U3387 (N_3387,N_3226,N_3231);
and U3388 (N_3388,N_3230,N_3271);
nor U3389 (N_3389,N_3218,N_3217);
nand U3390 (N_3390,N_3243,N_3295);
or U3391 (N_3391,N_3292,N_3289);
and U3392 (N_3392,N_3207,N_3268);
and U3393 (N_3393,N_3282,N_3268);
nand U3394 (N_3394,N_3239,N_3232);
nor U3395 (N_3395,N_3292,N_3217);
and U3396 (N_3396,N_3263,N_3260);
or U3397 (N_3397,N_3218,N_3221);
nand U3398 (N_3398,N_3210,N_3272);
nand U3399 (N_3399,N_3207,N_3202);
and U3400 (N_3400,N_3394,N_3355);
nand U3401 (N_3401,N_3376,N_3343);
or U3402 (N_3402,N_3349,N_3374);
nor U3403 (N_3403,N_3337,N_3361);
xor U3404 (N_3404,N_3371,N_3306);
and U3405 (N_3405,N_3388,N_3399);
and U3406 (N_3406,N_3300,N_3304);
nand U3407 (N_3407,N_3312,N_3354);
nand U3408 (N_3408,N_3327,N_3366);
nand U3409 (N_3409,N_3334,N_3310);
and U3410 (N_3410,N_3369,N_3329);
xnor U3411 (N_3411,N_3314,N_3379);
nor U3412 (N_3412,N_3356,N_3338);
nand U3413 (N_3413,N_3317,N_3320);
or U3414 (N_3414,N_3363,N_3389);
nand U3415 (N_3415,N_3307,N_3392);
or U3416 (N_3416,N_3345,N_3383);
or U3417 (N_3417,N_3302,N_3393);
or U3418 (N_3418,N_3336,N_3321);
and U3419 (N_3419,N_3378,N_3368);
nor U3420 (N_3420,N_3390,N_3347);
or U3421 (N_3421,N_3372,N_3359);
or U3422 (N_3422,N_3311,N_3331);
xor U3423 (N_3423,N_3332,N_3301);
and U3424 (N_3424,N_3330,N_3396);
xor U3425 (N_3425,N_3391,N_3380);
xor U3426 (N_3426,N_3348,N_3364);
or U3427 (N_3427,N_3365,N_3386);
and U3428 (N_3428,N_3344,N_3322);
or U3429 (N_3429,N_3353,N_3362);
nand U3430 (N_3430,N_3340,N_3382);
xor U3431 (N_3431,N_3360,N_3381);
or U3432 (N_3432,N_3323,N_3342);
or U3433 (N_3433,N_3324,N_3316);
nand U3434 (N_3434,N_3352,N_3325);
nor U3435 (N_3435,N_3397,N_3319);
nor U3436 (N_3436,N_3309,N_3350);
nor U3437 (N_3437,N_3385,N_3313);
or U3438 (N_3438,N_3333,N_3387);
or U3439 (N_3439,N_3335,N_3328);
nor U3440 (N_3440,N_3308,N_3384);
or U3441 (N_3441,N_3315,N_3358);
or U3442 (N_3442,N_3339,N_3398);
nor U3443 (N_3443,N_3303,N_3346);
or U3444 (N_3444,N_3341,N_3377);
and U3445 (N_3445,N_3373,N_3375);
nor U3446 (N_3446,N_3305,N_3370);
nand U3447 (N_3447,N_3367,N_3395);
nand U3448 (N_3448,N_3318,N_3351);
xor U3449 (N_3449,N_3326,N_3357);
or U3450 (N_3450,N_3389,N_3396);
nand U3451 (N_3451,N_3368,N_3336);
nand U3452 (N_3452,N_3312,N_3320);
and U3453 (N_3453,N_3391,N_3312);
nor U3454 (N_3454,N_3302,N_3389);
nor U3455 (N_3455,N_3354,N_3360);
or U3456 (N_3456,N_3336,N_3367);
nor U3457 (N_3457,N_3338,N_3315);
and U3458 (N_3458,N_3395,N_3380);
and U3459 (N_3459,N_3349,N_3348);
nand U3460 (N_3460,N_3326,N_3319);
nor U3461 (N_3461,N_3344,N_3345);
and U3462 (N_3462,N_3380,N_3309);
and U3463 (N_3463,N_3377,N_3356);
xor U3464 (N_3464,N_3338,N_3371);
nor U3465 (N_3465,N_3386,N_3370);
nand U3466 (N_3466,N_3325,N_3329);
nand U3467 (N_3467,N_3316,N_3333);
or U3468 (N_3468,N_3372,N_3363);
or U3469 (N_3469,N_3335,N_3322);
nor U3470 (N_3470,N_3376,N_3300);
or U3471 (N_3471,N_3342,N_3307);
nor U3472 (N_3472,N_3301,N_3358);
or U3473 (N_3473,N_3371,N_3353);
or U3474 (N_3474,N_3324,N_3376);
xnor U3475 (N_3475,N_3391,N_3332);
nor U3476 (N_3476,N_3334,N_3376);
xor U3477 (N_3477,N_3358,N_3378);
or U3478 (N_3478,N_3343,N_3397);
nand U3479 (N_3479,N_3399,N_3319);
or U3480 (N_3480,N_3337,N_3336);
nor U3481 (N_3481,N_3374,N_3356);
or U3482 (N_3482,N_3300,N_3348);
xor U3483 (N_3483,N_3394,N_3310);
or U3484 (N_3484,N_3369,N_3339);
or U3485 (N_3485,N_3307,N_3388);
and U3486 (N_3486,N_3302,N_3387);
or U3487 (N_3487,N_3314,N_3393);
and U3488 (N_3488,N_3334,N_3301);
nand U3489 (N_3489,N_3371,N_3341);
nor U3490 (N_3490,N_3358,N_3321);
and U3491 (N_3491,N_3383,N_3380);
nor U3492 (N_3492,N_3376,N_3308);
nor U3493 (N_3493,N_3382,N_3383);
or U3494 (N_3494,N_3333,N_3393);
nand U3495 (N_3495,N_3348,N_3366);
or U3496 (N_3496,N_3311,N_3322);
nand U3497 (N_3497,N_3315,N_3388);
nand U3498 (N_3498,N_3328,N_3382);
nand U3499 (N_3499,N_3382,N_3341);
and U3500 (N_3500,N_3491,N_3487);
or U3501 (N_3501,N_3432,N_3435);
nor U3502 (N_3502,N_3482,N_3489);
nor U3503 (N_3503,N_3443,N_3472);
nor U3504 (N_3504,N_3493,N_3463);
and U3505 (N_3505,N_3466,N_3430);
or U3506 (N_3506,N_3429,N_3457);
or U3507 (N_3507,N_3448,N_3461);
and U3508 (N_3508,N_3428,N_3407);
nor U3509 (N_3509,N_3476,N_3445);
and U3510 (N_3510,N_3437,N_3498);
nand U3511 (N_3511,N_3416,N_3492);
xor U3512 (N_3512,N_3483,N_3409);
or U3513 (N_3513,N_3488,N_3486);
or U3514 (N_3514,N_3431,N_3454);
xnor U3515 (N_3515,N_3411,N_3494);
and U3516 (N_3516,N_3497,N_3405);
nand U3517 (N_3517,N_3421,N_3480);
xnor U3518 (N_3518,N_3420,N_3406);
and U3519 (N_3519,N_3485,N_3475);
xnor U3520 (N_3520,N_3478,N_3477);
and U3521 (N_3521,N_3417,N_3419);
nand U3522 (N_3522,N_3455,N_3499);
and U3523 (N_3523,N_3460,N_3400);
nor U3524 (N_3524,N_3462,N_3456);
or U3525 (N_3525,N_3414,N_3402);
or U3526 (N_3526,N_3444,N_3458);
and U3527 (N_3527,N_3452,N_3439);
nor U3528 (N_3528,N_3474,N_3408);
or U3529 (N_3529,N_3418,N_3410);
or U3530 (N_3530,N_3401,N_3451);
or U3531 (N_3531,N_3479,N_3413);
and U3532 (N_3532,N_3422,N_3436);
nand U3533 (N_3533,N_3434,N_3467);
and U3534 (N_3534,N_3441,N_3459);
nor U3535 (N_3535,N_3481,N_3425);
nand U3536 (N_3536,N_3469,N_3426);
or U3537 (N_3537,N_3496,N_3447);
xnor U3538 (N_3538,N_3424,N_3465);
or U3539 (N_3539,N_3470,N_3415);
and U3540 (N_3540,N_3495,N_3446);
xnor U3541 (N_3541,N_3427,N_3449);
and U3542 (N_3542,N_3453,N_3438);
nand U3543 (N_3543,N_3468,N_3404);
nand U3544 (N_3544,N_3464,N_3450);
xor U3545 (N_3545,N_3403,N_3440);
and U3546 (N_3546,N_3490,N_3433);
xor U3547 (N_3547,N_3471,N_3412);
or U3548 (N_3548,N_3473,N_3484);
or U3549 (N_3549,N_3423,N_3442);
nor U3550 (N_3550,N_3416,N_3496);
and U3551 (N_3551,N_3488,N_3466);
xnor U3552 (N_3552,N_3490,N_3459);
nand U3553 (N_3553,N_3435,N_3458);
xor U3554 (N_3554,N_3469,N_3465);
or U3555 (N_3555,N_3432,N_3417);
xor U3556 (N_3556,N_3412,N_3486);
or U3557 (N_3557,N_3468,N_3469);
nand U3558 (N_3558,N_3428,N_3478);
or U3559 (N_3559,N_3474,N_3441);
nor U3560 (N_3560,N_3445,N_3479);
nor U3561 (N_3561,N_3477,N_3407);
and U3562 (N_3562,N_3420,N_3412);
nand U3563 (N_3563,N_3477,N_3450);
nand U3564 (N_3564,N_3440,N_3492);
nand U3565 (N_3565,N_3476,N_3462);
or U3566 (N_3566,N_3438,N_3456);
nor U3567 (N_3567,N_3404,N_3474);
and U3568 (N_3568,N_3406,N_3405);
nand U3569 (N_3569,N_3472,N_3459);
nor U3570 (N_3570,N_3414,N_3440);
nor U3571 (N_3571,N_3467,N_3420);
nand U3572 (N_3572,N_3407,N_3491);
nand U3573 (N_3573,N_3418,N_3495);
nand U3574 (N_3574,N_3493,N_3414);
or U3575 (N_3575,N_3498,N_3404);
and U3576 (N_3576,N_3423,N_3403);
nand U3577 (N_3577,N_3447,N_3464);
and U3578 (N_3578,N_3449,N_3461);
xnor U3579 (N_3579,N_3448,N_3432);
and U3580 (N_3580,N_3448,N_3486);
nand U3581 (N_3581,N_3425,N_3432);
nand U3582 (N_3582,N_3454,N_3467);
nor U3583 (N_3583,N_3421,N_3427);
and U3584 (N_3584,N_3472,N_3484);
nor U3585 (N_3585,N_3404,N_3460);
or U3586 (N_3586,N_3434,N_3496);
or U3587 (N_3587,N_3496,N_3450);
nand U3588 (N_3588,N_3426,N_3441);
and U3589 (N_3589,N_3407,N_3418);
or U3590 (N_3590,N_3480,N_3466);
and U3591 (N_3591,N_3467,N_3487);
xnor U3592 (N_3592,N_3469,N_3401);
and U3593 (N_3593,N_3460,N_3482);
nor U3594 (N_3594,N_3461,N_3408);
and U3595 (N_3595,N_3411,N_3402);
and U3596 (N_3596,N_3469,N_3410);
or U3597 (N_3597,N_3490,N_3447);
xnor U3598 (N_3598,N_3440,N_3465);
nand U3599 (N_3599,N_3462,N_3443);
and U3600 (N_3600,N_3507,N_3591);
or U3601 (N_3601,N_3576,N_3557);
nand U3602 (N_3602,N_3548,N_3519);
and U3603 (N_3603,N_3593,N_3518);
or U3604 (N_3604,N_3559,N_3555);
or U3605 (N_3605,N_3570,N_3586);
and U3606 (N_3606,N_3537,N_3522);
or U3607 (N_3607,N_3592,N_3534);
and U3608 (N_3608,N_3565,N_3514);
and U3609 (N_3609,N_3530,N_3533);
and U3610 (N_3610,N_3516,N_3567);
or U3611 (N_3611,N_3595,N_3525);
and U3612 (N_3612,N_3573,N_3552);
nor U3613 (N_3613,N_3503,N_3540);
or U3614 (N_3614,N_3523,N_3582);
nand U3615 (N_3615,N_3572,N_3521);
nor U3616 (N_3616,N_3527,N_3532);
or U3617 (N_3617,N_3583,N_3554);
nand U3618 (N_3618,N_3538,N_3505);
and U3619 (N_3619,N_3547,N_3551);
and U3620 (N_3620,N_3571,N_3528);
and U3621 (N_3621,N_3597,N_3531);
and U3622 (N_3622,N_3561,N_3590);
and U3623 (N_3623,N_3520,N_3545);
xnor U3624 (N_3624,N_3506,N_3524);
nand U3625 (N_3625,N_3543,N_3558);
or U3626 (N_3626,N_3563,N_3584);
nor U3627 (N_3627,N_3585,N_3580);
and U3628 (N_3628,N_3535,N_3536);
nand U3629 (N_3629,N_3549,N_3553);
or U3630 (N_3630,N_3542,N_3579);
nand U3631 (N_3631,N_3574,N_3529);
and U3632 (N_3632,N_3596,N_3581);
xnor U3633 (N_3633,N_3509,N_3599);
nand U3634 (N_3634,N_3504,N_3566);
xnor U3635 (N_3635,N_3517,N_3589);
and U3636 (N_3636,N_3511,N_3510);
or U3637 (N_3637,N_3569,N_3598);
nor U3638 (N_3638,N_3560,N_3502);
nand U3639 (N_3639,N_3578,N_3515);
or U3640 (N_3640,N_3577,N_3546);
nor U3641 (N_3641,N_3588,N_3501);
nand U3642 (N_3642,N_3526,N_3556);
nor U3643 (N_3643,N_3508,N_3568);
or U3644 (N_3644,N_3564,N_3513);
nand U3645 (N_3645,N_3550,N_3544);
or U3646 (N_3646,N_3539,N_3541);
and U3647 (N_3647,N_3512,N_3500);
and U3648 (N_3648,N_3594,N_3562);
nor U3649 (N_3649,N_3575,N_3587);
nor U3650 (N_3650,N_3551,N_3507);
xnor U3651 (N_3651,N_3590,N_3534);
nor U3652 (N_3652,N_3582,N_3514);
or U3653 (N_3653,N_3582,N_3566);
or U3654 (N_3654,N_3563,N_3583);
nand U3655 (N_3655,N_3510,N_3537);
or U3656 (N_3656,N_3523,N_3519);
or U3657 (N_3657,N_3519,N_3591);
and U3658 (N_3658,N_3587,N_3588);
or U3659 (N_3659,N_3596,N_3598);
or U3660 (N_3660,N_3579,N_3509);
or U3661 (N_3661,N_3580,N_3512);
or U3662 (N_3662,N_3536,N_3525);
nand U3663 (N_3663,N_3549,N_3513);
and U3664 (N_3664,N_3554,N_3532);
and U3665 (N_3665,N_3538,N_3572);
xnor U3666 (N_3666,N_3530,N_3579);
or U3667 (N_3667,N_3508,N_3546);
nor U3668 (N_3668,N_3585,N_3511);
nor U3669 (N_3669,N_3573,N_3570);
or U3670 (N_3670,N_3557,N_3587);
nand U3671 (N_3671,N_3592,N_3590);
and U3672 (N_3672,N_3572,N_3518);
nand U3673 (N_3673,N_3543,N_3534);
nor U3674 (N_3674,N_3567,N_3513);
and U3675 (N_3675,N_3589,N_3551);
and U3676 (N_3676,N_3526,N_3576);
and U3677 (N_3677,N_3501,N_3594);
or U3678 (N_3678,N_3554,N_3516);
or U3679 (N_3679,N_3597,N_3542);
xor U3680 (N_3680,N_3590,N_3571);
nand U3681 (N_3681,N_3535,N_3576);
nand U3682 (N_3682,N_3501,N_3591);
nor U3683 (N_3683,N_3594,N_3566);
and U3684 (N_3684,N_3562,N_3505);
xnor U3685 (N_3685,N_3583,N_3523);
nor U3686 (N_3686,N_3548,N_3589);
nor U3687 (N_3687,N_3581,N_3574);
or U3688 (N_3688,N_3517,N_3574);
nand U3689 (N_3689,N_3544,N_3532);
and U3690 (N_3690,N_3564,N_3549);
xnor U3691 (N_3691,N_3523,N_3526);
or U3692 (N_3692,N_3573,N_3567);
or U3693 (N_3693,N_3550,N_3596);
or U3694 (N_3694,N_3501,N_3561);
nor U3695 (N_3695,N_3557,N_3571);
nor U3696 (N_3696,N_3539,N_3513);
nor U3697 (N_3697,N_3502,N_3575);
or U3698 (N_3698,N_3553,N_3556);
and U3699 (N_3699,N_3531,N_3510);
and U3700 (N_3700,N_3666,N_3650);
and U3701 (N_3701,N_3680,N_3603);
nand U3702 (N_3702,N_3668,N_3627);
xnor U3703 (N_3703,N_3679,N_3667);
or U3704 (N_3704,N_3678,N_3618);
and U3705 (N_3705,N_3670,N_3631);
and U3706 (N_3706,N_3672,N_3608);
or U3707 (N_3707,N_3693,N_3674);
nand U3708 (N_3708,N_3636,N_3632);
nand U3709 (N_3709,N_3614,N_3663);
nand U3710 (N_3710,N_3626,N_3613);
and U3711 (N_3711,N_3600,N_3683);
and U3712 (N_3712,N_3620,N_3684);
nand U3713 (N_3713,N_3610,N_3639);
and U3714 (N_3714,N_3675,N_3662);
or U3715 (N_3715,N_3628,N_3697);
nand U3716 (N_3716,N_3681,N_3698);
or U3717 (N_3717,N_3685,N_3689);
and U3718 (N_3718,N_3602,N_3601);
and U3719 (N_3719,N_3615,N_3690);
nor U3720 (N_3720,N_3621,N_3676);
and U3721 (N_3721,N_3664,N_3637);
nand U3722 (N_3722,N_3606,N_3629);
nor U3723 (N_3723,N_3607,N_3633);
or U3724 (N_3724,N_3604,N_3695);
nor U3725 (N_3725,N_3655,N_3635);
nor U3726 (N_3726,N_3665,N_3696);
nand U3727 (N_3727,N_3643,N_3611);
and U3728 (N_3728,N_3651,N_3656);
nor U3729 (N_3729,N_3619,N_3699);
or U3730 (N_3730,N_3646,N_3673);
nand U3731 (N_3731,N_3612,N_3653);
or U3732 (N_3732,N_3661,N_3645);
nor U3733 (N_3733,N_3657,N_3649);
nor U3734 (N_3734,N_3634,N_3671);
nand U3735 (N_3735,N_3624,N_3625);
nand U3736 (N_3736,N_3640,N_3644);
or U3737 (N_3737,N_3660,N_3642);
xnor U3738 (N_3738,N_3682,N_3641);
nand U3739 (N_3739,N_3686,N_3677);
or U3740 (N_3740,N_3694,N_3659);
nor U3741 (N_3741,N_3609,N_3669);
nand U3742 (N_3742,N_3658,N_3605);
and U3743 (N_3743,N_3647,N_3691);
nand U3744 (N_3744,N_3616,N_3692);
or U3745 (N_3745,N_3622,N_3638);
and U3746 (N_3746,N_3617,N_3688);
or U3747 (N_3747,N_3630,N_3648);
xor U3748 (N_3748,N_3654,N_3652);
nand U3749 (N_3749,N_3687,N_3623);
nor U3750 (N_3750,N_3600,N_3670);
and U3751 (N_3751,N_3663,N_3659);
nand U3752 (N_3752,N_3655,N_3664);
nor U3753 (N_3753,N_3628,N_3656);
or U3754 (N_3754,N_3681,N_3663);
and U3755 (N_3755,N_3635,N_3633);
nand U3756 (N_3756,N_3608,N_3602);
or U3757 (N_3757,N_3623,N_3667);
nor U3758 (N_3758,N_3616,N_3678);
or U3759 (N_3759,N_3678,N_3657);
and U3760 (N_3760,N_3691,N_3666);
xor U3761 (N_3761,N_3648,N_3662);
xnor U3762 (N_3762,N_3647,N_3657);
nor U3763 (N_3763,N_3656,N_3698);
and U3764 (N_3764,N_3640,N_3600);
or U3765 (N_3765,N_3615,N_3618);
and U3766 (N_3766,N_3669,N_3675);
xnor U3767 (N_3767,N_3630,N_3644);
and U3768 (N_3768,N_3655,N_3684);
or U3769 (N_3769,N_3674,N_3665);
xor U3770 (N_3770,N_3653,N_3623);
nand U3771 (N_3771,N_3669,N_3661);
nand U3772 (N_3772,N_3625,N_3626);
or U3773 (N_3773,N_3654,N_3677);
or U3774 (N_3774,N_3682,N_3642);
xor U3775 (N_3775,N_3689,N_3643);
nor U3776 (N_3776,N_3661,N_3607);
nor U3777 (N_3777,N_3602,N_3647);
nand U3778 (N_3778,N_3648,N_3602);
and U3779 (N_3779,N_3688,N_3610);
and U3780 (N_3780,N_3680,N_3652);
nand U3781 (N_3781,N_3668,N_3693);
nor U3782 (N_3782,N_3658,N_3618);
xor U3783 (N_3783,N_3612,N_3635);
nand U3784 (N_3784,N_3613,N_3683);
and U3785 (N_3785,N_3675,N_3617);
or U3786 (N_3786,N_3601,N_3635);
nor U3787 (N_3787,N_3636,N_3658);
nand U3788 (N_3788,N_3629,N_3608);
nor U3789 (N_3789,N_3683,N_3602);
nand U3790 (N_3790,N_3621,N_3604);
and U3791 (N_3791,N_3606,N_3631);
or U3792 (N_3792,N_3669,N_3648);
nand U3793 (N_3793,N_3634,N_3640);
nor U3794 (N_3794,N_3699,N_3666);
xnor U3795 (N_3795,N_3602,N_3672);
and U3796 (N_3796,N_3605,N_3664);
nand U3797 (N_3797,N_3604,N_3661);
nor U3798 (N_3798,N_3670,N_3645);
nor U3799 (N_3799,N_3675,N_3688);
or U3800 (N_3800,N_3749,N_3768);
nor U3801 (N_3801,N_3777,N_3706);
and U3802 (N_3802,N_3751,N_3782);
nor U3803 (N_3803,N_3721,N_3735);
xor U3804 (N_3804,N_3704,N_3707);
and U3805 (N_3805,N_3755,N_3718);
or U3806 (N_3806,N_3795,N_3779);
or U3807 (N_3807,N_3781,N_3709);
or U3808 (N_3808,N_3731,N_3712);
nand U3809 (N_3809,N_3744,N_3739);
nor U3810 (N_3810,N_3741,N_3766);
or U3811 (N_3811,N_3719,N_3708);
or U3812 (N_3812,N_3759,N_3717);
or U3813 (N_3813,N_3769,N_3720);
nor U3814 (N_3814,N_3799,N_3774);
xnor U3815 (N_3815,N_3778,N_3715);
nor U3816 (N_3816,N_3723,N_3737);
and U3817 (N_3817,N_3767,N_3793);
xor U3818 (N_3818,N_3716,N_3761);
or U3819 (N_3819,N_3722,N_3745);
nor U3820 (N_3820,N_3746,N_3772);
nor U3821 (N_3821,N_3750,N_3730);
nor U3822 (N_3822,N_3728,N_3703);
nand U3823 (N_3823,N_3763,N_3754);
nor U3824 (N_3824,N_3794,N_3729);
or U3825 (N_3825,N_3760,N_3762);
nand U3826 (N_3826,N_3701,N_3773);
nor U3827 (N_3827,N_3726,N_3736);
and U3828 (N_3828,N_3702,N_3747);
nor U3829 (N_3829,N_3798,N_3748);
nand U3830 (N_3830,N_3789,N_3724);
or U3831 (N_3831,N_3797,N_3753);
and U3832 (N_3832,N_3713,N_3734);
and U3833 (N_3833,N_3765,N_3796);
nand U3834 (N_3834,N_3784,N_3714);
nor U3835 (N_3835,N_3788,N_3790);
xor U3836 (N_3836,N_3738,N_3752);
xnor U3837 (N_3837,N_3711,N_3742);
or U3838 (N_3838,N_3780,N_3725);
nand U3839 (N_3839,N_3756,N_3787);
and U3840 (N_3840,N_3783,N_3786);
or U3841 (N_3841,N_3710,N_3727);
nor U3842 (N_3842,N_3700,N_3740);
nand U3843 (N_3843,N_3732,N_3764);
xor U3844 (N_3844,N_3743,N_3785);
and U3845 (N_3845,N_3705,N_3733);
nand U3846 (N_3846,N_3791,N_3776);
nand U3847 (N_3847,N_3757,N_3758);
or U3848 (N_3848,N_3770,N_3775);
or U3849 (N_3849,N_3771,N_3792);
and U3850 (N_3850,N_3733,N_3795);
and U3851 (N_3851,N_3766,N_3742);
nor U3852 (N_3852,N_3744,N_3717);
nand U3853 (N_3853,N_3778,N_3720);
xor U3854 (N_3854,N_3740,N_3763);
and U3855 (N_3855,N_3756,N_3765);
xor U3856 (N_3856,N_3782,N_3770);
nand U3857 (N_3857,N_3721,N_3794);
nor U3858 (N_3858,N_3762,N_3722);
nand U3859 (N_3859,N_3785,N_3712);
and U3860 (N_3860,N_3778,N_3757);
nor U3861 (N_3861,N_3755,N_3735);
xor U3862 (N_3862,N_3787,N_3781);
and U3863 (N_3863,N_3724,N_3790);
and U3864 (N_3864,N_3702,N_3729);
or U3865 (N_3865,N_3775,N_3742);
nand U3866 (N_3866,N_3735,N_3713);
nand U3867 (N_3867,N_3732,N_3797);
nor U3868 (N_3868,N_3771,N_3722);
nand U3869 (N_3869,N_3719,N_3764);
nor U3870 (N_3870,N_3705,N_3737);
or U3871 (N_3871,N_3732,N_3792);
nor U3872 (N_3872,N_3712,N_3795);
and U3873 (N_3873,N_3781,N_3716);
and U3874 (N_3874,N_3747,N_3726);
nor U3875 (N_3875,N_3723,N_3755);
nor U3876 (N_3876,N_3796,N_3753);
nor U3877 (N_3877,N_3758,N_3714);
or U3878 (N_3878,N_3701,N_3794);
nor U3879 (N_3879,N_3752,N_3765);
and U3880 (N_3880,N_3797,N_3703);
nor U3881 (N_3881,N_3766,N_3786);
nor U3882 (N_3882,N_3704,N_3776);
nor U3883 (N_3883,N_3769,N_3737);
nand U3884 (N_3884,N_3716,N_3795);
and U3885 (N_3885,N_3717,N_3705);
nor U3886 (N_3886,N_3798,N_3756);
xor U3887 (N_3887,N_3705,N_3758);
and U3888 (N_3888,N_3725,N_3703);
xor U3889 (N_3889,N_3723,N_3766);
and U3890 (N_3890,N_3791,N_3775);
or U3891 (N_3891,N_3782,N_3709);
and U3892 (N_3892,N_3763,N_3703);
xor U3893 (N_3893,N_3734,N_3704);
xnor U3894 (N_3894,N_3785,N_3753);
or U3895 (N_3895,N_3783,N_3774);
nor U3896 (N_3896,N_3777,N_3756);
nor U3897 (N_3897,N_3776,N_3714);
or U3898 (N_3898,N_3798,N_3799);
or U3899 (N_3899,N_3746,N_3775);
nor U3900 (N_3900,N_3812,N_3873);
nand U3901 (N_3901,N_3830,N_3888);
nor U3902 (N_3902,N_3869,N_3859);
or U3903 (N_3903,N_3828,N_3822);
nand U3904 (N_3904,N_3877,N_3887);
and U3905 (N_3905,N_3892,N_3890);
or U3906 (N_3906,N_3858,N_3818);
and U3907 (N_3907,N_3817,N_3852);
nand U3908 (N_3908,N_3850,N_3860);
and U3909 (N_3909,N_3870,N_3847);
or U3910 (N_3910,N_3863,N_3861);
nand U3911 (N_3911,N_3884,N_3879);
or U3912 (N_3912,N_3886,N_3857);
nor U3913 (N_3913,N_3805,N_3853);
and U3914 (N_3914,N_3881,N_3827);
nor U3915 (N_3915,N_3823,N_3851);
and U3916 (N_3916,N_3854,N_3845);
and U3917 (N_3917,N_3813,N_3893);
and U3918 (N_3918,N_3804,N_3815);
nor U3919 (N_3919,N_3814,N_3810);
or U3920 (N_3920,N_3842,N_3824);
or U3921 (N_3921,N_3872,N_3807);
and U3922 (N_3922,N_3816,N_3855);
and U3923 (N_3923,N_3848,N_3802);
and U3924 (N_3924,N_3803,N_3808);
nand U3925 (N_3925,N_3898,N_3801);
xor U3926 (N_3926,N_3897,N_3880);
nor U3927 (N_3927,N_3846,N_3875);
nor U3928 (N_3928,N_3866,N_3891);
nand U3929 (N_3929,N_3821,N_3811);
and U3930 (N_3930,N_3839,N_3868);
nor U3931 (N_3931,N_3800,N_3831);
nand U3932 (N_3932,N_3837,N_3899);
xnor U3933 (N_3933,N_3894,N_3809);
nand U3934 (N_3934,N_3856,N_3862);
or U3935 (N_3935,N_3825,N_3889);
xnor U3936 (N_3936,N_3833,N_3836);
and U3937 (N_3937,N_3871,N_3867);
nand U3938 (N_3938,N_3896,N_3876);
nand U3939 (N_3939,N_3835,N_3841);
nor U3940 (N_3940,N_3819,N_3874);
xnor U3941 (N_3941,N_3838,N_3885);
xor U3942 (N_3942,N_3864,N_3820);
xnor U3943 (N_3943,N_3843,N_3834);
xor U3944 (N_3944,N_3826,N_3840);
and U3945 (N_3945,N_3878,N_3882);
nor U3946 (N_3946,N_3829,N_3883);
and U3947 (N_3947,N_3806,N_3895);
and U3948 (N_3948,N_3865,N_3832);
and U3949 (N_3949,N_3844,N_3849);
nor U3950 (N_3950,N_3882,N_3867);
nand U3951 (N_3951,N_3868,N_3872);
xnor U3952 (N_3952,N_3871,N_3813);
or U3953 (N_3953,N_3881,N_3815);
or U3954 (N_3954,N_3818,N_3882);
nor U3955 (N_3955,N_3813,N_3839);
nand U3956 (N_3956,N_3890,N_3823);
nor U3957 (N_3957,N_3867,N_3883);
and U3958 (N_3958,N_3845,N_3850);
or U3959 (N_3959,N_3888,N_3831);
nand U3960 (N_3960,N_3886,N_3820);
xor U3961 (N_3961,N_3876,N_3837);
nand U3962 (N_3962,N_3838,N_3839);
nand U3963 (N_3963,N_3871,N_3881);
or U3964 (N_3964,N_3804,N_3822);
nor U3965 (N_3965,N_3844,N_3830);
or U3966 (N_3966,N_3842,N_3838);
and U3967 (N_3967,N_3892,N_3853);
nand U3968 (N_3968,N_3803,N_3858);
nor U3969 (N_3969,N_3896,N_3851);
and U3970 (N_3970,N_3809,N_3889);
or U3971 (N_3971,N_3815,N_3842);
and U3972 (N_3972,N_3885,N_3833);
xor U3973 (N_3973,N_3850,N_3814);
and U3974 (N_3974,N_3846,N_3834);
nor U3975 (N_3975,N_3848,N_3843);
or U3976 (N_3976,N_3871,N_3880);
or U3977 (N_3977,N_3896,N_3815);
and U3978 (N_3978,N_3830,N_3828);
nor U3979 (N_3979,N_3818,N_3896);
nor U3980 (N_3980,N_3840,N_3881);
nand U3981 (N_3981,N_3874,N_3848);
and U3982 (N_3982,N_3875,N_3810);
or U3983 (N_3983,N_3896,N_3858);
nand U3984 (N_3984,N_3831,N_3805);
or U3985 (N_3985,N_3839,N_3896);
nor U3986 (N_3986,N_3823,N_3876);
nand U3987 (N_3987,N_3859,N_3857);
and U3988 (N_3988,N_3879,N_3852);
nor U3989 (N_3989,N_3811,N_3886);
or U3990 (N_3990,N_3890,N_3835);
and U3991 (N_3991,N_3829,N_3800);
nand U3992 (N_3992,N_3875,N_3837);
nor U3993 (N_3993,N_3869,N_3867);
or U3994 (N_3994,N_3827,N_3835);
nor U3995 (N_3995,N_3897,N_3833);
nand U3996 (N_3996,N_3837,N_3855);
and U3997 (N_3997,N_3893,N_3823);
and U3998 (N_3998,N_3816,N_3883);
nor U3999 (N_3999,N_3812,N_3809);
xor U4000 (N_4000,N_3901,N_3962);
nand U4001 (N_4001,N_3980,N_3987);
nor U4002 (N_4002,N_3936,N_3904);
nand U4003 (N_4003,N_3967,N_3951);
nand U4004 (N_4004,N_3970,N_3937);
nand U4005 (N_4005,N_3992,N_3926);
and U4006 (N_4006,N_3906,N_3976);
nand U4007 (N_4007,N_3978,N_3958);
or U4008 (N_4008,N_3946,N_3902);
xnor U4009 (N_4009,N_3973,N_3908);
nand U4010 (N_4010,N_3950,N_3903);
nand U4011 (N_4011,N_3944,N_3954);
or U4012 (N_4012,N_3974,N_3933);
xnor U4013 (N_4013,N_3941,N_3984);
or U4014 (N_4014,N_3917,N_3905);
nand U4015 (N_4015,N_3940,N_3989);
or U4016 (N_4016,N_3916,N_3910);
nor U4017 (N_4017,N_3953,N_3909);
nor U4018 (N_4018,N_3945,N_3995);
nor U4019 (N_4019,N_3935,N_3907);
or U4020 (N_4020,N_3900,N_3948);
or U4021 (N_4021,N_3994,N_3920);
xnor U4022 (N_4022,N_3983,N_3959);
xnor U4023 (N_4023,N_3975,N_3972);
or U4024 (N_4024,N_3932,N_3928);
nand U4025 (N_4025,N_3918,N_3938);
nor U4026 (N_4026,N_3911,N_3952);
or U4027 (N_4027,N_3991,N_3914);
xnor U4028 (N_4028,N_3960,N_3913);
nor U4029 (N_4029,N_3955,N_3957);
xor U4030 (N_4030,N_3919,N_3966);
nand U4031 (N_4031,N_3993,N_3981);
and U4032 (N_4032,N_3969,N_3956);
and U4033 (N_4033,N_3971,N_3939);
or U4034 (N_4034,N_3931,N_3929);
nand U4035 (N_4035,N_3988,N_3982);
and U4036 (N_4036,N_3912,N_3943);
and U4037 (N_4037,N_3965,N_3924);
nor U4038 (N_4038,N_3996,N_3977);
and U4039 (N_4039,N_3949,N_3923);
and U4040 (N_4040,N_3985,N_3921);
or U4041 (N_4041,N_3990,N_3979);
and U4042 (N_4042,N_3998,N_3925);
or U4043 (N_4043,N_3927,N_3961);
or U4044 (N_4044,N_3922,N_3963);
or U4045 (N_4045,N_3964,N_3968);
and U4046 (N_4046,N_3986,N_3999);
nor U4047 (N_4047,N_3915,N_3934);
or U4048 (N_4048,N_3947,N_3942);
or U4049 (N_4049,N_3930,N_3997);
nor U4050 (N_4050,N_3930,N_3962);
nor U4051 (N_4051,N_3952,N_3907);
and U4052 (N_4052,N_3987,N_3915);
nor U4053 (N_4053,N_3938,N_3992);
xnor U4054 (N_4054,N_3933,N_3947);
nor U4055 (N_4055,N_3923,N_3958);
nor U4056 (N_4056,N_3984,N_3919);
or U4057 (N_4057,N_3956,N_3943);
xor U4058 (N_4058,N_3940,N_3928);
nor U4059 (N_4059,N_3910,N_3948);
or U4060 (N_4060,N_3932,N_3966);
or U4061 (N_4061,N_3978,N_3987);
and U4062 (N_4062,N_3907,N_3917);
and U4063 (N_4063,N_3971,N_3967);
nand U4064 (N_4064,N_3917,N_3904);
and U4065 (N_4065,N_3982,N_3950);
or U4066 (N_4066,N_3943,N_3964);
or U4067 (N_4067,N_3952,N_3927);
nor U4068 (N_4068,N_3907,N_3950);
nor U4069 (N_4069,N_3917,N_3980);
nor U4070 (N_4070,N_3953,N_3925);
or U4071 (N_4071,N_3945,N_3994);
nor U4072 (N_4072,N_3923,N_3967);
and U4073 (N_4073,N_3956,N_3987);
nor U4074 (N_4074,N_3965,N_3944);
nor U4075 (N_4075,N_3995,N_3907);
xnor U4076 (N_4076,N_3946,N_3983);
or U4077 (N_4077,N_3972,N_3924);
and U4078 (N_4078,N_3931,N_3961);
nand U4079 (N_4079,N_3935,N_3918);
or U4080 (N_4080,N_3949,N_3952);
or U4081 (N_4081,N_3926,N_3911);
or U4082 (N_4082,N_3937,N_3994);
nor U4083 (N_4083,N_3955,N_3987);
and U4084 (N_4084,N_3913,N_3928);
and U4085 (N_4085,N_3964,N_3937);
xor U4086 (N_4086,N_3912,N_3987);
nor U4087 (N_4087,N_3941,N_3971);
or U4088 (N_4088,N_3915,N_3933);
xor U4089 (N_4089,N_3911,N_3982);
xnor U4090 (N_4090,N_3916,N_3911);
and U4091 (N_4091,N_3988,N_3947);
nor U4092 (N_4092,N_3983,N_3928);
nand U4093 (N_4093,N_3955,N_3944);
and U4094 (N_4094,N_3938,N_3900);
and U4095 (N_4095,N_3944,N_3968);
nand U4096 (N_4096,N_3914,N_3973);
nand U4097 (N_4097,N_3988,N_3943);
and U4098 (N_4098,N_3928,N_3993);
nand U4099 (N_4099,N_3922,N_3976);
nor U4100 (N_4100,N_4021,N_4027);
and U4101 (N_4101,N_4071,N_4057);
nand U4102 (N_4102,N_4020,N_4099);
nand U4103 (N_4103,N_4010,N_4034);
or U4104 (N_4104,N_4022,N_4044);
and U4105 (N_4105,N_4047,N_4015);
nor U4106 (N_4106,N_4088,N_4023);
and U4107 (N_4107,N_4030,N_4063);
and U4108 (N_4108,N_4009,N_4006);
xnor U4109 (N_4109,N_4028,N_4074);
xor U4110 (N_4110,N_4042,N_4081);
xnor U4111 (N_4111,N_4094,N_4026);
nor U4112 (N_4112,N_4096,N_4017);
nand U4113 (N_4113,N_4011,N_4084);
or U4114 (N_4114,N_4052,N_4004);
nor U4115 (N_4115,N_4083,N_4065);
xor U4116 (N_4116,N_4005,N_4072);
and U4117 (N_4117,N_4029,N_4060);
nand U4118 (N_4118,N_4070,N_4068);
nor U4119 (N_4119,N_4091,N_4077);
and U4120 (N_4120,N_4043,N_4098);
nor U4121 (N_4121,N_4075,N_4035);
xnor U4122 (N_4122,N_4018,N_4073);
nor U4123 (N_4123,N_4062,N_4036);
nor U4124 (N_4124,N_4003,N_4086);
nand U4125 (N_4125,N_4039,N_4024);
nand U4126 (N_4126,N_4076,N_4085);
and U4127 (N_4127,N_4095,N_4064);
nand U4128 (N_4128,N_4037,N_4014);
or U4129 (N_4129,N_4079,N_4050);
or U4130 (N_4130,N_4048,N_4045);
or U4131 (N_4131,N_4041,N_4016);
nand U4132 (N_4132,N_4056,N_4032);
xor U4133 (N_4133,N_4066,N_4002);
or U4134 (N_4134,N_4001,N_4082);
nor U4135 (N_4135,N_4019,N_4059);
xnor U4136 (N_4136,N_4053,N_4031);
nand U4137 (N_4137,N_4012,N_4061);
nand U4138 (N_4138,N_4080,N_4013);
nand U4139 (N_4139,N_4051,N_4055);
or U4140 (N_4140,N_4033,N_4067);
and U4141 (N_4141,N_4078,N_4038);
and U4142 (N_4142,N_4008,N_4000);
and U4143 (N_4143,N_4049,N_4090);
or U4144 (N_4144,N_4040,N_4097);
and U4145 (N_4145,N_4092,N_4054);
xnor U4146 (N_4146,N_4087,N_4046);
nor U4147 (N_4147,N_4093,N_4025);
nand U4148 (N_4148,N_4089,N_4058);
nand U4149 (N_4149,N_4069,N_4007);
nand U4150 (N_4150,N_4049,N_4046);
nand U4151 (N_4151,N_4094,N_4049);
and U4152 (N_4152,N_4094,N_4079);
and U4153 (N_4153,N_4099,N_4047);
nor U4154 (N_4154,N_4064,N_4049);
nor U4155 (N_4155,N_4084,N_4093);
nor U4156 (N_4156,N_4078,N_4021);
xnor U4157 (N_4157,N_4055,N_4028);
nand U4158 (N_4158,N_4079,N_4081);
or U4159 (N_4159,N_4053,N_4042);
nor U4160 (N_4160,N_4085,N_4003);
nor U4161 (N_4161,N_4049,N_4060);
and U4162 (N_4162,N_4075,N_4039);
nor U4163 (N_4163,N_4057,N_4044);
nand U4164 (N_4164,N_4089,N_4035);
nor U4165 (N_4165,N_4066,N_4080);
xor U4166 (N_4166,N_4007,N_4055);
or U4167 (N_4167,N_4074,N_4018);
nand U4168 (N_4168,N_4057,N_4048);
and U4169 (N_4169,N_4000,N_4071);
or U4170 (N_4170,N_4042,N_4043);
nor U4171 (N_4171,N_4092,N_4000);
nor U4172 (N_4172,N_4098,N_4061);
and U4173 (N_4173,N_4015,N_4067);
nand U4174 (N_4174,N_4088,N_4070);
xor U4175 (N_4175,N_4080,N_4008);
nand U4176 (N_4176,N_4025,N_4070);
xor U4177 (N_4177,N_4036,N_4077);
or U4178 (N_4178,N_4043,N_4032);
xnor U4179 (N_4179,N_4062,N_4012);
nor U4180 (N_4180,N_4047,N_4088);
xor U4181 (N_4181,N_4001,N_4049);
or U4182 (N_4182,N_4092,N_4011);
nor U4183 (N_4183,N_4073,N_4029);
or U4184 (N_4184,N_4098,N_4027);
nor U4185 (N_4185,N_4086,N_4058);
and U4186 (N_4186,N_4004,N_4054);
nand U4187 (N_4187,N_4076,N_4084);
and U4188 (N_4188,N_4014,N_4040);
nor U4189 (N_4189,N_4028,N_4040);
xnor U4190 (N_4190,N_4065,N_4007);
and U4191 (N_4191,N_4072,N_4061);
or U4192 (N_4192,N_4093,N_4051);
and U4193 (N_4193,N_4055,N_4056);
or U4194 (N_4194,N_4058,N_4040);
nand U4195 (N_4195,N_4024,N_4001);
nand U4196 (N_4196,N_4024,N_4099);
and U4197 (N_4197,N_4015,N_4046);
xor U4198 (N_4198,N_4056,N_4054);
nor U4199 (N_4199,N_4017,N_4055);
xor U4200 (N_4200,N_4156,N_4160);
and U4201 (N_4201,N_4139,N_4170);
nand U4202 (N_4202,N_4196,N_4115);
nor U4203 (N_4203,N_4197,N_4185);
and U4204 (N_4204,N_4103,N_4187);
nor U4205 (N_4205,N_4102,N_4136);
or U4206 (N_4206,N_4171,N_4122);
or U4207 (N_4207,N_4107,N_4106);
nor U4208 (N_4208,N_4148,N_4142);
and U4209 (N_4209,N_4191,N_4165);
nor U4210 (N_4210,N_4182,N_4134);
or U4211 (N_4211,N_4155,N_4132);
nand U4212 (N_4212,N_4147,N_4118);
and U4213 (N_4213,N_4138,N_4166);
and U4214 (N_4214,N_4125,N_4195);
nand U4215 (N_4215,N_4188,N_4157);
xor U4216 (N_4216,N_4105,N_4177);
nor U4217 (N_4217,N_4130,N_4110);
nor U4218 (N_4218,N_4183,N_4117);
nand U4219 (N_4219,N_4108,N_4113);
nand U4220 (N_4220,N_4194,N_4146);
or U4221 (N_4221,N_4131,N_4192);
xnor U4222 (N_4222,N_4168,N_4119);
or U4223 (N_4223,N_4184,N_4154);
nand U4224 (N_4224,N_4140,N_4135);
and U4225 (N_4225,N_4120,N_4124);
nor U4226 (N_4226,N_4169,N_4199);
nor U4227 (N_4227,N_4153,N_4144);
or U4228 (N_4228,N_4143,N_4193);
and U4229 (N_4229,N_4133,N_4172);
or U4230 (N_4230,N_4179,N_4116);
nand U4231 (N_4231,N_4127,N_4161);
xnor U4232 (N_4232,N_4181,N_4167);
nor U4233 (N_4233,N_4158,N_4175);
xor U4234 (N_4234,N_4159,N_4163);
xnor U4235 (N_4235,N_4173,N_4104);
nor U4236 (N_4236,N_4186,N_4109);
nor U4237 (N_4237,N_4126,N_4121);
nor U4238 (N_4238,N_4176,N_4150);
or U4239 (N_4239,N_4111,N_4129);
and U4240 (N_4240,N_4178,N_4149);
nor U4241 (N_4241,N_4164,N_4100);
or U4242 (N_4242,N_4151,N_4180);
nor U4243 (N_4243,N_4128,N_4152);
nor U4244 (N_4244,N_4112,N_4174);
or U4245 (N_4245,N_4101,N_4137);
nand U4246 (N_4246,N_4189,N_4162);
and U4247 (N_4247,N_4145,N_4198);
nor U4248 (N_4248,N_4141,N_4190);
and U4249 (N_4249,N_4114,N_4123);
or U4250 (N_4250,N_4156,N_4194);
or U4251 (N_4251,N_4165,N_4128);
nor U4252 (N_4252,N_4109,N_4192);
nor U4253 (N_4253,N_4141,N_4151);
nand U4254 (N_4254,N_4116,N_4130);
nor U4255 (N_4255,N_4148,N_4125);
or U4256 (N_4256,N_4172,N_4152);
nor U4257 (N_4257,N_4176,N_4114);
and U4258 (N_4258,N_4165,N_4148);
nand U4259 (N_4259,N_4131,N_4153);
or U4260 (N_4260,N_4182,N_4143);
nor U4261 (N_4261,N_4112,N_4123);
or U4262 (N_4262,N_4146,N_4142);
nor U4263 (N_4263,N_4142,N_4170);
and U4264 (N_4264,N_4110,N_4194);
nand U4265 (N_4265,N_4182,N_4167);
nand U4266 (N_4266,N_4105,N_4101);
nand U4267 (N_4267,N_4173,N_4157);
nand U4268 (N_4268,N_4177,N_4119);
nor U4269 (N_4269,N_4157,N_4198);
xor U4270 (N_4270,N_4196,N_4190);
or U4271 (N_4271,N_4192,N_4196);
nand U4272 (N_4272,N_4152,N_4189);
or U4273 (N_4273,N_4189,N_4176);
nor U4274 (N_4274,N_4108,N_4162);
xnor U4275 (N_4275,N_4172,N_4145);
or U4276 (N_4276,N_4123,N_4116);
nor U4277 (N_4277,N_4149,N_4152);
and U4278 (N_4278,N_4104,N_4126);
and U4279 (N_4279,N_4172,N_4115);
nor U4280 (N_4280,N_4187,N_4166);
nand U4281 (N_4281,N_4108,N_4149);
nor U4282 (N_4282,N_4188,N_4196);
nand U4283 (N_4283,N_4166,N_4174);
xor U4284 (N_4284,N_4125,N_4132);
and U4285 (N_4285,N_4140,N_4119);
and U4286 (N_4286,N_4109,N_4172);
nand U4287 (N_4287,N_4144,N_4195);
nor U4288 (N_4288,N_4195,N_4132);
nand U4289 (N_4289,N_4163,N_4171);
and U4290 (N_4290,N_4122,N_4121);
and U4291 (N_4291,N_4125,N_4152);
nand U4292 (N_4292,N_4109,N_4164);
or U4293 (N_4293,N_4183,N_4178);
nor U4294 (N_4294,N_4194,N_4131);
nand U4295 (N_4295,N_4177,N_4174);
and U4296 (N_4296,N_4156,N_4104);
nor U4297 (N_4297,N_4175,N_4152);
or U4298 (N_4298,N_4192,N_4189);
nand U4299 (N_4299,N_4119,N_4154);
and U4300 (N_4300,N_4285,N_4202);
nand U4301 (N_4301,N_4264,N_4206);
nor U4302 (N_4302,N_4227,N_4284);
or U4303 (N_4303,N_4204,N_4282);
xnor U4304 (N_4304,N_4236,N_4241);
and U4305 (N_4305,N_4299,N_4271);
nor U4306 (N_4306,N_4278,N_4224);
xor U4307 (N_4307,N_4210,N_4261);
xnor U4308 (N_4308,N_4280,N_4268);
or U4309 (N_4309,N_4291,N_4238);
and U4310 (N_4310,N_4290,N_4255);
nor U4311 (N_4311,N_4251,N_4211);
or U4312 (N_4312,N_4297,N_4266);
nor U4313 (N_4313,N_4257,N_4272);
or U4314 (N_4314,N_4229,N_4298);
nor U4315 (N_4315,N_4208,N_4287);
and U4316 (N_4316,N_4263,N_4267);
or U4317 (N_4317,N_4239,N_4270);
and U4318 (N_4318,N_4218,N_4233);
or U4319 (N_4319,N_4205,N_4212);
nor U4320 (N_4320,N_4223,N_4234);
and U4321 (N_4321,N_4295,N_4242);
or U4322 (N_4322,N_4260,N_4214);
or U4323 (N_4323,N_4245,N_4209);
nand U4324 (N_4324,N_4273,N_4248);
nand U4325 (N_4325,N_4213,N_4262);
nor U4326 (N_4326,N_4293,N_4279);
or U4327 (N_4327,N_4254,N_4276);
nor U4328 (N_4328,N_4249,N_4275);
xor U4329 (N_4329,N_4217,N_4252);
nor U4330 (N_4330,N_4296,N_4243);
and U4331 (N_4331,N_4244,N_4250);
or U4332 (N_4332,N_4231,N_4288);
or U4333 (N_4333,N_4232,N_4274);
and U4334 (N_4334,N_4258,N_4215);
nor U4335 (N_4335,N_4221,N_4226);
xor U4336 (N_4336,N_4265,N_4283);
nor U4337 (N_4337,N_4259,N_4203);
and U4338 (N_4338,N_4200,N_4240);
and U4339 (N_4339,N_4289,N_4201);
xnor U4340 (N_4340,N_4230,N_4235);
nor U4341 (N_4341,N_4228,N_4225);
or U4342 (N_4342,N_4294,N_4237);
and U4343 (N_4343,N_4219,N_4207);
and U4344 (N_4344,N_4246,N_4222);
or U4345 (N_4345,N_4253,N_4247);
nand U4346 (N_4346,N_4281,N_4220);
xor U4347 (N_4347,N_4269,N_4292);
or U4348 (N_4348,N_4286,N_4256);
nor U4349 (N_4349,N_4277,N_4216);
and U4350 (N_4350,N_4281,N_4273);
and U4351 (N_4351,N_4297,N_4268);
and U4352 (N_4352,N_4223,N_4231);
nor U4353 (N_4353,N_4238,N_4260);
and U4354 (N_4354,N_4220,N_4289);
nand U4355 (N_4355,N_4200,N_4249);
or U4356 (N_4356,N_4263,N_4226);
and U4357 (N_4357,N_4250,N_4294);
nor U4358 (N_4358,N_4246,N_4230);
and U4359 (N_4359,N_4235,N_4224);
nand U4360 (N_4360,N_4220,N_4277);
or U4361 (N_4361,N_4265,N_4226);
nor U4362 (N_4362,N_4224,N_4263);
and U4363 (N_4363,N_4294,N_4258);
nor U4364 (N_4364,N_4296,N_4225);
and U4365 (N_4365,N_4254,N_4203);
nor U4366 (N_4366,N_4260,N_4221);
xor U4367 (N_4367,N_4296,N_4259);
xor U4368 (N_4368,N_4237,N_4293);
xnor U4369 (N_4369,N_4250,N_4210);
nand U4370 (N_4370,N_4287,N_4214);
xnor U4371 (N_4371,N_4212,N_4262);
xor U4372 (N_4372,N_4281,N_4233);
and U4373 (N_4373,N_4261,N_4266);
nand U4374 (N_4374,N_4279,N_4261);
nor U4375 (N_4375,N_4255,N_4252);
xor U4376 (N_4376,N_4215,N_4295);
nand U4377 (N_4377,N_4257,N_4230);
nand U4378 (N_4378,N_4233,N_4286);
nor U4379 (N_4379,N_4299,N_4220);
nand U4380 (N_4380,N_4277,N_4280);
and U4381 (N_4381,N_4240,N_4264);
nor U4382 (N_4382,N_4215,N_4223);
and U4383 (N_4383,N_4209,N_4207);
nand U4384 (N_4384,N_4205,N_4202);
or U4385 (N_4385,N_4232,N_4239);
or U4386 (N_4386,N_4272,N_4246);
nor U4387 (N_4387,N_4283,N_4270);
and U4388 (N_4388,N_4279,N_4225);
nor U4389 (N_4389,N_4213,N_4210);
xor U4390 (N_4390,N_4254,N_4225);
nand U4391 (N_4391,N_4273,N_4245);
or U4392 (N_4392,N_4227,N_4294);
nand U4393 (N_4393,N_4291,N_4236);
xnor U4394 (N_4394,N_4235,N_4264);
nand U4395 (N_4395,N_4248,N_4230);
nor U4396 (N_4396,N_4238,N_4249);
and U4397 (N_4397,N_4241,N_4233);
xor U4398 (N_4398,N_4243,N_4245);
or U4399 (N_4399,N_4200,N_4238);
or U4400 (N_4400,N_4398,N_4396);
nand U4401 (N_4401,N_4394,N_4348);
xnor U4402 (N_4402,N_4322,N_4309);
nor U4403 (N_4403,N_4339,N_4382);
or U4404 (N_4404,N_4301,N_4375);
nor U4405 (N_4405,N_4391,N_4393);
nor U4406 (N_4406,N_4366,N_4369);
and U4407 (N_4407,N_4353,N_4359);
nand U4408 (N_4408,N_4390,N_4327);
nor U4409 (N_4409,N_4328,N_4317);
or U4410 (N_4410,N_4316,N_4312);
nand U4411 (N_4411,N_4344,N_4305);
or U4412 (N_4412,N_4323,N_4329);
nor U4413 (N_4413,N_4374,N_4395);
nand U4414 (N_4414,N_4372,N_4343);
nor U4415 (N_4415,N_4357,N_4365);
or U4416 (N_4416,N_4304,N_4387);
nand U4417 (N_4417,N_4378,N_4385);
nor U4418 (N_4418,N_4318,N_4345);
nor U4419 (N_4419,N_4388,N_4303);
and U4420 (N_4420,N_4381,N_4306);
or U4421 (N_4421,N_4370,N_4354);
xnor U4422 (N_4422,N_4389,N_4333);
nor U4423 (N_4423,N_4352,N_4371);
and U4424 (N_4424,N_4325,N_4355);
nor U4425 (N_4425,N_4361,N_4302);
xor U4426 (N_4426,N_4346,N_4349);
xnor U4427 (N_4427,N_4300,N_4386);
nor U4428 (N_4428,N_4350,N_4399);
nor U4429 (N_4429,N_4330,N_4373);
or U4430 (N_4430,N_4332,N_4397);
nor U4431 (N_4431,N_4341,N_4331);
nor U4432 (N_4432,N_4358,N_4336);
nor U4433 (N_4433,N_4368,N_4340);
or U4434 (N_4434,N_4310,N_4311);
or U4435 (N_4435,N_4364,N_4379);
and U4436 (N_4436,N_4380,N_4338);
and U4437 (N_4437,N_4362,N_4314);
nor U4438 (N_4438,N_4356,N_4337);
nor U4439 (N_4439,N_4308,N_4351);
or U4440 (N_4440,N_4384,N_4335);
or U4441 (N_4441,N_4334,N_4367);
or U4442 (N_4442,N_4319,N_4377);
and U4443 (N_4443,N_4347,N_4313);
and U4444 (N_4444,N_4307,N_4315);
nor U4445 (N_4445,N_4342,N_4360);
nand U4446 (N_4446,N_4326,N_4363);
nand U4447 (N_4447,N_4321,N_4383);
or U4448 (N_4448,N_4320,N_4376);
and U4449 (N_4449,N_4392,N_4324);
nor U4450 (N_4450,N_4305,N_4356);
nand U4451 (N_4451,N_4332,N_4387);
or U4452 (N_4452,N_4322,N_4380);
or U4453 (N_4453,N_4387,N_4327);
nand U4454 (N_4454,N_4323,N_4320);
xnor U4455 (N_4455,N_4343,N_4387);
and U4456 (N_4456,N_4340,N_4325);
or U4457 (N_4457,N_4321,N_4382);
and U4458 (N_4458,N_4315,N_4325);
nor U4459 (N_4459,N_4398,N_4389);
nand U4460 (N_4460,N_4342,N_4385);
nand U4461 (N_4461,N_4346,N_4396);
xnor U4462 (N_4462,N_4375,N_4349);
and U4463 (N_4463,N_4310,N_4396);
and U4464 (N_4464,N_4396,N_4353);
or U4465 (N_4465,N_4390,N_4357);
nor U4466 (N_4466,N_4353,N_4395);
or U4467 (N_4467,N_4338,N_4327);
and U4468 (N_4468,N_4341,N_4379);
nor U4469 (N_4469,N_4349,N_4376);
xor U4470 (N_4470,N_4392,N_4339);
and U4471 (N_4471,N_4315,N_4314);
nor U4472 (N_4472,N_4388,N_4301);
nor U4473 (N_4473,N_4317,N_4382);
and U4474 (N_4474,N_4314,N_4317);
and U4475 (N_4475,N_4399,N_4372);
and U4476 (N_4476,N_4329,N_4316);
xor U4477 (N_4477,N_4343,N_4348);
and U4478 (N_4478,N_4378,N_4393);
nand U4479 (N_4479,N_4360,N_4305);
nor U4480 (N_4480,N_4341,N_4326);
nor U4481 (N_4481,N_4314,N_4306);
nand U4482 (N_4482,N_4372,N_4376);
or U4483 (N_4483,N_4334,N_4310);
nand U4484 (N_4484,N_4315,N_4305);
or U4485 (N_4485,N_4355,N_4310);
and U4486 (N_4486,N_4391,N_4382);
and U4487 (N_4487,N_4313,N_4314);
and U4488 (N_4488,N_4311,N_4350);
xor U4489 (N_4489,N_4300,N_4374);
and U4490 (N_4490,N_4389,N_4379);
nand U4491 (N_4491,N_4369,N_4319);
nor U4492 (N_4492,N_4366,N_4374);
nor U4493 (N_4493,N_4385,N_4321);
and U4494 (N_4494,N_4317,N_4303);
nor U4495 (N_4495,N_4398,N_4334);
and U4496 (N_4496,N_4325,N_4345);
xnor U4497 (N_4497,N_4338,N_4387);
and U4498 (N_4498,N_4323,N_4307);
and U4499 (N_4499,N_4344,N_4333);
and U4500 (N_4500,N_4494,N_4477);
nor U4501 (N_4501,N_4462,N_4434);
nand U4502 (N_4502,N_4418,N_4459);
nand U4503 (N_4503,N_4411,N_4452);
nor U4504 (N_4504,N_4488,N_4416);
nand U4505 (N_4505,N_4438,N_4430);
xnor U4506 (N_4506,N_4410,N_4433);
or U4507 (N_4507,N_4482,N_4417);
and U4508 (N_4508,N_4439,N_4454);
and U4509 (N_4509,N_4443,N_4475);
or U4510 (N_4510,N_4442,N_4421);
xnor U4511 (N_4511,N_4474,N_4468);
nand U4512 (N_4512,N_4425,N_4455);
xor U4513 (N_4513,N_4435,N_4490);
or U4514 (N_4514,N_4437,N_4448);
nor U4515 (N_4515,N_4473,N_4465);
nand U4516 (N_4516,N_4424,N_4481);
nor U4517 (N_4517,N_4491,N_4420);
and U4518 (N_4518,N_4471,N_4485);
or U4519 (N_4519,N_4414,N_4478);
nor U4520 (N_4520,N_4401,N_4466);
nor U4521 (N_4521,N_4453,N_4460);
or U4522 (N_4522,N_4498,N_4487);
nor U4523 (N_4523,N_4402,N_4444);
nand U4524 (N_4524,N_4457,N_4461);
and U4525 (N_4525,N_4451,N_4486);
nand U4526 (N_4526,N_4495,N_4483);
and U4527 (N_4527,N_4415,N_4492);
nor U4528 (N_4528,N_4404,N_4464);
or U4529 (N_4529,N_4458,N_4479);
nand U4530 (N_4530,N_4413,N_4445);
and U4531 (N_4531,N_4441,N_4456);
nand U4532 (N_4532,N_4428,N_4450);
or U4533 (N_4533,N_4440,N_4470);
nand U4534 (N_4534,N_4407,N_4449);
nand U4535 (N_4535,N_4403,N_4408);
or U4536 (N_4536,N_4427,N_4469);
nor U4537 (N_4537,N_4405,N_4422);
nand U4538 (N_4538,N_4447,N_4446);
and U4539 (N_4539,N_4476,N_4489);
or U4540 (N_4540,N_4436,N_4423);
or U4541 (N_4541,N_4467,N_4409);
and U4542 (N_4542,N_4431,N_4472);
nand U4543 (N_4543,N_4480,N_4426);
nor U4544 (N_4544,N_4493,N_4499);
or U4545 (N_4545,N_4419,N_4432);
or U4546 (N_4546,N_4429,N_4496);
and U4547 (N_4547,N_4400,N_4412);
xnor U4548 (N_4548,N_4497,N_4463);
or U4549 (N_4549,N_4484,N_4406);
or U4550 (N_4550,N_4455,N_4457);
xnor U4551 (N_4551,N_4435,N_4470);
or U4552 (N_4552,N_4470,N_4452);
nor U4553 (N_4553,N_4412,N_4473);
nand U4554 (N_4554,N_4463,N_4487);
and U4555 (N_4555,N_4413,N_4489);
or U4556 (N_4556,N_4468,N_4476);
nand U4557 (N_4557,N_4400,N_4417);
and U4558 (N_4558,N_4433,N_4485);
nor U4559 (N_4559,N_4431,N_4461);
nor U4560 (N_4560,N_4459,N_4499);
nand U4561 (N_4561,N_4411,N_4450);
nand U4562 (N_4562,N_4448,N_4404);
or U4563 (N_4563,N_4467,N_4454);
or U4564 (N_4564,N_4415,N_4489);
or U4565 (N_4565,N_4419,N_4449);
nand U4566 (N_4566,N_4493,N_4490);
nor U4567 (N_4567,N_4435,N_4482);
xor U4568 (N_4568,N_4483,N_4427);
and U4569 (N_4569,N_4461,N_4443);
nor U4570 (N_4570,N_4494,N_4460);
nor U4571 (N_4571,N_4461,N_4426);
nand U4572 (N_4572,N_4411,N_4481);
nand U4573 (N_4573,N_4498,N_4418);
xnor U4574 (N_4574,N_4438,N_4486);
and U4575 (N_4575,N_4429,N_4405);
nand U4576 (N_4576,N_4468,N_4469);
nand U4577 (N_4577,N_4420,N_4417);
and U4578 (N_4578,N_4406,N_4414);
nand U4579 (N_4579,N_4414,N_4485);
and U4580 (N_4580,N_4440,N_4402);
or U4581 (N_4581,N_4451,N_4491);
and U4582 (N_4582,N_4435,N_4478);
and U4583 (N_4583,N_4423,N_4474);
nand U4584 (N_4584,N_4436,N_4434);
or U4585 (N_4585,N_4463,N_4469);
and U4586 (N_4586,N_4432,N_4425);
or U4587 (N_4587,N_4413,N_4494);
nand U4588 (N_4588,N_4482,N_4401);
xnor U4589 (N_4589,N_4422,N_4469);
nand U4590 (N_4590,N_4459,N_4482);
or U4591 (N_4591,N_4428,N_4471);
or U4592 (N_4592,N_4484,N_4481);
nor U4593 (N_4593,N_4495,N_4401);
nor U4594 (N_4594,N_4480,N_4461);
or U4595 (N_4595,N_4433,N_4454);
nor U4596 (N_4596,N_4475,N_4477);
and U4597 (N_4597,N_4452,N_4401);
or U4598 (N_4598,N_4498,N_4461);
xnor U4599 (N_4599,N_4428,N_4494);
nor U4600 (N_4600,N_4559,N_4547);
and U4601 (N_4601,N_4555,N_4538);
nor U4602 (N_4602,N_4507,N_4508);
and U4603 (N_4603,N_4585,N_4568);
and U4604 (N_4604,N_4552,N_4500);
nand U4605 (N_4605,N_4548,N_4516);
nand U4606 (N_4606,N_4567,N_4519);
and U4607 (N_4607,N_4566,N_4578);
nand U4608 (N_4608,N_4520,N_4532);
nand U4609 (N_4609,N_4599,N_4565);
nor U4610 (N_4610,N_4534,N_4583);
nor U4611 (N_4611,N_4587,N_4522);
or U4612 (N_4612,N_4561,N_4521);
or U4613 (N_4613,N_4506,N_4582);
and U4614 (N_4614,N_4560,N_4594);
and U4615 (N_4615,N_4571,N_4576);
xor U4616 (N_4616,N_4581,N_4509);
nand U4617 (N_4617,N_4524,N_4535);
nor U4618 (N_4618,N_4528,N_4510);
and U4619 (N_4619,N_4588,N_4536);
nand U4620 (N_4620,N_4531,N_4580);
and U4621 (N_4621,N_4541,N_4586);
nor U4622 (N_4622,N_4550,N_4544);
or U4623 (N_4623,N_4572,N_4579);
or U4624 (N_4624,N_4517,N_4590);
or U4625 (N_4625,N_4533,N_4529);
nand U4626 (N_4626,N_4598,N_4526);
or U4627 (N_4627,N_4527,N_4545);
or U4628 (N_4628,N_4551,N_4557);
and U4629 (N_4629,N_4556,N_4575);
and U4630 (N_4630,N_4596,N_4592);
nand U4631 (N_4631,N_4597,N_4584);
or U4632 (N_4632,N_4505,N_4542);
or U4633 (N_4633,N_4569,N_4501);
or U4634 (N_4634,N_4591,N_4562);
nor U4635 (N_4635,N_4502,N_4546);
and U4636 (N_4636,N_4577,N_4523);
xor U4637 (N_4637,N_4539,N_4513);
nand U4638 (N_4638,N_4518,N_4589);
nor U4639 (N_4639,N_4514,N_4540);
xor U4640 (N_4640,N_4595,N_4553);
or U4641 (N_4641,N_4511,N_4563);
xor U4642 (N_4642,N_4573,N_4549);
or U4643 (N_4643,N_4512,N_4593);
and U4644 (N_4644,N_4515,N_4504);
and U4645 (N_4645,N_4537,N_4564);
and U4646 (N_4646,N_4554,N_4558);
nor U4647 (N_4647,N_4503,N_4530);
or U4648 (N_4648,N_4570,N_4525);
nor U4649 (N_4649,N_4574,N_4543);
or U4650 (N_4650,N_4569,N_4593);
nor U4651 (N_4651,N_4566,N_4598);
nand U4652 (N_4652,N_4522,N_4527);
nand U4653 (N_4653,N_4526,N_4564);
xor U4654 (N_4654,N_4533,N_4549);
and U4655 (N_4655,N_4576,N_4580);
nand U4656 (N_4656,N_4500,N_4558);
nor U4657 (N_4657,N_4574,N_4528);
nand U4658 (N_4658,N_4520,N_4547);
or U4659 (N_4659,N_4572,N_4588);
nor U4660 (N_4660,N_4550,N_4543);
xor U4661 (N_4661,N_4539,N_4585);
nor U4662 (N_4662,N_4574,N_4570);
nand U4663 (N_4663,N_4502,N_4501);
nor U4664 (N_4664,N_4568,N_4560);
or U4665 (N_4665,N_4534,N_4543);
nor U4666 (N_4666,N_4532,N_4513);
nand U4667 (N_4667,N_4535,N_4576);
nand U4668 (N_4668,N_4514,N_4552);
or U4669 (N_4669,N_4554,N_4548);
nand U4670 (N_4670,N_4571,N_4552);
and U4671 (N_4671,N_4523,N_4571);
and U4672 (N_4672,N_4595,N_4531);
xor U4673 (N_4673,N_4502,N_4532);
nand U4674 (N_4674,N_4573,N_4560);
and U4675 (N_4675,N_4519,N_4521);
or U4676 (N_4676,N_4597,N_4535);
or U4677 (N_4677,N_4523,N_4593);
nor U4678 (N_4678,N_4543,N_4506);
or U4679 (N_4679,N_4562,N_4516);
nand U4680 (N_4680,N_4577,N_4576);
or U4681 (N_4681,N_4575,N_4511);
and U4682 (N_4682,N_4549,N_4506);
nor U4683 (N_4683,N_4597,N_4538);
nor U4684 (N_4684,N_4571,N_4592);
xor U4685 (N_4685,N_4514,N_4535);
or U4686 (N_4686,N_4574,N_4537);
or U4687 (N_4687,N_4542,N_4534);
or U4688 (N_4688,N_4512,N_4565);
nor U4689 (N_4689,N_4581,N_4551);
or U4690 (N_4690,N_4504,N_4522);
nor U4691 (N_4691,N_4508,N_4588);
nor U4692 (N_4692,N_4578,N_4596);
and U4693 (N_4693,N_4557,N_4519);
nand U4694 (N_4694,N_4512,N_4544);
or U4695 (N_4695,N_4583,N_4573);
and U4696 (N_4696,N_4571,N_4511);
and U4697 (N_4697,N_4537,N_4569);
nor U4698 (N_4698,N_4557,N_4544);
nand U4699 (N_4699,N_4527,N_4518);
or U4700 (N_4700,N_4657,N_4604);
and U4701 (N_4701,N_4667,N_4648);
or U4702 (N_4702,N_4668,N_4679);
nand U4703 (N_4703,N_4611,N_4613);
xnor U4704 (N_4704,N_4670,N_4690);
or U4705 (N_4705,N_4699,N_4685);
nor U4706 (N_4706,N_4622,N_4632);
nand U4707 (N_4707,N_4612,N_4655);
nand U4708 (N_4708,N_4600,N_4620);
xnor U4709 (N_4709,N_4636,N_4650);
or U4710 (N_4710,N_4676,N_4605);
nand U4711 (N_4711,N_4601,N_4630);
or U4712 (N_4712,N_4602,N_4689);
and U4713 (N_4713,N_4642,N_4618);
or U4714 (N_4714,N_4686,N_4691);
and U4715 (N_4715,N_4663,N_4695);
nor U4716 (N_4716,N_4631,N_4608);
and U4717 (N_4717,N_4654,N_4672);
and U4718 (N_4718,N_4675,N_4687);
and U4719 (N_4719,N_4678,N_4606);
or U4720 (N_4720,N_4662,N_4637);
or U4721 (N_4721,N_4614,N_4640);
nand U4722 (N_4722,N_4683,N_4625);
nor U4723 (N_4723,N_4665,N_4666);
nor U4724 (N_4724,N_4693,N_4633);
or U4725 (N_4725,N_4610,N_4643);
and U4726 (N_4726,N_4692,N_4653);
nand U4727 (N_4727,N_4615,N_4639);
nand U4728 (N_4728,N_4624,N_4697);
xor U4729 (N_4729,N_4644,N_4629);
nand U4730 (N_4730,N_4628,N_4673);
nand U4731 (N_4731,N_4609,N_4641);
nor U4732 (N_4732,N_4696,N_4669);
and U4733 (N_4733,N_4638,N_4698);
and U4734 (N_4734,N_4658,N_4661);
nor U4735 (N_4735,N_4647,N_4616);
nand U4736 (N_4736,N_4680,N_4634);
and U4737 (N_4737,N_4671,N_4677);
or U4738 (N_4738,N_4681,N_4664);
or U4739 (N_4739,N_4603,N_4682);
nand U4740 (N_4740,N_4656,N_4627);
nor U4741 (N_4741,N_4659,N_4688);
or U4742 (N_4742,N_4635,N_4607);
or U4743 (N_4743,N_4617,N_4646);
xnor U4744 (N_4744,N_4621,N_4651);
nand U4745 (N_4745,N_4649,N_4684);
nand U4746 (N_4746,N_4660,N_4619);
and U4747 (N_4747,N_4674,N_4623);
xor U4748 (N_4748,N_4652,N_4645);
nand U4749 (N_4749,N_4626,N_4694);
or U4750 (N_4750,N_4636,N_4697);
nor U4751 (N_4751,N_4664,N_4603);
xor U4752 (N_4752,N_4615,N_4627);
nor U4753 (N_4753,N_4625,N_4629);
and U4754 (N_4754,N_4660,N_4638);
or U4755 (N_4755,N_4650,N_4684);
nand U4756 (N_4756,N_4653,N_4681);
nor U4757 (N_4757,N_4627,N_4687);
and U4758 (N_4758,N_4669,N_4671);
and U4759 (N_4759,N_4684,N_4676);
nor U4760 (N_4760,N_4645,N_4685);
nand U4761 (N_4761,N_4695,N_4623);
or U4762 (N_4762,N_4675,N_4638);
or U4763 (N_4763,N_4641,N_4637);
or U4764 (N_4764,N_4624,N_4661);
nand U4765 (N_4765,N_4630,N_4648);
and U4766 (N_4766,N_4614,N_4672);
nor U4767 (N_4767,N_4671,N_4696);
nand U4768 (N_4768,N_4697,N_4638);
and U4769 (N_4769,N_4677,N_4652);
nor U4770 (N_4770,N_4698,N_4620);
nand U4771 (N_4771,N_4670,N_4647);
and U4772 (N_4772,N_4662,N_4683);
nor U4773 (N_4773,N_4622,N_4696);
xnor U4774 (N_4774,N_4641,N_4608);
and U4775 (N_4775,N_4646,N_4682);
and U4776 (N_4776,N_4696,N_4648);
nor U4777 (N_4777,N_4697,N_4639);
nor U4778 (N_4778,N_4694,N_4600);
or U4779 (N_4779,N_4688,N_4682);
and U4780 (N_4780,N_4606,N_4626);
nand U4781 (N_4781,N_4674,N_4655);
and U4782 (N_4782,N_4646,N_4637);
nor U4783 (N_4783,N_4686,N_4600);
nand U4784 (N_4784,N_4689,N_4626);
nor U4785 (N_4785,N_4646,N_4676);
nor U4786 (N_4786,N_4678,N_4636);
and U4787 (N_4787,N_4677,N_4628);
nor U4788 (N_4788,N_4635,N_4624);
or U4789 (N_4789,N_4641,N_4678);
or U4790 (N_4790,N_4646,N_4669);
or U4791 (N_4791,N_4672,N_4638);
nand U4792 (N_4792,N_4633,N_4687);
nor U4793 (N_4793,N_4618,N_4611);
nor U4794 (N_4794,N_4656,N_4686);
or U4795 (N_4795,N_4665,N_4657);
and U4796 (N_4796,N_4669,N_4637);
nand U4797 (N_4797,N_4681,N_4645);
and U4798 (N_4798,N_4662,N_4640);
and U4799 (N_4799,N_4631,N_4634);
or U4800 (N_4800,N_4741,N_4715);
and U4801 (N_4801,N_4735,N_4792);
or U4802 (N_4802,N_4733,N_4752);
nand U4803 (N_4803,N_4760,N_4744);
nor U4804 (N_4804,N_4725,N_4761);
nor U4805 (N_4805,N_4762,N_4782);
and U4806 (N_4806,N_4780,N_4729);
nand U4807 (N_4807,N_4703,N_4784);
and U4808 (N_4808,N_4702,N_4786);
nand U4809 (N_4809,N_4788,N_4739);
nand U4810 (N_4810,N_4730,N_4740);
nor U4811 (N_4811,N_4724,N_4790);
nand U4812 (N_4812,N_4700,N_4764);
nand U4813 (N_4813,N_4771,N_4781);
or U4814 (N_4814,N_4705,N_4765);
nand U4815 (N_4815,N_4794,N_4768);
or U4816 (N_4816,N_4791,N_4754);
nor U4817 (N_4817,N_4701,N_4745);
and U4818 (N_4818,N_4717,N_4720);
or U4819 (N_4819,N_4787,N_4713);
nand U4820 (N_4820,N_4726,N_4757);
xnor U4821 (N_4821,N_4759,N_4769);
nor U4822 (N_4822,N_4770,N_4779);
and U4823 (N_4823,N_4756,N_4710);
nand U4824 (N_4824,N_4793,N_4711);
nor U4825 (N_4825,N_4751,N_4743);
xnor U4826 (N_4826,N_4712,N_4748);
nor U4827 (N_4827,N_4773,N_4758);
xor U4828 (N_4828,N_4723,N_4749);
and U4829 (N_4829,N_4777,N_4734);
and U4830 (N_4830,N_4783,N_4798);
or U4831 (N_4831,N_4742,N_4796);
nor U4832 (N_4832,N_4706,N_4774);
and U4833 (N_4833,N_4797,N_4767);
nor U4834 (N_4834,N_4738,N_4776);
xor U4835 (N_4835,N_4766,N_4716);
or U4836 (N_4836,N_4753,N_4727);
nor U4837 (N_4837,N_4731,N_4737);
nor U4838 (N_4838,N_4750,N_4704);
or U4839 (N_4839,N_4707,N_4709);
nor U4840 (N_4840,N_4719,N_4732);
and U4841 (N_4841,N_4799,N_4772);
nand U4842 (N_4842,N_4736,N_4789);
and U4843 (N_4843,N_4721,N_4785);
or U4844 (N_4844,N_4775,N_4746);
nand U4845 (N_4845,N_4755,N_4747);
and U4846 (N_4846,N_4795,N_4778);
nand U4847 (N_4847,N_4718,N_4708);
nor U4848 (N_4848,N_4714,N_4763);
nand U4849 (N_4849,N_4722,N_4728);
nor U4850 (N_4850,N_4737,N_4720);
nand U4851 (N_4851,N_4747,N_4778);
nand U4852 (N_4852,N_4766,N_4720);
nand U4853 (N_4853,N_4738,N_4744);
or U4854 (N_4854,N_4770,N_4734);
nor U4855 (N_4855,N_4707,N_4769);
and U4856 (N_4856,N_4701,N_4793);
nor U4857 (N_4857,N_4720,N_4745);
and U4858 (N_4858,N_4796,N_4719);
nor U4859 (N_4859,N_4713,N_4793);
nor U4860 (N_4860,N_4771,N_4707);
or U4861 (N_4861,N_4786,N_4726);
and U4862 (N_4862,N_4769,N_4755);
and U4863 (N_4863,N_4794,N_4756);
nand U4864 (N_4864,N_4761,N_4722);
or U4865 (N_4865,N_4795,N_4712);
nand U4866 (N_4866,N_4766,N_4752);
or U4867 (N_4867,N_4704,N_4765);
nor U4868 (N_4868,N_4714,N_4799);
or U4869 (N_4869,N_4760,N_4723);
nor U4870 (N_4870,N_4722,N_4748);
and U4871 (N_4871,N_4752,N_4710);
nor U4872 (N_4872,N_4716,N_4761);
nand U4873 (N_4873,N_4740,N_4703);
nor U4874 (N_4874,N_4741,N_4722);
xor U4875 (N_4875,N_4782,N_4771);
xnor U4876 (N_4876,N_4789,N_4725);
nand U4877 (N_4877,N_4745,N_4791);
xnor U4878 (N_4878,N_4710,N_4725);
and U4879 (N_4879,N_4736,N_4735);
xor U4880 (N_4880,N_4796,N_4754);
nor U4881 (N_4881,N_4714,N_4761);
xnor U4882 (N_4882,N_4748,N_4761);
nand U4883 (N_4883,N_4730,N_4746);
nand U4884 (N_4884,N_4710,N_4718);
nor U4885 (N_4885,N_4768,N_4745);
nor U4886 (N_4886,N_4702,N_4752);
nor U4887 (N_4887,N_4768,N_4723);
or U4888 (N_4888,N_4717,N_4703);
and U4889 (N_4889,N_4779,N_4716);
nand U4890 (N_4890,N_4783,N_4785);
nor U4891 (N_4891,N_4778,N_4716);
nand U4892 (N_4892,N_4763,N_4743);
xnor U4893 (N_4893,N_4768,N_4785);
nand U4894 (N_4894,N_4777,N_4745);
and U4895 (N_4895,N_4767,N_4745);
or U4896 (N_4896,N_4721,N_4782);
nand U4897 (N_4897,N_4749,N_4745);
or U4898 (N_4898,N_4755,N_4706);
nand U4899 (N_4899,N_4779,N_4784);
and U4900 (N_4900,N_4831,N_4898);
or U4901 (N_4901,N_4839,N_4848);
or U4902 (N_4902,N_4852,N_4818);
and U4903 (N_4903,N_4820,N_4816);
nand U4904 (N_4904,N_4802,N_4876);
or U4905 (N_4905,N_4886,N_4811);
nand U4906 (N_4906,N_4897,N_4833);
nand U4907 (N_4907,N_4869,N_4849);
and U4908 (N_4908,N_4861,N_4803);
nor U4909 (N_4909,N_4858,N_4815);
and U4910 (N_4910,N_4856,N_4819);
nor U4911 (N_4911,N_4836,N_4873);
and U4912 (N_4912,N_4881,N_4883);
xnor U4913 (N_4913,N_4850,N_4842);
and U4914 (N_4914,N_4859,N_4853);
and U4915 (N_4915,N_4810,N_4829);
or U4916 (N_4916,N_4809,N_4824);
nor U4917 (N_4917,N_4892,N_4828);
and U4918 (N_4918,N_4800,N_4834);
nand U4919 (N_4919,N_4843,N_4855);
nand U4920 (N_4920,N_4879,N_4806);
nor U4921 (N_4921,N_4804,N_4895);
nand U4922 (N_4922,N_4805,N_4817);
nor U4923 (N_4923,N_4899,N_4888);
nor U4924 (N_4924,N_4837,N_4877);
and U4925 (N_4925,N_4891,N_4846);
xor U4926 (N_4926,N_4889,N_4854);
and U4927 (N_4927,N_4887,N_4808);
nor U4928 (N_4928,N_4801,N_4845);
nor U4929 (N_4929,N_4812,N_4860);
or U4930 (N_4930,N_4825,N_4872);
or U4931 (N_4931,N_4896,N_4862);
nand U4932 (N_4932,N_4885,N_4857);
and U4933 (N_4933,N_4875,N_4813);
nand U4934 (N_4934,N_4807,N_4838);
nor U4935 (N_4935,N_4874,N_4864);
and U4936 (N_4936,N_4844,N_4826);
nor U4937 (N_4937,N_4893,N_4865);
xnor U4938 (N_4938,N_4866,N_4814);
nand U4939 (N_4939,N_4867,N_4890);
and U4940 (N_4940,N_4822,N_4884);
nand U4941 (N_4941,N_4882,N_4821);
nand U4942 (N_4942,N_4863,N_4841);
xnor U4943 (N_4943,N_4827,N_4870);
nand U4944 (N_4944,N_4830,N_4840);
nor U4945 (N_4945,N_4868,N_4880);
nor U4946 (N_4946,N_4835,N_4871);
nor U4947 (N_4947,N_4847,N_4894);
or U4948 (N_4948,N_4878,N_4851);
and U4949 (N_4949,N_4823,N_4832);
nand U4950 (N_4950,N_4848,N_4867);
nor U4951 (N_4951,N_4869,N_4802);
nand U4952 (N_4952,N_4808,N_4871);
nor U4953 (N_4953,N_4877,N_4892);
nor U4954 (N_4954,N_4803,N_4855);
nor U4955 (N_4955,N_4810,N_4868);
or U4956 (N_4956,N_4891,N_4865);
or U4957 (N_4957,N_4880,N_4889);
or U4958 (N_4958,N_4869,N_4859);
and U4959 (N_4959,N_4873,N_4853);
and U4960 (N_4960,N_4880,N_4821);
nor U4961 (N_4961,N_4852,N_4843);
nor U4962 (N_4962,N_4824,N_4892);
or U4963 (N_4963,N_4800,N_4837);
nand U4964 (N_4964,N_4898,N_4807);
and U4965 (N_4965,N_4880,N_4827);
nand U4966 (N_4966,N_4816,N_4897);
nor U4967 (N_4967,N_4870,N_4826);
nor U4968 (N_4968,N_4883,N_4841);
nand U4969 (N_4969,N_4881,N_4817);
and U4970 (N_4970,N_4808,N_4846);
nor U4971 (N_4971,N_4809,N_4833);
or U4972 (N_4972,N_4871,N_4832);
and U4973 (N_4973,N_4813,N_4888);
nor U4974 (N_4974,N_4808,N_4888);
xnor U4975 (N_4975,N_4821,N_4897);
and U4976 (N_4976,N_4888,N_4841);
nor U4977 (N_4977,N_4807,N_4805);
and U4978 (N_4978,N_4811,N_4819);
nor U4979 (N_4979,N_4823,N_4837);
or U4980 (N_4980,N_4870,N_4896);
nor U4981 (N_4981,N_4867,N_4868);
or U4982 (N_4982,N_4888,N_4802);
xor U4983 (N_4983,N_4851,N_4881);
xnor U4984 (N_4984,N_4877,N_4800);
or U4985 (N_4985,N_4873,N_4858);
or U4986 (N_4986,N_4857,N_4868);
and U4987 (N_4987,N_4853,N_4845);
or U4988 (N_4988,N_4883,N_4859);
and U4989 (N_4989,N_4851,N_4827);
or U4990 (N_4990,N_4862,N_4884);
nand U4991 (N_4991,N_4899,N_4828);
or U4992 (N_4992,N_4838,N_4894);
nand U4993 (N_4993,N_4830,N_4804);
and U4994 (N_4994,N_4861,N_4807);
xor U4995 (N_4995,N_4829,N_4893);
or U4996 (N_4996,N_4809,N_4897);
nor U4997 (N_4997,N_4854,N_4853);
nor U4998 (N_4998,N_4862,N_4887);
or U4999 (N_4999,N_4871,N_4863);
nor UO_0 (O_0,N_4989,N_4965);
and UO_1 (O_1,N_4912,N_4971);
and UO_2 (O_2,N_4930,N_4937);
nand UO_3 (O_3,N_4947,N_4903);
and UO_4 (O_4,N_4948,N_4934);
xnor UO_5 (O_5,N_4975,N_4921);
nand UO_6 (O_6,N_4914,N_4924);
or UO_7 (O_7,N_4900,N_4920);
nand UO_8 (O_8,N_4972,N_4940);
nand UO_9 (O_9,N_4908,N_4968);
nand UO_10 (O_10,N_4977,N_4929);
and UO_11 (O_11,N_4902,N_4976);
or UO_12 (O_12,N_4973,N_4993);
and UO_13 (O_13,N_4907,N_4981);
xor UO_14 (O_14,N_4922,N_4955);
xnor UO_15 (O_15,N_4941,N_4994);
xor UO_16 (O_16,N_4913,N_4978);
and UO_17 (O_17,N_4919,N_4961);
nor UO_18 (O_18,N_4910,N_4969);
nand UO_19 (O_19,N_4998,N_4970);
nor UO_20 (O_20,N_4925,N_4936);
xor UO_21 (O_21,N_4957,N_4928);
and UO_22 (O_22,N_4999,N_4963);
and UO_23 (O_23,N_4954,N_4938);
or UO_24 (O_24,N_4905,N_4933);
and UO_25 (O_25,N_4990,N_4992);
and UO_26 (O_26,N_4939,N_4951);
nand UO_27 (O_27,N_4935,N_4943);
or UO_28 (O_28,N_4956,N_4915);
xor UO_29 (O_29,N_4980,N_4958);
or UO_30 (O_30,N_4906,N_4982);
and UO_31 (O_31,N_4987,N_4944);
and UO_32 (O_32,N_4986,N_4931);
nand UO_33 (O_33,N_4985,N_4946);
and UO_34 (O_34,N_4974,N_4911);
and UO_35 (O_35,N_4952,N_4953);
xor UO_36 (O_36,N_4901,N_4979);
nor UO_37 (O_37,N_4927,N_4909);
nor UO_38 (O_38,N_4988,N_4996);
xor UO_39 (O_39,N_4904,N_4942);
or UO_40 (O_40,N_4964,N_4984);
nor UO_41 (O_41,N_4945,N_4991);
and UO_42 (O_42,N_4916,N_4949);
or UO_43 (O_43,N_4967,N_4997);
nor UO_44 (O_44,N_4926,N_4923);
xnor UO_45 (O_45,N_4932,N_4966);
nor UO_46 (O_46,N_4950,N_4960);
nand UO_47 (O_47,N_4995,N_4959);
xor UO_48 (O_48,N_4962,N_4918);
nand UO_49 (O_49,N_4917,N_4983);
or UO_50 (O_50,N_4926,N_4989);
nand UO_51 (O_51,N_4901,N_4937);
nand UO_52 (O_52,N_4988,N_4900);
and UO_53 (O_53,N_4937,N_4932);
nor UO_54 (O_54,N_4917,N_4971);
and UO_55 (O_55,N_4978,N_4967);
and UO_56 (O_56,N_4929,N_4917);
nand UO_57 (O_57,N_4967,N_4983);
nand UO_58 (O_58,N_4959,N_4902);
xnor UO_59 (O_59,N_4950,N_4924);
or UO_60 (O_60,N_4969,N_4968);
nand UO_61 (O_61,N_4902,N_4930);
and UO_62 (O_62,N_4994,N_4927);
or UO_63 (O_63,N_4976,N_4961);
nand UO_64 (O_64,N_4944,N_4905);
nor UO_65 (O_65,N_4913,N_4971);
and UO_66 (O_66,N_4937,N_4972);
and UO_67 (O_67,N_4977,N_4990);
nor UO_68 (O_68,N_4908,N_4981);
and UO_69 (O_69,N_4988,N_4972);
xnor UO_70 (O_70,N_4904,N_4945);
nor UO_71 (O_71,N_4963,N_4931);
nand UO_72 (O_72,N_4993,N_4903);
nor UO_73 (O_73,N_4967,N_4912);
or UO_74 (O_74,N_4946,N_4958);
nor UO_75 (O_75,N_4956,N_4977);
nor UO_76 (O_76,N_4962,N_4909);
nor UO_77 (O_77,N_4995,N_4964);
or UO_78 (O_78,N_4944,N_4914);
nor UO_79 (O_79,N_4970,N_4984);
nor UO_80 (O_80,N_4953,N_4966);
xnor UO_81 (O_81,N_4931,N_4951);
and UO_82 (O_82,N_4995,N_4976);
nor UO_83 (O_83,N_4982,N_4908);
nor UO_84 (O_84,N_4930,N_4952);
or UO_85 (O_85,N_4966,N_4964);
nand UO_86 (O_86,N_4909,N_4951);
nor UO_87 (O_87,N_4925,N_4993);
or UO_88 (O_88,N_4946,N_4966);
and UO_89 (O_89,N_4981,N_4972);
nor UO_90 (O_90,N_4919,N_4993);
nor UO_91 (O_91,N_4970,N_4977);
and UO_92 (O_92,N_4963,N_4958);
nor UO_93 (O_93,N_4943,N_4957);
and UO_94 (O_94,N_4925,N_4961);
nand UO_95 (O_95,N_4914,N_4935);
nand UO_96 (O_96,N_4907,N_4921);
nor UO_97 (O_97,N_4979,N_4902);
and UO_98 (O_98,N_4955,N_4965);
nor UO_99 (O_99,N_4995,N_4900);
and UO_100 (O_100,N_4992,N_4974);
or UO_101 (O_101,N_4967,N_4940);
or UO_102 (O_102,N_4978,N_4928);
nand UO_103 (O_103,N_4959,N_4998);
and UO_104 (O_104,N_4975,N_4980);
xnor UO_105 (O_105,N_4998,N_4933);
nand UO_106 (O_106,N_4986,N_4939);
or UO_107 (O_107,N_4960,N_4996);
nand UO_108 (O_108,N_4912,N_4985);
and UO_109 (O_109,N_4912,N_4969);
or UO_110 (O_110,N_4963,N_4949);
nand UO_111 (O_111,N_4998,N_4938);
and UO_112 (O_112,N_4988,N_4901);
or UO_113 (O_113,N_4988,N_4932);
and UO_114 (O_114,N_4991,N_4999);
or UO_115 (O_115,N_4998,N_4971);
nor UO_116 (O_116,N_4978,N_4939);
and UO_117 (O_117,N_4950,N_4905);
nor UO_118 (O_118,N_4902,N_4998);
nand UO_119 (O_119,N_4964,N_4982);
and UO_120 (O_120,N_4956,N_4923);
and UO_121 (O_121,N_4951,N_4938);
nand UO_122 (O_122,N_4936,N_4989);
nor UO_123 (O_123,N_4908,N_4929);
or UO_124 (O_124,N_4920,N_4948);
nand UO_125 (O_125,N_4915,N_4921);
nor UO_126 (O_126,N_4927,N_4967);
or UO_127 (O_127,N_4909,N_4915);
or UO_128 (O_128,N_4974,N_4966);
and UO_129 (O_129,N_4933,N_4976);
nand UO_130 (O_130,N_4996,N_4931);
nand UO_131 (O_131,N_4963,N_4919);
and UO_132 (O_132,N_4977,N_4974);
or UO_133 (O_133,N_4988,N_4908);
or UO_134 (O_134,N_4964,N_4925);
nand UO_135 (O_135,N_4946,N_4937);
and UO_136 (O_136,N_4955,N_4967);
and UO_137 (O_137,N_4976,N_4987);
and UO_138 (O_138,N_4976,N_4942);
and UO_139 (O_139,N_4950,N_4997);
or UO_140 (O_140,N_4928,N_4983);
and UO_141 (O_141,N_4986,N_4940);
and UO_142 (O_142,N_4966,N_4926);
or UO_143 (O_143,N_4982,N_4978);
nand UO_144 (O_144,N_4900,N_4971);
nand UO_145 (O_145,N_4949,N_4998);
nor UO_146 (O_146,N_4945,N_4988);
nor UO_147 (O_147,N_4993,N_4927);
nor UO_148 (O_148,N_4949,N_4975);
nand UO_149 (O_149,N_4945,N_4996);
and UO_150 (O_150,N_4937,N_4947);
or UO_151 (O_151,N_4913,N_4995);
nand UO_152 (O_152,N_4966,N_4978);
or UO_153 (O_153,N_4969,N_4922);
nor UO_154 (O_154,N_4939,N_4956);
or UO_155 (O_155,N_4942,N_4916);
nor UO_156 (O_156,N_4956,N_4955);
or UO_157 (O_157,N_4995,N_4966);
or UO_158 (O_158,N_4976,N_4922);
and UO_159 (O_159,N_4951,N_4977);
or UO_160 (O_160,N_4945,N_4923);
nor UO_161 (O_161,N_4910,N_4979);
nor UO_162 (O_162,N_4980,N_4933);
nor UO_163 (O_163,N_4917,N_4928);
nand UO_164 (O_164,N_4924,N_4929);
or UO_165 (O_165,N_4911,N_4904);
or UO_166 (O_166,N_4935,N_4955);
nand UO_167 (O_167,N_4991,N_4939);
and UO_168 (O_168,N_4982,N_4914);
and UO_169 (O_169,N_4996,N_4949);
and UO_170 (O_170,N_4964,N_4908);
xnor UO_171 (O_171,N_4938,N_4932);
nor UO_172 (O_172,N_4964,N_4985);
nand UO_173 (O_173,N_4952,N_4908);
or UO_174 (O_174,N_4992,N_4943);
or UO_175 (O_175,N_4929,N_4983);
nand UO_176 (O_176,N_4990,N_4936);
and UO_177 (O_177,N_4941,N_4980);
and UO_178 (O_178,N_4953,N_4965);
and UO_179 (O_179,N_4935,N_4976);
nor UO_180 (O_180,N_4962,N_4977);
nand UO_181 (O_181,N_4952,N_4904);
nand UO_182 (O_182,N_4947,N_4959);
nor UO_183 (O_183,N_4929,N_4912);
and UO_184 (O_184,N_4956,N_4947);
nor UO_185 (O_185,N_4927,N_4920);
nor UO_186 (O_186,N_4977,N_4997);
nand UO_187 (O_187,N_4934,N_4958);
nor UO_188 (O_188,N_4916,N_4990);
nand UO_189 (O_189,N_4928,N_4939);
and UO_190 (O_190,N_4928,N_4988);
xnor UO_191 (O_191,N_4949,N_4919);
and UO_192 (O_192,N_4927,N_4981);
and UO_193 (O_193,N_4903,N_4907);
nand UO_194 (O_194,N_4964,N_4967);
and UO_195 (O_195,N_4980,N_4947);
nand UO_196 (O_196,N_4930,N_4979);
nor UO_197 (O_197,N_4968,N_4998);
or UO_198 (O_198,N_4950,N_4989);
nand UO_199 (O_199,N_4970,N_4990);
nor UO_200 (O_200,N_4991,N_4980);
and UO_201 (O_201,N_4900,N_4939);
or UO_202 (O_202,N_4989,N_4931);
xor UO_203 (O_203,N_4951,N_4910);
nand UO_204 (O_204,N_4967,N_4984);
and UO_205 (O_205,N_4902,N_4977);
or UO_206 (O_206,N_4903,N_4934);
nor UO_207 (O_207,N_4983,N_4998);
nor UO_208 (O_208,N_4976,N_4955);
nor UO_209 (O_209,N_4938,N_4967);
nor UO_210 (O_210,N_4992,N_4946);
xnor UO_211 (O_211,N_4955,N_4962);
nand UO_212 (O_212,N_4981,N_4998);
and UO_213 (O_213,N_4916,N_4954);
xnor UO_214 (O_214,N_4904,N_4963);
nor UO_215 (O_215,N_4954,N_4963);
or UO_216 (O_216,N_4972,N_4919);
and UO_217 (O_217,N_4915,N_4904);
or UO_218 (O_218,N_4955,N_4999);
or UO_219 (O_219,N_4979,N_4947);
nand UO_220 (O_220,N_4954,N_4925);
nor UO_221 (O_221,N_4975,N_4932);
and UO_222 (O_222,N_4989,N_4928);
and UO_223 (O_223,N_4978,N_4916);
nand UO_224 (O_224,N_4929,N_4937);
and UO_225 (O_225,N_4980,N_4935);
nor UO_226 (O_226,N_4941,N_4925);
or UO_227 (O_227,N_4946,N_4951);
and UO_228 (O_228,N_4932,N_4961);
or UO_229 (O_229,N_4910,N_4956);
and UO_230 (O_230,N_4915,N_4946);
or UO_231 (O_231,N_4962,N_4957);
nand UO_232 (O_232,N_4968,N_4985);
nor UO_233 (O_233,N_4936,N_4921);
or UO_234 (O_234,N_4913,N_4989);
nor UO_235 (O_235,N_4959,N_4996);
or UO_236 (O_236,N_4989,N_4969);
and UO_237 (O_237,N_4943,N_4914);
and UO_238 (O_238,N_4928,N_4945);
and UO_239 (O_239,N_4909,N_4924);
nand UO_240 (O_240,N_4945,N_4960);
and UO_241 (O_241,N_4935,N_4986);
xor UO_242 (O_242,N_4961,N_4942);
nor UO_243 (O_243,N_4906,N_4954);
nor UO_244 (O_244,N_4911,N_4980);
or UO_245 (O_245,N_4940,N_4905);
and UO_246 (O_246,N_4945,N_4980);
nand UO_247 (O_247,N_4938,N_4912);
nand UO_248 (O_248,N_4921,N_4928);
nor UO_249 (O_249,N_4931,N_4917);
or UO_250 (O_250,N_4906,N_4935);
nand UO_251 (O_251,N_4909,N_4949);
or UO_252 (O_252,N_4927,N_4908);
and UO_253 (O_253,N_4923,N_4970);
and UO_254 (O_254,N_4978,N_4968);
nor UO_255 (O_255,N_4973,N_4919);
or UO_256 (O_256,N_4951,N_4976);
nand UO_257 (O_257,N_4944,N_4910);
and UO_258 (O_258,N_4996,N_4983);
and UO_259 (O_259,N_4991,N_4926);
nand UO_260 (O_260,N_4914,N_4921);
nand UO_261 (O_261,N_4934,N_4974);
nand UO_262 (O_262,N_4971,N_4943);
nand UO_263 (O_263,N_4956,N_4959);
nand UO_264 (O_264,N_4924,N_4932);
xnor UO_265 (O_265,N_4925,N_4958);
nor UO_266 (O_266,N_4928,N_4901);
nor UO_267 (O_267,N_4917,N_4934);
nand UO_268 (O_268,N_4965,N_4962);
nand UO_269 (O_269,N_4947,N_4999);
and UO_270 (O_270,N_4940,N_4995);
nor UO_271 (O_271,N_4932,N_4994);
and UO_272 (O_272,N_4900,N_4918);
and UO_273 (O_273,N_4905,N_4993);
or UO_274 (O_274,N_4935,N_4968);
nand UO_275 (O_275,N_4905,N_4915);
nand UO_276 (O_276,N_4989,N_4930);
nand UO_277 (O_277,N_4973,N_4933);
nor UO_278 (O_278,N_4905,N_4927);
and UO_279 (O_279,N_4951,N_4964);
nand UO_280 (O_280,N_4996,N_4963);
and UO_281 (O_281,N_4925,N_4977);
xnor UO_282 (O_282,N_4987,N_4954);
nand UO_283 (O_283,N_4977,N_4983);
nand UO_284 (O_284,N_4962,N_4992);
or UO_285 (O_285,N_4976,N_4914);
nor UO_286 (O_286,N_4990,N_4910);
and UO_287 (O_287,N_4950,N_4998);
and UO_288 (O_288,N_4950,N_4991);
nand UO_289 (O_289,N_4944,N_4936);
nor UO_290 (O_290,N_4912,N_4966);
nand UO_291 (O_291,N_4934,N_4989);
or UO_292 (O_292,N_4923,N_4939);
or UO_293 (O_293,N_4996,N_4994);
nor UO_294 (O_294,N_4997,N_4949);
or UO_295 (O_295,N_4944,N_4943);
nand UO_296 (O_296,N_4918,N_4902);
or UO_297 (O_297,N_4997,N_4959);
or UO_298 (O_298,N_4961,N_4975);
nand UO_299 (O_299,N_4974,N_4969);
nand UO_300 (O_300,N_4918,N_4940);
nand UO_301 (O_301,N_4976,N_4962);
and UO_302 (O_302,N_4919,N_4982);
or UO_303 (O_303,N_4954,N_4970);
nor UO_304 (O_304,N_4925,N_4929);
xnor UO_305 (O_305,N_4994,N_4981);
nand UO_306 (O_306,N_4968,N_4911);
nand UO_307 (O_307,N_4985,N_4918);
or UO_308 (O_308,N_4994,N_4939);
or UO_309 (O_309,N_4950,N_4966);
and UO_310 (O_310,N_4950,N_4942);
nor UO_311 (O_311,N_4931,N_4992);
nand UO_312 (O_312,N_4919,N_4906);
nor UO_313 (O_313,N_4917,N_4927);
xor UO_314 (O_314,N_4908,N_4995);
nand UO_315 (O_315,N_4939,N_4936);
nor UO_316 (O_316,N_4949,N_4928);
xnor UO_317 (O_317,N_4908,N_4916);
nor UO_318 (O_318,N_4992,N_4933);
or UO_319 (O_319,N_4908,N_4901);
or UO_320 (O_320,N_4901,N_4927);
xnor UO_321 (O_321,N_4975,N_4969);
nor UO_322 (O_322,N_4969,N_4943);
and UO_323 (O_323,N_4917,N_4932);
or UO_324 (O_324,N_4967,N_4949);
or UO_325 (O_325,N_4920,N_4972);
nand UO_326 (O_326,N_4911,N_4918);
or UO_327 (O_327,N_4951,N_4981);
nand UO_328 (O_328,N_4977,N_4998);
and UO_329 (O_329,N_4977,N_4959);
nand UO_330 (O_330,N_4975,N_4948);
and UO_331 (O_331,N_4995,N_4955);
and UO_332 (O_332,N_4961,N_4929);
nand UO_333 (O_333,N_4908,N_4924);
nand UO_334 (O_334,N_4952,N_4981);
nor UO_335 (O_335,N_4984,N_4923);
nor UO_336 (O_336,N_4998,N_4963);
or UO_337 (O_337,N_4932,N_4900);
and UO_338 (O_338,N_4969,N_4902);
nor UO_339 (O_339,N_4922,N_4923);
and UO_340 (O_340,N_4946,N_4963);
nor UO_341 (O_341,N_4963,N_4955);
or UO_342 (O_342,N_4914,N_4942);
and UO_343 (O_343,N_4934,N_4905);
or UO_344 (O_344,N_4959,N_4989);
or UO_345 (O_345,N_4918,N_4990);
nor UO_346 (O_346,N_4954,N_4964);
nor UO_347 (O_347,N_4936,N_4997);
nor UO_348 (O_348,N_4947,N_4958);
nor UO_349 (O_349,N_4963,N_4990);
nand UO_350 (O_350,N_4908,N_4998);
xor UO_351 (O_351,N_4949,N_4924);
or UO_352 (O_352,N_4961,N_4917);
nor UO_353 (O_353,N_4970,N_4912);
nor UO_354 (O_354,N_4930,N_4969);
nand UO_355 (O_355,N_4933,N_4935);
nor UO_356 (O_356,N_4963,N_4937);
nand UO_357 (O_357,N_4903,N_4989);
nand UO_358 (O_358,N_4913,N_4925);
or UO_359 (O_359,N_4996,N_4935);
and UO_360 (O_360,N_4976,N_4991);
and UO_361 (O_361,N_4948,N_4930);
nand UO_362 (O_362,N_4950,N_4996);
or UO_363 (O_363,N_4944,N_4904);
nor UO_364 (O_364,N_4920,N_4973);
and UO_365 (O_365,N_4935,N_4984);
nor UO_366 (O_366,N_4910,N_4962);
and UO_367 (O_367,N_4966,N_4994);
and UO_368 (O_368,N_4982,N_4934);
nand UO_369 (O_369,N_4944,N_4964);
and UO_370 (O_370,N_4939,N_4969);
nand UO_371 (O_371,N_4927,N_4989);
nor UO_372 (O_372,N_4913,N_4938);
and UO_373 (O_373,N_4960,N_4921);
and UO_374 (O_374,N_4972,N_4941);
and UO_375 (O_375,N_4975,N_4981);
nand UO_376 (O_376,N_4949,N_4957);
or UO_377 (O_377,N_4923,N_4951);
nor UO_378 (O_378,N_4969,N_4938);
nor UO_379 (O_379,N_4951,N_4962);
nand UO_380 (O_380,N_4959,N_4932);
nand UO_381 (O_381,N_4907,N_4912);
nand UO_382 (O_382,N_4988,N_4998);
xor UO_383 (O_383,N_4933,N_4903);
nand UO_384 (O_384,N_4940,N_4987);
xnor UO_385 (O_385,N_4966,N_4982);
and UO_386 (O_386,N_4947,N_4941);
or UO_387 (O_387,N_4978,N_4905);
and UO_388 (O_388,N_4975,N_4984);
nand UO_389 (O_389,N_4901,N_4914);
or UO_390 (O_390,N_4917,N_4902);
nor UO_391 (O_391,N_4924,N_4997);
or UO_392 (O_392,N_4911,N_4996);
and UO_393 (O_393,N_4973,N_4924);
and UO_394 (O_394,N_4921,N_4972);
or UO_395 (O_395,N_4955,N_4910);
nor UO_396 (O_396,N_4999,N_4943);
and UO_397 (O_397,N_4944,N_4960);
or UO_398 (O_398,N_4968,N_4963);
nand UO_399 (O_399,N_4966,N_4985);
and UO_400 (O_400,N_4992,N_4937);
or UO_401 (O_401,N_4971,N_4920);
and UO_402 (O_402,N_4911,N_4999);
and UO_403 (O_403,N_4922,N_4954);
or UO_404 (O_404,N_4904,N_4946);
nand UO_405 (O_405,N_4993,N_4967);
nand UO_406 (O_406,N_4908,N_4966);
nand UO_407 (O_407,N_4941,N_4906);
nand UO_408 (O_408,N_4981,N_4990);
and UO_409 (O_409,N_4936,N_4998);
nor UO_410 (O_410,N_4976,N_4974);
nand UO_411 (O_411,N_4911,N_4947);
xnor UO_412 (O_412,N_4997,N_4903);
nor UO_413 (O_413,N_4995,N_4916);
and UO_414 (O_414,N_4998,N_4926);
nor UO_415 (O_415,N_4920,N_4970);
and UO_416 (O_416,N_4912,N_4928);
and UO_417 (O_417,N_4938,N_4929);
nor UO_418 (O_418,N_4940,N_4965);
nand UO_419 (O_419,N_4903,N_4950);
nor UO_420 (O_420,N_4937,N_4957);
nand UO_421 (O_421,N_4992,N_4995);
nor UO_422 (O_422,N_4921,N_4905);
and UO_423 (O_423,N_4927,N_4961);
or UO_424 (O_424,N_4981,N_4942);
nand UO_425 (O_425,N_4997,N_4994);
nor UO_426 (O_426,N_4989,N_4941);
xor UO_427 (O_427,N_4935,N_4911);
nor UO_428 (O_428,N_4960,N_4952);
nand UO_429 (O_429,N_4981,N_4940);
or UO_430 (O_430,N_4943,N_4909);
or UO_431 (O_431,N_4909,N_4955);
and UO_432 (O_432,N_4905,N_4967);
nand UO_433 (O_433,N_4978,N_4907);
nand UO_434 (O_434,N_4970,N_4933);
and UO_435 (O_435,N_4951,N_4940);
nor UO_436 (O_436,N_4958,N_4935);
or UO_437 (O_437,N_4938,N_4966);
nor UO_438 (O_438,N_4983,N_4944);
nor UO_439 (O_439,N_4992,N_4975);
and UO_440 (O_440,N_4981,N_4993);
and UO_441 (O_441,N_4958,N_4927);
nor UO_442 (O_442,N_4931,N_4995);
or UO_443 (O_443,N_4999,N_4949);
nor UO_444 (O_444,N_4937,N_4984);
and UO_445 (O_445,N_4994,N_4999);
and UO_446 (O_446,N_4917,N_4975);
or UO_447 (O_447,N_4917,N_4984);
or UO_448 (O_448,N_4927,N_4922);
nand UO_449 (O_449,N_4995,N_4967);
xor UO_450 (O_450,N_4988,N_4971);
nand UO_451 (O_451,N_4968,N_4932);
nor UO_452 (O_452,N_4953,N_4974);
or UO_453 (O_453,N_4931,N_4997);
and UO_454 (O_454,N_4921,N_4908);
or UO_455 (O_455,N_4979,N_4939);
nor UO_456 (O_456,N_4989,N_4955);
and UO_457 (O_457,N_4938,N_4942);
nand UO_458 (O_458,N_4922,N_4920);
or UO_459 (O_459,N_4952,N_4902);
nor UO_460 (O_460,N_4949,N_4960);
or UO_461 (O_461,N_4986,N_4984);
nor UO_462 (O_462,N_4990,N_4902);
or UO_463 (O_463,N_4969,N_4948);
nand UO_464 (O_464,N_4995,N_4930);
xnor UO_465 (O_465,N_4924,N_4996);
or UO_466 (O_466,N_4950,N_4968);
or UO_467 (O_467,N_4973,N_4958);
nand UO_468 (O_468,N_4984,N_4922);
nor UO_469 (O_469,N_4938,N_4944);
or UO_470 (O_470,N_4967,N_4976);
nor UO_471 (O_471,N_4985,N_4986);
xor UO_472 (O_472,N_4999,N_4933);
nand UO_473 (O_473,N_4907,N_4930);
and UO_474 (O_474,N_4982,N_4951);
nand UO_475 (O_475,N_4905,N_4989);
and UO_476 (O_476,N_4903,N_4984);
or UO_477 (O_477,N_4955,N_4927);
xor UO_478 (O_478,N_4914,N_4915);
nand UO_479 (O_479,N_4998,N_4906);
and UO_480 (O_480,N_4980,N_4954);
nand UO_481 (O_481,N_4988,N_4985);
and UO_482 (O_482,N_4958,N_4976);
or UO_483 (O_483,N_4916,N_4992);
nor UO_484 (O_484,N_4934,N_4960);
nor UO_485 (O_485,N_4988,N_4969);
xor UO_486 (O_486,N_4906,N_4924);
nor UO_487 (O_487,N_4973,N_4906);
nor UO_488 (O_488,N_4963,N_4960);
or UO_489 (O_489,N_4990,N_4903);
or UO_490 (O_490,N_4912,N_4997);
or UO_491 (O_491,N_4923,N_4909);
nand UO_492 (O_492,N_4941,N_4911);
xor UO_493 (O_493,N_4918,N_4978);
nor UO_494 (O_494,N_4984,N_4994);
and UO_495 (O_495,N_4909,N_4936);
nand UO_496 (O_496,N_4975,N_4950);
nand UO_497 (O_497,N_4907,N_4953);
and UO_498 (O_498,N_4929,N_4978);
nor UO_499 (O_499,N_4967,N_4943);
nor UO_500 (O_500,N_4911,N_4979);
or UO_501 (O_501,N_4968,N_4975);
and UO_502 (O_502,N_4986,N_4921);
nor UO_503 (O_503,N_4923,N_4999);
and UO_504 (O_504,N_4935,N_4925);
nor UO_505 (O_505,N_4936,N_4950);
nor UO_506 (O_506,N_4937,N_4997);
or UO_507 (O_507,N_4994,N_4965);
nor UO_508 (O_508,N_4950,N_4900);
and UO_509 (O_509,N_4933,N_4917);
and UO_510 (O_510,N_4948,N_4989);
or UO_511 (O_511,N_4915,N_4983);
nand UO_512 (O_512,N_4938,N_4941);
nor UO_513 (O_513,N_4903,N_4952);
nand UO_514 (O_514,N_4964,N_4903);
or UO_515 (O_515,N_4989,N_4953);
or UO_516 (O_516,N_4983,N_4920);
nand UO_517 (O_517,N_4991,N_4952);
nand UO_518 (O_518,N_4955,N_4988);
or UO_519 (O_519,N_4996,N_4955);
nand UO_520 (O_520,N_4954,N_4948);
nor UO_521 (O_521,N_4966,N_4927);
and UO_522 (O_522,N_4919,N_4981);
nor UO_523 (O_523,N_4919,N_4908);
or UO_524 (O_524,N_4943,N_4904);
or UO_525 (O_525,N_4927,N_4969);
and UO_526 (O_526,N_4914,N_4965);
xnor UO_527 (O_527,N_4959,N_4973);
or UO_528 (O_528,N_4931,N_4982);
or UO_529 (O_529,N_4987,N_4986);
and UO_530 (O_530,N_4936,N_4970);
nor UO_531 (O_531,N_4977,N_4933);
or UO_532 (O_532,N_4914,N_4920);
nor UO_533 (O_533,N_4966,N_4955);
or UO_534 (O_534,N_4984,N_4957);
nor UO_535 (O_535,N_4996,N_4929);
and UO_536 (O_536,N_4945,N_4914);
nand UO_537 (O_537,N_4922,N_4991);
nor UO_538 (O_538,N_4958,N_4987);
or UO_539 (O_539,N_4962,N_4921);
and UO_540 (O_540,N_4969,N_4997);
nor UO_541 (O_541,N_4914,N_4997);
xor UO_542 (O_542,N_4918,N_4952);
and UO_543 (O_543,N_4975,N_4965);
nand UO_544 (O_544,N_4964,N_4957);
nand UO_545 (O_545,N_4997,N_4920);
and UO_546 (O_546,N_4944,N_4970);
or UO_547 (O_547,N_4952,N_4927);
nor UO_548 (O_548,N_4945,N_4986);
and UO_549 (O_549,N_4923,N_4912);
xor UO_550 (O_550,N_4971,N_4975);
xnor UO_551 (O_551,N_4994,N_4909);
nand UO_552 (O_552,N_4979,N_4914);
xnor UO_553 (O_553,N_4921,N_4973);
and UO_554 (O_554,N_4916,N_4970);
or UO_555 (O_555,N_4972,N_4914);
and UO_556 (O_556,N_4945,N_4998);
nand UO_557 (O_557,N_4958,N_4970);
and UO_558 (O_558,N_4979,N_4956);
or UO_559 (O_559,N_4947,N_4901);
nor UO_560 (O_560,N_4948,N_4999);
and UO_561 (O_561,N_4944,N_4916);
nand UO_562 (O_562,N_4967,N_4992);
or UO_563 (O_563,N_4971,N_4948);
xor UO_564 (O_564,N_4911,N_4945);
nor UO_565 (O_565,N_4921,N_4991);
or UO_566 (O_566,N_4901,N_4942);
and UO_567 (O_567,N_4938,N_4957);
nor UO_568 (O_568,N_4901,N_4965);
nand UO_569 (O_569,N_4927,N_4932);
nand UO_570 (O_570,N_4935,N_4957);
or UO_571 (O_571,N_4998,N_4927);
nand UO_572 (O_572,N_4955,N_4942);
nor UO_573 (O_573,N_4981,N_4978);
or UO_574 (O_574,N_4972,N_4932);
nor UO_575 (O_575,N_4946,N_4932);
nand UO_576 (O_576,N_4975,N_4954);
nand UO_577 (O_577,N_4972,N_4944);
xnor UO_578 (O_578,N_4941,N_4936);
or UO_579 (O_579,N_4936,N_4965);
xnor UO_580 (O_580,N_4942,N_4900);
or UO_581 (O_581,N_4982,N_4900);
or UO_582 (O_582,N_4918,N_4934);
nand UO_583 (O_583,N_4928,N_4920);
and UO_584 (O_584,N_4966,N_4941);
nand UO_585 (O_585,N_4922,N_4957);
and UO_586 (O_586,N_4951,N_4956);
and UO_587 (O_587,N_4903,N_4945);
and UO_588 (O_588,N_4924,N_4967);
and UO_589 (O_589,N_4908,N_4922);
nor UO_590 (O_590,N_4903,N_4971);
xor UO_591 (O_591,N_4954,N_4934);
nand UO_592 (O_592,N_4926,N_4924);
xnor UO_593 (O_593,N_4920,N_4924);
nand UO_594 (O_594,N_4941,N_4974);
nor UO_595 (O_595,N_4958,N_4928);
or UO_596 (O_596,N_4944,N_4955);
or UO_597 (O_597,N_4994,N_4903);
nor UO_598 (O_598,N_4915,N_4961);
and UO_599 (O_599,N_4953,N_4926);
or UO_600 (O_600,N_4943,N_4923);
or UO_601 (O_601,N_4990,N_4968);
and UO_602 (O_602,N_4984,N_4974);
and UO_603 (O_603,N_4971,N_4979);
and UO_604 (O_604,N_4946,N_4976);
or UO_605 (O_605,N_4937,N_4952);
or UO_606 (O_606,N_4933,N_4951);
and UO_607 (O_607,N_4918,N_4910);
or UO_608 (O_608,N_4960,N_4908);
xor UO_609 (O_609,N_4938,N_4996);
xor UO_610 (O_610,N_4993,N_4952);
xor UO_611 (O_611,N_4949,N_4990);
nand UO_612 (O_612,N_4912,N_4920);
xnor UO_613 (O_613,N_4918,N_4957);
nor UO_614 (O_614,N_4940,N_4959);
nand UO_615 (O_615,N_4920,N_4994);
xor UO_616 (O_616,N_4919,N_4997);
nand UO_617 (O_617,N_4938,N_4909);
xnor UO_618 (O_618,N_4969,N_4900);
nand UO_619 (O_619,N_4973,N_4948);
nand UO_620 (O_620,N_4968,N_4949);
nor UO_621 (O_621,N_4993,N_4947);
or UO_622 (O_622,N_4991,N_4938);
and UO_623 (O_623,N_4952,N_4907);
and UO_624 (O_624,N_4932,N_4958);
nand UO_625 (O_625,N_4939,N_4952);
or UO_626 (O_626,N_4967,N_4936);
nand UO_627 (O_627,N_4929,N_4909);
nand UO_628 (O_628,N_4926,N_4921);
or UO_629 (O_629,N_4992,N_4986);
xor UO_630 (O_630,N_4912,N_4901);
and UO_631 (O_631,N_4944,N_4935);
nand UO_632 (O_632,N_4998,N_4907);
and UO_633 (O_633,N_4923,N_4993);
or UO_634 (O_634,N_4925,N_4909);
xnor UO_635 (O_635,N_4964,N_4955);
nor UO_636 (O_636,N_4904,N_4971);
nand UO_637 (O_637,N_4916,N_4984);
nand UO_638 (O_638,N_4974,N_4912);
nand UO_639 (O_639,N_4960,N_4922);
or UO_640 (O_640,N_4970,N_4993);
and UO_641 (O_641,N_4907,N_4963);
xnor UO_642 (O_642,N_4959,N_4950);
nand UO_643 (O_643,N_4909,N_4902);
nor UO_644 (O_644,N_4980,N_4950);
nor UO_645 (O_645,N_4920,N_4936);
nand UO_646 (O_646,N_4928,N_4982);
and UO_647 (O_647,N_4955,N_4998);
xor UO_648 (O_648,N_4958,N_4918);
nor UO_649 (O_649,N_4928,N_4946);
or UO_650 (O_650,N_4986,N_4909);
and UO_651 (O_651,N_4975,N_4963);
xor UO_652 (O_652,N_4942,N_4944);
nor UO_653 (O_653,N_4994,N_4929);
nor UO_654 (O_654,N_4969,N_4970);
xor UO_655 (O_655,N_4952,N_4959);
nand UO_656 (O_656,N_4995,N_4948);
nand UO_657 (O_657,N_4968,N_4999);
nand UO_658 (O_658,N_4969,N_4987);
or UO_659 (O_659,N_4932,N_4906);
xnor UO_660 (O_660,N_4994,N_4995);
xor UO_661 (O_661,N_4901,N_4918);
nor UO_662 (O_662,N_4953,N_4968);
xor UO_663 (O_663,N_4916,N_4920);
nor UO_664 (O_664,N_4962,N_4922);
and UO_665 (O_665,N_4909,N_4916);
nor UO_666 (O_666,N_4917,N_4967);
or UO_667 (O_667,N_4996,N_4974);
xnor UO_668 (O_668,N_4980,N_4972);
nor UO_669 (O_669,N_4930,N_4927);
or UO_670 (O_670,N_4997,N_4984);
xnor UO_671 (O_671,N_4984,N_4929);
nor UO_672 (O_672,N_4949,N_4931);
nand UO_673 (O_673,N_4928,N_4925);
or UO_674 (O_674,N_4959,N_4915);
nor UO_675 (O_675,N_4939,N_4995);
xor UO_676 (O_676,N_4938,N_4933);
nand UO_677 (O_677,N_4952,N_4987);
nor UO_678 (O_678,N_4943,N_4955);
nor UO_679 (O_679,N_4937,N_4938);
nor UO_680 (O_680,N_4953,N_4975);
xnor UO_681 (O_681,N_4981,N_4965);
or UO_682 (O_682,N_4999,N_4905);
nand UO_683 (O_683,N_4912,N_4973);
and UO_684 (O_684,N_4975,N_4909);
and UO_685 (O_685,N_4954,N_4953);
and UO_686 (O_686,N_4980,N_4920);
or UO_687 (O_687,N_4984,N_4998);
xnor UO_688 (O_688,N_4997,N_4943);
nand UO_689 (O_689,N_4950,N_4944);
or UO_690 (O_690,N_4959,N_4999);
and UO_691 (O_691,N_4997,N_4922);
nor UO_692 (O_692,N_4943,N_4947);
nor UO_693 (O_693,N_4954,N_4926);
xor UO_694 (O_694,N_4967,N_4915);
nand UO_695 (O_695,N_4960,N_4932);
and UO_696 (O_696,N_4943,N_4972);
nor UO_697 (O_697,N_4958,N_4913);
nor UO_698 (O_698,N_4913,N_4930);
xnor UO_699 (O_699,N_4966,N_4970);
nor UO_700 (O_700,N_4929,N_4980);
xnor UO_701 (O_701,N_4988,N_4956);
nand UO_702 (O_702,N_4905,N_4970);
or UO_703 (O_703,N_4949,N_4946);
nor UO_704 (O_704,N_4931,N_4945);
and UO_705 (O_705,N_4914,N_4994);
or UO_706 (O_706,N_4951,N_4907);
or UO_707 (O_707,N_4941,N_4960);
nand UO_708 (O_708,N_4991,N_4984);
and UO_709 (O_709,N_4904,N_4961);
and UO_710 (O_710,N_4988,N_4978);
nand UO_711 (O_711,N_4978,N_4938);
nand UO_712 (O_712,N_4990,N_4938);
nand UO_713 (O_713,N_4930,N_4903);
nor UO_714 (O_714,N_4979,N_4978);
nand UO_715 (O_715,N_4958,N_4974);
nand UO_716 (O_716,N_4927,N_4915);
nor UO_717 (O_717,N_4913,N_4961);
nand UO_718 (O_718,N_4995,N_4927);
nor UO_719 (O_719,N_4952,N_4932);
and UO_720 (O_720,N_4979,N_4900);
xnor UO_721 (O_721,N_4924,N_4960);
and UO_722 (O_722,N_4962,N_4997);
nor UO_723 (O_723,N_4975,N_4943);
nand UO_724 (O_724,N_4983,N_4909);
nand UO_725 (O_725,N_4907,N_4984);
or UO_726 (O_726,N_4904,N_4949);
nand UO_727 (O_727,N_4938,N_4901);
xnor UO_728 (O_728,N_4909,N_4988);
xnor UO_729 (O_729,N_4947,N_4961);
nor UO_730 (O_730,N_4958,N_4969);
nand UO_731 (O_731,N_4911,N_4981);
or UO_732 (O_732,N_4936,N_4934);
xor UO_733 (O_733,N_4992,N_4963);
or UO_734 (O_734,N_4933,N_4908);
or UO_735 (O_735,N_4939,N_4983);
nor UO_736 (O_736,N_4934,N_4933);
nor UO_737 (O_737,N_4973,N_4998);
or UO_738 (O_738,N_4953,N_4945);
or UO_739 (O_739,N_4909,N_4907);
and UO_740 (O_740,N_4950,N_4941);
and UO_741 (O_741,N_4902,N_4929);
and UO_742 (O_742,N_4946,N_4908);
nand UO_743 (O_743,N_4950,N_4957);
and UO_744 (O_744,N_4947,N_4921);
or UO_745 (O_745,N_4985,N_4937);
nor UO_746 (O_746,N_4993,N_4974);
nor UO_747 (O_747,N_4993,N_4988);
and UO_748 (O_748,N_4911,N_4924);
nor UO_749 (O_749,N_4947,N_4923);
nand UO_750 (O_750,N_4995,N_4961);
nor UO_751 (O_751,N_4990,N_4991);
nor UO_752 (O_752,N_4910,N_4942);
and UO_753 (O_753,N_4910,N_4983);
or UO_754 (O_754,N_4969,N_4984);
nor UO_755 (O_755,N_4966,N_4922);
xor UO_756 (O_756,N_4929,N_4958);
and UO_757 (O_757,N_4997,N_4998);
and UO_758 (O_758,N_4973,N_4962);
or UO_759 (O_759,N_4997,N_4956);
nor UO_760 (O_760,N_4945,N_4981);
nand UO_761 (O_761,N_4900,N_4947);
nor UO_762 (O_762,N_4941,N_4902);
nor UO_763 (O_763,N_4938,N_4982);
nor UO_764 (O_764,N_4966,N_4973);
or UO_765 (O_765,N_4951,N_4993);
nor UO_766 (O_766,N_4907,N_4957);
nor UO_767 (O_767,N_4956,N_4986);
and UO_768 (O_768,N_4918,N_4904);
and UO_769 (O_769,N_4954,N_4921);
and UO_770 (O_770,N_4975,N_4976);
nand UO_771 (O_771,N_4960,N_4983);
nor UO_772 (O_772,N_4917,N_4994);
and UO_773 (O_773,N_4932,N_4943);
or UO_774 (O_774,N_4907,N_4977);
or UO_775 (O_775,N_4970,N_4909);
or UO_776 (O_776,N_4974,N_4907);
nand UO_777 (O_777,N_4994,N_4913);
and UO_778 (O_778,N_4980,N_4953);
nor UO_779 (O_779,N_4908,N_4948);
nand UO_780 (O_780,N_4972,N_4975);
and UO_781 (O_781,N_4954,N_4972);
nand UO_782 (O_782,N_4944,N_4988);
nor UO_783 (O_783,N_4933,N_4957);
nand UO_784 (O_784,N_4985,N_4958);
nand UO_785 (O_785,N_4949,N_4911);
or UO_786 (O_786,N_4920,N_4931);
or UO_787 (O_787,N_4944,N_4995);
nor UO_788 (O_788,N_4918,N_4913);
or UO_789 (O_789,N_4990,N_4912);
nand UO_790 (O_790,N_4916,N_4921);
nor UO_791 (O_791,N_4999,N_4979);
and UO_792 (O_792,N_4981,N_4974);
nor UO_793 (O_793,N_4933,N_4911);
or UO_794 (O_794,N_4995,N_4960);
and UO_795 (O_795,N_4913,N_4975);
nor UO_796 (O_796,N_4972,N_4951);
nor UO_797 (O_797,N_4981,N_4931);
and UO_798 (O_798,N_4933,N_4944);
nor UO_799 (O_799,N_4909,N_4919);
and UO_800 (O_800,N_4981,N_4973);
and UO_801 (O_801,N_4995,N_4978);
nor UO_802 (O_802,N_4965,N_4977);
nand UO_803 (O_803,N_4949,N_4977);
or UO_804 (O_804,N_4992,N_4918);
nor UO_805 (O_805,N_4977,N_4918);
and UO_806 (O_806,N_4978,N_4973);
and UO_807 (O_807,N_4957,N_4910);
and UO_808 (O_808,N_4956,N_4933);
nand UO_809 (O_809,N_4916,N_4963);
and UO_810 (O_810,N_4925,N_4934);
or UO_811 (O_811,N_4932,N_4953);
xnor UO_812 (O_812,N_4962,N_4940);
xor UO_813 (O_813,N_4921,N_4980);
nor UO_814 (O_814,N_4911,N_4916);
nand UO_815 (O_815,N_4912,N_4965);
or UO_816 (O_816,N_4935,N_4940);
xor UO_817 (O_817,N_4953,N_4983);
or UO_818 (O_818,N_4902,N_4955);
nor UO_819 (O_819,N_4927,N_4965);
and UO_820 (O_820,N_4963,N_4926);
nor UO_821 (O_821,N_4933,N_4954);
and UO_822 (O_822,N_4948,N_4959);
nand UO_823 (O_823,N_4908,N_4945);
and UO_824 (O_824,N_4900,N_4992);
nand UO_825 (O_825,N_4972,N_4996);
nor UO_826 (O_826,N_4911,N_4976);
and UO_827 (O_827,N_4957,N_4939);
nor UO_828 (O_828,N_4905,N_4975);
or UO_829 (O_829,N_4961,N_4968);
nand UO_830 (O_830,N_4902,N_4940);
and UO_831 (O_831,N_4985,N_4916);
or UO_832 (O_832,N_4999,N_4998);
and UO_833 (O_833,N_4967,N_4906);
and UO_834 (O_834,N_4980,N_4938);
nand UO_835 (O_835,N_4964,N_4987);
nor UO_836 (O_836,N_4948,N_4994);
and UO_837 (O_837,N_4936,N_4903);
and UO_838 (O_838,N_4950,N_4908);
or UO_839 (O_839,N_4992,N_4908);
nand UO_840 (O_840,N_4932,N_4941);
xnor UO_841 (O_841,N_4986,N_4957);
nand UO_842 (O_842,N_4984,N_4945);
and UO_843 (O_843,N_4914,N_4968);
and UO_844 (O_844,N_4918,N_4991);
and UO_845 (O_845,N_4909,N_4985);
and UO_846 (O_846,N_4911,N_4915);
nor UO_847 (O_847,N_4954,N_4990);
nand UO_848 (O_848,N_4927,N_4990);
or UO_849 (O_849,N_4967,N_4911);
or UO_850 (O_850,N_4911,N_4983);
nor UO_851 (O_851,N_4991,N_4983);
and UO_852 (O_852,N_4959,N_4967);
and UO_853 (O_853,N_4923,N_4908);
nor UO_854 (O_854,N_4949,N_4908);
nand UO_855 (O_855,N_4936,N_4916);
xnor UO_856 (O_856,N_4943,N_4968);
nand UO_857 (O_857,N_4938,N_4985);
or UO_858 (O_858,N_4972,N_4922);
nand UO_859 (O_859,N_4924,N_4912);
and UO_860 (O_860,N_4922,N_4948);
nand UO_861 (O_861,N_4989,N_4944);
or UO_862 (O_862,N_4902,N_4995);
nand UO_863 (O_863,N_4911,N_4922);
nor UO_864 (O_864,N_4933,N_4983);
or UO_865 (O_865,N_4936,N_4979);
xor UO_866 (O_866,N_4926,N_4946);
or UO_867 (O_867,N_4949,N_4932);
or UO_868 (O_868,N_4907,N_4908);
and UO_869 (O_869,N_4986,N_4928);
nor UO_870 (O_870,N_4990,N_4982);
and UO_871 (O_871,N_4982,N_4905);
and UO_872 (O_872,N_4931,N_4922);
and UO_873 (O_873,N_4922,N_4963);
and UO_874 (O_874,N_4970,N_4942);
or UO_875 (O_875,N_4945,N_4972);
xor UO_876 (O_876,N_4933,N_4945);
and UO_877 (O_877,N_4941,N_4903);
and UO_878 (O_878,N_4981,N_4957);
nor UO_879 (O_879,N_4970,N_4961);
nand UO_880 (O_880,N_4974,N_4935);
and UO_881 (O_881,N_4934,N_4927);
xor UO_882 (O_882,N_4910,N_4966);
and UO_883 (O_883,N_4993,N_4939);
and UO_884 (O_884,N_4945,N_4958);
nor UO_885 (O_885,N_4946,N_4912);
nand UO_886 (O_886,N_4989,N_4957);
nand UO_887 (O_887,N_4943,N_4905);
nand UO_888 (O_888,N_4996,N_4904);
nor UO_889 (O_889,N_4962,N_4969);
nand UO_890 (O_890,N_4970,N_4989);
and UO_891 (O_891,N_4958,N_4975);
nor UO_892 (O_892,N_4942,N_4979);
nand UO_893 (O_893,N_4917,N_4910);
xor UO_894 (O_894,N_4960,N_4942);
xor UO_895 (O_895,N_4917,N_4908);
or UO_896 (O_896,N_4921,N_4922);
nand UO_897 (O_897,N_4905,N_4963);
and UO_898 (O_898,N_4997,N_4985);
nand UO_899 (O_899,N_4912,N_4984);
and UO_900 (O_900,N_4913,N_4927);
and UO_901 (O_901,N_4985,N_4975);
and UO_902 (O_902,N_4954,N_4932);
xor UO_903 (O_903,N_4991,N_4997);
nor UO_904 (O_904,N_4906,N_4969);
and UO_905 (O_905,N_4913,N_4996);
or UO_906 (O_906,N_4954,N_4942);
nor UO_907 (O_907,N_4988,N_4974);
nand UO_908 (O_908,N_4988,N_4942);
nand UO_909 (O_909,N_4920,N_4996);
or UO_910 (O_910,N_4913,N_4974);
nand UO_911 (O_911,N_4968,N_4972);
and UO_912 (O_912,N_4980,N_4951);
and UO_913 (O_913,N_4923,N_4917);
nor UO_914 (O_914,N_4980,N_4983);
and UO_915 (O_915,N_4900,N_4999);
nand UO_916 (O_916,N_4939,N_4909);
nor UO_917 (O_917,N_4994,N_4908);
xnor UO_918 (O_918,N_4929,N_4939);
nand UO_919 (O_919,N_4985,N_4970);
or UO_920 (O_920,N_4934,N_4972);
nor UO_921 (O_921,N_4962,N_4978);
and UO_922 (O_922,N_4994,N_4954);
nand UO_923 (O_923,N_4990,N_4985);
nand UO_924 (O_924,N_4900,N_4994);
nor UO_925 (O_925,N_4931,N_4900);
or UO_926 (O_926,N_4932,N_4957);
xnor UO_927 (O_927,N_4975,N_4970);
or UO_928 (O_928,N_4978,N_4914);
and UO_929 (O_929,N_4930,N_4932);
nand UO_930 (O_930,N_4937,N_4922);
or UO_931 (O_931,N_4920,N_4935);
or UO_932 (O_932,N_4954,N_4997);
or UO_933 (O_933,N_4907,N_4962);
or UO_934 (O_934,N_4958,N_4912);
xor UO_935 (O_935,N_4911,N_4930);
nor UO_936 (O_936,N_4939,N_4987);
and UO_937 (O_937,N_4929,N_4936);
and UO_938 (O_938,N_4986,N_4904);
nor UO_939 (O_939,N_4958,N_4942);
nand UO_940 (O_940,N_4980,N_4981);
nor UO_941 (O_941,N_4929,N_4928);
and UO_942 (O_942,N_4902,N_4920);
or UO_943 (O_943,N_4928,N_4952);
nand UO_944 (O_944,N_4902,N_4957);
nand UO_945 (O_945,N_4983,N_4949);
and UO_946 (O_946,N_4998,N_4964);
nor UO_947 (O_947,N_4979,N_4944);
and UO_948 (O_948,N_4961,N_4972);
or UO_949 (O_949,N_4918,N_4941);
or UO_950 (O_950,N_4978,N_4919);
and UO_951 (O_951,N_4947,N_4978);
and UO_952 (O_952,N_4996,N_4906);
nand UO_953 (O_953,N_4946,N_4972);
and UO_954 (O_954,N_4956,N_4949);
nand UO_955 (O_955,N_4976,N_4940);
or UO_956 (O_956,N_4913,N_4969);
xnor UO_957 (O_957,N_4984,N_4942);
nor UO_958 (O_958,N_4928,N_4926);
nor UO_959 (O_959,N_4910,N_4905);
and UO_960 (O_960,N_4988,N_4940);
or UO_961 (O_961,N_4937,N_4970);
xnor UO_962 (O_962,N_4974,N_4980);
nand UO_963 (O_963,N_4958,N_4971);
nor UO_964 (O_964,N_4939,N_4968);
and UO_965 (O_965,N_4905,N_4983);
nand UO_966 (O_966,N_4904,N_4998);
xnor UO_967 (O_967,N_4955,N_4930);
or UO_968 (O_968,N_4950,N_4999);
nor UO_969 (O_969,N_4957,N_4966);
or UO_970 (O_970,N_4977,N_4967);
xnor UO_971 (O_971,N_4981,N_4943);
nor UO_972 (O_972,N_4942,N_4905);
or UO_973 (O_973,N_4935,N_4978);
nand UO_974 (O_974,N_4964,N_4932);
or UO_975 (O_975,N_4968,N_4994);
nor UO_976 (O_976,N_4947,N_4915);
or UO_977 (O_977,N_4926,N_4911);
nand UO_978 (O_978,N_4970,N_4939);
nand UO_979 (O_979,N_4927,N_4983);
nand UO_980 (O_980,N_4942,N_4953);
xor UO_981 (O_981,N_4907,N_4942);
xnor UO_982 (O_982,N_4946,N_4978);
and UO_983 (O_983,N_4955,N_4925);
nand UO_984 (O_984,N_4975,N_4952);
and UO_985 (O_985,N_4975,N_4944);
nor UO_986 (O_986,N_4992,N_4973);
or UO_987 (O_987,N_4942,N_4911);
or UO_988 (O_988,N_4943,N_4996);
and UO_989 (O_989,N_4939,N_4950);
nor UO_990 (O_990,N_4980,N_4969);
and UO_991 (O_991,N_4974,N_4905);
and UO_992 (O_992,N_4977,N_4900);
or UO_993 (O_993,N_4929,N_4971);
nand UO_994 (O_994,N_4956,N_4921);
or UO_995 (O_995,N_4968,N_4984);
nand UO_996 (O_996,N_4961,N_4971);
or UO_997 (O_997,N_4943,N_4930);
and UO_998 (O_998,N_4964,N_4956);
nand UO_999 (O_999,N_4936,N_4984);
endmodule