module basic_3000_30000_3500_60_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_2994,In_2839);
and U1 (N_1,In_2898,In_2387);
xor U2 (N_2,In_324,In_1408);
nor U3 (N_3,In_650,In_692);
or U4 (N_4,In_1761,In_815);
xor U5 (N_5,In_771,In_327);
nor U6 (N_6,In_1936,In_2763);
xnor U7 (N_7,In_1698,In_2629);
nand U8 (N_8,In_1289,In_2381);
xnor U9 (N_9,In_1798,In_2847);
nand U10 (N_10,In_2097,In_2125);
xor U11 (N_11,In_2045,In_2832);
nor U12 (N_12,In_1590,In_2592);
or U13 (N_13,In_1328,In_2121);
nor U14 (N_14,In_940,In_1640);
or U15 (N_15,In_5,In_2162);
and U16 (N_16,In_206,In_1536);
nor U17 (N_17,In_2697,In_200);
xor U18 (N_18,In_2671,In_2090);
nor U19 (N_19,In_833,In_2730);
xnor U20 (N_20,In_797,In_2739);
xnor U21 (N_21,In_1876,In_632);
xnor U22 (N_22,In_1025,In_1589);
nand U23 (N_23,In_757,In_1304);
nand U24 (N_24,In_686,In_223);
nand U25 (N_25,In_1276,In_1967);
nand U26 (N_26,In_398,In_1181);
nand U27 (N_27,In_256,In_777);
xnor U28 (N_28,In_1800,In_2618);
nand U29 (N_29,In_994,In_2063);
nand U30 (N_30,In_787,In_1460);
xnor U31 (N_31,In_2767,In_456);
nor U32 (N_32,In_847,In_1909);
nand U33 (N_33,In_441,In_1065);
nand U34 (N_34,In_2738,In_919);
and U35 (N_35,In_2712,In_2153);
nand U36 (N_36,In_2519,In_1133);
xnor U37 (N_37,In_460,In_1960);
and U38 (N_38,In_187,In_458);
or U39 (N_39,In_2988,In_512);
and U40 (N_40,In_720,In_1817);
or U41 (N_41,In_684,In_1485);
xnor U42 (N_42,In_338,In_80);
xor U43 (N_43,In_2585,In_2656);
nand U44 (N_44,In_1937,In_1769);
or U45 (N_45,In_190,In_390);
nand U46 (N_46,In_2302,In_953);
xnor U47 (N_47,In_2882,In_1185);
xnor U48 (N_48,In_936,In_774);
xnor U49 (N_49,In_2559,In_1418);
nand U50 (N_50,In_2423,In_1260);
or U51 (N_51,In_2251,In_2345);
and U52 (N_52,In_1802,In_471);
nor U53 (N_53,In_1400,In_1495);
or U54 (N_54,In_993,In_1131);
nor U55 (N_55,In_1988,In_128);
xor U56 (N_56,In_1084,In_1700);
xnor U57 (N_57,In_1374,In_2610);
nor U58 (N_58,In_1666,In_1746);
and U59 (N_59,In_1452,In_1480);
xnor U60 (N_60,In_149,In_2427);
or U61 (N_61,In_1193,In_153);
nor U62 (N_62,In_1704,In_1266);
nor U63 (N_63,In_1015,In_2052);
and U64 (N_64,In_1337,In_2866);
and U65 (N_65,In_615,In_2737);
nor U66 (N_66,In_1339,In_2714);
xor U67 (N_67,In_17,In_600);
xnor U68 (N_68,In_1413,In_385);
and U69 (N_69,In_1101,In_843);
xnor U70 (N_70,In_860,In_595);
or U71 (N_71,In_932,In_467);
xnor U72 (N_72,In_13,In_2367);
or U73 (N_73,In_53,In_2682);
nand U74 (N_74,In_2782,In_322);
and U75 (N_75,In_1865,In_895);
nor U76 (N_76,In_2711,In_2893);
xnor U77 (N_77,In_1889,In_2088);
nor U78 (N_78,In_2932,In_2168);
xnor U79 (N_79,In_2337,In_1257);
or U80 (N_80,In_1173,In_1394);
or U81 (N_81,In_782,In_689);
or U82 (N_82,In_363,In_2013);
or U83 (N_83,In_1362,In_75);
xnor U84 (N_84,In_427,In_301);
and U85 (N_85,In_52,In_640);
and U86 (N_86,In_1166,In_2999);
and U87 (N_87,In_359,In_2580);
or U88 (N_88,In_2201,In_2222);
and U89 (N_89,In_1252,In_1285);
xor U90 (N_90,In_67,In_1161);
xnor U91 (N_91,In_59,In_1931);
and U92 (N_92,In_1110,In_1508);
and U93 (N_93,In_1493,In_2742);
xnor U94 (N_94,In_1719,In_243);
and U95 (N_95,In_2323,In_1728);
and U96 (N_96,In_1669,In_924);
and U97 (N_97,In_493,In_2528);
nor U98 (N_98,In_1831,In_2516);
nor U99 (N_99,In_2616,In_2385);
xor U100 (N_100,In_1896,In_2785);
nor U101 (N_101,In_2129,In_2281);
nor U102 (N_102,In_150,In_145);
nor U103 (N_103,In_2224,In_391);
and U104 (N_104,In_2192,In_1690);
xnor U105 (N_105,In_1016,In_821);
xnor U106 (N_106,In_412,In_1273);
xor U107 (N_107,In_2664,In_2725);
nand U108 (N_108,In_1355,In_1816);
and U109 (N_109,In_1819,In_22);
xor U110 (N_110,In_1612,In_660);
nor U111 (N_111,In_1447,In_1781);
and U112 (N_112,In_725,In_534);
nand U113 (N_113,In_2700,In_930);
or U114 (N_114,In_1822,In_2996);
nor U115 (N_115,In_1435,In_231);
nand U116 (N_116,In_742,In_2661);
and U117 (N_117,In_2987,In_2388);
nor U118 (N_118,In_2096,In_1987);
nand U119 (N_119,In_2641,In_1233);
nor U120 (N_120,In_1673,In_64);
nor U121 (N_121,In_942,In_2284);
or U122 (N_122,In_244,In_1384);
and U123 (N_123,In_1727,In_2023);
nand U124 (N_124,In_869,In_2010);
nand U125 (N_125,In_1202,In_2394);
xnor U126 (N_126,In_446,In_197);
nand U127 (N_127,In_2309,In_2139);
nor U128 (N_128,In_482,In_587);
nand U129 (N_129,In_1887,In_1620);
xor U130 (N_130,In_550,In_1363);
nand U131 (N_131,In_1299,In_66);
xnor U132 (N_132,In_1614,In_1130);
and U133 (N_133,In_872,In_2546);
and U134 (N_134,In_2921,In_681);
xnor U135 (N_135,In_2867,In_1208);
or U136 (N_136,In_2726,In_2286);
and U137 (N_137,In_2484,In_879);
nor U138 (N_138,In_2499,In_189);
nor U139 (N_139,In_1848,In_1102);
xnor U140 (N_140,In_2326,In_2699);
and U141 (N_141,In_1550,In_1340);
or U142 (N_142,In_2231,In_735);
or U143 (N_143,In_1502,In_960);
nor U144 (N_144,In_367,In_1079);
nor U145 (N_145,In_839,In_2608);
or U146 (N_146,In_2566,In_2415);
and U147 (N_147,In_1228,In_2420);
or U148 (N_148,In_1440,In_1419);
and U149 (N_149,In_965,In_2517);
and U150 (N_150,In_1058,In_750);
xnor U151 (N_151,In_1200,In_644);
or U152 (N_152,In_1224,In_2215);
or U153 (N_153,In_1389,In_366);
nand U154 (N_154,In_603,In_1854);
nor U155 (N_155,In_414,In_1617);
and U156 (N_156,In_2878,In_1671);
and U157 (N_157,In_811,In_1098);
nor U158 (N_158,In_1136,In_2896);
or U159 (N_159,In_858,In_2486);
nor U160 (N_160,In_2851,In_570);
and U161 (N_161,In_2718,In_1057);
xnor U162 (N_162,In_996,In_1907);
nand U163 (N_163,In_2735,In_46);
xor U164 (N_164,In_1870,In_95);
xnor U165 (N_165,In_1470,In_1106);
nor U166 (N_166,In_2689,In_1085);
xor U167 (N_167,In_2011,In_2218);
or U168 (N_168,In_61,In_2498);
nor U169 (N_169,In_3,In_580);
or U170 (N_170,In_753,In_1488);
and U171 (N_171,In_152,In_2329);
nand U172 (N_172,In_1078,In_2172);
xor U173 (N_173,In_2173,In_2873);
nor U174 (N_174,In_2209,In_237);
or U175 (N_175,In_2626,In_2705);
nand U176 (N_176,In_28,In_1120);
xnor U177 (N_177,In_2716,In_1128);
nand U178 (N_178,In_1365,In_1542);
nand U179 (N_179,In_1545,In_1343);
nor U180 (N_180,In_2630,In_1454);
xor U181 (N_181,In_2156,In_522);
xnor U182 (N_182,In_877,In_1223);
and U183 (N_183,In_1665,In_1066);
nand U184 (N_184,In_393,In_1326);
nand U185 (N_185,In_2169,In_1577);
and U186 (N_186,In_2356,In_1529);
or U187 (N_187,In_48,In_325);
xnor U188 (N_188,In_1707,In_2743);
xor U189 (N_189,In_1039,In_1047);
and U190 (N_190,In_1427,In_1972);
and U191 (N_191,In_2961,In_2463);
nand U192 (N_192,In_118,In_2755);
nand U193 (N_193,In_1197,In_1563);
xor U194 (N_194,In_2469,In_2124);
nor U195 (N_195,In_204,In_1451);
and U196 (N_196,In_577,In_1891);
nand U197 (N_197,In_975,In_2609);
nor U198 (N_198,In_1026,In_2531);
nor U199 (N_199,In_2354,In_1407);
and U200 (N_200,In_1358,In_2478);
xor U201 (N_201,In_1511,In_1631);
and U202 (N_202,In_1618,In_934);
and U203 (N_203,In_192,In_2272);
xnor U204 (N_204,In_2651,In_1794);
nand U205 (N_205,In_2698,In_1649);
or U206 (N_206,In_948,In_410);
xor U207 (N_207,In_544,In_2158);
xor U208 (N_208,In_2181,In_333);
or U209 (N_209,In_831,In_1115);
xor U210 (N_210,In_1095,In_1482);
or U211 (N_211,In_516,In_2946);
nand U212 (N_212,In_210,In_383);
xor U213 (N_213,In_1417,In_1119);
or U214 (N_214,In_1581,In_1230);
nand U215 (N_215,In_2142,In_2678);
nand U216 (N_216,In_622,In_2213);
and U217 (N_217,In_1472,In_1812);
xor U218 (N_218,In_2319,In_1040);
xor U219 (N_219,In_115,In_1718);
nand U220 (N_220,In_840,In_313);
and U221 (N_221,In_384,In_2617);
xor U222 (N_222,In_268,In_1920);
xor U223 (N_223,In_65,In_1356);
xnor U224 (N_224,In_1246,In_1443);
xnor U225 (N_225,In_38,In_910);
nor U226 (N_226,In_2565,In_1297);
or U227 (N_227,In_2395,In_312);
or U228 (N_228,In_1191,In_1955);
nand U229 (N_229,In_1533,In_1320);
xor U230 (N_230,In_2008,In_2840);
xor U231 (N_231,In_485,In_1976);
nor U232 (N_232,In_2247,In_1853);
xnor U233 (N_233,In_1744,In_2133);
and U234 (N_234,In_1562,In_1998);
nand U235 (N_235,In_1636,In_1828);
xor U236 (N_236,In_1585,In_2545);
xnor U237 (N_237,In_2553,In_2362);
or U238 (N_238,In_1683,In_2862);
and U239 (N_239,In_1432,In_225);
or U240 (N_240,In_2501,In_1232);
xor U241 (N_241,In_2110,In_1656);
xor U242 (N_242,In_2310,In_664);
and U243 (N_243,In_2514,In_2050);
and U244 (N_244,In_2692,In_2452);
xnor U245 (N_245,In_2370,In_2227);
or U246 (N_246,In_481,In_1989);
xor U247 (N_247,In_1271,In_981);
and U248 (N_248,In_2871,In_2037);
xor U249 (N_249,In_2804,In_259);
xor U250 (N_250,In_2645,In_792);
nand U251 (N_251,In_549,In_678);
and U252 (N_252,In_1006,In_2959);
nand U253 (N_253,In_776,In_154);
xnor U254 (N_254,In_2530,In_2496);
nand U255 (N_255,In_643,In_258);
nor U256 (N_256,In_1926,In_955);
or U257 (N_257,In_1159,In_1105);
and U258 (N_258,In_937,In_477);
nor U259 (N_259,In_2265,In_260);
nand U260 (N_260,In_1555,In_762);
and U261 (N_261,In_2967,In_10);
nand U262 (N_262,In_489,In_814);
nor U263 (N_263,In_1143,In_1035);
xnor U264 (N_264,In_1862,In_2647);
xnor U265 (N_265,In_1806,In_1014);
or U266 (N_266,In_2648,In_625);
nand U267 (N_267,In_2637,In_760);
xor U268 (N_268,In_1044,In_68);
or U269 (N_269,In_2095,In_2891);
nand U270 (N_270,In_513,In_2600);
and U271 (N_271,In_129,In_466);
nand U272 (N_272,In_183,In_1902);
and U273 (N_273,In_362,In_1022);
xnor U274 (N_274,In_1530,In_452);
and U275 (N_275,In_2057,In_1314);
and U276 (N_276,In_2586,In_1993);
or U277 (N_277,In_2859,In_1783);
and U278 (N_278,In_532,In_2317);
and U279 (N_279,In_386,In_1940);
nor U280 (N_280,In_709,In_677);
and U281 (N_281,In_2453,In_2405);
nor U282 (N_282,In_1123,In_1772);
nand U283 (N_283,In_347,In_1834);
and U284 (N_284,In_2071,In_926);
and U285 (N_285,In_2760,In_1375);
nand U286 (N_286,In_747,In_661);
xnor U287 (N_287,In_1559,In_2243);
nor U288 (N_288,In_11,In_1730);
nand U289 (N_289,In_943,In_2673);
xnor U290 (N_290,In_1207,In_2253);
nand U291 (N_291,In_1626,In_1256);
or U292 (N_292,In_2099,In_1415);
xor U293 (N_293,In_1033,In_465);
nor U294 (N_294,In_1650,In_1027);
xor U295 (N_295,In_2536,In_888);
or U296 (N_296,In_1948,In_2803);
and U297 (N_297,In_2925,In_392);
nor U298 (N_298,In_582,In_2033);
nand U299 (N_299,In_1724,In_927);
nor U300 (N_300,In_2606,In_2677);
nor U301 (N_301,In_598,In_388);
nor U302 (N_302,In_1606,In_508);
xnor U303 (N_303,In_1011,In_1234);
nand U304 (N_304,In_1259,In_2249);
nor U305 (N_305,In_1385,In_723);
and U306 (N_306,In_2311,In_2965);
or U307 (N_307,In_2359,In_2557);
nand U308 (N_308,In_2784,In_576);
xor U309 (N_309,In_275,In_2098);
and U310 (N_310,In_395,In_1053);
nand U311 (N_311,In_809,In_416);
xnor U312 (N_312,In_1168,In_2307);
xnor U313 (N_313,In_1056,In_1849);
or U314 (N_314,In_315,In_2141);
or U315 (N_315,In_2721,In_1588);
nor U316 (N_316,In_2038,In_1333);
xnor U317 (N_317,In_665,In_705);
nand U318 (N_318,In_1146,In_1913);
xor U319 (N_319,In_419,In_1457);
or U320 (N_320,In_1564,In_806);
nand U321 (N_321,In_1567,In_2685);
and U322 (N_322,In_2238,In_1911);
nor U323 (N_323,In_2022,In_239);
nor U324 (N_324,In_317,In_2049);
xor U325 (N_325,In_1416,In_1941);
and U326 (N_326,In_2591,In_369);
and U327 (N_327,In_1553,In_1388);
nor U328 (N_328,In_2457,In_864);
or U329 (N_329,In_2444,In_794);
or U330 (N_330,In_179,In_2199);
nand U331 (N_331,In_2849,In_2219);
nand U332 (N_332,In_1348,In_2954);
nand U333 (N_333,In_124,In_1857);
or U334 (N_334,In_2225,In_810);
or U335 (N_335,In_2160,In_751);
nor U336 (N_336,In_8,In_517);
or U337 (N_337,In_1722,In_647);
and U338 (N_338,In_1565,In_1206);
nor U339 (N_339,In_344,In_2295);
or U340 (N_340,In_866,In_1490);
or U341 (N_341,In_880,In_1103);
and U342 (N_342,In_2687,In_2561);
xor U343 (N_343,In_2019,In_1927);
nor U344 (N_344,In_2384,In_2910);
or U345 (N_345,In_2534,In_509);
or U346 (N_346,In_2492,In_980);
or U347 (N_347,In_1436,In_1113);
nand U348 (N_348,In_307,In_121);
or U349 (N_349,In_1438,In_498);
nand U350 (N_350,In_2462,In_2250);
xor U351 (N_351,In_1134,In_1046);
xnor U352 (N_352,In_1426,In_2773);
xnor U353 (N_353,In_2917,In_524);
nand U354 (N_354,In_900,In_266);
xnor U355 (N_355,In_683,In_2476);
xnor U356 (N_356,In_372,In_430);
nor U357 (N_357,In_2290,In_1695);
xor U358 (N_358,In_1904,In_827);
nor U359 (N_359,In_2596,In_1322);
nor U360 (N_360,In_1652,In_759);
or U361 (N_361,In_1126,In_656);
nor U362 (N_362,In_1226,In_2056);
or U363 (N_363,In_618,In_518);
nand U364 (N_364,In_155,In_2633);
or U365 (N_365,In_1944,In_1213);
nand U366 (N_366,In_1752,In_2450);
xor U367 (N_367,In_2555,In_2436);
and U368 (N_368,In_1604,In_931);
xnor U369 (N_369,In_133,In_1028);
or U370 (N_370,In_2720,In_2643);
nand U371 (N_371,In_106,In_2489);
xnor U372 (N_372,In_726,In_1122);
and U373 (N_373,In_1963,In_1306);
nand U374 (N_374,In_2695,In_613);
nor U375 (N_375,In_2666,In_1075);
nand U376 (N_376,In_194,In_2652);
nand U377 (N_377,In_878,In_562);
nand U378 (N_378,In_712,In_36);
nor U379 (N_379,In_1117,In_904);
xor U380 (N_380,In_280,In_796);
or U381 (N_381,In_703,In_314);
nor U382 (N_382,In_2715,In_2978);
nor U383 (N_383,In_1463,In_1681);
nand U384 (N_384,In_2481,In_876);
xnor U385 (N_385,In_990,In_752);
nand U386 (N_386,In_1858,In_2207);
and U387 (N_387,In_1952,In_2150);
or U388 (N_388,In_1264,In_2106);
xnor U389 (N_389,In_2183,In_708);
nor U390 (N_390,In_2401,In_2245);
nor U391 (N_391,In_464,In_533);
or U392 (N_392,In_2582,In_1089);
nand U393 (N_393,In_2200,In_2654);
and U394 (N_394,In_1754,In_2771);
nor U395 (N_395,In_790,In_165);
nor U396 (N_396,In_2263,In_2527);
nor U397 (N_397,In_1778,In_345);
or U398 (N_398,In_355,In_161);
nor U399 (N_399,In_1151,In_2781);
xor U400 (N_400,In_1192,In_2400);
nand U401 (N_401,In_1600,In_2830);
and U402 (N_402,In_1787,In_2653);
nor U403 (N_403,In_1593,In_2740);
nand U404 (N_404,In_1815,In_1517);
xnor U405 (N_405,In_156,In_185);
or U406 (N_406,In_1843,In_1186);
xnor U407 (N_407,In_1428,In_556);
or U408 (N_408,In_1127,In_915);
and U409 (N_409,In_1402,In_1576);
or U410 (N_410,In_2936,In_350);
and U411 (N_411,In_81,In_1635);
nand U412 (N_412,In_1265,In_1634);
nor U413 (N_413,In_403,In_1648);
and U414 (N_414,In_729,In_221);
xnor U415 (N_415,In_2460,In_1531);
or U416 (N_416,In_2338,In_54);
xnor U417 (N_417,In_1483,In_1357);
xor U418 (N_418,In_1194,In_2375);
or U419 (N_419,In_368,In_2065);
nor U420 (N_420,In_2167,In_2728);
and U421 (N_421,In_1327,In_1270);
or U422 (N_422,In_2030,In_922);
nand U423 (N_423,In_574,In_1654);
nand U424 (N_424,In_894,In_612);
nand U425 (N_425,In_2552,In_160);
xnor U426 (N_426,In_832,In_1740);
and U427 (N_427,In_35,In_2937);
or U428 (N_428,In_2389,In_303);
and U429 (N_429,In_2177,In_2897);
nor U430 (N_430,In_2597,In_1799);
nand U431 (N_431,In_2935,In_1540);
nand U432 (N_432,In_1874,In_671);
xnor U433 (N_433,In_2915,In_589);
and U434 (N_434,In_164,In_2355);
xnor U435 (N_435,In_1811,In_2845);
or U436 (N_436,In_1885,In_1269);
nand U437 (N_437,In_535,In_1062);
nor U438 (N_438,In_887,In_125);
nand U439 (N_439,In_2846,In_173);
nor U440 (N_440,In_911,In_284);
nand U441 (N_441,In_407,In_2117);
or U442 (N_442,In_2942,In_1467);
nor U443 (N_443,In_413,In_718);
or U444 (N_444,In_893,In_1733);
or U445 (N_445,In_130,In_2900);
nand U446 (N_446,In_2590,In_408);
or U447 (N_447,In_1214,In_1294);
or U448 (N_448,In_2467,In_2161);
xor U449 (N_449,In_370,In_1693);
and U450 (N_450,In_2691,In_2703);
nand U451 (N_451,In_1278,In_2679);
nor U452 (N_452,In_2285,In_2475);
or U453 (N_453,In_1059,In_1945);
and U454 (N_454,In_1099,In_783);
nor U455 (N_455,In_917,In_2468);
nand U456 (N_456,In_1586,In_434);
or U457 (N_457,In_956,In_1009);
or U458 (N_458,In_555,In_1019);
and U459 (N_459,In_2837,In_1906);
xor U460 (N_460,In_1431,In_1311);
and U461 (N_461,In_2053,In_1295);
or U462 (N_462,In_2217,In_2506);
and U463 (N_463,In_1331,In_995);
and U464 (N_464,In_1759,In_1720);
xor U465 (N_465,In_2175,In_1421);
and U466 (N_466,In_1336,In_2870);
or U467 (N_467,In_2335,In_588);
xor U468 (N_468,In_1994,In_1444);
or U469 (N_469,In_2458,In_2854);
nor U470 (N_470,In_431,In_2443);
and U471 (N_471,In_1082,In_285);
nand U472 (N_472,In_2086,In_436);
nand U473 (N_473,In_1717,In_2690);
xnor U474 (N_474,In_2903,In_741);
and U475 (N_475,In_1167,In_1144);
xnor U476 (N_476,In_1305,In_2541);
nor U477 (N_477,In_1745,In_1709);
and U478 (N_478,In_1282,In_2916);
and U479 (N_479,In_2731,In_2283);
or U480 (N_480,In_1174,In_2918);
and U481 (N_481,In_1371,In_916);
and U482 (N_482,In_704,In_178);
nor U483 (N_483,In_1360,In_2801);
nand U484 (N_484,In_1814,In_2995);
or U485 (N_485,In_2390,In_144);
and U486 (N_486,In_375,In_2931);
xnor U487 (N_487,In_1532,In_1074);
xor U488 (N_488,In_571,In_1953);
nor U489 (N_489,In_2301,In_2602);
and U490 (N_490,In_2210,In_1163);
or U491 (N_491,In_320,In_1466);
and U492 (N_492,In_2477,In_2683);
nand U493 (N_493,In_813,In_72);
or U494 (N_494,In_1446,In_585);
xnor U495 (N_495,In_1183,In_824);
xor U496 (N_496,In_1198,In_621);
xor U497 (N_497,In_480,In_30);
nor U498 (N_498,In_2834,In_361);
or U499 (N_499,In_2576,In_208);
nand U500 (N_500,In_2408,In_1569);
xnor U501 (N_501,N_96,In_2257);
xnor U502 (N_502,In_492,In_2391);
nand U503 (N_503,In_834,In_205);
nor U504 (N_504,In_2581,In_529);
nand U505 (N_505,In_2662,In_1797);
xnor U506 (N_506,In_1393,In_1121);
or U507 (N_507,In_235,In_2363);
nand U508 (N_508,In_2879,In_1179);
or U509 (N_509,In_2208,N_419);
xor U510 (N_510,In_1155,In_1296);
or U511 (N_511,N_318,In_462);
xnor U512 (N_512,In_1869,In_1129);
xnor U513 (N_513,N_415,In_2093);
and U514 (N_514,In_2520,In_1928);
xnor U515 (N_515,In_1052,In_2733);
nand U516 (N_516,In_711,In_958);
nor U517 (N_517,In_1729,N_488);
nand U518 (N_518,In_202,In_2958);
xnor U519 (N_519,In_675,In_487);
nor U520 (N_520,In_2884,In_1049);
nand U521 (N_521,In_1300,In_499);
nand U522 (N_522,In_1662,In_2021);
and U523 (N_523,In_2237,N_130);
and U524 (N_524,In_1932,In_1882);
and U525 (N_525,In_1646,In_2969);
nand U526 (N_526,In_2638,In_1971);
or U527 (N_527,In_1108,In_1915);
xnor U528 (N_528,N_253,In_793);
nor U529 (N_529,In_2853,In_2799);
nand U530 (N_530,In_112,In_1292);
xnor U531 (N_531,N_86,In_881);
nand U532 (N_532,In_1789,In_918);
or U533 (N_533,In_2075,In_1851);
xnor U534 (N_534,In_1279,In_2454);
or U535 (N_535,N_370,In_2122);
or U536 (N_536,N_67,N_424);
or U537 (N_537,In_214,In_1788);
nand U538 (N_538,In_494,N_341);
nand U539 (N_539,N_377,In_1411);
nor U540 (N_540,N_211,In_2914);
and U541 (N_541,N_244,In_1760);
xor U542 (N_542,N_396,In_1900);
nor U543 (N_543,In_1225,In_1676);
or U544 (N_544,In_136,In_293);
nor U545 (N_545,N_179,In_382);
nor U546 (N_546,In_2861,In_2328);
and U547 (N_547,In_2426,In_1308);
nor U548 (N_548,In_1366,In_377);
nor U549 (N_549,In_2791,In_1977);
or U550 (N_550,N_361,In_2313);
or U551 (N_551,In_2863,In_1023);
or U552 (N_552,In_1574,N_152);
nand U553 (N_553,In_2431,In_2171);
and U554 (N_554,In_1275,In_1793);
nor U555 (N_555,N_343,In_2105);
nand U556 (N_556,N_277,In_1491);
xor U557 (N_557,In_2852,In_964);
xnor U558 (N_558,In_2059,In_406);
and U559 (N_559,In_1475,N_441);
or U560 (N_560,In_2430,In_199);
and U561 (N_561,In_969,N_371);
nor U562 (N_562,In_2298,In_680);
and U563 (N_563,In_2076,In_983);
nor U564 (N_564,In_863,In_1354);
and U565 (N_565,In_766,N_26);
nor U566 (N_566,In_1832,In_113);
or U567 (N_567,In_2660,In_2944);
xnor U568 (N_568,In_619,N_428);
or U569 (N_569,In_1689,In_1017);
or U570 (N_570,In_218,In_727);
nor U571 (N_571,In_2204,In_1969);
and U572 (N_572,In_1494,N_283);
and U573 (N_573,N_352,N_224);
nand U574 (N_574,N_254,In_2174);
nor U575 (N_575,In_637,N_76);
and U576 (N_576,In_469,In_2291);
xor U577 (N_577,In_2722,N_367);
xnor U578 (N_578,In_1496,In_1782);
or U579 (N_579,N_258,In_254);
nand U580 (N_580,In_2667,In_2233);
nand U581 (N_581,In_255,In_2);
and U582 (N_582,In_567,In_868);
xor U583 (N_583,In_1551,In_2403);
nand U584 (N_584,In_99,In_402);
or U585 (N_585,In_497,In_2472);
nand U586 (N_586,In_2860,In_1196);
nand U587 (N_587,In_1677,In_2196);
and U588 (N_588,In_1007,In_1464);
nor U589 (N_589,In_2924,N_479);
nor U590 (N_590,In_1087,In_2762);
nand U591 (N_591,In_2085,In_2482);
and U592 (N_592,N_5,In_558);
or U593 (N_593,In_2713,In_2342);
nor U594 (N_594,In_1838,N_84);
or U595 (N_595,N_338,In_635);
or U596 (N_596,N_413,In_332);
xor U597 (N_597,In_2628,In_2361);
nor U598 (N_598,In_2264,In_2881);
and U599 (N_599,N_498,In_802);
nor U600 (N_600,In_2132,In_1158);
or U601 (N_601,In_2658,In_2675);
xor U602 (N_602,In_1453,N_450);
xnor U603 (N_603,In_2064,In_1764);
and U604 (N_604,In_659,In_2166);
nand U605 (N_605,In_546,In_86);
and U606 (N_606,N_237,In_2424);
or U607 (N_607,In_691,In_2907);
nand U608 (N_608,In_443,In_1755);
or U609 (N_609,In_2278,N_390);
xor U610 (N_610,In_799,In_2814);
xnor U611 (N_611,N_112,N_51);
and U612 (N_612,In_2991,In_447);
or U613 (N_613,In_1204,In_1883);
nor U614 (N_614,N_382,In_123);
xnor U615 (N_615,In_2823,In_687);
and U616 (N_616,In_569,In_2894);
and U617 (N_617,In_429,In_1008);
and U618 (N_618,In_1522,N_374);
and U619 (N_619,N_83,In_2069);
xor U620 (N_620,In_2396,In_216);
nor U621 (N_621,In_2276,N_398);
or U622 (N_622,In_2560,In_2140);
and U623 (N_623,In_1268,In_1868);
or U624 (N_624,In_859,In_1425);
or U625 (N_625,In_2544,In_2047);
or U626 (N_626,In_1154,N_39);
nor U627 (N_627,In_882,In_2757);
nand U628 (N_628,In_2657,In_352);
and U629 (N_629,In_1791,In_1312);
or U630 (N_630,In_2759,In_1382);
nor U631 (N_631,In_495,In_553);
xnor U632 (N_632,In_2101,In_816);
and U633 (N_633,In_2102,In_1227);
nor U634 (N_634,In_340,In_270);
and U635 (N_635,In_1934,In_2776);
and U636 (N_636,In_1499,In_1548);
xnor U637 (N_637,N_80,In_2919);
nor U638 (N_638,N_150,In_2672);
or U639 (N_639,N_329,In_2805);
xor U640 (N_640,In_758,In_2625);
nand U641 (N_641,N_326,In_309);
xor U642 (N_642,In_559,In_1679);
nor U643 (N_643,N_140,In_1471);
or U644 (N_644,In_2303,In_706);
nor U645 (N_645,In_2525,In_2577);
or U646 (N_646,In_1524,N_136);
or U647 (N_647,In_2964,In_669);
nand U648 (N_648,N_105,In_1439);
nor U649 (N_649,N_165,N_68);
or U650 (N_650,N_121,In_1539);
or U651 (N_651,In_1386,N_28);
xor U652 (N_652,In_923,In_1469);
nor U653 (N_653,N_119,In_2039);
nand U654 (N_654,In_252,In_1430);
xor U655 (N_655,In_668,In_2951);
and U656 (N_656,In_1578,N_134);
and U657 (N_657,In_1373,In_1030);
or U658 (N_658,In_2018,N_135);
xnor U659 (N_659,In_433,N_109);
xnor U660 (N_660,In_2905,In_1217);
or U661 (N_661,N_3,In_2214);
nand U662 (N_662,In_527,N_132);
xor U663 (N_663,N_303,In_914);
and U664 (N_664,N_108,In_92);
nand U665 (N_665,In_2876,N_193);
nand U666 (N_666,N_418,In_2084);
nand U667 (N_667,N_161,In_2774);
nor U668 (N_668,In_1041,In_426);
or U669 (N_669,In_1002,In_1073);
nand U670 (N_670,In_699,N_291);
nand U671 (N_671,In_380,In_1525);
xor U672 (N_672,N_154,In_1871);
and U673 (N_673,In_2442,In_1383);
and U674 (N_674,In_2558,In_343);
xnor U675 (N_675,In_1964,In_2466);
or U676 (N_676,In_455,In_265);
nand U677 (N_677,In_2277,N_218);
or U678 (N_678,In_1543,In_1484);
and U679 (N_679,In_2511,N_70);
xor U680 (N_680,N_93,In_944);
nand U681 (N_681,In_186,In_2532);
nand U682 (N_682,N_483,In_57);
nand U683 (N_683,In_789,N_63);
nor U684 (N_684,In_1997,In_2548);
and U685 (N_685,In_685,In_2701);
xor U686 (N_686,In_599,N_23);
xor U687 (N_687,In_2441,In_1450);
xnor U688 (N_688,In_2686,In_418);
nor U689 (N_689,In_334,In_2727);
and U690 (N_690,N_156,N_113);
and U691 (N_691,N_142,N_71);
nor U692 (N_692,In_14,N_485);
nor U693 (N_693,In_2843,In_2598);
nor U694 (N_694,N_310,In_1826);
and U695 (N_695,N_223,N_217);
and U696 (N_696,N_118,In_19);
nor U697 (N_697,In_605,In_1086);
nor U698 (N_698,In_674,In_775);
and U699 (N_699,In_2729,In_2254);
nand U700 (N_700,In_2821,In_506);
nand U701 (N_701,In_2202,In_1114);
and U702 (N_702,In_2226,In_69);
xor U703 (N_703,In_1512,In_1894);
nor U704 (N_704,N_280,In_1088);
and U705 (N_705,In_2640,In_2943);
or U706 (N_706,In_1624,In_2524);
nor U707 (N_707,In_733,In_2320);
or U708 (N_708,In_1573,In_829);
and U709 (N_709,In_1979,In_1509);
and U710 (N_710,In_2220,In_283);
and U711 (N_711,In_304,In_2710);
xnor U712 (N_712,In_2811,In_1060);
xnor U713 (N_713,In_1153,In_1036);
and U714 (N_714,In_1097,In_563);
or U715 (N_715,In_104,N_321);
xnor U716 (N_716,In_1261,In_1714);
or U717 (N_717,In_1623,In_1424);
and U718 (N_718,In_769,In_2184);
or U719 (N_719,In_1486,In_2933);
nand U720 (N_720,In_2130,In_1757);
nor U721 (N_721,In_2461,In_1021);
nand U722 (N_722,In_310,N_473);
xor U723 (N_723,N_103,In_1739);
nand U724 (N_724,In_2820,In_60);
nand U725 (N_725,N_308,In_41);
xor U726 (N_726,In_319,In_2574);
nand U727 (N_727,In_2000,In_862);
nand U728 (N_728,In_70,N_376);
nand U729 (N_729,In_169,In_346);
and U730 (N_730,In_761,In_137);
nand U731 (N_731,In_2131,N_19);
or U732 (N_732,In_2299,In_1005);
and U733 (N_733,In_682,In_1107);
and U734 (N_734,In_222,N_477);
or U735 (N_735,In_2950,In_1165);
xor U736 (N_736,In_1594,In_1687);
nor U737 (N_737,In_2016,In_116);
nor U738 (N_738,In_1209,N_474);
nand U739 (N_739,In_2636,In_998);
and U740 (N_740,N_171,In_1391);
nor U741 (N_741,In_2244,In_1462);
xnor U742 (N_742,In_1175,In_2982);
nor U743 (N_743,N_233,N_368);
or U744 (N_744,N_127,N_385);
and U745 (N_745,In_1786,In_2198);
and U746 (N_746,In_468,N_74);
xnor U747 (N_747,In_1575,In_2732);
nor U748 (N_748,N_206,N_366);
or U749 (N_749,N_469,In_496);
or U750 (N_750,In_291,In_1910);
or U751 (N_751,In_2835,In_2564);
and U752 (N_752,In_1672,N_316);
nor U753 (N_753,In_1780,N_190);
nand U754 (N_754,In_1912,N_73);
or U755 (N_755,In_415,N_276);
nand U756 (N_756,In_913,In_2480);
nand U757 (N_757,In_1773,In_749);
nor U758 (N_758,In_82,In_1302);
and U759 (N_759,In_1369,In_826);
xor U760 (N_760,In_2537,N_222);
xnor U761 (N_761,N_467,N_345);
nand U762 (N_762,In_425,In_405);
nor U763 (N_763,In_213,In_2904);
nand U764 (N_764,In_597,N_102);
nor U765 (N_765,In_548,In_229);
xnor U766 (N_766,In_2205,In_2144);
xnor U767 (N_767,N_402,N_461);
or U768 (N_768,In_2126,In_1301);
or U769 (N_769,In_1956,In_1905);
or U770 (N_770,N_281,In_2089);
and U771 (N_771,In_1630,In_24);
nor U772 (N_772,In_2471,In_1688);
nand U773 (N_773,In_2563,In_2372);
and U774 (N_774,In_857,N_304);
xnor U775 (N_775,In_2223,N_476);
and U776 (N_776,In_1267,In_2939);
nand U777 (N_777,In_2885,In_1602);
or U778 (N_778,In_353,In_1231);
or U779 (N_779,N_430,In_2072);
and U780 (N_780,In_666,In_422);
and U781 (N_781,In_2824,N_234);
xor U782 (N_782,In_184,N_245);
nor U783 (N_783,In_44,In_32);
or U784 (N_784,In_1061,In_1592);
nand U785 (N_785,In_227,In_451);
xor U786 (N_786,In_2787,In_2984);
nor U787 (N_787,In_177,In_2688);
and U788 (N_788,N_275,N_208);
nand U789 (N_789,In_724,N_69);
xnor U790 (N_790,In_1506,In_1768);
or U791 (N_791,N_261,In_122);
nor U792 (N_792,In_1981,N_54);
and U793 (N_793,In_40,In_1970);
nor U794 (N_794,In_2521,N_182);
nand U795 (N_795,In_1653,In_690);
nor U796 (N_796,In_404,In_49);
and U797 (N_797,In_63,In_631);
or U798 (N_798,In_1070,In_1182);
xnor U799 (N_799,N_494,In_138);
nand U800 (N_800,In_1229,In_274);
and U801 (N_801,In_2451,In_201);
nor U802 (N_802,In_1315,In_626);
or U803 (N_803,In_1603,N_314);
nand U804 (N_804,N_181,N_356);
nor U805 (N_805,In_1749,N_496);
nand U806 (N_806,N_481,In_1520);
or U807 (N_807,N_339,In_2780);
or U808 (N_808,In_1903,In_1319);
nand U809 (N_809,In_212,In_745);
and U810 (N_810,In_772,N_263);
and U811 (N_811,In_1244,In_2922);
or U812 (N_812,In_636,In_2819);
or U813 (N_813,N_454,In_0);
nand U814 (N_814,In_174,In_1212);
xnor U815 (N_815,N_236,In_1621);
nor U816 (N_816,In_979,In_2055);
nand U817 (N_817,In_2393,In_662);
nand U818 (N_818,N_348,In_1093);
nand U819 (N_819,N_123,In_2402);
xnor U820 (N_820,N_330,N_383);
nor U821 (N_821,In_1899,In_2956);
and U822 (N_822,N_267,N_492);
xnor U823 (N_823,In_2014,In_1613);
or U824 (N_824,In_2807,N_111);
nand U825 (N_825,In_2448,In_1674);
and U826 (N_826,In_1664,In_74);
and U827 (N_827,In_1657,In_1954);
or U828 (N_828,In_861,In_2815);
nand U829 (N_829,N_420,In_2779);
and U830 (N_830,In_541,In_2092);
xnor U831 (N_831,In_867,In_2336);
nor U832 (N_832,In_2670,In_731);
nand U833 (N_833,N_447,In_1552);
and U834 (N_834,N_448,In_300);
xor U835 (N_835,In_837,In_1827);
or U836 (N_836,N_357,In_238);
nand U837 (N_837,In_1112,In_1243);
or U838 (N_838,In_1190,N_168);
xnor U839 (N_839,In_294,In_2696);
xnor U840 (N_840,In_1329,In_1071);
or U841 (N_841,In_2966,In_267);
xnor U842 (N_842,In_1678,In_2483);
nand U843 (N_843,In_271,In_2410);
xor U844 (N_844,In_42,In_1497);
and U845 (N_845,In_1951,In_34);
nor U846 (N_846,In_226,In_1751);
nor U847 (N_847,In_2145,In_2043);
xnor U848 (N_848,In_2813,In_504);
nand U849 (N_849,In_2083,In_568);
or U850 (N_850,In_1923,N_124);
and U851 (N_851,In_399,In_648);
and U852 (N_852,In_2087,In_2875);
or U853 (N_853,In_2485,In_1042);
or U854 (N_854,In_611,In_530);
or U855 (N_855,N_452,In_1697);
nor U856 (N_856,N_472,In_1561);
nor U857 (N_857,In_2826,In_2674);
xnor U858 (N_858,In_1974,In_2605);
nor U859 (N_859,In_1537,In_1986);
xor U860 (N_860,In_2082,In_1184);
nand U861 (N_861,In_18,In_627);
or U862 (N_862,In_891,In_1325);
and U863 (N_863,In_1682,In_2322);
or U864 (N_864,In_263,In_2383);
xor U865 (N_865,N_101,In_2398);
nor U866 (N_866,In_819,N_31);
xnor U867 (N_867,In_545,In_337);
xnor U868 (N_868,In_2035,In_999);
nand U869 (N_869,In_2549,In_732);
or U870 (N_870,N_300,N_151);
nand U871 (N_871,In_1850,N_359);
nor U872 (N_872,In_2259,In_1959);
nand U873 (N_873,In_2306,In_2724);
nand U874 (N_874,In_1094,In_207);
or U875 (N_875,N_213,N_317);
or U876 (N_876,In_1807,In_311);
or U877 (N_877,N_381,N_372);
and U878 (N_878,In_938,In_2957);
xnor U879 (N_879,In_2314,In_148);
nand U880 (N_880,In_1668,In_1221);
or U881 (N_881,In_1924,In_502);
or U882 (N_882,In_1422,In_2888);
and U883 (N_883,In_119,In_281);
or U884 (N_884,In_264,In_2154);
xor U885 (N_885,In_1732,In_2332);
xor U886 (N_886,In_808,N_365);
xnor U887 (N_887,N_342,In_505);
and U888 (N_888,In_1298,In_1334);
nor U889 (N_889,N_174,In_2497);
nor U890 (N_890,In_1473,In_2449);
or U891 (N_891,In_335,In_211);
nand U892 (N_892,In_1538,In_2274);
and U893 (N_893,In_1157,In_543);
nor U894 (N_894,In_801,N_439);
nor U895 (N_895,In_269,In_1829);
or U896 (N_896,In_1872,In_2293);
nand U897 (N_897,N_219,In_1091);
nor U898 (N_898,In_203,In_2134);
nand U899 (N_899,In_2455,In_2344);
or U900 (N_900,In_2758,In_1441);
and U901 (N_901,In_2027,In_1568);
nand U902 (N_902,N_42,In_1835);
nand U903 (N_903,N_97,In_1949);
and U904 (N_904,N_25,In_984);
nand U905 (N_905,In_1961,N_451);
or U906 (N_906,In_764,In_929);
or U907 (N_907,In_1544,In_592);
and U908 (N_908,In_84,N_455);
nor U909 (N_909,In_432,N_315);
xor U910 (N_910,In_55,In_394);
nor U911 (N_911,N_57,In_2542);
and U912 (N_912,In_1855,N_10);
xnor U913 (N_913,In_2304,In_1104);
xor U914 (N_914,N_212,In_162);
xnor U915 (N_915,In_1442,In_1795);
nor U916 (N_916,In_620,In_2366);
or U917 (N_917,In_358,In_617);
and U918 (N_918,In_1933,In_784);
nand U919 (N_919,N_416,In_2751);
xnor U920 (N_920,In_273,In_2112);
nand U921 (N_921,N_148,In_1598);
nand U922 (N_922,In_1353,N_169);
nor U923 (N_923,In_1601,In_1595);
xor U924 (N_924,In_755,In_2892);
nor U925 (N_925,N_394,In_1045);
nand U926 (N_926,N_395,In_873);
nand U927 (N_927,In_1670,In_2374);
nor U928 (N_928,In_2316,In_1685);
xnor U929 (N_929,In_886,N_296);
xnor U930 (N_930,In_2487,N_497);
and U931 (N_931,In_172,In_952);
and U932 (N_932,N_290,N_157);
nor U933 (N_933,In_1138,In_507);
nand U934 (N_934,In_1852,In_2746);
and U935 (N_935,In_181,In_2352);
nor U936 (N_936,N_248,N_72);
and U937 (N_937,In_2920,N_49);
nand U938 (N_938,In_1991,In_2842);
xnor U939 (N_939,In_2985,In_2938);
nor U940 (N_940,In_2503,In_126);
nor U941 (N_941,In_2040,N_292);
nor U942 (N_942,In_1187,In_2765);
xor U943 (N_943,N_243,In_2912);
nand U944 (N_944,In_1966,In_224);
or U945 (N_945,In_2392,In_2635);
or U946 (N_946,In_1943,In_330);
xnor U947 (N_947,In_2456,In_841);
and U948 (N_948,In_2376,In_1118);
or U949 (N_949,In_2170,In_1338);
or U950 (N_950,In_1215,In_196);
or U951 (N_951,In_905,In_2070);
or U952 (N_952,In_2649,In_848);
nor U953 (N_953,In_800,In_717);
and U954 (N_954,In_2015,In_2330);
or U955 (N_955,In_719,In_2203);
and U956 (N_956,In_1706,In_2783);
and U957 (N_957,N_273,In_1950);
or U958 (N_958,N_198,In_191);
and U959 (N_959,N_444,N_307);
nor U960 (N_960,In_898,In_1476);
or U961 (N_961,In_360,N_78);
and U962 (N_962,In_374,In_2655);
nand U963 (N_963,In_2066,In_695);
nand U964 (N_964,N_278,In_288);
or U965 (N_965,In_261,N_87);
and U966 (N_966,In_2054,N_33);
nor U967 (N_967,In_2646,In_2750);
nor U968 (N_968,N_458,N_4);
xor U969 (N_969,In_912,In_1796);
xnor U970 (N_970,In_2079,In_2836);
xnor U971 (N_971,In_1734,In_2024);
nor U972 (N_972,In_1705,In_2800);
nand U973 (N_973,In_573,N_302);
and U974 (N_974,In_1489,In_100);
nand U975 (N_975,In_1999,N_88);
xnor U976 (N_976,In_1990,In_767);
nor U977 (N_977,In_2435,N_220);
and U978 (N_978,In_2753,In_2440);
nand U979 (N_979,In_1738,In_609);
or U980 (N_980,In_1765,N_216);
and U981 (N_981,In_817,In_1813);
nor U982 (N_982,In_2269,In_2273);
nor U983 (N_983,In_2868,In_1072);
nor U984 (N_984,In_27,In_2343);
nand U985 (N_985,N_238,In_1083);
and U986 (N_986,In_778,In_1205);
nor U987 (N_987,In_2627,N_14);
and U988 (N_988,In_1461,In_2887);
nor U989 (N_989,In_12,N_489);
nor U990 (N_990,N_470,In_2371);
and U991 (N_991,In_1579,In_1898);
xnor U992 (N_992,In_1742,In_85);
nor U993 (N_993,In_2953,In_2971);
and U994 (N_994,In_1141,In_295);
and U995 (N_995,In_2952,In_428);
or U996 (N_996,In_2412,N_298);
xnor U997 (N_997,In_411,In_2947);
xnor U998 (N_998,In_2147,In_2186);
nor U999 (N_999,In_722,In_2556);
nor U1000 (N_1000,In_2305,N_965);
and U1001 (N_1001,N_948,In_2074);
xor U1002 (N_1002,In_1317,N_210);
nand U1003 (N_1003,In_1433,In_2754);
xor U1004 (N_1004,In_1762,In_1546);
or U1005 (N_1005,In_770,In_850);
nor U1006 (N_1006,In_2911,In_2165);
and U1007 (N_1007,N_883,In_409);
nand U1008 (N_1008,N_838,In_2663);
xor U1009 (N_1009,N_407,In_2123);
nor U1010 (N_1010,N_762,In_2386);
xor U1011 (N_1011,In_1694,In_29);
nand U1012 (N_1012,N_99,In_215);
nand U1013 (N_1013,N_346,In_246);
or U1014 (N_1014,In_908,In_795);
xor U1015 (N_1015,N_480,N_906);
or U1016 (N_1016,In_1629,In_1747);
xor U1017 (N_1017,In_282,In_2508);
xor U1018 (N_1018,In_786,In_2137);
and U1019 (N_1019,In_1237,N_594);
nor U1020 (N_1020,N_89,In_1335);
xor U1021 (N_1021,In_538,N_689);
nand U1022 (N_1022,In_1236,N_66);
nand U1023 (N_1023,N_691,In_714);
and U1024 (N_1024,In_1980,N_683);
nand U1025 (N_1025,In_96,In_2360);
nor U1026 (N_1026,In_2681,In_1401);
nand U1027 (N_1027,N_153,N_331);
nand U1028 (N_1028,In_2488,N_799);
nand U1029 (N_1029,N_631,In_47);
nor U1030 (N_1030,N_531,In_557);
and U1031 (N_1031,In_1242,In_364);
nor U1032 (N_1032,In_1445,In_855);
or U1033 (N_1033,In_697,In_805);
and U1034 (N_1034,In_2841,In_561);
or U1035 (N_1035,N_579,N_903);
nor U1036 (N_1036,In_2357,In_31);
xnor U1037 (N_1037,In_2604,In_77);
or U1038 (N_1038,N_533,In_1863);
or U1039 (N_1039,N_286,N_644);
and U1040 (N_1040,N_804,In_1779);
nand U1041 (N_1041,N_279,N_774);
nor U1042 (N_1042,N_710,In_245);
or U1043 (N_1043,In_629,In_2136);
and U1044 (N_1044,In_2368,In_540);
and U1045 (N_1045,In_4,In_1710);
or U1046 (N_1046,In_1995,In_1978);
nor U1047 (N_1047,N_612,N_274);
nor U1048 (N_1048,In_2934,N_646);
nand U1049 (N_1049,In_1808,In_798);
xor U1050 (N_1050,In_2752,In_1051);
xnor U1051 (N_1051,N_981,In_2709);
or U1052 (N_1052,N_556,N_403);
and U1053 (N_1053,In_2607,N_755);
nand U1054 (N_1054,In_306,N_94);
or U1055 (N_1055,In_1459,In_1591);
nand U1056 (N_1056,N_611,In_2507);
and U1057 (N_1057,In_159,N_602);
nand U1058 (N_1058,In_182,N_177);
nor U1059 (N_1059,N_733,In_93);
xor U1060 (N_1060,N_411,In_584);
and U1061 (N_1061,N_610,In_1096);
or U1062 (N_1062,In_2748,N_697);
and U1063 (N_1063,In_331,In_1172);
or U1064 (N_1064,N_748,N_564);
and U1065 (N_1065,In_397,In_1930);
nor U1066 (N_1066,In_39,In_519);
nand U1067 (N_1067,N_538,N_334);
or U1068 (N_1068,N_650,N_695);
or U1069 (N_1069,In_2833,N_881);
nor U1070 (N_1070,In_242,In_1048);
and U1071 (N_1071,In_2296,In_1518);
nand U1072 (N_1072,N_185,N_872);
nand U1073 (N_1073,N_878,In_1873);
or U1074 (N_1074,In_417,N_199);
and U1075 (N_1075,N_836,In_756);
xnor U1076 (N_1076,In_448,In_654);
or U1077 (N_1077,In_2067,In_1699);
or U1078 (N_1078,In_2906,N_162);
xor U1079 (N_1079,In_1888,In_2831);
and U1080 (N_1080,N_848,In_2230);
nor U1081 (N_1081,N_840,N_860);
nand U1082 (N_1082,In_1547,In_2997);
and U1083 (N_1083,In_299,In_1263);
or U1084 (N_1084,In_2890,In_2595);
or U1085 (N_1085,In_2493,In_2240);
or U1086 (N_1086,In_1818,In_2432);
xor U1087 (N_1087,In_2621,In_1245);
or U1088 (N_1088,N_551,In_233);
nor U1089 (N_1089,In_1504,In_1867);
xnor U1090 (N_1090,In_1638,In_2221);
xnor U1091 (N_1091,In_2406,N_160);
nor U1092 (N_1092,N_885,In_2194);
or U1093 (N_1093,N_241,In_2143);
nand U1094 (N_1094,In_601,N_77);
or U1095 (N_1095,N_431,N_994);
or U1096 (N_1096,In_167,N_684);
and U1097 (N_1097,In_435,N_48);
and U1098 (N_1098,N_499,In_1316);
nand U1099 (N_1099,N_761,N_355);
nor U1100 (N_1100,N_828,In_1281);
xnor U1101 (N_1101,N_350,In_959);
nor U1102 (N_1102,In_440,In_2080);
and U1103 (N_1103,N_328,In_539);
nand U1104 (N_1104,In_590,N_410);
or U1105 (N_1105,In_1080,In_2930);
nand U1106 (N_1106,In_1984,In_1272);
and U1107 (N_1107,In_986,In_2260);
nand U1108 (N_1108,In_962,In_91);
or U1109 (N_1109,N_621,N_145);
and U1110 (N_1110,In_1171,N_306);
nand U1111 (N_1111,N_522,In_2613);
and U1112 (N_1112,N_574,N_983);
and U1113 (N_1113,In_423,N_517);
nor U1114 (N_1114,N_905,In_1054);
or U1115 (N_1115,N_240,In_696);
xor U1116 (N_1116,In_1622,In_2998);
nand U1117 (N_1117,In_2188,N_325);
nor U1118 (N_1118,In_1342,N_806);
nor U1119 (N_1119,In_670,In_2333);
xnor U1120 (N_1120,In_1050,In_2572);
or U1121 (N_1121,In_748,N_546);
or U1122 (N_1122,N_221,N_147);
and U1123 (N_1123,N_271,N_841);
nor U1124 (N_1124,In_1639,In_2119);
nor U1125 (N_1125,In_2409,N_627);
and U1126 (N_1126,In_1235,In_175);
nand U1127 (N_1127,In_2421,In_1641);
nand U1128 (N_1128,N_849,In_920);
nor U1129 (N_1129,N_751,In_1519);
nand U1130 (N_1130,N_580,N_516);
or U1131 (N_1131,N_781,In_251);
and U1132 (N_1132,N_62,In_1092);
nand U1133 (N_1133,N_766,N_6);
and U1134 (N_1134,In_2325,In_1258);
nor U1135 (N_1135,N_809,N_715);
xor U1136 (N_1136,N_863,N_877);
xor U1137 (N_1137,In_1655,In_444);
xor U1138 (N_1138,In_1996,In_2775);
xor U1139 (N_1139,In_2981,In_454);
or U1140 (N_1140,In_108,In_2148);
nor U1141 (N_1141,N_754,In_2788);
xor U1142 (N_1142,In_351,N_652);
xnor U1143 (N_1143,N_951,In_804);
nor U1144 (N_1144,In_1528,N_788);
nand U1145 (N_1145,N_625,In_874);
xor U1146 (N_1146,In_2377,In_2003);
xor U1147 (N_1147,In_2880,In_257);
or U1148 (N_1148,N_597,N_719);
nor U1149 (N_1149,N_909,N_945);
and U1150 (N_1150,N_40,In_2972);
xor U1151 (N_1151,In_1809,In_2414);
xor U1152 (N_1152,In_1376,In_1111);
nor U1153 (N_1153,In_1031,In_1474);
nor U1154 (N_1154,N_197,N_837);
nand U1155 (N_1155,In_1859,N_18);
or U1156 (N_1156,In_1013,N_974);
and U1157 (N_1157,In_788,In_623);
nand U1158 (N_1158,N_15,In_2806);
xnor U1159 (N_1159,In_1239,In_2578);
nor U1160 (N_1160,In_168,In_1434);
nor U1161 (N_1161,In_2797,In_1189);
xnor U1162 (N_1162,N_599,In_2857);
nand U1163 (N_1163,In_2152,In_1409);
xor U1164 (N_1164,N_16,N_668);
and U1165 (N_1165,N_525,In_2789);
or U1166 (N_1166,In_652,In_1587);
nor U1167 (N_1167,N_138,In_1985);
nand U1168 (N_1168,N_249,N_705);
nand U1169 (N_1169,In_1503,N_351);
or U1170 (N_1170,N_874,In_88);
xor U1171 (N_1171,In_1501,N_137);
and U1172 (N_1172,In_328,In_2115);
and U1173 (N_1173,N_117,N_626);
or U1174 (N_1174,In_2347,In_1324);
nand U1175 (N_1175,In_2292,In_2808);
xnor U1176 (N_1176,N_731,N_686);
xor U1177 (N_1177,N_796,N_963);
and U1178 (N_1178,N_250,In_2433);
nand U1179 (N_1179,In_781,In_1405);
or U1180 (N_1180,In_693,N_58);
or U1181 (N_1181,In_2769,N_90);
xnor U1182 (N_1182,In_2601,In_2976);
or U1183 (N_1183,In_1716,N_167);
nor U1184 (N_1184,In_2447,N_558);
nand U1185 (N_1185,In_1507,N_82);
and U1186 (N_1186,In_628,In_151);
or U1187 (N_1187,In_1392,N_632);
and U1188 (N_1188,In_278,In_2940);
or U1189 (N_1189,N_362,In_2615);
and U1190 (N_1190,N_506,N_453);
or U1191 (N_1191,N_756,N_435);
xnor U1192 (N_1192,In_1864,N_400);
xor U1193 (N_1193,In_2397,N_607);
nand U1194 (N_1194,In_679,In_2267);
xor U1195 (N_1195,In_1696,In_1420);
and U1196 (N_1196,In_2419,N_432);
or U1197 (N_1197,N_313,In_1847);
nand U1198 (N_1198,N_693,In_2747);
or U1199 (N_1199,N_200,In_1351);
nor U1200 (N_1200,In_1397,N_50);
xnor U1201 (N_1201,In_2017,In_490);
or U1202 (N_1202,N_463,N_386);
xor U1203 (N_1203,N_976,In_736);
xor U1204 (N_1204,N_264,In_1766);
nand U1205 (N_1205,In_1897,In_421);
and U1206 (N_1206,In_976,In_253);
nor U1207 (N_1207,In_1034,In_997);
nor U1208 (N_1208,N_462,In_1169);
xor U1209 (N_1209,In_707,N_500);
xnor U1210 (N_1210,N_666,N_714);
or U1211 (N_1211,N_45,In_45);
and U1212 (N_1212,N_793,In_2510);
xor U1213 (N_1213,In_1010,N_991);
nand U1214 (N_1214,In_2955,N_779);
xnor U1215 (N_1215,In_1616,N_586);
and U1216 (N_1216,N_864,N_524);
xor U1217 (N_1217,In_1919,N_189);
nor U1218 (N_1218,N_392,In_2340);
xor U1219 (N_1219,In_2380,In_2588);
or U1220 (N_1220,In_1667,In_249);
or U1221 (N_1221,In_2622,In_1753);
nand U1222 (N_1222,In_1684,In_610);
nor U1223 (N_1223,N_353,In_143);
or U1224 (N_1224,In_947,In_2113);
or U1225 (N_1225,N_920,In_2048);
or U1226 (N_1226,In_1627,In_484);
nor U1227 (N_1227,In_1139,N_896);
nand U1228 (N_1228,In_1290,In_89);
nand U1229 (N_1229,N_552,In_1390);
xor U1230 (N_1230,N_887,In_2028);
or U1231 (N_1231,In_949,N_466);
nor U1232 (N_1232,In_2297,In_566);
and U1233 (N_1233,N_776,In_1965);
or U1234 (N_1234,In_2111,N_685);
nor U1235 (N_1235,In_2179,N_662);
nand U1236 (N_1236,In_2668,N_482);
or U1237 (N_1237,N_634,In_1935);
xnor U1238 (N_1238,In_853,In_379);
xnor U1239 (N_1239,In_277,In_1777);
or U1240 (N_1240,In_2533,N_785);
nor U1241 (N_1241,In_989,N_511);
nand U1242 (N_1242,N_268,N_854);
nor U1243 (N_1243,In_321,N_706);
or U1244 (N_1244,N_933,In_779);
nand U1245 (N_1245,In_2504,N_437);
nor U1246 (N_1246,N_510,In_2324);
nor U1247 (N_1247,In_2792,In_2242);
nor U1248 (N_1248,In_2694,In_971);
nand U1249 (N_1249,In_2927,In_1663);
xor U1250 (N_1250,In_305,In_2551);
nand U1251 (N_1251,In_977,N_792);
nand U1252 (N_1252,N_543,In_2109);
nor U1253 (N_1253,In_2777,N_617);
nor U1254 (N_1254,In_978,In_1370);
nand U1255 (N_1255,In_2228,In_2970);
or U1256 (N_1256,In_1240,In_2289);
nand U1257 (N_1257,N_717,N_989);
nand U1258 (N_1258,N_375,In_954);
nor U1259 (N_1259,In_2587,N_591);
xnor U1260 (N_1260,N_7,In_1637);
nor U1261 (N_1261,N_95,In_2540);
xnor U1262 (N_1262,In_992,N_819);
xor U1263 (N_1263,In_2118,N_868);
and U1264 (N_1264,In_230,N_170);
nor U1265 (N_1265,N_958,N_800);
and U1266 (N_1266,In_1611,In_289);
and U1267 (N_1267,N_812,In_371);
nand U1268 (N_1268,N_449,In_1609);
and U1269 (N_1269,In_2926,N_915);
xnor U1270 (N_1270,N_126,In_734);
and U1271 (N_1271,In_1918,N_562);
nand U1272 (N_1272,N_590,N_327);
or U1273 (N_1273,In_2650,N_183);
xnor U1274 (N_1274,In_1515,N_520);
xor U1275 (N_1275,N_704,N_899);
xor U1276 (N_1276,In_2869,In_1962);
nor U1277 (N_1277,N_561,In_2872);
nor U1278 (N_1278,In_483,In_2980);
and U1279 (N_1279,N_834,In_1170);
nor U1280 (N_1280,N_459,N_242);
nand U1281 (N_1281,In_1361,N_323);
nand U1282 (N_1282,In_710,In_2796);
and U1283 (N_1283,In_651,N_545);
or U1284 (N_1284,In_2378,N_824);
nand U1285 (N_1285,In_2975,N_604);
nand U1286 (N_1286,In_2275,In_883);
or U1287 (N_1287,N_425,In_2334);
and U1288 (N_1288,In_2212,N_56);
or U1289 (N_1289,In_581,N_643);
xnor U1290 (N_1290,N_133,N_335);
and U1291 (N_1291,N_270,N_9);
or U1292 (N_1292,N_79,In_445);
xor U1293 (N_1293,N_681,In_2280);
and U1294 (N_1294,N_973,In_907);
xor U1295 (N_1295,In_1280,In_2279);
nand U1296 (N_1296,N_803,N_584);
and U1297 (N_1297,In_1736,In_2373);
and U1298 (N_1298,N_729,In_1770);
nand U1299 (N_1299,In_2786,N_942);
or U1300 (N_1300,In_2163,In_2036);
nor U1301 (N_1301,In_2599,In_854);
nor U1302 (N_1302,N_542,In_2495);
nand U1303 (N_1303,In_21,In_1599);
or U1304 (N_1304,N_851,In_2073);
nor U1305 (N_1305,In_2707,In_236);
nand U1306 (N_1306,N_129,In_376);
nand U1307 (N_1307,N_711,In_845);
and U1308 (N_1308,In_1572,N_701);
xor U1309 (N_1309,In_1708,In_2180);
nand U1310 (N_1310,In_140,N_596);
nor U1311 (N_1311,N_866,In_2044);
nand U1312 (N_1312,In_1359,In_2429);
xnor U1313 (N_1313,In_43,N_934);
or U1314 (N_1314,In_1743,N_422);
or U1315 (N_1315,In_2062,N_947);
xor U1316 (N_1316,In_2736,N_143);
or U1317 (N_1317,N_699,In_830);
nor U1318 (N_1318,N_436,N_324);
and U1319 (N_1319,In_2593,In_1643);
nor U1320 (N_1320,N_457,In_2979);
nor U1321 (N_1321,In_624,In_2644);
xnor U1322 (N_1322,In_1830,In_608);
and U1323 (N_1323,N_847,N_777);
or U1324 (N_1324,N_257,In_2108);
nor U1325 (N_1325,In_1344,In_457);
or U1326 (N_1326,In_171,In_925);
xnor U1327 (N_1327,In_1608,In_2500);
nor U1328 (N_1328,In_2744,In_1580);
or U1329 (N_1329,N_925,N_759);
or U1330 (N_1330,In_2399,N_624);
or U1331 (N_1331,In_1642,In_2512);
or U1332 (N_1332,In_871,In_2413);
nor U1333 (N_1333,In_594,N_867);
nand U1334 (N_1334,In_2584,In_1004);
nor U1335 (N_1335,In_2829,In_2974);
xor U1336 (N_1336,In_1661,In_607);
and U1337 (N_1337,N_735,N_664);
nor U1338 (N_1338,In_2157,N_537);
or U1339 (N_1339,N_576,In_1554);
and U1340 (N_1340,In_2465,N_709);
and U1341 (N_1341,N_913,In_1908);
nand U1342 (N_1342,In_1968,N_679);
nor U1343 (N_1343,In_1805,In_279);
xor U1344 (N_1344,In_823,In_354);
xnor U1345 (N_1345,In_1478,N_585);
nand U1346 (N_1346,In_950,N_671);
or U1347 (N_1347,In_968,In_2241);
and U1348 (N_1348,In_2206,In_1277);
or U1349 (N_1349,In_2107,In_835);
and U1350 (N_1350,In_2051,N_260);
or U1351 (N_1351,In_551,In_1222);
and U1352 (N_1352,N_205,N_227);
nor U1353 (N_1353,N_37,In_1403);
nor U1354 (N_1354,In_1077,N_445);
and U1355 (N_1355,In_1703,In_1249);
nor U1356 (N_1356,In_1660,In_401);
nor U1357 (N_1357,N_259,In_1481);
or U1358 (N_1358,In_2321,In_2676);
or U1359 (N_1359,In_2009,In_2236);
and U1360 (N_1360,N_125,In_2159);
and U1361 (N_1361,N_529,N_898);
nor U1362 (N_1362,In_2437,N_320);
xnor U1363 (N_1363,In_1675,In_2992);
nor U1364 (N_1364,In_1199,In_220);
nor U1365 (N_1365,In_163,N_826);
xnor U1366 (N_1366,N_563,In_812);
nand U1367 (N_1367,N_85,In_2191);
nor U1368 (N_1368,N_912,In_2407);
nor U1369 (N_1369,In_560,In_2745);
nand U1370 (N_1370,N_544,N_215);
and U1371 (N_1371,In_2068,In_2473);
nor U1372 (N_1372,In_2770,N_740);
and U1373 (N_1373,In_389,N_889);
xnor U1374 (N_1374,N_648,In_2659);
nor U1375 (N_1375,In_2002,In_2768);
or U1376 (N_1376,N_27,In_856);
nand U1377 (N_1377,In_2060,In_400);
nand U1378 (N_1378,In_1922,In_700);
nand U1379 (N_1379,In_528,N_369);
nor U1380 (N_1380,In_387,In_2445);
xnor U1381 (N_1381,In_1803,In_290);
xnor U1382 (N_1382,In_2026,In_109);
nand U1383 (N_1383,In_604,N_364);
nand U1384 (N_1384,In_2416,N_38);
and U1385 (N_1385,In_1164,In_649);
or U1386 (N_1386,In_2248,N_870);
xnor U1387 (N_1387,N_540,In_2766);
xor U1388 (N_1388,In_1566,N_813);
and U1389 (N_1389,In_298,In_472);
and U1390 (N_1390,In_828,In_928);
nor U1391 (N_1391,In_248,N_797);
nor U1392 (N_1392,In_1090,N_725);
and U1393 (N_1393,In_537,In_1178);
nand U1394 (N_1394,In_453,In_1560);
or U1395 (N_1395,N_831,In_1410);
nand U1396 (N_1396,In_1063,In_846);
xor U1397 (N_1397,In_1116,N_589);
nand U1398 (N_1398,In_2877,N_830);
xor U1399 (N_1399,N_846,In_2764);
or U1400 (N_1400,In_1291,N_468);
nand U1401 (N_1401,In_844,In_2318);
nor U1402 (N_1402,In_763,In_1658);
nand U1403 (N_1403,N_289,N_979);
or U1404 (N_1404,In_2874,In_2350);
nand U1405 (N_1405,N_943,N_282);
nand U1406 (N_1406,In_2962,N_993);
and U1407 (N_1407,N_565,N_265);
xnor U1408 (N_1408,In_2509,In_146);
nor U1409 (N_1409,N_43,N_775);
nor U1410 (N_1410,In_2827,N_954);
nand U1411 (N_1411,In_2012,In_209);
or U1412 (N_1412,N_676,In_2734);
nand U1413 (N_1413,N_918,N_81);
or U1414 (N_1414,N_713,In_1942);
xnor U1415 (N_1415,In_2865,N_654);
and U1416 (N_1416,N_347,N_787);
xor U1417 (N_1417,In_1983,N_661);
and U1418 (N_1418,In_2986,N_601);
nand U1419 (N_1419,In_2229,In_1785);
nand U1420 (N_1420,In_247,In_142);
nor U1421 (N_1421,In_698,In_501);
xnor U1422 (N_1422,N_742,In_1241);
nand U1423 (N_1423,In_715,N_938);
and U1424 (N_1424,N_115,N_293);
nand U1425 (N_1425,In_292,N_91);
and U1426 (N_1426,N_266,N_344);
or U1427 (N_1427,In_2522,N_128);
or U1428 (N_1428,In_2061,N_914);
nor U1429 (N_1429,In_2828,N_784);
or U1430 (N_1430,In_349,In_2004);
xor U1431 (N_1431,In_1341,In_2620);
and U1432 (N_1432,N_978,In_339);
and U1433 (N_1433,In_892,In_2268);
and U1434 (N_1434,In_2899,In_87);
nand U1435 (N_1435,In_195,In_2977);
nand U1436 (N_1436,In_459,In_2358);
nor U1437 (N_1437,In_702,N_568);
nand U1438 (N_1438,N_904,In_1535);
and U1439 (N_1439,In_1823,In_1596);
or U1440 (N_1440,In_102,N_52);
xnor U1441 (N_1441,N_464,In_768);
or U1442 (N_1442,N_997,In_2895);
nand U1443 (N_1443,N_937,In_1372);
xor U1444 (N_1444,N_110,In_2554);
nor U1445 (N_1445,In_1318,N_158);
nand U1446 (N_1446,In_1064,In_217);
nor U1447 (N_1447,N_931,In_2312);
xor U1448 (N_1448,N_187,N_659);
nor U1449 (N_1449,N_554,In_1881);
nand U1450 (N_1450,N_902,In_2968);
and U1451 (N_1451,In_1583,N_491);
xor U1452 (N_1452,In_973,N_647);
nand U1453 (N_1453,In_2817,In_2135);
nand U1454 (N_1454,N_269,In_341);
or U1455 (N_1455,In_642,In_2569);
nor U1456 (N_1456,In_2428,N_623);
xor U1457 (N_1457,In_2032,In_2741);
or U1458 (N_1458,In_2114,N_986);
or U1459 (N_1459,In_1584,In_1352);
nor U1460 (N_1460,In_2031,N_737);
nor U1461 (N_1461,N_337,In_117);
nand U1462 (N_1462,N_821,In_1145);
xnor U1463 (N_1463,N_21,In_716);
xor U1464 (N_1464,In_1510,N_907);
or U1465 (N_1465,In_1498,In_479);
or U1466 (N_1466,In_836,In_262);
xor U1467 (N_1467,In_7,In_83);
or U1468 (N_1468,N_406,In_870);
or U1469 (N_1469,N_502,In_461);
nand U1470 (N_1470,In_56,In_2793);
xnor U1471 (N_1471,In_2042,In_1645);
nor U1472 (N_1472,In_906,In_1821);
and U1473 (N_1473,N_744,N_295);
nor U1474 (N_1474,In_147,N_745);
xor U1475 (N_1475,N_682,N_932);
and U1476 (N_1476,N_707,N_960);
nor U1477 (N_1477,N_614,N_688);
and U1478 (N_1478,In_1825,N_732);
and U1479 (N_1479,In_1274,N_959);
nand U1480 (N_1480,N_843,N_358);
and U1481 (N_1481,In_1886,In_1001);
or U1482 (N_1482,In_1713,In_2579);
xor U1483 (N_1483,N_823,In_884);
or U1484 (N_1484,N_940,In_1404);
nand U1485 (N_1485,N_600,N_184);
xor U1486 (N_1486,N_852,In_2246);
nand U1487 (N_1487,In_2339,N_401);
nor U1488 (N_1488,N_301,N_998);
nand U1489 (N_1489,N_332,In_2680);
and U1490 (N_1490,N_294,In_2164);
nor U1491 (N_1491,In_188,In_1725);
nand U1492 (N_1492,N_507,In_2178);
or U1493 (N_1493,In_2948,In_1380);
nand U1494 (N_1494,N_603,In_1124);
nand U1495 (N_1495,N_288,N_930);
and U1496 (N_1496,N_333,In_1137);
xnor U1497 (N_1497,N_559,In_2369);
xnor U1498 (N_1498,In_135,N_890);
or U1499 (N_1499,N_638,In_318);
nor U1500 (N_1500,In_1914,In_2494);
or U1501 (N_1501,N_1400,N_515);
xnor U1502 (N_1502,In_655,In_2567);
or U1503 (N_1503,N_1201,N_1120);
nand U1504 (N_1504,In_170,N_1405);
or U1505 (N_1505,In_2459,N_256);
nor U1506 (N_1506,In_2928,N_700);
or U1507 (N_1507,In_1516,N_1000);
xnor U1508 (N_1508,N_1310,In_744);
xor U1509 (N_1509,In_1804,N_1493);
and U1510 (N_1510,N_120,N_490);
nor U1511 (N_1511,N_822,N_560);
xor U1512 (N_1512,N_753,N_1409);
nand U1513 (N_1513,In_1406,N_675);
nand U1514 (N_1514,In_1479,N_1267);
xnor U1515 (N_1515,In_1068,N_1160);
nor U1516 (N_1516,In_51,N_1088);
and U1517 (N_1517,In_2189,In_1188);
xnor U1518 (N_1518,N_1018,N_592);
and U1519 (N_1519,N_606,N_528);
and U1520 (N_1520,In_198,In_9);
and U1521 (N_1521,In_1003,N_1312);
nand U1522 (N_1522,N_1073,In_2193);
nand U1523 (N_1523,N_1016,N_1417);
and U1524 (N_1524,N_703,N_1389);
nand U1525 (N_1525,N_64,In_639);
nand U1526 (N_1526,In_2704,N_1206);
or U1527 (N_1527,N_1198,N_1357);
and U1528 (N_1528,In_342,N_1347);
nor U1529 (N_1529,In_1925,In_1686);
nor U1530 (N_1530,N_1011,N_1114);
or U1531 (N_1531,N_988,N_855);
or U1532 (N_1532,N_921,In_1140);
nor U1533 (N_1533,N_924,In_653);
nor U1534 (N_1534,N_1433,N_741);
nor U1535 (N_1535,N_1141,N_1308);
nor U1536 (N_1536,In_1893,In_241);
and U1537 (N_1537,N_214,In_1878);
xnor U1538 (N_1538,In_1029,N_880);
nand U1539 (N_1539,N_1442,N_615);
xnor U1540 (N_1540,In_1721,N_1344);
xnor U1541 (N_1541,In_2818,N_493);
nor U1542 (N_1542,N_1338,In_1731);
xnor U1543 (N_1543,In_475,N_1421);
xor U1544 (N_1544,N_1460,N_746);
and U1545 (N_1545,N_1177,In_463);
and U1546 (N_1546,In_730,N_980);
and U1547 (N_1547,In_2603,N_734);
nand U1548 (N_1548,N_408,N_1032);
or U1549 (N_1549,N_116,N_1487);
and U1550 (N_1550,N_1358,N_1249);
or U1551 (N_1551,N_235,In_2756);
nand U1552 (N_1552,N_1025,In_79);
xnor U1553 (N_1553,N_923,In_2798);
or U1554 (N_1554,N_1169,N_1285);
nor U1555 (N_1555,In_1845,N_191);
nand U1556 (N_1556,N_1029,In_1364);
nor U1557 (N_1557,N_888,N_1070);
and U1558 (N_1558,In_2104,N_1225);
or U1559 (N_1559,N_1386,In_2502);
xor U1560 (N_1560,N_1227,N_12);
nand U1561 (N_1561,N_1475,N_827);
or U1562 (N_1562,N_1179,N_955);
xnor U1563 (N_1563,N_505,N_977);
nor U1564 (N_1564,N_1036,N_1383);
and U1565 (N_1565,In_2614,In_316);
nor U1566 (N_1566,In_2288,N_1272);
nand U1567 (N_1567,In_1381,N_1403);
nor U1568 (N_1568,N_1331,In_134);
and U1569 (N_1569,N_144,In_1973);
nor U1570 (N_1570,N_1246,N_882);
nor U1571 (N_1571,N_1350,In_1081);
nor U1572 (N_1572,In_491,In_1628);
nand U1573 (N_1573,N_17,In_2772);
nor U1574 (N_1574,N_388,In_73);
xnor U1575 (N_1575,N_518,In_1890);
xnor U1576 (N_1576,In_1149,In_1938);
nand U1577 (N_1577,In_348,N_1336);
nand U1578 (N_1578,N_990,N_1123);
or U1579 (N_1579,N_1498,N_1489);
or U1580 (N_1580,N_1112,N_670);
nand U1581 (N_1581,In_1958,N_1298);
xor U1582 (N_1582,N_1373,In_701);
and U1583 (N_1583,N_61,N_1283);
nor U1584 (N_1584,N_577,N_1499);
nand U1585 (N_1585,N_1062,In_1100);
nor U1586 (N_1586,In_2351,N_555);
nand U1587 (N_1587,N_672,N_1218);
nand U1588 (N_1588,N_1172,N_1325);
and U1589 (N_1589,In_420,N_1327);
and U1590 (N_1590,In_2239,N_975);
and U1591 (N_1591,N_272,In_97);
and U1592 (N_1592,In_2631,N_1232);
or U1593 (N_1593,In_1921,N_956);
nand U1594 (N_1594,N_1393,N_1037);
or U1595 (N_1595,N_723,N_1271);
and U1596 (N_1596,N_891,In_2909);
or U1597 (N_1597,In_658,In_578);
xor U1598 (N_1598,N_673,N_429);
nand U1599 (N_1599,N_1273,N_1049);
nor U1600 (N_1600,In_2308,N_818);
or U1601 (N_1601,In_1715,In_951);
xor U1602 (N_1602,In_1465,N_1387);
nand U1603 (N_1603,In_131,N_11);
nor U1604 (N_1604,In_822,N_378);
and U1605 (N_1605,N_1146,N_1332);
or U1606 (N_1606,N_917,N_1152);
and U1607 (N_1607,N_438,N_1248);
xnor U1608 (N_1608,N_1268,N_1316);
nor U1609 (N_1609,N_1128,N_228);
or U1610 (N_1610,N_1470,N_1352);
or U1611 (N_1611,N_722,N_1001);
nor U1612 (N_1612,N_724,In_2262);
and U1613 (N_1613,N_1439,In_1412);
and U1614 (N_1614,In_1203,In_2005);
nor U1615 (N_1615,N_201,In_2120);
xnor U1616 (N_1616,N_363,In_1748);
xnor U1617 (N_1617,In_1414,N_1065);
nor U1618 (N_1618,In_1210,In_2594);
and U1619 (N_1619,In_1387,In_2761);
or U1620 (N_1620,N_1121,In_575);
and U1621 (N_1621,In_1216,N_566);
nand U1622 (N_1622,N_1279,In_127);
and U1623 (N_1623,N_1086,In_1541);
nor U1624 (N_1624,N_1481,N_239);
xor U1625 (N_1625,In_1211,In_941);
and U1626 (N_1626,In_885,In_2889);
or U1627 (N_1627,In_1947,N_1445);
xnor U1628 (N_1628,N_1461,In_1895);
xor U1629 (N_1629,In_739,N_908);
nor U1630 (N_1630,N_30,In_688);
or U1631 (N_1631,N_504,N_1183);
nand U1632 (N_1632,N_547,In_2058);
nor U1633 (N_1633,N_982,In_851);
or U1634 (N_1634,In_326,In_1032);
nand U1635 (N_1635,N_1038,In_2583);
nor U1636 (N_1636,N_513,In_1323);
nand U1637 (N_1637,In_1712,In_1284);
and U1638 (N_1638,In_2346,N_421);
nand U1639 (N_1639,In_2128,N_1022);
or U1640 (N_1640,In_596,In_754);
or U1641 (N_1641,In_1346,N_916);
or U1642 (N_1642,In_2993,N_373);
nor U1643 (N_1643,N_1260,In_785);
nor U1644 (N_1644,In_1771,In_180);
nor U1645 (N_1645,N_992,N_1446);
nor U1646 (N_1646,In_1492,In_2719);
and U1647 (N_1647,In_1449,In_972);
or U1648 (N_1648,N_262,In_2989);
or U1649 (N_1649,N_1287,N_949);
xnor U1650 (N_1650,N_588,N_1115);
or U1651 (N_1651,N_1281,In_240);
xor U1652 (N_1652,In_2794,In_1332);
or U1653 (N_1653,In_1076,N_203);
or U1654 (N_1654,N_1153,N_557);
nor U1655 (N_1655,N_512,N_478);
xor U1656 (N_1656,N_1189,N_1414);
or U1657 (N_1657,In_2642,N_1182);
nor U1658 (N_1658,In_921,In_1368);
and U1659 (N_1659,N_637,N_1217);
xnor U1660 (N_1660,N_789,N_1447);
and U1661 (N_1661,In_2706,In_1820);
and U1662 (N_1662,N_391,N_1297);
xor U1663 (N_1663,In_1619,N_892);
xnor U1664 (N_1664,N_527,In_1293);
nand U1665 (N_1665,N_749,In_336);
or U1666 (N_1666,N_1300,In_1396);
or U1667 (N_1667,N_771,In_974);
nor U1668 (N_1668,In_765,In_94);
xor U1669 (N_1669,N_1072,In_176);
nand U1670 (N_1670,In_2929,N_92);
and U1671 (N_1671,N_853,In_470);
nand U1672 (N_1672,N_620,N_1052);
nand U1673 (N_1673,N_687,In_1558);
and U1674 (N_1674,N_1137,N_1349);
or U1675 (N_1675,In_1726,In_957);
nand U1676 (N_1676,In_276,N_712);
or U1677 (N_1677,In_101,N_721);
nor U1678 (N_1678,N_1377,N_1051);
or U1679 (N_1679,In_901,N_953);
nor U1680 (N_1680,N_1410,N_1192);
xor U1681 (N_1681,N_1092,N_1173);
nand U1682 (N_1682,In_1633,In_838);
nor U1683 (N_1683,N_571,N_1103);
and U1684 (N_1684,In_961,N_708);
nor U1685 (N_1685,N_750,In_357);
nand U1686 (N_1686,N_509,N_1107);
and U1687 (N_1687,N_131,In_638);
or U1688 (N_1688,N_1313,N_1007);
nand U1689 (N_1689,N_835,N_412);
nand U1690 (N_1690,N_1462,N_1216);
xnor U1691 (N_1691,In_2886,N_297);
nand U1692 (N_1692,N_663,N_1135);
or U1693 (N_1693,N_336,In_1610);
or U1694 (N_1694,N_164,N_1419);
or U1695 (N_1695,N_1209,In_2261);
nor U1696 (N_1696,In_158,In_1156);
nor U1697 (N_1697,In_2474,N_727);
nand U1698 (N_1698,N_1060,In_1255);
nand U1699 (N_1699,In_26,N_635);
and U1700 (N_1700,N_536,In_2006);
xnor U1701 (N_1701,N_972,In_1916);
xnor U1702 (N_1702,In_1527,N_1130);
or U1703 (N_1703,In_2138,In_2348);
nand U1704 (N_1704,N_593,N_910);
nor U1705 (N_1705,In_2151,In_939);
xor U1706 (N_1706,In_2232,N_655);
nor U1707 (N_1707,In_2547,N_379);
and U1708 (N_1708,N_1305,N_1256);
or U1709 (N_1709,N_1054,N_1496);
nor U1710 (N_1710,In_2094,N_832);
nor U1711 (N_1711,N_1004,In_780);
nand U1712 (N_1712,N_844,N_1427);
nor U1713 (N_1713,N_783,In_2091);
nand U1714 (N_1714,In_297,In_1455);
nand U1715 (N_1715,In_1659,In_1162);
nor U1716 (N_1716,N_1089,N_760);
nor U1717 (N_1717,In_2573,N_1398);
nor U1718 (N_1718,N_1399,In_76);
and U1719 (N_1719,N_1323,N_1031);
or U1720 (N_1720,N_767,In_62);
nor U1721 (N_1721,In_1625,N_791);
nand U1722 (N_1722,N_180,N_36);
or U1723 (N_1723,N_1212,In_2902);
nand U1724 (N_1724,In_1248,In_773);
nor U1725 (N_1725,In_673,In_1691);
and U1726 (N_1726,N_22,N_801);
nand U1727 (N_1727,N_952,N_957);
nor U1728 (N_1728,In_1571,N_961);
xor U1729 (N_1729,N_1015,In_1330);
xnor U1730 (N_1730,N_1291,N_1196);
nor U1731 (N_1731,N_1230,In_2575);
or U1732 (N_1732,In_2810,N_790);
nand U1733 (N_1733,In_2723,In_645);
nand U1734 (N_1734,In_1468,N_1156);
or U1735 (N_1735,In_2825,N_1364);
xnor U1736 (N_1736,N_1381,In_2515);
xor U1737 (N_1737,N_1020,In_2568);
xnor U1738 (N_1738,N_1228,In_1879);
nor U1739 (N_1739,N_922,N_1471);
or U1740 (N_1740,N_20,N_1483);
nor U1741 (N_1741,N_2,In_510);
nor U1742 (N_1742,In_1767,In_488);
nor U1743 (N_1743,N_1353,N_1275);
nor U1744 (N_1744,N_720,N_252);
nand U1745 (N_1745,N_1455,N_1286);
nand U1746 (N_1746,N_1415,N_501);
and U1747 (N_1747,In_1238,N_1339);
and U1748 (N_1748,In_740,N_166);
and U1749 (N_1749,N_770,In_1917);
and U1750 (N_1750,N_149,N_969);
xnor U1751 (N_1751,In_1647,N_1057);
or U1752 (N_1752,In_2353,In_903);
nor U1753 (N_1753,In_2838,N_814);
or U1754 (N_1754,N_1058,N_1486);
or U1755 (N_1755,In_2973,In_2702);
nand U1756 (N_1756,N_1341,N_1186);
or U1757 (N_1757,In_1201,In_2417);
nand U1758 (N_1758,N_1093,In_473);
xnor U1759 (N_1759,N_1175,N_1394);
nand U1760 (N_1760,In_232,In_2665);
xor U1761 (N_1761,N_442,In_2195);
nand U1762 (N_1762,N_1485,N_195);
nor U1763 (N_1763,In_2526,In_2103);
nand U1764 (N_1764,In_902,N_24);
or U1765 (N_1765,In_1856,N_1282);
xnor U1766 (N_1766,N_534,N_1237);
xnor U1767 (N_1767,N_446,In_33);
nand U1768 (N_1768,In_1250,N_98);
or U1769 (N_1769,N_1314,N_1397);
nand U1770 (N_1770,N_1203,In_2619);
nor U1771 (N_1771,In_2270,In_1557);
xnor U1772 (N_1772,N_1366,N_1380);
and U1773 (N_1773,N_1416,N_862);
nor U1774 (N_1774,In_2252,N_1045);
nand U1775 (N_1775,N_1317,In_1756);
xor U1776 (N_1776,N_1407,N_897);
nor U1777 (N_1777,N_1042,N_1180);
or U1778 (N_1778,N_319,N_641);
or U1779 (N_1779,N_1028,N_1371);
nand U1780 (N_1780,In_1982,N_657);
xnor U1781 (N_1781,N_46,N_1252);
xnor U1782 (N_1782,In_1024,N_188);
and U1783 (N_1783,In_2883,N_1082);
xnor U1784 (N_1784,N_642,In_1350);
xor U1785 (N_1785,N_548,In_602);
xnor U1786 (N_1786,N_798,N_1269);
and U1787 (N_1787,N_769,In_2749);
and U1788 (N_1788,In_1836,N_163);
nand U1789 (N_1789,In_2624,In_1349);
nor U1790 (N_1790,In_523,N_1185);
and U1791 (N_1791,N_1118,In_579);
or U1792 (N_1792,N_833,In_1012);
or U1793 (N_1793,N_1492,N_1178);
and U1794 (N_1794,In_2778,N_1207);
nand U1795 (N_1795,In_329,In_2234);
nand U1796 (N_1796,N_1098,N_1465);
nand U1797 (N_1797,In_2864,N_726);
nor U1798 (N_1798,N_730,In_2684);
xnor U1799 (N_1799,N_1063,N_1302);
and U1800 (N_1800,In_606,In_2539);
xnor U1801 (N_1801,N_950,In_1505);
nand U1802 (N_1802,N_653,In_663);
and U1803 (N_1803,In_1784,N_471);
nor U1804 (N_1804,In_1307,In_1615);
and U1805 (N_1805,N_1376,N_575);
or U1806 (N_1806,N_1318,N_44);
nand U1807 (N_1807,N_1116,In_2081);
or U1808 (N_1808,In_2491,In_2046);
nor U1809 (N_1809,N_752,In_738);
and U1810 (N_1810,N_1342,N_639);
and U1811 (N_1811,In_737,In_234);
and U1812 (N_1812,In_1939,In_1437);
nand U1813 (N_1813,N_194,N_1259);
xnor U1814 (N_1814,N_1438,N_1133);
and U1815 (N_1815,N_1497,In_2941);
xnor U1816 (N_1816,N_1404,N_1048);
xnor U1817 (N_1817,In_2300,N_1125);
nor U1818 (N_1818,N_1210,N_1162);
xor U1819 (N_1819,N_172,N_1233);
nor U1820 (N_1820,N_1043,In_743);
nor U1821 (N_1821,N_41,In_450);
and U1822 (N_1822,In_2809,N_875);
nand U1823 (N_1823,In_1303,N_884);
nand U1824 (N_1824,In_515,In_20);
nand U1825 (N_1825,N_893,N_1145);
and U1826 (N_1826,N_255,N_1469);
nor U1827 (N_1827,In_2945,N_1330);
nor U1828 (N_1828,In_1321,N_1213);
xnor U1829 (N_1829,In_1737,N_1041);
xnor U1830 (N_1830,N_209,N_1333);
nor U1831 (N_1831,N_207,N_399);
or U1832 (N_1832,N_1161,In_1148);
xor U1833 (N_1833,N_1384,In_23);
xnor U1834 (N_1834,N_1046,N_1309);
nor U1835 (N_1835,In_2562,N_764);
and U1836 (N_1836,In_2632,In_667);
nand U1837 (N_1837,In_476,N_1124);
nor U1838 (N_1838,N_1432,In_111);
nand U1839 (N_1839,N_879,N_1085);
nand U1840 (N_1840,N_1155,N_1214);
xnor U1841 (N_1841,N_583,N_1477);
xnor U1842 (N_1842,N_1019,In_552);
and U1843 (N_1843,N_202,In_865);
nor U1844 (N_1844,N_861,N_287);
or U1845 (N_1845,N_146,N_1301);
or U1846 (N_1846,N_106,N_1494);
and U1847 (N_1847,N_680,N_1335);
nor U1848 (N_1848,In_250,N_532);
nand U1849 (N_1849,In_634,In_107);
or U1850 (N_1850,N_1385,N_1110);
and U1851 (N_1851,N_1289,N_845);
nand U1852 (N_1852,N_1033,N_0);
and U1853 (N_1853,N_595,N_658);
and U1854 (N_1854,In_2127,In_105);
nand U1855 (N_1855,N_1066,N_743);
xnor U1856 (N_1856,N_34,N_1080);
and U1857 (N_1857,In_554,N_1221);
or U1858 (N_1858,N_1311,N_1343);
nand U1859 (N_1859,In_2434,N_1429);
or U1860 (N_1860,N_581,N_340);
nor U1861 (N_1861,In_1741,N_1102);
xor U1862 (N_1862,N_1307,In_897);
nand U1863 (N_1863,In_1929,In_2490);
xor U1864 (N_1864,N_1117,In_875);
xnor U1865 (N_1865,N_1355,In_849);
xor U1866 (N_1866,In_2020,N_1367);
or U1867 (N_1867,N_886,In_356);
nand U1868 (N_1868,N_1219,N_251);
xnor U1869 (N_1869,N_1143,N_1);
nor U1870 (N_1870,In_1680,N_159);
or U1871 (N_1871,N_1194,N_1490);
and U1872 (N_1872,N_587,In_2790);
or U1873 (N_1873,N_817,N_929);
nor U1874 (N_1874,N_894,N_1370);
nand U1875 (N_1875,In_970,In_1125);
or U1876 (N_1876,In_287,N_858);
nor U1877 (N_1877,N_569,N_1132);
and U1878 (N_1878,In_2439,In_2327);
and U1879 (N_1879,N_696,N_608);
nor U1880 (N_1880,N_1056,N_971);
nor U1881 (N_1881,N_1104,N_1356);
and U1882 (N_1882,N_59,In_2379);
or U1883 (N_1883,N_1422,N_598);
xnor U1884 (N_1884,In_6,N_967);
nand U1885 (N_1885,In_909,In_2100);
and U1886 (N_1886,N_1142,In_500);
nor U1887 (N_1887,In_1513,N_1412);
and U1888 (N_1888,N_460,N_1204);
nor U1889 (N_1889,N_1106,N_1138);
xnor U1890 (N_1890,N_1328,N_1149);
nor U1891 (N_1891,N_13,In_2816);
nand U1892 (N_1892,N_859,In_2623);
nor U1893 (N_1893,N_1109,In_791);
xnor U1894 (N_1894,In_803,N_1096);
or U1895 (N_1895,N_1165,N_384);
xnor U1896 (N_1896,N_434,N_1478);
xor U1897 (N_1897,In_526,N_1476);
nor U1898 (N_1898,In_1801,In_58);
or U1899 (N_1899,In_1514,N_1220);
nand U1900 (N_1900,N_1108,In_373);
xor U1901 (N_1901,N_1435,N_1495);
nor U1902 (N_1902,In_1288,In_586);
xnor U1903 (N_1903,N_1097,N_692);
nand U1904 (N_1904,N_514,N_1395);
or U1905 (N_1905,N_869,In_1975);
or U1906 (N_1906,N_1200,In_2001);
nor U1907 (N_1907,In_1347,In_641);
nand U1908 (N_1908,N_397,In_1);
and U1909 (N_1909,N_1068,In_2315);
nand U1910 (N_1910,N_1147,In_98);
xor U1911 (N_1911,In_2382,N_1284);
and U1912 (N_1912,N_618,In_820);
or U1913 (N_1913,In_1846,N_857);
nor U1914 (N_1914,N_1488,In_1377);
nor U1915 (N_1915,In_1877,In_1448);
or U1916 (N_1916,N_1482,N_619);
xnor U1917 (N_1917,N_984,N_1127);
or U1918 (N_1918,In_1195,N_1340);
nand U1919 (N_1919,N_1039,In_439);
nand U1920 (N_1920,N_1265,N_865);
nand U1921 (N_1921,N_226,In_1176);
and U1922 (N_1922,N_8,N_186);
xor U1923 (N_1923,N_1205,N_484);
nor U1924 (N_1924,In_946,In_157);
nor U1925 (N_1925,N_1017,In_2149);
nand U1926 (N_1926,In_1521,In_2963);
nand U1927 (N_1927,In_2256,N_1199);
xor U1928 (N_1928,In_987,In_2190);
xnor U1929 (N_1929,N_1484,N_535);
or U1930 (N_1930,In_547,In_1632);
nor U1931 (N_1931,N_1164,N_1294);
xnor U1932 (N_1932,In_2349,N_1244);
nand U1933 (N_1933,In_1500,N_1134);
nor U1934 (N_1934,In_2258,N_829);
xor U1935 (N_1935,N_605,N_1466);
and U1936 (N_1936,N_1129,N_1157);
and U1937 (N_1937,N_678,N_176);
and U1938 (N_1938,N_738,N_1374);
and U1939 (N_1939,In_1218,N_630);
nand U1940 (N_1940,In_2923,In_219);
xnor U1941 (N_1941,In_478,In_2570);
or U1942 (N_1942,N_139,In_1702);
and U1943 (N_1943,N_677,N_1392);
xnor U1944 (N_1944,N_32,N_694);
and U1945 (N_1945,N_629,In_2266);
nor U1946 (N_1946,In_2812,N_609);
nor U1947 (N_1947,In_2550,In_1597);
and U1948 (N_1948,In_899,N_1276);
nor U1949 (N_1949,N_1296,In_449);
and U1950 (N_1950,N_1428,N_778);
xor U1951 (N_1951,N_285,In_1723);
and U1952 (N_1952,N_941,N_1079);
and U1953 (N_1953,N_1030,N_178);
or U1954 (N_1954,N_1288,In_521);
xnor U1955 (N_1955,N_1444,N_1420);
and U1956 (N_1956,N_360,In_676);
or U1957 (N_1957,N_1159,N_1148);
xnor U1958 (N_1958,N_1050,In_890);
or U1959 (N_1959,N_553,N_698);
nor U1960 (N_1960,N_1434,In_1701);
and U1961 (N_1961,In_2294,N_1261);
nand U1962 (N_1962,N_1458,In_78);
and U1963 (N_1963,N_716,In_2331);
xor U1964 (N_1964,N_1348,In_114);
and U1965 (N_1965,N_582,N_1094);
nor U1966 (N_1966,N_1197,In_593);
nand U1967 (N_1967,N_1239,N_443);
nor U1968 (N_1968,N_1351,N_423);
nand U1969 (N_1969,N_926,N_1467);
or U1970 (N_1970,N_839,N_1168);
xor U1971 (N_1971,In_1423,In_71);
xor U1972 (N_1972,In_1644,N_1436);
and U1973 (N_1973,In_1142,In_2025);
nor U1974 (N_1974,In_50,In_721);
xor U1975 (N_1975,N_1379,N_850);
nor U1976 (N_1976,N_1083,N_1354);
and U1977 (N_1977,N_1191,In_2529);
nand U1978 (N_1978,N_622,N_1236);
and U1979 (N_1979,In_1135,In_166);
nand U1980 (N_1980,In_141,N_349);
or U1981 (N_1981,N_526,In_966);
nor U1982 (N_1982,N_1396,In_2422);
and U1983 (N_1983,N_1424,In_2960);
or U1984 (N_1984,In_1043,In_1875);
and U1985 (N_1985,In_1992,In_2543);
and U1986 (N_1986,N_935,N_1167);
or U1987 (N_1987,N_1270,In_2611);
nor U1988 (N_1988,In_1775,N_1035);
nand U1989 (N_1989,N_322,N_389);
nand U1990 (N_1990,N_1208,In_1957);
nand U1991 (N_1991,N_780,N_1163);
and U1992 (N_1992,N_204,In_1837);
nor U1993 (N_1993,N_1324,N_757);
nand U1994 (N_1994,In_694,N_805);
xor U1995 (N_1995,In_1287,N_1224);
nor U1996 (N_1996,In_807,N_1450);
xor U1997 (N_1997,In_2589,In_365);
and U1998 (N_1998,In_139,In_90);
nor U1999 (N_1999,N_1078,In_1220);
or U2000 (N_2000,N_928,N_936);
and U2001 (N_2001,In_935,N_1747);
or U2002 (N_2002,N_1617,N_1423);
and U2003 (N_2003,N_1969,N_1874);
and U2004 (N_2004,N_1235,N_1695);
nor U2005 (N_2005,In_1378,N_1826);
or U2006 (N_2006,N_1568,N_1520);
or U2007 (N_2007,N_1543,N_1945);
xnor U2008 (N_2008,N_75,In_503);
or U2009 (N_2009,N_1095,N_312);
nor U2010 (N_2010,N_1594,In_2908);
or U2011 (N_2011,N_919,N_1696);
xnor U2012 (N_2012,N_1660,N_1136);
or U2013 (N_2013,N_944,N_1508);
and U2014 (N_2014,N_1457,N_1955);
or U2015 (N_2015,N_1805,N_1840);
and U2016 (N_2016,In_982,N_1962);
xnor U2017 (N_2017,N_1686,N_763);
or U2018 (N_2018,N_1292,N_1613);
nand U2019 (N_2019,N_1382,In_825);
or U2020 (N_2020,N_1507,N_175);
or U2021 (N_2021,N_1013,N_1977);
and U2022 (N_2022,N_1801,N_1992);
nand U2023 (N_2023,N_1634,N_1578);
xor U2024 (N_2024,In_308,N_1010);
or U2025 (N_2025,N_1334,N_1770);
or U2026 (N_2026,N_1583,N_1648);
nor U2027 (N_2027,N_1732,N_1949);
or U2028 (N_2028,N_1061,N_1774);
xnor U2029 (N_2029,N_1642,N_1827);
and U2030 (N_2030,N_1337,In_1067);
and U2031 (N_2031,N_1069,N_810);
or U2032 (N_2032,N_1876,N_433);
or U2033 (N_2033,In_16,N_1555);
nand U2034 (N_2034,N_1527,N_1599);
and U2035 (N_2035,N_1504,N_1505);
xnor U2036 (N_2036,N_1965,N_1939);
nand U2037 (N_2037,In_474,N_1615);
nand U2038 (N_2038,In_1399,N_1119);
nor U2039 (N_2039,N_486,N_567);
and U2040 (N_2040,N_1649,N_1914);
xor U2041 (N_2041,N_1783,N_1658);
xor U2042 (N_2042,N_786,N_1074);
or U2043 (N_2043,N_1580,N_1961);
or U2044 (N_2044,N_1786,In_2669);
or U2045 (N_2045,N_1454,In_228);
nor U2046 (N_2046,N_739,N_1766);
nand U2047 (N_2047,N_1587,N_1087);
and U2048 (N_2048,N_651,N_856);
nor U2049 (N_2049,N_1884,N_1739);
nand U2050 (N_2050,In_2146,N_1867);
nand U2051 (N_2051,N_1712,N_1877);
or U2052 (N_2052,In_1037,N_808);
nand U2053 (N_2053,In_2182,N_1645);
nor U2054 (N_2054,N_35,N_523);
xnor U2055 (N_2055,N_1591,N_768);
nand U2056 (N_2056,N_1953,N_1315);
xor U2057 (N_2057,N_1612,N_1998);
nand U2058 (N_2058,N_1665,N_1790);
and U2059 (N_2059,N_305,In_2446);
nand U2060 (N_2060,N_802,N_1807);
nor U2061 (N_2061,N_1863,N_1973);
nor U2062 (N_2062,N_1988,N_1948);
nand U2063 (N_2063,N_1793,N_1595);
nor U2064 (N_2064,N_996,N_1818);
nor U2065 (N_2065,N_1873,N_1077);
and U2066 (N_2066,N_1559,N_1630);
nand U2067 (N_2067,N_811,N_1720);
nand U2068 (N_2068,N_1139,In_2282);
nor U2069 (N_2069,In_2029,N_1554);
and U2070 (N_2070,N_465,In_1345);
xor U2071 (N_2071,N_1602,N_1549);
and U2072 (N_2072,N_1544,In_1109);
nand U2073 (N_2073,N_1718,N_1105);
xnor U2074 (N_2074,In_1810,N_440);
xor U2075 (N_2075,In_1283,N_1845);
nand U2076 (N_2076,N_229,N_1750);
and U2077 (N_2077,N_1245,N_1907);
nand U2078 (N_2078,N_995,N_1808);
xor U2079 (N_2079,N_1859,N_1709);
nand U2080 (N_2080,N_1878,In_1456);
nand U2081 (N_2081,N_1740,N_1569);
nor U2082 (N_2082,N_47,N_1653);
xor U2083 (N_2083,N_1822,N_1576);
and U2084 (N_2084,N_1474,In_1152);
nor U2085 (N_2085,N_1368,N_1902);
nor U2086 (N_2086,N_1525,N_1655);
nor U2087 (N_2087,N_1550,In_2197);
or U2088 (N_2088,N_1837,N_1875);
nand U2089 (N_2089,In_1379,N_1306);
and U2090 (N_2090,N_1008,N_1593);
xor U2091 (N_2091,In_1880,In_2365);
and U2092 (N_2092,N_539,In_1398);
xnor U2093 (N_2093,In_424,In_2034);
and U2094 (N_2094,N_1034,In_1069);
nor U2095 (N_2095,N_1683,N_1663);
nor U2096 (N_2096,In_1841,N_1603);
nor U2097 (N_2097,In_1477,N_1908);
and U2098 (N_2098,N_1150,N_519);
nor U2099 (N_2099,In_2538,N_1980);
and U2100 (N_2100,In_1605,In_2255);
xnor U2101 (N_2101,N_1743,N_1262);
and U2102 (N_2102,N_640,In_2235);
and U2103 (N_2103,In_2116,N_1459);
nand U2104 (N_2104,In_193,In_1147);
nor U2105 (N_2105,N_1441,N_901);
xor U2106 (N_2106,N_1211,N_1503);
nand U2107 (N_2107,N_405,N_1763);
and U2108 (N_2108,N_1629,In_1310);
or U2109 (N_2109,In_2341,In_1866);
or U2110 (N_2110,N_1053,N_1705);
nand U2111 (N_2111,N_1664,N_1745);
nor U2112 (N_2112,N_1813,N_1851);
xor U2113 (N_2113,N_1622,N_1778);
nor U2114 (N_2114,N_196,N_1754);
xor U2115 (N_2115,In_728,N_962);
nor U2116 (N_2116,N_1676,N_660);
and U2117 (N_2117,N_1848,In_2176);
or U2118 (N_2118,In_1219,N_1999);
or U2119 (N_2119,N_1473,N_1426);
or U2120 (N_2120,N_1151,In_967);
nand U2121 (N_2121,N_1391,N_1943);
or U2122 (N_2122,N_1654,N_1855);
xnor U2123 (N_2123,N_613,N_1985);
nor U2124 (N_2124,N_1556,N_1994);
and U2125 (N_2125,N_1677,N_104);
nand U2126 (N_2126,N_1295,N_1979);
or U2127 (N_2127,In_1020,N_1730);
or U2128 (N_2128,In_531,N_1987);
nor U2129 (N_2129,N_636,N_999);
nor U2130 (N_2130,N_1453,N_1044);
nor U2131 (N_2131,N_795,N_1952);
xnor U2132 (N_2132,In_2078,N_1264);
nor U2133 (N_2133,In_2850,N_900);
xnor U2134 (N_2134,In_2438,N_503);
nor U2135 (N_2135,N_1574,N_966);
nand U2136 (N_2136,N_1853,N_1891);
or U2137 (N_2137,N_1263,N_1944);
nor U2138 (N_2138,N_1755,N_1865);
and U2139 (N_2139,In_2693,N_1247);
xnor U2140 (N_2140,In_1180,N_1843);
xor U2141 (N_2141,N_1862,N_1917);
and U2142 (N_2142,N_1684,In_438);
nand U2143 (N_2143,N_426,N_1322);
or U2144 (N_2144,N_1215,N_1700);
and U2145 (N_2145,N_1997,In_1395);
xor U2146 (N_2146,N_1806,N_1250);
and U2147 (N_2147,N_1685,N_1942);
xnor U2148 (N_2148,N_1021,In_1758);
nand U2149 (N_2149,N_1360,In_2708);
nand U2150 (N_2150,N_1579,N_1668);
and U2151 (N_2151,N_1586,N_1632);
xor U2152 (N_2152,N_728,N_1794);
nand U2153 (N_2153,N_1611,N_718);
xnor U2154 (N_2154,N_1834,N_1738);
or U2155 (N_2155,N_736,N_1737);
and U2156 (N_2156,N_1537,In_2271);
or U2157 (N_2157,N_1798,N_1644);
nand U2158 (N_2158,N_247,N_1925);
nor U2159 (N_2159,N_1547,N_1577);
nor U2160 (N_2160,N_1989,N_1717);
nand U2161 (N_2161,In_296,N_1690);
xnor U2162 (N_2162,N_633,N_1882);
xnor U2163 (N_2163,N_1701,N_1518);
and U2164 (N_2164,N_1858,N_1601);
xor U2165 (N_2165,N_1931,In_437);
and U2166 (N_2166,N_1976,In_2639);
and U2167 (N_2167,N_1536,In_1824);
nand U2168 (N_2168,N_667,N_1009);
xor U2169 (N_2169,N_1761,N_1620);
nand U2170 (N_2170,In_852,N_1736);
xnor U2171 (N_2171,N_107,In_1177);
nand U2172 (N_2172,N_1290,N_772);
nand U2173 (N_2173,N_1637,N_1675);
nor U2174 (N_2174,In_103,N_1959);
or U2175 (N_2175,N_1759,N_1975);
xnor U2176 (N_2176,N_1266,N_1006);
nand U2177 (N_2177,N_1363,In_1160);
xnor U2178 (N_2178,In_2513,N_508);
and U2179 (N_2179,N_1627,N_1562);
or U2180 (N_2180,N_1780,N_1598);
nand U2181 (N_2181,N_1014,N_1934);
and U2182 (N_2182,N_1304,In_1526);
nand U2183 (N_2183,N_1919,N_1929);
nor U2184 (N_2184,In_1309,N_1693);
nand U2185 (N_2185,N_1829,N_1506);
and U2186 (N_2186,In_564,N_1661);
nand U2187 (N_2187,In_520,In_2364);
xnor U2188 (N_2188,N_1772,N_968);
and U2189 (N_2189,N_309,N_1480);
nand U2190 (N_2190,In_1570,N_1408);
nand U2191 (N_2191,N_114,N_1369);
or U2192 (N_2192,N_1861,N_541);
xnor U2193 (N_2193,In_2634,N_1918);
or U2194 (N_2194,In_2418,In_630);
or U2195 (N_2195,In_991,N_1464);
nor U2196 (N_2196,N_475,N_1938);
or U2197 (N_2197,N_1625,N_1539);
and U2198 (N_2198,N_1892,In_988);
or U2199 (N_2199,N_1767,N_1560);
nor U2200 (N_2200,N_1864,N_521);
nor U2201 (N_2201,In_323,N_231);
xor U2202 (N_2202,N_1511,N_1243);
xor U2203 (N_2203,N_1456,N_1940);
and U2204 (N_2204,N_985,N_495);
nor U2205 (N_2205,N_65,N_1023);
nand U2206 (N_2206,N_1697,N_1669);
or U2207 (N_2207,N_1760,N_1468);
nand U2208 (N_2208,In_672,N_387);
or U2209 (N_2209,N_1691,In_272);
or U2210 (N_2210,In_1251,N_1903);
nor U2211 (N_2211,N_1756,N_173);
xnor U2212 (N_2212,N_690,N_1901);
nand U2213 (N_2213,N_1836,In_2007);
and U2214 (N_2214,N_1657,N_1707);
nand U2215 (N_2215,N_1623,In_1711);
and U2216 (N_2216,In_2155,In_2983);
nor U2217 (N_2217,In_633,N_1240);
nor U2218 (N_2218,N_1698,N_1781);
and U2219 (N_2219,N_1472,N_1523);
nor U2220 (N_2220,N_816,In_1946);
nor U2221 (N_2221,N_1242,N_1880);
nor U2222 (N_2222,In_1901,N_53);
and U2223 (N_2223,N_674,N_1346);
nor U2224 (N_2224,N_1514,N_225);
nand U2225 (N_2225,In_2901,N_1764);
or U2226 (N_2226,N_1084,N_1894);
nand U2227 (N_2227,N_1910,N_649);
nand U2228 (N_2228,N_1890,N_1624);
xnor U2229 (N_2229,N_1889,N_1752);
or U2230 (N_2230,N_1463,In_2216);
nand U2231 (N_2231,N_842,N_1534);
or U2232 (N_2232,N_573,N_1795);
xor U2233 (N_2233,N_232,In_1556);
and U2234 (N_2234,N_1553,N_1565);
nand U2235 (N_2235,N_1638,In_1150);
nor U2236 (N_2236,N_530,N_1831);
or U2237 (N_2237,In_1833,N_1558);
and U2238 (N_2238,In_2470,N_1689);
xnor U2239 (N_2239,N_987,N_1957);
or U2240 (N_2240,N_1926,N_1597);
and U2241 (N_2241,N_1223,N_1868);
nand U2242 (N_2242,N_1222,N_1608);
and U2243 (N_2243,N_1659,In_2795);
and U2244 (N_2244,N_1303,N_1815);
nor U2245 (N_2245,N_1274,N_1983);
nand U2246 (N_2246,N_1704,N_1437);
nand U2247 (N_2247,N_1724,N_1872);
nor U2248 (N_2248,N_1140,N_1616);
nor U2249 (N_2249,N_1320,N_1835);
nand U2250 (N_2250,N_1538,N_1231);
and U2251 (N_2251,N_1866,In_1839);
nor U2252 (N_2252,N_1401,N_1734);
and U2253 (N_2253,N_1621,N_1832);
nand U2254 (N_2254,N_1258,N_1913);
or U2255 (N_2255,N_1792,N_939);
nor U2256 (N_2256,N_1375,N_1887);
nand U2257 (N_2257,N_1626,N_1365);
or U2258 (N_2258,N_122,In_2187);
or U2259 (N_2259,N_1321,N_1922);
nor U2260 (N_2260,In_1840,In_1582);
nor U2261 (N_2261,N_1131,In_565);
or U2262 (N_2262,N_1757,N_1561);
nand U2263 (N_2263,N_1946,N_1762);
or U2264 (N_2264,N_1768,N_758);
xnor U2265 (N_2265,N_702,N_1176);
xor U2266 (N_2266,N_1448,N_1639);
nor U2267 (N_2267,N_1964,In_1651);
nor U2268 (N_2268,N_1886,N_354);
xnor U2269 (N_2269,N_1651,N_1099);
nand U2270 (N_2270,N_1610,N_1452);
xnor U2271 (N_2271,N_1581,In_896);
or U2272 (N_2272,In_2185,N_1706);
and U2273 (N_2273,In_1429,In_511);
xor U2274 (N_2274,N_1111,N_1071);
xnor U2275 (N_2275,N_1803,N_1255);
and U2276 (N_2276,N_1443,N_1510);
and U2277 (N_2277,In_1884,N_1986);
xor U2278 (N_2278,N_1993,N_782);
or U2279 (N_2279,N_100,N_1751);
nand U2280 (N_2280,N_1895,In_818);
and U2281 (N_2281,N_1631,In_2571);
and U2282 (N_2282,N_570,N_1592);
nor U2283 (N_2283,N_873,N_1928);
xnor U2284 (N_2284,N_1905,In_1262);
and U2285 (N_2285,N_1526,N_1824);
and U2286 (N_2286,In_2211,N_1609);
xor U2287 (N_2287,In_15,N_1171);
and U2288 (N_2288,N_1681,N_1633);
xnor U2289 (N_2289,N_1911,N_1814);
and U2290 (N_2290,N_1726,In_1892);
nor U2291 (N_2291,N_1936,N_1195);
xor U2292 (N_2292,N_1796,N_1047);
nand U2293 (N_2293,N_1571,N_1674);
nand U2294 (N_2294,In_286,N_1885);
nor U2295 (N_2295,N_1055,N_1839);
nor U2296 (N_2296,N_1238,N_1870);
nand U2297 (N_2297,N_1567,N_1775);
or U2298 (N_2298,In_2287,N_1519);
nor U2299 (N_2299,N_1372,N_1727);
nand U2300 (N_2300,N_1906,N_1517);
or U2301 (N_2301,N_230,In_1000);
or U2302 (N_2302,N_1817,N_1646);
xnor U2303 (N_2303,N_1995,N_1670);
and U2304 (N_2304,N_876,N_1411);
and U2305 (N_2305,N_1181,N_1551);
nor U2306 (N_2306,N_669,In_2822);
nand U2307 (N_2307,In_657,In_1750);
xor U2308 (N_2308,N_1254,N_1521);
nor U2309 (N_2309,N_1956,In_25);
or U2310 (N_2310,N_1860,N_1897);
or U2311 (N_2311,N_1040,N_1711);
xor U2312 (N_2312,N_1721,N_1733);
nor U2313 (N_2313,N_1425,N_1688);
nand U2314 (N_2314,N_1971,N_820);
nand U2315 (N_2315,N_1968,N_1921);
and U2316 (N_2316,N_1024,N_1777);
xor U2317 (N_2317,N_1059,In_2523);
or U2318 (N_2318,N_1970,N_794);
nand U2319 (N_2319,N_1800,N_1854);
nor U2320 (N_2320,N_1064,N_1362);
xnor U2321 (N_2321,N_1823,In_1018);
and U2322 (N_2322,In_614,N_665);
and U2323 (N_2323,In_2425,N_1954);
xor U2324 (N_2324,N_1524,N_1673);
xor U2325 (N_2325,N_1731,N_311);
nor U2326 (N_2326,N_1406,In_381);
xor U2327 (N_2327,N_1982,In_2518);
nand U2328 (N_2328,N_1749,N_1802);
nand U2329 (N_2329,N_1930,In_1861);
nor U2330 (N_2330,In_1253,In_646);
nand U2331 (N_2331,In_486,N_1947);
and U2332 (N_2332,N_1671,In_933);
nor U2333 (N_2333,N_1779,N_964);
nand U2334 (N_2334,N_1820,N_1531);
nor U2335 (N_2335,N_1782,N_1804);
and U2336 (N_2336,N_1842,N_1319);
xor U2337 (N_2337,N_1257,In_985);
nand U2338 (N_2338,N_1361,N_1981);
and U2339 (N_2339,N_1996,N_1846);
nand U2340 (N_2340,N_1154,N_1647);
and U2341 (N_2341,N_1773,N_1819);
nor U2342 (N_2342,In_889,N_1530);
and U2343 (N_2343,N_1984,In_1534);
and U2344 (N_2344,N_1277,N_1241);
xor U2345 (N_2345,N_1522,N_1692);
xnor U2346 (N_2346,N_1679,In_2612);
xor U2347 (N_2347,N_1122,N_1573);
nand U2348 (N_2348,N_1491,In_1487);
nor U2349 (N_2349,N_1166,In_1247);
xnor U2350 (N_2350,N_1725,N_1869);
nand U2351 (N_2351,N_1542,N_773);
or U2352 (N_2352,N_1966,N_1251);
or U2353 (N_2353,N_1329,N_1002);
and U2354 (N_2354,In_572,N_1799);
or U2355 (N_2355,N_1359,N_1026);
or U2356 (N_2356,In_2855,In_746);
nand U2357 (N_2357,N_1769,N_1188);
nor U2358 (N_2358,In_2848,N_1856);
nor U2359 (N_2359,N_927,N_1787);
xnor U2360 (N_2360,N_1430,N_1784);
and U2361 (N_2361,In_1860,In_1313);
or U2362 (N_2362,N_1719,N_1742);
xnor U2363 (N_2363,N_1636,N_1900);
xnor U2364 (N_2364,N_414,N_1012);
nor U2365 (N_2365,N_1847,N_1729);
nor U2366 (N_2366,N_1516,N_1978);
or U2367 (N_2367,N_1776,In_1055);
and U2368 (N_2368,N_1589,In_616);
nand U2369 (N_2369,N_1174,In_120);
nor U2370 (N_2370,N_1904,In_110);
or U2371 (N_2371,N_1923,In_2535);
xor U2372 (N_2372,N_1666,N_1326);
xnor U2373 (N_2373,In_302,N_1293);
nand U2374 (N_2374,N_1585,N_1797);
or U2375 (N_2375,N_1003,N_1935);
nor U2376 (N_2376,N_1541,In_2858);
nor U2377 (N_2377,N_1687,N_1741);
and U2378 (N_2378,N_1605,N_1226);
xnor U2379 (N_2379,N_1963,N_1888);
and U2380 (N_2380,N_141,N_1515);
nor U2381 (N_2381,N_572,N_1081);
xor U2382 (N_2382,In_1523,N_549);
or U2383 (N_2383,N_1027,N_1575);
or U2384 (N_2384,N_970,N_1744);
and U2385 (N_2385,N_1418,N_765);
xor U2386 (N_2386,N_1234,N_1378);
nor U2387 (N_2387,N_1278,N_1548);
and U2388 (N_2388,N_1280,In_713);
nor U2389 (N_2389,N_1596,N_1715);
nor U2390 (N_2390,N_1933,In_842);
nor U2391 (N_2391,N_417,N_946);
or U2392 (N_2392,In_2505,N_1540);
or U2393 (N_2393,N_1501,N_1607);
nand U2394 (N_2394,N_825,N_1563);
nand U2395 (N_2395,N_1821,In_2464);
xnor U2396 (N_2396,N_1187,N_1402);
and U2397 (N_2397,N_1652,N_1896);
xnor U2398 (N_2398,N_1728,N_1713);
nand U2399 (N_2399,N_1810,N_1229);
nand U2400 (N_2400,N_1852,N_1678);
nor U2401 (N_2401,N_895,In_1792);
nand U2402 (N_2402,N_1828,N_299);
nor U2403 (N_2403,N_1528,N_1871);
nand U2404 (N_2404,N_1590,N_1722);
nand U2405 (N_2405,In_2990,N_1703);
xnor U2406 (N_2406,N_1451,In_2717);
and U2407 (N_2407,N_578,In_442);
nor U2408 (N_2408,N_1785,N_1838);
nand U2409 (N_2409,N_456,N_1388);
and U2410 (N_2410,N_1967,N_1566);
or U2411 (N_2411,N_1075,N_1572);
or U2412 (N_2412,In_1844,N_1958);
xnor U2413 (N_2413,N_1920,In_2041);
or U2414 (N_2414,N_1972,N_1702);
or U2415 (N_2415,N_1440,N_1529);
nor U2416 (N_2416,N_1990,N_1126);
nor U2417 (N_2417,N_1825,In_2802);
nand U2418 (N_2418,N_1883,N_1513);
xor U2419 (N_2419,N_1765,N_1950);
nand U2420 (N_2420,N_1667,N_1758);
and U2421 (N_2421,N_404,N_1753);
or U2422 (N_2422,N_1850,N_1915);
xor U2423 (N_2423,N_1584,N_1546);
or U2424 (N_2424,In_132,N_1899);
xor U2425 (N_2425,N_1588,N_1746);
or U2426 (N_2426,In_514,N_1932);
nand U2427 (N_2427,In_1790,N_1190);
or U2428 (N_2428,N_1184,N_1881);
nor U2429 (N_2429,In_1549,N_1619);
and U2430 (N_2430,N_1680,In_1763);
or U2431 (N_2431,In_378,In_1367);
nand U2432 (N_2432,N_1816,N_1076);
or U2433 (N_2433,N_1532,N_1600);
and U2434 (N_2434,N_1723,In_1038);
nor U2435 (N_2435,N_1604,N_1512);
xnor U2436 (N_2436,N_1937,N_1449);
nand U2437 (N_2437,N_1545,N_1912);
nor U2438 (N_2438,N_1699,N_1735);
nand U2439 (N_2439,In_396,N_1714);
or U2440 (N_2440,N_284,N_1650);
nand U2441 (N_2441,In_1842,N_1844);
or U2442 (N_2442,N_747,N_1345);
nand U2443 (N_2443,N_1951,N_1682);
nor U2444 (N_2444,N_1809,N_1570);
or U2445 (N_2445,In_963,N_911);
nor U2446 (N_2446,N_1960,N_1618);
xor U2447 (N_2447,N_1635,N_1628);
nand U2448 (N_2448,N_1502,N_1144);
nor U2449 (N_2449,N_1789,N_1833);
and U2450 (N_2450,N_1643,N_1694);
or U2451 (N_2451,N_1564,N_1090);
or U2452 (N_2452,N_487,N_1413);
and U2453 (N_2453,N_616,N_1710);
nor U2454 (N_2454,N_29,In_1132);
nand U2455 (N_2455,N_1170,In_2077);
nor U2456 (N_2456,N_1253,N_427);
nand U2457 (N_2457,N_1879,N_1893);
nand U2458 (N_2458,N_1067,N_1916);
and U2459 (N_2459,In_1607,In_2404);
or U2460 (N_2460,In_1735,N_1431);
nand U2461 (N_2461,N_1101,N_1557);
nor U2462 (N_2462,N_645,N_1811);
or U2463 (N_2463,N_409,N_656);
xnor U2464 (N_2464,N_1974,N_1672);
nand U2465 (N_2465,In_2844,N_550);
nor U2466 (N_2466,N_393,N_1091);
and U2467 (N_2467,N_1552,N_1771);
nand U2468 (N_2468,N_1641,N_1898);
or U2469 (N_2469,N_807,N_1857);
xnor U2470 (N_2470,In_37,N_1662);
xor U2471 (N_2471,N_1941,N_1582);
nand U2472 (N_2472,In_583,N_628);
nand U2473 (N_2473,N_1656,In_2949);
xnor U2474 (N_2474,N_1193,In_542);
nand U2475 (N_2475,N_1005,N_871);
and U2476 (N_2476,In_2411,N_1500);
and U2477 (N_2477,In_2913,N_1788);
or U2478 (N_2478,N_815,N_1927);
and U2479 (N_2479,N_1158,N_1606);
and U2480 (N_2480,N_1390,N_1479);
nor U2481 (N_2481,In_1286,N_1535);
and U2482 (N_2482,N_1202,N_1924);
or U2483 (N_2483,In_1254,N_1841);
xor U2484 (N_2484,In_945,N_1849);
and U2485 (N_2485,N_1533,In_2856);
and U2486 (N_2486,In_536,N_1100);
xor U2487 (N_2487,N_1748,In_1458);
and U2488 (N_2488,N_1812,In_591);
or U2489 (N_2489,N_1909,N_1991);
nand U2490 (N_2490,N_155,In_1774);
and U2491 (N_2491,N_1113,N_1830);
or U2492 (N_2492,In_1692,N_1708);
nand U2493 (N_2493,N_1640,N_246);
and U2494 (N_2494,N_1299,N_380);
xnor U2495 (N_2495,N_192,N_1509);
nand U2496 (N_2496,N_1614,N_1791);
nor U2497 (N_2497,In_1776,In_525);
or U2498 (N_2498,N_60,In_2479);
xor U2499 (N_2499,N_55,N_1716);
nor U2500 (N_2500,N_2400,N_2441);
nand U2501 (N_2501,N_2172,N_2287);
nor U2502 (N_2502,N_2075,N_2464);
or U2503 (N_2503,N_2164,N_2371);
nor U2504 (N_2504,N_2459,N_2025);
nor U2505 (N_2505,N_2000,N_2083);
xnor U2506 (N_2506,N_2357,N_2012);
xor U2507 (N_2507,N_2184,N_2079);
and U2508 (N_2508,N_2261,N_2349);
or U2509 (N_2509,N_2159,N_2355);
and U2510 (N_2510,N_2238,N_2390);
nand U2511 (N_2511,N_2448,N_2145);
or U2512 (N_2512,N_2253,N_2340);
and U2513 (N_2513,N_2466,N_2150);
nor U2514 (N_2514,N_2486,N_2136);
and U2515 (N_2515,N_2035,N_2498);
and U2516 (N_2516,N_2382,N_2343);
nor U2517 (N_2517,N_2208,N_2101);
nor U2518 (N_2518,N_2258,N_2140);
nor U2519 (N_2519,N_2060,N_2338);
and U2520 (N_2520,N_2137,N_2076);
nand U2521 (N_2521,N_2367,N_2142);
nand U2522 (N_2522,N_2389,N_2011);
and U2523 (N_2523,N_2353,N_2452);
nand U2524 (N_2524,N_2018,N_2255);
and U2525 (N_2525,N_2002,N_2308);
and U2526 (N_2526,N_2201,N_2458);
or U2527 (N_2527,N_2420,N_2050);
nor U2528 (N_2528,N_2369,N_2176);
nor U2529 (N_2529,N_2005,N_2028);
and U2530 (N_2530,N_2288,N_2320);
xnor U2531 (N_2531,N_2364,N_2386);
nor U2532 (N_2532,N_2190,N_2213);
or U2533 (N_2533,N_2268,N_2451);
and U2534 (N_2534,N_2051,N_2312);
or U2535 (N_2535,N_2203,N_2211);
xor U2536 (N_2536,N_2148,N_2395);
and U2537 (N_2537,N_2071,N_2405);
and U2538 (N_2538,N_2331,N_2026);
and U2539 (N_2539,N_2197,N_2327);
or U2540 (N_2540,N_2476,N_2455);
and U2541 (N_2541,N_2059,N_2038);
and U2542 (N_2542,N_2483,N_2216);
xnor U2543 (N_2543,N_2198,N_2354);
xnor U2544 (N_2544,N_2068,N_2157);
nand U2545 (N_2545,N_2438,N_2110);
xor U2546 (N_2546,N_2422,N_2300);
or U2547 (N_2547,N_2127,N_2014);
or U2548 (N_2548,N_2251,N_2162);
nand U2549 (N_2549,N_2392,N_2381);
nand U2550 (N_2550,N_2099,N_2315);
nor U2551 (N_2551,N_2131,N_2105);
xor U2552 (N_2552,N_2094,N_2022);
xor U2553 (N_2553,N_2385,N_2450);
nor U2554 (N_2554,N_2348,N_2040);
nor U2555 (N_2555,N_2352,N_2016);
nor U2556 (N_2556,N_2301,N_2309);
nand U2557 (N_2557,N_2388,N_2158);
nand U2558 (N_2558,N_2092,N_2477);
and U2559 (N_2559,N_2256,N_2096);
and U2560 (N_2560,N_2319,N_2478);
and U2561 (N_2561,N_2491,N_2036);
nor U2562 (N_2562,N_2174,N_2363);
nor U2563 (N_2563,N_2270,N_2493);
xnor U2564 (N_2564,N_2154,N_2324);
nand U2565 (N_2565,N_2200,N_2454);
nor U2566 (N_2566,N_2437,N_2134);
and U2567 (N_2567,N_2103,N_2244);
and U2568 (N_2568,N_2228,N_2274);
nand U2569 (N_2569,N_2078,N_2045);
and U2570 (N_2570,N_2304,N_2419);
and U2571 (N_2571,N_2032,N_2209);
xor U2572 (N_2572,N_2084,N_2100);
nor U2573 (N_2573,N_2297,N_2229);
xnor U2574 (N_2574,N_2104,N_2088);
xor U2575 (N_2575,N_2008,N_2226);
nor U2576 (N_2576,N_2168,N_2425);
xnor U2577 (N_2577,N_2281,N_2398);
or U2578 (N_2578,N_2368,N_2116);
nor U2579 (N_2579,N_2171,N_2433);
or U2580 (N_2580,N_2144,N_2043);
nor U2581 (N_2581,N_2254,N_2219);
xnor U2582 (N_2582,N_2298,N_2163);
nor U2583 (N_2583,N_2399,N_2492);
and U2584 (N_2584,N_2202,N_2414);
nor U2585 (N_2585,N_2418,N_2463);
and U2586 (N_2586,N_2417,N_2410);
nand U2587 (N_2587,N_2462,N_2409);
nand U2588 (N_2588,N_2241,N_2047);
and U2589 (N_2589,N_2387,N_2443);
xnor U2590 (N_2590,N_2471,N_2264);
nor U2591 (N_2591,N_2378,N_2436);
and U2592 (N_2592,N_2021,N_2423);
xor U2593 (N_2593,N_2210,N_2191);
nor U2594 (N_2594,N_2033,N_2293);
xnor U2595 (N_2595,N_2024,N_2081);
and U2596 (N_2596,N_2372,N_2095);
nor U2597 (N_2597,N_2236,N_2231);
or U2598 (N_2598,N_2063,N_2487);
or U2599 (N_2599,N_2117,N_2266);
xor U2600 (N_2600,N_2342,N_2020);
nand U2601 (N_2601,N_2182,N_2499);
and U2602 (N_2602,N_2339,N_2166);
nor U2603 (N_2603,N_2130,N_2265);
or U2604 (N_2604,N_2453,N_2013);
xnor U2605 (N_2605,N_2126,N_2004);
nand U2606 (N_2606,N_2447,N_2461);
xnor U2607 (N_2607,N_2376,N_2321);
and U2608 (N_2608,N_2046,N_2027);
and U2609 (N_2609,N_2082,N_2192);
or U2610 (N_2610,N_2360,N_2102);
nand U2611 (N_2611,N_2058,N_2223);
or U2612 (N_2612,N_2235,N_2085);
and U2613 (N_2613,N_2207,N_2222);
xor U2614 (N_2614,N_2054,N_2179);
xor U2615 (N_2615,N_2359,N_2034);
nor U2616 (N_2616,N_2122,N_2053);
nand U2617 (N_2617,N_2183,N_2001);
nor U2618 (N_2618,N_2175,N_2052);
or U2619 (N_2619,N_2193,N_2344);
or U2620 (N_2620,N_2449,N_2139);
and U2621 (N_2621,N_2429,N_2073);
and U2622 (N_2622,N_2296,N_2432);
xnor U2623 (N_2623,N_2243,N_2276);
or U2624 (N_2624,N_2457,N_2278);
and U2625 (N_2625,N_2484,N_2430);
nand U2626 (N_2626,N_2039,N_2233);
and U2627 (N_2627,N_2080,N_2494);
nor U2628 (N_2628,N_2488,N_2056);
xnor U2629 (N_2629,N_2273,N_2257);
and U2630 (N_2630,N_2347,N_2291);
and U2631 (N_2631,N_2467,N_2497);
or U2632 (N_2632,N_2442,N_2470);
and U2633 (N_2633,N_2093,N_2440);
nand U2634 (N_2634,N_2106,N_2397);
xor U2635 (N_2635,N_2125,N_2181);
or U2636 (N_2636,N_2472,N_2377);
xnor U2637 (N_2637,N_2220,N_2177);
nand U2638 (N_2638,N_2087,N_2234);
xnor U2639 (N_2639,N_2048,N_2062);
and U2640 (N_2640,N_2187,N_2224);
nand U2641 (N_2641,N_2275,N_2240);
and U2642 (N_2642,N_2318,N_2394);
nand U2643 (N_2643,N_2350,N_2070);
xor U2644 (N_2644,N_2481,N_2407);
or U2645 (N_2645,N_2465,N_2129);
nor U2646 (N_2646,N_2269,N_2115);
or U2647 (N_2647,N_2124,N_2090);
or U2648 (N_2648,N_2042,N_2237);
xor U2649 (N_2649,N_2218,N_2061);
or U2650 (N_2650,N_2249,N_2416);
nand U2651 (N_2651,N_2285,N_2245);
or U2652 (N_2652,N_2260,N_2290);
nor U2653 (N_2653,N_2199,N_2474);
xnor U2654 (N_2654,N_2160,N_2023);
nor U2655 (N_2655,N_2188,N_2345);
nor U2656 (N_2656,N_2314,N_2393);
nor U2657 (N_2657,N_2325,N_2204);
xor U2658 (N_2658,N_2180,N_2495);
or U2659 (N_2659,N_2445,N_2185);
or U2660 (N_2660,N_2446,N_2311);
nor U2661 (N_2661,N_2310,N_2091);
or U2662 (N_2662,N_2468,N_2143);
and U2663 (N_2663,N_2456,N_2326);
nand U2664 (N_2664,N_2402,N_2307);
xnor U2665 (N_2665,N_2317,N_2316);
and U2666 (N_2666,N_2284,N_2138);
nand U2667 (N_2667,N_2313,N_2373);
xnor U2668 (N_2668,N_2109,N_2217);
xnor U2669 (N_2669,N_2151,N_2247);
or U2670 (N_2670,N_2206,N_2370);
and U2671 (N_2671,N_2375,N_2248);
or U2672 (N_2672,N_2282,N_2064);
and U2673 (N_2673,N_2194,N_2156);
xor U2674 (N_2674,N_2239,N_2279);
and U2675 (N_2675,N_2186,N_2286);
nor U2676 (N_2676,N_2411,N_2401);
and U2677 (N_2677,N_2074,N_2120);
nand U2678 (N_2678,N_2055,N_2406);
xor U2679 (N_2679,N_2169,N_2329);
and U2680 (N_2680,N_2173,N_2351);
or U2681 (N_2681,N_2098,N_2408);
nand U2682 (N_2682,N_2155,N_2132);
nor U2683 (N_2683,N_2412,N_2108);
nand U2684 (N_2684,N_2009,N_2112);
nand U2685 (N_2685,N_2067,N_2427);
and U2686 (N_2686,N_2232,N_2489);
or U2687 (N_2687,N_2336,N_2149);
nand U2688 (N_2688,N_2366,N_2029);
or U2689 (N_2689,N_2469,N_2121);
nor U2690 (N_2690,N_2230,N_2089);
and U2691 (N_2691,N_2242,N_2114);
xor U2692 (N_2692,N_2119,N_2413);
nor U2693 (N_2693,N_2272,N_2041);
and U2694 (N_2694,N_2069,N_2365);
nand U2695 (N_2695,N_2299,N_2017);
xnor U2696 (N_2696,N_2403,N_2271);
nand U2697 (N_2697,N_2111,N_2107);
nand U2698 (N_2698,N_2133,N_2333);
nor U2699 (N_2699,N_2170,N_2267);
and U2700 (N_2700,N_2379,N_2049);
nand U2701 (N_2701,N_2346,N_2019);
and U2702 (N_2702,N_2196,N_2252);
nand U2703 (N_2703,N_2031,N_2215);
and U2704 (N_2704,N_2482,N_2323);
and U2705 (N_2705,N_2227,N_2003);
nor U2706 (N_2706,N_2330,N_2421);
or U2707 (N_2707,N_2305,N_2262);
nor U2708 (N_2708,N_2010,N_2302);
nor U2709 (N_2709,N_2460,N_2259);
nor U2710 (N_2710,N_2167,N_2328);
xor U2711 (N_2711,N_2030,N_2221);
nor U2712 (N_2712,N_2303,N_2015);
nor U2713 (N_2713,N_2415,N_2306);
and U2714 (N_2714,N_2294,N_2341);
nor U2715 (N_2715,N_2295,N_2289);
xor U2716 (N_2716,N_2135,N_2374);
xnor U2717 (N_2717,N_2383,N_2485);
nand U2718 (N_2718,N_2384,N_2263);
xor U2719 (N_2719,N_2434,N_2391);
and U2720 (N_2720,N_2473,N_2292);
nand U2721 (N_2721,N_2189,N_2128);
xor U2722 (N_2722,N_2426,N_2057);
or U2723 (N_2723,N_2146,N_2214);
nand U2724 (N_2724,N_2225,N_2044);
and U2725 (N_2725,N_2066,N_2152);
xor U2726 (N_2726,N_2332,N_2424);
xor U2727 (N_2727,N_2358,N_2212);
nand U2728 (N_2728,N_2475,N_2428);
xor U2729 (N_2729,N_2006,N_2147);
nand U2730 (N_2730,N_2123,N_2195);
nand U2731 (N_2731,N_2283,N_2250);
nor U2732 (N_2732,N_2178,N_2037);
nor U2733 (N_2733,N_2334,N_2165);
nand U2734 (N_2734,N_2007,N_2356);
or U2735 (N_2735,N_2161,N_2337);
nand U2736 (N_2736,N_2439,N_2380);
nor U2737 (N_2737,N_2479,N_2431);
xnor U2738 (N_2738,N_2153,N_2113);
or U2739 (N_2739,N_2404,N_2362);
xor U2740 (N_2740,N_2141,N_2496);
and U2741 (N_2741,N_2490,N_2246);
xor U2742 (N_2742,N_2077,N_2065);
and U2743 (N_2743,N_2118,N_2205);
xnor U2744 (N_2744,N_2480,N_2280);
nor U2745 (N_2745,N_2444,N_2435);
xnor U2746 (N_2746,N_2072,N_2361);
nand U2747 (N_2747,N_2322,N_2335);
nor U2748 (N_2748,N_2277,N_2097);
and U2749 (N_2749,N_2396,N_2086);
nor U2750 (N_2750,N_2191,N_2355);
and U2751 (N_2751,N_2400,N_2396);
and U2752 (N_2752,N_2345,N_2372);
and U2753 (N_2753,N_2008,N_2062);
xnor U2754 (N_2754,N_2426,N_2006);
and U2755 (N_2755,N_2220,N_2003);
nand U2756 (N_2756,N_2268,N_2297);
nand U2757 (N_2757,N_2264,N_2464);
nor U2758 (N_2758,N_2337,N_2076);
and U2759 (N_2759,N_2153,N_2306);
and U2760 (N_2760,N_2071,N_2356);
nand U2761 (N_2761,N_2437,N_2096);
or U2762 (N_2762,N_2287,N_2111);
xnor U2763 (N_2763,N_2422,N_2344);
xor U2764 (N_2764,N_2030,N_2397);
nor U2765 (N_2765,N_2044,N_2068);
xor U2766 (N_2766,N_2329,N_2465);
nor U2767 (N_2767,N_2028,N_2038);
or U2768 (N_2768,N_2144,N_2114);
nand U2769 (N_2769,N_2033,N_2336);
nand U2770 (N_2770,N_2114,N_2338);
nand U2771 (N_2771,N_2115,N_2143);
nand U2772 (N_2772,N_2244,N_2141);
nand U2773 (N_2773,N_2370,N_2279);
nand U2774 (N_2774,N_2474,N_2117);
and U2775 (N_2775,N_2213,N_2299);
nand U2776 (N_2776,N_2159,N_2065);
nor U2777 (N_2777,N_2010,N_2202);
and U2778 (N_2778,N_2246,N_2248);
nand U2779 (N_2779,N_2440,N_2461);
nand U2780 (N_2780,N_2434,N_2239);
nor U2781 (N_2781,N_2241,N_2400);
xnor U2782 (N_2782,N_2161,N_2136);
and U2783 (N_2783,N_2144,N_2199);
nor U2784 (N_2784,N_2189,N_2476);
nand U2785 (N_2785,N_2046,N_2062);
nand U2786 (N_2786,N_2240,N_2121);
nor U2787 (N_2787,N_2245,N_2358);
nand U2788 (N_2788,N_2157,N_2352);
nand U2789 (N_2789,N_2385,N_2317);
and U2790 (N_2790,N_2279,N_2080);
xnor U2791 (N_2791,N_2180,N_2311);
nand U2792 (N_2792,N_2495,N_2225);
nand U2793 (N_2793,N_2444,N_2427);
nor U2794 (N_2794,N_2326,N_2478);
nand U2795 (N_2795,N_2364,N_2392);
nor U2796 (N_2796,N_2274,N_2176);
or U2797 (N_2797,N_2269,N_2336);
or U2798 (N_2798,N_2342,N_2261);
nand U2799 (N_2799,N_2099,N_2201);
or U2800 (N_2800,N_2002,N_2393);
nand U2801 (N_2801,N_2170,N_2469);
xor U2802 (N_2802,N_2294,N_2274);
nand U2803 (N_2803,N_2391,N_2009);
xor U2804 (N_2804,N_2303,N_2307);
nand U2805 (N_2805,N_2012,N_2013);
nand U2806 (N_2806,N_2356,N_2433);
nand U2807 (N_2807,N_2466,N_2452);
or U2808 (N_2808,N_2497,N_2101);
or U2809 (N_2809,N_2121,N_2082);
or U2810 (N_2810,N_2333,N_2469);
nor U2811 (N_2811,N_2083,N_2123);
nand U2812 (N_2812,N_2380,N_2133);
xnor U2813 (N_2813,N_2304,N_2003);
or U2814 (N_2814,N_2459,N_2374);
and U2815 (N_2815,N_2309,N_2312);
xnor U2816 (N_2816,N_2484,N_2155);
nor U2817 (N_2817,N_2460,N_2316);
xor U2818 (N_2818,N_2087,N_2026);
nor U2819 (N_2819,N_2023,N_2060);
and U2820 (N_2820,N_2166,N_2096);
nand U2821 (N_2821,N_2377,N_2422);
nor U2822 (N_2822,N_2185,N_2466);
xnor U2823 (N_2823,N_2123,N_2058);
nand U2824 (N_2824,N_2370,N_2303);
nor U2825 (N_2825,N_2499,N_2387);
or U2826 (N_2826,N_2240,N_2378);
or U2827 (N_2827,N_2198,N_2106);
xnor U2828 (N_2828,N_2245,N_2257);
xor U2829 (N_2829,N_2447,N_2451);
nand U2830 (N_2830,N_2166,N_2477);
or U2831 (N_2831,N_2006,N_2243);
xor U2832 (N_2832,N_2226,N_2039);
or U2833 (N_2833,N_2292,N_2000);
xor U2834 (N_2834,N_2247,N_2257);
or U2835 (N_2835,N_2284,N_2170);
nor U2836 (N_2836,N_2038,N_2342);
xnor U2837 (N_2837,N_2356,N_2082);
or U2838 (N_2838,N_2141,N_2316);
nor U2839 (N_2839,N_2182,N_2060);
xnor U2840 (N_2840,N_2053,N_2471);
and U2841 (N_2841,N_2311,N_2232);
nor U2842 (N_2842,N_2454,N_2245);
nor U2843 (N_2843,N_2322,N_2165);
and U2844 (N_2844,N_2006,N_2094);
nor U2845 (N_2845,N_2483,N_2381);
and U2846 (N_2846,N_2394,N_2465);
nand U2847 (N_2847,N_2141,N_2295);
nand U2848 (N_2848,N_2314,N_2341);
or U2849 (N_2849,N_2226,N_2079);
nor U2850 (N_2850,N_2016,N_2174);
nor U2851 (N_2851,N_2370,N_2041);
or U2852 (N_2852,N_2044,N_2366);
xnor U2853 (N_2853,N_2106,N_2388);
nor U2854 (N_2854,N_2367,N_2125);
or U2855 (N_2855,N_2449,N_2029);
xnor U2856 (N_2856,N_2046,N_2373);
xnor U2857 (N_2857,N_2001,N_2188);
or U2858 (N_2858,N_2261,N_2462);
nor U2859 (N_2859,N_2488,N_2072);
and U2860 (N_2860,N_2443,N_2333);
or U2861 (N_2861,N_2243,N_2223);
and U2862 (N_2862,N_2412,N_2106);
or U2863 (N_2863,N_2057,N_2132);
and U2864 (N_2864,N_2235,N_2219);
or U2865 (N_2865,N_2440,N_2495);
or U2866 (N_2866,N_2381,N_2350);
or U2867 (N_2867,N_2343,N_2208);
or U2868 (N_2868,N_2390,N_2174);
and U2869 (N_2869,N_2224,N_2382);
and U2870 (N_2870,N_2032,N_2010);
nor U2871 (N_2871,N_2212,N_2440);
nor U2872 (N_2872,N_2435,N_2068);
xnor U2873 (N_2873,N_2436,N_2160);
or U2874 (N_2874,N_2309,N_2264);
nand U2875 (N_2875,N_2434,N_2358);
xnor U2876 (N_2876,N_2233,N_2099);
nand U2877 (N_2877,N_2379,N_2102);
nor U2878 (N_2878,N_2357,N_2214);
and U2879 (N_2879,N_2078,N_2039);
or U2880 (N_2880,N_2435,N_2410);
nand U2881 (N_2881,N_2402,N_2142);
or U2882 (N_2882,N_2208,N_2037);
nor U2883 (N_2883,N_2297,N_2493);
and U2884 (N_2884,N_2395,N_2463);
nand U2885 (N_2885,N_2178,N_2124);
nand U2886 (N_2886,N_2143,N_2394);
or U2887 (N_2887,N_2121,N_2052);
xnor U2888 (N_2888,N_2299,N_2263);
and U2889 (N_2889,N_2285,N_2222);
or U2890 (N_2890,N_2215,N_2484);
or U2891 (N_2891,N_2341,N_2410);
and U2892 (N_2892,N_2426,N_2193);
xnor U2893 (N_2893,N_2359,N_2050);
nor U2894 (N_2894,N_2009,N_2288);
or U2895 (N_2895,N_2043,N_2411);
nor U2896 (N_2896,N_2256,N_2161);
and U2897 (N_2897,N_2485,N_2189);
nor U2898 (N_2898,N_2218,N_2157);
or U2899 (N_2899,N_2065,N_2022);
or U2900 (N_2900,N_2299,N_2175);
nor U2901 (N_2901,N_2463,N_2186);
nor U2902 (N_2902,N_2074,N_2050);
or U2903 (N_2903,N_2234,N_2085);
nor U2904 (N_2904,N_2323,N_2438);
nand U2905 (N_2905,N_2007,N_2205);
and U2906 (N_2906,N_2465,N_2117);
nor U2907 (N_2907,N_2065,N_2455);
or U2908 (N_2908,N_2101,N_2148);
or U2909 (N_2909,N_2135,N_2392);
or U2910 (N_2910,N_2224,N_2284);
and U2911 (N_2911,N_2443,N_2151);
nor U2912 (N_2912,N_2488,N_2362);
and U2913 (N_2913,N_2431,N_2131);
xor U2914 (N_2914,N_2266,N_2210);
nand U2915 (N_2915,N_2030,N_2304);
nand U2916 (N_2916,N_2498,N_2419);
nand U2917 (N_2917,N_2311,N_2275);
or U2918 (N_2918,N_2057,N_2363);
nor U2919 (N_2919,N_2326,N_2182);
xnor U2920 (N_2920,N_2043,N_2075);
nor U2921 (N_2921,N_2152,N_2068);
xor U2922 (N_2922,N_2125,N_2172);
and U2923 (N_2923,N_2410,N_2095);
and U2924 (N_2924,N_2101,N_2068);
nor U2925 (N_2925,N_2167,N_2193);
nor U2926 (N_2926,N_2226,N_2383);
or U2927 (N_2927,N_2434,N_2232);
nand U2928 (N_2928,N_2435,N_2069);
nand U2929 (N_2929,N_2328,N_2338);
or U2930 (N_2930,N_2284,N_2155);
or U2931 (N_2931,N_2226,N_2472);
nor U2932 (N_2932,N_2189,N_2302);
and U2933 (N_2933,N_2346,N_2335);
xnor U2934 (N_2934,N_2453,N_2049);
xor U2935 (N_2935,N_2300,N_2255);
xor U2936 (N_2936,N_2118,N_2404);
and U2937 (N_2937,N_2300,N_2332);
nor U2938 (N_2938,N_2113,N_2143);
nor U2939 (N_2939,N_2183,N_2156);
and U2940 (N_2940,N_2301,N_2079);
and U2941 (N_2941,N_2244,N_2006);
nand U2942 (N_2942,N_2164,N_2187);
nor U2943 (N_2943,N_2023,N_2361);
nor U2944 (N_2944,N_2191,N_2206);
xnor U2945 (N_2945,N_2259,N_2385);
or U2946 (N_2946,N_2316,N_2136);
nand U2947 (N_2947,N_2228,N_2258);
and U2948 (N_2948,N_2318,N_2184);
and U2949 (N_2949,N_2212,N_2382);
xor U2950 (N_2950,N_2202,N_2312);
xnor U2951 (N_2951,N_2084,N_2306);
or U2952 (N_2952,N_2391,N_2260);
and U2953 (N_2953,N_2381,N_2147);
or U2954 (N_2954,N_2497,N_2351);
or U2955 (N_2955,N_2258,N_2495);
nand U2956 (N_2956,N_2479,N_2350);
nor U2957 (N_2957,N_2253,N_2396);
xor U2958 (N_2958,N_2272,N_2021);
nand U2959 (N_2959,N_2415,N_2429);
nand U2960 (N_2960,N_2448,N_2328);
and U2961 (N_2961,N_2454,N_2386);
xor U2962 (N_2962,N_2259,N_2473);
nor U2963 (N_2963,N_2209,N_2077);
nor U2964 (N_2964,N_2491,N_2271);
and U2965 (N_2965,N_2387,N_2454);
or U2966 (N_2966,N_2273,N_2070);
nor U2967 (N_2967,N_2388,N_2320);
nand U2968 (N_2968,N_2419,N_2200);
xnor U2969 (N_2969,N_2000,N_2285);
or U2970 (N_2970,N_2130,N_2085);
xor U2971 (N_2971,N_2213,N_2095);
or U2972 (N_2972,N_2333,N_2208);
or U2973 (N_2973,N_2077,N_2251);
and U2974 (N_2974,N_2467,N_2358);
or U2975 (N_2975,N_2107,N_2391);
nor U2976 (N_2976,N_2108,N_2168);
nand U2977 (N_2977,N_2125,N_2136);
or U2978 (N_2978,N_2320,N_2062);
and U2979 (N_2979,N_2355,N_2291);
and U2980 (N_2980,N_2193,N_2413);
xor U2981 (N_2981,N_2131,N_2090);
xnor U2982 (N_2982,N_2118,N_2432);
or U2983 (N_2983,N_2107,N_2145);
xor U2984 (N_2984,N_2193,N_2488);
xor U2985 (N_2985,N_2360,N_2239);
and U2986 (N_2986,N_2321,N_2387);
nor U2987 (N_2987,N_2474,N_2169);
nor U2988 (N_2988,N_2402,N_2458);
nor U2989 (N_2989,N_2493,N_2424);
xor U2990 (N_2990,N_2183,N_2056);
and U2991 (N_2991,N_2481,N_2367);
nand U2992 (N_2992,N_2007,N_2442);
and U2993 (N_2993,N_2175,N_2061);
xnor U2994 (N_2994,N_2205,N_2474);
and U2995 (N_2995,N_2345,N_2133);
and U2996 (N_2996,N_2375,N_2431);
xnor U2997 (N_2997,N_2453,N_2057);
xor U2998 (N_2998,N_2463,N_2492);
xor U2999 (N_2999,N_2015,N_2282);
nand U3000 (N_3000,N_2567,N_2586);
or U3001 (N_3001,N_2903,N_2651);
nor U3002 (N_3002,N_2845,N_2604);
xor U3003 (N_3003,N_2791,N_2956);
nor U3004 (N_3004,N_2983,N_2659);
or U3005 (N_3005,N_2821,N_2838);
xnor U3006 (N_3006,N_2554,N_2697);
nand U3007 (N_3007,N_2787,N_2891);
and U3008 (N_3008,N_2633,N_2518);
or U3009 (N_3009,N_2915,N_2966);
nand U3010 (N_3010,N_2827,N_2943);
xor U3011 (N_3011,N_2835,N_2779);
and U3012 (N_3012,N_2816,N_2857);
nor U3013 (N_3013,N_2847,N_2799);
nor U3014 (N_3014,N_2675,N_2951);
or U3015 (N_3015,N_2877,N_2579);
or U3016 (N_3016,N_2905,N_2707);
or U3017 (N_3017,N_2866,N_2907);
xor U3018 (N_3018,N_2686,N_2679);
nor U3019 (N_3019,N_2617,N_2597);
or U3020 (N_3020,N_2513,N_2657);
nor U3021 (N_3021,N_2591,N_2912);
nor U3022 (N_3022,N_2739,N_2806);
or U3023 (N_3023,N_2771,N_2998);
nor U3024 (N_3024,N_2761,N_2802);
and U3025 (N_3025,N_2742,N_2927);
nor U3026 (N_3026,N_2616,N_2911);
and U3027 (N_3027,N_2996,N_2812);
or U3028 (N_3028,N_2517,N_2605);
nand U3029 (N_3029,N_2904,N_2972);
nand U3030 (N_3030,N_2696,N_2590);
and U3031 (N_3031,N_2886,N_2741);
or U3032 (N_3032,N_2815,N_2797);
nor U3033 (N_3033,N_2995,N_2618);
nor U3034 (N_3034,N_2786,N_2602);
nor U3035 (N_3035,N_2833,N_2843);
nor U3036 (N_3036,N_2701,N_2755);
nand U3037 (N_3037,N_2546,N_2710);
nand U3038 (N_3038,N_2563,N_2778);
and U3039 (N_3039,N_2773,N_2814);
nor U3040 (N_3040,N_2576,N_2603);
nand U3041 (N_3041,N_2528,N_2846);
nand U3042 (N_3042,N_2676,N_2527);
nor U3043 (N_3043,N_2746,N_2980);
nor U3044 (N_3044,N_2543,N_2990);
or U3045 (N_3045,N_2977,N_2844);
xor U3046 (N_3046,N_2716,N_2861);
or U3047 (N_3047,N_2937,N_2705);
or U3048 (N_3048,N_2685,N_2934);
or U3049 (N_3049,N_2794,N_2561);
nand U3050 (N_3050,N_2982,N_2627);
nor U3051 (N_3051,N_2639,N_2539);
nor U3052 (N_3052,N_2783,N_2774);
and U3053 (N_3053,N_2785,N_2569);
or U3054 (N_3054,N_2993,N_2665);
or U3055 (N_3055,N_2764,N_2643);
nand U3056 (N_3056,N_2926,N_2737);
nor U3057 (N_3057,N_2889,N_2708);
and U3058 (N_3058,N_2624,N_2621);
nor U3059 (N_3059,N_2818,N_2535);
nand U3060 (N_3060,N_2540,N_2673);
nor U3061 (N_3061,N_2671,N_2735);
and U3062 (N_3062,N_2628,N_2867);
nand U3063 (N_3063,N_2669,N_2693);
and U3064 (N_3064,N_2813,N_2558);
or U3065 (N_3065,N_2792,N_2524);
xnor U3066 (N_3066,N_2890,N_2704);
xnor U3067 (N_3067,N_2747,N_2900);
nor U3068 (N_3068,N_2876,N_2992);
or U3069 (N_3069,N_2512,N_2531);
or U3070 (N_3070,N_2544,N_2978);
nand U3071 (N_3071,N_2578,N_2928);
nand U3072 (N_3072,N_2840,N_2551);
xor U3073 (N_3073,N_2803,N_2655);
and U3074 (N_3074,N_2690,N_2830);
and U3075 (N_3075,N_2500,N_2714);
xnor U3076 (N_3076,N_2706,N_2784);
or U3077 (N_3077,N_2650,N_2975);
nor U3078 (N_3078,N_2506,N_2553);
xor U3079 (N_3079,N_2820,N_2849);
nor U3080 (N_3080,N_2589,N_2932);
xnor U3081 (N_3081,N_2807,N_2880);
nor U3082 (N_3082,N_2793,N_2511);
nor U3083 (N_3083,N_2729,N_2939);
or U3084 (N_3084,N_2896,N_2950);
xor U3085 (N_3085,N_2647,N_2678);
xor U3086 (N_3086,N_2908,N_2788);
nand U3087 (N_3087,N_2985,N_2585);
or U3088 (N_3088,N_2879,N_2727);
nor U3089 (N_3089,N_2858,N_2573);
or U3090 (N_3090,N_2749,N_2895);
and U3091 (N_3091,N_2836,N_2970);
or U3092 (N_3092,N_2981,N_2930);
and U3093 (N_3093,N_2622,N_2887);
or U3094 (N_3094,N_2526,N_2947);
nor U3095 (N_3095,N_2760,N_2949);
or U3096 (N_3096,N_2684,N_2522);
and U3097 (N_3097,N_2906,N_2984);
nor U3098 (N_3098,N_2571,N_2775);
nand U3099 (N_3099,N_2552,N_2831);
or U3100 (N_3100,N_2560,N_2922);
or U3101 (N_3101,N_2635,N_2945);
nand U3102 (N_3102,N_2881,N_2557);
nand U3103 (N_3103,N_2766,N_2822);
nor U3104 (N_3104,N_2712,N_2600);
xor U3105 (N_3105,N_2682,N_2940);
xor U3106 (N_3106,N_2948,N_2859);
nor U3107 (N_3107,N_2999,N_2958);
or U3108 (N_3108,N_2968,N_2960);
nor U3109 (N_3109,N_2864,N_2523);
nor U3110 (N_3110,N_2645,N_2798);
xor U3111 (N_3111,N_2751,N_2709);
or U3112 (N_3112,N_2961,N_2566);
xor U3113 (N_3113,N_2612,N_2962);
and U3114 (N_3114,N_2965,N_2620);
or U3115 (N_3115,N_2568,N_2629);
xor U3116 (N_3116,N_2899,N_2933);
xor U3117 (N_3117,N_2888,N_2574);
nor U3118 (N_3118,N_2801,N_2795);
nor U3119 (N_3119,N_2711,N_2893);
nand U3120 (N_3120,N_2583,N_2593);
and U3121 (N_3121,N_2681,N_2507);
or U3122 (N_3122,N_2796,N_2575);
xnor U3123 (N_3123,N_2728,N_2997);
and U3124 (N_3124,N_2957,N_2687);
nor U3125 (N_3125,N_2763,N_2520);
nand U3126 (N_3126,N_2834,N_2863);
or U3127 (N_3127,N_2850,N_2658);
nor U3128 (N_3128,N_2594,N_2626);
nor U3129 (N_3129,N_2610,N_2611);
or U3130 (N_3130,N_2782,N_2752);
xor U3131 (N_3131,N_2614,N_2810);
nor U3132 (N_3132,N_2577,N_2545);
xor U3133 (N_3133,N_2854,N_2661);
nand U3134 (N_3134,N_2868,N_2514);
xor U3135 (N_3135,N_2919,N_2765);
and U3136 (N_3136,N_2653,N_2555);
nor U3137 (N_3137,N_2580,N_2525);
or U3138 (N_3138,N_2703,N_2757);
xor U3139 (N_3139,N_2852,N_2536);
nor U3140 (N_3140,N_2811,N_2971);
xnor U3141 (N_3141,N_2756,N_2641);
nand U3142 (N_3142,N_2663,N_2750);
and U3143 (N_3143,N_2884,N_2588);
nor U3144 (N_3144,N_2768,N_2601);
nor U3145 (N_3145,N_2666,N_2994);
nor U3146 (N_3146,N_2564,N_2636);
nor U3147 (N_3147,N_2963,N_2924);
nand U3148 (N_3148,N_2509,N_2664);
xor U3149 (N_3149,N_2855,N_2515);
or U3150 (N_3150,N_2776,N_2865);
or U3151 (N_3151,N_2640,N_2914);
xnor U3152 (N_3152,N_2936,N_2946);
nand U3153 (N_3153,N_2608,N_2829);
nor U3154 (N_3154,N_2670,N_2825);
nand U3155 (N_3155,N_2550,N_2606);
or U3156 (N_3156,N_2767,N_2800);
or U3157 (N_3157,N_2715,N_2929);
and U3158 (N_3158,N_2790,N_2758);
and U3159 (N_3159,N_2955,N_2953);
xor U3160 (N_3160,N_2689,N_2878);
nand U3161 (N_3161,N_2944,N_2780);
nor U3162 (N_3162,N_2702,N_2549);
or U3163 (N_3163,N_2516,N_2587);
or U3164 (N_3164,N_2691,N_2521);
xnor U3165 (N_3165,N_2632,N_2503);
xor U3166 (N_3166,N_2967,N_2519);
nor U3167 (N_3167,N_2826,N_2772);
and U3168 (N_3168,N_2959,N_2913);
and U3169 (N_3169,N_2988,N_2853);
nand U3170 (N_3170,N_2819,N_2832);
nor U3171 (N_3171,N_2630,N_2672);
or U3172 (N_3172,N_2808,N_2730);
nand U3173 (N_3173,N_2733,N_2916);
and U3174 (N_3174,N_2851,N_2942);
and U3175 (N_3175,N_2649,N_2860);
or U3176 (N_3176,N_2723,N_2894);
nand U3177 (N_3177,N_2724,N_2987);
nor U3178 (N_3178,N_2917,N_2824);
xor U3179 (N_3179,N_2738,N_2969);
nor U3180 (N_3180,N_2743,N_2921);
xor U3181 (N_3181,N_2631,N_2873);
nand U3182 (N_3182,N_2910,N_2648);
nand U3183 (N_3183,N_2609,N_2976);
nor U3184 (N_3184,N_2935,N_2762);
nand U3185 (N_3185,N_2582,N_2744);
nand U3186 (N_3186,N_2615,N_2581);
xor U3187 (N_3187,N_2722,N_2638);
xnor U3188 (N_3188,N_2902,N_2918);
nor U3189 (N_3189,N_2979,N_2570);
nand U3190 (N_3190,N_2748,N_2619);
and U3191 (N_3191,N_2599,N_2719);
xnor U3192 (N_3192,N_2923,N_2505);
and U3193 (N_3193,N_2870,N_2789);
or U3194 (N_3194,N_2547,N_2841);
nand U3195 (N_3195,N_2882,N_2726);
xor U3196 (N_3196,N_2607,N_2938);
or U3197 (N_3197,N_2885,N_2548);
and U3198 (N_3198,N_2694,N_2668);
xor U3199 (N_3199,N_2642,N_2740);
and U3200 (N_3200,N_2952,N_2637);
and U3201 (N_3201,N_2501,N_2872);
nand U3202 (N_3202,N_2925,N_2713);
xor U3203 (N_3203,N_2683,N_2596);
and U3204 (N_3204,N_2986,N_2754);
or U3205 (N_3205,N_2745,N_2532);
nand U3206 (N_3206,N_2504,N_2805);
nor U3207 (N_3207,N_2674,N_2804);
nor U3208 (N_3208,N_2646,N_2734);
xnor U3209 (N_3209,N_2856,N_2874);
nor U3210 (N_3210,N_2529,N_2909);
or U3211 (N_3211,N_2530,N_2989);
nor U3212 (N_3212,N_2718,N_2595);
or U3213 (N_3213,N_2538,N_2920);
and U3214 (N_3214,N_2897,N_2502);
nand U3215 (N_3215,N_2721,N_2901);
xor U3216 (N_3216,N_2839,N_2625);
xor U3217 (N_3217,N_2875,N_2680);
nor U3218 (N_3218,N_2781,N_2848);
and U3219 (N_3219,N_2660,N_2823);
and U3220 (N_3220,N_2510,N_2892);
and U3221 (N_3221,N_2828,N_2562);
nor U3222 (N_3222,N_2817,N_2656);
nand U3223 (N_3223,N_2898,N_2542);
and U3224 (N_3224,N_2598,N_2809);
or U3225 (N_3225,N_2753,N_2667);
or U3226 (N_3226,N_2654,N_2973);
nand U3227 (N_3227,N_2731,N_2964);
nand U3228 (N_3228,N_2623,N_2556);
nor U3229 (N_3229,N_2613,N_2559);
xnor U3230 (N_3230,N_2695,N_2634);
or U3231 (N_3231,N_2732,N_2584);
and U3232 (N_3232,N_2698,N_2770);
or U3233 (N_3233,N_2592,N_2508);
nand U3234 (N_3234,N_2662,N_2842);
xnor U3235 (N_3235,N_2769,N_2541);
xor U3236 (N_3236,N_2777,N_2677);
or U3237 (N_3237,N_2537,N_2869);
and U3238 (N_3238,N_2871,N_2565);
xor U3239 (N_3239,N_2991,N_2759);
nor U3240 (N_3240,N_2862,N_2717);
and U3241 (N_3241,N_2700,N_2725);
or U3242 (N_3242,N_2699,N_2688);
nand U3243 (N_3243,N_2954,N_2652);
nand U3244 (N_3244,N_2534,N_2533);
or U3245 (N_3245,N_2572,N_2692);
nor U3246 (N_3246,N_2720,N_2883);
xnor U3247 (N_3247,N_2837,N_2941);
nand U3248 (N_3248,N_2931,N_2974);
or U3249 (N_3249,N_2736,N_2644);
nand U3250 (N_3250,N_2538,N_2660);
xor U3251 (N_3251,N_2913,N_2549);
nand U3252 (N_3252,N_2707,N_2845);
nor U3253 (N_3253,N_2667,N_2812);
or U3254 (N_3254,N_2604,N_2989);
nand U3255 (N_3255,N_2761,N_2958);
xor U3256 (N_3256,N_2599,N_2948);
xor U3257 (N_3257,N_2657,N_2731);
xnor U3258 (N_3258,N_2613,N_2977);
nor U3259 (N_3259,N_2948,N_2696);
or U3260 (N_3260,N_2633,N_2818);
and U3261 (N_3261,N_2740,N_2617);
and U3262 (N_3262,N_2882,N_2679);
xnor U3263 (N_3263,N_2822,N_2801);
and U3264 (N_3264,N_2713,N_2656);
xnor U3265 (N_3265,N_2837,N_2549);
and U3266 (N_3266,N_2898,N_2849);
nor U3267 (N_3267,N_2824,N_2731);
and U3268 (N_3268,N_2661,N_2651);
xnor U3269 (N_3269,N_2578,N_2688);
nor U3270 (N_3270,N_2686,N_2580);
xor U3271 (N_3271,N_2950,N_2557);
nand U3272 (N_3272,N_2932,N_2798);
nor U3273 (N_3273,N_2656,N_2718);
xor U3274 (N_3274,N_2788,N_2867);
nor U3275 (N_3275,N_2510,N_2831);
nand U3276 (N_3276,N_2586,N_2559);
and U3277 (N_3277,N_2780,N_2954);
nor U3278 (N_3278,N_2519,N_2707);
and U3279 (N_3279,N_2928,N_2930);
nor U3280 (N_3280,N_2932,N_2831);
xnor U3281 (N_3281,N_2907,N_2773);
nor U3282 (N_3282,N_2816,N_2987);
nor U3283 (N_3283,N_2672,N_2877);
nor U3284 (N_3284,N_2865,N_2518);
xor U3285 (N_3285,N_2560,N_2817);
nor U3286 (N_3286,N_2776,N_2711);
nor U3287 (N_3287,N_2776,N_2891);
nand U3288 (N_3288,N_2579,N_2613);
nor U3289 (N_3289,N_2942,N_2571);
and U3290 (N_3290,N_2539,N_2850);
xor U3291 (N_3291,N_2704,N_2838);
and U3292 (N_3292,N_2514,N_2963);
nand U3293 (N_3293,N_2881,N_2772);
nand U3294 (N_3294,N_2507,N_2864);
xor U3295 (N_3295,N_2719,N_2840);
nand U3296 (N_3296,N_2560,N_2531);
nor U3297 (N_3297,N_2502,N_2553);
or U3298 (N_3298,N_2849,N_2852);
nor U3299 (N_3299,N_2917,N_2726);
nor U3300 (N_3300,N_2559,N_2845);
nor U3301 (N_3301,N_2976,N_2585);
nand U3302 (N_3302,N_2953,N_2539);
nor U3303 (N_3303,N_2756,N_2534);
nor U3304 (N_3304,N_2858,N_2684);
and U3305 (N_3305,N_2854,N_2990);
xor U3306 (N_3306,N_2671,N_2944);
and U3307 (N_3307,N_2628,N_2597);
nand U3308 (N_3308,N_2701,N_2518);
nand U3309 (N_3309,N_2646,N_2638);
or U3310 (N_3310,N_2941,N_2723);
nand U3311 (N_3311,N_2876,N_2771);
nor U3312 (N_3312,N_2581,N_2914);
and U3313 (N_3313,N_2680,N_2782);
or U3314 (N_3314,N_2643,N_2664);
and U3315 (N_3315,N_2633,N_2858);
xor U3316 (N_3316,N_2571,N_2972);
or U3317 (N_3317,N_2656,N_2824);
nor U3318 (N_3318,N_2609,N_2630);
or U3319 (N_3319,N_2584,N_2543);
and U3320 (N_3320,N_2685,N_2947);
xor U3321 (N_3321,N_2745,N_2695);
and U3322 (N_3322,N_2565,N_2750);
xnor U3323 (N_3323,N_2573,N_2505);
nor U3324 (N_3324,N_2960,N_2685);
and U3325 (N_3325,N_2677,N_2700);
and U3326 (N_3326,N_2932,N_2750);
nand U3327 (N_3327,N_2646,N_2794);
and U3328 (N_3328,N_2917,N_2548);
nand U3329 (N_3329,N_2596,N_2804);
nand U3330 (N_3330,N_2774,N_2568);
xnor U3331 (N_3331,N_2518,N_2914);
or U3332 (N_3332,N_2998,N_2848);
or U3333 (N_3333,N_2979,N_2634);
nor U3334 (N_3334,N_2761,N_2776);
nor U3335 (N_3335,N_2659,N_2607);
or U3336 (N_3336,N_2949,N_2950);
xor U3337 (N_3337,N_2728,N_2810);
and U3338 (N_3338,N_2714,N_2543);
nand U3339 (N_3339,N_2719,N_2956);
or U3340 (N_3340,N_2988,N_2527);
and U3341 (N_3341,N_2974,N_2685);
and U3342 (N_3342,N_2520,N_2900);
nand U3343 (N_3343,N_2917,N_2581);
xor U3344 (N_3344,N_2831,N_2828);
xor U3345 (N_3345,N_2918,N_2548);
xnor U3346 (N_3346,N_2560,N_2718);
xnor U3347 (N_3347,N_2870,N_2583);
xnor U3348 (N_3348,N_2929,N_2793);
or U3349 (N_3349,N_2795,N_2842);
or U3350 (N_3350,N_2816,N_2524);
xor U3351 (N_3351,N_2666,N_2990);
nor U3352 (N_3352,N_2752,N_2948);
and U3353 (N_3353,N_2926,N_2896);
xor U3354 (N_3354,N_2542,N_2782);
or U3355 (N_3355,N_2545,N_2967);
xor U3356 (N_3356,N_2734,N_2541);
nor U3357 (N_3357,N_2674,N_2618);
xor U3358 (N_3358,N_2617,N_2904);
or U3359 (N_3359,N_2546,N_2883);
xor U3360 (N_3360,N_2758,N_2713);
and U3361 (N_3361,N_2717,N_2875);
or U3362 (N_3362,N_2888,N_2909);
or U3363 (N_3363,N_2725,N_2688);
or U3364 (N_3364,N_2694,N_2863);
and U3365 (N_3365,N_2975,N_2529);
nor U3366 (N_3366,N_2881,N_2691);
and U3367 (N_3367,N_2613,N_2896);
xor U3368 (N_3368,N_2637,N_2540);
nor U3369 (N_3369,N_2840,N_2759);
nand U3370 (N_3370,N_2754,N_2954);
or U3371 (N_3371,N_2572,N_2521);
or U3372 (N_3372,N_2925,N_2578);
nor U3373 (N_3373,N_2824,N_2769);
xnor U3374 (N_3374,N_2823,N_2939);
xnor U3375 (N_3375,N_2918,N_2886);
or U3376 (N_3376,N_2689,N_2501);
nand U3377 (N_3377,N_2672,N_2928);
nor U3378 (N_3378,N_2968,N_2727);
or U3379 (N_3379,N_2777,N_2568);
xor U3380 (N_3380,N_2787,N_2742);
nand U3381 (N_3381,N_2859,N_2586);
or U3382 (N_3382,N_2979,N_2836);
or U3383 (N_3383,N_2948,N_2960);
nor U3384 (N_3384,N_2743,N_2864);
nand U3385 (N_3385,N_2549,N_2911);
nor U3386 (N_3386,N_2761,N_2678);
and U3387 (N_3387,N_2742,N_2650);
nand U3388 (N_3388,N_2662,N_2779);
and U3389 (N_3389,N_2610,N_2834);
or U3390 (N_3390,N_2705,N_2891);
nand U3391 (N_3391,N_2644,N_2773);
xnor U3392 (N_3392,N_2698,N_2750);
nor U3393 (N_3393,N_2848,N_2607);
xnor U3394 (N_3394,N_2921,N_2986);
nand U3395 (N_3395,N_2849,N_2665);
xnor U3396 (N_3396,N_2527,N_2834);
or U3397 (N_3397,N_2974,N_2684);
and U3398 (N_3398,N_2942,N_2727);
xnor U3399 (N_3399,N_2541,N_2807);
nand U3400 (N_3400,N_2811,N_2799);
nor U3401 (N_3401,N_2959,N_2861);
nor U3402 (N_3402,N_2917,N_2546);
xor U3403 (N_3403,N_2835,N_2944);
and U3404 (N_3404,N_2662,N_2704);
nand U3405 (N_3405,N_2611,N_2988);
nand U3406 (N_3406,N_2780,N_2869);
or U3407 (N_3407,N_2611,N_2742);
xnor U3408 (N_3408,N_2861,N_2628);
or U3409 (N_3409,N_2923,N_2591);
or U3410 (N_3410,N_2660,N_2706);
nand U3411 (N_3411,N_2762,N_2836);
xnor U3412 (N_3412,N_2606,N_2725);
nor U3413 (N_3413,N_2895,N_2949);
or U3414 (N_3414,N_2770,N_2607);
xor U3415 (N_3415,N_2768,N_2883);
or U3416 (N_3416,N_2627,N_2873);
and U3417 (N_3417,N_2654,N_2868);
and U3418 (N_3418,N_2947,N_2963);
nor U3419 (N_3419,N_2511,N_2796);
nand U3420 (N_3420,N_2852,N_2960);
and U3421 (N_3421,N_2557,N_2758);
nand U3422 (N_3422,N_2597,N_2973);
xnor U3423 (N_3423,N_2735,N_2951);
nand U3424 (N_3424,N_2797,N_2748);
nor U3425 (N_3425,N_2515,N_2743);
and U3426 (N_3426,N_2807,N_2993);
xnor U3427 (N_3427,N_2790,N_2895);
nand U3428 (N_3428,N_2911,N_2771);
nand U3429 (N_3429,N_2871,N_2806);
xnor U3430 (N_3430,N_2678,N_2662);
or U3431 (N_3431,N_2572,N_2992);
and U3432 (N_3432,N_2614,N_2634);
nand U3433 (N_3433,N_2631,N_2584);
xnor U3434 (N_3434,N_2878,N_2888);
and U3435 (N_3435,N_2788,N_2925);
nand U3436 (N_3436,N_2583,N_2758);
nor U3437 (N_3437,N_2853,N_2974);
nand U3438 (N_3438,N_2632,N_2671);
nor U3439 (N_3439,N_2857,N_2923);
or U3440 (N_3440,N_2722,N_2956);
nor U3441 (N_3441,N_2741,N_2627);
nor U3442 (N_3442,N_2704,N_2670);
xnor U3443 (N_3443,N_2740,N_2906);
nand U3444 (N_3444,N_2796,N_2923);
nand U3445 (N_3445,N_2768,N_2663);
or U3446 (N_3446,N_2527,N_2837);
or U3447 (N_3447,N_2890,N_2534);
xor U3448 (N_3448,N_2777,N_2659);
or U3449 (N_3449,N_2704,N_2888);
xnor U3450 (N_3450,N_2756,N_2645);
nor U3451 (N_3451,N_2945,N_2616);
nand U3452 (N_3452,N_2821,N_2518);
and U3453 (N_3453,N_2562,N_2952);
and U3454 (N_3454,N_2832,N_2697);
nand U3455 (N_3455,N_2665,N_2562);
and U3456 (N_3456,N_2786,N_2503);
or U3457 (N_3457,N_2536,N_2517);
and U3458 (N_3458,N_2828,N_2987);
nor U3459 (N_3459,N_2925,N_2500);
and U3460 (N_3460,N_2517,N_2703);
nand U3461 (N_3461,N_2883,N_2601);
nand U3462 (N_3462,N_2671,N_2710);
and U3463 (N_3463,N_2986,N_2911);
nand U3464 (N_3464,N_2955,N_2651);
xor U3465 (N_3465,N_2866,N_2843);
xnor U3466 (N_3466,N_2603,N_2839);
nand U3467 (N_3467,N_2783,N_2541);
xor U3468 (N_3468,N_2691,N_2848);
xor U3469 (N_3469,N_2570,N_2561);
and U3470 (N_3470,N_2786,N_2787);
nand U3471 (N_3471,N_2554,N_2624);
and U3472 (N_3472,N_2582,N_2753);
xor U3473 (N_3473,N_2758,N_2681);
nor U3474 (N_3474,N_2577,N_2578);
and U3475 (N_3475,N_2827,N_2888);
nand U3476 (N_3476,N_2982,N_2698);
and U3477 (N_3477,N_2611,N_2873);
and U3478 (N_3478,N_2604,N_2525);
or U3479 (N_3479,N_2836,N_2861);
nand U3480 (N_3480,N_2958,N_2820);
xnor U3481 (N_3481,N_2709,N_2860);
or U3482 (N_3482,N_2691,N_2784);
and U3483 (N_3483,N_2665,N_2548);
or U3484 (N_3484,N_2703,N_2966);
nor U3485 (N_3485,N_2625,N_2803);
nor U3486 (N_3486,N_2519,N_2690);
nor U3487 (N_3487,N_2528,N_2934);
nand U3488 (N_3488,N_2992,N_2820);
nand U3489 (N_3489,N_2848,N_2588);
xnor U3490 (N_3490,N_2979,N_2567);
or U3491 (N_3491,N_2804,N_2874);
xnor U3492 (N_3492,N_2706,N_2869);
nor U3493 (N_3493,N_2538,N_2783);
nor U3494 (N_3494,N_2878,N_2583);
nand U3495 (N_3495,N_2773,N_2652);
nand U3496 (N_3496,N_2727,N_2519);
nor U3497 (N_3497,N_2877,N_2870);
nor U3498 (N_3498,N_2691,N_2748);
or U3499 (N_3499,N_2622,N_2843);
nand U3500 (N_3500,N_3479,N_3258);
nor U3501 (N_3501,N_3034,N_3336);
nand U3502 (N_3502,N_3011,N_3036);
xnor U3503 (N_3503,N_3261,N_3384);
nor U3504 (N_3504,N_3499,N_3014);
nand U3505 (N_3505,N_3076,N_3108);
xnor U3506 (N_3506,N_3144,N_3337);
and U3507 (N_3507,N_3421,N_3066);
xor U3508 (N_3508,N_3425,N_3130);
nand U3509 (N_3509,N_3098,N_3018);
nand U3510 (N_3510,N_3168,N_3266);
nand U3511 (N_3511,N_3041,N_3118);
xor U3512 (N_3512,N_3075,N_3062);
xor U3513 (N_3513,N_3338,N_3087);
and U3514 (N_3514,N_3442,N_3228);
and U3515 (N_3515,N_3486,N_3453);
xnor U3516 (N_3516,N_3020,N_3471);
or U3517 (N_3517,N_3398,N_3434);
nor U3518 (N_3518,N_3224,N_3200);
nand U3519 (N_3519,N_3423,N_3368);
nand U3520 (N_3520,N_3121,N_3422);
nand U3521 (N_3521,N_3182,N_3220);
or U3522 (N_3522,N_3031,N_3305);
nor U3523 (N_3523,N_3063,N_3099);
nand U3524 (N_3524,N_3458,N_3400);
and U3525 (N_3525,N_3177,N_3496);
or U3526 (N_3526,N_3444,N_3288);
xnor U3527 (N_3527,N_3126,N_3179);
and U3528 (N_3528,N_3407,N_3164);
nand U3529 (N_3529,N_3404,N_3236);
or U3530 (N_3530,N_3498,N_3279);
and U3531 (N_3531,N_3232,N_3351);
or U3532 (N_3532,N_3257,N_3049);
xor U3533 (N_3533,N_3326,N_3252);
and U3534 (N_3534,N_3133,N_3078);
nand U3535 (N_3535,N_3270,N_3097);
nor U3536 (N_3536,N_3308,N_3419);
and U3537 (N_3537,N_3125,N_3072);
nand U3538 (N_3538,N_3093,N_3095);
and U3539 (N_3539,N_3264,N_3199);
and U3540 (N_3540,N_3008,N_3007);
nand U3541 (N_3541,N_3291,N_3058);
xor U3542 (N_3542,N_3023,N_3208);
or U3543 (N_3543,N_3188,N_3235);
nand U3544 (N_3544,N_3156,N_3229);
or U3545 (N_3545,N_3094,N_3077);
and U3546 (N_3546,N_3013,N_3119);
or U3547 (N_3547,N_3397,N_3390);
or U3548 (N_3548,N_3113,N_3280);
or U3549 (N_3549,N_3355,N_3473);
nand U3550 (N_3550,N_3495,N_3477);
nor U3551 (N_3551,N_3433,N_3403);
nor U3552 (N_3552,N_3205,N_3316);
nand U3553 (N_3553,N_3490,N_3203);
or U3554 (N_3554,N_3186,N_3101);
and U3555 (N_3555,N_3366,N_3493);
nand U3556 (N_3556,N_3448,N_3440);
or U3557 (N_3557,N_3492,N_3080);
and U3558 (N_3558,N_3114,N_3281);
and U3559 (N_3559,N_3174,N_3251);
nand U3560 (N_3560,N_3055,N_3475);
or U3561 (N_3561,N_3255,N_3104);
xor U3562 (N_3562,N_3210,N_3382);
nand U3563 (N_3563,N_3047,N_3141);
nand U3564 (N_3564,N_3106,N_3143);
and U3565 (N_3565,N_3309,N_3107);
nor U3566 (N_3566,N_3334,N_3386);
nand U3567 (N_3567,N_3081,N_3438);
or U3568 (N_3568,N_3171,N_3197);
and U3569 (N_3569,N_3370,N_3105);
nand U3570 (N_3570,N_3231,N_3183);
or U3571 (N_3571,N_3322,N_3482);
nand U3572 (N_3572,N_3388,N_3122);
nor U3573 (N_3573,N_3006,N_3226);
and U3574 (N_3574,N_3292,N_3064);
or U3575 (N_3575,N_3132,N_3243);
and U3576 (N_3576,N_3256,N_3227);
or U3577 (N_3577,N_3016,N_3299);
nor U3578 (N_3578,N_3411,N_3116);
and U3579 (N_3579,N_3033,N_3103);
nor U3580 (N_3580,N_3052,N_3408);
xnor U3581 (N_3581,N_3470,N_3165);
or U3582 (N_3582,N_3206,N_3462);
nand U3583 (N_3583,N_3409,N_3367);
or U3584 (N_3584,N_3412,N_3332);
nor U3585 (N_3585,N_3110,N_3348);
nand U3586 (N_3586,N_3166,N_3100);
nand U3587 (N_3587,N_3464,N_3115);
nor U3588 (N_3588,N_3145,N_3276);
xor U3589 (N_3589,N_3304,N_3219);
or U3590 (N_3590,N_3474,N_3497);
nor U3591 (N_3591,N_3446,N_3260);
nand U3592 (N_3592,N_3181,N_3435);
nor U3593 (N_3593,N_3429,N_3185);
and U3594 (N_3594,N_3465,N_3214);
and U3595 (N_3595,N_3040,N_3092);
xnor U3596 (N_3596,N_3417,N_3413);
or U3597 (N_3597,N_3420,N_3494);
xnor U3598 (N_3598,N_3238,N_3472);
nor U3599 (N_3599,N_3259,N_3102);
or U3600 (N_3600,N_3466,N_3035);
nand U3601 (N_3601,N_3415,N_3037);
xnor U3602 (N_3602,N_3377,N_3039);
and U3603 (N_3603,N_3485,N_3149);
xor U3604 (N_3604,N_3216,N_3406);
and U3605 (N_3605,N_3269,N_3050);
or U3606 (N_3606,N_3155,N_3242);
or U3607 (N_3607,N_3053,N_3339);
nor U3608 (N_3608,N_3414,N_3467);
nand U3609 (N_3609,N_3004,N_3287);
nor U3610 (N_3610,N_3191,N_3333);
nor U3611 (N_3611,N_3449,N_3392);
and U3612 (N_3612,N_3432,N_3001);
nand U3613 (N_3613,N_3030,N_3278);
nor U3614 (N_3614,N_3396,N_3300);
xor U3615 (N_3615,N_3074,N_3140);
nor U3616 (N_3616,N_3153,N_3109);
or U3617 (N_3617,N_3330,N_3005);
xor U3618 (N_3618,N_3357,N_3443);
and U3619 (N_3619,N_3211,N_3056);
or U3620 (N_3620,N_3491,N_3002);
nor U3621 (N_3621,N_3343,N_3374);
nor U3622 (N_3622,N_3154,N_3138);
and U3623 (N_3623,N_3057,N_3265);
and U3624 (N_3624,N_3298,N_3213);
or U3625 (N_3625,N_3312,N_3068);
and U3626 (N_3626,N_3321,N_3489);
xor U3627 (N_3627,N_3241,N_3418);
xnor U3628 (N_3628,N_3358,N_3437);
xnor U3629 (N_3629,N_3430,N_3302);
nor U3630 (N_3630,N_3196,N_3246);
nand U3631 (N_3631,N_3083,N_3146);
nor U3632 (N_3632,N_3441,N_3247);
nor U3633 (N_3633,N_3285,N_3431);
and U3634 (N_3634,N_3488,N_3012);
and U3635 (N_3635,N_3178,N_3344);
or U3636 (N_3636,N_3277,N_3051);
and U3637 (N_3637,N_3207,N_3375);
and U3638 (N_3638,N_3328,N_3184);
and U3639 (N_3639,N_3424,N_3478);
or U3640 (N_3640,N_3327,N_3022);
and U3641 (N_3641,N_3283,N_3294);
nand U3642 (N_3642,N_3148,N_3142);
nor U3643 (N_3643,N_3381,N_3027);
and U3644 (N_3644,N_3373,N_3457);
xor U3645 (N_3645,N_3230,N_3065);
and U3646 (N_3646,N_3459,N_3253);
nand U3647 (N_3647,N_3268,N_3352);
and U3648 (N_3648,N_3192,N_3369);
or U3649 (N_3649,N_3376,N_3009);
xor U3650 (N_3650,N_3159,N_3389);
xor U3651 (N_3651,N_3317,N_3239);
xor U3652 (N_3652,N_3029,N_3223);
nor U3653 (N_3653,N_3387,N_3111);
and U3654 (N_3654,N_3198,N_3160);
and U3655 (N_3655,N_3134,N_3271);
nor U3656 (N_3656,N_3028,N_3315);
nor U3657 (N_3657,N_3293,N_3329);
or U3658 (N_3658,N_3372,N_3120);
xor U3659 (N_3659,N_3071,N_3346);
or U3660 (N_3660,N_3451,N_3152);
nor U3661 (N_3661,N_3380,N_3085);
nand U3662 (N_3662,N_3193,N_3324);
nor U3663 (N_3663,N_3139,N_3218);
xnor U3664 (N_3664,N_3314,N_3162);
xor U3665 (N_3665,N_3362,N_3073);
or U3666 (N_3666,N_3342,N_3303);
nor U3667 (N_3667,N_3297,N_3249);
nand U3668 (N_3668,N_3263,N_3383);
xor U3669 (N_3669,N_3289,N_3331);
xnor U3670 (N_3670,N_3395,N_3069);
xnor U3671 (N_3671,N_3086,N_3371);
nand U3672 (N_3672,N_3379,N_3234);
xor U3673 (N_3673,N_3262,N_3117);
xnor U3674 (N_3674,N_3021,N_3436);
or U3675 (N_3675,N_3032,N_3452);
nand U3676 (N_3676,N_3222,N_3468);
nand U3677 (N_3677,N_3127,N_3454);
or U3678 (N_3678,N_3169,N_3067);
and U3679 (N_3679,N_3364,N_3461);
xor U3680 (N_3680,N_3318,N_3157);
and U3681 (N_3681,N_3137,N_3135);
or U3682 (N_3682,N_3447,N_3082);
nand U3683 (N_3683,N_3170,N_3175);
xor U3684 (N_3684,N_3019,N_3254);
or U3685 (N_3685,N_3173,N_3079);
xor U3686 (N_3686,N_3301,N_3089);
and U3687 (N_3687,N_3426,N_3393);
nand U3688 (N_3688,N_3399,N_3167);
and U3689 (N_3689,N_3084,N_3463);
and U3690 (N_3690,N_3319,N_3217);
or U3691 (N_3691,N_3320,N_3003);
or U3692 (N_3692,N_3313,N_3060);
nor U3693 (N_3693,N_3401,N_3307);
nor U3694 (N_3694,N_3090,N_3311);
nor U3695 (N_3695,N_3365,N_3088);
nor U3696 (N_3696,N_3469,N_3354);
xnor U3697 (N_3697,N_3150,N_3195);
nand U3698 (N_3698,N_3024,N_3248);
and U3699 (N_3699,N_3476,N_3353);
nor U3700 (N_3700,N_3483,N_3340);
and U3701 (N_3701,N_3043,N_3295);
and U3702 (N_3702,N_3290,N_3025);
and U3703 (N_3703,N_3445,N_3275);
nor U3704 (N_3704,N_3274,N_3048);
and U3705 (N_3705,N_3487,N_3136);
nor U3706 (N_3706,N_3070,N_3428);
nor U3707 (N_3707,N_3212,N_3410);
or U3708 (N_3708,N_3061,N_3112);
nand U3709 (N_3709,N_3054,N_3042);
nand U3710 (N_3710,N_3296,N_3347);
nand U3711 (N_3711,N_3361,N_3349);
nand U3712 (N_3712,N_3335,N_3310);
or U3713 (N_3713,N_3202,N_3402);
or U3714 (N_3714,N_3484,N_3123);
xor U3715 (N_3715,N_3015,N_3190);
xor U3716 (N_3716,N_3394,N_3245);
and U3717 (N_3717,N_3455,N_3151);
nor U3718 (N_3718,N_3325,N_3350);
xnor U3719 (N_3719,N_3147,N_3359);
nor U3720 (N_3720,N_3385,N_3201);
and U3721 (N_3721,N_3128,N_3163);
or U3722 (N_3722,N_3176,N_3378);
nand U3723 (N_3723,N_3306,N_3194);
xnor U3724 (N_3724,N_3460,N_3046);
nand U3725 (N_3725,N_3017,N_3284);
or U3726 (N_3726,N_3405,N_3323);
and U3727 (N_3727,N_3045,N_3044);
nor U3728 (N_3728,N_3272,N_3391);
nand U3729 (N_3729,N_3026,N_3161);
and U3730 (N_3730,N_3059,N_3189);
and U3731 (N_3731,N_3038,N_3480);
nand U3732 (N_3732,N_3233,N_3250);
nor U3733 (N_3733,N_3124,N_3131);
nor U3734 (N_3734,N_3341,N_3282);
nor U3735 (N_3735,N_3360,N_3356);
nand U3736 (N_3736,N_3267,N_3240);
nor U3737 (N_3737,N_3091,N_3427);
nand U3738 (N_3738,N_3187,N_3204);
and U3739 (N_3739,N_3273,N_3481);
xnor U3740 (N_3740,N_3172,N_3416);
nor U3741 (N_3741,N_3215,N_3244);
and U3742 (N_3742,N_3000,N_3439);
and U3743 (N_3743,N_3345,N_3450);
nor U3744 (N_3744,N_3180,N_3096);
and U3745 (N_3745,N_3237,N_3456);
or U3746 (N_3746,N_3286,N_3158);
nor U3747 (N_3747,N_3363,N_3209);
nor U3748 (N_3748,N_3225,N_3010);
nor U3749 (N_3749,N_3221,N_3129);
xnor U3750 (N_3750,N_3129,N_3212);
nor U3751 (N_3751,N_3403,N_3275);
nand U3752 (N_3752,N_3098,N_3157);
and U3753 (N_3753,N_3497,N_3273);
nand U3754 (N_3754,N_3244,N_3342);
nor U3755 (N_3755,N_3496,N_3329);
xnor U3756 (N_3756,N_3290,N_3419);
and U3757 (N_3757,N_3167,N_3232);
nand U3758 (N_3758,N_3186,N_3444);
xor U3759 (N_3759,N_3444,N_3317);
nand U3760 (N_3760,N_3229,N_3477);
or U3761 (N_3761,N_3396,N_3133);
or U3762 (N_3762,N_3452,N_3268);
nand U3763 (N_3763,N_3473,N_3320);
xor U3764 (N_3764,N_3486,N_3489);
or U3765 (N_3765,N_3268,N_3254);
or U3766 (N_3766,N_3256,N_3164);
nand U3767 (N_3767,N_3317,N_3153);
nor U3768 (N_3768,N_3281,N_3161);
xor U3769 (N_3769,N_3014,N_3070);
and U3770 (N_3770,N_3203,N_3334);
and U3771 (N_3771,N_3151,N_3119);
nand U3772 (N_3772,N_3282,N_3441);
nand U3773 (N_3773,N_3180,N_3140);
or U3774 (N_3774,N_3328,N_3168);
nand U3775 (N_3775,N_3219,N_3362);
and U3776 (N_3776,N_3059,N_3226);
or U3777 (N_3777,N_3155,N_3214);
xnor U3778 (N_3778,N_3461,N_3378);
nand U3779 (N_3779,N_3457,N_3369);
nand U3780 (N_3780,N_3294,N_3062);
nor U3781 (N_3781,N_3145,N_3314);
xor U3782 (N_3782,N_3093,N_3138);
xor U3783 (N_3783,N_3070,N_3272);
nor U3784 (N_3784,N_3269,N_3117);
nand U3785 (N_3785,N_3473,N_3073);
xnor U3786 (N_3786,N_3092,N_3217);
or U3787 (N_3787,N_3431,N_3291);
and U3788 (N_3788,N_3295,N_3187);
or U3789 (N_3789,N_3318,N_3022);
xnor U3790 (N_3790,N_3143,N_3193);
nand U3791 (N_3791,N_3286,N_3054);
nor U3792 (N_3792,N_3115,N_3020);
nand U3793 (N_3793,N_3197,N_3113);
nand U3794 (N_3794,N_3288,N_3052);
and U3795 (N_3795,N_3005,N_3371);
xnor U3796 (N_3796,N_3023,N_3217);
and U3797 (N_3797,N_3441,N_3419);
or U3798 (N_3798,N_3032,N_3364);
nand U3799 (N_3799,N_3190,N_3224);
nand U3800 (N_3800,N_3285,N_3062);
and U3801 (N_3801,N_3251,N_3324);
and U3802 (N_3802,N_3425,N_3329);
nor U3803 (N_3803,N_3142,N_3056);
nor U3804 (N_3804,N_3290,N_3385);
xor U3805 (N_3805,N_3099,N_3187);
nand U3806 (N_3806,N_3055,N_3276);
nand U3807 (N_3807,N_3001,N_3175);
xor U3808 (N_3808,N_3248,N_3480);
or U3809 (N_3809,N_3291,N_3404);
or U3810 (N_3810,N_3299,N_3197);
nor U3811 (N_3811,N_3405,N_3464);
nand U3812 (N_3812,N_3455,N_3313);
nand U3813 (N_3813,N_3364,N_3203);
xor U3814 (N_3814,N_3135,N_3393);
nor U3815 (N_3815,N_3121,N_3459);
nand U3816 (N_3816,N_3059,N_3496);
and U3817 (N_3817,N_3307,N_3003);
xnor U3818 (N_3818,N_3362,N_3028);
or U3819 (N_3819,N_3029,N_3483);
xor U3820 (N_3820,N_3128,N_3306);
or U3821 (N_3821,N_3196,N_3283);
xnor U3822 (N_3822,N_3347,N_3012);
nor U3823 (N_3823,N_3273,N_3469);
xnor U3824 (N_3824,N_3395,N_3025);
xor U3825 (N_3825,N_3110,N_3288);
xor U3826 (N_3826,N_3168,N_3120);
and U3827 (N_3827,N_3469,N_3200);
or U3828 (N_3828,N_3468,N_3362);
nor U3829 (N_3829,N_3215,N_3405);
xor U3830 (N_3830,N_3425,N_3341);
nor U3831 (N_3831,N_3203,N_3370);
nand U3832 (N_3832,N_3446,N_3224);
nand U3833 (N_3833,N_3061,N_3191);
nor U3834 (N_3834,N_3155,N_3027);
nand U3835 (N_3835,N_3435,N_3166);
nor U3836 (N_3836,N_3106,N_3087);
or U3837 (N_3837,N_3452,N_3200);
or U3838 (N_3838,N_3371,N_3478);
nand U3839 (N_3839,N_3083,N_3013);
nand U3840 (N_3840,N_3128,N_3014);
and U3841 (N_3841,N_3428,N_3367);
and U3842 (N_3842,N_3310,N_3474);
xor U3843 (N_3843,N_3041,N_3181);
and U3844 (N_3844,N_3195,N_3382);
xor U3845 (N_3845,N_3300,N_3376);
nand U3846 (N_3846,N_3221,N_3100);
and U3847 (N_3847,N_3054,N_3398);
or U3848 (N_3848,N_3312,N_3185);
or U3849 (N_3849,N_3370,N_3009);
or U3850 (N_3850,N_3375,N_3371);
or U3851 (N_3851,N_3200,N_3215);
nand U3852 (N_3852,N_3084,N_3153);
nand U3853 (N_3853,N_3430,N_3064);
nor U3854 (N_3854,N_3367,N_3269);
nand U3855 (N_3855,N_3439,N_3221);
nor U3856 (N_3856,N_3011,N_3057);
and U3857 (N_3857,N_3348,N_3393);
nand U3858 (N_3858,N_3299,N_3467);
or U3859 (N_3859,N_3485,N_3352);
and U3860 (N_3860,N_3216,N_3176);
and U3861 (N_3861,N_3471,N_3206);
nor U3862 (N_3862,N_3016,N_3096);
nand U3863 (N_3863,N_3067,N_3452);
or U3864 (N_3864,N_3486,N_3294);
and U3865 (N_3865,N_3438,N_3456);
xnor U3866 (N_3866,N_3043,N_3218);
xor U3867 (N_3867,N_3468,N_3498);
nand U3868 (N_3868,N_3068,N_3254);
xor U3869 (N_3869,N_3054,N_3022);
xnor U3870 (N_3870,N_3481,N_3357);
nor U3871 (N_3871,N_3472,N_3430);
xor U3872 (N_3872,N_3391,N_3238);
and U3873 (N_3873,N_3173,N_3422);
xnor U3874 (N_3874,N_3341,N_3197);
nor U3875 (N_3875,N_3063,N_3082);
nor U3876 (N_3876,N_3268,N_3146);
and U3877 (N_3877,N_3422,N_3124);
and U3878 (N_3878,N_3297,N_3474);
or U3879 (N_3879,N_3000,N_3024);
xor U3880 (N_3880,N_3490,N_3493);
nor U3881 (N_3881,N_3143,N_3466);
and U3882 (N_3882,N_3468,N_3171);
xor U3883 (N_3883,N_3087,N_3417);
nand U3884 (N_3884,N_3458,N_3066);
xnor U3885 (N_3885,N_3295,N_3298);
and U3886 (N_3886,N_3066,N_3232);
nand U3887 (N_3887,N_3356,N_3455);
xor U3888 (N_3888,N_3051,N_3404);
xor U3889 (N_3889,N_3483,N_3125);
nor U3890 (N_3890,N_3261,N_3406);
xor U3891 (N_3891,N_3067,N_3230);
nor U3892 (N_3892,N_3336,N_3154);
and U3893 (N_3893,N_3177,N_3447);
or U3894 (N_3894,N_3170,N_3432);
nand U3895 (N_3895,N_3379,N_3426);
nor U3896 (N_3896,N_3021,N_3349);
xor U3897 (N_3897,N_3428,N_3471);
and U3898 (N_3898,N_3461,N_3224);
and U3899 (N_3899,N_3103,N_3452);
xnor U3900 (N_3900,N_3074,N_3107);
or U3901 (N_3901,N_3079,N_3359);
nand U3902 (N_3902,N_3464,N_3254);
and U3903 (N_3903,N_3248,N_3027);
and U3904 (N_3904,N_3193,N_3196);
nand U3905 (N_3905,N_3487,N_3380);
nor U3906 (N_3906,N_3225,N_3364);
or U3907 (N_3907,N_3207,N_3210);
nor U3908 (N_3908,N_3171,N_3046);
and U3909 (N_3909,N_3365,N_3356);
nor U3910 (N_3910,N_3291,N_3429);
nand U3911 (N_3911,N_3423,N_3007);
and U3912 (N_3912,N_3030,N_3294);
xnor U3913 (N_3913,N_3227,N_3343);
nand U3914 (N_3914,N_3100,N_3026);
and U3915 (N_3915,N_3231,N_3381);
nand U3916 (N_3916,N_3143,N_3482);
nand U3917 (N_3917,N_3443,N_3243);
xnor U3918 (N_3918,N_3478,N_3365);
xnor U3919 (N_3919,N_3375,N_3013);
nand U3920 (N_3920,N_3304,N_3487);
nor U3921 (N_3921,N_3058,N_3039);
or U3922 (N_3922,N_3254,N_3381);
and U3923 (N_3923,N_3304,N_3328);
xnor U3924 (N_3924,N_3349,N_3280);
or U3925 (N_3925,N_3012,N_3173);
xnor U3926 (N_3926,N_3039,N_3001);
nand U3927 (N_3927,N_3422,N_3076);
nor U3928 (N_3928,N_3479,N_3111);
xnor U3929 (N_3929,N_3033,N_3200);
nor U3930 (N_3930,N_3114,N_3352);
or U3931 (N_3931,N_3320,N_3025);
nor U3932 (N_3932,N_3012,N_3362);
or U3933 (N_3933,N_3382,N_3076);
nor U3934 (N_3934,N_3155,N_3463);
xor U3935 (N_3935,N_3463,N_3081);
or U3936 (N_3936,N_3497,N_3353);
nor U3937 (N_3937,N_3439,N_3276);
xnor U3938 (N_3938,N_3009,N_3356);
and U3939 (N_3939,N_3487,N_3307);
xnor U3940 (N_3940,N_3197,N_3337);
or U3941 (N_3941,N_3011,N_3460);
and U3942 (N_3942,N_3145,N_3091);
nand U3943 (N_3943,N_3186,N_3336);
or U3944 (N_3944,N_3431,N_3155);
nand U3945 (N_3945,N_3310,N_3187);
and U3946 (N_3946,N_3111,N_3291);
nor U3947 (N_3947,N_3405,N_3347);
nor U3948 (N_3948,N_3487,N_3081);
nor U3949 (N_3949,N_3265,N_3156);
nand U3950 (N_3950,N_3028,N_3412);
xor U3951 (N_3951,N_3498,N_3235);
nor U3952 (N_3952,N_3383,N_3134);
or U3953 (N_3953,N_3107,N_3348);
or U3954 (N_3954,N_3061,N_3411);
and U3955 (N_3955,N_3050,N_3237);
and U3956 (N_3956,N_3354,N_3171);
or U3957 (N_3957,N_3154,N_3279);
xor U3958 (N_3958,N_3094,N_3351);
or U3959 (N_3959,N_3091,N_3252);
nor U3960 (N_3960,N_3163,N_3219);
and U3961 (N_3961,N_3016,N_3246);
xnor U3962 (N_3962,N_3098,N_3089);
and U3963 (N_3963,N_3138,N_3294);
nand U3964 (N_3964,N_3359,N_3412);
nor U3965 (N_3965,N_3277,N_3497);
nor U3966 (N_3966,N_3475,N_3384);
or U3967 (N_3967,N_3390,N_3402);
or U3968 (N_3968,N_3165,N_3085);
and U3969 (N_3969,N_3464,N_3194);
xor U3970 (N_3970,N_3466,N_3255);
xnor U3971 (N_3971,N_3385,N_3454);
or U3972 (N_3972,N_3110,N_3461);
xnor U3973 (N_3973,N_3429,N_3486);
nand U3974 (N_3974,N_3400,N_3260);
and U3975 (N_3975,N_3042,N_3256);
or U3976 (N_3976,N_3297,N_3035);
xor U3977 (N_3977,N_3406,N_3378);
nand U3978 (N_3978,N_3109,N_3220);
nor U3979 (N_3979,N_3237,N_3152);
xnor U3980 (N_3980,N_3417,N_3315);
or U3981 (N_3981,N_3094,N_3340);
xor U3982 (N_3982,N_3259,N_3338);
nand U3983 (N_3983,N_3302,N_3044);
xnor U3984 (N_3984,N_3268,N_3225);
xnor U3985 (N_3985,N_3310,N_3473);
and U3986 (N_3986,N_3368,N_3060);
nor U3987 (N_3987,N_3307,N_3400);
nor U3988 (N_3988,N_3278,N_3305);
nor U3989 (N_3989,N_3372,N_3251);
nor U3990 (N_3990,N_3444,N_3472);
or U3991 (N_3991,N_3101,N_3123);
and U3992 (N_3992,N_3463,N_3359);
and U3993 (N_3993,N_3339,N_3212);
xnor U3994 (N_3994,N_3293,N_3357);
xnor U3995 (N_3995,N_3319,N_3496);
nand U3996 (N_3996,N_3207,N_3341);
nor U3997 (N_3997,N_3439,N_3400);
and U3998 (N_3998,N_3274,N_3317);
xor U3999 (N_3999,N_3208,N_3462);
and U4000 (N_4000,N_3738,N_3932);
or U4001 (N_4001,N_3643,N_3717);
nand U4002 (N_4002,N_3746,N_3968);
nor U4003 (N_4003,N_3922,N_3780);
nand U4004 (N_4004,N_3830,N_3974);
and U4005 (N_4005,N_3826,N_3610);
nand U4006 (N_4006,N_3851,N_3550);
nor U4007 (N_4007,N_3973,N_3852);
xor U4008 (N_4008,N_3701,N_3556);
xor U4009 (N_4009,N_3946,N_3981);
and U4010 (N_4010,N_3602,N_3934);
nor U4011 (N_4011,N_3528,N_3588);
nand U4012 (N_4012,N_3545,N_3658);
nor U4013 (N_4013,N_3950,N_3599);
nand U4014 (N_4014,N_3933,N_3984);
nor U4015 (N_4015,N_3652,N_3989);
nand U4016 (N_4016,N_3657,N_3634);
or U4017 (N_4017,N_3882,N_3879);
nand U4018 (N_4018,N_3894,N_3996);
xnor U4019 (N_4019,N_3690,N_3706);
nor U4020 (N_4020,N_3878,N_3900);
or U4021 (N_4021,N_3551,N_3540);
xor U4022 (N_4022,N_3563,N_3763);
and U4023 (N_4023,N_3951,N_3565);
or U4024 (N_4024,N_3539,N_3770);
and U4025 (N_4025,N_3507,N_3579);
nand U4026 (N_4026,N_3881,N_3749);
and U4027 (N_4027,N_3559,N_3664);
or U4028 (N_4028,N_3532,N_3735);
nor U4029 (N_4029,N_3605,N_3784);
nand U4030 (N_4030,N_3511,N_3668);
or U4031 (N_4031,N_3673,N_3694);
nor U4032 (N_4032,N_3831,N_3815);
and U4033 (N_4033,N_3713,N_3838);
and U4034 (N_4034,N_3716,N_3936);
nand U4035 (N_4035,N_3502,N_3943);
nor U4036 (N_4036,N_3697,N_3889);
nor U4037 (N_4037,N_3589,N_3834);
nand U4038 (N_4038,N_3986,N_3920);
and U4039 (N_4039,N_3711,N_3574);
and U4040 (N_4040,N_3525,N_3843);
nor U4041 (N_4041,N_3773,N_3526);
nand U4042 (N_4042,N_3793,N_3764);
nand U4043 (N_4043,N_3681,N_3560);
and U4044 (N_4044,N_3613,N_3742);
nand U4045 (N_4045,N_3999,N_3504);
nand U4046 (N_4046,N_3725,N_3662);
or U4047 (N_4047,N_3655,N_3594);
nor U4048 (N_4048,N_3731,N_3855);
xor U4049 (N_4049,N_3582,N_3521);
xor U4050 (N_4050,N_3959,N_3872);
xor U4051 (N_4051,N_3935,N_3978);
nor U4052 (N_4052,N_3781,N_3642);
nor U4053 (N_4053,N_3638,N_3863);
nor U4054 (N_4054,N_3908,N_3672);
xnor U4055 (N_4055,N_3636,N_3783);
nor U4056 (N_4056,N_3769,N_3810);
nand U4057 (N_4057,N_3699,N_3649);
nor U4058 (N_4058,N_3670,N_3543);
and U4059 (N_4059,N_3956,N_3760);
xnor U4060 (N_4060,N_3527,N_3917);
or U4061 (N_4061,N_3500,N_3869);
nand U4062 (N_4062,N_3992,N_3693);
and U4063 (N_4063,N_3848,N_3629);
xor U4064 (N_4064,N_3534,N_3802);
nand U4065 (N_4065,N_3627,N_3756);
nor U4066 (N_4066,N_3789,N_3535);
xnor U4067 (N_4067,N_3569,N_3666);
xnor U4068 (N_4068,N_3859,N_3975);
and U4069 (N_4069,N_3868,N_3597);
and U4070 (N_4070,N_3741,N_3998);
nor U4071 (N_4071,N_3876,N_3656);
and U4072 (N_4072,N_3604,N_3586);
xnor U4073 (N_4073,N_3625,N_3779);
xor U4074 (N_4074,N_3547,N_3575);
and U4075 (N_4075,N_3921,N_3555);
or U4076 (N_4076,N_3990,N_3850);
xnor U4077 (N_4077,N_3628,N_3519);
nand U4078 (N_4078,N_3970,N_3748);
xnor U4079 (N_4079,N_3570,N_3911);
xnor U4080 (N_4080,N_3653,N_3710);
nand U4081 (N_4081,N_3660,N_3776);
and U4082 (N_4082,N_3614,N_3651);
and U4083 (N_4083,N_3997,N_3727);
nor U4084 (N_4084,N_3606,N_3558);
nor U4085 (N_4085,N_3562,N_3768);
xor U4086 (N_4086,N_3825,N_3944);
xor U4087 (N_4087,N_3544,N_3958);
or U4088 (N_4088,N_3700,N_3583);
nor U4089 (N_4089,N_3966,N_3593);
xnor U4090 (N_4090,N_3506,N_3572);
or U4091 (N_4091,N_3603,N_3795);
or U4092 (N_4092,N_3592,N_3632);
and U4093 (N_4093,N_3899,N_3745);
nor U4094 (N_4094,N_3661,N_3775);
nor U4095 (N_4095,N_3953,N_3962);
and U4096 (N_4096,N_3564,N_3611);
and U4097 (N_4097,N_3718,N_3704);
or U4098 (N_4098,N_3983,N_3596);
xor U4099 (N_4099,N_3880,N_3621);
or U4100 (N_4100,N_3669,N_3788);
nand U4101 (N_4101,N_3542,N_3686);
nor U4102 (N_4102,N_3679,N_3840);
nor U4103 (N_4103,N_3907,N_3898);
nand U4104 (N_4104,N_3674,N_3685);
nor U4105 (N_4105,N_3541,N_3884);
xnor U4106 (N_4106,N_3811,N_3837);
nand U4107 (N_4107,N_3720,N_3622);
or U4108 (N_4108,N_3896,N_3552);
nor U4109 (N_4109,N_3940,N_3576);
or U4110 (N_4110,N_3639,N_3833);
or U4111 (N_4111,N_3941,N_3906);
nor U4112 (N_4112,N_3754,N_3767);
nor U4113 (N_4113,N_3865,N_3965);
nand U4114 (N_4114,N_3994,N_3626);
nand U4115 (N_4115,N_3696,N_3991);
xor U4116 (N_4116,N_3722,N_3961);
nand U4117 (N_4117,N_3520,N_3530);
nor U4118 (N_4118,N_3601,N_3512);
and U4119 (N_4119,N_3708,N_3912);
xnor U4120 (N_4120,N_3501,N_3942);
or U4121 (N_4121,N_3938,N_3744);
nor U4122 (N_4122,N_3891,N_3967);
xnor U4123 (N_4123,N_3698,N_3772);
nand U4124 (N_4124,N_3774,N_3856);
xor U4125 (N_4125,N_3667,N_3905);
xnor U4126 (N_4126,N_3712,N_3918);
nor U4127 (N_4127,N_3952,N_3835);
xor U4128 (N_4128,N_3609,N_3916);
and U4129 (N_4129,N_3567,N_3612);
nor U4130 (N_4130,N_3791,N_3949);
nand U4131 (N_4131,N_3926,N_3915);
nor U4132 (N_4132,N_3832,N_3647);
or U4133 (N_4133,N_3578,N_3870);
and U4134 (N_4134,N_3929,N_3671);
and U4135 (N_4135,N_3987,N_3573);
nor U4136 (N_4136,N_3822,N_3792);
and U4137 (N_4137,N_3893,N_3729);
or U4138 (N_4138,N_3529,N_3842);
nand U4139 (N_4139,N_3620,N_3508);
or U4140 (N_4140,N_3857,N_3595);
or U4141 (N_4141,N_3641,N_3719);
nand U4142 (N_4142,N_3762,N_3800);
or U4143 (N_4143,N_3703,N_3849);
nor U4144 (N_4144,N_3937,N_3904);
or U4145 (N_4145,N_3515,N_3919);
or U4146 (N_4146,N_3778,N_3549);
or U4147 (N_4147,N_3721,N_3635);
or U4148 (N_4148,N_3633,N_3566);
nor U4149 (N_4149,N_3554,N_3948);
nand U4150 (N_4150,N_3750,N_3568);
xor U4151 (N_4151,N_3980,N_3957);
nor U4152 (N_4152,N_3964,N_3873);
nor U4153 (N_4153,N_3707,N_3702);
or U4154 (N_4154,N_3883,N_3805);
xnor U4155 (N_4155,N_3841,N_3931);
nand U4156 (N_4156,N_3514,N_3839);
and U4157 (N_4157,N_3736,N_3887);
nor U4158 (N_4158,N_3677,N_3737);
nor U4159 (N_4159,N_3797,N_3853);
nand U4160 (N_4160,N_3533,N_3969);
nand U4161 (N_4161,N_3753,N_3523);
nand U4162 (N_4162,N_3709,N_3692);
nand U4163 (N_4163,N_3571,N_3858);
nand U4164 (N_4164,N_3854,N_3799);
nor U4165 (N_4165,N_3874,N_3637);
xor U4166 (N_4166,N_3923,N_3536);
and U4167 (N_4167,N_3758,N_3624);
nor U4168 (N_4168,N_3801,N_3960);
and U4169 (N_4169,N_3650,N_3902);
and U4170 (N_4170,N_3518,N_3765);
nand U4171 (N_4171,N_3927,N_3730);
nor U4172 (N_4172,N_3864,N_3947);
and U4173 (N_4173,N_3819,N_3688);
and U4174 (N_4174,N_3537,N_3646);
or U4175 (N_4175,N_3814,N_3590);
nand U4176 (N_4176,N_3924,N_3875);
nor U4177 (N_4177,N_3695,N_3751);
or U4178 (N_4178,N_3818,N_3977);
or U4179 (N_4179,N_3752,N_3682);
and U4180 (N_4180,N_3598,N_3757);
xnor U4181 (N_4181,N_3732,N_3993);
and U4182 (N_4182,N_3561,N_3786);
and U4183 (N_4183,N_3734,N_3631);
nand U4184 (N_4184,N_3678,N_3971);
nor U4185 (N_4185,N_3548,N_3577);
and U4186 (N_4186,N_3680,N_3743);
xor U4187 (N_4187,N_3817,N_3954);
or U4188 (N_4188,N_3587,N_3824);
and U4189 (N_4189,N_3867,N_3823);
nand U4190 (N_4190,N_3890,N_3985);
nand U4191 (N_4191,N_3726,N_3689);
xnor U4192 (N_4192,N_3691,N_3510);
nand U4193 (N_4193,N_3659,N_3820);
xor U4194 (N_4194,N_3623,N_3546);
or U4195 (N_4195,N_3665,N_3914);
nor U4196 (N_4196,N_3684,N_3617);
and U4197 (N_4197,N_3630,N_3648);
xnor U4198 (N_4198,N_3759,N_3888);
nor U4199 (N_4199,N_3723,N_3538);
nor U4200 (N_4200,N_3581,N_3715);
and U4201 (N_4201,N_3644,N_3844);
and U4202 (N_4202,N_3600,N_3903);
nand U4203 (N_4203,N_3862,N_3930);
nand U4204 (N_4204,N_3683,N_3860);
nor U4205 (N_4205,N_3584,N_3925);
nor U4206 (N_4206,N_3901,N_3733);
nor U4207 (N_4207,N_3976,N_3740);
nand U4208 (N_4208,N_3503,N_3816);
or U4209 (N_4209,N_3829,N_3988);
nand U4210 (N_4210,N_3796,N_3804);
xor U4211 (N_4211,N_3836,N_3798);
nor U4212 (N_4212,N_3963,N_3995);
and U4213 (N_4213,N_3585,N_3813);
xnor U4214 (N_4214,N_3806,N_3982);
nor U4215 (N_4215,N_3885,N_3892);
xor U4216 (N_4216,N_3828,N_3808);
nand U4217 (N_4217,N_3812,N_3616);
and U4218 (N_4218,N_3803,N_3618);
or U4219 (N_4219,N_3714,N_3663);
xor U4220 (N_4220,N_3761,N_3640);
xor U4221 (N_4221,N_3909,N_3787);
and U4222 (N_4222,N_3845,N_3619);
xnor U4223 (N_4223,N_3553,N_3728);
and U4224 (N_4224,N_3782,N_3747);
xor U4225 (N_4225,N_3766,N_3645);
nand U4226 (N_4226,N_3886,N_3846);
xnor U4227 (N_4227,N_3972,N_3522);
and U4228 (N_4228,N_3827,N_3790);
nand U4229 (N_4229,N_3580,N_3739);
xnor U4230 (N_4230,N_3809,N_3531);
xnor U4231 (N_4231,N_3771,N_3807);
and U4232 (N_4232,N_3524,N_3687);
nand U4233 (N_4233,N_3724,N_3505);
nand U4234 (N_4234,N_3557,N_3928);
and U4235 (N_4235,N_3777,N_3945);
xnor U4236 (N_4236,N_3955,N_3785);
and U4237 (N_4237,N_3910,N_3675);
xor U4238 (N_4238,N_3615,N_3755);
nor U4239 (N_4239,N_3913,N_3607);
and U4240 (N_4240,N_3877,N_3895);
nand U4241 (N_4241,N_3821,N_3705);
nand U4242 (N_4242,N_3861,N_3979);
nor U4243 (N_4243,N_3608,N_3866);
and U4244 (N_4244,N_3676,N_3509);
nor U4245 (N_4245,N_3513,N_3591);
xnor U4246 (N_4246,N_3654,N_3897);
and U4247 (N_4247,N_3847,N_3516);
and U4248 (N_4248,N_3517,N_3939);
or U4249 (N_4249,N_3794,N_3871);
or U4250 (N_4250,N_3836,N_3855);
nand U4251 (N_4251,N_3832,N_3826);
xor U4252 (N_4252,N_3599,N_3544);
or U4253 (N_4253,N_3709,N_3752);
xnor U4254 (N_4254,N_3662,N_3543);
and U4255 (N_4255,N_3840,N_3918);
and U4256 (N_4256,N_3912,N_3974);
xnor U4257 (N_4257,N_3651,N_3702);
nand U4258 (N_4258,N_3986,N_3869);
nand U4259 (N_4259,N_3526,N_3912);
or U4260 (N_4260,N_3523,N_3807);
xnor U4261 (N_4261,N_3522,N_3698);
and U4262 (N_4262,N_3909,N_3506);
nand U4263 (N_4263,N_3982,N_3995);
or U4264 (N_4264,N_3852,N_3560);
nand U4265 (N_4265,N_3875,N_3960);
and U4266 (N_4266,N_3874,N_3750);
and U4267 (N_4267,N_3640,N_3840);
xor U4268 (N_4268,N_3986,N_3876);
and U4269 (N_4269,N_3586,N_3934);
or U4270 (N_4270,N_3725,N_3832);
nand U4271 (N_4271,N_3535,N_3573);
xor U4272 (N_4272,N_3848,N_3789);
nor U4273 (N_4273,N_3874,N_3857);
nor U4274 (N_4274,N_3560,N_3848);
or U4275 (N_4275,N_3654,N_3986);
and U4276 (N_4276,N_3715,N_3902);
xnor U4277 (N_4277,N_3965,N_3514);
nor U4278 (N_4278,N_3581,N_3585);
xor U4279 (N_4279,N_3661,N_3962);
xor U4280 (N_4280,N_3618,N_3855);
nand U4281 (N_4281,N_3688,N_3731);
nor U4282 (N_4282,N_3730,N_3559);
or U4283 (N_4283,N_3820,N_3912);
nand U4284 (N_4284,N_3508,N_3971);
or U4285 (N_4285,N_3655,N_3657);
nand U4286 (N_4286,N_3843,N_3628);
xnor U4287 (N_4287,N_3772,N_3739);
or U4288 (N_4288,N_3961,N_3515);
nor U4289 (N_4289,N_3519,N_3786);
and U4290 (N_4290,N_3609,N_3967);
xnor U4291 (N_4291,N_3599,N_3820);
nor U4292 (N_4292,N_3963,N_3726);
and U4293 (N_4293,N_3886,N_3859);
or U4294 (N_4294,N_3940,N_3876);
xor U4295 (N_4295,N_3677,N_3586);
nand U4296 (N_4296,N_3621,N_3840);
nor U4297 (N_4297,N_3861,N_3787);
nand U4298 (N_4298,N_3749,N_3952);
or U4299 (N_4299,N_3723,N_3785);
xor U4300 (N_4300,N_3959,N_3794);
xor U4301 (N_4301,N_3758,N_3895);
and U4302 (N_4302,N_3839,N_3769);
xnor U4303 (N_4303,N_3940,N_3901);
nor U4304 (N_4304,N_3851,N_3951);
and U4305 (N_4305,N_3754,N_3566);
nand U4306 (N_4306,N_3627,N_3957);
nand U4307 (N_4307,N_3783,N_3907);
nor U4308 (N_4308,N_3557,N_3725);
or U4309 (N_4309,N_3957,N_3668);
nand U4310 (N_4310,N_3694,N_3645);
nor U4311 (N_4311,N_3905,N_3791);
and U4312 (N_4312,N_3821,N_3969);
nor U4313 (N_4313,N_3694,N_3592);
xor U4314 (N_4314,N_3800,N_3526);
nand U4315 (N_4315,N_3937,N_3769);
and U4316 (N_4316,N_3881,N_3529);
xnor U4317 (N_4317,N_3812,N_3957);
and U4318 (N_4318,N_3823,N_3988);
nor U4319 (N_4319,N_3752,N_3862);
and U4320 (N_4320,N_3893,N_3607);
nand U4321 (N_4321,N_3811,N_3823);
and U4322 (N_4322,N_3850,N_3636);
and U4323 (N_4323,N_3762,N_3950);
xnor U4324 (N_4324,N_3557,N_3800);
or U4325 (N_4325,N_3504,N_3556);
or U4326 (N_4326,N_3537,N_3824);
nand U4327 (N_4327,N_3665,N_3956);
and U4328 (N_4328,N_3821,N_3924);
nor U4329 (N_4329,N_3573,N_3761);
or U4330 (N_4330,N_3911,N_3750);
or U4331 (N_4331,N_3960,N_3706);
nand U4332 (N_4332,N_3908,N_3728);
nor U4333 (N_4333,N_3682,N_3929);
or U4334 (N_4334,N_3780,N_3897);
xnor U4335 (N_4335,N_3547,N_3510);
nand U4336 (N_4336,N_3655,N_3936);
xnor U4337 (N_4337,N_3786,N_3548);
or U4338 (N_4338,N_3764,N_3609);
or U4339 (N_4339,N_3909,N_3966);
or U4340 (N_4340,N_3711,N_3878);
nand U4341 (N_4341,N_3939,N_3833);
or U4342 (N_4342,N_3923,N_3572);
and U4343 (N_4343,N_3646,N_3618);
and U4344 (N_4344,N_3731,N_3752);
nor U4345 (N_4345,N_3610,N_3881);
xor U4346 (N_4346,N_3922,N_3859);
nor U4347 (N_4347,N_3552,N_3985);
nand U4348 (N_4348,N_3623,N_3930);
xor U4349 (N_4349,N_3918,N_3992);
nor U4350 (N_4350,N_3950,N_3771);
and U4351 (N_4351,N_3791,N_3645);
xnor U4352 (N_4352,N_3599,N_3764);
nand U4353 (N_4353,N_3827,N_3859);
nor U4354 (N_4354,N_3899,N_3846);
xnor U4355 (N_4355,N_3874,N_3971);
nand U4356 (N_4356,N_3821,N_3629);
nor U4357 (N_4357,N_3885,N_3780);
nor U4358 (N_4358,N_3794,N_3533);
or U4359 (N_4359,N_3744,N_3596);
and U4360 (N_4360,N_3560,N_3713);
nand U4361 (N_4361,N_3619,N_3857);
nand U4362 (N_4362,N_3733,N_3956);
nand U4363 (N_4363,N_3885,N_3971);
nand U4364 (N_4364,N_3571,N_3726);
and U4365 (N_4365,N_3864,N_3962);
nand U4366 (N_4366,N_3573,N_3975);
xor U4367 (N_4367,N_3997,N_3575);
xnor U4368 (N_4368,N_3610,N_3581);
and U4369 (N_4369,N_3988,N_3670);
and U4370 (N_4370,N_3965,N_3508);
or U4371 (N_4371,N_3923,N_3885);
and U4372 (N_4372,N_3924,N_3934);
xor U4373 (N_4373,N_3748,N_3565);
nor U4374 (N_4374,N_3599,N_3970);
nand U4375 (N_4375,N_3822,N_3528);
xnor U4376 (N_4376,N_3877,N_3591);
nand U4377 (N_4377,N_3513,N_3595);
nand U4378 (N_4378,N_3990,N_3970);
or U4379 (N_4379,N_3769,N_3702);
xnor U4380 (N_4380,N_3745,N_3740);
and U4381 (N_4381,N_3802,N_3579);
xor U4382 (N_4382,N_3699,N_3859);
nor U4383 (N_4383,N_3875,N_3650);
or U4384 (N_4384,N_3816,N_3894);
and U4385 (N_4385,N_3588,N_3954);
xnor U4386 (N_4386,N_3679,N_3530);
nor U4387 (N_4387,N_3989,N_3525);
nand U4388 (N_4388,N_3651,N_3523);
xor U4389 (N_4389,N_3856,N_3632);
and U4390 (N_4390,N_3904,N_3846);
nand U4391 (N_4391,N_3809,N_3738);
xnor U4392 (N_4392,N_3814,N_3889);
nand U4393 (N_4393,N_3689,N_3956);
xnor U4394 (N_4394,N_3689,N_3967);
xnor U4395 (N_4395,N_3875,N_3776);
and U4396 (N_4396,N_3794,N_3870);
or U4397 (N_4397,N_3697,N_3587);
and U4398 (N_4398,N_3864,N_3534);
nand U4399 (N_4399,N_3618,N_3589);
nand U4400 (N_4400,N_3625,N_3958);
xnor U4401 (N_4401,N_3818,N_3775);
and U4402 (N_4402,N_3845,N_3875);
and U4403 (N_4403,N_3863,N_3741);
and U4404 (N_4404,N_3816,N_3877);
xor U4405 (N_4405,N_3918,N_3821);
nor U4406 (N_4406,N_3729,N_3813);
and U4407 (N_4407,N_3617,N_3587);
and U4408 (N_4408,N_3946,N_3985);
and U4409 (N_4409,N_3912,N_3827);
nand U4410 (N_4410,N_3809,N_3716);
nand U4411 (N_4411,N_3519,N_3800);
nor U4412 (N_4412,N_3941,N_3586);
nor U4413 (N_4413,N_3672,N_3627);
nor U4414 (N_4414,N_3962,N_3771);
nand U4415 (N_4415,N_3636,N_3819);
nor U4416 (N_4416,N_3601,N_3686);
xnor U4417 (N_4417,N_3529,N_3959);
or U4418 (N_4418,N_3731,N_3561);
and U4419 (N_4419,N_3554,N_3853);
nor U4420 (N_4420,N_3855,N_3709);
and U4421 (N_4421,N_3506,N_3806);
nor U4422 (N_4422,N_3748,N_3995);
or U4423 (N_4423,N_3849,N_3589);
xnor U4424 (N_4424,N_3924,N_3917);
nor U4425 (N_4425,N_3517,N_3870);
or U4426 (N_4426,N_3942,N_3576);
xnor U4427 (N_4427,N_3742,N_3744);
xnor U4428 (N_4428,N_3632,N_3962);
and U4429 (N_4429,N_3721,N_3529);
xnor U4430 (N_4430,N_3809,N_3912);
and U4431 (N_4431,N_3889,N_3919);
nor U4432 (N_4432,N_3514,N_3701);
xor U4433 (N_4433,N_3580,N_3974);
and U4434 (N_4434,N_3954,N_3523);
or U4435 (N_4435,N_3769,N_3532);
nand U4436 (N_4436,N_3520,N_3901);
xnor U4437 (N_4437,N_3558,N_3969);
and U4438 (N_4438,N_3659,N_3616);
nand U4439 (N_4439,N_3909,N_3918);
xnor U4440 (N_4440,N_3660,N_3892);
and U4441 (N_4441,N_3868,N_3971);
or U4442 (N_4442,N_3549,N_3927);
or U4443 (N_4443,N_3780,N_3540);
nor U4444 (N_4444,N_3732,N_3517);
xor U4445 (N_4445,N_3583,N_3806);
nor U4446 (N_4446,N_3993,N_3755);
nand U4447 (N_4447,N_3677,N_3738);
nor U4448 (N_4448,N_3558,N_3704);
or U4449 (N_4449,N_3689,N_3810);
nand U4450 (N_4450,N_3992,N_3676);
or U4451 (N_4451,N_3773,N_3813);
or U4452 (N_4452,N_3759,N_3823);
xor U4453 (N_4453,N_3804,N_3760);
and U4454 (N_4454,N_3825,N_3549);
nor U4455 (N_4455,N_3514,N_3879);
nor U4456 (N_4456,N_3702,N_3733);
xnor U4457 (N_4457,N_3548,N_3787);
nand U4458 (N_4458,N_3971,N_3826);
nand U4459 (N_4459,N_3992,N_3854);
nor U4460 (N_4460,N_3669,N_3875);
and U4461 (N_4461,N_3558,N_3881);
or U4462 (N_4462,N_3533,N_3690);
nand U4463 (N_4463,N_3733,N_3583);
nand U4464 (N_4464,N_3987,N_3752);
and U4465 (N_4465,N_3970,N_3543);
or U4466 (N_4466,N_3961,N_3573);
xor U4467 (N_4467,N_3917,N_3538);
xor U4468 (N_4468,N_3536,N_3528);
or U4469 (N_4469,N_3545,N_3893);
and U4470 (N_4470,N_3747,N_3612);
and U4471 (N_4471,N_3801,N_3752);
nand U4472 (N_4472,N_3637,N_3853);
or U4473 (N_4473,N_3864,N_3913);
or U4474 (N_4474,N_3567,N_3684);
xnor U4475 (N_4475,N_3752,N_3851);
xnor U4476 (N_4476,N_3501,N_3737);
nor U4477 (N_4477,N_3865,N_3959);
nor U4478 (N_4478,N_3633,N_3536);
nand U4479 (N_4479,N_3704,N_3526);
nand U4480 (N_4480,N_3834,N_3826);
or U4481 (N_4481,N_3607,N_3917);
nor U4482 (N_4482,N_3718,N_3511);
or U4483 (N_4483,N_3710,N_3525);
nor U4484 (N_4484,N_3693,N_3549);
or U4485 (N_4485,N_3900,N_3812);
xnor U4486 (N_4486,N_3886,N_3745);
xor U4487 (N_4487,N_3824,N_3909);
and U4488 (N_4488,N_3743,N_3839);
nand U4489 (N_4489,N_3714,N_3937);
nor U4490 (N_4490,N_3633,N_3997);
or U4491 (N_4491,N_3988,N_3755);
nand U4492 (N_4492,N_3526,N_3662);
or U4493 (N_4493,N_3618,N_3892);
xnor U4494 (N_4494,N_3631,N_3953);
nand U4495 (N_4495,N_3571,N_3520);
xor U4496 (N_4496,N_3501,N_3704);
nor U4497 (N_4497,N_3959,N_3503);
nand U4498 (N_4498,N_3796,N_3872);
xnor U4499 (N_4499,N_3885,N_3731);
xnor U4500 (N_4500,N_4315,N_4196);
nand U4501 (N_4501,N_4421,N_4161);
and U4502 (N_4502,N_4252,N_4336);
nand U4503 (N_4503,N_4121,N_4066);
nor U4504 (N_4504,N_4133,N_4167);
nor U4505 (N_4505,N_4023,N_4046);
nand U4506 (N_4506,N_4459,N_4188);
xnor U4507 (N_4507,N_4223,N_4217);
nor U4508 (N_4508,N_4091,N_4227);
nand U4509 (N_4509,N_4187,N_4195);
nor U4510 (N_4510,N_4224,N_4116);
nor U4511 (N_4511,N_4286,N_4221);
nor U4512 (N_4512,N_4237,N_4498);
and U4513 (N_4513,N_4083,N_4175);
nor U4514 (N_4514,N_4174,N_4086);
or U4515 (N_4515,N_4367,N_4151);
or U4516 (N_4516,N_4104,N_4429);
or U4517 (N_4517,N_4369,N_4481);
or U4518 (N_4518,N_4006,N_4404);
and U4519 (N_4519,N_4106,N_4071);
and U4520 (N_4520,N_4433,N_4359);
nand U4521 (N_4521,N_4181,N_4263);
or U4522 (N_4522,N_4290,N_4009);
nand U4523 (N_4523,N_4031,N_4453);
and U4524 (N_4524,N_4138,N_4222);
nor U4525 (N_4525,N_4279,N_4392);
or U4526 (N_4526,N_4406,N_4305);
nor U4527 (N_4527,N_4037,N_4247);
or U4528 (N_4528,N_4059,N_4328);
xnor U4529 (N_4529,N_4028,N_4027);
nand U4530 (N_4530,N_4266,N_4487);
or U4531 (N_4531,N_4233,N_4025);
or U4532 (N_4532,N_4370,N_4403);
xnor U4533 (N_4533,N_4136,N_4039);
nand U4534 (N_4534,N_4372,N_4354);
nand U4535 (N_4535,N_4441,N_4358);
or U4536 (N_4536,N_4013,N_4268);
or U4537 (N_4537,N_4199,N_4388);
nor U4538 (N_4538,N_4271,N_4148);
or U4539 (N_4539,N_4464,N_4493);
or U4540 (N_4540,N_4343,N_4140);
and U4541 (N_4541,N_4134,N_4042);
nand U4542 (N_4542,N_4490,N_4093);
nand U4543 (N_4543,N_4128,N_4381);
nand U4544 (N_4544,N_4455,N_4332);
and U4545 (N_4545,N_4225,N_4312);
and U4546 (N_4546,N_4194,N_4488);
or U4547 (N_4547,N_4415,N_4007);
xor U4548 (N_4548,N_4072,N_4430);
or U4549 (N_4549,N_4055,N_4172);
and U4550 (N_4550,N_4241,N_4178);
and U4551 (N_4551,N_4064,N_4211);
nand U4552 (N_4552,N_4463,N_4101);
and U4553 (N_4553,N_4496,N_4057);
and U4554 (N_4554,N_4362,N_4373);
and U4555 (N_4555,N_4452,N_4314);
and U4556 (N_4556,N_4287,N_4125);
and U4557 (N_4557,N_4230,N_4061);
nand U4558 (N_4558,N_4000,N_4232);
and U4559 (N_4559,N_4448,N_4226);
nor U4560 (N_4560,N_4288,N_4143);
and U4561 (N_4561,N_4327,N_4095);
or U4562 (N_4562,N_4020,N_4052);
xnor U4563 (N_4563,N_4215,N_4016);
xnor U4564 (N_4564,N_4119,N_4479);
or U4565 (N_4565,N_4352,N_4130);
and U4566 (N_4566,N_4077,N_4219);
nand U4567 (N_4567,N_4147,N_4473);
and U4568 (N_4568,N_4274,N_4258);
or U4569 (N_4569,N_4350,N_4337);
xnor U4570 (N_4570,N_4228,N_4160);
nand U4571 (N_4571,N_4108,N_4179);
nor U4572 (N_4572,N_4102,N_4003);
xnor U4573 (N_4573,N_4303,N_4065);
nand U4574 (N_4574,N_4345,N_4084);
or U4575 (N_4575,N_4468,N_4386);
nand U4576 (N_4576,N_4238,N_4280);
xor U4577 (N_4577,N_4159,N_4425);
nand U4578 (N_4578,N_4236,N_4400);
or U4579 (N_4579,N_4396,N_4250);
nor U4580 (N_4580,N_4026,N_4293);
and U4581 (N_4581,N_4063,N_4357);
xor U4582 (N_4582,N_4257,N_4475);
and U4583 (N_4583,N_4262,N_4017);
and U4584 (N_4584,N_4409,N_4109);
nor U4585 (N_4585,N_4088,N_4438);
and U4586 (N_4586,N_4351,N_4371);
nand U4587 (N_4587,N_4024,N_4335);
or U4588 (N_4588,N_4348,N_4096);
and U4589 (N_4589,N_4365,N_4255);
or U4590 (N_4590,N_4368,N_4480);
or U4591 (N_4591,N_4304,N_4176);
xor U4592 (N_4592,N_4030,N_4110);
nor U4593 (N_4593,N_4321,N_4146);
nor U4594 (N_4594,N_4156,N_4244);
nor U4595 (N_4595,N_4465,N_4051);
nor U4596 (N_4596,N_4380,N_4135);
nand U4597 (N_4597,N_4246,N_4001);
xor U4598 (N_4598,N_4193,N_4344);
xnor U4599 (N_4599,N_4150,N_4427);
and U4600 (N_4600,N_4300,N_4416);
nand U4601 (N_4601,N_4398,N_4054);
and U4602 (N_4602,N_4056,N_4137);
nor U4603 (N_4603,N_4454,N_4387);
nand U4604 (N_4604,N_4318,N_4089);
nor U4605 (N_4605,N_4002,N_4495);
nor U4606 (N_4606,N_4360,N_4379);
nor U4607 (N_4607,N_4131,N_4302);
and U4608 (N_4608,N_4442,N_4278);
xnor U4609 (N_4609,N_4053,N_4395);
nor U4610 (N_4610,N_4322,N_4486);
or U4611 (N_4611,N_4333,N_4316);
and U4612 (N_4612,N_4289,N_4005);
or U4613 (N_4613,N_4308,N_4450);
nor U4614 (N_4614,N_4177,N_4434);
and U4615 (N_4615,N_4437,N_4098);
and U4616 (N_4616,N_4440,N_4213);
nand U4617 (N_4617,N_4447,N_4375);
xnor U4618 (N_4618,N_4218,N_4382);
nand U4619 (N_4619,N_4165,N_4426);
and U4620 (N_4620,N_4040,N_4112);
nor U4621 (N_4621,N_4256,N_4184);
or U4622 (N_4622,N_4127,N_4324);
nor U4623 (N_4623,N_4100,N_4259);
and U4624 (N_4624,N_4021,N_4331);
nor U4625 (N_4625,N_4129,N_4377);
xnor U4626 (N_4626,N_4295,N_4389);
nor U4627 (N_4627,N_4347,N_4260);
xnor U4628 (N_4628,N_4422,N_4018);
nand U4629 (N_4629,N_4044,N_4163);
or U4630 (N_4630,N_4466,N_4418);
or U4631 (N_4631,N_4231,N_4067);
xor U4632 (N_4632,N_4203,N_4154);
xnor U4633 (N_4633,N_4043,N_4275);
nor U4634 (N_4634,N_4074,N_4180);
or U4635 (N_4635,N_4298,N_4338);
and U4636 (N_4636,N_4008,N_4451);
xnor U4637 (N_4637,N_4402,N_4277);
and U4638 (N_4638,N_4190,N_4197);
or U4639 (N_4639,N_4182,N_4097);
or U4640 (N_4640,N_4124,N_4309);
xnor U4641 (N_4641,N_4145,N_4294);
nand U4642 (N_4642,N_4253,N_4458);
nand U4643 (N_4643,N_4269,N_4323);
nand U4644 (N_4644,N_4385,N_4022);
xor U4645 (N_4645,N_4366,N_4050);
and U4646 (N_4646,N_4378,N_4114);
or U4647 (N_4647,N_4317,N_4446);
or U4648 (N_4648,N_4405,N_4411);
xnor U4649 (N_4649,N_4393,N_4126);
and U4650 (N_4650,N_4132,N_4113);
nand U4651 (N_4651,N_4094,N_4254);
xor U4652 (N_4652,N_4192,N_4273);
and U4653 (N_4653,N_4157,N_4342);
or U4654 (N_4654,N_4270,N_4149);
and U4655 (N_4655,N_4183,N_4204);
or U4656 (N_4656,N_4346,N_4449);
or U4657 (N_4657,N_4423,N_4220);
and U4658 (N_4658,N_4281,N_4082);
or U4659 (N_4659,N_4472,N_4339);
and U4660 (N_4660,N_4329,N_4185);
xor U4661 (N_4661,N_4060,N_4436);
or U4662 (N_4662,N_4469,N_4435);
nor U4663 (N_4663,N_4341,N_4410);
xnor U4664 (N_4664,N_4240,N_4474);
or U4665 (N_4665,N_4296,N_4153);
nor U4666 (N_4666,N_4364,N_4048);
xnor U4667 (N_4667,N_4122,N_4186);
xor U4668 (N_4668,N_4099,N_4297);
xor U4669 (N_4669,N_4394,N_4092);
or U4670 (N_4670,N_4210,N_4170);
and U4671 (N_4671,N_4115,N_4047);
nand U4672 (N_4672,N_4325,N_4103);
or U4673 (N_4673,N_4205,N_4216);
nor U4674 (N_4674,N_4477,N_4045);
or U4675 (N_4675,N_4189,N_4162);
and U4676 (N_4676,N_4310,N_4497);
xnor U4677 (N_4677,N_4212,N_4191);
nor U4678 (N_4678,N_4340,N_4070);
xor U4679 (N_4679,N_4141,N_4432);
nor U4680 (N_4680,N_4471,N_4173);
and U4681 (N_4681,N_4408,N_4489);
nand U4682 (N_4682,N_4390,N_4476);
or U4683 (N_4683,N_4363,N_4120);
nand U4684 (N_4684,N_4248,N_4424);
and U4685 (N_4685,N_4090,N_4249);
nand U4686 (N_4686,N_4142,N_4158);
or U4687 (N_4687,N_4326,N_4164);
and U4688 (N_4688,N_4062,N_4209);
or U4689 (N_4689,N_4330,N_4198);
nand U4690 (N_4690,N_4033,N_4035);
or U4691 (N_4691,N_4374,N_4267);
or U4692 (N_4692,N_4272,N_4041);
nand U4693 (N_4693,N_4292,N_4011);
or U4694 (N_4694,N_4492,N_4264);
and U4695 (N_4695,N_4123,N_4361);
or U4696 (N_4696,N_4038,N_4313);
and U4697 (N_4697,N_4384,N_4235);
nand U4698 (N_4698,N_4032,N_4311);
xnor U4699 (N_4699,N_4420,N_4201);
xor U4700 (N_4700,N_4306,N_4456);
nand U4701 (N_4701,N_4319,N_4107);
xor U4702 (N_4702,N_4208,N_4111);
xnor U4703 (N_4703,N_4320,N_4484);
xor U4704 (N_4704,N_4012,N_4355);
xnor U4705 (N_4705,N_4284,N_4261);
nand U4706 (N_4706,N_4036,N_4291);
or U4707 (N_4707,N_4407,N_4049);
nor U4708 (N_4708,N_4207,N_4282);
and U4709 (N_4709,N_4397,N_4245);
and U4710 (N_4710,N_4087,N_4229);
nand U4711 (N_4711,N_4349,N_4285);
nor U4712 (N_4712,N_4353,N_4080);
or U4713 (N_4713,N_4058,N_4118);
xnor U4714 (N_4714,N_4478,N_4383);
or U4715 (N_4715,N_4417,N_4034);
nor U4716 (N_4716,N_4485,N_4019);
nand U4717 (N_4717,N_4015,N_4073);
and U4718 (N_4718,N_4243,N_4470);
xnor U4719 (N_4719,N_4029,N_4068);
nor U4720 (N_4720,N_4069,N_4171);
xor U4721 (N_4721,N_4356,N_4168);
and U4722 (N_4722,N_4139,N_4307);
nor U4723 (N_4723,N_4200,N_4169);
nor U4724 (N_4724,N_4239,N_4414);
nand U4725 (N_4725,N_4391,N_4460);
nand U4726 (N_4726,N_4445,N_4401);
and U4727 (N_4727,N_4491,N_4004);
nor U4728 (N_4728,N_4265,N_4010);
nor U4729 (N_4729,N_4144,N_4166);
or U4730 (N_4730,N_4242,N_4079);
nor U4731 (N_4731,N_4413,N_4444);
and U4732 (N_4732,N_4152,N_4467);
nand U4733 (N_4733,N_4081,N_4461);
or U4734 (N_4734,N_4206,N_4443);
and U4735 (N_4735,N_4499,N_4251);
and U4736 (N_4736,N_4457,N_4419);
xnor U4737 (N_4737,N_4105,N_4399);
nor U4738 (N_4738,N_4482,N_4376);
xnor U4739 (N_4739,N_4299,N_4076);
nor U4740 (N_4740,N_4202,N_4276);
and U4741 (N_4741,N_4301,N_4334);
xor U4742 (N_4742,N_4078,N_4412);
and U4743 (N_4743,N_4462,N_4283);
nand U4744 (N_4744,N_4075,N_4155);
xor U4745 (N_4745,N_4428,N_4014);
nor U4746 (N_4746,N_4439,N_4234);
or U4747 (N_4747,N_4483,N_4494);
and U4748 (N_4748,N_4214,N_4431);
xor U4749 (N_4749,N_4085,N_4117);
nand U4750 (N_4750,N_4416,N_4312);
or U4751 (N_4751,N_4406,N_4380);
xnor U4752 (N_4752,N_4119,N_4172);
and U4753 (N_4753,N_4353,N_4073);
and U4754 (N_4754,N_4346,N_4281);
nand U4755 (N_4755,N_4353,N_4346);
and U4756 (N_4756,N_4366,N_4221);
and U4757 (N_4757,N_4492,N_4012);
xor U4758 (N_4758,N_4377,N_4035);
nor U4759 (N_4759,N_4084,N_4211);
nor U4760 (N_4760,N_4116,N_4102);
xor U4761 (N_4761,N_4194,N_4461);
xnor U4762 (N_4762,N_4005,N_4213);
nor U4763 (N_4763,N_4253,N_4075);
nand U4764 (N_4764,N_4044,N_4376);
or U4765 (N_4765,N_4156,N_4090);
or U4766 (N_4766,N_4369,N_4104);
xnor U4767 (N_4767,N_4486,N_4381);
nor U4768 (N_4768,N_4364,N_4235);
nor U4769 (N_4769,N_4003,N_4408);
nand U4770 (N_4770,N_4260,N_4466);
nand U4771 (N_4771,N_4154,N_4288);
or U4772 (N_4772,N_4226,N_4365);
nor U4773 (N_4773,N_4283,N_4316);
nand U4774 (N_4774,N_4224,N_4251);
or U4775 (N_4775,N_4403,N_4201);
and U4776 (N_4776,N_4065,N_4333);
xnor U4777 (N_4777,N_4308,N_4073);
nor U4778 (N_4778,N_4198,N_4043);
and U4779 (N_4779,N_4193,N_4055);
nor U4780 (N_4780,N_4352,N_4411);
or U4781 (N_4781,N_4370,N_4192);
and U4782 (N_4782,N_4053,N_4459);
xor U4783 (N_4783,N_4232,N_4303);
nand U4784 (N_4784,N_4217,N_4089);
nand U4785 (N_4785,N_4332,N_4324);
and U4786 (N_4786,N_4494,N_4166);
or U4787 (N_4787,N_4319,N_4247);
nor U4788 (N_4788,N_4020,N_4213);
nand U4789 (N_4789,N_4490,N_4105);
or U4790 (N_4790,N_4065,N_4093);
nor U4791 (N_4791,N_4152,N_4174);
nand U4792 (N_4792,N_4028,N_4168);
nor U4793 (N_4793,N_4308,N_4496);
nor U4794 (N_4794,N_4440,N_4126);
or U4795 (N_4795,N_4495,N_4023);
nor U4796 (N_4796,N_4470,N_4393);
and U4797 (N_4797,N_4300,N_4373);
and U4798 (N_4798,N_4228,N_4029);
xnor U4799 (N_4799,N_4419,N_4141);
and U4800 (N_4800,N_4127,N_4317);
xor U4801 (N_4801,N_4377,N_4339);
or U4802 (N_4802,N_4055,N_4093);
nor U4803 (N_4803,N_4146,N_4454);
xnor U4804 (N_4804,N_4143,N_4194);
xor U4805 (N_4805,N_4334,N_4203);
nand U4806 (N_4806,N_4467,N_4496);
nand U4807 (N_4807,N_4369,N_4489);
xor U4808 (N_4808,N_4128,N_4491);
and U4809 (N_4809,N_4296,N_4315);
xnor U4810 (N_4810,N_4147,N_4032);
and U4811 (N_4811,N_4083,N_4242);
and U4812 (N_4812,N_4206,N_4018);
nand U4813 (N_4813,N_4123,N_4171);
xnor U4814 (N_4814,N_4382,N_4142);
and U4815 (N_4815,N_4278,N_4134);
nand U4816 (N_4816,N_4199,N_4140);
or U4817 (N_4817,N_4184,N_4455);
xnor U4818 (N_4818,N_4399,N_4342);
nand U4819 (N_4819,N_4361,N_4174);
or U4820 (N_4820,N_4115,N_4039);
nand U4821 (N_4821,N_4411,N_4052);
or U4822 (N_4822,N_4447,N_4476);
nor U4823 (N_4823,N_4360,N_4400);
xnor U4824 (N_4824,N_4146,N_4038);
xnor U4825 (N_4825,N_4341,N_4202);
nand U4826 (N_4826,N_4279,N_4121);
nand U4827 (N_4827,N_4003,N_4018);
xor U4828 (N_4828,N_4249,N_4307);
nor U4829 (N_4829,N_4280,N_4131);
xnor U4830 (N_4830,N_4455,N_4138);
and U4831 (N_4831,N_4085,N_4302);
xnor U4832 (N_4832,N_4272,N_4435);
nor U4833 (N_4833,N_4172,N_4031);
and U4834 (N_4834,N_4264,N_4090);
xnor U4835 (N_4835,N_4196,N_4085);
nor U4836 (N_4836,N_4419,N_4223);
nor U4837 (N_4837,N_4450,N_4004);
nor U4838 (N_4838,N_4265,N_4103);
and U4839 (N_4839,N_4496,N_4115);
xor U4840 (N_4840,N_4098,N_4494);
or U4841 (N_4841,N_4017,N_4015);
and U4842 (N_4842,N_4242,N_4121);
nor U4843 (N_4843,N_4307,N_4039);
nor U4844 (N_4844,N_4076,N_4135);
or U4845 (N_4845,N_4081,N_4370);
and U4846 (N_4846,N_4118,N_4211);
and U4847 (N_4847,N_4296,N_4300);
or U4848 (N_4848,N_4402,N_4113);
nand U4849 (N_4849,N_4270,N_4004);
or U4850 (N_4850,N_4151,N_4088);
or U4851 (N_4851,N_4125,N_4026);
nor U4852 (N_4852,N_4401,N_4469);
or U4853 (N_4853,N_4323,N_4000);
nor U4854 (N_4854,N_4010,N_4115);
or U4855 (N_4855,N_4396,N_4379);
or U4856 (N_4856,N_4075,N_4313);
nor U4857 (N_4857,N_4348,N_4292);
or U4858 (N_4858,N_4064,N_4296);
nor U4859 (N_4859,N_4402,N_4472);
nand U4860 (N_4860,N_4420,N_4114);
xor U4861 (N_4861,N_4200,N_4039);
xor U4862 (N_4862,N_4257,N_4262);
nor U4863 (N_4863,N_4117,N_4069);
nand U4864 (N_4864,N_4152,N_4204);
nand U4865 (N_4865,N_4483,N_4071);
nor U4866 (N_4866,N_4376,N_4325);
nand U4867 (N_4867,N_4356,N_4286);
nand U4868 (N_4868,N_4480,N_4483);
or U4869 (N_4869,N_4221,N_4013);
xor U4870 (N_4870,N_4285,N_4232);
and U4871 (N_4871,N_4013,N_4048);
and U4872 (N_4872,N_4237,N_4210);
nand U4873 (N_4873,N_4055,N_4016);
or U4874 (N_4874,N_4482,N_4061);
or U4875 (N_4875,N_4200,N_4235);
nor U4876 (N_4876,N_4287,N_4181);
nand U4877 (N_4877,N_4124,N_4329);
or U4878 (N_4878,N_4082,N_4130);
nor U4879 (N_4879,N_4420,N_4087);
or U4880 (N_4880,N_4321,N_4204);
xnor U4881 (N_4881,N_4489,N_4254);
xnor U4882 (N_4882,N_4283,N_4496);
xnor U4883 (N_4883,N_4483,N_4391);
nor U4884 (N_4884,N_4167,N_4426);
and U4885 (N_4885,N_4439,N_4295);
and U4886 (N_4886,N_4485,N_4365);
xor U4887 (N_4887,N_4212,N_4101);
xnor U4888 (N_4888,N_4120,N_4362);
or U4889 (N_4889,N_4204,N_4471);
or U4890 (N_4890,N_4040,N_4457);
nand U4891 (N_4891,N_4065,N_4475);
xnor U4892 (N_4892,N_4162,N_4195);
and U4893 (N_4893,N_4049,N_4082);
and U4894 (N_4894,N_4092,N_4468);
nor U4895 (N_4895,N_4068,N_4201);
or U4896 (N_4896,N_4341,N_4260);
nor U4897 (N_4897,N_4349,N_4174);
xor U4898 (N_4898,N_4430,N_4499);
or U4899 (N_4899,N_4473,N_4036);
xnor U4900 (N_4900,N_4454,N_4480);
and U4901 (N_4901,N_4316,N_4486);
nor U4902 (N_4902,N_4143,N_4203);
and U4903 (N_4903,N_4358,N_4027);
nor U4904 (N_4904,N_4047,N_4421);
nor U4905 (N_4905,N_4077,N_4148);
nor U4906 (N_4906,N_4286,N_4409);
nor U4907 (N_4907,N_4068,N_4203);
nand U4908 (N_4908,N_4086,N_4019);
nand U4909 (N_4909,N_4104,N_4309);
nand U4910 (N_4910,N_4494,N_4442);
xnor U4911 (N_4911,N_4156,N_4220);
and U4912 (N_4912,N_4168,N_4090);
nor U4913 (N_4913,N_4241,N_4343);
xor U4914 (N_4914,N_4293,N_4397);
or U4915 (N_4915,N_4171,N_4213);
and U4916 (N_4916,N_4216,N_4207);
or U4917 (N_4917,N_4313,N_4181);
or U4918 (N_4918,N_4020,N_4370);
nor U4919 (N_4919,N_4228,N_4109);
or U4920 (N_4920,N_4084,N_4272);
and U4921 (N_4921,N_4129,N_4359);
and U4922 (N_4922,N_4378,N_4157);
and U4923 (N_4923,N_4012,N_4294);
nand U4924 (N_4924,N_4314,N_4341);
or U4925 (N_4925,N_4092,N_4381);
or U4926 (N_4926,N_4210,N_4496);
and U4927 (N_4927,N_4227,N_4326);
nand U4928 (N_4928,N_4377,N_4280);
xor U4929 (N_4929,N_4290,N_4399);
xnor U4930 (N_4930,N_4286,N_4122);
nand U4931 (N_4931,N_4147,N_4439);
nand U4932 (N_4932,N_4203,N_4077);
and U4933 (N_4933,N_4397,N_4315);
and U4934 (N_4934,N_4396,N_4226);
or U4935 (N_4935,N_4456,N_4277);
xnor U4936 (N_4936,N_4133,N_4027);
xor U4937 (N_4937,N_4031,N_4408);
and U4938 (N_4938,N_4158,N_4218);
or U4939 (N_4939,N_4409,N_4010);
nor U4940 (N_4940,N_4055,N_4023);
nor U4941 (N_4941,N_4354,N_4423);
and U4942 (N_4942,N_4436,N_4493);
xor U4943 (N_4943,N_4129,N_4069);
or U4944 (N_4944,N_4351,N_4065);
nor U4945 (N_4945,N_4026,N_4348);
or U4946 (N_4946,N_4424,N_4119);
nand U4947 (N_4947,N_4088,N_4017);
or U4948 (N_4948,N_4149,N_4482);
and U4949 (N_4949,N_4278,N_4068);
nor U4950 (N_4950,N_4456,N_4065);
or U4951 (N_4951,N_4218,N_4194);
and U4952 (N_4952,N_4433,N_4096);
nor U4953 (N_4953,N_4007,N_4295);
or U4954 (N_4954,N_4058,N_4305);
and U4955 (N_4955,N_4457,N_4334);
and U4956 (N_4956,N_4015,N_4088);
xnor U4957 (N_4957,N_4207,N_4457);
nor U4958 (N_4958,N_4394,N_4073);
and U4959 (N_4959,N_4240,N_4010);
nor U4960 (N_4960,N_4246,N_4108);
xor U4961 (N_4961,N_4236,N_4166);
nor U4962 (N_4962,N_4391,N_4344);
and U4963 (N_4963,N_4272,N_4024);
nor U4964 (N_4964,N_4354,N_4028);
or U4965 (N_4965,N_4406,N_4450);
or U4966 (N_4966,N_4001,N_4091);
nand U4967 (N_4967,N_4400,N_4458);
and U4968 (N_4968,N_4419,N_4104);
and U4969 (N_4969,N_4252,N_4206);
or U4970 (N_4970,N_4160,N_4220);
and U4971 (N_4971,N_4102,N_4249);
and U4972 (N_4972,N_4026,N_4196);
xor U4973 (N_4973,N_4220,N_4048);
nand U4974 (N_4974,N_4038,N_4495);
nor U4975 (N_4975,N_4307,N_4494);
nand U4976 (N_4976,N_4487,N_4062);
nand U4977 (N_4977,N_4499,N_4375);
nand U4978 (N_4978,N_4413,N_4323);
or U4979 (N_4979,N_4093,N_4480);
nor U4980 (N_4980,N_4436,N_4496);
or U4981 (N_4981,N_4054,N_4471);
nor U4982 (N_4982,N_4013,N_4489);
nand U4983 (N_4983,N_4148,N_4167);
xnor U4984 (N_4984,N_4048,N_4329);
nor U4985 (N_4985,N_4371,N_4446);
and U4986 (N_4986,N_4245,N_4124);
or U4987 (N_4987,N_4050,N_4030);
nor U4988 (N_4988,N_4456,N_4424);
or U4989 (N_4989,N_4296,N_4038);
or U4990 (N_4990,N_4015,N_4240);
nand U4991 (N_4991,N_4249,N_4001);
xnor U4992 (N_4992,N_4459,N_4117);
xor U4993 (N_4993,N_4455,N_4253);
and U4994 (N_4994,N_4219,N_4350);
nor U4995 (N_4995,N_4089,N_4331);
xor U4996 (N_4996,N_4252,N_4139);
or U4997 (N_4997,N_4232,N_4221);
or U4998 (N_4998,N_4131,N_4213);
xnor U4999 (N_4999,N_4425,N_4324);
and U5000 (N_5000,N_4511,N_4598);
nand U5001 (N_5001,N_4543,N_4951);
xnor U5002 (N_5002,N_4952,N_4644);
xnor U5003 (N_5003,N_4504,N_4651);
or U5004 (N_5004,N_4891,N_4601);
nand U5005 (N_5005,N_4917,N_4958);
nand U5006 (N_5006,N_4707,N_4596);
xor U5007 (N_5007,N_4607,N_4531);
nor U5008 (N_5008,N_4815,N_4557);
or U5009 (N_5009,N_4565,N_4969);
or U5010 (N_5010,N_4701,N_4911);
nor U5011 (N_5011,N_4714,N_4791);
xor U5012 (N_5012,N_4930,N_4666);
xor U5013 (N_5013,N_4756,N_4896);
nor U5014 (N_5014,N_4932,N_4840);
xnor U5015 (N_5015,N_4956,N_4757);
or U5016 (N_5016,N_4819,N_4551);
xnor U5017 (N_5017,N_4509,N_4984);
or U5018 (N_5018,N_4905,N_4540);
xnor U5019 (N_5019,N_4670,N_4763);
and U5020 (N_5020,N_4992,N_4805);
nor U5021 (N_5021,N_4765,N_4977);
or U5022 (N_5022,N_4910,N_4667);
xor U5023 (N_5023,N_4500,N_4944);
xnor U5024 (N_5024,N_4697,N_4597);
nor U5025 (N_5025,N_4909,N_4722);
or U5026 (N_5026,N_4586,N_4547);
xor U5027 (N_5027,N_4580,N_4945);
nand U5028 (N_5028,N_4664,N_4548);
nor U5029 (N_5029,N_4904,N_4690);
and U5030 (N_5030,N_4792,N_4934);
nor U5031 (N_5031,N_4704,N_4529);
and U5032 (N_5032,N_4686,N_4927);
or U5033 (N_5033,N_4518,N_4674);
and U5034 (N_5034,N_4589,N_4936);
nor U5035 (N_5035,N_4859,N_4535);
nor U5036 (N_5036,N_4829,N_4705);
and U5037 (N_5037,N_4894,N_4938);
xnor U5038 (N_5038,N_4620,N_4654);
or U5039 (N_5039,N_4700,N_4549);
and U5040 (N_5040,N_4542,N_4685);
or U5041 (N_5041,N_4827,N_4550);
nand U5042 (N_5042,N_4659,N_4991);
and U5043 (N_5043,N_4861,N_4862);
nor U5044 (N_5044,N_4788,N_4652);
nor U5045 (N_5045,N_4799,N_4955);
nor U5046 (N_5046,N_4858,N_4983);
nand U5047 (N_5047,N_4773,N_4972);
or U5048 (N_5048,N_4880,N_4558);
nand U5049 (N_5049,N_4512,N_4692);
nor U5050 (N_5050,N_4820,N_4957);
or U5051 (N_5051,N_4808,N_4741);
nor U5052 (N_5052,N_4650,N_4860);
or U5053 (N_5053,N_4678,N_4689);
xnor U5054 (N_5054,N_4618,N_4522);
xor U5055 (N_5055,N_4948,N_4585);
xor U5056 (N_5056,N_4903,N_4530);
nand U5057 (N_5057,N_4662,N_4886);
xnor U5058 (N_5058,N_4574,N_4502);
or U5059 (N_5059,N_4754,N_4834);
nand U5060 (N_5060,N_4831,N_4570);
xor U5061 (N_5061,N_4852,N_4780);
nand U5062 (N_5062,N_4617,N_4559);
or U5063 (N_5063,N_4723,N_4821);
and U5064 (N_5064,N_4682,N_4939);
and U5065 (N_5065,N_4793,N_4514);
nand U5066 (N_5066,N_4605,N_4889);
and U5067 (N_5067,N_4643,N_4761);
and U5068 (N_5068,N_4978,N_4851);
nand U5069 (N_5069,N_4606,N_4625);
xnor U5070 (N_5070,N_4516,N_4536);
and U5071 (N_5071,N_4642,N_4968);
and U5072 (N_5072,N_4645,N_4582);
nand U5073 (N_5073,N_4712,N_4553);
and U5074 (N_5074,N_4874,N_4520);
nor U5075 (N_5075,N_4916,N_4668);
or U5076 (N_5076,N_4676,N_4818);
nand U5077 (N_5077,N_4735,N_4881);
xor U5078 (N_5078,N_4912,N_4836);
nand U5079 (N_5079,N_4844,N_4869);
nand U5080 (N_5080,N_4753,N_4814);
or U5081 (N_5081,N_4672,N_4593);
xnor U5082 (N_5082,N_4615,N_4898);
or U5083 (N_5083,N_4716,N_4564);
or U5084 (N_5084,N_4947,N_4552);
and U5085 (N_5085,N_4738,N_4680);
nor U5086 (N_5086,N_4866,N_4508);
xor U5087 (N_5087,N_4506,N_4648);
and U5088 (N_5088,N_4568,N_4647);
or U5089 (N_5089,N_4503,N_4528);
nor U5090 (N_5090,N_4973,N_4519);
nand U5091 (N_5091,N_4865,N_4892);
nor U5092 (N_5092,N_4742,N_4687);
and U5093 (N_5093,N_4640,N_4538);
xor U5094 (N_5094,N_4628,N_4800);
nand U5095 (N_5095,N_4863,N_4781);
and U5096 (N_5096,N_4604,N_4962);
and U5097 (N_5097,N_4942,N_4671);
nor U5098 (N_5098,N_4710,N_4846);
nand U5099 (N_5099,N_4525,N_4822);
xor U5100 (N_5100,N_4760,N_4796);
or U5101 (N_5101,N_4609,N_4751);
and U5102 (N_5102,N_4750,N_4599);
and U5103 (N_5103,N_4576,N_4539);
nor U5104 (N_5104,N_4825,N_4885);
xnor U5105 (N_5105,N_4941,N_4766);
xnor U5106 (N_5106,N_4785,N_4595);
or U5107 (N_5107,N_4635,N_4949);
nand U5108 (N_5108,N_4933,N_4849);
nor U5109 (N_5109,N_4720,N_4675);
xnor U5110 (N_5110,N_4613,N_4940);
xor U5111 (N_5111,N_4867,N_4526);
or U5112 (N_5112,N_4787,N_4556);
xnor U5113 (N_5113,N_4993,N_4994);
xor U5114 (N_5114,N_4807,N_4581);
or U5115 (N_5115,N_4673,N_4562);
or U5116 (N_5116,N_4711,N_4816);
nand U5117 (N_5117,N_4563,N_4771);
or U5118 (N_5118,N_4677,N_4870);
or U5119 (N_5119,N_4517,N_4501);
nor U5120 (N_5120,N_4578,N_4812);
nor U5121 (N_5121,N_4986,N_4876);
nand U5122 (N_5122,N_4946,N_4975);
nor U5123 (N_5123,N_4926,N_4826);
xnor U5124 (N_5124,N_4830,N_4713);
or U5125 (N_5125,N_4626,N_4541);
xnor U5126 (N_5126,N_4641,N_4657);
xnor U5127 (N_5127,N_4708,N_4967);
nand U5128 (N_5128,N_4612,N_4614);
or U5129 (N_5129,N_4928,N_4832);
xnor U5130 (N_5130,N_4848,N_4669);
nor U5131 (N_5131,N_4706,N_4798);
nand U5132 (N_5132,N_4505,N_4809);
nor U5133 (N_5133,N_4923,N_4663);
nor U5134 (N_5134,N_4767,N_4739);
nor U5135 (N_5135,N_4914,N_4619);
or U5136 (N_5136,N_4545,N_4950);
or U5137 (N_5137,N_4913,N_4696);
and U5138 (N_5138,N_4731,N_4684);
or U5139 (N_5139,N_4890,N_4811);
or U5140 (N_5140,N_4527,N_4954);
xor U5141 (N_5141,N_4532,N_4510);
xnor U5142 (N_5142,N_4931,N_4721);
and U5143 (N_5143,N_4694,N_4699);
or U5144 (N_5144,N_4729,N_4824);
and U5145 (N_5145,N_4665,N_4769);
nor U5146 (N_5146,N_4806,N_4728);
and U5147 (N_5147,N_4797,N_4681);
and U5148 (N_5148,N_4744,N_4918);
xnor U5149 (N_5149,N_4843,N_4600);
nor U5150 (N_5150,N_4872,N_4871);
and U5151 (N_5151,N_4772,N_4649);
xnor U5152 (N_5152,N_4971,N_4507);
nand U5153 (N_5153,N_4884,N_4554);
nor U5154 (N_5154,N_4718,N_4810);
nand U5155 (N_5155,N_4887,N_4786);
or U5156 (N_5156,N_4996,N_4813);
and U5157 (N_5157,N_4976,N_4734);
or U5158 (N_5158,N_4775,N_4803);
and U5159 (N_5159,N_4856,N_4778);
nand U5160 (N_5160,N_4835,N_4634);
or U5161 (N_5161,N_4864,N_4515);
nor U5162 (N_5162,N_4842,N_4770);
nor U5163 (N_5163,N_4733,N_4925);
nand U5164 (N_5164,N_4658,N_4745);
nor U5165 (N_5165,N_4857,N_4988);
and U5166 (N_5166,N_4782,N_4583);
and U5167 (N_5167,N_4998,N_4985);
or U5168 (N_5168,N_4762,N_4592);
xor U5169 (N_5169,N_4883,N_4660);
xor U5170 (N_5170,N_4732,N_4833);
or U5171 (N_5171,N_4779,N_4655);
nand U5172 (N_5172,N_4736,N_4629);
nand U5173 (N_5173,N_4747,N_4603);
nand U5174 (N_5174,N_4725,N_4639);
xnor U5175 (N_5175,N_4995,N_4758);
and U5176 (N_5176,N_4590,N_4979);
xor U5177 (N_5177,N_4661,N_4960);
or U5178 (N_5178,N_4524,N_4997);
nand U5179 (N_5179,N_4743,N_4573);
nor U5180 (N_5180,N_4823,N_4567);
xor U5181 (N_5181,N_4521,N_4577);
xor U5182 (N_5182,N_4873,N_4627);
xnor U5183 (N_5183,N_4555,N_4943);
nand U5184 (N_5184,N_4841,N_4566);
nand U5185 (N_5185,N_4953,N_4828);
or U5186 (N_5186,N_4879,N_4924);
xnor U5187 (N_5187,N_4533,N_4882);
xnor U5188 (N_5188,N_4919,N_4877);
or U5189 (N_5189,N_4688,N_4980);
and U5190 (N_5190,N_4715,N_4776);
and U5191 (N_5191,N_4937,N_4569);
or U5192 (N_5192,N_4907,N_4717);
nand U5193 (N_5193,N_4847,N_4587);
and U5194 (N_5194,N_4560,N_4746);
nand U5195 (N_5195,N_4768,N_4632);
and U5196 (N_5196,N_4989,N_4591);
and U5197 (N_5197,N_4817,N_4868);
or U5198 (N_5198,N_4878,N_4637);
and U5199 (N_5199,N_4638,N_4893);
nand U5200 (N_5200,N_4683,N_4959);
nor U5201 (N_5201,N_4624,N_4752);
nand U5202 (N_5202,N_4794,N_4915);
xor U5203 (N_5203,N_4902,N_4534);
nand U5204 (N_5204,N_4964,N_4982);
or U5205 (N_5205,N_4774,N_4724);
and U5206 (N_5206,N_4875,N_4895);
nor U5207 (N_5207,N_4572,N_4588);
and U5208 (N_5208,N_4630,N_4777);
or U5209 (N_5209,N_4921,N_4839);
and U5210 (N_5210,N_4608,N_4804);
and U5211 (N_5211,N_4575,N_4730);
nor U5212 (N_5212,N_4748,N_4790);
xor U5213 (N_5213,N_4963,N_4691);
nand U5214 (N_5214,N_4611,N_4656);
xor U5215 (N_5215,N_4726,N_4789);
nor U5216 (N_5216,N_4653,N_4709);
nand U5217 (N_5217,N_4900,N_4537);
nand U5218 (N_5218,N_4679,N_4523);
nand U5219 (N_5219,N_4693,N_4801);
nand U5220 (N_5220,N_4929,N_4571);
nand U5221 (N_5221,N_4719,N_4631);
xnor U5222 (N_5222,N_4854,N_4795);
nand U5223 (N_5223,N_4633,N_4561);
nand U5224 (N_5224,N_4755,N_4513);
or U5225 (N_5225,N_4784,N_4837);
nor U5226 (N_5226,N_4899,N_4802);
nor U5227 (N_5227,N_4702,N_4698);
and U5228 (N_5228,N_4855,N_4616);
or U5229 (N_5229,N_4740,N_4737);
nor U5230 (N_5230,N_4646,N_4546);
nor U5231 (N_5231,N_4544,N_4579);
and U5232 (N_5232,N_4961,N_4935);
nor U5233 (N_5233,N_4897,N_4623);
xor U5234 (N_5234,N_4922,N_4727);
nand U5235 (N_5235,N_4906,N_4602);
nand U5236 (N_5236,N_4594,N_4584);
and U5237 (N_5237,N_4764,N_4783);
nor U5238 (N_5238,N_4990,N_4908);
nand U5239 (N_5239,N_4703,N_4920);
nor U5240 (N_5240,N_4974,N_4970);
nand U5241 (N_5241,N_4610,N_4853);
or U5242 (N_5242,N_4838,N_4759);
and U5243 (N_5243,N_4981,N_4966);
or U5244 (N_5244,N_4622,N_4749);
nand U5245 (N_5245,N_4695,N_4987);
nor U5246 (N_5246,N_4621,N_4888);
or U5247 (N_5247,N_4636,N_4965);
nor U5248 (N_5248,N_4901,N_4850);
nor U5249 (N_5249,N_4999,N_4845);
nor U5250 (N_5250,N_4860,N_4734);
and U5251 (N_5251,N_4616,N_4831);
nand U5252 (N_5252,N_4856,N_4978);
nor U5253 (N_5253,N_4712,N_4608);
xnor U5254 (N_5254,N_4834,N_4698);
or U5255 (N_5255,N_4899,N_4557);
or U5256 (N_5256,N_4754,N_4914);
nand U5257 (N_5257,N_4830,N_4711);
or U5258 (N_5258,N_4826,N_4514);
and U5259 (N_5259,N_4916,N_4759);
and U5260 (N_5260,N_4984,N_4712);
or U5261 (N_5261,N_4818,N_4813);
or U5262 (N_5262,N_4899,N_4542);
nor U5263 (N_5263,N_4756,N_4739);
and U5264 (N_5264,N_4720,N_4510);
and U5265 (N_5265,N_4730,N_4917);
xnor U5266 (N_5266,N_4672,N_4623);
xor U5267 (N_5267,N_4572,N_4981);
or U5268 (N_5268,N_4573,N_4856);
xor U5269 (N_5269,N_4887,N_4637);
and U5270 (N_5270,N_4625,N_4701);
or U5271 (N_5271,N_4654,N_4802);
and U5272 (N_5272,N_4959,N_4883);
nor U5273 (N_5273,N_4823,N_4557);
and U5274 (N_5274,N_4710,N_4617);
xnor U5275 (N_5275,N_4779,N_4541);
nor U5276 (N_5276,N_4549,N_4886);
nor U5277 (N_5277,N_4985,N_4996);
nand U5278 (N_5278,N_4783,N_4637);
or U5279 (N_5279,N_4887,N_4645);
nand U5280 (N_5280,N_4987,N_4628);
xnor U5281 (N_5281,N_4666,N_4841);
and U5282 (N_5282,N_4742,N_4810);
or U5283 (N_5283,N_4624,N_4826);
and U5284 (N_5284,N_4978,N_4600);
nand U5285 (N_5285,N_4891,N_4804);
nand U5286 (N_5286,N_4772,N_4782);
nand U5287 (N_5287,N_4606,N_4862);
nand U5288 (N_5288,N_4895,N_4572);
xor U5289 (N_5289,N_4699,N_4702);
xor U5290 (N_5290,N_4959,N_4717);
or U5291 (N_5291,N_4991,N_4735);
nand U5292 (N_5292,N_4997,N_4999);
or U5293 (N_5293,N_4608,N_4754);
nand U5294 (N_5294,N_4801,N_4845);
xor U5295 (N_5295,N_4854,N_4785);
nor U5296 (N_5296,N_4751,N_4884);
or U5297 (N_5297,N_4656,N_4590);
xor U5298 (N_5298,N_4951,N_4590);
xor U5299 (N_5299,N_4616,N_4675);
or U5300 (N_5300,N_4801,N_4873);
xor U5301 (N_5301,N_4571,N_4875);
and U5302 (N_5302,N_4871,N_4705);
or U5303 (N_5303,N_4742,N_4862);
and U5304 (N_5304,N_4870,N_4860);
xnor U5305 (N_5305,N_4649,N_4644);
nor U5306 (N_5306,N_4712,N_4697);
or U5307 (N_5307,N_4520,N_4571);
or U5308 (N_5308,N_4586,N_4681);
nor U5309 (N_5309,N_4770,N_4568);
xor U5310 (N_5310,N_4664,N_4931);
or U5311 (N_5311,N_4861,N_4914);
or U5312 (N_5312,N_4609,N_4781);
and U5313 (N_5313,N_4919,N_4796);
or U5314 (N_5314,N_4928,N_4848);
nand U5315 (N_5315,N_4705,N_4790);
and U5316 (N_5316,N_4647,N_4977);
or U5317 (N_5317,N_4905,N_4842);
nand U5318 (N_5318,N_4843,N_4947);
nand U5319 (N_5319,N_4682,N_4659);
xor U5320 (N_5320,N_4864,N_4761);
nor U5321 (N_5321,N_4979,N_4507);
nor U5322 (N_5322,N_4817,N_4679);
nor U5323 (N_5323,N_4892,N_4651);
or U5324 (N_5324,N_4692,N_4544);
or U5325 (N_5325,N_4928,N_4560);
or U5326 (N_5326,N_4896,N_4794);
or U5327 (N_5327,N_4761,N_4880);
nand U5328 (N_5328,N_4541,N_4571);
nor U5329 (N_5329,N_4674,N_4927);
and U5330 (N_5330,N_4759,N_4574);
nand U5331 (N_5331,N_4795,N_4645);
xor U5332 (N_5332,N_4998,N_4547);
nand U5333 (N_5333,N_4718,N_4706);
nand U5334 (N_5334,N_4888,N_4606);
nor U5335 (N_5335,N_4904,N_4636);
nand U5336 (N_5336,N_4860,N_4665);
and U5337 (N_5337,N_4830,N_4512);
nor U5338 (N_5338,N_4740,N_4786);
or U5339 (N_5339,N_4951,N_4732);
nor U5340 (N_5340,N_4791,N_4511);
nand U5341 (N_5341,N_4779,N_4961);
and U5342 (N_5342,N_4997,N_4597);
nand U5343 (N_5343,N_4553,N_4627);
and U5344 (N_5344,N_4825,N_4845);
nor U5345 (N_5345,N_4966,N_4912);
and U5346 (N_5346,N_4898,N_4812);
or U5347 (N_5347,N_4611,N_4706);
and U5348 (N_5348,N_4736,N_4562);
xnor U5349 (N_5349,N_4769,N_4953);
and U5350 (N_5350,N_4796,N_4683);
or U5351 (N_5351,N_4591,N_4573);
xor U5352 (N_5352,N_4990,N_4839);
xor U5353 (N_5353,N_4811,N_4881);
or U5354 (N_5354,N_4953,N_4632);
nand U5355 (N_5355,N_4983,N_4518);
or U5356 (N_5356,N_4759,N_4599);
or U5357 (N_5357,N_4819,N_4982);
nand U5358 (N_5358,N_4699,N_4871);
or U5359 (N_5359,N_4820,N_4572);
and U5360 (N_5360,N_4943,N_4852);
and U5361 (N_5361,N_4530,N_4637);
xor U5362 (N_5362,N_4788,N_4866);
xnor U5363 (N_5363,N_4540,N_4770);
nor U5364 (N_5364,N_4615,N_4868);
or U5365 (N_5365,N_4807,N_4517);
or U5366 (N_5366,N_4852,N_4858);
and U5367 (N_5367,N_4897,N_4993);
xor U5368 (N_5368,N_4776,N_4857);
and U5369 (N_5369,N_4618,N_4801);
and U5370 (N_5370,N_4573,N_4597);
or U5371 (N_5371,N_4873,N_4698);
or U5372 (N_5372,N_4575,N_4880);
or U5373 (N_5373,N_4610,N_4699);
or U5374 (N_5374,N_4836,N_4522);
and U5375 (N_5375,N_4655,N_4783);
or U5376 (N_5376,N_4694,N_4723);
nor U5377 (N_5377,N_4606,N_4938);
or U5378 (N_5378,N_4836,N_4693);
nor U5379 (N_5379,N_4905,N_4927);
nand U5380 (N_5380,N_4581,N_4690);
or U5381 (N_5381,N_4532,N_4583);
nor U5382 (N_5382,N_4971,N_4837);
nor U5383 (N_5383,N_4904,N_4515);
xnor U5384 (N_5384,N_4663,N_4731);
and U5385 (N_5385,N_4727,N_4808);
nand U5386 (N_5386,N_4721,N_4576);
or U5387 (N_5387,N_4852,N_4640);
nor U5388 (N_5388,N_4526,N_4752);
and U5389 (N_5389,N_4920,N_4801);
or U5390 (N_5390,N_4834,N_4722);
xor U5391 (N_5391,N_4572,N_4819);
or U5392 (N_5392,N_4759,N_4938);
and U5393 (N_5393,N_4544,N_4742);
nor U5394 (N_5394,N_4600,N_4848);
xor U5395 (N_5395,N_4824,N_4699);
nor U5396 (N_5396,N_4626,N_4621);
nand U5397 (N_5397,N_4896,N_4515);
nor U5398 (N_5398,N_4803,N_4656);
nor U5399 (N_5399,N_4587,N_4500);
or U5400 (N_5400,N_4835,N_4829);
or U5401 (N_5401,N_4852,N_4655);
xnor U5402 (N_5402,N_4886,N_4806);
nand U5403 (N_5403,N_4971,N_4905);
nand U5404 (N_5404,N_4910,N_4937);
nor U5405 (N_5405,N_4976,N_4750);
and U5406 (N_5406,N_4517,N_4805);
nor U5407 (N_5407,N_4755,N_4695);
and U5408 (N_5408,N_4680,N_4704);
or U5409 (N_5409,N_4510,N_4557);
nor U5410 (N_5410,N_4900,N_4891);
nand U5411 (N_5411,N_4824,N_4794);
and U5412 (N_5412,N_4999,N_4662);
nor U5413 (N_5413,N_4783,N_4735);
xor U5414 (N_5414,N_4624,N_4786);
nand U5415 (N_5415,N_4924,N_4717);
nor U5416 (N_5416,N_4683,N_4626);
or U5417 (N_5417,N_4995,N_4623);
or U5418 (N_5418,N_4682,N_4635);
and U5419 (N_5419,N_4787,N_4770);
nand U5420 (N_5420,N_4545,N_4619);
or U5421 (N_5421,N_4928,N_4556);
nand U5422 (N_5422,N_4884,N_4507);
or U5423 (N_5423,N_4675,N_4695);
and U5424 (N_5424,N_4877,N_4697);
xnor U5425 (N_5425,N_4809,N_4600);
and U5426 (N_5426,N_4637,N_4961);
xor U5427 (N_5427,N_4873,N_4681);
and U5428 (N_5428,N_4751,N_4552);
xor U5429 (N_5429,N_4992,N_4788);
xor U5430 (N_5430,N_4610,N_4614);
and U5431 (N_5431,N_4600,N_4816);
or U5432 (N_5432,N_4675,N_4601);
nand U5433 (N_5433,N_4699,N_4556);
nand U5434 (N_5434,N_4845,N_4524);
or U5435 (N_5435,N_4715,N_4998);
nor U5436 (N_5436,N_4889,N_4952);
or U5437 (N_5437,N_4614,N_4987);
or U5438 (N_5438,N_4667,N_4509);
or U5439 (N_5439,N_4793,N_4891);
and U5440 (N_5440,N_4791,N_4673);
nor U5441 (N_5441,N_4838,N_4537);
and U5442 (N_5442,N_4997,N_4648);
xnor U5443 (N_5443,N_4671,N_4876);
and U5444 (N_5444,N_4637,N_4514);
nand U5445 (N_5445,N_4559,N_4675);
nor U5446 (N_5446,N_4991,N_4856);
and U5447 (N_5447,N_4546,N_4615);
nand U5448 (N_5448,N_4582,N_4847);
nor U5449 (N_5449,N_4785,N_4718);
or U5450 (N_5450,N_4720,N_4725);
xnor U5451 (N_5451,N_4846,N_4916);
nand U5452 (N_5452,N_4547,N_4560);
nor U5453 (N_5453,N_4778,N_4590);
xnor U5454 (N_5454,N_4878,N_4717);
or U5455 (N_5455,N_4727,N_4906);
nor U5456 (N_5456,N_4751,N_4955);
nor U5457 (N_5457,N_4789,N_4765);
nand U5458 (N_5458,N_4746,N_4747);
nor U5459 (N_5459,N_4506,N_4925);
xor U5460 (N_5460,N_4648,N_4538);
and U5461 (N_5461,N_4564,N_4515);
xnor U5462 (N_5462,N_4770,N_4588);
nand U5463 (N_5463,N_4944,N_4553);
or U5464 (N_5464,N_4612,N_4691);
nand U5465 (N_5465,N_4571,N_4635);
or U5466 (N_5466,N_4574,N_4611);
or U5467 (N_5467,N_4773,N_4589);
nor U5468 (N_5468,N_4554,N_4771);
nand U5469 (N_5469,N_4947,N_4719);
nor U5470 (N_5470,N_4593,N_4712);
and U5471 (N_5471,N_4586,N_4560);
nor U5472 (N_5472,N_4808,N_4666);
xnor U5473 (N_5473,N_4789,N_4700);
nor U5474 (N_5474,N_4782,N_4727);
and U5475 (N_5475,N_4866,N_4846);
nor U5476 (N_5476,N_4695,N_4705);
xor U5477 (N_5477,N_4534,N_4998);
nand U5478 (N_5478,N_4513,N_4821);
and U5479 (N_5479,N_4582,N_4935);
nor U5480 (N_5480,N_4784,N_4985);
nand U5481 (N_5481,N_4563,N_4991);
xnor U5482 (N_5482,N_4860,N_4528);
nor U5483 (N_5483,N_4707,N_4628);
xor U5484 (N_5484,N_4752,N_4780);
and U5485 (N_5485,N_4733,N_4958);
nor U5486 (N_5486,N_4709,N_4544);
xnor U5487 (N_5487,N_4583,N_4855);
or U5488 (N_5488,N_4950,N_4663);
xnor U5489 (N_5489,N_4556,N_4910);
or U5490 (N_5490,N_4648,N_4564);
nand U5491 (N_5491,N_4677,N_4625);
or U5492 (N_5492,N_4742,N_4680);
and U5493 (N_5493,N_4786,N_4635);
nand U5494 (N_5494,N_4726,N_4888);
nor U5495 (N_5495,N_4983,N_4874);
nand U5496 (N_5496,N_4593,N_4529);
and U5497 (N_5497,N_4582,N_4838);
xnor U5498 (N_5498,N_4846,N_4537);
and U5499 (N_5499,N_4823,N_4586);
nor U5500 (N_5500,N_5267,N_5184);
xor U5501 (N_5501,N_5358,N_5375);
nor U5502 (N_5502,N_5260,N_5286);
nand U5503 (N_5503,N_5187,N_5317);
xnor U5504 (N_5504,N_5203,N_5193);
nand U5505 (N_5505,N_5298,N_5185);
nand U5506 (N_5506,N_5023,N_5295);
nand U5507 (N_5507,N_5109,N_5439);
xor U5508 (N_5508,N_5173,N_5389);
or U5509 (N_5509,N_5336,N_5388);
xor U5510 (N_5510,N_5199,N_5441);
and U5511 (N_5511,N_5150,N_5430);
nor U5512 (N_5512,N_5299,N_5106);
xnor U5513 (N_5513,N_5281,N_5280);
nand U5514 (N_5514,N_5138,N_5357);
nand U5515 (N_5515,N_5059,N_5294);
xor U5516 (N_5516,N_5119,N_5425);
or U5517 (N_5517,N_5355,N_5458);
and U5518 (N_5518,N_5255,N_5137);
and U5519 (N_5519,N_5334,N_5016);
or U5520 (N_5520,N_5379,N_5321);
nor U5521 (N_5521,N_5026,N_5302);
or U5522 (N_5522,N_5052,N_5035);
and U5523 (N_5523,N_5333,N_5475);
and U5524 (N_5524,N_5019,N_5010);
nand U5525 (N_5525,N_5311,N_5253);
xnor U5526 (N_5526,N_5102,N_5380);
nor U5527 (N_5527,N_5285,N_5248);
xor U5528 (N_5528,N_5161,N_5291);
xnor U5529 (N_5529,N_5340,N_5217);
xor U5530 (N_5530,N_5367,N_5022);
nand U5531 (N_5531,N_5178,N_5120);
nand U5532 (N_5532,N_5081,N_5142);
and U5533 (N_5533,N_5435,N_5180);
xnor U5534 (N_5534,N_5172,N_5235);
and U5535 (N_5535,N_5247,N_5234);
or U5536 (N_5536,N_5211,N_5196);
nand U5537 (N_5537,N_5098,N_5432);
nand U5538 (N_5538,N_5316,N_5058);
nand U5539 (N_5539,N_5040,N_5224);
xnor U5540 (N_5540,N_5467,N_5214);
nor U5541 (N_5541,N_5320,N_5393);
nor U5542 (N_5542,N_5404,N_5384);
and U5543 (N_5543,N_5129,N_5112);
nand U5544 (N_5544,N_5126,N_5075);
nand U5545 (N_5545,N_5139,N_5155);
and U5546 (N_5546,N_5485,N_5216);
and U5547 (N_5547,N_5352,N_5319);
nand U5548 (N_5548,N_5031,N_5373);
and U5549 (N_5549,N_5497,N_5104);
nand U5550 (N_5550,N_5376,N_5084);
xor U5551 (N_5551,N_5390,N_5082);
nor U5552 (N_5552,N_5371,N_5400);
nand U5553 (N_5553,N_5314,N_5479);
nor U5554 (N_5554,N_5232,N_5141);
nand U5555 (N_5555,N_5190,N_5060);
or U5556 (N_5556,N_5306,N_5396);
and U5557 (N_5557,N_5077,N_5230);
nand U5558 (N_5558,N_5381,N_5192);
or U5559 (N_5559,N_5378,N_5325);
or U5560 (N_5560,N_5301,N_5169);
nand U5561 (N_5561,N_5153,N_5240);
nor U5562 (N_5562,N_5460,N_5287);
or U5563 (N_5563,N_5252,N_5015);
or U5564 (N_5564,N_5265,N_5055);
or U5565 (N_5565,N_5043,N_5428);
and U5566 (N_5566,N_5246,N_5480);
xor U5567 (N_5567,N_5110,N_5154);
or U5568 (N_5568,N_5495,N_5383);
nor U5569 (N_5569,N_5231,N_5067);
or U5570 (N_5570,N_5000,N_5338);
or U5571 (N_5571,N_5163,N_5128);
or U5572 (N_5572,N_5354,N_5341);
nand U5573 (N_5573,N_5484,N_5222);
or U5574 (N_5574,N_5447,N_5477);
xnor U5575 (N_5575,N_5125,N_5365);
xnor U5576 (N_5576,N_5177,N_5027);
nand U5577 (N_5577,N_5144,N_5453);
nor U5578 (N_5578,N_5419,N_5118);
nor U5579 (N_5579,N_5263,N_5100);
xor U5580 (N_5580,N_5201,N_5471);
or U5581 (N_5581,N_5003,N_5002);
nor U5582 (N_5582,N_5127,N_5420);
nand U5583 (N_5583,N_5174,N_5449);
xor U5584 (N_5584,N_5021,N_5028);
xor U5585 (N_5585,N_5445,N_5088);
or U5586 (N_5586,N_5158,N_5342);
xor U5587 (N_5587,N_5005,N_5271);
nor U5588 (N_5588,N_5152,N_5042);
xor U5589 (N_5589,N_5437,N_5078);
and U5590 (N_5590,N_5045,N_5496);
or U5591 (N_5591,N_5366,N_5322);
or U5592 (N_5592,N_5391,N_5001);
nor U5593 (N_5593,N_5053,N_5036);
nor U5594 (N_5594,N_5243,N_5087);
and U5595 (N_5595,N_5037,N_5181);
xor U5596 (N_5596,N_5033,N_5147);
nand U5597 (N_5597,N_5269,N_5489);
and U5598 (N_5598,N_5283,N_5490);
nor U5599 (N_5599,N_5239,N_5412);
nor U5600 (N_5600,N_5051,N_5148);
and U5601 (N_5601,N_5047,N_5250);
nor U5602 (N_5602,N_5123,N_5094);
or U5603 (N_5603,N_5064,N_5443);
xnor U5604 (N_5604,N_5188,N_5399);
xnor U5605 (N_5605,N_5450,N_5071);
or U5606 (N_5606,N_5262,N_5436);
nor U5607 (N_5607,N_5249,N_5009);
or U5608 (N_5608,N_5208,N_5149);
and U5609 (N_5609,N_5070,N_5346);
xor U5610 (N_5610,N_5057,N_5370);
nand U5611 (N_5611,N_5498,N_5275);
or U5612 (N_5612,N_5395,N_5162);
and U5613 (N_5613,N_5401,N_5258);
nor U5614 (N_5614,N_5486,N_5284);
nor U5615 (N_5615,N_5062,N_5305);
and U5616 (N_5616,N_5303,N_5213);
nand U5617 (N_5617,N_5440,N_5124);
xnor U5618 (N_5618,N_5166,N_5417);
xor U5619 (N_5619,N_5034,N_5259);
nor U5620 (N_5620,N_5220,N_5494);
xor U5621 (N_5621,N_5274,N_5297);
and U5622 (N_5622,N_5332,N_5344);
nand U5623 (N_5623,N_5113,N_5288);
nand U5624 (N_5624,N_5013,N_5063);
nand U5625 (N_5625,N_5397,N_5309);
and U5626 (N_5626,N_5242,N_5093);
or U5627 (N_5627,N_5226,N_5159);
xnor U5628 (N_5628,N_5251,N_5382);
nand U5629 (N_5629,N_5423,N_5014);
xor U5630 (N_5630,N_5223,N_5135);
and U5631 (N_5631,N_5061,N_5377);
nor U5632 (N_5632,N_5069,N_5096);
xnor U5633 (N_5633,N_5029,N_5228);
or U5634 (N_5634,N_5372,N_5422);
xor U5635 (N_5635,N_5160,N_5469);
nor U5636 (N_5636,N_5134,N_5090);
nand U5637 (N_5637,N_5066,N_5293);
nand U5638 (N_5638,N_5461,N_5356);
or U5639 (N_5639,N_5241,N_5499);
nand U5640 (N_5640,N_5261,N_5433);
and U5641 (N_5641,N_5219,N_5481);
nand U5642 (N_5642,N_5394,N_5410);
and U5643 (N_5643,N_5464,N_5151);
or U5644 (N_5644,N_5402,N_5183);
nand U5645 (N_5645,N_5218,N_5318);
nand U5646 (N_5646,N_5289,N_5343);
xnor U5647 (N_5647,N_5363,N_5170);
or U5648 (N_5648,N_5326,N_5121);
xnor U5649 (N_5649,N_5431,N_5227);
nand U5650 (N_5650,N_5012,N_5337);
or U5651 (N_5651,N_5312,N_5238);
or U5652 (N_5652,N_5429,N_5083);
or U5653 (N_5653,N_5300,N_5080);
nand U5654 (N_5654,N_5054,N_5491);
and U5655 (N_5655,N_5133,N_5350);
xor U5656 (N_5656,N_5103,N_5438);
and U5657 (N_5657,N_5006,N_5175);
xnor U5658 (N_5658,N_5105,N_5074);
and U5659 (N_5659,N_5132,N_5268);
nand U5660 (N_5660,N_5330,N_5176);
nand U5661 (N_5661,N_5487,N_5292);
or U5662 (N_5662,N_5463,N_5385);
and U5663 (N_5663,N_5099,N_5277);
or U5664 (N_5664,N_5264,N_5386);
and U5665 (N_5665,N_5156,N_5018);
nand U5666 (N_5666,N_5179,N_5362);
or U5667 (N_5667,N_5323,N_5198);
or U5668 (N_5668,N_5046,N_5493);
nor U5669 (N_5669,N_5407,N_5424);
nand U5670 (N_5670,N_5004,N_5446);
or U5671 (N_5671,N_5278,N_5245);
nand U5672 (N_5672,N_5413,N_5454);
nor U5673 (N_5673,N_5473,N_5416);
and U5674 (N_5674,N_5168,N_5195);
nand U5675 (N_5675,N_5307,N_5345);
or U5676 (N_5676,N_5092,N_5296);
and U5677 (N_5677,N_5331,N_5313);
and U5678 (N_5678,N_5442,N_5038);
xor U5679 (N_5679,N_5221,N_5111);
nand U5680 (N_5680,N_5465,N_5024);
or U5681 (N_5681,N_5349,N_5089);
nand U5682 (N_5682,N_5091,N_5143);
nand U5683 (N_5683,N_5451,N_5415);
xnor U5684 (N_5684,N_5116,N_5270);
nor U5685 (N_5685,N_5072,N_5470);
nor U5686 (N_5686,N_5368,N_5418);
xor U5687 (N_5687,N_5369,N_5210);
and U5688 (N_5688,N_5020,N_5324);
nand U5689 (N_5689,N_5488,N_5117);
and U5690 (N_5690,N_5229,N_5076);
nor U5691 (N_5691,N_5310,N_5068);
or U5692 (N_5692,N_5459,N_5421);
or U5693 (N_5693,N_5236,N_5025);
and U5694 (N_5694,N_5276,N_5403);
nor U5695 (N_5695,N_5364,N_5200);
and U5696 (N_5696,N_5482,N_5164);
xnor U5697 (N_5697,N_5353,N_5032);
nand U5698 (N_5698,N_5468,N_5044);
nor U5699 (N_5699,N_5048,N_5191);
nand U5700 (N_5700,N_5207,N_5359);
or U5701 (N_5701,N_5348,N_5374);
nand U5702 (N_5702,N_5049,N_5167);
and U5703 (N_5703,N_5492,N_5073);
xnor U5704 (N_5704,N_5279,N_5205);
and U5705 (N_5705,N_5140,N_5448);
nand U5706 (N_5706,N_5197,N_5233);
nand U5707 (N_5707,N_5165,N_5186);
and U5708 (N_5708,N_5360,N_5315);
xnor U5709 (N_5709,N_5206,N_5065);
and U5710 (N_5710,N_5472,N_5466);
nand U5711 (N_5711,N_5329,N_5056);
xor U5712 (N_5712,N_5204,N_5130);
nor U5713 (N_5713,N_5189,N_5351);
nand U5714 (N_5714,N_5414,N_5387);
and U5715 (N_5715,N_5145,N_5455);
nand U5716 (N_5716,N_5406,N_5011);
xor U5717 (N_5717,N_5282,N_5476);
xnor U5718 (N_5718,N_5225,N_5409);
nand U5719 (N_5719,N_5452,N_5237);
and U5720 (N_5720,N_5008,N_5050);
nor U5721 (N_5721,N_5007,N_5427);
or U5722 (N_5722,N_5122,N_5101);
and U5723 (N_5723,N_5244,N_5017);
xnor U5724 (N_5724,N_5209,N_5254);
xor U5725 (N_5725,N_5115,N_5405);
or U5726 (N_5726,N_5212,N_5108);
and U5727 (N_5727,N_5041,N_5456);
nor U5728 (N_5728,N_5107,N_5483);
and U5729 (N_5729,N_5266,N_5434);
or U5730 (N_5730,N_5039,N_5171);
or U5731 (N_5731,N_5079,N_5131);
nor U5732 (N_5732,N_5392,N_5194);
and U5733 (N_5733,N_5328,N_5256);
and U5734 (N_5734,N_5030,N_5361);
xor U5735 (N_5735,N_5157,N_5290);
or U5736 (N_5736,N_5462,N_5202);
xnor U5737 (N_5737,N_5146,N_5304);
and U5738 (N_5738,N_5182,N_5273);
or U5739 (N_5739,N_5339,N_5408);
and U5740 (N_5740,N_5272,N_5114);
or U5741 (N_5741,N_5095,N_5335);
or U5742 (N_5742,N_5398,N_5474);
and U5743 (N_5743,N_5215,N_5444);
or U5744 (N_5744,N_5478,N_5097);
or U5745 (N_5745,N_5457,N_5085);
nand U5746 (N_5746,N_5327,N_5426);
xor U5747 (N_5747,N_5257,N_5086);
xor U5748 (N_5748,N_5411,N_5347);
xnor U5749 (N_5749,N_5136,N_5308);
nor U5750 (N_5750,N_5224,N_5223);
or U5751 (N_5751,N_5037,N_5403);
nand U5752 (N_5752,N_5133,N_5326);
or U5753 (N_5753,N_5034,N_5250);
or U5754 (N_5754,N_5396,N_5436);
nand U5755 (N_5755,N_5150,N_5328);
xor U5756 (N_5756,N_5151,N_5433);
or U5757 (N_5757,N_5033,N_5159);
xor U5758 (N_5758,N_5174,N_5137);
and U5759 (N_5759,N_5212,N_5036);
or U5760 (N_5760,N_5440,N_5326);
or U5761 (N_5761,N_5011,N_5322);
nor U5762 (N_5762,N_5099,N_5327);
and U5763 (N_5763,N_5348,N_5017);
nor U5764 (N_5764,N_5184,N_5109);
or U5765 (N_5765,N_5479,N_5473);
xor U5766 (N_5766,N_5238,N_5131);
or U5767 (N_5767,N_5359,N_5146);
nand U5768 (N_5768,N_5092,N_5009);
xnor U5769 (N_5769,N_5362,N_5350);
or U5770 (N_5770,N_5285,N_5310);
nor U5771 (N_5771,N_5209,N_5427);
or U5772 (N_5772,N_5132,N_5059);
xor U5773 (N_5773,N_5353,N_5134);
xor U5774 (N_5774,N_5378,N_5142);
xor U5775 (N_5775,N_5021,N_5265);
nor U5776 (N_5776,N_5103,N_5414);
or U5777 (N_5777,N_5069,N_5339);
xnor U5778 (N_5778,N_5430,N_5075);
nand U5779 (N_5779,N_5233,N_5072);
or U5780 (N_5780,N_5422,N_5047);
nor U5781 (N_5781,N_5268,N_5113);
or U5782 (N_5782,N_5101,N_5491);
xnor U5783 (N_5783,N_5266,N_5411);
xor U5784 (N_5784,N_5122,N_5011);
or U5785 (N_5785,N_5045,N_5289);
xor U5786 (N_5786,N_5082,N_5194);
and U5787 (N_5787,N_5325,N_5120);
nand U5788 (N_5788,N_5176,N_5320);
and U5789 (N_5789,N_5314,N_5156);
or U5790 (N_5790,N_5002,N_5161);
or U5791 (N_5791,N_5378,N_5206);
nor U5792 (N_5792,N_5184,N_5261);
xor U5793 (N_5793,N_5089,N_5231);
and U5794 (N_5794,N_5236,N_5438);
nor U5795 (N_5795,N_5442,N_5052);
and U5796 (N_5796,N_5087,N_5153);
and U5797 (N_5797,N_5075,N_5268);
xnor U5798 (N_5798,N_5406,N_5145);
or U5799 (N_5799,N_5184,N_5377);
or U5800 (N_5800,N_5095,N_5154);
xnor U5801 (N_5801,N_5402,N_5005);
nand U5802 (N_5802,N_5115,N_5359);
nand U5803 (N_5803,N_5137,N_5474);
or U5804 (N_5804,N_5497,N_5077);
xor U5805 (N_5805,N_5455,N_5487);
nand U5806 (N_5806,N_5230,N_5496);
nand U5807 (N_5807,N_5434,N_5234);
nor U5808 (N_5808,N_5266,N_5033);
nand U5809 (N_5809,N_5157,N_5229);
xor U5810 (N_5810,N_5448,N_5282);
and U5811 (N_5811,N_5380,N_5496);
and U5812 (N_5812,N_5493,N_5084);
and U5813 (N_5813,N_5020,N_5337);
or U5814 (N_5814,N_5315,N_5366);
xor U5815 (N_5815,N_5041,N_5066);
xor U5816 (N_5816,N_5293,N_5363);
nor U5817 (N_5817,N_5207,N_5187);
nor U5818 (N_5818,N_5286,N_5460);
and U5819 (N_5819,N_5220,N_5474);
or U5820 (N_5820,N_5322,N_5087);
nand U5821 (N_5821,N_5044,N_5266);
nand U5822 (N_5822,N_5442,N_5153);
or U5823 (N_5823,N_5269,N_5405);
xnor U5824 (N_5824,N_5063,N_5426);
nor U5825 (N_5825,N_5304,N_5052);
xnor U5826 (N_5826,N_5486,N_5375);
nand U5827 (N_5827,N_5125,N_5072);
nand U5828 (N_5828,N_5363,N_5320);
or U5829 (N_5829,N_5448,N_5160);
nand U5830 (N_5830,N_5149,N_5304);
or U5831 (N_5831,N_5391,N_5158);
or U5832 (N_5832,N_5418,N_5107);
and U5833 (N_5833,N_5286,N_5062);
or U5834 (N_5834,N_5258,N_5112);
or U5835 (N_5835,N_5376,N_5105);
nor U5836 (N_5836,N_5166,N_5268);
nor U5837 (N_5837,N_5299,N_5354);
xnor U5838 (N_5838,N_5428,N_5170);
xnor U5839 (N_5839,N_5149,N_5336);
nor U5840 (N_5840,N_5099,N_5471);
nand U5841 (N_5841,N_5186,N_5437);
nor U5842 (N_5842,N_5232,N_5413);
and U5843 (N_5843,N_5450,N_5124);
nand U5844 (N_5844,N_5378,N_5365);
or U5845 (N_5845,N_5394,N_5184);
nand U5846 (N_5846,N_5365,N_5296);
and U5847 (N_5847,N_5354,N_5315);
nand U5848 (N_5848,N_5475,N_5103);
or U5849 (N_5849,N_5365,N_5255);
nor U5850 (N_5850,N_5193,N_5126);
nand U5851 (N_5851,N_5098,N_5139);
nor U5852 (N_5852,N_5229,N_5066);
or U5853 (N_5853,N_5021,N_5258);
xnor U5854 (N_5854,N_5368,N_5413);
and U5855 (N_5855,N_5119,N_5384);
nor U5856 (N_5856,N_5079,N_5239);
nand U5857 (N_5857,N_5183,N_5107);
and U5858 (N_5858,N_5360,N_5100);
nor U5859 (N_5859,N_5352,N_5303);
nand U5860 (N_5860,N_5267,N_5384);
or U5861 (N_5861,N_5449,N_5280);
nor U5862 (N_5862,N_5159,N_5301);
and U5863 (N_5863,N_5120,N_5278);
nand U5864 (N_5864,N_5396,N_5162);
nor U5865 (N_5865,N_5335,N_5161);
nor U5866 (N_5866,N_5455,N_5222);
xnor U5867 (N_5867,N_5000,N_5376);
xnor U5868 (N_5868,N_5246,N_5456);
nand U5869 (N_5869,N_5342,N_5474);
or U5870 (N_5870,N_5255,N_5445);
nor U5871 (N_5871,N_5075,N_5067);
xnor U5872 (N_5872,N_5006,N_5200);
nand U5873 (N_5873,N_5181,N_5358);
and U5874 (N_5874,N_5255,N_5078);
xor U5875 (N_5875,N_5411,N_5157);
nor U5876 (N_5876,N_5154,N_5099);
and U5877 (N_5877,N_5076,N_5289);
nand U5878 (N_5878,N_5476,N_5494);
or U5879 (N_5879,N_5383,N_5231);
or U5880 (N_5880,N_5263,N_5495);
or U5881 (N_5881,N_5134,N_5166);
xnor U5882 (N_5882,N_5426,N_5199);
nor U5883 (N_5883,N_5471,N_5029);
and U5884 (N_5884,N_5420,N_5022);
nand U5885 (N_5885,N_5114,N_5479);
xnor U5886 (N_5886,N_5497,N_5305);
nor U5887 (N_5887,N_5098,N_5191);
or U5888 (N_5888,N_5117,N_5386);
xnor U5889 (N_5889,N_5032,N_5266);
and U5890 (N_5890,N_5273,N_5079);
xnor U5891 (N_5891,N_5319,N_5339);
nand U5892 (N_5892,N_5386,N_5000);
nor U5893 (N_5893,N_5147,N_5023);
nand U5894 (N_5894,N_5194,N_5342);
xnor U5895 (N_5895,N_5381,N_5070);
and U5896 (N_5896,N_5117,N_5044);
nor U5897 (N_5897,N_5000,N_5100);
or U5898 (N_5898,N_5319,N_5007);
nand U5899 (N_5899,N_5023,N_5424);
nor U5900 (N_5900,N_5193,N_5194);
nor U5901 (N_5901,N_5403,N_5484);
xor U5902 (N_5902,N_5436,N_5473);
nor U5903 (N_5903,N_5230,N_5377);
or U5904 (N_5904,N_5076,N_5198);
nand U5905 (N_5905,N_5442,N_5454);
nor U5906 (N_5906,N_5198,N_5457);
xnor U5907 (N_5907,N_5341,N_5191);
nand U5908 (N_5908,N_5456,N_5201);
nor U5909 (N_5909,N_5338,N_5488);
and U5910 (N_5910,N_5082,N_5422);
nor U5911 (N_5911,N_5281,N_5156);
or U5912 (N_5912,N_5064,N_5029);
nor U5913 (N_5913,N_5024,N_5358);
nor U5914 (N_5914,N_5390,N_5283);
or U5915 (N_5915,N_5290,N_5111);
xnor U5916 (N_5916,N_5327,N_5464);
nand U5917 (N_5917,N_5142,N_5224);
xnor U5918 (N_5918,N_5315,N_5110);
or U5919 (N_5919,N_5321,N_5076);
or U5920 (N_5920,N_5245,N_5189);
nand U5921 (N_5921,N_5476,N_5239);
and U5922 (N_5922,N_5118,N_5490);
xnor U5923 (N_5923,N_5425,N_5397);
xnor U5924 (N_5924,N_5336,N_5399);
xor U5925 (N_5925,N_5221,N_5401);
or U5926 (N_5926,N_5026,N_5413);
and U5927 (N_5927,N_5432,N_5146);
nand U5928 (N_5928,N_5326,N_5024);
or U5929 (N_5929,N_5377,N_5191);
xnor U5930 (N_5930,N_5291,N_5155);
nor U5931 (N_5931,N_5135,N_5264);
nand U5932 (N_5932,N_5164,N_5072);
or U5933 (N_5933,N_5043,N_5480);
and U5934 (N_5934,N_5208,N_5292);
and U5935 (N_5935,N_5314,N_5110);
or U5936 (N_5936,N_5144,N_5428);
nand U5937 (N_5937,N_5010,N_5112);
or U5938 (N_5938,N_5288,N_5056);
and U5939 (N_5939,N_5262,N_5015);
nor U5940 (N_5940,N_5177,N_5179);
and U5941 (N_5941,N_5038,N_5469);
and U5942 (N_5942,N_5329,N_5064);
nand U5943 (N_5943,N_5209,N_5285);
xor U5944 (N_5944,N_5326,N_5037);
or U5945 (N_5945,N_5393,N_5207);
and U5946 (N_5946,N_5023,N_5426);
nand U5947 (N_5947,N_5198,N_5310);
nor U5948 (N_5948,N_5334,N_5378);
nor U5949 (N_5949,N_5139,N_5362);
xor U5950 (N_5950,N_5222,N_5378);
nor U5951 (N_5951,N_5331,N_5121);
and U5952 (N_5952,N_5401,N_5300);
xor U5953 (N_5953,N_5040,N_5356);
and U5954 (N_5954,N_5100,N_5080);
or U5955 (N_5955,N_5485,N_5086);
xnor U5956 (N_5956,N_5485,N_5278);
nor U5957 (N_5957,N_5280,N_5057);
or U5958 (N_5958,N_5465,N_5044);
and U5959 (N_5959,N_5028,N_5327);
xor U5960 (N_5960,N_5083,N_5412);
or U5961 (N_5961,N_5000,N_5244);
nand U5962 (N_5962,N_5057,N_5401);
and U5963 (N_5963,N_5419,N_5450);
nor U5964 (N_5964,N_5298,N_5393);
nor U5965 (N_5965,N_5209,N_5477);
and U5966 (N_5966,N_5240,N_5064);
or U5967 (N_5967,N_5245,N_5466);
xor U5968 (N_5968,N_5206,N_5490);
nand U5969 (N_5969,N_5203,N_5272);
or U5970 (N_5970,N_5156,N_5487);
nand U5971 (N_5971,N_5007,N_5264);
xor U5972 (N_5972,N_5043,N_5170);
nor U5973 (N_5973,N_5475,N_5420);
nand U5974 (N_5974,N_5448,N_5016);
and U5975 (N_5975,N_5424,N_5210);
nor U5976 (N_5976,N_5123,N_5159);
or U5977 (N_5977,N_5152,N_5155);
xnor U5978 (N_5978,N_5052,N_5084);
xor U5979 (N_5979,N_5465,N_5236);
and U5980 (N_5980,N_5254,N_5176);
and U5981 (N_5981,N_5220,N_5452);
and U5982 (N_5982,N_5313,N_5238);
and U5983 (N_5983,N_5164,N_5272);
xnor U5984 (N_5984,N_5299,N_5139);
or U5985 (N_5985,N_5416,N_5061);
and U5986 (N_5986,N_5483,N_5410);
or U5987 (N_5987,N_5049,N_5109);
nand U5988 (N_5988,N_5327,N_5298);
nand U5989 (N_5989,N_5444,N_5322);
or U5990 (N_5990,N_5170,N_5427);
xnor U5991 (N_5991,N_5124,N_5496);
or U5992 (N_5992,N_5302,N_5333);
or U5993 (N_5993,N_5203,N_5230);
and U5994 (N_5994,N_5214,N_5265);
nand U5995 (N_5995,N_5162,N_5046);
and U5996 (N_5996,N_5237,N_5356);
nand U5997 (N_5997,N_5491,N_5313);
nand U5998 (N_5998,N_5038,N_5382);
xnor U5999 (N_5999,N_5014,N_5137);
nor U6000 (N_6000,N_5666,N_5849);
and U6001 (N_6001,N_5521,N_5805);
and U6002 (N_6002,N_5946,N_5551);
nand U6003 (N_6003,N_5510,N_5619);
xnor U6004 (N_6004,N_5823,N_5637);
and U6005 (N_6005,N_5999,N_5958);
and U6006 (N_6006,N_5871,N_5866);
nor U6007 (N_6007,N_5682,N_5635);
or U6008 (N_6008,N_5664,N_5741);
nand U6009 (N_6009,N_5624,N_5723);
nand U6010 (N_6010,N_5712,N_5868);
and U6011 (N_6011,N_5529,N_5651);
and U6012 (N_6012,N_5766,N_5612);
and U6013 (N_6013,N_5901,N_5907);
xnor U6014 (N_6014,N_5675,N_5532);
xnor U6015 (N_6015,N_5998,N_5967);
nor U6016 (N_6016,N_5520,N_5772);
nand U6017 (N_6017,N_5530,N_5860);
and U6018 (N_6018,N_5917,N_5523);
nor U6019 (N_6019,N_5894,N_5918);
and U6020 (N_6020,N_5945,N_5938);
nor U6021 (N_6021,N_5586,N_5813);
or U6022 (N_6022,N_5955,N_5507);
and U6023 (N_6023,N_5748,N_5736);
or U6024 (N_6024,N_5626,N_5591);
xnor U6025 (N_6025,N_5862,N_5522);
or U6026 (N_6026,N_5787,N_5713);
nor U6027 (N_6027,N_5798,N_5926);
nor U6028 (N_6028,N_5714,N_5954);
nand U6029 (N_6029,N_5639,N_5581);
xnor U6030 (N_6030,N_5789,N_5982);
or U6031 (N_6031,N_5590,N_5597);
or U6032 (N_6032,N_5824,N_5984);
nand U6033 (N_6033,N_5972,N_5891);
nor U6034 (N_6034,N_5928,N_5839);
and U6035 (N_6035,N_5807,N_5568);
nand U6036 (N_6036,N_5986,N_5742);
xnor U6037 (N_6037,N_5773,N_5977);
nor U6038 (N_6038,N_5856,N_5820);
nand U6039 (N_6039,N_5662,N_5983);
nor U6040 (N_6040,N_5631,N_5923);
nor U6041 (N_6041,N_5659,N_5501);
nor U6042 (N_6042,N_5847,N_5557);
and U6043 (N_6043,N_5916,N_5774);
nor U6044 (N_6044,N_5504,N_5726);
or U6045 (N_6045,N_5873,N_5980);
or U6046 (N_6046,N_5806,N_5692);
or U6047 (N_6047,N_5758,N_5780);
and U6048 (N_6048,N_5660,N_5796);
nor U6049 (N_6049,N_5833,N_5888);
or U6050 (N_6050,N_5710,N_5690);
and U6051 (N_6051,N_5695,N_5782);
nand U6052 (N_6052,N_5625,N_5815);
nand U6053 (N_6053,N_5562,N_5699);
and U6054 (N_6054,N_5587,N_5864);
nand U6055 (N_6055,N_5895,N_5846);
nor U6056 (N_6056,N_5852,N_5623);
nor U6057 (N_6057,N_5908,N_5640);
xnor U6058 (N_6058,N_5605,N_5974);
or U6059 (N_6059,N_5575,N_5953);
and U6060 (N_6060,N_5589,N_5519);
or U6061 (N_6061,N_5584,N_5733);
and U6062 (N_6062,N_5697,N_5865);
and U6063 (N_6063,N_5727,N_5768);
nand U6064 (N_6064,N_5564,N_5831);
and U6065 (N_6065,N_5512,N_5711);
and U6066 (N_6066,N_5859,N_5598);
nand U6067 (N_6067,N_5737,N_5593);
and U6068 (N_6068,N_5744,N_5722);
nand U6069 (N_6069,N_5904,N_5960);
nand U6070 (N_6070,N_5541,N_5817);
and U6071 (N_6071,N_5990,N_5648);
or U6072 (N_6072,N_5686,N_5875);
xnor U6073 (N_6073,N_5542,N_5554);
xor U6074 (N_6074,N_5604,N_5611);
xor U6075 (N_6075,N_5838,N_5616);
or U6076 (N_6076,N_5992,N_5567);
and U6077 (N_6077,N_5534,N_5845);
nand U6078 (N_6078,N_5515,N_5588);
nand U6079 (N_6079,N_5655,N_5968);
and U6080 (N_6080,N_5663,N_5889);
nand U6081 (N_6081,N_5751,N_5665);
nand U6082 (N_6082,N_5931,N_5786);
or U6083 (N_6083,N_5776,N_5957);
nor U6084 (N_6084,N_5518,N_5566);
and U6085 (N_6085,N_5580,N_5544);
xor U6086 (N_6086,N_5652,N_5969);
or U6087 (N_6087,N_5985,N_5964);
nor U6088 (N_6088,N_5735,N_5578);
xnor U6089 (N_6089,N_5514,N_5739);
xor U6090 (N_6090,N_5851,N_5618);
nand U6091 (N_6091,N_5854,N_5696);
and U6092 (N_6092,N_5558,N_5561);
nand U6093 (N_6093,N_5730,N_5821);
or U6094 (N_6094,N_5935,N_5853);
nor U6095 (N_6095,N_5775,N_5961);
and U6096 (N_6096,N_5784,N_5996);
and U6097 (N_6097,N_5747,N_5676);
xnor U6098 (N_6098,N_5988,N_5814);
xnor U6099 (N_6099,N_5533,N_5850);
or U6100 (N_6100,N_5603,N_5654);
nor U6101 (N_6101,N_5799,N_5677);
and U6102 (N_6102,N_5535,N_5565);
nand U6103 (N_6103,N_5756,N_5914);
and U6104 (N_6104,N_5753,N_5767);
xor U6105 (N_6105,N_5740,N_5777);
nand U6106 (N_6106,N_5678,N_5702);
and U6107 (N_6107,N_5927,N_5634);
xnor U6108 (N_6108,N_5876,N_5505);
and U6109 (N_6109,N_5645,N_5606);
or U6110 (N_6110,N_5620,N_5790);
nand U6111 (N_6111,N_5802,N_5738);
nand U6112 (N_6112,N_5915,N_5912);
and U6113 (N_6113,N_5900,N_5704);
xor U6114 (N_6114,N_5638,N_5609);
xor U6115 (N_6115,N_5684,N_5718);
xnor U6116 (N_6116,N_5801,N_5804);
or U6117 (N_6117,N_5617,N_5808);
and U6118 (N_6118,N_5538,N_5970);
nor U6119 (N_6119,N_5668,N_5810);
and U6120 (N_6120,N_5720,N_5670);
and U6121 (N_6121,N_5880,N_5658);
nor U6122 (N_6122,N_5552,N_5641);
xnor U6123 (N_6123,N_5537,N_5791);
xor U6124 (N_6124,N_5759,N_5878);
nor U6125 (N_6125,N_5771,N_5933);
or U6126 (N_6126,N_5650,N_5882);
xnor U6127 (N_6127,N_5516,N_5672);
nor U6128 (N_6128,N_5921,N_5800);
xor U6129 (N_6129,N_5649,N_5947);
and U6130 (N_6130,N_5600,N_5576);
xor U6131 (N_6131,N_5896,N_5841);
nand U6132 (N_6132,N_5949,N_5979);
and U6133 (N_6133,N_5531,N_5994);
nor U6134 (N_6134,N_5610,N_5929);
or U6135 (N_6135,N_5981,N_5892);
xor U6136 (N_6136,N_5940,N_5596);
nor U6137 (N_6137,N_5646,N_5886);
or U6138 (N_6138,N_5903,N_5779);
and U6139 (N_6139,N_5539,N_5572);
or U6140 (N_6140,N_5976,N_5936);
nor U6141 (N_6141,N_5698,N_5577);
and U6142 (N_6142,N_5585,N_5797);
and U6143 (N_6143,N_5794,N_5528);
or U6144 (N_6144,N_5559,N_5897);
nor U6145 (N_6145,N_5685,N_5669);
or U6146 (N_6146,N_5653,N_5822);
nor U6147 (N_6147,N_5793,N_5869);
xnor U6148 (N_6148,N_5509,N_5836);
xor U6149 (N_6149,N_5879,N_5540);
nand U6150 (N_6150,N_5781,N_5819);
xnor U6151 (N_6151,N_5546,N_5837);
and U6152 (N_6152,N_5829,N_5573);
nand U6153 (N_6153,N_5622,N_5890);
or U6154 (N_6154,N_5857,N_5700);
xnor U6155 (N_6155,N_5732,N_5956);
nand U6156 (N_6156,N_5855,N_5614);
xnor U6157 (N_6157,N_5687,N_5762);
nor U6158 (N_6158,N_5693,N_5536);
nor U6159 (N_6159,N_5765,N_5569);
nor U6160 (N_6160,N_5863,N_5592);
and U6161 (N_6161,N_5830,N_5508);
and U6162 (N_6162,N_5842,N_5749);
and U6163 (N_6163,N_5703,N_5832);
xnor U6164 (N_6164,N_5525,N_5524);
and U6165 (N_6165,N_5870,N_5987);
and U6166 (N_6166,N_5526,N_5919);
nand U6167 (N_6167,N_5673,N_5601);
or U6168 (N_6168,N_5694,N_5997);
xnor U6169 (N_6169,N_5574,N_5769);
nand U6170 (N_6170,N_5995,N_5527);
nor U6171 (N_6171,N_5607,N_5761);
nand U6172 (N_6172,N_5770,N_5834);
xor U6173 (N_6173,N_5642,N_5632);
nand U6174 (N_6174,N_5731,N_5547);
and U6175 (N_6175,N_5543,N_5502);
xnor U6176 (N_6176,N_5719,N_5848);
nand U6177 (N_6177,N_5689,N_5911);
nand U6178 (N_6178,N_5555,N_5978);
nor U6179 (N_6179,N_5734,N_5828);
nor U6180 (N_6180,N_5975,N_5656);
or U6181 (N_6181,N_5725,N_5630);
xnor U6182 (N_6182,N_5881,N_5884);
xnor U6183 (N_6183,N_5706,N_5715);
nand U6184 (N_6184,N_5973,N_5583);
xor U6185 (N_6185,N_5550,N_5825);
or U6186 (N_6186,N_5883,N_5743);
and U6187 (N_6187,N_5571,N_5991);
or U6188 (N_6188,N_5840,N_5595);
and U6189 (N_6189,N_5948,N_5843);
xor U6190 (N_6190,N_5877,N_5755);
or U6191 (N_6191,N_5708,N_5844);
nor U6192 (N_6192,N_5922,N_5760);
nor U6193 (N_6193,N_5644,N_5657);
or U6194 (N_6194,N_5966,N_5925);
xor U6195 (N_6195,N_5788,N_5963);
nor U6196 (N_6196,N_5628,N_5671);
nor U6197 (N_6197,N_5680,N_5709);
nand U6198 (N_6198,N_5661,N_5809);
or U6199 (N_6199,N_5965,N_5826);
nand U6200 (N_6200,N_5939,N_5941);
nor U6201 (N_6201,N_5545,N_5959);
and U6202 (N_6202,N_5989,N_5679);
nor U6203 (N_6203,N_5707,N_5615);
nand U6204 (N_6204,N_5548,N_5563);
xnor U6205 (N_6205,N_5885,N_5716);
nor U6206 (N_6206,N_5930,N_5899);
and U6207 (N_6207,N_5728,N_5944);
nor U6208 (N_6208,N_5792,N_5902);
and U6209 (N_6209,N_5754,N_5570);
and U6210 (N_6210,N_5909,N_5785);
and U6211 (N_6211,N_5803,N_5910);
nand U6212 (N_6212,N_5783,N_5745);
and U6213 (N_6213,N_5934,N_5887);
and U6214 (N_6214,N_5874,N_5503);
nor U6215 (N_6215,N_5511,N_5691);
and U6216 (N_6216,N_5681,N_5905);
or U6217 (N_6217,N_5608,N_5674);
and U6218 (N_6218,N_5942,N_5560);
nor U6219 (N_6219,N_5932,N_5913);
xnor U6220 (N_6220,N_5627,N_5513);
and U6221 (N_6221,N_5993,N_5517);
or U6222 (N_6222,N_5861,N_5920);
xor U6223 (N_6223,N_5688,N_5721);
nand U6224 (N_6224,N_5724,N_5643);
xor U6225 (N_6225,N_5579,N_5717);
xor U6226 (N_6226,N_5613,N_5633);
or U6227 (N_6227,N_5924,N_5667);
or U6228 (N_6228,N_5867,N_5621);
nand U6229 (N_6229,N_5906,N_5962);
nor U6230 (N_6230,N_5898,N_5683);
and U6231 (N_6231,N_5556,N_5858);
nand U6232 (N_6232,N_5818,N_5835);
and U6233 (N_6233,N_5778,N_5750);
nand U6234 (N_6234,N_5553,N_5701);
nor U6235 (N_6235,N_5943,N_5971);
xnor U6236 (N_6236,N_5647,N_5599);
nand U6237 (N_6237,N_5549,N_5795);
xor U6238 (N_6238,N_5763,N_5827);
and U6239 (N_6239,N_5746,N_5764);
nor U6240 (N_6240,N_5893,N_5594);
or U6241 (N_6241,N_5812,N_5952);
nand U6242 (N_6242,N_5636,N_5602);
nand U6243 (N_6243,N_5937,N_5705);
xnor U6244 (N_6244,N_5752,N_5757);
and U6245 (N_6245,N_5582,N_5816);
or U6246 (N_6246,N_5629,N_5811);
nand U6247 (N_6247,N_5951,N_5872);
or U6248 (N_6248,N_5950,N_5729);
nor U6249 (N_6249,N_5500,N_5506);
nand U6250 (N_6250,N_5663,N_5985);
nand U6251 (N_6251,N_5799,N_5696);
or U6252 (N_6252,N_5783,N_5763);
xnor U6253 (N_6253,N_5571,N_5833);
and U6254 (N_6254,N_5661,N_5995);
nor U6255 (N_6255,N_5527,N_5621);
or U6256 (N_6256,N_5963,N_5581);
or U6257 (N_6257,N_5585,N_5999);
and U6258 (N_6258,N_5643,N_5516);
xor U6259 (N_6259,N_5639,N_5908);
xnor U6260 (N_6260,N_5916,N_5687);
nand U6261 (N_6261,N_5576,N_5603);
nand U6262 (N_6262,N_5524,N_5943);
and U6263 (N_6263,N_5896,N_5936);
and U6264 (N_6264,N_5703,N_5547);
nor U6265 (N_6265,N_5874,N_5901);
xnor U6266 (N_6266,N_5935,N_5844);
nor U6267 (N_6267,N_5907,N_5717);
xor U6268 (N_6268,N_5668,N_5817);
nor U6269 (N_6269,N_5680,N_5794);
and U6270 (N_6270,N_5510,N_5553);
nand U6271 (N_6271,N_5912,N_5901);
and U6272 (N_6272,N_5970,N_5686);
nor U6273 (N_6273,N_5536,N_5675);
nand U6274 (N_6274,N_5513,N_5800);
and U6275 (N_6275,N_5993,N_5607);
or U6276 (N_6276,N_5608,N_5872);
and U6277 (N_6277,N_5649,N_5617);
nand U6278 (N_6278,N_5524,N_5710);
and U6279 (N_6279,N_5766,N_5651);
xor U6280 (N_6280,N_5903,N_5950);
and U6281 (N_6281,N_5603,N_5822);
xor U6282 (N_6282,N_5824,N_5583);
xor U6283 (N_6283,N_5977,N_5670);
and U6284 (N_6284,N_5657,N_5852);
xor U6285 (N_6285,N_5826,N_5747);
and U6286 (N_6286,N_5971,N_5700);
and U6287 (N_6287,N_5686,N_5800);
nand U6288 (N_6288,N_5647,N_5516);
xor U6289 (N_6289,N_5893,N_5852);
xor U6290 (N_6290,N_5585,N_5965);
xnor U6291 (N_6291,N_5677,N_5548);
or U6292 (N_6292,N_5973,N_5877);
xor U6293 (N_6293,N_5817,N_5910);
xnor U6294 (N_6294,N_5794,N_5778);
nor U6295 (N_6295,N_5788,N_5965);
nand U6296 (N_6296,N_5860,N_5901);
nand U6297 (N_6297,N_5716,N_5898);
nor U6298 (N_6298,N_5583,N_5666);
xnor U6299 (N_6299,N_5649,N_5682);
xor U6300 (N_6300,N_5707,N_5934);
nor U6301 (N_6301,N_5708,N_5797);
or U6302 (N_6302,N_5955,N_5636);
or U6303 (N_6303,N_5812,N_5625);
xnor U6304 (N_6304,N_5872,N_5635);
xor U6305 (N_6305,N_5976,N_5586);
xor U6306 (N_6306,N_5737,N_5503);
nor U6307 (N_6307,N_5818,N_5790);
and U6308 (N_6308,N_5889,N_5677);
and U6309 (N_6309,N_5622,N_5873);
and U6310 (N_6310,N_5545,N_5834);
or U6311 (N_6311,N_5919,N_5954);
or U6312 (N_6312,N_5720,N_5815);
xnor U6313 (N_6313,N_5510,N_5673);
and U6314 (N_6314,N_5971,N_5797);
nand U6315 (N_6315,N_5657,N_5760);
and U6316 (N_6316,N_5879,N_5675);
nor U6317 (N_6317,N_5973,N_5702);
xnor U6318 (N_6318,N_5665,N_5670);
nor U6319 (N_6319,N_5585,N_5543);
nand U6320 (N_6320,N_5582,N_5590);
nand U6321 (N_6321,N_5557,N_5785);
nor U6322 (N_6322,N_5943,N_5919);
xor U6323 (N_6323,N_5624,N_5625);
or U6324 (N_6324,N_5916,N_5527);
nand U6325 (N_6325,N_5667,N_5978);
or U6326 (N_6326,N_5630,N_5621);
xnor U6327 (N_6327,N_5727,N_5859);
and U6328 (N_6328,N_5652,N_5565);
and U6329 (N_6329,N_5857,N_5710);
and U6330 (N_6330,N_5533,N_5663);
or U6331 (N_6331,N_5866,N_5742);
nand U6332 (N_6332,N_5997,N_5531);
nor U6333 (N_6333,N_5675,N_5821);
xnor U6334 (N_6334,N_5639,N_5932);
nor U6335 (N_6335,N_5846,N_5857);
nor U6336 (N_6336,N_5966,N_5993);
nor U6337 (N_6337,N_5675,N_5565);
or U6338 (N_6338,N_5697,N_5854);
nor U6339 (N_6339,N_5710,N_5887);
nand U6340 (N_6340,N_5594,N_5663);
nand U6341 (N_6341,N_5704,N_5664);
nor U6342 (N_6342,N_5561,N_5586);
or U6343 (N_6343,N_5546,N_5770);
nand U6344 (N_6344,N_5990,N_5885);
nor U6345 (N_6345,N_5896,N_5645);
and U6346 (N_6346,N_5734,N_5706);
xor U6347 (N_6347,N_5927,N_5868);
xnor U6348 (N_6348,N_5791,N_5637);
nor U6349 (N_6349,N_5820,N_5573);
nor U6350 (N_6350,N_5558,N_5906);
and U6351 (N_6351,N_5830,N_5815);
or U6352 (N_6352,N_5646,N_5706);
or U6353 (N_6353,N_5610,N_5918);
or U6354 (N_6354,N_5689,N_5961);
and U6355 (N_6355,N_5635,N_5809);
and U6356 (N_6356,N_5583,N_5674);
xnor U6357 (N_6357,N_5500,N_5564);
nor U6358 (N_6358,N_5640,N_5975);
xor U6359 (N_6359,N_5839,N_5555);
and U6360 (N_6360,N_5548,N_5573);
or U6361 (N_6361,N_5875,N_5729);
and U6362 (N_6362,N_5848,N_5977);
xnor U6363 (N_6363,N_5974,N_5764);
and U6364 (N_6364,N_5541,N_5537);
or U6365 (N_6365,N_5922,N_5972);
nand U6366 (N_6366,N_5677,N_5744);
nor U6367 (N_6367,N_5877,N_5520);
and U6368 (N_6368,N_5624,N_5720);
and U6369 (N_6369,N_5857,N_5691);
and U6370 (N_6370,N_5893,N_5910);
nor U6371 (N_6371,N_5822,N_5507);
xnor U6372 (N_6372,N_5827,N_5912);
nor U6373 (N_6373,N_5663,N_5591);
nand U6374 (N_6374,N_5904,N_5655);
xnor U6375 (N_6375,N_5823,N_5913);
nor U6376 (N_6376,N_5936,N_5529);
nor U6377 (N_6377,N_5815,N_5932);
and U6378 (N_6378,N_5741,N_5774);
or U6379 (N_6379,N_5908,N_5571);
nand U6380 (N_6380,N_5542,N_5603);
or U6381 (N_6381,N_5995,N_5679);
or U6382 (N_6382,N_5575,N_5742);
xnor U6383 (N_6383,N_5924,N_5747);
or U6384 (N_6384,N_5539,N_5577);
or U6385 (N_6385,N_5505,N_5742);
nor U6386 (N_6386,N_5555,N_5742);
and U6387 (N_6387,N_5763,N_5667);
nor U6388 (N_6388,N_5903,N_5569);
and U6389 (N_6389,N_5886,N_5847);
xor U6390 (N_6390,N_5756,N_5837);
or U6391 (N_6391,N_5960,N_5891);
nor U6392 (N_6392,N_5554,N_5558);
or U6393 (N_6393,N_5917,N_5630);
nand U6394 (N_6394,N_5729,N_5885);
nor U6395 (N_6395,N_5893,N_5754);
nor U6396 (N_6396,N_5813,N_5724);
xor U6397 (N_6397,N_5635,N_5844);
and U6398 (N_6398,N_5827,N_5730);
and U6399 (N_6399,N_5721,N_5764);
nand U6400 (N_6400,N_5767,N_5820);
xnor U6401 (N_6401,N_5706,N_5716);
xor U6402 (N_6402,N_5964,N_5901);
xnor U6403 (N_6403,N_5623,N_5713);
nand U6404 (N_6404,N_5847,N_5873);
nor U6405 (N_6405,N_5998,N_5665);
nand U6406 (N_6406,N_5750,N_5948);
or U6407 (N_6407,N_5731,N_5696);
xor U6408 (N_6408,N_5681,N_5642);
or U6409 (N_6409,N_5729,N_5936);
xor U6410 (N_6410,N_5985,N_5636);
xnor U6411 (N_6411,N_5987,N_5804);
xor U6412 (N_6412,N_5842,N_5699);
xnor U6413 (N_6413,N_5751,N_5882);
and U6414 (N_6414,N_5775,N_5675);
and U6415 (N_6415,N_5925,N_5652);
or U6416 (N_6416,N_5974,N_5711);
xnor U6417 (N_6417,N_5619,N_5716);
or U6418 (N_6418,N_5904,N_5993);
nor U6419 (N_6419,N_5715,N_5863);
nand U6420 (N_6420,N_5732,N_5644);
nor U6421 (N_6421,N_5748,N_5958);
and U6422 (N_6422,N_5766,N_5669);
nor U6423 (N_6423,N_5840,N_5585);
and U6424 (N_6424,N_5689,N_5806);
nand U6425 (N_6425,N_5731,N_5958);
and U6426 (N_6426,N_5837,N_5555);
nor U6427 (N_6427,N_5639,N_5680);
and U6428 (N_6428,N_5758,N_5520);
or U6429 (N_6429,N_5731,N_5906);
nand U6430 (N_6430,N_5589,N_5528);
xnor U6431 (N_6431,N_5679,N_5976);
nand U6432 (N_6432,N_5535,N_5847);
and U6433 (N_6433,N_5769,N_5727);
and U6434 (N_6434,N_5532,N_5536);
or U6435 (N_6435,N_5734,N_5555);
nor U6436 (N_6436,N_5890,N_5951);
nor U6437 (N_6437,N_5810,N_5888);
nor U6438 (N_6438,N_5829,N_5567);
xor U6439 (N_6439,N_5842,N_5591);
nand U6440 (N_6440,N_5842,N_5764);
nor U6441 (N_6441,N_5769,N_5603);
and U6442 (N_6442,N_5516,N_5749);
and U6443 (N_6443,N_5994,N_5939);
nand U6444 (N_6444,N_5937,N_5740);
and U6445 (N_6445,N_5840,N_5556);
or U6446 (N_6446,N_5634,N_5728);
and U6447 (N_6447,N_5688,N_5991);
xnor U6448 (N_6448,N_5615,N_5653);
nand U6449 (N_6449,N_5813,N_5975);
and U6450 (N_6450,N_5725,N_5781);
and U6451 (N_6451,N_5692,N_5986);
or U6452 (N_6452,N_5577,N_5688);
or U6453 (N_6453,N_5508,N_5770);
or U6454 (N_6454,N_5918,N_5631);
and U6455 (N_6455,N_5522,N_5766);
xor U6456 (N_6456,N_5847,N_5641);
and U6457 (N_6457,N_5758,N_5925);
and U6458 (N_6458,N_5663,N_5761);
nand U6459 (N_6459,N_5917,N_5966);
xor U6460 (N_6460,N_5786,N_5773);
xor U6461 (N_6461,N_5827,N_5711);
and U6462 (N_6462,N_5786,N_5916);
and U6463 (N_6463,N_5893,N_5945);
and U6464 (N_6464,N_5645,N_5737);
xor U6465 (N_6465,N_5771,N_5809);
nand U6466 (N_6466,N_5656,N_5910);
and U6467 (N_6467,N_5954,N_5573);
xor U6468 (N_6468,N_5645,N_5839);
or U6469 (N_6469,N_5885,N_5518);
nand U6470 (N_6470,N_5626,N_5690);
xor U6471 (N_6471,N_5985,N_5818);
xor U6472 (N_6472,N_5772,N_5688);
xnor U6473 (N_6473,N_5677,N_5749);
xnor U6474 (N_6474,N_5524,N_5507);
nor U6475 (N_6475,N_5549,N_5562);
or U6476 (N_6476,N_5766,N_5919);
nand U6477 (N_6477,N_5628,N_5515);
xnor U6478 (N_6478,N_5546,N_5812);
nand U6479 (N_6479,N_5694,N_5875);
nor U6480 (N_6480,N_5812,N_5520);
or U6481 (N_6481,N_5699,N_5531);
and U6482 (N_6482,N_5654,N_5533);
nand U6483 (N_6483,N_5868,N_5561);
and U6484 (N_6484,N_5757,N_5897);
and U6485 (N_6485,N_5959,N_5872);
nand U6486 (N_6486,N_5792,N_5840);
nand U6487 (N_6487,N_5771,N_5653);
or U6488 (N_6488,N_5559,N_5760);
or U6489 (N_6489,N_5905,N_5674);
nand U6490 (N_6490,N_5592,N_5588);
nor U6491 (N_6491,N_5604,N_5625);
nand U6492 (N_6492,N_5766,N_5876);
and U6493 (N_6493,N_5656,N_5679);
xnor U6494 (N_6494,N_5589,N_5821);
or U6495 (N_6495,N_5851,N_5592);
and U6496 (N_6496,N_5559,N_5615);
or U6497 (N_6497,N_5792,N_5707);
and U6498 (N_6498,N_5810,N_5910);
and U6499 (N_6499,N_5835,N_5817);
xnor U6500 (N_6500,N_6326,N_6277);
xnor U6501 (N_6501,N_6306,N_6454);
xnor U6502 (N_6502,N_6276,N_6217);
xor U6503 (N_6503,N_6013,N_6052);
nand U6504 (N_6504,N_6265,N_6432);
nand U6505 (N_6505,N_6300,N_6411);
nand U6506 (N_6506,N_6246,N_6288);
and U6507 (N_6507,N_6285,N_6315);
xor U6508 (N_6508,N_6114,N_6191);
nand U6509 (N_6509,N_6385,N_6163);
nor U6510 (N_6510,N_6496,N_6290);
nand U6511 (N_6511,N_6005,N_6424);
xnor U6512 (N_6512,N_6193,N_6001);
nand U6513 (N_6513,N_6110,N_6268);
xnor U6514 (N_6514,N_6229,N_6425);
nor U6515 (N_6515,N_6490,N_6412);
xnor U6516 (N_6516,N_6477,N_6120);
xnor U6517 (N_6517,N_6206,N_6377);
nor U6518 (N_6518,N_6497,N_6108);
nor U6519 (N_6519,N_6488,N_6089);
xnor U6520 (N_6520,N_6062,N_6494);
xor U6521 (N_6521,N_6054,N_6117);
nand U6522 (N_6522,N_6298,N_6463);
xnor U6523 (N_6523,N_6393,N_6018);
nor U6524 (N_6524,N_6157,N_6338);
or U6525 (N_6525,N_6106,N_6003);
nand U6526 (N_6526,N_6261,N_6325);
xnor U6527 (N_6527,N_6014,N_6395);
nand U6528 (N_6528,N_6440,N_6188);
nor U6529 (N_6529,N_6213,N_6445);
and U6530 (N_6530,N_6242,N_6205);
and U6531 (N_6531,N_6384,N_6186);
nand U6532 (N_6532,N_6452,N_6070);
nand U6533 (N_6533,N_6389,N_6324);
and U6534 (N_6534,N_6124,N_6269);
and U6535 (N_6535,N_6155,N_6446);
xor U6536 (N_6536,N_6164,N_6207);
and U6537 (N_6537,N_6127,N_6467);
nor U6538 (N_6538,N_6015,N_6319);
nor U6539 (N_6539,N_6140,N_6274);
nand U6540 (N_6540,N_6299,N_6085);
or U6541 (N_6541,N_6112,N_6159);
and U6542 (N_6542,N_6403,N_6037);
nor U6543 (N_6543,N_6266,N_6255);
nand U6544 (N_6544,N_6078,N_6273);
xor U6545 (N_6545,N_6391,N_6336);
or U6546 (N_6546,N_6233,N_6133);
xnor U6547 (N_6547,N_6388,N_6184);
nand U6548 (N_6548,N_6378,N_6296);
xnor U6549 (N_6549,N_6495,N_6182);
and U6550 (N_6550,N_6209,N_6286);
xor U6551 (N_6551,N_6080,N_6252);
nand U6552 (N_6552,N_6101,N_6221);
nor U6553 (N_6553,N_6475,N_6485);
nand U6554 (N_6554,N_6308,N_6489);
or U6555 (N_6555,N_6121,N_6421);
nand U6556 (N_6556,N_6000,N_6459);
nand U6557 (N_6557,N_6358,N_6406);
or U6558 (N_6558,N_6382,N_6020);
and U6559 (N_6559,N_6270,N_6498);
or U6560 (N_6560,N_6444,N_6220);
and U6561 (N_6561,N_6478,N_6334);
xnor U6562 (N_6562,N_6098,N_6125);
nor U6563 (N_6563,N_6086,N_6049);
nor U6564 (N_6564,N_6064,N_6333);
nand U6565 (N_6565,N_6203,N_6038);
nand U6566 (N_6566,N_6431,N_6027);
nand U6567 (N_6567,N_6416,N_6046);
and U6568 (N_6568,N_6359,N_6142);
xor U6569 (N_6569,N_6017,N_6219);
or U6570 (N_6570,N_6257,N_6430);
nor U6571 (N_6571,N_6198,N_6415);
nand U6572 (N_6572,N_6011,N_6006);
nand U6573 (N_6573,N_6441,N_6063);
nor U6574 (N_6574,N_6151,N_6036);
xor U6575 (N_6575,N_6032,N_6429);
nand U6576 (N_6576,N_6464,N_6280);
xnor U6577 (N_6577,N_6414,N_6177);
nand U6578 (N_6578,N_6212,N_6022);
and U6579 (N_6579,N_6343,N_6116);
xor U6580 (N_6580,N_6012,N_6087);
and U6581 (N_6581,N_6442,N_6465);
nand U6582 (N_6582,N_6404,N_6060);
nor U6583 (N_6583,N_6312,N_6185);
and U6584 (N_6584,N_6313,N_6480);
and U6585 (N_6585,N_6433,N_6158);
nor U6586 (N_6586,N_6084,N_6316);
or U6587 (N_6587,N_6167,N_6335);
and U6588 (N_6588,N_6035,N_6437);
or U6589 (N_6589,N_6079,N_6225);
and U6590 (N_6590,N_6051,N_6428);
or U6591 (N_6591,N_6066,N_6448);
xnor U6592 (N_6592,N_6386,N_6251);
nor U6593 (N_6593,N_6435,N_6173);
or U6594 (N_6594,N_6392,N_6271);
and U6595 (N_6595,N_6281,N_6072);
nor U6596 (N_6596,N_6123,N_6234);
and U6597 (N_6597,N_6387,N_6249);
xor U6598 (N_6598,N_6195,N_6152);
xnor U6599 (N_6599,N_6239,N_6202);
nand U6600 (N_6600,N_6238,N_6287);
nand U6601 (N_6601,N_6449,N_6232);
nand U6602 (N_6602,N_6342,N_6109);
nor U6603 (N_6603,N_6081,N_6374);
nor U6604 (N_6604,N_6486,N_6199);
and U6605 (N_6605,N_6002,N_6367);
nor U6606 (N_6606,N_6210,N_6409);
xnor U6607 (N_6607,N_6473,N_6248);
and U6608 (N_6608,N_6043,N_6065);
nand U6609 (N_6609,N_6350,N_6471);
xnor U6610 (N_6610,N_6194,N_6344);
nor U6611 (N_6611,N_6126,N_6189);
nor U6612 (N_6612,N_6162,N_6351);
or U6613 (N_6613,N_6100,N_6460);
or U6614 (N_6614,N_6067,N_6154);
xnor U6615 (N_6615,N_6201,N_6456);
or U6616 (N_6616,N_6244,N_6147);
nand U6617 (N_6617,N_6399,N_6016);
or U6618 (N_6618,N_6137,N_6362);
nor U6619 (N_6619,N_6082,N_6420);
or U6620 (N_6620,N_6278,N_6128);
and U6621 (N_6621,N_6383,N_6056);
and U6622 (N_6622,N_6153,N_6057);
or U6623 (N_6623,N_6283,N_6474);
nor U6624 (N_6624,N_6092,N_6138);
nor U6625 (N_6625,N_6113,N_6090);
xnor U6626 (N_6626,N_6169,N_6224);
or U6627 (N_6627,N_6487,N_6472);
xor U6628 (N_6628,N_6439,N_6438);
or U6629 (N_6629,N_6462,N_6230);
nor U6630 (N_6630,N_6317,N_6118);
nand U6631 (N_6631,N_6307,N_6275);
nor U6632 (N_6632,N_6394,N_6007);
nand U6633 (N_6633,N_6115,N_6176);
or U6634 (N_6634,N_6434,N_6029);
nor U6635 (N_6635,N_6427,N_6131);
xor U6636 (N_6636,N_6226,N_6094);
nand U6637 (N_6637,N_6262,N_6492);
and U6638 (N_6638,N_6410,N_6339);
and U6639 (N_6639,N_6041,N_6245);
or U6640 (N_6640,N_6426,N_6341);
xnor U6641 (N_6641,N_6470,N_6160);
and U6642 (N_6642,N_6030,N_6039);
nor U6643 (N_6643,N_6004,N_6111);
or U6644 (N_6644,N_6197,N_6447);
nor U6645 (N_6645,N_6107,N_6103);
or U6646 (N_6646,N_6119,N_6216);
and U6647 (N_6647,N_6129,N_6150);
nand U6648 (N_6648,N_6413,N_6055);
or U6649 (N_6649,N_6284,N_6320);
nand U6650 (N_6650,N_6294,N_6321);
xor U6651 (N_6651,N_6301,N_6345);
nand U6652 (N_6652,N_6376,N_6491);
or U6653 (N_6653,N_6059,N_6024);
or U6654 (N_6654,N_6357,N_6305);
or U6655 (N_6655,N_6381,N_6293);
or U6656 (N_6656,N_6398,N_6122);
nor U6657 (N_6657,N_6348,N_6282);
nor U6658 (N_6658,N_6405,N_6483);
and U6659 (N_6659,N_6097,N_6025);
xnor U6660 (N_6660,N_6364,N_6061);
xor U6661 (N_6661,N_6396,N_6077);
xor U6662 (N_6662,N_6304,N_6401);
nor U6663 (N_6663,N_6372,N_6419);
nand U6664 (N_6664,N_6161,N_6019);
nand U6665 (N_6665,N_6250,N_6422);
and U6666 (N_6666,N_6149,N_6457);
xnor U6667 (N_6667,N_6310,N_6068);
nor U6668 (N_6668,N_6145,N_6190);
nor U6669 (N_6669,N_6314,N_6175);
xnor U6670 (N_6670,N_6400,N_6484);
nand U6671 (N_6671,N_6363,N_6267);
nor U6672 (N_6672,N_6228,N_6045);
nor U6673 (N_6673,N_6165,N_6170);
xnor U6674 (N_6674,N_6332,N_6379);
xor U6675 (N_6675,N_6214,N_6455);
nand U6676 (N_6676,N_6166,N_6071);
and U6677 (N_6677,N_6292,N_6258);
nor U6678 (N_6678,N_6337,N_6223);
and U6679 (N_6679,N_6243,N_6366);
or U6680 (N_6680,N_6026,N_6171);
xor U6681 (N_6681,N_6028,N_6371);
nor U6682 (N_6682,N_6204,N_6323);
and U6683 (N_6683,N_6443,N_6417);
xor U6684 (N_6684,N_6303,N_6256);
nor U6685 (N_6685,N_6134,N_6289);
xor U6686 (N_6686,N_6240,N_6347);
xnor U6687 (N_6687,N_6047,N_6048);
nand U6688 (N_6688,N_6178,N_6168);
or U6689 (N_6689,N_6453,N_6380);
xor U6690 (N_6690,N_6368,N_6156);
nand U6691 (N_6691,N_6192,N_6479);
or U6692 (N_6692,N_6075,N_6436);
and U6693 (N_6693,N_6076,N_6466);
or U6694 (N_6694,N_6095,N_6263);
nand U6695 (N_6695,N_6136,N_6318);
nand U6696 (N_6696,N_6143,N_6135);
xor U6697 (N_6697,N_6402,N_6236);
nand U6698 (N_6698,N_6196,N_6461);
nor U6699 (N_6699,N_6104,N_6218);
and U6700 (N_6700,N_6356,N_6481);
nor U6701 (N_6701,N_6264,N_6222);
nor U6702 (N_6702,N_6260,N_6349);
xnor U6703 (N_6703,N_6105,N_6352);
and U6704 (N_6704,N_6340,N_6328);
nand U6705 (N_6705,N_6099,N_6468);
xor U6706 (N_6706,N_6291,N_6361);
xor U6707 (N_6707,N_6272,N_6329);
nand U6708 (N_6708,N_6297,N_6181);
xnor U6709 (N_6709,N_6227,N_6040);
and U6710 (N_6710,N_6469,N_6088);
nor U6711 (N_6711,N_6309,N_6010);
xnor U6712 (N_6712,N_6390,N_6139);
or U6713 (N_6713,N_6295,N_6083);
and U6714 (N_6714,N_6208,N_6370);
and U6715 (N_6715,N_6353,N_6074);
or U6716 (N_6716,N_6021,N_6418);
nor U6717 (N_6717,N_6354,N_6130);
nand U6718 (N_6718,N_6458,N_6102);
nand U6719 (N_6719,N_6330,N_6322);
or U6720 (N_6720,N_6053,N_6327);
or U6721 (N_6721,N_6247,N_6397);
xnor U6722 (N_6722,N_6331,N_6034);
or U6723 (N_6723,N_6172,N_6174);
and U6724 (N_6724,N_6375,N_6423);
or U6725 (N_6725,N_6096,N_6365);
or U6726 (N_6726,N_6008,N_6451);
nor U6727 (N_6727,N_6259,N_6499);
nor U6728 (N_6728,N_6346,N_6302);
xnor U6729 (N_6729,N_6144,N_6355);
nand U6730 (N_6730,N_6211,N_6369);
nor U6731 (N_6731,N_6215,N_6482);
xnor U6732 (N_6732,N_6093,N_6254);
xor U6733 (N_6733,N_6373,N_6141);
and U6734 (N_6734,N_6031,N_6058);
and U6735 (N_6735,N_6042,N_6279);
xor U6736 (N_6736,N_6360,N_6146);
or U6737 (N_6737,N_6450,N_6073);
nor U6738 (N_6738,N_6023,N_6033);
and U6739 (N_6739,N_6235,N_6009);
and U6740 (N_6740,N_6069,N_6241);
nor U6741 (N_6741,N_6407,N_6200);
or U6742 (N_6742,N_6408,N_6179);
and U6743 (N_6743,N_6183,N_6091);
nor U6744 (N_6744,N_6044,N_6253);
and U6745 (N_6745,N_6132,N_6187);
nor U6746 (N_6746,N_6180,N_6231);
xnor U6747 (N_6747,N_6148,N_6311);
nor U6748 (N_6748,N_6050,N_6493);
nor U6749 (N_6749,N_6476,N_6237);
nor U6750 (N_6750,N_6301,N_6010);
and U6751 (N_6751,N_6131,N_6063);
or U6752 (N_6752,N_6235,N_6495);
xor U6753 (N_6753,N_6233,N_6341);
or U6754 (N_6754,N_6266,N_6256);
nor U6755 (N_6755,N_6013,N_6232);
nand U6756 (N_6756,N_6390,N_6101);
nand U6757 (N_6757,N_6248,N_6158);
nand U6758 (N_6758,N_6336,N_6394);
xnor U6759 (N_6759,N_6103,N_6260);
nor U6760 (N_6760,N_6383,N_6074);
and U6761 (N_6761,N_6143,N_6286);
xnor U6762 (N_6762,N_6053,N_6115);
nor U6763 (N_6763,N_6038,N_6177);
or U6764 (N_6764,N_6249,N_6383);
and U6765 (N_6765,N_6354,N_6365);
nor U6766 (N_6766,N_6368,N_6400);
nor U6767 (N_6767,N_6165,N_6121);
or U6768 (N_6768,N_6429,N_6417);
and U6769 (N_6769,N_6282,N_6437);
nor U6770 (N_6770,N_6277,N_6191);
nor U6771 (N_6771,N_6254,N_6213);
or U6772 (N_6772,N_6308,N_6301);
xor U6773 (N_6773,N_6450,N_6326);
nor U6774 (N_6774,N_6451,N_6166);
or U6775 (N_6775,N_6140,N_6441);
nor U6776 (N_6776,N_6492,N_6491);
nand U6777 (N_6777,N_6481,N_6379);
or U6778 (N_6778,N_6259,N_6374);
xnor U6779 (N_6779,N_6470,N_6372);
xor U6780 (N_6780,N_6271,N_6266);
nand U6781 (N_6781,N_6161,N_6170);
nand U6782 (N_6782,N_6367,N_6432);
xor U6783 (N_6783,N_6122,N_6136);
and U6784 (N_6784,N_6384,N_6069);
or U6785 (N_6785,N_6283,N_6161);
nand U6786 (N_6786,N_6096,N_6132);
nor U6787 (N_6787,N_6453,N_6213);
or U6788 (N_6788,N_6465,N_6141);
nor U6789 (N_6789,N_6139,N_6017);
and U6790 (N_6790,N_6068,N_6473);
or U6791 (N_6791,N_6258,N_6052);
or U6792 (N_6792,N_6025,N_6283);
or U6793 (N_6793,N_6150,N_6313);
nand U6794 (N_6794,N_6101,N_6250);
xnor U6795 (N_6795,N_6304,N_6356);
nand U6796 (N_6796,N_6078,N_6278);
nand U6797 (N_6797,N_6171,N_6468);
nor U6798 (N_6798,N_6355,N_6397);
nand U6799 (N_6799,N_6097,N_6026);
and U6800 (N_6800,N_6038,N_6438);
nand U6801 (N_6801,N_6037,N_6006);
and U6802 (N_6802,N_6114,N_6100);
nor U6803 (N_6803,N_6436,N_6057);
nand U6804 (N_6804,N_6297,N_6316);
xor U6805 (N_6805,N_6144,N_6213);
and U6806 (N_6806,N_6109,N_6159);
and U6807 (N_6807,N_6072,N_6140);
xnor U6808 (N_6808,N_6303,N_6127);
xor U6809 (N_6809,N_6057,N_6396);
and U6810 (N_6810,N_6481,N_6183);
and U6811 (N_6811,N_6027,N_6453);
nor U6812 (N_6812,N_6293,N_6052);
nor U6813 (N_6813,N_6255,N_6392);
or U6814 (N_6814,N_6486,N_6454);
nor U6815 (N_6815,N_6048,N_6009);
nand U6816 (N_6816,N_6086,N_6486);
or U6817 (N_6817,N_6494,N_6100);
nand U6818 (N_6818,N_6371,N_6052);
nor U6819 (N_6819,N_6153,N_6006);
and U6820 (N_6820,N_6180,N_6370);
xnor U6821 (N_6821,N_6162,N_6286);
nor U6822 (N_6822,N_6305,N_6104);
and U6823 (N_6823,N_6031,N_6471);
or U6824 (N_6824,N_6037,N_6298);
and U6825 (N_6825,N_6262,N_6004);
nand U6826 (N_6826,N_6267,N_6270);
nand U6827 (N_6827,N_6451,N_6172);
nand U6828 (N_6828,N_6065,N_6175);
xnor U6829 (N_6829,N_6197,N_6477);
and U6830 (N_6830,N_6091,N_6162);
nor U6831 (N_6831,N_6262,N_6285);
or U6832 (N_6832,N_6020,N_6461);
xnor U6833 (N_6833,N_6163,N_6239);
xor U6834 (N_6834,N_6280,N_6013);
nor U6835 (N_6835,N_6454,N_6080);
and U6836 (N_6836,N_6434,N_6389);
nand U6837 (N_6837,N_6330,N_6278);
or U6838 (N_6838,N_6007,N_6179);
nand U6839 (N_6839,N_6355,N_6466);
and U6840 (N_6840,N_6389,N_6478);
xor U6841 (N_6841,N_6157,N_6203);
nand U6842 (N_6842,N_6070,N_6145);
and U6843 (N_6843,N_6156,N_6086);
nand U6844 (N_6844,N_6077,N_6375);
or U6845 (N_6845,N_6285,N_6191);
or U6846 (N_6846,N_6266,N_6394);
xor U6847 (N_6847,N_6238,N_6367);
nand U6848 (N_6848,N_6383,N_6467);
nor U6849 (N_6849,N_6339,N_6140);
or U6850 (N_6850,N_6238,N_6475);
or U6851 (N_6851,N_6131,N_6444);
xor U6852 (N_6852,N_6240,N_6104);
xor U6853 (N_6853,N_6338,N_6173);
nand U6854 (N_6854,N_6416,N_6041);
and U6855 (N_6855,N_6293,N_6244);
xor U6856 (N_6856,N_6408,N_6050);
xor U6857 (N_6857,N_6054,N_6490);
and U6858 (N_6858,N_6129,N_6191);
nand U6859 (N_6859,N_6005,N_6131);
or U6860 (N_6860,N_6146,N_6353);
xnor U6861 (N_6861,N_6474,N_6046);
and U6862 (N_6862,N_6005,N_6148);
or U6863 (N_6863,N_6084,N_6431);
xor U6864 (N_6864,N_6193,N_6332);
xnor U6865 (N_6865,N_6119,N_6112);
xnor U6866 (N_6866,N_6376,N_6359);
nor U6867 (N_6867,N_6294,N_6160);
xor U6868 (N_6868,N_6147,N_6199);
xor U6869 (N_6869,N_6381,N_6291);
and U6870 (N_6870,N_6023,N_6079);
nand U6871 (N_6871,N_6496,N_6371);
nor U6872 (N_6872,N_6332,N_6306);
nor U6873 (N_6873,N_6047,N_6435);
and U6874 (N_6874,N_6039,N_6397);
nand U6875 (N_6875,N_6004,N_6353);
and U6876 (N_6876,N_6185,N_6091);
xnor U6877 (N_6877,N_6213,N_6330);
xnor U6878 (N_6878,N_6015,N_6244);
and U6879 (N_6879,N_6135,N_6132);
nand U6880 (N_6880,N_6358,N_6112);
nand U6881 (N_6881,N_6476,N_6144);
nand U6882 (N_6882,N_6045,N_6004);
or U6883 (N_6883,N_6287,N_6031);
nor U6884 (N_6884,N_6299,N_6338);
or U6885 (N_6885,N_6320,N_6184);
nand U6886 (N_6886,N_6461,N_6203);
nor U6887 (N_6887,N_6038,N_6259);
or U6888 (N_6888,N_6264,N_6401);
and U6889 (N_6889,N_6429,N_6000);
nand U6890 (N_6890,N_6186,N_6038);
xnor U6891 (N_6891,N_6342,N_6391);
and U6892 (N_6892,N_6337,N_6408);
or U6893 (N_6893,N_6075,N_6284);
or U6894 (N_6894,N_6101,N_6409);
nor U6895 (N_6895,N_6180,N_6045);
and U6896 (N_6896,N_6020,N_6414);
nor U6897 (N_6897,N_6077,N_6480);
or U6898 (N_6898,N_6358,N_6430);
nand U6899 (N_6899,N_6170,N_6369);
xnor U6900 (N_6900,N_6009,N_6187);
or U6901 (N_6901,N_6246,N_6385);
xnor U6902 (N_6902,N_6412,N_6223);
and U6903 (N_6903,N_6200,N_6060);
nor U6904 (N_6904,N_6220,N_6459);
nor U6905 (N_6905,N_6079,N_6107);
xor U6906 (N_6906,N_6133,N_6112);
and U6907 (N_6907,N_6294,N_6045);
xor U6908 (N_6908,N_6367,N_6124);
nor U6909 (N_6909,N_6322,N_6000);
nand U6910 (N_6910,N_6119,N_6138);
or U6911 (N_6911,N_6168,N_6240);
or U6912 (N_6912,N_6097,N_6260);
nand U6913 (N_6913,N_6287,N_6395);
xor U6914 (N_6914,N_6435,N_6198);
and U6915 (N_6915,N_6169,N_6387);
nor U6916 (N_6916,N_6203,N_6037);
nand U6917 (N_6917,N_6071,N_6239);
or U6918 (N_6918,N_6450,N_6453);
or U6919 (N_6919,N_6374,N_6092);
nand U6920 (N_6920,N_6318,N_6480);
nand U6921 (N_6921,N_6014,N_6266);
nor U6922 (N_6922,N_6323,N_6374);
nor U6923 (N_6923,N_6478,N_6155);
xor U6924 (N_6924,N_6196,N_6314);
xor U6925 (N_6925,N_6154,N_6204);
or U6926 (N_6926,N_6439,N_6348);
nor U6927 (N_6927,N_6070,N_6076);
and U6928 (N_6928,N_6282,N_6084);
nor U6929 (N_6929,N_6402,N_6183);
or U6930 (N_6930,N_6401,N_6337);
xor U6931 (N_6931,N_6068,N_6184);
nand U6932 (N_6932,N_6275,N_6034);
and U6933 (N_6933,N_6052,N_6132);
and U6934 (N_6934,N_6310,N_6019);
or U6935 (N_6935,N_6360,N_6155);
and U6936 (N_6936,N_6446,N_6023);
and U6937 (N_6937,N_6279,N_6498);
nor U6938 (N_6938,N_6440,N_6187);
nor U6939 (N_6939,N_6331,N_6495);
and U6940 (N_6940,N_6330,N_6457);
or U6941 (N_6941,N_6367,N_6185);
nand U6942 (N_6942,N_6103,N_6423);
or U6943 (N_6943,N_6143,N_6463);
or U6944 (N_6944,N_6291,N_6499);
xor U6945 (N_6945,N_6411,N_6287);
xnor U6946 (N_6946,N_6461,N_6057);
nand U6947 (N_6947,N_6265,N_6126);
nand U6948 (N_6948,N_6479,N_6205);
or U6949 (N_6949,N_6167,N_6365);
nor U6950 (N_6950,N_6395,N_6321);
or U6951 (N_6951,N_6170,N_6047);
nor U6952 (N_6952,N_6465,N_6353);
and U6953 (N_6953,N_6065,N_6145);
xnor U6954 (N_6954,N_6121,N_6403);
nand U6955 (N_6955,N_6351,N_6170);
or U6956 (N_6956,N_6163,N_6104);
xor U6957 (N_6957,N_6250,N_6399);
xnor U6958 (N_6958,N_6098,N_6057);
nand U6959 (N_6959,N_6168,N_6224);
nand U6960 (N_6960,N_6324,N_6401);
nand U6961 (N_6961,N_6006,N_6104);
nor U6962 (N_6962,N_6066,N_6421);
xor U6963 (N_6963,N_6392,N_6017);
xor U6964 (N_6964,N_6001,N_6456);
and U6965 (N_6965,N_6221,N_6325);
nand U6966 (N_6966,N_6011,N_6060);
nand U6967 (N_6967,N_6291,N_6108);
or U6968 (N_6968,N_6274,N_6380);
nand U6969 (N_6969,N_6479,N_6255);
and U6970 (N_6970,N_6487,N_6074);
nand U6971 (N_6971,N_6456,N_6211);
nand U6972 (N_6972,N_6179,N_6152);
nand U6973 (N_6973,N_6042,N_6478);
and U6974 (N_6974,N_6485,N_6368);
xor U6975 (N_6975,N_6165,N_6109);
xnor U6976 (N_6976,N_6392,N_6432);
nand U6977 (N_6977,N_6096,N_6094);
and U6978 (N_6978,N_6380,N_6003);
and U6979 (N_6979,N_6197,N_6362);
or U6980 (N_6980,N_6300,N_6358);
and U6981 (N_6981,N_6357,N_6255);
and U6982 (N_6982,N_6270,N_6210);
xnor U6983 (N_6983,N_6289,N_6252);
and U6984 (N_6984,N_6335,N_6388);
nor U6985 (N_6985,N_6372,N_6390);
xor U6986 (N_6986,N_6209,N_6385);
xor U6987 (N_6987,N_6458,N_6353);
xor U6988 (N_6988,N_6086,N_6363);
or U6989 (N_6989,N_6385,N_6328);
nand U6990 (N_6990,N_6028,N_6360);
xnor U6991 (N_6991,N_6293,N_6472);
and U6992 (N_6992,N_6473,N_6275);
or U6993 (N_6993,N_6257,N_6024);
nand U6994 (N_6994,N_6158,N_6173);
nor U6995 (N_6995,N_6250,N_6432);
or U6996 (N_6996,N_6361,N_6248);
nor U6997 (N_6997,N_6392,N_6377);
nor U6998 (N_6998,N_6100,N_6351);
and U6999 (N_6999,N_6086,N_6361);
or U7000 (N_7000,N_6532,N_6700);
nand U7001 (N_7001,N_6855,N_6626);
and U7002 (N_7002,N_6678,N_6932);
nor U7003 (N_7003,N_6738,N_6995);
nand U7004 (N_7004,N_6925,N_6865);
xnor U7005 (N_7005,N_6592,N_6597);
nor U7006 (N_7006,N_6546,N_6934);
nand U7007 (N_7007,N_6685,N_6548);
and U7008 (N_7008,N_6924,N_6543);
and U7009 (N_7009,N_6745,N_6535);
nor U7010 (N_7010,N_6968,N_6945);
nor U7011 (N_7011,N_6591,N_6607);
xnor U7012 (N_7012,N_6692,N_6832);
and U7013 (N_7013,N_6820,N_6755);
nor U7014 (N_7014,N_6710,N_6796);
nor U7015 (N_7015,N_6754,N_6926);
or U7016 (N_7016,N_6653,N_6578);
nor U7017 (N_7017,N_6879,N_6654);
nor U7018 (N_7018,N_6861,N_6839);
xor U7019 (N_7019,N_6523,N_6978);
or U7020 (N_7020,N_6937,N_6791);
and U7021 (N_7021,N_6731,N_6531);
nor U7022 (N_7022,N_6665,N_6849);
or U7023 (N_7023,N_6793,N_6562);
and U7024 (N_7024,N_6711,N_6641);
or U7025 (N_7025,N_6911,N_6743);
and U7026 (N_7026,N_6867,N_6646);
nor U7027 (N_7027,N_6724,N_6957);
or U7028 (N_7028,N_6918,N_6903);
or U7029 (N_7029,N_6545,N_6746);
and U7030 (N_7030,N_6555,N_6589);
nor U7031 (N_7031,N_6949,N_6519);
nand U7032 (N_7032,N_6517,N_6502);
and U7033 (N_7033,N_6857,N_6844);
and U7034 (N_7034,N_6884,N_6987);
nand U7035 (N_7035,N_6506,N_6912);
xnor U7036 (N_7036,N_6979,N_6583);
xnor U7037 (N_7037,N_6803,N_6668);
nor U7038 (N_7038,N_6969,N_6584);
nand U7039 (N_7039,N_6602,N_6947);
or U7040 (N_7040,N_6614,N_6670);
or U7041 (N_7041,N_6950,N_6890);
or U7042 (N_7042,N_6909,N_6778);
or U7043 (N_7043,N_6656,N_6784);
nand U7044 (N_7044,N_6822,N_6615);
or U7045 (N_7045,N_6958,N_6818);
or U7046 (N_7046,N_6919,N_6913);
and U7047 (N_7047,N_6579,N_6892);
xnor U7048 (N_7048,N_6734,N_6612);
or U7049 (N_7049,N_6792,N_6732);
and U7050 (N_7050,N_6671,N_6853);
xor U7051 (N_7051,N_6994,N_6600);
nor U7052 (N_7052,N_6898,N_6908);
nor U7053 (N_7053,N_6975,N_6508);
nand U7054 (N_7054,N_6885,N_6974);
xnor U7055 (N_7055,N_6776,N_6888);
or U7056 (N_7056,N_6990,N_6611);
nor U7057 (N_7057,N_6681,N_6633);
or U7058 (N_7058,N_6833,N_6554);
nand U7059 (N_7059,N_6730,N_6511);
and U7060 (N_7060,N_6787,N_6774);
nand U7061 (N_7061,N_6953,N_6902);
xnor U7062 (N_7062,N_6630,N_6663);
or U7063 (N_7063,N_6538,N_6624);
nand U7064 (N_7064,N_6827,N_6807);
nor U7065 (N_7065,N_6765,N_6799);
and U7066 (N_7066,N_6625,N_6946);
nor U7067 (N_7067,N_6920,N_6571);
or U7068 (N_7068,N_6749,N_6878);
nor U7069 (N_7069,N_6870,N_6860);
nor U7070 (N_7070,N_6530,N_6631);
or U7071 (N_7071,N_6553,N_6580);
or U7072 (N_7072,N_6736,N_6815);
nor U7073 (N_7073,N_6739,N_6882);
nor U7074 (N_7074,N_6526,N_6836);
and U7075 (N_7075,N_6610,N_6603);
nor U7076 (N_7076,N_6564,N_6690);
xor U7077 (N_7077,N_6775,N_6856);
or U7078 (N_7078,N_6988,N_6748);
or U7079 (N_7079,N_6706,N_6843);
or U7080 (N_7080,N_6936,N_6770);
and U7081 (N_7081,N_6921,N_6956);
xnor U7082 (N_7082,N_6542,N_6834);
xnor U7083 (N_7083,N_6507,N_6735);
or U7084 (N_7084,N_6842,N_6698);
or U7085 (N_7085,N_6740,N_6773);
xnor U7086 (N_7086,N_6989,N_6725);
nand U7087 (N_7087,N_6874,N_6664);
xnor U7088 (N_7088,N_6951,N_6719);
xor U7089 (N_7089,N_6621,N_6915);
or U7090 (N_7090,N_6565,N_6804);
nand U7091 (N_7091,N_6782,N_6869);
and U7092 (N_7092,N_6723,N_6797);
nor U7093 (N_7093,N_6941,N_6572);
xor U7094 (N_7094,N_6753,N_6635);
or U7095 (N_7095,N_6588,N_6914);
or U7096 (N_7096,N_6986,N_6751);
nor U7097 (N_7097,N_6872,N_6858);
or U7098 (N_7098,N_6595,N_6650);
xnor U7099 (N_7099,N_6707,N_6848);
xnor U7100 (N_7100,N_6805,N_6733);
nand U7101 (N_7101,N_6613,N_6960);
xor U7102 (N_7102,N_6559,N_6647);
nor U7103 (N_7103,N_6574,N_6606);
or U7104 (N_7104,N_6862,N_6504);
or U7105 (N_7105,N_6819,N_6666);
nor U7106 (N_7106,N_6906,N_6540);
nand U7107 (N_7107,N_6917,N_6800);
xor U7108 (N_7108,N_6769,N_6944);
xnor U7109 (N_7109,N_6510,N_6720);
and U7110 (N_7110,N_6761,N_6756);
xnor U7111 (N_7111,N_6752,N_6729);
xnor U7112 (N_7112,N_6712,N_6891);
or U7113 (N_7113,N_6826,N_6599);
nor U7114 (N_7114,N_6705,N_6965);
xnor U7115 (N_7115,N_6806,N_6901);
xnor U7116 (N_7116,N_6929,N_6655);
or U7117 (N_7117,N_6967,N_6868);
and U7118 (N_7118,N_6628,N_6515);
and U7119 (N_7119,N_6840,N_6964);
nand U7120 (N_7120,N_6557,N_6977);
nand U7121 (N_7121,N_6766,N_6943);
or U7122 (N_7122,N_6899,N_6777);
xor U7123 (N_7123,N_6623,N_6718);
and U7124 (N_7124,N_6781,N_6881);
nor U7125 (N_7125,N_6616,N_6636);
xor U7126 (N_7126,N_6648,N_6505);
and U7127 (N_7127,N_6566,N_6586);
nand U7128 (N_7128,N_6859,N_6852);
and U7129 (N_7129,N_6737,N_6846);
xnor U7130 (N_7130,N_6795,N_6701);
or U7131 (N_7131,N_6930,N_6823);
and U7132 (N_7132,N_6722,N_6577);
and U7133 (N_7133,N_6651,N_6696);
or U7134 (N_7134,N_6959,N_6939);
and U7135 (N_7135,N_6644,N_6598);
nor U7136 (N_7136,N_6889,N_6713);
xor U7137 (N_7137,N_6760,N_6617);
xnor U7138 (N_7138,N_6813,N_6672);
and U7139 (N_7139,N_6829,N_6618);
or U7140 (N_7140,N_6927,N_6871);
and U7141 (N_7141,N_6998,N_6916);
nor U7142 (N_7142,N_6667,N_6601);
nand U7143 (N_7143,N_6933,N_6841);
or U7144 (N_7144,N_6809,N_6680);
nor U7145 (N_7145,N_6802,N_6981);
nand U7146 (N_7146,N_6972,N_6593);
xnor U7147 (N_7147,N_6980,N_6768);
nand U7148 (N_7148,N_6721,N_6716);
or U7149 (N_7149,N_6767,N_6652);
xor U7150 (N_7150,N_6609,N_6691);
nand U7151 (N_7151,N_6684,N_6544);
nor U7152 (N_7152,N_6786,N_6703);
xor U7153 (N_7153,N_6556,N_6997);
and U7154 (N_7154,N_6500,N_6824);
nand U7155 (N_7155,N_6552,N_6771);
xor U7156 (N_7156,N_6715,N_6895);
or U7157 (N_7157,N_6970,N_6558);
xnor U7158 (N_7158,N_6886,N_6582);
and U7159 (N_7159,N_6780,N_6568);
nor U7160 (N_7160,N_6640,N_6744);
nand U7161 (N_7161,N_6509,N_6539);
nand U7162 (N_7162,N_6596,N_6900);
xnor U7163 (N_7163,N_6928,N_6785);
nor U7164 (N_7164,N_6940,N_6534);
or U7165 (N_7165,N_6764,N_6687);
nand U7166 (N_7166,N_6637,N_6717);
nor U7167 (N_7167,N_6605,N_6828);
xnor U7168 (N_7168,N_6904,N_6570);
nand U7169 (N_7169,N_6541,N_6661);
nor U7170 (N_7170,N_6576,N_6962);
or U7171 (N_7171,N_6693,N_6503);
nor U7172 (N_7172,N_6838,N_6873);
nand U7173 (N_7173,N_6708,N_6963);
nand U7174 (N_7174,N_6847,N_6938);
nand U7175 (N_7175,N_6875,N_6854);
or U7176 (N_7176,N_6573,N_6851);
and U7177 (N_7177,N_6877,N_6643);
or U7178 (N_7178,N_6547,N_6677);
xnor U7179 (N_7179,N_6525,N_6537);
nor U7180 (N_7180,N_6520,N_6669);
nor U7181 (N_7181,N_6984,N_6931);
xnor U7182 (N_7182,N_6627,N_6830);
xor U7183 (N_7183,N_6608,N_6971);
and U7184 (N_7184,N_6682,N_6704);
xnor U7185 (N_7185,N_6763,N_6801);
xnor U7186 (N_7186,N_6935,N_6560);
xor U7187 (N_7187,N_6662,N_6821);
or U7188 (N_7188,N_6955,N_6694);
and U7189 (N_7189,N_6728,N_6587);
or U7190 (N_7190,N_6894,N_6522);
nand U7191 (N_7191,N_6845,N_6695);
and U7192 (N_7192,N_6619,N_6996);
or U7193 (N_7193,N_6702,N_6622);
and U7194 (N_7194,N_6810,N_6549);
and U7195 (N_7195,N_6590,N_6741);
and U7196 (N_7196,N_6714,N_6524);
or U7197 (N_7197,N_6659,N_6660);
nand U7198 (N_7198,N_6893,N_6699);
xnor U7199 (N_7199,N_6529,N_6658);
nand U7200 (N_7200,N_6910,N_6762);
or U7201 (N_7201,N_6518,N_6569);
or U7202 (N_7202,N_6814,N_6866);
or U7203 (N_7203,N_6789,N_6788);
nand U7204 (N_7204,N_6533,N_6727);
nor U7205 (N_7205,N_6897,N_6521);
or U7206 (N_7206,N_6649,N_6516);
and U7207 (N_7207,N_6992,N_6620);
xnor U7208 (N_7208,N_6999,N_6863);
nor U7209 (N_7209,N_6657,N_6513);
and U7210 (N_7210,N_6629,N_6790);
nor U7211 (N_7211,N_6816,N_6837);
nor U7212 (N_7212,N_6501,N_6575);
and U7213 (N_7213,N_6581,N_6674);
nor U7214 (N_7214,N_6683,N_6676);
and U7215 (N_7215,N_6905,N_6634);
xor U7216 (N_7216,N_6952,N_6907);
or U7217 (N_7217,N_6942,N_6779);
or U7218 (N_7218,N_6679,N_6645);
xor U7219 (N_7219,N_6585,N_6750);
and U7220 (N_7220,N_6675,N_6864);
nor U7221 (N_7221,N_6551,N_6689);
or U7222 (N_7222,N_6604,N_6567);
nor U7223 (N_7223,N_6880,N_6561);
xnor U7224 (N_7224,N_6563,N_6726);
and U7225 (N_7225,N_6817,N_6673);
or U7226 (N_7226,N_6747,N_6923);
nor U7227 (N_7227,N_6811,N_6876);
nor U7228 (N_7228,N_6514,N_6594);
and U7229 (N_7229,N_6983,N_6512);
or U7230 (N_7230,N_6922,N_6825);
nor U7231 (N_7231,N_6697,N_6757);
or U7232 (N_7232,N_6993,N_6632);
or U7233 (N_7233,N_6973,N_6686);
or U7234 (N_7234,N_6976,N_6896);
or U7235 (N_7235,N_6985,N_6688);
and U7236 (N_7236,N_6982,N_6642);
xnor U7237 (N_7237,N_6794,N_6948);
nand U7238 (N_7238,N_6961,N_6783);
and U7239 (N_7239,N_6835,N_6954);
or U7240 (N_7240,N_6991,N_6639);
nor U7241 (N_7241,N_6772,N_6759);
xnor U7242 (N_7242,N_6798,N_6887);
and U7243 (N_7243,N_6528,N_6812);
nand U7244 (N_7244,N_6638,N_6536);
and U7245 (N_7245,N_6709,N_6550);
xor U7246 (N_7246,N_6966,N_6850);
nand U7247 (N_7247,N_6808,N_6831);
or U7248 (N_7248,N_6883,N_6742);
or U7249 (N_7249,N_6527,N_6758);
and U7250 (N_7250,N_6951,N_6849);
nand U7251 (N_7251,N_6893,N_6852);
and U7252 (N_7252,N_6761,N_6904);
xor U7253 (N_7253,N_6552,N_6629);
nand U7254 (N_7254,N_6689,N_6834);
xor U7255 (N_7255,N_6885,N_6835);
and U7256 (N_7256,N_6874,N_6944);
nor U7257 (N_7257,N_6963,N_6864);
nor U7258 (N_7258,N_6962,N_6620);
or U7259 (N_7259,N_6509,N_6642);
xnor U7260 (N_7260,N_6827,N_6541);
and U7261 (N_7261,N_6963,N_6733);
xnor U7262 (N_7262,N_6992,N_6740);
nand U7263 (N_7263,N_6801,N_6915);
nand U7264 (N_7264,N_6749,N_6818);
or U7265 (N_7265,N_6712,N_6642);
nor U7266 (N_7266,N_6574,N_6716);
nor U7267 (N_7267,N_6774,N_6650);
xnor U7268 (N_7268,N_6850,N_6706);
or U7269 (N_7269,N_6781,N_6733);
xnor U7270 (N_7270,N_6606,N_6627);
xnor U7271 (N_7271,N_6748,N_6695);
xnor U7272 (N_7272,N_6686,N_6914);
or U7273 (N_7273,N_6708,N_6722);
and U7274 (N_7274,N_6653,N_6510);
nand U7275 (N_7275,N_6518,N_6549);
xor U7276 (N_7276,N_6851,N_6987);
and U7277 (N_7277,N_6796,N_6537);
and U7278 (N_7278,N_6531,N_6527);
xor U7279 (N_7279,N_6603,N_6664);
xor U7280 (N_7280,N_6875,N_6728);
and U7281 (N_7281,N_6539,N_6510);
and U7282 (N_7282,N_6531,N_6720);
nor U7283 (N_7283,N_6606,N_6974);
or U7284 (N_7284,N_6966,N_6986);
xnor U7285 (N_7285,N_6831,N_6833);
or U7286 (N_7286,N_6707,N_6815);
xnor U7287 (N_7287,N_6890,N_6561);
nand U7288 (N_7288,N_6910,N_6850);
and U7289 (N_7289,N_6963,N_6921);
xnor U7290 (N_7290,N_6670,N_6851);
nand U7291 (N_7291,N_6624,N_6768);
and U7292 (N_7292,N_6740,N_6968);
xor U7293 (N_7293,N_6738,N_6683);
or U7294 (N_7294,N_6659,N_6865);
nor U7295 (N_7295,N_6858,N_6931);
nand U7296 (N_7296,N_6758,N_6644);
or U7297 (N_7297,N_6561,N_6792);
xor U7298 (N_7298,N_6696,N_6775);
xnor U7299 (N_7299,N_6690,N_6784);
nor U7300 (N_7300,N_6641,N_6784);
and U7301 (N_7301,N_6858,N_6545);
xnor U7302 (N_7302,N_6912,N_6969);
xnor U7303 (N_7303,N_6833,N_6564);
and U7304 (N_7304,N_6893,N_6980);
xnor U7305 (N_7305,N_6964,N_6744);
and U7306 (N_7306,N_6529,N_6606);
or U7307 (N_7307,N_6642,N_6656);
xnor U7308 (N_7308,N_6520,N_6628);
nand U7309 (N_7309,N_6636,N_6576);
or U7310 (N_7310,N_6608,N_6535);
or U7311 (N_7311,N_6617,N_6535);
nor U7312 (N_7312,N_6838,N_6980);
nor U7313 (N_7313,N_6938,N_6849);
xor U7314 (N_7314,N_6921,N_6873);
nand U7315 (N_7315,N_6784,N_6557);
xor U7316 (N_7316,N_6604,N_6963);
or U7317 (N_7317,N_6756,N_6654);
and U7318 (N_7318,N_6916,N_6737);
or U7319 (N_7319,N_6547,N_6752);
xnor U7320 (N_7320,N_6853,N_6979);
xor U7321 (N_7321,N_6964,N_6778);
nand U7322 (N_7322,N_6593,N_6541);
and U7323 (N_7323,N_6509,N_6827);
nor U7324 (N_7324,N_6831,N_6571);
nand U7325 (N_7325,N_6708,N_6690);
nor U7326 (N_7326,N_6711,N_6672);
xor U7327 (N_7327,N_6591,N_6942);
or U7328 (N_7328,N_6935,N_6746);
or U7329 (N_7329,N_6507,N_6809);
nor U7330 (N_7330,N_6529,N_6705);
nand U7331 (N_7331,N_6901,N_6848);
and U7332 (N_7332,N_6532,N_6863);
and U7333 (N_7333,N_6868,N_6971);
xor U7334 (N_7334,N_6821,N_6672);
xor U7335 (N_7335,N_6687,N_6729);
and U7336 (N_7336,N_6788,N_6861);
or U7337 (N_7337,N_6822,N_6957);
or U7338 (N_7338,N_6538,N_6932);
xor U7339 (N_7339,N_6768,N_6829);
nor U7340 (N_7340,N_6714,N_6884);
or U7341 (N_7341,N_6718,N_6929);
or U7342 (N_7342,N_6524,N_6691);
xnor U7343 (N_7343,N_6833,N_6980);
nand U7344 (N_7344,N_6874,N_6668);
or U7345 (N_7345,N_6758,N_6714);
and U7346 (N_7346,N_6763,N_6972);
xnor U7347 (N_7347,N_6984,N_6769);
nor U7348 (N_7348,N_6641,N_6701);
or U7349 (N_7349,N_6646,N_6846);
xnor U7350 (N_7350,N_6836,N_6948);
and U7351 (N_7351,N_6918,N_6553);
xor U7352 (N_7352,N_6752,N_6727);
xor U7353 (N_7353,N_6567,N_6772);
nor U7354 (N_7354,N_6514,N_6748);
and U7355 (N_7355,N_6989,N_6902);
nor U7356 (N_7356,N_6680,N_6705);
xnor U7357 (N_7357,N_6692,N_6860);
nand U7358 (N_7358,N_6607,N_6539);
nand U7359 (N_7359,N_6623,N_6617);
xnor U7360 (N_7360,N_6755,N_6771);
xnor U7361 (N_7361,N_6717,N_6831);
nor U7362 (N_7362,N_6983,N_6875);
and U7363 (N_7363,N_6625,N_6920);
nor U7364 (N_7364,N_6961,N_6715);
nor U7365 (N_7365,N_6633,N_6635);
xor U7366 (N_7366,N_6903,N_6811);
xor U7367 (N_7367,N_6890,N_6739);
nor U7368 (N_7368,N_6813,N_6569);
nor U7369 (N_7369,N_6998,N_6586);
xor U7370 (N_7370,N_6828,N_6873);
and U7371 (N_7371,N_6826,N_6507);
nand U7372 (N_7372,N_6618,N_6522);
nor U7373 (N_7373,N_6962,N_6694);
nand U7374 (N_7374,N_6936,N_6994);
or U7375 (N_7375,N_6674,N_6694);
xor U7376 (N_7376,N_6546,N_6714);
and U7377 (N_7377,N_6651,N_6968);
xor U7378 (N_7378,N_6554,N_6941);
xnor U7379 (N_7379,N_6569,N_6765);
nand U7380 (N_7380,N_6840,N_6773);
or U7381 (N_7381,N_6708,N_6542);
nand U7382 (N_7382,N_6953,N_6825);
nand U7383 (N_7383,N_6762,N_6885);
nor U7384 (N_7384,N_6848,N_6902);
or U7385 (N_7385,N_6857,N_6548);
and U7386 (N_7386,N_6924,N_6755);
nand U7387 (N_7387,N_6742,N_6571);
or U7388 (N_7388,N_6776,N_6731);
and U7389 (N_7389,N_6511,N_6910);
or U7390 (N_7390,N_6551,N_6678);
or U7391 (N_7391,N_6696,N_6732);
nand U7392 (N_7392,N_6587,N_6747);
xor U7393 (N_7393,N_6614,N_6945);
nand U7394 (N_7394,N_6980,N_6804);
nor U7395 (N_7395,N_6776,N_6501);
and U7396 (N_7396,N_6646,N_6699);
and U7397 (N_7397,N_6680,N_6632);
xor U7398 (N_7398,N_6786,N_6686);
xor U7399 (N_7399,N_6754,N_6944);
nor U7400 (N_7400,N_6624,N_6810);
nor U7401 (N_7401,N_6987,N_6806);
nor U7402 (N_7402,N_6511,N_6908);
xor U7403 (N_7403,N_6720,N_6663);
and U7404 (N_7404,N_6684,N_6605);
nor U7405 (N_7405,N_6798,N_6530);
xnor U7406 (N_7406,N_6957,N_6829);
or U7407 (N_7407,N_6876,N_6526);
nor U7408 (N_7408,N_6529,N_6945);
xnor U7409 (N_7409,N_6965,N_6831);
nor U7410 (N_7410,N_6884,N_6812);
nor U7411 (N_7411,N_6873,N_6603);
nor U7412 (N_7412,N_6870,N_6525);
xnor U7413 (N_7413,N_6679,N_6747);
nand U7414 (N_7414,N_6940,N_6728);
and U7415 (N_7415,N_6948,N_6934);
nand U7416 (N_7416,N_6728,N_6737);
and U7417 (N_7417,N_6512,N_6782);
and U7418 (N_7418,N_6863,N_6746);
or U7419 (N_7419,N_6897,N_6905);
and U7420 (N_7420,N_6709,N_6986);
xor U7421 (N_7421,N_6582,N_6527);
and U7422 (N_7422,N_6605,N_6680);
nor U7423 (N_7423,N_6881,N_6747);
nor U7424 (N_7424,N_6984,N_6646);
nor U7425 (N_7425,N_6577,N_6915);
and U7426 (N_7426,N_6892,N_6739);
and U7427 (N_7427,N_6756,N_6785);
nand U7428 (N_7428,N_6594,N_6576);
or U7429 (N_7429,N_6916,N_6785);
nor U7430 (N_7430,N_6623,N_6772);
nor U7431 (N_7431,N_6704,N_6504);
nor U7432 (N_7432,N_6821,N_6682);
nor U7433 (N_7433,N_6539,N_6553);
nand U7434 (N_7434,N_6592,N_6635);
and U7435 (N_7435,N_6950,N_6876);
nor U7436 (N_7436,N_6948,N_6517);
nor U7437 (N_7437,N_6664,N_6870);
nand U7438 (N_7438,N_6751,N_6593);
nand U7439 (N_7439,N_6875,N_6917);
nor U7440 (N_7440,N_6970,N_6749);
nand U7441 (N_7441,N_6805,N_6724);
nor U7442 (N_7442,N_6716,N_6693);
and U7443 (N_7443,N_6909,N_6883);
and U7444 (N_7444,N_6635,N_6725);
and U7445 (N_7445,N_6580,N_6771);
and U7446 (N_7446,N_6783,N_6895);
and U7447 (N_7447,N_6730,N_6833);
nor U7448 (N_7448,N_6684,N_6812);
nand U7449 (N_7449,N_6672,N_6773);
nand U7450 (N_7450,N_6573,N_6525);
and U7451 (N_7451,N_6827,N_6629);
nand U7452 (N_7452,N_6753,N_6538);
nor U7453 (N_7453,N_6570,N_6815);
xnor U7454 (N_7454,N_6990,N_6726);
or U7455 (N_7455,N_6872,N_6894);
xnor U7456 (N_7456,N_6752,N_6943);
nor U7457 (N_7457,N_6768,N_6762);
nand U7458 (N_7458,N_6666,N_6737);
and U7459 (N_7459,N_6837,N_6625);
nor U7460 (N_7460,N_6930,N_6634);
or U7461 (N_7461,N_6603,N_6707);
nor U7462 (N_7462,N_6994,N_6968);
xor U7463 (N_7463,N_6849,N_6646);
nor U7464 (N_7464,N_6735,N_6782);
or U7465 (N_7465,N_6784,N_6947);
xor U7466 (N_7466,N_6740,N_6755);
or U7467 (N_7467,N_6668,N_6879);
nor U7468 (N_7468,N_6640,N_6564);
nand U7469 (N_7469,N_6638,N_6698);
nor U7470 (N_7470,N_6724,N_6880);
xnor U7471 (N_7471,N_6618,N_6660);
nor U7472 (N_7472,N_6592,N_6925);
xnor U7473 (N_7473,N_6514,N_6911);
or U7474 (N_7474,N_6954,N_6877);
nor U7475 (N_7475,N_6629,N_6901);
and U7476 (N_7476,N_6706,N_6724);
and U7477 (N_7477,N_6505,N_6671);
and U7478 (N_7478,N_6726,N_6775);
and U7479 (N_7479,N_6689,N_6720);
nor U7480 (N_7480,N_6943,N_6955);
xnor U7481 (N_7481,N_6507,N_6671);
xor U7482 (N_7482,N_6660,N_6576);
nand U7483 (N_7483,N_6759,N_6813);
nand U7484 (N_7484,N_6844,N_6879);
nand U7485 (N_7485,N_6821,N_6556);
nor U7486 (N_7486,N_6648,N_6908);
xor U7487 (N_7487,N_6746,N_6834);
or U7488 (N_7488,N_6721,N_6871);
or U7489 (N_7489,N_6749,N_6981);
nor U7490 (N_7490,N_6856,N_6668);
and U7491 (N_7491,N_6774,N_6855);
or U7492 (N_7492,N_6665,N_6801);
and U7493 (N_7493,N_6840,N_6686);
and U7494 (N_7494,N_6910,N_6723);
xnor U7495 (N_7495,N_6590,N_6503);
nor U7496 (N_7496,N_6782,N_6639);
xor U7497 (N_7497,N_6585,N_6828);
and U7498 (N_7498,N_6578,N_6957);
nor U7499 (N_7499,N_6604,N_6585);
or U7500 (N_7500,N_7421,N_7389);
and U7501 (N_7501,N_7257,N_7364);
xnor U7502 (N_7502,N_7113,N_7050);
nand U7503 (N_7503,N_7101,N_7100);
xor U7504 (N_7504,N_7462,N_7020);
nor U7505 (N_7505,N_7036,N_7185);
or U7506 (N_7506,N_7133,N_7245);
or U7507 (N_7507,N_7067,N_7229);
nand U7508 (N_7508,N_7108,N_7070);
nor U7509 (N_7509,N_7329,N_7148);
or U7510 (N_7510,N_7207,N_7028);
nand U7511 (N_7511,N_7188,N_7231);
or U7512 (N_7512,N_7446,N_7497);
xor U7513 (N_7513,N_7397,N_7477);
nand U7514 (N_7514,N_7013,N_7496);
nand U7515 (N_7515,N_7365,N_7270);
nor U7516 (N_7516,N_7293,N_7177);
nor U7517 (N_7517,N_7000,N_7203);
or U7518 (N_7518,N_7349,N_7415);
nand U7519 (N_7519,N_7011,N_7346);
and U7520 (N_7520,N_7112,N_7413);
nor U7521 (N_7521,N_7247,N_7157);
nand U7522 (N_7522,N_7126,N_7200);
and U7523 (N_7523,N_7033,N_7417);
or U7524 (N_7524,N_7493,N_7407);
and U7525 (N_7525,N_7221,N_7208);
or U7526 (N_7526,N_7281,N_7178);
and U7527 (N_7527,N_7438,N_7353);
or U7528 (N_7528,N_7427,N_7412);
or U7529 (N_7529,N_7102,N_7117);
and U7530 (N_7530,N_7204,N_7418);
xor U7531 (N_7531,N_7330,N_7189);
nor U7532 (N_7532,N_7456,N_7314);
xnor U7533 (N_7533,N_7035,N_7219);
nand U7534 (N_7534,N_7088,N_7287);
xnor U7535 (N_7535,N_7080,N_7408);
and U7536 (N_7536,N_7479,N_7236);
nor U7537 (N_7537,N_7114,N_7468);
nor U7538 (N_7538,N_7403,N_7455);
or U7539 (N_7539,N_7424,N_7395);
or U7540 (N_7540,N_7411,N_7095);
and U7541 (N_7541,N_7366,N_7433);
xor U7542 (N_7542,N_7109,N_7195);
and U7543 (N_7543,N_7288,N_7384);
nand U7544 (N_7544,N_7129,N_7046);
nand U7545 (N_7545,N_7077,N_7124);
nor U7546 (N_7546,N_7472,N_7448);
and U7547 (N_7547,N_7173,N_7171);
or U7548 (N_7548,N_7385,N_7027);
xor U7549 (N_7549,N_7104,N_7425);
or U7550 (N_7550,N_7368,N_7338);
nand U7551 (N_7551,N_7009,N_7322);
and U7552 (N_7552,N_7144,N_7122);
xor U7553 (N_7553,N_7461,N_7409);
or U7554 (N_7554,N_7164,N_7278);
xnor U7555 (N_7555,N_7030,N_7319);
nor U7556 (N_7556,N_7008,N_7042);
and U7557 (N_7557,N_7084,N_7258);
and U7558 (N_7558,N_7280,N_7498);
nor U7559 (N_7559,N_7194,N_7379);
or U7560 (N_7560,N_7051,N_7440);
xor U7561 (N_7561,N_7213,N_7453);
nand U7562 (N_7562,N_7243,N_7037);
and U7563 (N_7563,N_7165,N_7457);
or U7564 (N_7564,N_7224,N_7414);
and U7565 (N_7565,N_7359,N_7056);
xnor U7566 (N_7566,N_7431,N_7169);
nand U7567 (N_7567,N_7459,N_7473);
nand U7568 (N_7568,N_7436,N_7048);
and U7569 (N_7569,N_7172,N_7463);
and U7570 (N_7570,N_7145,N_7449);
xor U7571 (N_7571,N_7094,N_7063);
nor U7572 (N_7572,N_7361,N_7119);
or U7573 (N_7573,N_7211,N_7201);
and U7574 (N_7574,N_7375,N_7140);
nand U7575 (N_7575,N_7347,N_7210);
nand U7576 (N_7576,N_7064,N_7485);
nand U7577 (N_7577,N_7294,N_7125);
and U7578 (N_7578,N_7460,N_7378);
nand U7579 (N_7579,N_7158,N_7218);
nand U7580 (N_7580,N_7285,N_7032);
nor U7581 (N_7581,N_7391,N_7386);
and U7582 (N_7582,N_7167,N_7429);
nor U7583 (N_7583,N_7404,N_7399);
and U7584 (N_7584,N_7297,N_7255);
nand U7585 (N_7585,N_7267,N_7420);
or U7586 (N_7586,N_7494,N_7435);
nand U7587 (N_7587,N_7197,N_7162);
and U7588 (N_7588,N_7332,N_7487);
or U7589 (N_7589,N_7049,N_7107);
and U7590 (N_7590,N_7256,N_7432);
nor U7591 (N_7591,N_7381,N_7470);
or U7592 (N_7592,N_7324,N_7123);
or U7593 (N_7593,N_7437,N_7166);
nand U7594 (N_7594,N_7476,N_7334);
nor U7595 (N_7595,N_7066,N_7301);
xor U7596 (N_7596,N_7342,N_7295);
xnor U7597 (N_7597,N_7458,N_7394);
nor U7598 (N_7598,N_7367,N_7031);
and U7599 (N_7599,N_7306,N_7057);
or U7600 (N_7600,N_7328,N_7223);
and U7601 (N_7601,N_7040,N_7344);
and U7602 (N_7602,N_7303,N_7268);
xor U7603 (N_7603,N_7490,N_7136);
xnor U7604 (N_7604,N_7052,N_7249);
or U7605 (N_7605,N_7312,N_7059);
and U7606 (N_7606,N_7382,N_7376);
nor U7607 (N_7607,N_7333,N_7087);
and U7608 (N_7608,N_7244,N_7209);
and U7609 (N_7609,N_7192,N_7355);
xnor U7610 (N_7610,N_7350,N_7022);
nand U7611 (N_7611,N_7327,N_7043);
nor U7612 (N_7612,N_7062,N_7396);
xnor U7613 (N_7613,N_7469,N_7180);
xor U7614 (N_7614,N_7110,N_7341);
xnor U7615 (N_7615,N_7015,N_7151);
nand U7616 (N_7616,N_7153,N_7152);
nand U7617 (N_7617,N_7098,N_7250);
and U7618 (N_7618,N_7422,N_7426);
xnor U7619 (N_7619,N_7044,N_7454);
nor U7620 (N_7620,N_7358,N_7357);
nor U7621 (N_7621,N_7161,N_7047);
xor U7622 (N_7622,N_7016,N_7186);
nand U7623 (N_7623,N_7466,N_7089);
nand U7624 (N_7624,N_7131,N_7370);
and U7625 (N_7625,N_7193,N_7305);
nor U7626 (N_7626,N_7002,N_7024);
or U7627 (N_7627,N_7121,N_7434);
or U7628 (N_7628,N_7491,N_7277);
or U7629 (N_7629,N_7234,N_7416);
or U7630 (N_7630,N_7082,N_7263);
nor U7631 (N_7631,N_7286,N_7168);
or U7632 (N_7632,N_7388,N_7004);
nor U7633 (N_7633,N_7356,N_7369);
or U7634 (N_7634,N_7387,N_7060);
nor U7635 (N_7635,N_7181,N_7118);
nor U7636 (N_7636,N_7103,N_7068);
nand U7637 (N_7637,N_7139,N_7400);
nor U7638 (N_7638,N_7351,N_7430);
or U7639 (N_7639,N_7091,N_7212);
and U7640 (N_7640,N_7184,N_7475);
nor U7641 (N_7641,N_7191,N_7307);
nor U7642 (N_7642,N_7292,N_7445);
or U7643 (N_7643,N_7354,N_7071);
and U7644 (N_7644,N_7137,N_7127);
and U7645 (N_7645,N_7374,N_7313);
and U7646 (N_7646,N_7105,N_7097);
nand U7647 (N_7647,N_7222,N_7337);
xnor U7648 (N_7648,N_7096,N_7362);
nor U7649 (N_7649,N_7474,N_7065);
or U7650 (N_7650,N_7134,N_7174);
and U7651 (N_7651,N_7111,N_7467);
xnor U7652 (N_7652,N_7183,N_7450);
and U7653 (N_7653,N_7447,N_7072);
xor U7654 (N_7654,N_7055,N_7402);
or U7655 (N_7655,N_7264,N_7239);
or U7656 (N_7656,N_7075,N_7296);
or U7657 (N_7657,N_7282,N_7142);
or U7658 (N_7658,N_7298,N_7225);
nor U7659 (N_7659,N_7340,N_7325);
nand U7660 (N_7660,N_7232,N_7230);
nand U7661 (N_7661,N_7300,N_7116);
and U7662 (N_7662,N_7182,N_7320);
and U7663 (N_7663,N_7423,N_7290);
nor U7664 (N_7664,N_7154,N_7086);
and U7665 (N_7665,N_7299,N_7310);
nor U7666 (N_7666,N_7318,N_7398);
nor U7667 (N_7667,N_7345,N_7138);
nand U7668 (N_7668,N_7315,N_7156);
xnor U7669 (N_7669,N_7214,N_7202);
and U7670 (N_7670,N_7215,N_7226);
nor U7671 (N_7671,N_7465,N_7441);
nor U7672 (N_7672,N_7014,N_7106);
nand U7673 (N_7673,N_7039,N_7343);
xor U7674 (N_7674,N_7034,N_7254);
nand U7675 (N_7675,N_7266,N_7115);
nand U7676 (N_7676,N_7489,N_7003);
nand U7677 (N_7677,N_7309,N_7227);
nor U7678 (N_7678,N_7336,N_7090);
and U7679 (N_7679,N_7316,N_7276);
xor U7680 (N_7680,N_7041,N_7248);
nor U7681 (N_7681,N_7480,N_7005);
nor U7682 (N_7682,N_7198,N_7029);
nor U7683 (N_7683,N_7272,N_7260);
xor U7684 (N_7684,N_7073,N_7007);
and U7685 (N_7685,N_7135,N_7061);
or U7686 (N_7686,N_7228,N_7377);
xor U7687 (N_7687,N_7252,N_7406);
or U7688 (N_7688,N_7099,N_7220);
and U7689 (N_7689,N_7492,N_7352);
nor U7690 (N_7690,N_7069,N_7078);
xnor U7691 (N_7691,N_7235,N_7076);
nor U7692 (N_7692,N_7326,N_7392);
xor U7693 (N_7693,N_7443,N_7196);
nor U7694 (N_7694,N_7241,N_7175);
nor U7695 (N_7695,N_7143,N_7372);
nand U7696 (N_7696,N_7323,N_7373);
nor U7697 (N_7697,N_7471,N_7187);
and U7698 (N_7698,N_7419,N_7302);
and U7699 (N_7699,N_7401,N_7483);
xnor U7700 (N_7700,N_7321,N_7348);
or U7701 (N_7701,N_7464,N_7451);
or U7702 (N_7702,N_7291,N_7311);
nand U7703 (N_7703,N_7289,N_7371);
xnor U7704 (N_7704,N_7120,N_7274);
and U7705 (N_7705,N_7199,N_7275);
and U7706 (N_7706,N_7132,N_7262);
nand U7707 (N_7707,N_7273,N_7006);
or U7708 (N_7708,N_7360,N_7428);
or U7709 (N_7709,N_7159,N_7141);
nand U7710 (N_7710,N_7233,N_7163);
or U7711 (N_7711,N_7246,N_7160);
or U7712 (N_7712,N_7074,N_7149);
nand U7713 (N_7713,N_7486,N_7242);
xor U7714 (N_7714,N_7259,N_7237);
and U7715 (N_7715,N_7058,N_7442);
xor U7716 (N_7716,N_7012,N_7128);
xnor U7717 (N_7717,N_7018,N_7053);
or U7718 (N_7718,N_7484,N_7054);
and U7719 (N_7719,N_7176,N_7083);
nor U7720 (N_7720,N_7216,N_7079);
xor U7721 (N_7721,N_7001,N_7279);
xor U7722 (N_7722,N_7393,N_7085);
xnor U7723 (N_7723,N_7495,N_7045);
and U7724 (N_7724,N_7439,N_7146);
or U7725 (N_7725,N_7025,N_7093);
or U7726 (N_7726,N_7339,N_7478);
nor U7727 (N_7727,N_7238,N_7308);
nor U7728 (N_7728,N_7405,N_7283);
xor U7729 (N_7729,N_7380,N_7410);
and U7730 (N_7730,N_7179,N_7304);
xnor U7731 (N_7731,N_7317,N_7444);
or U7732 (N_7732,N_7251,N_7081);
and U7733 (N_7733,N_7481,N_7452);
nand U7734 (N_7734,N_7261,N_7284);
nand U7735 (N_7735,N_7026,N_7170);
xnor U7736 (N_7736,N_7271,N_7331);
nor U7737 (N_7737,N_7390,N_7010);
nand U7738 (N_7738,N_7147,N_7265);
nor U7739 (N_7739,N_7019,N_7205);
and U7740 (N_7740,N_7269,N_7482);
nand U7741 (N_7741,N_7217,N_7021);
or U7742 (N_7742,N_7017,N_7150);
and U7743 (N_7743,N_7206,N_7092);
xnor U7744 (N_7744,N_7335,N_7190);
nor U7745 (N_7745,N_7155,N_7038);
xor U7746 (N_7746,N_7130,N_7363);
or U7747 (N_7747,N_7253,N_7240);
xnor U7748 (N_7748,N_7023,N_7499);
or U7749 (N_7749,N_7488,N_7383);
nor U7750 (N_7750,N_7413,N_7167);
nor U7751 (N_7751,N_7257,N_7175);
and U7752 (N_7752,N_7094,N_7113);
nor U7753 (N_7753,N_7171,N_7121);
nor U7754 (N_7754,N_7022,N_7444);
and U7755 (N_7755,N_7466,N_7127);
xnor U7756 (N_7756,N_7497,N_7228);
nor U7757 (N_7757,N_7057,N_7029);
or U7758 (N_7758,N_7293,N_7169);
xor U7759 (N_7759,N_7329,N_7326);
or U7760 (N_7760,N_7402,N_7464);
xor U7761 (N_7761,N_7070,N_7460);
nand U7762 (N_7762,N_7049,N_7050);
and U7763 (N_7763,N_7013,N_7088);
or U7764 (N_7764,N_7402,N_7235);
xor U7765 (N_7765,N_7482,N_7095);
and U7766 (N_7766,N_7228,N_7223);
and U7767 (N_7767,N_7310,N_7108);
nand U7768 (N_7768,N_7051,N_7154);
nand U7769 (N_7769,N_7109,N_7436);
nor U7770 (N_7770,N_7345,N_7404);
xnor U7771 (N_7771,N_7213,N_7011);
and U7772 (N_7772,N_7063,N_7272);
or U7773 (N_7773,N_7104,N_7229);
xor U7774 (N_7774,N_7472,N_7313);
nand U7775 (N_7775,N_7030,N_7298);
xor U7776 (N_7776,N_7439,N_7144);
or U7777 (N_7777,N_7444,N_7143);
nor U7778 (N_7778,N_7490,N_7338);
nand U7779 (N_7779,N_7264,N_7421);
nand U7780 (N_7780,N_7030,N_7314);
nand U7781 (N_7781,N_7050,N_7454);
nor U7782 (N_7782,N_7044,N_7205);
or U7783 (N_7783,N_7231,N_7175);
or U7784 (N_7784,N_7478,N_7077);
nand U7785 (N_7785,N_7118,N_7100);
nand U7786 (N_7786,N_7357,N_7263);
and U7787 (N_7787,N_7233,N_7422);
nor U7788 (N_7788,N_7430,N_7395);
nand U7789 (N_7789,N_7489,N_7058);
or U7790 (N_7790,N_7234,N_7206);
nor U7791 (N_7791,N_7254,N_7169);
nor U7792 (N_7792,N_7489,N_7354);
or U7793 (N_7793,N_7309,N_7112);
nand U7794 (N_7794,N_7395,N_7064);
nor U7795 (N_7795,N_7292,N_7135);
nand U7796 (N_7796,N_7285,N_7078);
or U7797 (N_7797,N_7121,N_7230);
xnor U7798 (N_7798,N_7222,N_7156);
nand U7799 (N_7799,N_7018,N_7001);
or U7800 (N_7800,N_7222,N_7164);
nand U7801 (N_7801,N_7060,N_7002);
nand U7802 (N_7802,N_7204,N_7457);
nand U7803 (N_7803,N_7249,N_7293);
nand U7804 (N_7804,N_7231,N_7225);
nand U7805 (N_7805,N_7348,N_7127);
nand U7806 (N_7806,N_7001,N_7036);
nor U7807 (N_7807,N_7094,N_7374);
or U7808 (N_7808,N_7319,N_7495);
and U7809 (N_7809,N_7324,N_7114);
and U7810 (N_7810,N_7393,N_7099);
or U7811 (N_7811,N_7081,N_7457);
xnor U7812 (N_7812,N_7052,N_7150);
xnor U7813 (N_7813,N_7420,N_7215);
nand U7814 (N_7814,N_7149,N_7332);
or U7815 (N_7815,N_7430,N_7228);
and U7816 (N_7816,N_7457,N_7029);
nor U7817 (N_7817,N_7121,N_7317);
nor U7818 (N_7818,N_7474,N_7231);
or U7819 (N_7819,N_7070,N_7340);
nor U7820 (N_7820,N_7337,N_7493);
nor U7821 (N_7821,N_7249,N_7283);
and U7822 (N_7822,N_7276,N_7261);
nor U7823 (N_7823,N_7197,N_7038);
xnor U7824 (N_7824,N_7230,N_7119);
and U7825 (N_7825,N_7029,N_7343);
or U7826 (N_7826,N_7315,N_7292);
xnor U7827 (N_7827,N_7297,N_7305);
or U7828 (N_7828,N_7165,N_7049);
xor U7829 (N_7829,N_7399,N_7388);
nand U7830 (N_7830,N_7149,N_7477);
nand U7831 (N_7831,N_7249,N_7171);
nor U7832 (N_7832,N_7087,N_7470);
nor U7833 (N_7833,N_7346,N_7376);
and U7834 (N_7834,N_7317,N_7346);
xnor U7835 (N_7835,N_7457,N_7069);
or U7836 (N_7836,N_7237,N_7056);
nor U7837 (N_7837,N_7460,N_7385);
and U7838 (N_7838,N_7460,N_7015);
nor U7839 (N_7839,N_7477,N_7040);
and U7840 (N_7840,N_7154,N_7245);
nand U7841 (N_7841,N_7057,N_7216);
nor U7842 (N_7842,N_7352,N_7451);
nor U7843 (N_7843,N_7251,N_7152);
xnor U7844 (N_7844,N_7173,N_7029);
nand U7845 (N_7845,N_7417,N_7100);
nand U7846 (N_7846,N_7040,N_7016);
or U7847 (N_7847,N_7383,N_7082);
xnor U7848 (N_7848,N_7244,N_7103);
xnor U7849 (N_7849,N_7363,N_7175);
nor U7850 (N_7850,N_7310,N_7006);
xnor U7851 (N_7851,N_7305,N_7234);
nand U7852 (N_7852,N_7411,N_7156);
nor U7853 (N_7853,N_7019,N_7356);
or U7854 (N_7854,N_7097,N_7107);
or U7855 (N_7855,N_7353,N_7046);
nor U7856 (N_7856,N_7094,N_7499);
nor U7857 (N_7857,N_7240,N_7039);
nor U7858 (N_7858,N_7435,N_7289);
or U7859 (N_7859,N_7346,N_7368);
nor U7860 (N_7860,N_7381,N_7304);
nand U7861 (N_7861,N_7147,N_7030);
or U7862 (N_7862,N_7456,N_7196);
or U7863 (N_7863,N_7253,N_7477);
and U7864 (N_7864,N_7001,N_7388);
or U7865 (N_7865,N_7196,N_7301);
and U7866 (N_7866,N_7344,N_7401);
nand U7867 (N_7867,N_7221,N_7126);
or U7868 (N_7868,N_7222,N_7172);
nor U7869 (N_7869,N_7473,N_7260);
nor U7870 (N_7870,N_7390,N_7427);
nand U7871 (N_7871,N_7286,N_7022);
nand U7872 (N_7872,N_7060,N_7340);
nand U7873 (N_7873,N_7036,N_7333);
nor U7874 (N_7874,N_7300,N_7123);
nand U7875 (N_7875,N_7083,N_7175);
nand U7876 (N_7876,N_7302,N_7039);
nor U7877 (N_7877,N_7203,N_7454);
nor U7878 (N_7878,N_7457,N_7164);
xor U7879 (N_7879,N_7086,N_7200);
nand U7880 (N_7880,N_7089,N_7080);
or U7881 (N_7881,N_7203,N_7160);
and U7882 (N_7882,N_7266,N_7260);
nand U7883 (N_7883,N_7484,N_7228);
and U7884 (N_7884,N_7239,N_7317);
nand U7885 (N_7885,N_7226,N_7464);
nor U7886 (N_7886,N_7404,N_7351);
or U7887 (N_7887,N_7428,N_7316);
xor U7888 (N_7888,N_7073,N_7312);
xor U7889 (N_7889,N_7249,N_7164);
xor U7890 (N_7890,N_7471,N_7083);
or U7891 (N_7891,N_7337,N_7476);
nand U7892 (N_7892,N_7111,N_7328);
nand U7893 (N_7893,N_7488,N_7093);
nand U7894 (N_7894,N_7196,N_7467);
nor U7895 (N_7895,N_7416,N_7173);
xor U7896 (N_7896,N_7436,N_7035);
and U7897 (N_7897,N_7246,N_7082);
and U7898 (N_7898,N_7466,N_7169);
or U7899 (N_7899,N_7186,N_7317);
or U7900 (N_7900,N_7274,N_7050);
xor U7901 (N_7901,N_7381,N_7369);
or U7902 (N_7902,N_7156,N_7303);
or U7903 (N_7903,N_7188,N_7205);
nand U7904 (N_7904,N_7474,N_7487);
or U7905 (N_7905,N_7401,N_7178);
nand U7906 (N_7906,N_7028,N_7103);
and U7907 (N_7907,N_7191,N_7356);
xnor U7908 (N_7908,N_7284,N_7451);
nand U7909 (N_7909,N_7347,N_7075);
nand U7910 (N_7910,N_7355,N_7081);
and U7911 (N_7911,N_7166,N_7472);
xnor U7912 (N_7912,N_7300,N_7188);
nor U7913 (N_7913,N_7181,N_7094);
xnor U7914 (N_7914,N_7395,N_7440);
xor U7915 (N_7915,N_7390,N_7355);
nor U7916 (N_7916,N_7158,N_7146);
xnor U7917 (N_7917,N_7363,N_7147);
nor U7918 (N_7918,N_7388,N_7094);
and U7919 (N_7919,N_7297,N_7403);
nand U7920 (N_7920,N_7441,N_7197);
nor U7921 (N_7921,N_7342,N_7391);
xor U7922 (N_7922,N_7028,N_7417);
nand U7923 (N_7923,N_7317,N_7307);
xnor U7924 (N_7924,N_7305,N_7238);
nor U7925 (N_7925,N_7261,N_7212);
nand U7926 (N_7926,N_7451,N_7152);
nor U7927 (N_7927,N_7263,N_7322);
and U7928 (N_7928,N_7008,N_7241);
nand U7929 (N_7929,N_7208,N_7487);
nor U7930 (N_7930,N_7064,N_7375);
xnor U7931 (N_7931,N_7450,N_7279);
nand U7932 (N_7932,N_7343,N_7299);
nor U7933 (N_7933,N_7426,N_7237);
nor U7934 (N_7934,N_7286,N_7057);
nand U7935 (N_7935,N_7336,N_7155);
and U7936 (N_7936,N_7311,N_7391);
nor U7937 (N_7937,N_7062,N_7019);
nand U7938 (N_7938,N_7074,N_7133);
or U7939 (N_7939,N_7053,N_7297);
nor U7940 (N_7940,N_7434,N_7324);
xnor U7941 (N_7941,N_7017,N_7374);
xnor U7942 (N_7942,N_7470,N_7449);
or U7943 (N_7943,N_7287,N_7471);
nor U7944 (N_7944,N_7111,N_7072);
xnor U7945 (N_7945,N_7250,N_7376);
and U7946 (N_7946,N_7342,N_7104);
xor U7947 (N_7947,N_7282,N_7136);
nand U7948 (N_7948,N_7283,N_7327);
nor U7949 (N_7949,N_7349,N_7127);
xnor U7950 (N_7950,N_7452,N_7357);
nor U7951 (N_7951,N_7353,N_7262);
or U7952 (N_7952,N_7075,N_7046);
nand U7953 (N_7953,N_7094,N_7482);
xor U7954 (N_7954,N_7345,N_7336);
and U7955 (N_7955,N_7225,N_7218);
nand U7956 (N_7956,N_7327,N_7471);
xnor U7957 (N_7957,N_7213,N_7118);
xor U7958 (N_7958,N_7396,N_7239);
xor U7959 (N_7959,N_7425,N_7219);
nor U7960 (N_7960,N_7120,N_7171);
nand U7961 (N_7961,N_7303,N_7420);
nand U7962 (N_7962,N_7189,N_7451);
nand U7963 (N_7963,N_7325,N_7360);
and U7964 (N_7964,N_7394,N_7271);
nor U7965 (N_7965,N_7482,N_7405);
and U7966 (N_7966,N_7122,N_7060);
nand U7967 (N_7967,N_7315,N_7127);
and U7968 (N_7968,N_7132,N_7427);
xor U7969 (N_7969,N_7359,N_7445);
or U7970 (N_7970,N_7387,N_7111);
xor U7971 (N_7971,N_7009,N_7458);
and U7972 (N_7972,N_7318,N_7174);
nand U7973 (N_7973,N_7175,N_7226);
nor U7974 (N_7974,N_7385,N_7499);
and U7975 (N_7975,N_7473,N_7300);
nand U7976 (N_7976,N_7297,N_7132);
xor U7977 (N_7977,N_7010,N_7111);
nand U7978 (N_7978,N_7135,N_7253);
nand U7979 (N_7979,N_7428,N_7337);
and U7980 (N_7980,N_7023,N_7393);
nand U7981 (N_7981,N_7095,N_7202);
nand U7982 (N_7982,N_7146,N_7166);
and U7983 (N_7983,N_7495,N_7206);
and U7984 (N_7984,N_7244,N_7190);
nand U7985 (N_7985,N_7497,N_7472);
nand U7986 (N_7986,N_7156,N_7114);
nand U7987 (N_7987,N_7210,N_7044);
or U7988 (N_7988,N_7319,N_7313);
or U7989 (N_7989,N_7111,N_7490);
and U7990 (N_7990,N_7141,N_7475);
nand U7991 (N_7991,N_7250,N_7017);
nor U7992 (N_7992,N_7465,N_7365);
or U7993 (N_7993,N_7274,N_7442);
and U7994 (N_7994,N_7445,N_7220);
xnor U7995 (N_7995,N_7359,N_7238);
xor U7996 (N_7996,N_7246,N_7007);
nor U7997 (N_7997,N_7079,N_7318);
nand U7998 (N_7998,N_7241,N_7494);
and U7999 (N_7999,N_7301,N_7035);
and U8000 (N_8000,N_7922,N_7820);
or U8001 (N_8001,N_7905,N_7775);
or U8002 (N_8002,N_7974,N_7863);
nor U8003 (N_8003,N_7948,N_7949);
nand U8004 (N_8004,N_7995,N_7952);
nor U8005 (N_8005,N_7811,N_7998);
nor U8006 (N_8006,N_7515,N_7763);
nor U8007 (N_8007,N_7618,N_7885);
nor U8008 (N_8008,N_7703,N_7676);
or U8009 (N_8009,N_7631,N_7720);
xnor U8010 (N_8010,N_7533,N_7507);
nand U8011 (N_8011,N_7899,N_7656);
nor U8012 (N_8012,N_7535,N_7619);
nand U8013 (N_8013,N_7559,N_7932);
nor U8014 (N_8014,N_7518,N_7887);
nor U8015 (N_8015,N_7610,N_7543);
nor U8016 (N_8016,N_7827,N_7530);
and U8017 (N_8017,N_7510,N_7587);
nor U8018 (N_8018,N_7880,N_7555);
xnor U8019 (N_8019,N_7526,N_7601);
or U8020 (N_8020,N_7879,N_7664);
nor U8021 (N_8021,N_7690,N_7945);
and U8022 (N_8022,N_7910,N_7577);
and U8023 (N_8023,N_7517,N_7634);
and U8024 (N_8024,N_7751,N_7867);
or U8025 (N_8025,N_7911,N_7603);
nor U8026 (N_8026,N_7695,N_7570);
nand U8027 (N_8027,N_7663,N_7638);
xnor U8028 (N_8028,N_7862,N_7883);
xor U8029 (N_8029,N_7781,N_7571);
xor U8030 (N_8030,N_7909,N_7629);
or U8031 (N_8031,N_7602,N_7677);
nor U8032 (N_8032,N_7506,N_7944);
or U8033 (N_8033,N_7897,N_7991);
xor U8034 (N_8034,N_7511,N_7564);
nand U8035 (N_8035,N_7900,N_7585);
nor U8036 (N_8036,N_7693,N_7938);
nor U8037 (N_8037,N_7669,N_7519);
nor U8038 (N_8038,N_7583,N_7620);
xnor U8039 (N_8039,N_7737,N_7660);
nor U8040 (N_8040,N_7626,N_7590);
nand U8041 (N_8041,N_7606,N_7685);
and U8042 (N_8042,N_7710,N_7574);
xnor U8043 (N_8043,N_7914,N_7728);
and U8044 (N_8044,N_7760,N_7904);
nand U8045 (N_8045,N_7734,N_7704);
nor U8046 (N_8046,N_7970,N_7648);
or U8047 (N_8047,N_7962,N_7616);
nand U8048 (N_8048,N_7748,N_7805);
and U8049 (N_8049,N_7908,N_7786);
nor U8050 (N_8050,N_7823,N_7868);
nand U8051 (N_8051,N_7892,N_7836);
nor U8052 (N_8052,N_7912,N_7598);
xor U8053 (N_8053,N_7981,N_7953);
nor U8054 (N_8054,N_7833,N_7858);
and U8055 (N_8055,N_7550,N_7562);
nand U8056 (N_8056,N_7622,N_7803);
nor U8057 (N_8057,N_7984,N_7582);
xnor U8058 (N_8058,N_7770,N_7919);
nor U8059 (N_8059,N_7937,N_7651);
or U8060 (N_8060,N_7873,N_7527);
nor U8061 (N_8061,N_7870,N_7579);
nand U8062 (N_8062,N_7636,N_7850);
or U8063 (N_8063,N_7609,N_7975);
or U8064 (N_8064,N_7627,N_7942);
xor U8065 (N_8065,N_7864,N_7847);
xnor U8066 (N_8066,N_7783,N_7979);
nor U8067 (N_8067,N_7605,N_7642);
and U8068 (N_8068,N_7537,N_7674);
or U8069 (N_8069,N_7572,N_7758);
nand U8070 (N_8070,N_7921,N_7898);
and U8071 (N_8071,N_7988,N_7540);
xor U8072 (N_8072,N_7633,N_7785);
xnor U8073 (N_8073,N_7861,N_7814);
nand U8074 (N_8074,N_7776,N_7986);
xor U8075 (N_8075,N_7662,N_7985);
or U8076 (N_8076,N_7968,N_7874);
or U8077 (N_8077,N_7553,N_7792);
and U8078 (N_8078,N_7683,N_7712);
and U8079 (N_8079,N_7791,N_7554);
xnor U8080 (N_8080,N_7604,N_7790);
nor U8081 (N_8081,N_7966,N_7594);
and U8082 (N_8082,N_7624,N_7658);
nor U8083 (N_8083,N_7615,N_7521);
nand U8084 (N_8084,N_7757,N_7856);
nand U8085 (N_8085,N_7992,N_7614);
and U8086 (N_8086,N_7578,N_7830);
and U8087 (N_8087,N_7976,N_7745);
or U8088 (N_8088,N_7673,N_7713);
xor U8089 (N_8089,N_7933,N_7983);
nand U8090 (N_8090,N_7560,N_7701);
or U8091 (N_8091,N_7961,N_7804);
nor U8092 (N_8092,N_7769,N_7923);
or U8093 (N_8093,N_7520,N_7608);
xnor U8094 (N_8094,N_7588,N_7784);
nor U8095 (N_8095,N_7557,N_7567);
nand U8096 (N_8096,N_7738,N_7934);
nand U8097 (N_8097,N_7671,N_7668);
or U8098 (N_8098,N_7789,N_7741);
nor U8099 (N_8099,N_7566,N_7580);
and U8100 (N_8100,N_7706,N_7955);
or U8101 (N_8101,N_7718,N_7931);
nor U8102 (N_8102,N_7754,N_7581);
xnor U8103 (N_8103,N_7808,N_7759);
xnor U8104 (N_8104,N_7643,N_7607);
or U8105 (N_8105,N_7708,N_7742);
xor U8106 (N_8106,N_7573,N_7552);
and U8107 (N_8107,N_7732,N_7641);
and U8108 (N_8108,N_7716,N_7967);
nand U8109 (N_8109,N_7505,N_7855);
and U8110 (N_8110,N_7999,N_7707);
nand U8111 (N_8111,N_7524,N_7852);
xnor U8112 (N_8112,N_7930,N_7725);
nor U8113 (N_8113,N_7896,N_7628);
or U8114 (N_8114,N_7960,N_7972);
xnor U8115 (N_8115,N_7670,N_7743);
nor U8116 (N_8116,N_7928,N_7698);
nand U8117 (N_8117,N_7876,N_7702);
and U8118 (N_8118,N_7843,N_7508);
nand U8119 (N_8119,N_7592,N_7800);
or U8120 (N_8120,N_7679,N_7875);
xor U8121 (N_8121,N_7964,N_7749);
nor U8122 (N_8122,N_7735,N_7779);
xor U8123 (N_8123,N_7871,N_7584);
nand U8124 (N_8124,N_7514,N_7963);
nor U8125 (N_8125,N_7639,N_7694);
or U8126 (N_8126,N_7829,N_7838);
or U8127 (N_8127,N_7650,N_7652);
xor U8128 (N_8128,N_7840,N_7973);
nor U8129 (N_8129,N_7849,N_7696);
or U8130 (N_8130,N_7727,N_7516);
nor U8131 (N_8131,N_7532,N_7565);
nor U8132 (N_8132,N_7824,N_7882);
and U8133 (N_8133,N_7645,N_7918);
xnor U8134 (N_8134,N_7957,N_7661);
nand U8135 (N_8135,N_7802,N_7859);
and U8136 (N_8136,N_7767,N_7561);
nor U8137 (N_8137,N_7665,N_7913);
xnor U8138 (N_8138,N_7810,N_7680);
nand U8139 (N_8139,N_7726,N_7941);
or U8140 (N_8140,N_7657,N_7625);
or U8141 (N_8141,N_7589,N_7951);
or U8142 (N_8142,N_7649,N_7756);
nor U8143 (N_8143,N_7653,N_7834);
nand U8144 (N_8144,N_7542,N_7819);
nand U8145 (N_8145,N_7854,N_7700);
nand U8146 (N_8146,N_7798,N_7865);
nand U8147 (N_8147,N_7958,N_7746);
nor U8148 (N_8148,N_7654,N_7940);
or U8149 (N_8149,N_7845,N_7901);
nor U8150 (N_8150,N_7612,N_7538);
nand U8151 (N_8151,N_7640,N_7522);
xnor U8152 (N_8152,N_7655,N_7857);
and U8153 (N_8153,N_7807,N_7723);
nor U8154 (N_8154,N_7644,N_7946);
xnor U8155 (N_8155,N_7623,N_7717);
xnor U8156 (N_8156,N_7764,N_7826);
and U8157 (N_8157,N_7549,N_7793);
xor U8158 (N_8158,N_7994,N_7500);
nor U8159 (N_8159,N_7753,N_7780);
or U8160 (N_8160,N_7895,N_7687);
xor U8161 (N_8161,N_7755,N_7548);
or U8162 (N_8162,N_7835,N_7841);
nor U8163 (N_8163,N_7647,N_7886);
and U8164 (N_8164,N_7672,N_7774);
nor U8165 (N_8165,N_7766,N_7576);
nor U8166 (N_8166,N_7730,N_7541);
and U8167 (N_8167,N_7987,N_7722);
or U8168 (N_8168,N_7501,N_7523);
xor U8169 (N_8169,N_7996,N_7551);
and U8170 (N_8170,N_7832,N_7828);
nand U8171 (N_8171,N_7691,N_7632);
or U8172 (N_8172,N_7837,N_7744);
and U8173 (N_8173,N_7599,N_7969);
or U8174 (N_8174,N_7939,N_7545);
nand U8175 (N_8175,N_7721,N_7637);
xor U8176 (N_8176,N_7771,N_7556);
nor U8177 (N_8177,N_7529,N_7926);
nor U8178 (N_8178,N_7575,N_7815);
nand U8179 (N_8179,N_7596,N_7750);
or U8180 (N_8180,N_7684,N_7801);
or U8181 (N_8181,N_7936,N_7740);
nor U8182 (N_8182,N_7736,N_7724);
nand U8183 (N_8183,N_7525,N_7621);
xor U8184 (N_8184,N_7797,N_7893);
and U8185 (N_8185,N_7534,N_7977);
and U8186 (N_8186,N_7682,N_7872);
xor U8187 (N_8187,N_7692,N_7536);
or U8188 (N_8188,N_7697,N_7821);
or U8189 (N_8189,N_7822,N_7956);
or U8190 (N_8190,N_7709,N_7773);
and U8191 (N_8191,N_7890,N_7681);
nand U8192 (N_8192,N_7630,N_7877);
and U8193 (N_8193,N_7729,N_7563);
and U8194 (N_8194,N_7600,N_7782);
nand U8195 (N_8195,N_7711,N_7659);
xor U8196 (N_8196,N_7916,N_7635);
xor U8197 (N_8197,N_7646,N_7731);
nor U8198 (N_8198,N_7593,N_7965);
or U8199 (N_8199,N_7891,N_7569);
or U8200 (N_8200,N_7813,N_7678);
or U8201 (N_8201,N_7539,N_7765);
nand U8202 (N_8202,N_7943,N_7817);
nand U8203 (N_8203,N_7591,N_7611);
nor U8204 (N_8204,N_7839,N_7812);
and U8205 (N_8205,N_7761,N_7917);
or U8206 (N_8206,N_7768,N_7831);
nor U8207 (N_8207,N_7954,N_7795);
and U8208 (N_8208,N_7688,N_7597);
nand U8209 (N_8209,N_7544,N_7915);
nand U8210 (N_8210,N_7705,N_7971);
nand U8211 (N_8211,N_7925,N_7739);
nand U8212 (N_8212,N_7982,N_7686);
or U8213 (N_8213,N_7719,N_7924);
nand U8214 (N_8214,N_7509,N_7818);
nand U8215 (N_8215,N_7902,N_7714);
nand U8216 (N_8216,N_7666,N_7787);
and U8217 (N_8217,N_7950,N_7927);
nor U8218 (N_8218,N_7920,N_7989);
and U8219 (N_8219,N_7869,N_7881);
nor U8220 (N_8220,N_7504,N_7878);
nor U8221 (N_8221,N_7903,N_7667);
or U8222 (N_8222,N_7825,N_7558);
xor U8223 (N_8223,N_7978,N_7853);
xor U8224 (N_8224,N_7595,N_7993);
or U8225 (N_8225,N_7906,N_7947);
xnor U8226 (N_8226,N_7846,N_7513);
nor U8227 (N_8227,N_7568,N_7848);
nand U8228 (N_8228,N_7809,N_7788);
and U8229 (N_8229,N_7547,N_7617);
xor U8230 (N_8230,N_7935,N_7959);
or U8231 (N_8231,N_7546,N_7816);
or U8232 (N_8232,N_7699,N_7586);
and U8233 (N_8233,N_7889,N_7528);
nand U8234 (N_8234,N_7888,N_7777);
xor U8235 (N_8235,N_7715,N_7762);
or U8236 (N_8236,N_7997,N_7844);
xor U8237 (N_8237,N_7778,N_7860);
nand U8238 (N_8238,N_7929,N_7794);
nor U8239 (N_8239,N_7884,N_7733);
xnor U8240 (N_8240,N_7806,N_7866);
nor U8241 (N_8241,N_7796,N_7752);
and U8242 (N_8242,N_7894,N_7689);
or U8243 (N_8243,N_7531,N_7799);
nand U8244 (N_8244,N_7980,N_7675);
nand U8245 (N_8245,N_7747,N_7851);
xnor U8246 (N_8246,N_7613,N_7842);
or U8247 (N_8247,N_7502,N_7990);
or U8248 (N_8248,N_7512,N_7772);
nor U8249 (N_8249,N_7907,N_7503);
or U8250 (N_8250,N_7846,N_7782);
or U8251 (N_8251,N_7791,N_7802);
and U8252 (N_8252,N_7726,N_7826);
or U8253 (N_8253,N_7993,N_7765);
nor U8254 (N_8254,N_7630,N_7945);
nor U8255 (N_8255,N_7571,N_7903);
and U8256 (N_8256,N_7546,N_7997);
nand U8257 (N_8257,N_7594,N_7880);
and U8258 (N_8258,N_7699,N_7657);
and U8259 (N_8259,N_7592,N_7861);
nor U8260 (N_8260,N_7620,N_7896);
and U8261 (N_8261,N_7983,N_7531);
nor U8262 (N_8262,N_7859,N_7586);
nor U8263 (N_8263,N_7823,N_7509);
xor U8264 (N_8264,N_7876,N_7603);
xor U8265 (N_8265,N_7655,N_7964);
xor U8266 (N_8266,N_7867,N_7879);
nand U8267 (N_8267,N_7800,N_7938);
xnor U8268 (N_8268,N_7722,N_7731);
or U8269 (N_8269,N_7971,N_7552);
and U8270 (N_8270,N_7945,N_7774);
and U8271 (N_8271,N_7851,N_7952);
and U8272 (N_8272,N_7901,N_7695);
nand U8273 (N_8273,N_7582,N_7650);
or U8274 (N_8274,N_7863,N_7829);
nand U8275 (N_8275,N_7867,N_7758);
nand U8276 (N_8276,N_7605,N_7627);
xor U8277 (N_8277,N_7906,N_7588);
and U8278 (N_8278,N_7719,N_7881);
xnor U8279 (N_8279,N_7931,N_7752);
nand U8280 (N_8280,N_7538,N_7704);
nand U8281 (N_8281,N_7625,N_7515);
or U8282 (N_8282,N_7607,N_7587);
xor U8283 (N_8283,N_7754,N_7826);
nand U8284 (N_8284,N_7691,N_7908);
or U8285 (N_8285,N_7783,N_7801);
nor U8286 (N_8286,N_7712,N_7707);
and U8287 (N_8287,N_7699,N_7995);
or U8288 (N_8288,N_7773,N_7755);
and U8289 (N_8289,N_7593,N_7782);
or U8290 (N_8290,N_7933,N_7945);
or U8291 (N_8291,N_7715,N_7580);
nand U8292 (N_8292,N_7751,N_7950);
xor U8293 (N_8293,N_7876,N_7849);
or U8294 (N_8294,N_7900,N_7610);
nand U8295 (N_8295,N_7600,N_7726);
or U8296 (N_8296,N_7726,N_7639);
xor U8297 (N_8297,N_7705,N_7843);
or U8298 (N_8298,N_7657,N_7576);
and U8299 (N_8299,N_7682,N_7857);
nor U8300 (N_8300,N_7643,N_7616);
xor U8301 (N_8301,N_7541,N_7849);
and U8302 (N_8302,N_7946,N_7573);
nand U8303 (N_8303,N_7764,N_7590);
nor U8304 (N_8304,N_7647,N_7928);
nor U8305 (N_8305,N_7943,N_7816);
xnor U8306 (N_8306,N_7700,N_7926);
nand U8307 (N_8307,N_7812,N_7977);
xor U8308 (N_8308,N_7653,N_7532);
or U8309 (N_8309,N_7997,N_7653);
nand U8310 (N_8310,N_7823,N_7922);
or U8311 (N_8311,N_7844,N_7505);
and U8312 (N_8312,N_7512,N_7962);
nor U8313 (N_8313,N_7558,N_7856);
xnor U8314 (N_8314,N_7636,N_7692);
nand U8315 (N_8315,N_7851,N_7988);
nand U8316 (N_8316,N_7988,N_7770);
nor U8317 (N_8317,N_7984,N_7629);
and U8318 (N_8318,N_7941,N_7745);
nor U8319 (N_8319,N_7655,N_7846);
or U8320 (N_8320,N_7827,N_7695);
nor U8321 (N_8321,N_7692,N_7561);
xor U8322 (N_8322,N_7774,N_7568);
nor U8323 (N_8323,N_7856,N_7892);
and U8324 (N_8324,N_7948,N_7666);
or U8325 (N_8325,N_7618,N_7580);
and U8326 (N_8326,N_7583,N_7618);
nand U8327 (N_8327,N_7568,N_7920);
nor U8328 (N_8328,N_7578,N_7626);
xor U8329 (N_8329,N_7871,N_7646);
or U8330 (N_8330,N_7805,N_7957);
xnor U8331 (N_8331,N_7597,N_7786);
xnor U8332 (N_8332,N_7844,N_7722);
and U8333 (N_8333,N_7926,N_7848);
nor U8334 (N_8334,N_7993,N_7636);
xnor U8335 (N_8335,N_7631,N_7518);
or U8336 (N_8336,N_7559,N_7766);
and U8337 (N_8337,N_7749,N_7981);
and U8338 (N_8338,N_7714,N_7873);
nand U8339 (N_8339,N_7906,N_7724);
nor U8340 (N_8340,N_7814,N_7538);
or U8341 (N_8341,N_7785,N_7579);
or U8342 (N_8342,N_7678,N_7543);
nand U8343 (N_8343,N_7956,N_7878);
or U8344 (N_8344,N_7536,N_7591);
or U8345 (N_8345,N_7667,N_7657);
and U8346 (N_8346,N_7637,N_7948);
nor U8347 (N_8347,N_7768,N_7543);
and U8348 (N_8348,N_7713,N_7734);
or U8349 (N_8349,N_7659,N_7821);
nor U8350 (N_8350,N_7775,N_7802);
xor U8351 (N_8351,N_7522,N_7775);
and U8352 (N_8352,N_7663,N_7547);
nor U8353 (N_8353,N_7945,N_7961);
nor U8354 (N_8354,N_7522,N_7647);
nand U8355 (N_8355,N_7502,N_7770);
nor U8356 (N_8356,N_7613,N_7720);
nor U8357 (N_8357,N_7751,N_7511);
or U8358 (N_8358,N_7618,N_7986);
and U8359 (N_8359,N_7693,N_7827);
xnor U8360 (N_8360,N_7883,N_7655);
nand U8361 (N_8361,N_7523,N_7966);
or U8362 (N_8362,N_7926,N_7991);
or U8363 (N_8363,N_7713,N_7504);
and U8364 (N_8364,N_7974,N_7706);
nand U8365 (N_8365,N_7709,N_7887);
or U8366 (N_8366,N_7701,N_7621);
and U8367 (N_8367,N_7965,N_7530);
or U8368 (N_8368,N_7510,N_7600);
or U8369 (N_8369,N_7841,N_7712);
nor U8370 (N_8370,N_7936,N_7718);
nor U8371 (N_8371,N_7903,N_7590);
or U8372 (N_8372,N_7751,N_7622);
or U8373 (N_8373,N_7798,N_7976);
xor U8374 (N_8374,N_7868,N_7624);
or U8375 (N_8375,N_7580,N_7688);
or U8376 (N_8376,N_7827,N_7538);
and U8377 (N_8377,N_7930,N_7906);
nor U8378 (N_8378,N_7855,N_7818);
nor U8379 (N_8379,N_7675,N_7992);
xnor U8380 (N_8380,N_7510,N_7703);
or U8381 (N_8381,N_7599,N_7703);
nand U8382 (N_8382,N_7786,N_7613);
or U8383 (N_8383,N_7783,N_7769);
and U8384 (N_8384,N_7790,N_7987);
nor U8385 (N_8385,N_7575,N_7831);
and U8386 (N_8386,N_7579,N_7587);
and U8387 (N_8387,N_7811,N_7824);
or U8388 (N_8388,N_7645,N_7765);
xnor U8389 (N_8389,N_7839,N_7580);
or U8390 (N_8390,N_7705,N_7647);
xor U8391 (N_8391,N_7762,N_7688);
and U8392 (N_8392,N_7761,N_7536);
or U8393 (N_8393,N_7994,N_7941);
xnor U8394 (N_8394,N_7826,N_7920);
nor U8395 (N_8395,N_7558,N_7855);
nand U8396 (N_8396,N_7939,N_7807);
xor U8397 (N_8397,N_7611,N_7828);
xor U8398 (N_8398,N_7730,N_7789);
or U8399 (N_8399,N_7792,N_7797);
or U8400 (N_8400,N_7886,N_7834);
nand U8401 (N_8401,N_7723,N_7830);
nand U8402 (N_8402,N_7583,N_7640);
or U8403 (N_8403,N_7892,N_7796);
nor U8404 (N_8404,N_7608,N_7808);
nand U8405 (N_8405,N_7873,N_7628);
xnor U8406 (N_8406,N_7853,N_7532);
xnor U8407 (N_8407,N_7758,N_7811);
xor U8408 (N_8408,N_7925,N_7982);
xor U8409 (N_8409,N_7988,N_7949);
nand U8410 (N_8410,N_7520,N_7796);
xor U8411 (N_8411,N_7704,N_7788);
nor U8412 (N_8412,N_7652,N_7568);
xor U8413 (N_8413,N_7911,N_7817);
nand U8414 (N_8414,N_7547,N_7976);
nand U8415 (N_8415,N_7859,N_7978);
nand U8416 (N_8416,N_7770,N_7735);
nor U8417 (N_8417,N_7694,N_7825);
xor U8418 (N_8418,N_7880,N_7845);
nand U8419 (N_8419,N_7961,N_7767);
xnor U8420 (N_8420,N_7968,N_7779);
nand U8421 (N_8421,N_7541,N_7961);
xor U8422 (N_8422,N_7528,N_7827);
nor U8423 (N_8423,N_7889,N_7814);
nand U8424 (N_8424,N_7739,N_7666);
xnor U8425 (N_8425,N_7678,N_7811);
xor U8426 (N_8426,N_7655,N_7949);
and U8427 (N_8427,N_7674,N_7966);
xnor U8428 (N_8428,N_7539,N_7515);
nand U8429 (N_8429,N_7551,N_7886);
or U8430 (N_8430,N_7888,N_7535);
or U8431 (N_8431,N_7776,N_7993);
xor U8432 (N_8432,N_7801,N_7533);
xor U8433 (N_8433,N_7689,N_7700);
nand U8434 (N_8434,N_7952,N_7507);
or U8435 (N_8435,N_7628,N_7776);
and U8436 (N_8436,N_7743,N_7649);
nor U8437 (N_8437,N_7725,N_7903);
xor U8438 (N_8438,N_7963,N_7533);
nand U8439 (N_8439,N_7916,N_7652);
or U8440 (N_8440,N_7885,N_7899);
xor U8441 (N_8441,N_7612,N_7951);
nand U8442 (N_8442,N_7520,N_7541);
and U8443 (N_8443,N_7850,N_7564);
nand U8444 (N_8444,N_7984,N_7799);
nor U8445 (N_8445,N_7747,N_7846);
or U8446 (N_8446,N_7973,N_7991);
or U8447 (N_8447,N_7825,N_7515);
nand U8448 (N_8448,N_7535,N_7558);
and U8449 (N_8449,N_7974,N_7895);
xnor U8450 (N_8450,N_7768,N_7544);
nand U8451 (N_8451,N_7576,N_7913);
or U8452 (N_8452,N_7531,N_7688);
or U8453 (N_8453,N_7728,N_7912);
or U8454 (N_8454,N_7980,N_7631);
and U8455 (N_8455,N_7674,N_7518);
nand U8456 (N_8456,N_7690,N_7758);
and U8457 (N_8457,N_7919,N_7653);
and U8458 (N_8458,N_7958,N_7869);
nand U8459 (N_8459,N_7853,N_7684);
or U8460 (N_8460,N_7990,N_7824);
xnor U8461 (N_8461,N_7819,N_7844);
or U8462 (N_8462,N_7544,N_7621);
nor U8463 (N_8463,N_7723,N_7675);
and U8464 (N_8464,N_7629,N_7648);
nand U8465 (N_8465,N_7829,N_7842);
xor U8466 (N_8466,N_7838,N_7517);
or U8467 (N_8467,N_7815,N_7738);
xor U8468 (N_8468,N_7685,N_7849);
nor U8469 (N_8469,N_7702,N_7657);
nand U8470 (N_8470,N_7662,N_7965);
nand U8471 (N_8471,N_7954,N_7969);
and U8472 (N_8472,N_7771,N_7984);
xnor U8473 (N_8473,N_7962,N_7685);
nor U8474 (N_8474,N_7985,N_7698);
nor U8475 (N_8475,N_7729,N_7780);
xor U8476 (N_8476,N_7604,N_7555);
nor U8477 (N_8477,N_7536,N_7531);
nand U8478 (N_8478,N_7691,N_7564);
nand U8479 (N_8479,N_7502,N_7808);
or U8480 (N_8480,N_7588,N_7995);
and U8481 (N_8481,N_7843,N_7947);
and U8482 (N_8482,N_7980,N_7796);
nor U8483 (N_8483,N_7748,N_7548);
and U8484 (N_8484,N_7662,N_7647);
and U8485 (N_8485,N_7865,N_7818);
nor U8486 (N_8486,N_7916,N_7699);
or U8487 (N_8487,N_7594,N_7637);
xnor U8488 (N_8488,N_7733,N_7886);
or U8489 (N_8489,N_7500,N_7624);
nand U8490 (N_8490,N_7803,N_7781);
or U8491 (N_8491,N_7820,N_7794);
xnor U8492 (N_8492,N_7531,N_7917);
and U8493 (N_8493,N_7686,N_7818);
or U8494 (N_8494,N_7648,N_7839);
or U8495 (N_8495,N_7931,N_7577);
nand U8496 (N_8496,N_7898,N_7998);
and U8497 (N_8497,N_7921,N_7674);
nand U8498 (N_8498,N_7937,N_7595);
or U8499 (N_8499,N_7831,N_7879);
xor U8500 (N_8500,N_8319,N_8256);
or U8501 (N_8501,N_8291,N_8282);
xor U8502 (N_8502,N_8062,N_8204);
nand U8503 (N_8503,N_8158,N_8166);
xor U8504 (N_8504,N_8492,N_8181);
and U8505 (N_8505,N_8242,N_8091);
xor U8506 (N_8506,N_8023,N_8090);
nand U8507 (N_8507,N_8359,N_8097);
and U8508 (N_8508,N_8325,N_8132);
or U8509 (N_8509,N_8495,N_8483);
nand U8510 (N_8510,N_8419,N_8234);
nand U8511 (N_8511,N_8338,N_8077);
xor U8512 (N_8512,N_8043,N_8425);
nand U8513 (N_8513,N_8450,N_8306);
nand U8514 (N_8514,N_8134,N_8197);
and U8515 (N_8515,N_8330,N_8129);
xnor U8516 (N_8516,N_8124,N_8277);
nor U8517 (N_8517,N_8164,N_8210);
xor U8518 (N_8518,N_8001,N_8030);
nand U8519 (N_8519,N_8014,N_8012);
nor U8520 (N_8520,N_8060,N_8047);
or U8521 (N_8521,N_8460,N_8276);
nor U8522 (N_8522,N_8286,N_8408);
nor U8523 (N_8523,N_8052,N_8123);
nand U8524 (N_8524,N_8447,N_8035);
nand U8525 (N_8525,N_8120,N_8163);
and U8526 (N_8526,N_8195,N_8233);
nor U8527 (N_8527,N_8322,N_8037);
nand U8528 (N_8528,N_8323,N_8347);
nand U8529 (N_8529,N_8493,N_8315);
nand U8530 (N_8530,N_8041,N_8415);
or U8531 (N_8531,N_8212,N_8200);
nand U8532 (N_8532,N_8384,N_8290);
and U8533 (N_8533,N_8026,N_8364);
nor U8534 (N_8534,N_8059,N_8240);
nand U8535 (N_8535,N_8321,N_8292);
nor U8536 (N_8536,N_8346,N_8314);
and U8537 (N_8537,N_8183,N_8382);
or U8538 (N_8538,N_8002,N_8112);
nor U8539 (N_8539,N_8395,N_8165);
nor U8540 (N_8540,N_8236,N_8295);
nor U8541 (N_8541,N_8173,N_8377);
or U8542 (N_8542,N_8016,N_8497);
or U8543 (N_8543,N_8433,N_8046);
xor U8544 (N_8544,N_8003,N_8151);
or U8545 (N_8545,N_8273,N_8309);
and U8546 (N_8546,N_8318,N_8157);
xor U8547 (N_8547,N_8106,N_8435);
nand U8548 (N_8548,N_8288,N_8140);
and U8549 (N_8549,N_8413,N_8417);
nor U8550 (N_8550,N_8099,N_8180);
xor U8551 (N_8551,N_8471,N_8142);
and U8552 (N_8552,N_8403,N_8362);
nor U8553 (N_8553,N_8088,N_8156);
and U8554 (N_8554,N_8392,N_8011);
xnor U8555 (N_8555,N_8479,N_8018);
nand U8556 (N_8556,N_8264,N_8215);
xor U8557 (N_8557,N_8159,N_8462);
nand U8558 (N_8558,N_8044,N_8407);
and U8559 (N_8559,N_8125,N_8285);
nand U8560 (N_8560,N_8143,N_8228);
and U8561 (N_8561,N_8130,N_8485);
or U8562 (N_8562,N_8452,N_8335);
or U8563 (N_8563,N_8174,N_8207);
nand U8564 (N_8564,N_8464,N_8482);
xor U8565 (N_8565,N_8138,N_8101);
and U8566 (N_8566,N_8305,N_8353);
nand U8567 (N_8567,N_8310,N_8496);
xnor U8568 (N_8568,N_8094,N_8354);
or U8569 (N_8569,N_8071,N_8297);
xor U8570 (N_8570,N_8294,N_8127);
nand U8571 (N_8571,N_8349,N_8188);
xor U8572 (N_8572,N_8472,N_8186);
or U8573 (N_8573,N_8465,N_8056);
nand U8574 (N_8574,N_8401,N_8213);
and U8575 (N_8575,N_8487,N_8469);
nor U8576 (N_8576,N_8051,N_8214);
or U8577 (N_8577,N_8102,N_8316);
nor U8578 (N_8578,N_8024,N_8253);
and U8579 (N_8579,N_8061,N_8036);
nand U8580 (N_8580,N_8406,N_8383);
or U8581 (N_8581,N_8414,N_8182);
and U8582 (N_8582,N_8045,N_8474);
and U8583 (N_8583,N_8098,N_8089);
nand U8584 (N_8584,N_8266,N_8144);
and U8585 (N_8585,N_8378,N_8000);
or U8586 (N_8586,N_8070,N_8375);
nand U8587 (N_8587,N_8289,N_8179);
nand U8588 (N_8588,N_8201,N_8437);
and U8589 (N_8589,N_8410,N_8239);
nor U8590 (N_8590,N_8092,N_8491);
or U8591 (N_8591,N_8385,N_8248);
xor U8592 (N_8592,N_8176,N_8178);
nor U8593 (N_8593,N_8072,N_8454);
nand U8594 (N_8594,N_8154,N_8387);
xnor U8595 (N_8595,N_8170,N_8081);
xnor U8596 (N_8596,N_8287,N_8128);
nor U8597 (N_8597,N_8177,N_8416);
nor U8598 (N_8598,N_8146,N_8339);
and U8599 (N_8599,N_8326,N_8426);
xor U8600 (N_8600,N_8267,N_8303);
nand U8601 (N_8601,N_8396,N_8473);
nand U8602 (N_8602,N_8342,N_8107);
nand U8603 (N_8603,N_8459,N_8455);
or U8604 (N_8604,N_8031,N_8079);
and U8605 (N_8605,N_8033,N_8265);
or U8606 (N_8606,N_8246,N_8067);
or U8607 (N_8607,N_8196,N_8263);
nand U8608 (N_8608,N_8117,N_8149);
or U8609 (N_8609,N_8331,N_8320);
nand U8610 (N_8610,N_8367,N_8221);
and U8611 (N_8611,N_8225,N_8218);
nand U8612 (N_8612,N_8076,N_8463);
nand U8613 (N_8613,N_8069,N_8270);
and U8614 (N_8614,N_8086,N_8017);
xnor U8615 (N_8615,N_8252,N_8066);
xor U8616 (N_8616,N_8477,N_8442);
nand U8617 (N_8617,N_8422,N_8202);
or U8618 (N_8618,N_8481,N_8148);
xor U8619 (N_8619,N_8490,N_8006);
or U8620 (N_8620,N_8308,N_8343);
or U8621 (N_8621,N_8110,N_8039);
xor U8622 (N_8622,N_8301,N_8184);
or U8623 (N_8623,N_8451,N_8281);
nor U8624 (N_8624,N_8073,N_8013);
nand U8625 (N_8625,N_8255,N_8208);
xor U8626 (N_8626,N_8230,N_8082);
or U8627 (N_8627,N_8131,N_8393);
or U8628 (N_8628,N_8361,N_8488);
xnor U8629 (N_8629,N_8296,N_8366);
xor U8630 (N_8630,N_8074,N_8103);
xor U8631 (N_8631,N_8280,N_8025);
and U8632 (N_8632,N_8399,N_8299);
nand U8633 (N_8633,N_8475,N_8019);
or U8634 (N_8634,N_8008,N_8257);
and U8635 (N_8635,N_8429,N_8022);
xor U8636 (N_8636,N_8038,N_8358);
and U8637 (N_8637,N_8217,N_8205);
and U8638 (N_8638,N_8311,N_8411);
xor U8639 (N_8639,N_8021,N_8100);
nor U8640 (N_8640,N_8423,N_8075);
xor U8641 (N_8641,N_8443,N_8027);
nand U8642 (N_8642,N_8193,N_8004);
nand U8643 (N_8643,N_8055,N_8199);
xnor U8644 (N_8644,N_8211,N_8445);
or U8645 (N_8645,N_8268,N_8198);
xnor U8646 (N_8646,N_8484,N_8247);
nand U8647 (N_8647,N_8390,N_8085);
xor U8648 (N_8648,N_8348,N_8351);
nor U8649 (N_8649,N_8334,N_8337);
or U8650 (N_8650,N_8380,N_8336);
and U8651 (N_8651,N_8250,N_8093);
and U8652 (N_8652,N_8262,N_8145);
and U8653 (N_8653,N_8227,N_8409);
xor U8654 (N_8654,N_8114,N_8418);
nor U8655 (N_8655,N_8078,N_8350);
and U8656 (N_8656,N_8150,N_8456);
nor U8657 (N_8657,N_8175,N_8470);
and U8658 (N_8658,N_8424,N_8357);
nand U8659 (N_8659,N_8254,N_8137);
or U8660 (N_8660,N_8356,N_8376);
and U8661 (N_8661,N_8345,N_8064);
or U8662 (N_8662,N_8042,N_8034);
or U8663 (N_8663,N_8104,N_8440);
nor U8664 (N_8664,N_8293,N_8054);
and U8665 (N_8665,N_8152,N_8121);
nand U8666 (N_8666,N_8049,N_8048);
and U8667 (N_8667,N_8421,N_8083);
nand U8668 (N_8668,N_8096,N_8087);
xor U8669 (N_8669,N_8275,N_8448);
nand U8670 (N_8670,N_8369,N_8223);
xnor U8671 (N_8671,N_8122,N_8374);
nand U8672 (N_8672,N_8160,N_8352);
nand U8673 (N_8673,N_8084,N_8009);
or U8674 (N_8674,N_8189,N_8172);
or U8675 (N_8675,N_8269,N_8458);
nand U8676 (N_8676,N_8259,N_8381);
xnor U8677 (N_8677,N_8139,N_8206);
nand U8678 (N_8678,N_8260,N_8203);
and U8679 (N_8679,N_8489,N_8040);
nor U8680 (N_8680,N_8258,N_8105);
nor U8681 (N_8681,N_8371,N_8020);
and U8682 (N_8682,N_8224,N_8300);
nor U8683 (N_8683,N_8453,N_8115);
nor U8684 (N_8684,N_8058,N_8389);
or U8685 (N_8685,N_8355,N_8222);
or U8686 (N_8686,N_8340,N_8312);
or U8687 (N_8687,N_8427,N_8438);
and U8688 (N_8688,N_8015,N_8360);
nand U8689 (N_8689,N_8219,N_8141);
nand U8690 (N_8690,N_8232,N_8398);
or U8691 (N_8691,N_8284,N_8251);
nand U8692 (N_8692,N_8405,N_8153);
nand U8693 (N_8693,N_8431,N_8461);
nand U8694 (N_8694,N_8192,N_8397);
nor U8695 (N_8695,N_8190,N_8328);
or U8696 (N_8696,N_8185,N_8118);
or U8697 (N_8697,N_8368,N_8272);
nand U8698 (N_8698,N_8394,N_8313);
and U8699 (N_8699,N_8373,N_8231);
and U8700 (N_8700,N_8332,N_8444);
nand U8701 (N_8701,N_8053,N_8480);
nor U8702 (N_8702,N_8498,N_8029);
and U8703 (N_8703,N_8274,N_8057);
nor U8704 (N_8704,N_8109,N_8468);
or U8705 (N_8705,N_8344,N_8261);
nand U8706 (N_8706,N_8441,N_8333);
nand U8707 (N_8707,N_8111,N_8370);
nor U8708 (N_8708,N_8283,N_8449);
xnor U8709 (N_8709,N_8065,N_8028);
or U8710 (N_8710,N_8007,N_8317);
and U8711 (N_8711,N_8457,N_8155);
xor U8712 (N_8712,N_8327,N_8229);
and U8713 (N_8713,N_8278,N_8379);
and U8714 (N_8714,N_8068,N_8476);
xor U8715 (N_8715,N_8119,N_8432);
nand U8716 (N_8716,N_8271,N_8412);
or U8717 (N_8717,N_8436,N_8032);
or U8718 (N_8718,N_8428,N_8095);
and U8719 (N_8719,N_8279,N_8434);
xor U8720 (N_8720,N_8363,N_8220);
and U8721 (N_8721,N_8244,N_8402);
and U8722 (N_8722,N_8446,N_8167);
xnor U8723 (N_8723,N_8187,N_8400);
xnor U8724 (N_8724,N_8194,N_8245);
or U8725 (N_8725,N_8478,N_8050);
nor U8726 (N_8726,N_8171,N_8365);
and U8727 (N_8727,N_8386,N_8209);
nor U8728 (N_8728,N_8241,N_8191);
and U8729 (N_8729,N_8494,N_8126);
xnor U8730 (N_8730,N_8237,N_8168);
nand U8731 (N_8731,N_8216,N_8133);
nor U8732 (N_8732,N_8388,N_8302);
or U8733 (N_8733,N_8430,N_8169);
or U8734 (N_8734,N_8238,N_8439);
and U8735 (N_8735,N_8298,N_8486);
and U8736 (N_8736,N_8304,N_8329);
or U8737 (N_8737,N_8391,N_8226);
nand U8738 (N_8738,N_8499,N_8147);
nand U8739 (N_8739,N_8235,N_8467);
xnor U8740 (N_8740,N_8108,N_8372);
nand U8741 (N_8741,N_8113,N_8080);
nor U8742 (N_8742,N_8136,N_8249);
or U8743 (N_8743,N_8005,N_8307);
and U8744 (N_8744,N_8420,N_8404);
nand U8745 (N_8745,N_8135,N_8161);
or U8746 (N_8746,N_8162,N_8466);
nor U8747 (N_8747,N_8324,N_8063);
xor U8748 (N_8748,N_8010,N_8341);
xnor U8749 (N_8749,N_8116,N_8243);
and U8750 (N_8750,N_8448,N_8465);
xnor U8751 (N_8751,N_8134,N_8481);
xnor U8752 (N_8752,N_8197,N_8190);
nor U8753 (N_8753,N_8185,N_8353);
xor U8754 (N_8754,N_8210,N_8117);
nor U8755 (N_8755,N_8356,N_8475);
or U8756 (N_8756,N_8037,N_8064);
xor U8757 (N_8757,N_8489,N_8224);
nor U8758 (N_8758,N_8423,N_8086);
xor U8759 (N_8759,N_8423,N_8370);
or U8760 (N_8760,N_8281,N_8496);
or U8761 (N_8761,N_8357,N_8367);
xnor U8762 (N_8762,N_8368,N_8150);
nor U8763 (N_8763,N_8071,N_8220);
nor U8764 (N_8764,N_8230,N_8221);
or U8765 (N_8765,N_8403,N_8212);
or U8766 (N_8766,N_8016,N_8367);
or U8767 (N_8767,N_8046,N_8099);
nand U8768 (N_8768,N_8490,N_8319);
nand U8769 (N_8769,N_8337,N_8346);
nand U8770 (N_8770,N_8397,N_8337);
xnor U8771 (N_8771,N_8045,N_8350);
xnor U8772 (N_8772,N_8418,N_8046);
nand U8773 (N_8773,N_8382,N_8127);
or U8774 (N_8774,N_8487,N_8097);
nand U8775 (N_8775,N_8259,N_8179);
nand U8776 (N_8776,N_8311,N_8094);
or U8777 (N_8777,N_8488,N_8111);
and U8778 (N_8778,N_8364,N_8369);
or U8779 (N_8779,N_8005,N_8358);
nor U8780 (N_8780,N_8420,N_8304);
nand U8781 (N_8781,N_8317,N_8207);
nor U8782 (N_8782,N_8269,N_8355);
xor U8783 (N_8783,N_8311,N_8318);
xor U8784 (N_8784,N_8323,N_8384);
xnor U8785 (N_8785,N_8167,N_8485);
nand U8786 (N_8786,N_8406,N_8288);
or U8787 (N_8787,N_8228,N_8414);
nand U8788 (N_8788,N_8002,N_8462);
xor U8789 (N_8789,N_8333,N_8374);
xnor U8790 (N_8790,N_8148,N_8373);
and U8791 (N_8791,N_8082,N_8211);
or U8792 (N_8792,N_8301,N_8205);
or U8793 (N_8793,N_8439,N_8315);
and U8794 (N_8794,N_8026,N_8224);
nand U8795 (N_8795,N_8120,N_8365);
or U8796 (N_8796,N_8185,N_8404);
nand U8797 (N_8797,N_8351,N_8494);
xor U8798 (N_8798,N_8371,N_8390);
nor U8799 (N_8799,N_8281,N_8093);
nand U8800 (N_8800,N_8137,N_8370);
or U8801 (N_8801,N_8179,N_8181);
and U8802 (N_8802,N_8065,N_8210);
xor U8803 (N_8803,N_8200,N_8113);
nor U8804 (N_8804,N_8159,N_8311);
xor U8805 (N_8805,N_8491,N_8405);
and U8806 (N_8806,N_8370,N_8108);
nand U8807 (N_8807,N_8209,N_8258);
xnor U8808 (N_8808,N_8433,N_8189);
and U8809 (N_8809,N_8007,N_8334);
xor U8810 (N_8810,N_8154,N_8069);
or U8811 (N_8811,N_8427,N_8089);
and U8812 (N_8812,N_8125,N_8278);
or U8813 (N_8813,N_8468,N_8370);
xnor U8814 (N_8814,N_8048,N_8046);
nor U8815 (N_8815,N_8037,N_8153);
or U8816 (N_8816,N_8050,N_8170);
nor U8817 (N_8817,N_8267,N_8404);
nand U8818 (N_8818,N_8056,N_8499);
or U8819 (N_8819,N_8240,N_8174);
and U8820 (N_8820,N_8041,N_8358);
nand U8821 (N_8821,N_8358,N_8174);
xor U8822 (N_8822,N_8224,N_8462);
nor U8823 (N_8823,N_8300,N_8052);
nand U8824 (N_8824,N_8429,N_8205);
or U8825 (N_8825,N_8007,N_8145);
nor U8826 (N_8826,N_8180,N_8088);
or U8827 (N_8827,N_8122,N_8190);
xnor U8828 (N_8828,N_8233,N_8368);
or U8829 (N_8829,N_8423,N_8194);
or U8830 (N_8830,N_8496,N_8449);
nor U8831 (N_8831,N_8275,N_8475);
nand U8832 (N_8832,N_8219,N_8380);
nor U8833 (N_8833,N_8049,N_8072);
and U8834 (N_8834,N_8241,N_8083);
or U8835 (N_8835,N_8229,N_8087);
nor U8836 (N_8836,N_8056,N_8207);
and U8837 (N_8837,N_8393,N_8093);
xnor U8838 (N_8838,N_8411,N_8354);
and U8839 (N_8839,N_8144,N_8143);
nand U8840 (N_8840,N_8408,N_8005);
or U8841 (N_8841,N_8045,N_8087);
xnor U8842 (N_8842,N_8112,N_8330);
and U8843 (N_8843,N_8257,N_8062);
or U8844 (N_8844,N_8408,N_8469);
nor U8845 (N_8845,N_8034,N_8012);
xnor U8846 (N_8846,N_8362,N_8272);
nand U8847 (N_8847,N_8123,N_8283);
nand U8848 (N_8848,N_8128,N_8113);
or U8849 (N_8849,N_8048,N_8273);
or U8850 (N_8850,N_8212,N_8483);
or U8851 (N_8851,N_8227,N_8362);
xnor U8852 (N_8852,N_8450,N_8363);
or U8853 (N_8853,N_8290,N_8236);
and U8854 (N_8854,N_8405,N_8318);
and U8855 (N_8855,N_8077,N_8004);
nor U8856 (N_8856,N_8443,N_8177);
nor U8857 (N_8857,N_8455,N_8471);
or U8858 (N_8858,N_8103,N_8256);
nor U8859 (N_8859,N_8260,N_8137);
xnor U8860 (N_8860,N_8189,N_8305);
and U8861 (N_8861,N_8130,N_8218);
nor U8862 (N_8862,N_8043,N_8370);
nand U8863 (N_8863,N_8213,N_8327);
xnor U8864 (N_8864,N_8338,N_8155);
and U8865 (N_8865,N_8339,N_8376);
nand U8866 (N_8866,N_8096,N_8078);
xnor U8867 (N_8867,N_8483,N_8251);
and U8868 (N_8868,N_8105,N_8388);
or U8869 (N_8869,N_8325,N_8135);
or U8870 (N_8870,N_8368,N_8182);
and U8871 (N_8871,N_8207,N_8379);
nand U8872 (N_8872,N_8033,N_8199);
nand U8873 (N_8873,N_8234,N_8035);
and U8874 (N_8874,N_8222,N_8169);
nor U8875 (N_8875,N_8178,N_8188);
and U8876 (N_8876,N_8164,N_8008);
and U8877 (N_8877,N_8494,N_8435);
nand U8878 (N_8878,N_8073,N_8478);
and U8879 (N_8879,N_8270,N_8037);
nand U8880 (N_8880,N_8481,N_8374);
nor U8881 (N_8881,N_8283,N_8219);
xnor U8882 (N_8882,N_8165,N_8139);
nand U8883 (N_8883,N_8431,N_8394);
and U8884 (N_8884,N_8249,N_8277);
nand U8885 (N_8885,N_8253,N_8491);
nand U8886 (N_8886,N_8048,N_8255);
nand U8887 (N_8887,N_8011,N_8450);
xor U8888 (N_8888,N_8154,N_8306);
xor U8889 (N_8889,N_8196,N_8091);
nand U8890 (N_8890,N_8368,N_8018);
nand U8891 (N_8891,N_8127,N_8169);
xor U8892 (N_8892,N_8062,N_8440);
or U8893 (N_8893,N_8401,N_8282);
xnor U8894 (N_8894,N_8178,N_8185);
nor U8895 (N_8895,N_8290,N_8454);
nand U8896 (N_8896,N_8355,N_8356);
or U8897 (N_8897,N_8032,N_8196);
nand U8898 (N_8898,N_8067,N_8063);
xor U8899 (N_8899,N_8439,N_8203);
xnor U8900 (N_8900,N_8265,N_8104);
and U8901 (N_8901,N_8286,N_8426);
xnor U8902 (N_8902,N_8373,N_8462);
nor U8903 (N_8903,N_8090,N_8045);
nand U8904 (N_8904,N_8313,N_8090);
or U8905 (N_8905,N_8232,N_8153);
or U8906 (N_8906,N_8435,N_8132);
nand U8907 (N_8907,N_8261,N_8271);
nand U8908 (N_8908,N_8189,N_8250);
xor U8909 (N_8909,N_8154,N_8197);
nor U8910 (N_8910,N_8316,N_8275);
nor U8911 (N_8911,N_8325,N_8444);
or U8912 (N_8912,N_8022,N_8266);
xnor U8913 (N_8913,N_8275,N_8416);
and U8914 (N_8914,N_8273,N_8322);
nand U8915 (N_8915,N_8004,N_8231);
nand U8916 (N_8916,N_8277,N_8078);
nor U8917 (N_8917,N_8459,N_8143);
nor U8918 (N_8918,N_8229,N_8380);
nor U8919 (N_8919,N_8273,N_8372);
and U8920 (N_8920,N_8235,N_8312);
nor U8921 (N_8921,N_8071,N_8170);
or U8922 (N_8922,N_8385,N_8273);
nor U8923 (N_8923,N_8379,N_8236);
or U8924 (N_8924,N_8015,N_8319);
nand U8925 (N_8925,N_8083,N_8321);
nand U8926 (N_8926,N_8012,N_8234);
nor U8927 (N_8927,N_8442,N_8488);
or U8928 (N_8928,N_8435,N_8296);
and U8929 (N_8929,N_8074,N_8349);
or U8930 (N_8930,N_8124,N_8348);
nor U8931 (N_8931,N_8320,N_8043);
and U8932 (N_8932,N_8450,N_8021);
and U8933 (N_8933,N_8048,N_8434);
nor U8934 (N_8934,N_8181,N_8097);
and U8935 (N_8935,N_8313,N_8277);
xor U8936 (N_8936,N_8383,N_8036);
or U8937 (N_8937,N_8192,N_8430);
or U8938 (N_8938,N_8268,N_8476);
xnor U8939 (N_8939,N_8071,N_8053);
xor U8940 (N_8940,N_8105,N_8053);
nand U8941 (N_8941,N_8396,N_8419);
nor U8942 (N_8942,N_8349,N_8362);
xor U8943 (N_8943,N_8270,N_8295);
nor U8944 (N_8944,N_8217,N_8033);
nand U8945 (N_8945,N_8017,N_8195);
nor U8946 (N_8946,N_8268,N_8492);
xnor U8947 (N_8947,N_8435,N_8220);
and U8948 (N_8948,N_8172,N_8492);
nor U8949 (N_8949,N_8301,N_8036);
or U8950 (N_8950,N_8238,N_8212);
and U8951 (N_8951,N_8474,N_8355);
nand U8952 (N_8952,N_8467,N_8313);
and U8953 (N_8953,N_8409,N_8093);
or U8954 (N_8954,N_8443,N_8287);
or U8955 (N_8955,N_8188,N_8240);
nand U8956 (N_8956,N_8218,N_8433);
and U8957 (N_8957,N_8182,N_8102);
or U8958 (N_8958,N_8445,N_8069);
and U8959 (N_8959,N_8079,N_8162);
nand U8960 (N_8960,N_8256,N_8016);
nand U8961 (N_8961,N_8160,N_8302);
nand U8962 (N_8962,N_8141,N_8057);
nand U8963 (N_8963,N_8113,N_8443);
nand U8964 (N_8964,N_8032,N_8027);
and U8965 (N_8965,N_8433,N_8355);
nand U8966 (N_8966,N_8220,N_8294);
nor U8967 (N_8967,N_8343,N_8087);
or U8968 (N_8968,N_8171,N_8267);
nand U8969 (N_8969,N_8405,N_8246);
xnor U8970 (N_8970,N_8233,N_8271);
or U8971 (N_8971,N_8275,N_8462);
nand U8972 (N_8972,N_8023,N_8333);
nand U8973 (N_8973,N_8349,N_8250);
xnor U8974 (N_8974,N_8179,N_8299);
and U8975 (N_8975,N_8162,N_8194);
nor U8976 (N_8976,N_8187,N_8238);
xor U8977 (N_8977,N_8273,N_8159);
or U8978 (N_8978,N_8388,N_8486);
nor U8979 (N_8979,N_8305,N_8447);
or U8980 (N_8980,N_8421,N_8235);
or U8981 (N_8981,N_8014,N_8088);
xnor U8982 (N_8982,N_8470,N_8206);
or U8983 (N_8983,N_8253,N_8105);
and U8984 (N_8984,N_8135,N_8243);
and U8985 (N_8985,N_8403,N_8072);
xnor U8986 (N_8986,N_8341,N_8055);
or U8987 (N_8987,N_8179,N_8301);
nor U8988 (N_8988,N_8189,N_8202);
nor U8989 (N_8989,N_8132,N_8110);
and U8990 (N_8990,N_8184,N_8135);
and U8991 (N_8991,N_8388,N_8434);
xnor U8992 (N_8992,N_8363,N_8446);
and U8993 (N_8993,N_8132,N_8496);
or U8994 (N_8994,N_8495,N_8070);
nor U8995 (N_8995,N_8169,N_8000);
and U8996 (N_8996,N_8276,N_8237);
or U8997 (N_8997,N_8282,N_8399);
nor U8998 (N_8998,N_8013,N_8131);
nor U8999 (N_8999,N_8439,N_8226);
nand U9000 (N_9000,N_8735,N_8821);
nor U9001 (N_9001,N_8982,N_8541);
and U9002 (N_9002,N_8567,N_8525);
nand U9003 (N_9003,N_8657,N_8748);
and U9004 (N_9004,N_8823,N_8987);
nand U9005 (N_9005,N_8533,N_8863);
or U9006 (N_9006,N_8833,N_8648);
and U9007 (N_9007,N_8721,N_8711);
nand U9008 (N_9008,N_8936,N_8928);
nand U9009 (N_9009,N_8834,N_8555);
xor U9010 (N_9010,N_8803,N_8677);
or U9011 (N_9011,N_8736,N_8852);
xor U9012 (N_9012,N_8954,N_8764);
or U9013 (N_9013,N_8912,N_8841);
xor U9014 (N_9014,N_8884,N_8846);
nand U9015 (N_9015,N_8752,N_8911);
and U9016 (N_9016,N_8709,N_8767);
nand U9017 (N_9017,N_8808,N_8508);
or U9018 (N_9018,N_8603,N_8586);
nor U9019 (N_9019,N_8899,N_8717);
or U9020 (N_9020,N_8605,N_8835);
and U9021 (N_9021,N_8795,N_8630);
xnor U9022 (N_9022,N_8546,N_8923);
nand U9023 (N_9023,N_8608,N_8785);
and U9024 (N_9024,N_8639,N_8663);
nand U9025 (N_9025,N_8751,N_8642);
nand U9026 (N_9026,N_8553,N_8817);
and U9027 (N_9027,N_8990,N_8924);
or U9028 (N_9028,N_8726,N_8776);
and U9029 (N_9029,N_8755,N_8890);
nand U9030 (N_9030,N_8732,N_8964);
and U9031 (N_9031,N_8937,N_8920);
xnor U9032 (N_9032,N_8652,N_8958);
xnor U9033 (N_9033,N_8563,N_8845);
xnor U9034 (N_9034,N_8624,N_8626);
nand U9035 (N_9035,N_8504,N_8629);
nor U9036 (N_9036,N_8734,N_8668);
and U9037 (N_9037,N_8888,N_8976);
nor U9038 (N_9038,N_8713,N_8611);
or U9039 (N_9039,N_8750,N_8723);
xor U9040 (N_9040,N_8913,N_8665);
xor U9041 (N_9041,N_8649,N_8638);
or U9042 (N_9042,N_8820,N_8731);
nor U9043 (N_9043,N_8816,N_8822);
nand U9044 (N_9044,N_8951,N_8728);
or U9045 (N_9045,N_8685,N_8851);
nand U9046 (N_9046,N_8617,N_8646);
and U9047 (N_9047,N_8980,N_8962);
xor U9048 (N_9048,N_8749,N_8559);
and U9049 (N_9049,N_8840,N_8666);
or U9050 (N_9050,N_8584,N_8893);
and U9051 (N_9051,N_8931,N_8679);
or U9052 (N_9052,N_8545,N_8683);
nor U9053 (N_9053,N_8539,N_8623);
nor U9054 (N_9054,N_8975,N_8694);
and U9055 (N_9055,N_8556,N_8604);
or U9056 (N_9056,N_8988,N_8867);
nand U9057 (N_9057,N_8784,N_8826);
xor U9058 (N_9058,N_8781,N_8896);
and U9059 (N_9059,N_8871,N_8939);
nand U9060 (N_9060,N_8789,N_8837);
xnor U9061 (N_9061,N_8869,N_8947);
nor U9062 (N_9062,N_8957,N_8614);
xnor U9063 (N_9063,N_8885,N_8692);
or U9064 (N_9064,N_8682,N_8534);
and U9065 (N_9065,N_8777,N_8870);
xnor U9066 (N_9066,N_8632,N_8618);
nand U9067 (N_9067,N_8687,N_8872);
nand U9068 (N_9068,N_8577,N_8747);
and U9069 (N_9069,N_8500,N_8695);
and U9070 (N_9070,N_8842,N_8664);
and U9071 (N_9071,N_8944,N_8760);
xnor U9072 (N_9072,N_8763,N_8887);
nor U9073 (N_9073,N_8654,N_8991);
nand U9074 (N_9074,N_8971,N_8797);
and U9075 (N_9075,N_8529,N_8905);
nor U9076 (N_9076,N_8526,N_8866);
or U9077 (N_9077,N_8703,N_8774);
or U9078 (N_9078,N_8597,N_8719);
xnor U9079 (N_9079,N_8984,N_8849);
xnor U9080 (N_9080,N_8733,N_8758);
nor U9081 (N_9081,N_8836,N_8616);
nor U9082 (N_9082,N_8699,N_8875);
or U9083 (N_9083,N_8818,N_8942);
or U9084 (N_9084,N_8768,N_8513);
or U9085 (N_9085,N_8540,N_8620);
or U9086 (N_9086,N_8720,N_8933);
or U9087 (N_9087,N_8985,N_8909);
nand U9088 (N_9088,N_8537,N_8635);
and U9089 (N_9089,N_8828,N_8798);
xnor U9090 (N_9090,N_8855,N_8554);
xor U9091 (N_9091,N_8744,N_8932);
or U9092 (N_9092,N_8520,N_8598);
nand U9093 (N_9093,N_8714,N_8551);
nor U9094 (N_9094,N_8918,N_8970);
xnor U9095 (N_9095,N_8961,N_8656);
nor U9096 (N_9096,N_8974,N_8791);
and U9097 (N_9097,N_8792,N_8583);
nor U9098 (N_9098,N_8535,N_8847);
and U9099 (N_9099,N_8756,N_8641);
and U9100 (N_9100,N_8806,N_8861);
and U9101 (N_9101,N_8645,N_8673);
or U9102 (N_9102,N_8517,N_8956);
xor U9103 (N_9103,N_8590,N_8927);
xnor U9104 (N_9104,N_8519,N_8670);
and U9105 (N_9105,N_8946,N_8696);
and U9106 (N_9106,N_8515,N_8686);
and U9107 (N_9107,N_8883,N_8934);
nor U9108 (N_9108,N_8708,N_8602);
nor U9109 (N_9109,N_8702,N_8997);
or U9110 (N_9110,N_8521,N_8596);
nor U9111 (N_9111,N_8643,N_8972);
nand U9112 (N_9112,N_8707,N_8941);
xor U9113 (N_9113,N_8788,N_8585);
nand U9114 (N_9114,N_8610,N_8579);
nor U9115 (N_9115,N_8848,N_8929);
nor U9116 (N_9116,N_8651,N_8775);
nor U9117 (N_9117,N_8973,N_8790);
xnor U9118 (N_9118,N_8671,N_8940);
nor U9119 (N_9119,N_8783,N_8804);
nand U9120 (N_9120,N_8981,N_8514);
xnor U9121 (N_9121,N_8802,N_8729);
xor U9122 (N_9122,N_8876,N_8575);
or U9123 (N_9123,N_8880,N_8594);
or U9124 (N_9124,N_8674,N_8765);
or U9125 (N_9125,N_8593,N_8505);
or U9126 (N_9126,N_8977,N_8565);
nor U9127 (N_9127,N_8622,N_8903);
and U9128 (N_9128,N_8907,N_8589);
nand U9129 (N_9129,N_8576,N_8722);
or U9130 (N_9130,N_8704,N_8609);
and U9131 (N_9131,N_8945,N_8730);
nand U9132 (N_9132,N_8926,N_8968);
or U9133 (N_9133,N_8715,N_8672);
xnor U9134 (N_9134,N_8647,N_8572);
xnor U9135 (N_9135,N_8601,N_8938);
and U9136 (N_9136,N_8796,N_8669);
nand U9137 (N_9137,N_8658,N_8800);
or U9138 (N_9138,N_8915,N_8607);
nand U9139 (N_9139,N_8678,N_8766);
nor U9140 (N_9140,N_8550,N_8960);
xor U9141 (N_9141,N_8963,N_8854);
nor U9142 (N_9142,N_8782,N_8743);
xnor U9143 (N_9143,N_8627,N_8779);
or U9144 (N_9144,N_8773,N_8625);
xor U9145 (N_9145,N_8778,N_8621);
nor U9146 (N_9146,N_8689,N_8691);
nor U9147 (N_9147,N_8549,N_8561);
xor U9148 (N_9148,N_8700,N_8516);
or U9149 (N_9149,N_8547,N_8619);
or U9150 (N_9150,N_8599,N_8571);
xnor U9151 (N_9151,N_8509,N_8850);
xor U9152 (N_9152,N_8753,N_8588);
or U9153 (N_9153,N_8636,N_8983);
or U9154 (N_9154,N_8829,N_8580);
or U9155 (N_9155,N_8897,N_8564);
and U9156 (N_9156,N_8675,N_8873);
nor U9157 (N_9157,N_8655,N_8712);
nor U9158 (N_9158,N_8698,N_8681);
or U9159 (N_9159,N_8662,N_8511);
xor U9160 (N_9160,N_8538,N_8531);
or U9161 (N_9161,N_8548,N_8967);
nor U9162 (N_9162,N_8542,N_8814);
nor U9163 (N_9163,N_8952,N_8772);
nor U9164 (N_9164,N_8581,N_8543);
nor U9165 (N_9165,N_8771,N_8741);
nand U9166 (N_9166,N_8787,N_8660);
nor U9167 (N_9167,N_8891,N_8992);
nor U9168 (N_9168,N_8902,N_8557);
and U9169 (N_9169,N_8978,N_8996);
and U9170 (N_9170,N_8917,N_8562);
nor U9171 (N_9171,N_8793,N_8532);
and U9172 (N_9172,N_8864,N_8812);
xor U9173 (N_9173,N_8780,N_8914);
or U9174 (N_9174,N_8959,N_8879);
or U9175 (N_9175,N_8612,N_8653);
and U9176 (N_9176,N_8993,N_8819);
or U9177 (N_9177,N_8948,N_8799);
or U9178 (N_9178,N_8930,N_8943);
nand U9179 (N_9179,N_8587,N_8566);
or U9180 (N_9180,N_8680,N_8640);
nand U9181 (N_9181,N_8754,N_8965);
and U9182 (N_9182,N_8570,N_8886);
nor U9183 (N_9183,N_8831,N_8527);
xnor U9184 (N_9184,N_8536,N_8503);
or U9185 (N_9185,N_8856,N_8922);
nor U9186 (N_9186,N_8628,N_8953);
or U9187 (N_9187,N_8949,N_8904);
xor U9188 (N_9188,N_8659,N_8898);
or U9189 (N_9189,N_8600,N_8574);
xnor U9190 (N_9190,N_8794,N_8824);
and U9191 (N_9191,N_8844,N_8832);
and U9192 (N_9192,N_8894,N_8813);
xor U9193 (N_9193,N_8874,N_8573);
and U9194 (N_9194,N_8769,N_8710);
nor U9195 (N_9195,N_8979,N_8892);
and U9196 (N_9196,N_8815,N_8859);
nand U9197 (N_9197,N_8858,N_8615);
xnor U9198 (N_9198,N_8560,N_8999);
nand U9199 (N_9199,N_8558,N_8507);
nand U9200 (N_9200,N_8523,N_8759);
or U9201 (N_9201,N_8935,N_8634);
nor U9202 (N_9202,N_8552,N_8578);
or U9203 (N_9203,N_8809,N_8591);
nand U9204 (N_9204,N_8568,N_8510);
nor U9205 (N_9205,N_8862,N_8910);
xnor U9206 (N_9206,N_8518,N_8705);
xor U9207 (N_9207,N_8676,N_8805);
nor U9208 (N_9208,N_8801,N_8592);
nor U9209 (N_9209,N_8966,N_8746);
or U9210 (N_9210,N_8644,N_8811);
or U9211 (N_9211,N_8631,N_8637);
nor U9212 (N_9212,N_8853,N_8693);
and U9213 (N_9213,N_8969,N_8916);
xnor U9214 (N_9214,N_8725,N_8633);
nor U9215 (N_9215,N_8868,N_8528);
or U9216 (N_9216,N_8986,N_8569);
nand U9217 (N_9217,N_8522,N_8595);
or U9218 (N_9218,N_8919,N_8825);
nor U9219 (N_9219,N_8830,N_8502);
nor U9220 (N_9220,N_8718,N_8900);
nand U9221 (N_9221,N_8989,N_8762);
nand U9222 (N_9222,N_8724,N_8737);
nand U9223 (N_9223,N_8524,N_8582);
and U9224 (N_9224,N_8843,N_8667);
nor U9225 (N_9225,N_8506,N_8770);
or U9226 (N_9226,N_8757,N_8995);
xor U9227 (N_9227,N_8860,N_8877);
xnor U9228 (N_9228,N_8865,N_8606);
nand U9229 (N_9229,N_8684,N_8925);
and U9230 (N_9230,N_8661,N_8706);
nor U9231 (N_9231,N_8738,N_8613);
nor U9232 (N_9232,N_8810,N_8727);
nor U9233 (N_9233,N_8882,N_8742);
nor U9234 (N_9234,N_8761,N_8739);
and U9235 (N_9235,N_8512,N_8745);
or U9236 (N_9236,N_8650,N_8908);
and U9237 (N_9237,N_8501,N_8906);
nor U9238 (N_9238,N_8950,N_8701);
xor U9239 (N_9239,N_8955,N_8530);
nor U9240 (N_9240,N_8881,N_8889);
and U9241 (N_9241,N_8921,N_8895);
nor U9242 (N_9242,N_8827,N_8786);
nand U9243 (N_9243,N_8857,N_8998);
and U9244 (N_9244,N_8688,N_8839);
or U9245 (N_9245,N_8740,N_8838);
or U9246 (N_9246,N_8901,N_8994);
and U9247 (N_9247,N_8807,N_8544);
nand U9248 (N_9248,N_8690,N_8878);
xor U9249 (N_9249,N_8716,N_8697);
nor U9250 (N_9250,N_8739,N_8783);
nand U9251 (N_9251,N_8941,N_8737);
nand U9252 (N_9252,N_8615,N_8557);
xnor U9253 (N_9253,N_8943,N_8743);
xor U9254 (N_9254,N_8687,N_8780);
xnor U9255 (N_9255,N_8721,N_8625);
nor U9256 (N_9256,N_8598,N_8644);
xnor U9257 (N_9257,N_8858,N_8556);
or U9258 (N_9258,N_8724,N_8914);
xor U9259 (N_9259,N_8559,N_8645);
and U9260 (N_9260,N_8669,N_8973);
nor U9261 (N_9261,N_8918,N_8865);
xor U9262 (N_9262,N_8546,N_8676);
xor U9263 (N_9263,N_8823,N_8894);
nor U9264 (N_9264,N_8757,N_8556);
xnor U9265 (N_9265,N_8750,N_8678);
nand U9266 (N_9266,N_8681,N_8530);
nor U9267 (N_9267,N_8808,N_8800);
or U9268 (N_9268,N_8945,N_8524);
or U9269 (N_9269,N_8901,N_8979);
and U9270 (N_9270,N_8846,N_8527);
or U9271 (N_9271,N_8660,N_8538);
nor U9272 (N_9272,N_8646,N_8769);
nor U9273 (N_9273,N_8558,N_8749);
or U9274 (N_9274,N_8720,N_8819);
nor U9275 (N_9275,N_8815,N_8971);
or U9276 (N_9276,N_8862,N_8933);
xor U9277 (N_9277,N_8940,N_8966);
and U9278 (N_9278,N_8735,N_8723);
nand U9279 (N_9279,N_8742,N_8696);
and U9280 (N_9280,N_8763,N_8954);
xor U9281 (N_9281,N_8859,N_8735);
nand U9282 (N_9282,N_8534,N_8543);
and U9283 (N_9283,N_8836,N_8887);
xor U9284 (N_9284,N_8578,N_8874);
nor U9285 (N_9285,N_8561,N_8575);
or U9286 (N_9286,N_8971,N_8534);
or U9287 (N_9287,N_8744,N_8846);
nor U9288 (N_9288,N_8636,N_8854);
or U9289 (N_9289,N_8877,N_8585);
nand U9290 (N_9290,N_8936,N_8898);
and U9291 (N_9291,N_8794,N_8786);
and U9292 (N_9292,N_8561,N_8954);
or U9293 (N_9293,N_8609,N_8572);
nand U9294 (N_9294,N_8986,N_8718);
and U9295 (N_9295,N_8906,N_8894);
and U9296 (N_9296,N_8843,N_8933);
nor U9297 (N_9297,N_8941,N_8567);
or U9298 (N_9298,N_8986,N_8866);
nor U9299 (N_9299,N_8963,N_8699);
and U9300 (N_9300,N_8893,N_8838);
and U9301 (N_9301,N_8762,N_8675);
xor U9302 (N_9302,N_8585,N_8500);
or U9303 (N_9303,N_8654,N_8983);
or U9304 (N_9304,N_8739,N_8921);
or U9305 (N_9305,N_8991,N_8959);
nor U9306 (N_9306,N_8509,N_8627);
and U9307 (N_9307,N_8769,N_8966);
nor U9308 (N_9308,N_8560,N_8620);
and U9309 (N_9309,N_8658,N_8825);
xnor U9310 (N_9310,N_8863,N_8913);
or U9311 (N_9311,N_8669,N_8828);
nor U9312 (N_9312,N_8849,N_8928);
nand U9313 (N_9313,N_8535,N_8983);
or U9314 (N_9314,N_8940,N_8780);
nor U9315 (N_9315,N_8705,N_8829);
and U9316 (N_9316,N_8851,N_8994);
xor U9317 (N_9317,N_8515,N_8949);
nor U9318 (N_9318,N_8895,N_8973);
and U9319 (N_9319,N_8650,N_8947);
and U9320 (N_9320,N_8758,N_8897);
and U9321 (N_9321,N_8973,N_8975);
or U9322 (N_9322,N_8881,N_8894);
nand U9323 (N_9323,N_8666,N_8655);
and U9324 (N_9324,N_8646,N_8724);
or U9325 (N_9325,N_8834,N_8514);
and U9326 (N_9326,N_8676,N_8643);
nor U9327 (N_9327,N_8631,N_8684);
nand U9328 (N_9328,N_8902,N_8645);
xor U9329 (N_9329,N_8806,N_8792);
xor U9330 (N_9330,N_8699,N_8850);
and U9331 (N_9331,N_8668,N_8736);
or U9332 (N_9332,N_8741,N_8972);
nor U9333 (N_9333,N_8698,N_8752);
xor U9334 (N_9334,N_8552,N_8928);
or U9335 (N_9335,N_8678,N_8908);
or U9336 (N_9336,N_8695,N_8773);
and U9337 (N_9337,N_8852,N_8926);
nand U9338 (N_9338,N_8882,N_8951);
or U9339 (N_9339,N_8886,N_8582);
and U9340 (N_9340,N_8520,N_8955);
nand U9341 (N_9341,N_8978,N_8563);
xor U9342 (N_9342,N_8782,N_8989);
xor U9343 (N_9343,N_8845,N_8578);
nand U9344 (N_9344,N_8671,N_8758);
nor U9345 (N_9345,N_8528,N_8995);
nor U9346 (N_9346,N_8590,N_8572);
xnor U9347 (N_9347,N_8991,N_8611);
and U9348 (N_9348,N_8999,N_8973);
nand U9349 (N_9349,N_8501,N_8723);
or U9350 (N_9350,N_8757,N_8829);
and U9351 (N_9351,N_8885,N_8801);
and U9352 (N_9352,N_8620,N_8597);
and U9353 (N_9353,N_8567,N_8617);
nand U9354 (N_9354,N_8829,N_8976);
nor U9355 (N_9355,N_8624,N_8645);
nor U9356 (N_9356,N_8658,N_8746);
nor U9357 (N_9357,N_8827,N_8962);
and U9358 (N_9358,N_8985,N_8743);
or U9359 (N_9359,N_8995,N_8722);
xor U9360 (N_9360,N_8942,N_8991);
nor U9361 (N_9361,N_8608,N_8846);
or U9362 (N_9362,N_8751,N_8907);
nor U9363 (N_9363,N_8759,N_8896);
or U9364 (N_9364,N_8740,N_8803);
nor U9365 (N_9365,N_8754,N_8586);
and U9366 (N_9366,N_8986,N_8808);
nor U9367 (N_9367,N_8749,N_8960);
nand U9368 (N_9368,N_8597,N_8994);
and U9369 (N_9369,N_8718,N_8904);
xor U9370 (N_9370,N_8652,N_8830);
nand U9371 (N_9371,N_8740,N_8681);
nor U9372 (N_9372,N_8809,N_8541);
or U9373 (N_9373,N_8713,N_8850);
nand U9374 (N_9374,N_8569,N_8981);
nand U9375 (N_9375,N_8720,N_8969);
or U9376 (N_9376,N_8824,N_8731);
nor U9377 (N_9377,N_8665,N_8997);
or U9378 (N_9378,N_8837,N_8798);
or U9379 (N_9379,N_8870,N_8824);
and U9380 (N_9380,N_8943,N_8550);
xnor U9381 (N_9381,N_8508,N_8839);
xnor U9382 (N_9382,N_8589,N_8635);
nor U9383 (N_9383,N_8950,N_8680);
xor U9384 (N_9384,N_8683,N_8960);
nand U9385 (N_9385,N_8764,N_8644);
xor U9386 (N_9386,N_8593,N_8862);
or U9387 (N_9387,N_8999,N_8971);
or U9388 (N_9388,N_8651,N_8583);
nand U9389 (N_9389,N_8933,N_8665);
nor U9390 (N_9390,N_8674,N_8986);
nand U9391 (N_9391,N_8951,N_8501);
nor U9392 (N_9392,N_8864,N_8926);
or U9393 (N_9393,N_8783,N_8692);
nor U9394 (N_9394,N_8603,N_8746);
xnor U9395 (N_9395,N_8798,N_8615);
and U9396 (N_9396,N_8992,N_8544);
xnor U9397 (N_9397,N_8901,N_8880);
nor U9398 (N_9398,N_8543,N_8752);
nor U9399 (N_9399,N_8701,N_8707);
nand U9400 (N_9400,N_8561,N_8685);
nand U9401 (N_9401,N_8835,N_8625);
xor U9402 (N_9402,N_8731,N_8511);
xor U9403 (N_9403,N_8978,N_8946);
or U9404 (N_9404,N_8512,N_8782);
nand U9405 (N_9405,N_8578,N_8897);
and U9406 (N_9406,N_8525,N_8600);
nor U9407 (N_9407,N_8807,N_8707);
xor U9408 (N_9408,N_8632,N_8960);
nand U9409 (N_9409,N_8834,N_8611);
or U9410 (N_9410,N_8826,N_8708);
or U9411 (N_9411,N_8998,N_8910);
and U9412 (N_9412,N_8926,N_8823);
xor U9413 (N_9413,N_8733,N_8714);
xnor U9414 (N_9414,N_8521,N_8778);
nor U9415 (N_9415,N_8688,N_8772);
and U9416 (N_9416,N_8984,N_8669);
or U9417 (N_9417,N_8626,N_8915);
and U9418 (N_9418,N_8533,N_8773);
or U9419 (N_9419,N_8860,N_8964);
and U9420 (N_9420,N_8810,N_8504);
or U9421 (N_9421,N_8609,N_8942);
nor U9422 (N_9422,N_8702,N_8840);
or U9423 (N_9423,N_8654,N_8756);
or U9424 (N_9424,N_8910,N_8985);
or U9425 (N_9425,N_8937,N_8540);
or U9426 (N_9426,N_8663,N_8875);
or U9427 (N_9427,N_8564,N_8907);
nand U9428 (N_9428,N_8556,N_8674);
or U9429 (N_9429,N_8567,N_8738);
nor U9430 (N_9430,N_8771,N_8876);
nor U9431 (N_9431,N_8861,N_8520);
or U9432 (N_9432,N_8716,N_8612);
or U9433 (N_9433,N_8977,N_8634);
nand U9434 (N_9434,N_8949,N_8676);
nor U9435 (N_9435,N_8864,N_8668);
nor U9436 (N_9436,N_8524,N_8807);
xnor U9437 (N_9437,N_8710,N_8725);
nor U9438 (N_9438,N_8599,N_8533);
or U9439 (N_9439,N_8966,N_8533);
and U9440 (N_9440,N_8932,N_8743);
and U9441 (N_9441,N_8530,N_8520);
or U9442 (N_9442,N_8521,N_8990);
xnor U9443 (N_9443,N_8877,N_8548);
xor U9444 (N_9444,N_8545,N_8770);
and U9445 (N_9445,N_8917,N_8835);
nand U9446 (N_9446,N_8905,N_8538);
and U9447 (N_9447,N_8820,N_8781);
nor U9448 (N_9448,N_8939,N_8802);
xnor U9449 (N_9449,N_8948,N_8998);
nor U9450 (N_9450,N_8956,N_8687);
nand U9451 (N_9451,N_8599,N_8931);
or U9452 (N_9452,N_8582,N_8746);
xor U9453 (N_9453,N_8807,N_8964);
or U9454 (N_9454,N_8715,N_8957);
or U9455 (N_9455,N_8582,N_8953);
nor U9456 (N_9456,N_8658,N_8850);
nor U9457 (N_9457,N_8610,N_8547);
xnor U9458 (N_9458,N_8967,N_8545);
nor U9459 (N_9459,N_8602,N_8532);
nor U9460 (N_9460,N_8575,N_8814);
or U9461 (N_9461,N_8531,N_8519);
and U9462 (N_9462,N_8948,N_8522);
or U9463 (N_9463,N_8760,N_8508);
nor U9464 (N_9464,N_8893,N_8779);
xnor U9465 (N_9465,N_8904,N_8658);
nor U9466 (N_9466,N_8648,N_8878);
or U9467 (N_9467,N_8654,N_8701);
nor U9468 (N_9468,N_8704,N_8693);
nand U9469 (N_9469,N_8896,N_8782);
xnor U9470 (N_9470,N_8915,N_8506);
nor U9471 (N_9471,N_8855,N_8529);
or U9472 (N_9472,N_8975,N_8788);
nand U9473 (N_9473,N_8656,N_8730);
nand U9474 (N_9474,N_8647,N_8921);
or U9475 (N_9475,N_8738,N_8621);
xnor U9476 (N_9476,N_8867,N_8915);
and U9477 (N_9477,N_8922,N_8699);
and U9478 (N_9478,N_8858,N_8943);
nor U9479 (N_9479,N_8776,N_8591);
nor U9480 (N_9480,N_8826,N_8866);
nand U9481 (N_9481,N_8892,N_8784);
xnor U9482 (N_9482,N_8791,N_8886);
and U9483 (N_9483,N_8709,N_8568);
nand U9484 (N_9484,N_8593,N_8627);
and U9485 (N_9485,N_8943,N_8985);
and U9486 (N_9486,N_8906,N_8677);
nor U9487 (N_9487,N_8835,N_8694);
nor U9488 (N_9488,N_8990,N_8928);
nor U9489 (N_9489,N_8660,N_8798);
and U9490 (N_9490,N_8519,N_8619);
or U9491 (N_9491,N_8668,N_8837);
nor U9492 (N_9492,N_8631,N_8748);
and U9493 (N_9493,N_8724,N_8592);
and U9494 (N_9494,N_8941,N_8854);
nor U9495 (N_9495,N_8845,N_8727);
or U9496 (N_9496,N_8862,N_8690);
xnor U9497 (N_9497,N_8892,N_8522);
nand U9498 (N_9498,N_8637,N_8904);
nor U9499 (N_9499,N_8661,N_8845);
or U9500 (N_9500,N_9201,N_9483);
xor U9501 (N_9501,N_9077,N_9435);
nand U9502 (N_9502,N_9264,N_9219);
or U9503 (N_9503,N_9069,N_9099);
xor U9504 (N_9504,N_9260,N_9210);
or U9505 (N_9505,N_9112,N_9018);
and U9506 (N_9506,N_9228,N_9062);
and U9507 (N_9507,N_9408,N_9379);
xnor U9508 (N_9508,N_9440,N_9334);
nor U9509 (N_9509,N_9104,N_9293);
and U9510 (N_9510,N_9054,N_9469);
and U9511 (N_9511,N_9124,N_9158);
or U9512 (N_9512,N_9447,N_9399);
nor U9513 (N_9513,N_9006,N_9360);
and U9514 (N_9514,N_9449,N_9261);
and U9515 (N_9515,N_9345,N_9118);
nand U9516 (N_9516,N_9419,N_9056);
nor U9517 (N_9517,N_9336,N_9157);
and U9518 (N_9518,N_9381,N_9120);
and U9519 (N_9519,N_9254,N_9107);
nand U9520 (N_9520,N_9059,N_9078);
nand U9521 (N_9521,N_9032,N_9089);
nand U9522 (N_9522,N_9313,N_9259);
xnor U9523 (N_9523,N_9328,N_9213);
and U9524 (N_9524,N_9008,N_9288);
or U9525 (N_9525,N_9130,N_9320);
and U9526 (N_9526,N_9347,N_9387);
nand U9527 (N_9527,N_9177,N_9188);
xnor U9528 (N_9528,N_9473,N_9364);
and U9529 (N_9529,N_9131,N_9146);
xor U9530 (N_9530,N_9216,N_9214);
nor U9531 (N_9531,N_9138,N_9487);
or U9532 (N_9532,N_9178,N_9255);
nand U9533 (N_9533,N_9115,N_9133);
xor U9534 (N_9534,N_9372,N_9303);
or U9535 (N_9535,N_9171,N_9241);
nor U9536 (N_9536,N_9195,N_9411);
nand U9537 (N_9537,N_9226,N_9102);
xnor U9538 (N_9538,N_9472,N_9035);
nor U9539 (N_9539,N_9489,N_9395);
nand U9540 (N_9540,N_9355,N_9160);
nand U9541 (N_9541,N_9438,N_9442);
nand U9542 (N_9542,N_9304,N_9374);
nand U9543 (N_9543,N_9194,N_9244);
and U9544 (N_9544,N_9174,N_9396);
and U9545 (N_9545,N_9012,N_9481);
or U9546 (N_9546,N_9439,N_9256);
xnor U9547 (N_9547,N_9050,N_9116);
xnor U9548 (N_9548,N_9092,N_9308);
or U9549 (N_9549,N_9448,N_9266);
nor U9550 (N_9550,N_9240,N_9108);
nor U9551 (N_9551,N_9272,N_9033);
nor U9552 (N_9552,N_9477,N_9187);
nor U9553 (N_9553,N_9010,N_9239);
nor U9554 (N_9554,N_9060,N_9159);
and U9555 (N_9555,N_9103,N_9011);
or U9556 (N_9556,N_9096,N_9427);
nand U9557 (N_9557,N_9114,N_9192);
nor U9558 (N_9558,N_9446,N_9383);
and U9559 (N_9559,N_9267,N_9052);
xnor U9560 (N_9560,N_9172,N_9076);
nand U9561 (N_9561,N_9058,N_9329);
nand U9562 (N_9562,N_9352,N_9007);
nor U9563 (N_9563,N_9470,N_9257);
nand U9564 (N_9564,N_9414,N_9202);
nand U9565 (N_9565,N_9176,N_9068);
nor U9566 (N_9566,N_9363,N_9391);
nor U9567 (N_9567,N_9309,N_9167);
nand U9568 (N_9568,N_9406,N_9211);
or U9569 (N_9569,N_9085,N_9140);
nand U9570 (N_9570,N_9464,N_9183);
nand U9571 (N_9571,N_9258,N_9066);
nand U9572 (N_9572,N_9377,N_9038);
or U9573 (N_9573,N_9215,N_9495);
nor U9574 (N_9574,N_9073,N_9080);
nor U9575 (N_9575,N_9350,N_9340);
or U9576 (N_9576,N_9390,N_9436);
nor U9577 (N_9577,N_9394,N_9321);
and U9578 (N_9578,N_9361,N_9476);
nor U9579 (N_9579,N_9220,N_9450);
nor U9580 (N_9580,N_9110,N_9325);
xnor U9581 (N_9581,N_9422,N_9365);
nor U9582 (N_9582,N_9437,N_9029);
xnor U9583 (N_9583,N_9232,N_9225);
xor U9584 (N_9584,N_9065,N_9229);
or U9585 (N_9585,N_9298,N_9161);
or U9586 (N_9586,N_9386,N_9282);
nand U9587 (N_9587,N_9388,N_9333);
nor U9588 (N_9588,N_9248,N_9492);
nor U9589 (N_9589,N_9416,N_9203);
and U9590 (N_9590,N_9460,N_9004);
nor U9591 (N_9591,N_9407,N_9462);
nor U9592 (N_9592,N_9312,N_9016);
and U9593 (N_9593,N_9091,N_9231);
nor U9594 (N_9594,N_9278,N_9074);
or U9595 (N_9595,N_9478,N_9471);
nor U9596 (N_9596,N_9441,N_9430);
xnor U9597 (N_9597,N_9322,N_9262);
xor U9598 (N_9598,N_9067,N_9283);
xnor U9599 (N_9599,N_9064,N_9398);
nand U9600 (N_9600,N_9063,N_9370);
nor U9601 (N_9601,N_9046,N_9237);
xnor U9602 (N_9602,N_9344,N_9009);
xor U9603 (N_9603,N_9300,N_9358);
xnor U9604 (N_9604,N_9141,N_9467);
nor U9605 (N_9605,N_9337,N_9209);
or U9606 (N_9606,N_9097,N_9418);
or U9607 (N_9607,N_9238,N_9125);
nand U9608 (N_9608,N_9119,N_9389);
and U9609 (N_9609,N_9031,N_9431);
nand U9610 (N_9610,N_9181,N_9482);
xnor U9611 (N_9611,N_9385,N_9380);
or U9612 (N_9612,N_9421,N_9001);
and U9613 (N_9613,N_9015,N_9319);
nand U9614 (N_9614,N_9221,N_9276);
nor U9615 (N_9615,N_9315,N_9135);
nor U9616 (N_9616,N_9393,N_9299);
or U9617 (N_9617,N_9189,N_9485);
xnor U9618 (N_9618,N_9081,N_9417);
nand U9619 (N_9619,N_9454,N_9468);
and U9620 (N_9620,N_9456,N_9122);
nand U9621 (N_9621,N_9185,N_9093);
or U9622 (N_9622,N_9230,N_9233);
xnor U9623 (N_9623,N_9371,N_9024);
xnor U9624 (N_9624,N_9036,N_9098);
nor U9625 (N_9625,N_9072,N_9269);
nor U9626 (N_9626,N_9297,N_9271);
or U9627 (N_9627,N_9453,N_9455);
and U9628 (N_9628,N_9287,N_9316);
xnor U9629 (N_9629,N_9323,N_9292);
nand U9630 (N_9630,N_9376,N_9474);
xor U9631 (N_9631,N_9326,N_9433);
nor U9632 (N_9632,N_9279,N_9499);
and U9633 (N_9633,N_9252,N_9351);
nor U9634 (N_9634,N_9368,N_9429);
and U9635 (N_9635,N_9047,N_9494);
nand U9636 (N_9636,N_9070,N_9184);
xnor U9637 (N_9637,N_9402,N_9019);
nor U9638 (N_9638,N_9030,N_9397);
nand U9639 (N_9639,N_9335,N_9444);
xnor U9640 (N_9640,N_9034,N_9339);
and U9641 (N_9641,N_9137,N_9204);
and U9642 (N_9642,N_9366,N_9318);
xor U9643 (N_9643,N_9162,N_9490);
nand U9644 (N_9644,N_9224,N_9020);
nor U9645 (N_9645,N_9222,N_9082);
nand U9646 (N_9646,N_9413,N_9153);
and U9647 (N_9647,N_9002,N_9212);
xnor U9648 (N_9648,N_9061,N_9409);
and U9649 (N_9649,N_9169,N_9243);
nand U9650 (N_9650,N_9342,N_9205);
nand U9651 (N_9651,N_9049,N_9246);
nor U9652 (N_9652,N_9445,N_9486);
xnor U9653 (N_9653,N_9301,N_9281);
or U9654 (N_9654,N_9095,N_9236);
xor U9655 (N_9655,N_9180,N_9179);
or U9656 (N_9656,N_9041,N_9479);
nand U9657 (N_9657,N_9317,N_9042);
or U9658 (N_9658,N_9491,N_9055);
nand U9659 (N_9659,N_9463,N_9121);
xnor U9660 (N_9660,N_9139,N_9128);
nand U9661 (N_9661,N_9410,N_9142);
xor U9662 (N_9662,N_9190,N_9245);
and U9663 (N_9663,N_9362,N_9294);
or U9664 (N_9664,N_9498,N_9331);
nor U9665 (N_9665,N_9400,N_9143);
xnor U9666 (N_9666,N_9459,N_9028);
xor U9667 (N_9667,N_9079,N_9405);
or U9668 (N_9668,N_9296,N_9191);
nor U9669 (N_9669,N_9466,N_9057);
and U9670 (N_9670,N_9127,N_9275);
nand U9671 (N_9671,N_9136,N_9017);
xnor U9672 (N_9672,N_9148,N_9330);
nor U9673 (N_9673,N_9426,N_9310);
nor U9674 (N_9674,N_9346,N_9175);
or U9675 (N_9675,N_9193,N_9458);
nor U9676 (N_9676,N_9314,N_9132);
and U9677 (N_9677,N_9113,N_9109);
nor U9678 (N_9678,N_9307,N_9145);
and U9679 (N_9679,N_9434,N_9013);
xor U9680 (N_9680,N_9053,N_9000);
nor U9681 (N_9681,N_9265,N_9165);
nand U9682 (N_9682,N_9327,N_9186);
and U9683 (N_9683,N_9338,N_9401);
xnor U9684 (N_9684,N_9359,N_9423);
and U9685 (N_9685,N_9425,N_9349);
nor U9686 (N_9686,N_9324,N_9424);
nand U9687 (N_9687,N_9234,N_9270);
nor U9688 (N_9688,N_9451,N_9100);
xor U9689 (N_9689,N_9311,N_9249);
nor U9690 (N_9690,N_9086,N_9199);
and U9691 (N_9691,N_9123,N_9173);
or U9692 (N_9692,N_9022,N_9384);
and U9693 (N_9693,N_9218,N_9206);
nor U9694 (N_9694,N_9382,N_9353);
nor U9695 (N_9695,N_9200,N_9014);
xor U9696 (N_9696,N_9025,N_9026);
or U9697 (N_9697,N_9134,N_9037);
nor U9698 (N_9698,N_9378,N_9090);
and U9699 (N_9699,N_9182,N_9284);
and U9700 (N_9700,N_9147,N_9392);
and U9701 (N_9701,N_9274,N_9465);
or U9702 (N_9702,N_9126,N_9354);
xnor U9703 (N_9703,N_9291,N_9223);
nand U9704 (N_9704,N_9152,N_9150);
xnor U9705 (N_9705,N_9404,N_9088);
and U9706 (N_9706,N_9443,N_9428);
or U9707 (N_9707,N_9268,N_9277);
and U9708 (N_9708,N_9156,N_9087);
xor U9709 (N_9709,N_9197,N_9170);
nor U9710 (N_9710,N_9290,N_9003);
nor U9711 (N_9711,N_9247,N_9154);
and U9712 (N_9712,N_9045,N_9235);
or U9713 (N_9713,N_9075,N_9302);
and U9714 (N_9714,N_9196,N_9273);
or U9715 (N_9715,N_9420,N_9043);
nor U9716 (N_9716,N_9111,N_9005);
and U9717 (N_9717,N_9250,N_9051);
nand U9718 (N_9718,N_9280,N_9217);
or U9719 (N_9719,N_9488,N_9144);
and U9720 (N_9720,N_9198,N_9168);
or U9721 (N_9721,N_9285,N_9305);
or U9722 (N_9722,N_9457,N_9023);
and U9723 (N_9723,N_9117,N_9475);
xnor U9724 (N_9724,N_9105,N_9412);
xnor U9725 (N_9725,N_9163,N_9348);
xnor U9726 (N_9726,N_9129,N_9403);
and U9727 (N_9727,N_9306,N_9207);
and U9728 (N_9728,N_9289,N_9164);
nor U9729 (N_9729,N_9094,N_9242);
and U9730 (N_9730,N_9367,N_9027);
nand U9731 (N_9731,N_9452,N_9432);
xnor U9732 (N_9732,N_9071,N_9048);
xor U9733 (N_9733,N_9040,N_9496);
xnor U9734 (N_9734,N_9263,N_9039);
and U9735 (N_9735,N_9083,N_9493);
xor U9736 (N_9736,N_9343,N_9375);
xnor U9737 (N_9737,N_9149,N_9356);
xor U9738 (N_9738,N_9021,N_9166);
nand U9739 (N_9739,N_9155,N_9227);
nor U9740 (N_9740,N_9208,N_9253);
and U9741 (N_9741,N_9084,N_9295);
nand U9742 (N_9742,N_9341,N_9461);
or U9743 (N_9743,N_9251,N_9151);
xor U9744 (N_9744,N_9357,N_9480);
nand U9745 (N_9745,N_9369,N_9415);
and U9746 (N_9746,N_9044,N_9497);
and U9747 (N_9747,N_9286,N_9484);
xnor U9748 (N_9748,N_9373,N_9106);
nand U9749 (N_9749,N_9332,N_9101);
nand U9750 (N_9750,N_9247,N_9177);
or U9751 (N_9751,N_9306,N_9454);
xor U9752 (N_9752,N_9392,N_9290);
and U9753 (N_9753,N_9286,N_9478);
or U9754 (N_9754,N_9488,N_9160);
xor U9755 (N_9755,N_9326,N_9029);
xnor U9756 (N_9756,N_9038,N_9147);
xnor U9757 (N_9757,N_9205,N_9490);
xnor U9758 (N_9758,N_9458,N_9113);
and U9759 (N_9759,N_9027,N_9312);
nor U9760 (N_9760,N_9232,N_9107);
nor U9761 (N_9761,N_9337,N_9006);
nand U9762 (N_9762,N_9184,N_9040);
nand U9763 (N_9763,N_9428,N_9241);
or U9764 (N_9764,N_9241,N_9453);
xor U9765 (N_9765,N_9098,N_9032);
nor U9766 (N_9766,N_9462,N_9298);
or U9767 (N_9767,N_9148,N_9240);
nand U9768 (N_9768,N_9263,N_9169);
and U9769 (N_9769,N_9047,N_9307);
or U9770 (N_9770,N_9408,N_9221);
xor U9771 (N_9771,N_9379,N_9127);
nand U9772 (N_9772,N_9040,N_9109);
xnor U9773 (N_9773,N_9437,N_9313);
nor U9774 (N_9774,N_9102,N_9114);
or U9775 (N_9775,N_9066,N_9366);
or U9776 (N_9776,N_9221,N_9349);
xor U9777 (N_9777,N_9166,N_9443);
and U9778 (N_9778,N_9337,N_9297);
nor U9779 (N_9779,N_9173,N_9135);
nand U9780 (N_9780,N_9422,N_9212);
and U9781 (N_9781,N_9253,N_9486);
and U9782 (N_9782,N_9276,N_9012);
xnor U9783 (N_9783,N_9061,N_9379);
or U9784 (N_9784,N_9238,N_9171);
or U9785 (N_9785,N_9046,N_9011);
or U9786 (N_9786,N_9202,N_9443);
and U9787 (N_9787,N_9254,N_9423);
nor U9788 (N_9788,N_9365,N_9426);
xnor U9789 (N_9789,N_9352,N_9054);
and U9790 (N_9790,N_9065,N_9143);
or U9791 (N_9791,N_9152,N_9403);
and U9792 (N_9792,N_9364,N_9261);
nor U9793 (N_9793,N_9293,N_9199);
nand U9794 (N_9794,N_9345,N_9459);
and U9795 (N_9795,N_9272,N_9021);
nor U9796 (N_9796,N_9344,N_9383);
xnor U9797 (N_9797,N_9384,N_9110);
xnor U9798 (N_9798,N_9303,N_9038);
nand U9799 (N_9799,N_9459,N_9244);
xor U9800 (N_9800,N_9032,N_9255);
nand U9801 (N_9801,N_9250,N_9472);
nand U9802 (N_9802,N_9323,N_9386);
nor U9803 (N_9803,N_9160,N_9153);
xnor U9804 (N_9804,N_9444,N_9375);
and U9805 (N_9805,N_9080,N_9293);
nand U9806 (N_9806,N_9137,N_9478);
nand U9807 (N_9807,N_9409,N_9075);
xor U9808 (N_9808,N_9066,N_9306);
xor U9809 (N_9809,N_9326,N_9397);
xor U9810 (N_9810,N_9305,N_9256);
nor U9811 (N_9811,N_9247,N_9230);
xnor U9812 (N_9812,N_9037,N_9336);
nor U9813 (N_9813,N_9259,N_9484);
nor U9814 (N_9814,N_9262,N_9177);
nor U9815 (N_9815,N_9447,N_9402);
xnor U9816 (N_9816,N_9029,N_9389);
xnor U9817 (N_9817,N_9093,N_9100);
nand U9818 (N_9818,N_9027,N_9445);
and U9819 (N_9819,N_9343,N_9245);
and U9820 (N_9820,N_9256,N_9028);
nand U9821 (N_9821,N_9402,N_9221);
xor U9822 (N_9822,N_9388,N_9103);
and U9823 (N_9823,N_9240,N_9294);
or U9824 (N_9824,N_9024,N_9133);
xnor U9825 (N_9825,N_9211,N_9307);
nor U9826 (N_9826,N_9276,N_9327);
or U9827 (N_9827,N_9079,N_9212);
nand U9828 (N_9828,N_9134,N_9151);
or U9829 (N_9829,N_9294,N_9142);
nand U9830 (N_9830,N_9219,N_9086);
or U9831 (N_9831,N_9408,N_9295);
xnor U9832 (N_9832,N_9239,N_9234);
nor U9833 (N_9833,N_9481,N_9333);
and U9834 (N_9834,N_9147,N_9240);
nand U9835 (N_9835,N_9034,N_9482);
nor U9836 (N_9836,N_9453,N_9333);
xor U9837 (N_9837,N_9496,N_9376);
or U9838 (N_9838,N_9297,N_9287);
nand U9839 (N_9839,N_9066,N_9196);
xnor U9840 (N_9840,N_9309,N_9472);
nand U9841 (N_9841,N_9223,N_9146);
nor U9842 (N_9842,N_9307,N_9209);
nor U9843 (N_9843,N_9085,N_9126);
or U9844 (N_9844,N_9209,N_9437);
nand U9845 (N_9845,N_9092,N_9126);
xnor U9846 (N_9846,N_9175,N_9043);
and U9847 (N_9847,N_9439,N_9113);
or U9848 (N_9848,N_9103,N_9325);
or U9849 (N_9849,N_9198,N_9480);
or U9850 (N_9850,N_9341,N_9087);
and U9851 (N_9851,N_9026,N_9323);
xnor U9852 (N_9852,N_9235,N_9081);
and U9853 (N_9853,N_9341,N_9437);
nor U9854 (N_9854,N_9433,N_9140);
nor U9855 (N_9855,N_9352,N_9408);
and U9856 (N_9856,N_9449,N_9131);
or U9857 (N_9857,N_9227,N_9450);
nor U9858 (N_9858,N_9106,N_9377);
or U9859 (N_9859,N_9343,N_9331);
nor U9860 (N_9860,N_9377,N_9086);
nor U9861 (N_9861,N_9113,N_9081);
nor U9862 (N_9862,N_9034,N_9054);
nand U9863 (N_9863,N_9467,N_9478);
or U9864 (N_9864,N_9450,N_9308);
and U9865 (N_9865,N_9123,N_9040);
and U9866 (N_9866,N_9443,N_9213);
or U9867 (N_9867,N_9293,N_9141);
nand U9868 (N_9868,N_9337,N_9211);
xor U9869 (N_9869,N_9312,N_9222);
nor U9870 (N_9870,N_9323,N_9231);
nor U9871 (N_9871,N_9313,N_9469);
nor U9872 (N_9872,N_9153,N_9426);
or U9873 (N_9873,N_9279,N_9395);
nand U9874 (N_9874,N_9321,N_9059);
nor U9875 (N_9875,N_9253,N_9037);
nor U9876 (N_9876,N_9172,N_9479);
nand U9877 (N_9877,N_9002,N_9204);
or U9878 (N_9878,N_9278,N_9265);
and U9879 (N_9879,N_9012,N_9269);
and U9880 (N_9880,N_9256,N_9218);
or U9881 (N_9881,N_9403,N_9006);
xor U9882 (N_9882,N_9117,N_9018);
nor U9883 (N_9883,N_9292,N_9306);
and U9884 (N_9884,N_9420,N_9496);
xnor U9885 (N_9885,N_9264,N_9336);
and U9886 (N_9886,N_9141,N_9251);
and U9887 (N_9887,N_9363,N_9382);
or U9888 (N_9888,N_9375,N_9486);
xor U9889 (N_9889,N_9185,N_9005);
and U9890 (N_9890,N_9004,N_9351);
nand U9891 (N_9891,N_9171,N_9026);
nor U9892 (N_9892,N_9207,N_9019);
nand U9893 (N_9893,N_9399,N_9277);
or U9894 (N_9894,N_9455,N_9407);
nand U9895 (N_9895,N_9149,N_9233);
and U9896 (N_9896,N_9233,N_9277);
or U9897 (N_9897,N_9091,N_9312);
or U9898 (N_9898,N_9140,N_9166);
and U9899 (N_9899,N_9438,N_9113);
nor U9900 (N_9900,N_9215,N_9211);
xor U9901 (N_9901,N_9498,N_9257);
xor U9902 (N_9902,N_9195,N_9187);
or U9903 (N_9903,N_9428,N_9267);
nand U9904 (N_9904,N_9007,N_9130);
xnor U9905 (N_9905,N_9367,N_9369);
nand U9906 (N_9906,N_9160,N_9016);
xnor U9907 (N_9907,N_9310,N_9342);
nand U9908 (N_9908,N_9266,N_9180);
xnor U9909 (N_9909,N_9305,N_9408);
or U9910 (N_9910,N_9387,N_9190);
nor U9911 (N_9911,N_9400,N_9001);
nand U9912 (N_9912,N_9048,N_9042);
nand U9913 (N_9913,N_9121,N_9002);
nor U9914 (N_9914,N_9356,N_9183);
nor U9915 (N_9915,N_9309,N_9222);
xnor U9916 (N_9916,N_9380,N_9193);
nor U9917 (N_9917,N_9120,N_9020);
and U9918 (N_9918,N_9196,N_9301);
nand U9919 (N_9919,N_9226,N_9120);
xor U9920 (N_9920,N_9396,N_9034);
nor U9921 (N_9921,N_9176,N_9334);
nor U9922 (N_9922,N_9263,N_9449);
xor U9923 (N_9923,N_9401,N_9288);
and U9924 (N_9924,N_9003,N_9129);
xnor U9925 (N_9925,N_9462,N_9035);
or U9926 (N_9926,N_9277,N_9148);
nor U9927 (N_9927,N_9086,N_9130);
nand U9928 (N_9928,N_9480,N_9151);
xnor U9929 (N_9929,N_9299,N_9359);
and U9930 (N_9930,N_9091,N_9056);
xnor U9931 (N_9931,N_9421,N_9024);
nand U9932 (N_9932,N_9091,N_9398);
nor U9933 (N_9933,N_9414,N_9072);
or U9934 (N_9934,N_9070,N_9232);
nand U9935 (N_9935,N_9016,N_9470);
and U9936 (N_9936,N_9347,N_9164);
xor U9937 (N_9937,N_9082,N_9385);
nor U9938 (N_9938,N_9383,N_9393);
or U9939 (N_9939,N_9189,N_9234);
nor U9940 (N_9940,N_9422,N_9460);
or U9941 (N_9941,N_9446,N_9352);
xor U9942 (N_9942,N_9425,N_9257);
nor U9943 (N_9943,N_9005,N_9221);
nand U9944 (N_9944,N_9434,N_9324);
and U9945 (N_9945,N_9214,N_9401);
and U9946 (N_9946,N_9196,N_9267);
or U9947 (N_9947,N_9233,N_9418);
nor U9948 (N_9948,N_9496,N_9107);
xor U9949 (N_9949,N_9417,N_9454);
xnor U9950 (N_9950,N_9172,N_9473);
or U9951 (N_9951,N_9307,N_9291);
nor U9952 (N_9952,N_9263,N_9353);
nand U9953 (N_9953,N_9380,N_9130);
nand U9954 (N_9954,N_9067,N_9280);
xnor U9955 (N_9955,N_9253,N_9105);
or U9956 (N_9956,N_9113,N_9067);
or U9957 (N_9957,N_9390,N_9465);
nand U9958 (N_9958,N_9253,N_9475);
nor U9959 (N_9959,N_9380,N_9164);
and U9960 (N_9960,N_9014,N_9078);
nor U9961 (N_9961,N_9426,N_9127);
nand U9962 (N_9962,N_9493,N_9458);
nor U9963 (N_9963,N_9306,N_9159);
nand U9964 (N_9964,N_9100,N_9282);
xor U9965 (N_9965,N_9085,N_9115);
nor U9966 (N_9966,N_9323,N_9445);
nand U9967 (N_9967,N_9379,N_9135);
nor U9968 (N_9968,N_9190,N_9340);
and U9969 (N_9969,N_9285,N_9425);
nand U9970 (N_9970,N_9135,N_9149);
nand U9971 (N_9971,N_9385,N_9097);
xnor U9972 (N_9972,N_9062,N_9160);
nor U9973 (N_9973,N_9354,N_9317);
and U9974 (N_9974,N_9090,N_9350);
and U9975 (N_9975,N_9098,N_9105);
and U9976 (N_9976,N_9422,N_9057);
nand U9977 (N_9977,N_9235,N_9458);
nor U9978 (N_9978,N_9041,N_9177);
nand U9979 (N_9979,N_9421,N_9451);
or U9980 (N_9980,N_9086,N_9021);
nand U9981 (N_9981,N_9099,N_9252);
and U9982 (N_9982,N_9311,N_9066);
or U9983 (N_9983,N_9397,N_9034);
and U9984 (N_9984,N_9312,N_9416);
xnor U9985 (N_9985,N_9392,N_9060);
or U9986 (N_9986,N_9286,N_9404);
xnor U9987 (N_9987,N_9223,N_9367);
or U9988 (N_9988,N_9134,N_9272);
or U9989 (N_9989,N_9137,N_9425);
nor U9990 (N_9990,N_9080,N_9432);
nand U9991 (N_9991,N_9157,N_9122);
xnor U9992 (N_9992,N_9081,N_9013);
and U9993 (N_9993,N_9159,N_9449);
nand U9994 (N_9994,N_9175,N_9008);
nor U9995 (N_9995,N_9331,N_9081);
or U9996 (N_9996,N_9480,N_9015);
nor U9997 (N_9997,N_9250,N_9323);
or U9998 (N_9998,N_9024,N_9013);
xnor U9999 (N_9999,N_9274,N_9171);
or U10000 (N_10000,N_9539,N_9953);
or U10001 (N_10001,N_9889,N_9507);
nand U10002 (N_10002,N_9613,N_9956);
and U10003 (N_10003,N_9860,N_9564);
xnor U10004 (N_10004,N_9972,N_9810);
or U10005 (N_10005,N_9572,N_9812);
and U10006 (N_10006,N_9913,N_9798);
or U10007 (N_10007,N_9585,N_9894);
nor U10008 (N_10008,N_9664,N_9838);
nor U10009 (N_10009,N_9587,N_9588);
nor U10010 (N_10010,N_9684,N_9771);
nand U10011 (N_10011,N_9918,N_9908);
xnor U10012 (N_10012,N_9911,N_9517);
nand U10013 (N_10013,N_9523,N_9778);
and U10014 (N_10014,N_9891,N_9690);
nand U10015 (N_10015,N_9931,N_9824);
and U10016 (N_10016,N_9786,N_9694);
and U10017 (N_10017,N_9792,N_9733);
and U10018 (N_10018,N_9688,N_9712);
xnor U10019 (N_10019,N_9628,N_9974);
and U10020 (N_10020,N_9837,N_9502);
nand U10021 (N_10021,N_9979,N_9852);
or U10022 (N_10022,N_9759,N_9963);
nand U10023 (N_10023,N_9981,N_9900);
nor U10024 (N_10024,N_9506,N_9598);
and U10025 (N_10025,N_9532,N_9867);
nor U10026 (N_10026,N_9619,N_9925);
xnor U10027 (N_10027,N_9691,N_9817);
nor U10028 (N_10028,N_9647,N_9504);
nand U10029 (N_10029,N_9937,N_9580);
and U10030 (N_10030,N_9832,N_9750);
or U10031 (N_10031,N_9795,N_9967);
xnor U10032 (N_10032,N_9714,N_9801);
and U10033 (N_10033,N_9873,N_9534);
and U10034 (N_10034,N_9753,N_9548);
nor U10035 (N_10035,N_9849,N_9743);
nor U10036 (N_10036,N_9893,N_9758);
nand U10037 (N_10037,N_9610,N_9631);
nor U10038 (N_10038,N_9609,N_9643);
nand U10039 (N_10039,N_9607,N_9769);
xnor U10040 (N_10040,N_9790,N_9606);
nor U10041 (N_10041,N_9624,N_9671);
xnor U10042 (N_10042,N_9980,N_9739);
nor U10043 (N_10043,N_9802,N_9885);
or U10044 (N_10044,N_9579,N_9922);
nor U10045 (N_10045,N_9681,N_9819);
nor U10046 (N_10046,N_9546,N_9676);
nor U10047 (N_10047,N_9661,N_9708);
nor U10048 (N_10048,N_9562,N_9730);
or U10049 (N_10049,N_9905,N_9724);
nor U10050 (N_10050,N_9531,N_9594);
nand U10051 (N_10051,N_9719,N_9711);
nor U10052 (N_10052,N_9800,N_9655);
or U10053 (N_10053,N_9616,N_9907);
nand U10054 (N_10054,N_9674,N_9685);
or U10055 (N_10055,N_9505,N_9958);
and U10056 (N_10056,N_9544,N_9738);
nand U10057 (N_10057,N_9912,N_9768);
or U10058 (N_10058,N_9603,N_9622);
xor U10059 (N_10059,N_9592,N_9704);
nor U10060 (N_10060,N_9649,N_9949);
xnor U10061 (N_10061,N_9946,N_9951);
nand U10062 (N_10062,N_9635,N_9914);
and U10063 (N_10063,N_9565,N_9945);
or U10064 (N_10064,N_9927,N_9668);
nand U10065 (N_10065,N_9767,N_9672);
xnor U10066 (N_10066,N_9799,N_9542);
xnor U10067 (N_10067,N_9586,N_9856);
xnor U10068 (N_10068,N_9764,N_9716);
or U10069 (N_10069,N_9899,N_9825);
nor U10070 (N_10070,N_9600,N_9796);
or U10071 (N_10071,N_9556,N_9513);
and U10072 (N_10072,N_9783,N_9844);
nor U10073 (N_10073,N_9842,N_9848);
and U10074 (N_10074,N_9508,N_9954);
or U10075 (N_10075,N_9737,N_9735);
nor U10076 (N_10076,N_9923,N_9675);
nor U10077 (N_10077,N_9577,N_9503);
nand U10078 (N_10078,N_9841,N_9978);
nand U10079 (N_10079,N_9576,N_9970);
nand U10080 (N_10080,N_9843,N_9557);
and U10081 (N_10081,N_9669,N_9836);
xnor U10082 (N_10082,N_9667,N_9682);
nand U10083 (N_10083,N_9961,N_9687);
and U10084 (N_10084,N_9653,N_9645);
or U10085 (N_10085,N_9835,N_9698);
nand U10086 (N_10086,N_9995,N_9968);
nor U10087 (N_10087,N_9777,N_9988);
and U10088 (N_10088,N_9890,N_9525);
or U10089 (N_10089,N_9623,N_9756);
nand U10090 (N_10090,N_9754,N_9966);
nand U10091 (N_10091,N_9554,N_9906);
or U10092 (N_10092,N_9997,N_9991);
nand U10093 (N_10093,N_9590,N_9566);
nand U10094 (N_10094,N_9969,N_9757);
or U10095 (N_10095,N_9830,N_9510);
nor U10096 (N_10096,N_9870,N_9521);
and U10097 (N_10097,N_9550,N_9942);
nand U10098 (N_10098,N_9872,N_9597);
or U10099 (N_10099,N_9519,N_9732);
xor U10100 (N_10100,N_9977,N_9876);
nand U10101 (N_10101,N_9599,N_9741);
or U10102 (N_10102,N_9871,N_9904);
nor U10103 (N_10103,N_9866,N_9608);
xor U10104 (N_10104,N_9656,N_9765);
xor U10105 (N_10105,N_9840,N_9595);
xnor U10106 (N_10106,N_9903,N_9646);
nor U10107 (N_10107,N_9568,N_9779);
nor U10108 (N_10108,N_9855,N_9701);
nor U10109 (N_10109,N_9940,N_9697);
nand U10110 (N_10110,N_9571,N_9853);
nor U10111 (N_10111,N_9637,N_9593);
xor U10112 (N_10112,N_9658,N_9955);
nor U10113 (N_10113,N_9826,N_9858);
xnor U10114 (N_10114,N_9823,N_9702);
xor U10115 (N_10115,N_9540,N_9629);
and U10116 (N_10116,N_9522,N_9791);
xnor U10117 (N_10117,N_9785,N_9561);
nand U10118 (N_10118,N_9705,N_9990);
nor U10119 (N_10119,N_9581,N_9861);
xnor U10120 (N_10120,N_9950,N_9892);
nor U10121 (N_10121,N_9973,N_9511);
or U10122 (N_10122,N_9559,N_9887);
nand U10123 (N_10123,N_9957,N_9901);
nand U10124 (N_10124,N_9986,N_9549);
and U10125 (N_10125,N_9831,N_9527);
nand U10126 (N_10126,N_9558,N_9720);
nor U10127 (N_10127,N_9578,N_9882);
or U10128 (N_10128,N_9793,N_9934);
and U10129 (N_10129,N_9617,N_9663);
or U10130 (N_10130,N_9569,N_9816);
or U10131 (N_10131,N_9936,N_9696);
or U10132 (N_10132,N_9722,N_9784);
nand U10133 (N_10133,N_9703,N_9926);
or U10134 (N_10134,N_9570,N_9947);
xor U10135 (N_10135,N_9749,N_9788);
or U10136 (N_10136,N_9850,N_9884);
and U10137 (N_10137,N_9533,N_9627);
or U10138 (N_10138,N_9960,N_9917);
or U10139 (N_10139,N_9547,N_9660);
xor U10140 (N_10140,N_9805,N_9582);
nor U10141 (N_10141,N_9772,N_9710);
or U10142 (N_10142,N_9695,N_9761);
nor U10143 (N_10143,N_9747,N_9659);
nand U10144 (N_10144,N_9641,N_9998);
and U10145 (N_10145,N_9615,N_9648);
xnor U10146 (N_10146,N_9902,N_9933);
xor U10147 (N_10147,N_9992,N_9536);
and U10148 (N_10148,N_9602,N_9808);
and U10149 (N_10149,N_9545,N_9657);
nor U10150 (N_10150,N_9854,N_9939);
nor U10151 (N_10151,N_9971,N_9781);
nor U10152 (N_10152,N_9541,N_9679);
nand U10153 (N_10153,N_9721,N_9530);
nor U10154 (N_10154,N_9987,N_9804);
nor U10155 (N_10155,N_9596,N_9632);
or U10156 (N_10156,N_9584,N_9528);
nand U10157 (N_10157,N_9654,N_9797);
nand U10158 (N_10158,N_9774,N_9821);
xor U10159 (N_10159,N_9938,N_9736);
nand U10160 (N_10160,N_9746,N_9723);
nor U10161 (N_10161,N_9976,N_9692);
or U10162 (N_10162,N_9924,N_9878);
or U10163 (N_10163,N_9700,N_9989);
nand U10164 (N_10164,N_9762,N_9915);
nand U10165 (N_10165,N_9575,N_9706);
xor U10166 (N_10166,N_9851,N_9857);
nand U10167 (N_10167,N_9725,N_9638);
nor U10168 (N_10168,N_9982,N_9752);
nand U10169 (N_10169,N_9612,N_9729);
nor U10170 (N_10170,N_9589,N_9959);
nand U10171 (N_10171,N_9809,N_9726);
nand U10172 (N_10172,N_9651,N_9744);
and U10173 (N_10173,N_9996,N_9715);
nand U10174 (N_10174,N_9941,N_9766);
nor U10175 (N_10175,N_9748,N_9869);
xnor U10176 (N_10176,N_9814,N_9935);
xor U10177 (N_10177,N_9864,N_9644);
or U10178 (N_10178,N_9845,N_9745);
nand U10179 (N_10179,N_9516,N_9620);
or U10180 (N_10180,N_9879,N_9846);
or U10181 (N_10181,N_9693,N_9859);
and U10182 (N_10182,N_9776,N_9524);
nor U10183 (N_10183,N_9881,N_9815);
xnor U10184 (N_10184,N_9583,N_9909);
and U10185 (N_10185,N_9734,N_9740);
xnor U10186 (N_10186,N_9731,N_9834);
xor U10187 (N_10187,N_9932,N_9775);
xnor U10188 (N_10188,N_9964,N_9604);
or U10189 (N_10189,N_9709,N_9862);
or U10190 (N_10190,N_9630,N_9591);
and U10191 (N_10191,N_9803,N_9770);
xnor U10192 (N_10192,N_9994,N_9625);
nor U10193 (N_10193,N_9944,N_9670);
xor U10194 (N_10194,N_9662,N_9717);
nor U10195 (N_10195,N_9883,N_9555);
and U10196 (N_10196,N_9948,N_9811);
xor U10197 (N_10197,N_9965,N_9865);
or U10198 (N_10198,N_9962,N_9897);
nand U10199 (N_10199,N_9512,N_9829);
nor U10200 (N_10200,N_9895,N_9822);
nor U10201 (N_10201,N_9863,N_9560);
xor U10202 (N_10202,N_9920,N_9888);
nand U10203 (N_10203,N_9742,N_9921);
and U10204 (N_10204,N_9755,N_9886);
nor U10205 (N_10205,N_9618,N_9789);
and U10206 (N_10206,N_9553,N_9875);
and U10207 (N_10207,N_9898,N_9983);
nand U10208 (N_10208,N_9634,N_9543);
and U10209 (N_10209,N_9999,N_9782);
nand U10210 (N_10210,N_9818,N_9567);
nand U10211 (N_10211,N_9847,N_9839);
or U10212 (N_10212,N_9537,N_9718);
xnor U10213 (N_10213,N_9910,N_9642);
xor U10214 (N_10214,N_9880,N_9929);
xor U10215 (N_10215,N_9601,N_9728);
or U10216 (N_10216,N_9626,N_9984);
and U10217 (N_10217,N_9760,N_9727);
nand U10218 (N_10218,N_9896,N_9515);
nor U10219 (N_10219,N_9780,N_9551);
or U10220 (N_10220,N_9820,N_9751);
xnor U10221 (N_10221,N_9650,N_9520);
xnor U10222 (N_10222,N_9827,N_9526);
nand U10223 (N_10223,N_9678,N_9611);
nor U10224 (N_10224,N_9877,N_9680);
xor U10225 (N_10225,N_9563,N_9552);
nor U10226 (N_10226,N_9919,N_9833);
nand U10227 (N_10227,N_9529,N_9573);
nor U10228 (N_10228,N_9518,N_9673);
and U10229 (N_10229,N_9683,N_9763);
nand U10230 (N_10230,N_9514,N_9574);
xor U10231 (N_10231,N_9916,N_9773);
xnor U10232 (N_10232,N_9874,N_9535);
and U10233 (N_10233,N_9806,N_9500);
or U10234 (N_10234,N_9665,N_9640);
or U10235 (N_10235,N_9930,N_9538);
and U10236 (N_10236,N_9928,N_9787);
nand U10237 (N_10237,N_9689,N_9652);
or U10238 (N_10238,N_9813,N_9975);
xnor U10239 (N_10239,N_9794,N_9677);
xor U10240 (N_10240,N_9699,N_9639);
xor U10241 (N_10241,N_9868,N_9605);
and U10242 (N_10242,N_9943,N_9666);
or U10243 (N_10243,N_9713,N_9828);
and U10244 (N_10244,N_9807,N_9707);
and U10245 (N_10245,N_9686,N_9633);
and U10246 (N_10246,N_9501,N_9614);
nand U10247 (N_10247,N_9621,N_9952);
nor U10248 (N_10248,N_9993,N_9509);
nand U10249 (N_10249,N_9985,N_9636);
nor U10250 (N_10250,N_9660,N_9633);
nor U10251 (N_10251,N_9644,N_9685);
and U10252 (N_10252,N_9810,N_9670);
or U10253 (N_10253,N_9748,N_9605);
and U10254 (N_10254,N_9905,N_9656);
nor U10255 (N_10255,N_9769,N_9591);
nor U10256 (N_10256,N_9874,N_9759);
or U10257 (N_10257,N_9916,N_9809);
nor U10258 (N_10258,N_9522,N_9995);
and U10259 (N_10259,N_9569,N_9669);
nand U10260 (N_10260,N_9620,N_9791);
nand U10261 (N_10261,N_9684,N_9529);
xor U10262 (N_10262,N_9538,N_9628);
or U10263 (N_10263,N_9776,N_9681);
nand U10264 (N_10264,N_9730,N_9821);
nor U10265 (N_10265,N_9746,N_9565);
nand U10266 (N_10266,N_9885,N_9787);
nor U10267 (N_10267,N_9658,N_9945);
xor U10268 (N_10268,N_9628,N_9607);
xor U10269 (N_10269,N_9796,N_9811);
or U10270 (N_10270,N_9992,N_9966);
or U10271 (N_10271,N_9508,N_9728);
xnor U10272 (N_10272,N_9965,N_9695);
nor U10273 (N_10273,N_9686,N_9783);
or U10274 (N_10274,N_9970,N_9931);
nand U10275 (N_10275,N_9774,N_9685);
nand U10276 (N_10276,N_9537,N_9965);
nor U10277 (N_10277,N_9532,N_9865);
or U10278 (N_10278,N_9722,N_9962);
nand U10279 (N_10279,N_9877,N_9797);
or U10280 (N_10280,N_9639,N_9814);
xor U10281 (N_10281,N_9643,N_9714);
xnor U10282 (N_10282,N_9984,N_9532);
nand U10283 (N_10283,N_9550,N_9742);
xor U10284 (N_10284,N_9980,N_9599);
and U10285 (N_10285,N_9553,N_9813);
nand U10286 (N_10286,N_9771,N_9539);
and U10287 (N_10287,N_9565,N_9927);
and U10288 (N_10288,N_9894,N_9535);
and U10289 (N_10289,N_9742,N_9738);
and U10290 (N_10290,N_9708,N_9915);
or U10291 (N_10291,N_9918,N_9662);
or U10292 (N_10292,N_9960,N_9870);
xor U10293 (N_10293,N_9607,N_9511);
nand U10294 (N_10294,N_9829,N_9515);
and U10295 (N_10295,N_9747,N_9505);
and U10296 (N_10296,N_9765,N_9546);
nor U10297 (N_10297,N_9884,N_9670);
or U10298 (N_10298,N_9927,N_9809);
nand U10299 (N_10299,N_9752,N_9748);
nor U10300 (N_10300,N_9769,N_9545);
nor U10301 (N_10301,N_9620,N_9827);
or U10302 (N_10302,N_9968,N_9721);
xnor U10303 (N_10303,N_9819,N_9739);
nand U10304 (N_10304,N_9882,N_9642);
and U10305 (N_10305,N_9972,N_9502);
xor U10306 (N_10306,N_9642,N_9740);
xor U10307 (N_10307,N_9710,N_9826);
xor U10308 (N_10308,N_9658,N_9884);
or U10309 (N_10309,N_9673,N_9649);
or U10310 (N_10310,N_9986,N_9951);
xor U10311 (N_10311,N_9898,N_9856);
or U10312 (N_10312,N_9532,N_9848);
nand U10313 (N_10313,N_9905,N_9889);
nor U10314 (N_10314,N_9683,N_9648);
xor U10315 (N_10315,N_9717,N_9653);
nor U10316 (N_10316,N_9936,N_9868);
xnor U10317 (N_10317,N_9771,N_9803);
nand U10318 (N_10318,N_9839,N_9788);
xnor U10319 (N_10319,N_9903,N_9778);
nand U10320 (N_10320,N_9565,N_9668);
nand U10321 (N_10321,N_9913,N_9886);
or U10322 (N_10322,N_9568,N_9937);
and U10323 (N_10323,N_9993,N_9941);
or U10324 (N_10324,N_9703,N_9994);
nor U10325 (N_10325,N_9830,N_9961);
nand U10326 (N_10326,N_9736,N_9881);
or U10327 (N_10327,N_9644,N_9687);
and U10328 (N_10328,N_9642,N_9801);
nor U10329 (N_10329,N_9703,N_9806);
or U10330 (N_10330,N_9702,N_9773);
nand U10331 (N_10331,N_9886,N_9804);
or U10332 (N_10332,N_9976,N_9642);
xnor U10333 (N_10333,N_9728,N_9598);
and U10334 (N_10334,N_9873,N_9679);
nor U10335 (N_10335,N_9621,N_9930);
or U10336 (N_10336,N_9553,N_9565);
or U10337 (N_10337,N_9808,N_9635);
nand U10338 (N_10338,N_9981,N_9739);
nand U10339 (N_10339,N_9906,N_9997);
nand U10340 (N_10340,N_9803,N_9794);
and U10341 (N_10341,N_9709,N_9563);
nor U10342 (N_10342,N_9730,N_9767);
and U10343 (N_10343,N_9877,N_9972);
xnor U10344 (N_10344,N_9910,N_9748);
nor U10345 (N_10345,N_9553,N_9652);
and U10346 (N_10346,N_9832,N_9531);
xnor U10347 (N_10347,N_9821,N_9773);
and U10348 (N_10348,N_9757,N_9656);
and U10349 (N_10349,N_9863,N_9999);
xor U10350 (N_10350,N_9825,N_9997);
or U10351 (N_10351,N_9802,N_9688);
nor U10352 (N_10352,N_9572,N_9919);
or U10353 (N_10353,N_9692,N_9674);
or U10354 (N_10354,N_9813,N_9814);
nor U10355 (N_10355,N_9816,N_9829);
nand U10356 (N_10356,N_9528,N_9567);
and U10357 (N_10357,N_9815,N_9597);
or U10358 (N_10358,N_9918,N_9862);
xor U10359 (N_10359,N_9575,N_9900);
xnor U10360 (N_10360,N_9795,N_9939);
or U10361 (N_10361,N_9963,N_9798);
and U10362 (N_10362,N_9679,N_9825);
xor U10363 (N_10363,N_9589,N_9766);
and U10364 (N_10364,N_9890,N_9582);
nand U10365 (N_10365,N_9619,N_9755);
nor U10366 (N_10366,N_9554,N_9512);
or U10367 (N_10367,N_9587,N_9751);
nor U10368 (N_10368,N_9532,N_9571);
or U10369 (N_10369,N_9733,N_9897);
xnor U10370 (N_10370,N_9559,N_9994);
or U10371 (N_10371,N_9708,N_9521);
nor U10372 (N_10372,N_9692,N_9981);
and U10373 (N_10373,N_9959,N_9815);
nand U10374 (N_10374,N_9929,N_9755);
nand U10375 (N_10375,N_9766,N_9762);
xnor U10376 (N_10376,N_9674,N_9847);
xor U10377 (N_10377,N_9711,N_9511);
nor U10378 (N_10378,N_9627,N_9828);
xnor U10379 (N_10379,N_9812,N_9599);
and U10380 (N_10380,N_9913,N_9633);
xor U10381 (N_10381,N_9651,N_9722);
nor U10382 (N_10382,N_9516,N_9915);
nor U10383 (N_10383,N_9788,N_9829);
nor U10384 (N_10384,N_9861,N_9520);
and U10385 (N_10385,N_9838,N_9571);
or U10386 (N_10386,N_9923,N_9606);
nand U10387 (N_10387,N_9691,N_9544);
or U10388 (N_10388,N_9713,N_9510);
or U10389 (N_10389,N_9769,N_9750);
and U10390 (N_10390,N_9980,N_9864);
xor U10391 (N_10391,N_9690,N_9831);
or U10392 (N_10392,N_9829,N_9915);
and U10393 (N_10393,N_9803,N_9576);
nand U10394 (N_10394,N_9742,N_9807);
or U10395 (N_10395,N_9809,N_9958);
nand U10396 (N_10396,N_9922,N_9818);
nor U10397 (N_10397,N_9970,N_9672);
xnor U10398 (N_10398,N_9726,N_9615);
nand U10399 (N_10399,N_9979,N_9549);
nor U10400 (N_10400,N_9886,N_9668);
xor U10401 (N_10401,N_9578,N_9521);
nand U10402 (N_10402,N_9769,N_9516);
or U10403 (N_10403,N_9568,N_9579);
and U10404 (N_10404,N_9723,N_9999);
nor U10405 (N_10405,N_9575,N_9735);
xor U10406 (N_10406,N_9542,N_9643);
nor U10407 (N_10407,N_9802,N_9978);
or U10408 (N_10408,N_9984,N_9658);
nor U10409 (N_10409,N_9797,N_9970);
xor U10410 (N_10410,N_9620,N_9904);
or U10411 (N_10411,N_9936,N_9838);
and U10412 (N_10412,N_9752,N_9928);
and U10413 (N_10413,N_9713,N_9728);
nor U10414 (N_10414,N_9790,N_9804);
or U10415 (N_10415,N_9853,N_9779);
and U10416 (N_10416,N_9971,N_9811);
or U10417 (N_10417,N_9796,N_9725);
and U10418 (N_10418,N_9738,N_9735);
nor U10419 (N_10419,N_9791,N_9602);
nor U10420 (N_10420,N_9570,N_9998);
or U10421 (N_10421,N_9541,N_9968);
nand U10422 (N_10422,N_9749,N_9559);
nor U10423 (N_10423,N_9876,N_9887);
xor U10424 (N_10424,N_9557,N_9674);
and U10425 (N_10425,N_9987,N_9826);
nor U10426 (N_10426,N_9966,N_9816);
xor U10427 (N_10427,N_9897,N_9604);
xnor U10428 (N_10428,N_9575,N_9574);
nor U10429 (N_10429,N_9757,N_9879);
xor U10430 (N_10430,N_9971,N_9824);
xnor U10431 (N_10431,N_9939,N_9981);
xor U10432 (N_10432,N_9932,N_9802);
and U10433 (N_10433,N_9970,N_9839);
and U10434 (N_10434,N_9632,N_9695);
nor U10435 (N_10435,N_9762,N_9798);
and U10436 (N_10436,N_9897,N_9730);
nand U10437 (N_10437,N_9549,N_9753);
or U10438 (N_10438,N_9640,N_9526);
xor U10439 (N_10439,N_9673,N_9652);
nand U10440 (N_10440,N_9990,N_9666);
nor U10441 (N_10441,N_9979,N_9878);
xor U10442 (N_10442,N_9721,N_9982);
xor U10443 (N_10443,N_9581,N_9803);
xor U10444 (N_10444,N_9593,N_9566);
or U10445 (N_10445,N_9579,N_9559);
nand U10446 (N_10446,N_9794,N_9582);
nand U10447 (N_10447,N_9546,N_9937);
nand U10448 (N_10448,N_9989,N_9503);
nand U10449 (N_10449,N_9931,N_9563);
xnor U10450 (N_10450,N_9539,N_9587);
or U10451 (N_10451,N_9585,N_9599);
and U10452 (N_10452,N_9678,N_9772);
nor U10453 (N_10453,N_9981,N_9533);
or U10454 (N_10454,N_9604,N_9662);
nand U10455 (N_10455,N_9507,N_9554);
nand U10456 (N_10456,N_9536,N_9889);
nand U10457 (N_10457,N_9750,N_9540);
nand U10458 (N_10458,N_9603,N_9611);
nand U10459 (N_10459,N_9730,N_9800);
nand U10460 (N_10460,N_9811,N_9737);
and U10461 (N_10461,N_9985,N_9829);
xor U10462 (N_10462,N_9536,N_9762);
xor U10463 (N_10463,N_9943,N_9740);
nor U10464 (N_10464,N_9935,N_9561);
nand U10465 (N_10465,N_9798,N_9515);
and U10466 (N_10466,N_9990,N_9955);
or U10467 (N_10467,N_9643,N_9548);
or U10468 (N_10468,N_9602,N_9715);
nor U10469 (N_10469,N_9812,N_9763);
and U10470 (N_10470,N_9888,N_9863);
and U10471 (N_10471,N_9628,N_9728);
nand U10472 (N_10472,N_9730,N_9752);
nor U10473 (N_10473,N_9909,N_9952);
nand U10474 (N_10474,N_9971,N_9705);
or U10475 (N_10475,N_9939,N_9917);
and U10476 (N_10476,N_9818,N_9677);
nand U10477 (N_10477,N_9510,N_9568);
and U10478 (N_10478,N_9918,N_9602);
and U10479 (N_10479,N_9611,N_9867);
xor U10480 (N_10480,N_9838,N_9970);
nor U10481 (N_10481,N_9836,N_9505);
nor U10482 (N_10482,N_9550,N_9637);
nand U10483 (N_10483,N_9822,N_9932);
and U10484 (N_10484,N_9827,N_9987);
or U10485 (N_10485,N_9610,N_9871);
nand U10486 (N_10486,N_9582,N_9598);
or U10487 (N_10487,N_9632,N_9810);
xnor U10488 (N_10488,N_9502,N_9653);
nand U10489 (N_10489,N_9547,N_9910);
nor U10490 (N_10490,N_9617,N_9696);
nor U10491 (N_10491,N_9945,N_9513);
or U10492 (N_10492,N_9543,N_9632);
and U10493 (N_10493,N_9774,N_9832);
and U10494 (N_10494,N_9600,N_9673);
or U10495 (N_10495,N_9536,N_9972);
and U10496 (N_10496,N_9902,N_9517);
and U10497 (N_10497,N_9708,N_9947);
xnor U10498 (N_10498,N_9542,N_9691);
and U10499 (N_10499,N_9761,N_9768);
and U10500 (N_10500,N_10356,N_10490);
nand U10501 (N_10501,N_10331,N_10128);
nor U10502 (N_10502,N_10444,N_10120);
nand U10503 (N_10503,N_10153,N_10189);
nand U10504 (N_10504,N_10085,N_10381);
or U10505 (N_10505,N_10240,N_10148);
nor U10506 (N_10506,N_10141,N_10241);
nand U10507 (N_10507,N_10345,N_10338);
xnor U10508 (N_10508,N_10266,N_10212);
or U10509 (N_10509,N_10409,N_10040);
nand U10510 (N_10510,N_10497,N_10406);
and U10511 (N_10511,N_10021,N_10301);
or U10512 (N_10512,N_10306,N_10066);
nand U10513 (N_10513,N_10080,N_10006);
xnor U10514 (N_10514,N_10319,N_10395);
or U10515 (N_10515,N_10161,N_10015);
and U10516 (N_10516,N_10482,N_10320);
nor U10517 (N_10517,N_10317,N_10463);
and U10518 (N_10518,N_10048,N_10252);
nand U10519 (N_10519,N_10346,N_10344);
nand U10520 (N_10520,N_10350,N_10260);
and U10521 (N_10521,N_10451,N_10073);
xor U10522 (N_10522,N_10322,N_10079);
xor U10523 (N_10523,N_10465,N_10429);
and U10524 (N_10524,N_10475,N_10173);
or U10525 (N_10525,N_10480,N_10106);
or U10526 (N_10526,N_10283,N_10334);
or U10527 (N_10527,N_10432,N_10191);
and U10528 (N_10528,N_10385,N_10363);
or U10529 (N_10529,N_10370,N_10354);
xor U10530 (N_10530,N_10425,N_10010);
nor U10531 (N_10531,N_10330,N_10027);
and U10532 (N_10532,N_10300,N_10478);
nand U10533 (N_10533,N_10324,N_10336);
or U10534 (N_10534,N_10488,N_10454);
xor U10535 (N_10535,N_10180,N_10019);
and U10536 (N_10536,N_10046,N_10155);
nor U10537 (N_10537,N_10167,N_10438);
nor U10538 (N_10538,N_10479,N_10119);
or U10539 (N_10539,N_10127,N_10459);
nor U10540 (N_10540,N_10380,N_10215);
and U10541 (N_10541,N_10034,N_10211);
xnor U10542 (N_10542,N_10121,N_10263);
or U10543 (N_10543,N_10071,N_10284);
and U10544 (N_10544,N_10113,N_10043);
and U10545 (N_10545,N_10170,N_10485);
or U10546 (N_10546,N_10014,N_10225);
nor U10547 (N_10547,N_10471,N_10236);
and U10548 (N_10548,N_10011,N_10058);
nor U10549 (N_10549,N_10393,N_10064);
or U10550 (N_10550,N_10295,N_10233);
xnor U10551 (N_10551,N_10168,N_10188);
or U10552 (N_10552,N_10256,N_10415);
nor U10553 (N_10553,N_10313,N_10428);
or U10554 (N_10554,N_10414,N_10387);
xnor U10555 (N_10555,N_10224,N_10194);
and U10556 (N_10556,N_10181,N_10392);
or U10557 (N_10557,N_10361,N_10422);
nor U10558 (N_10558,N_10205,N_10455);
and U10559 (N_10559,N_10223,N_10061);
xnor U10560 (N_10560,N_10162,N_10424);
nor U10561 (N_10561,N_10376,N_10367);
nand U10562 (N_10562,N_10008,N_10159);
xor U10563 (N_10563,N_10464,N_10391);
nor U10564 (N_10564,N_10202,N_10469);
or U10565 (N_10565,N_10467,N_10124);
nor U10566 (N_10566,N_10003,N_10386);
xnor U10567 (N_10567,N_10164,N_10311);
nand U10568 (N_10568,N_10292,N_10342);
and U10569 (N_10569,N_10107,N_10435);
nand U10570 (N_10570,N_10190,N_10213);
nand U10571 (N_10571,N_10209,N_10453);
nand U10572 (N_10572,N_10031,N_10253);
nor U10573 (N_10573,N_10445,N_10243);
nor U10574 (N_10574,N_10166,N_10023);
or U10575 (N_10575,N_10374,N_10474);
xor U10576 (N_10576,N_10275,N_10053);
nor U10577 (N_10577,N_10498,N_10192);
and U10578 (N_10578,N_10144,N_10130);
xnor U10579 (N_10579,N_10030,N_10210);
nor U10580 (N_10580,N_10169,N_10217);
nor U10581 (N_10581,N_10355,N_10197);
xnor U10582 (N_10582,N_10443,N_10093);
or U10583 (N_10583,N_10232,N_10154);
and U10584 (N_10584,N_10137,N_10327);
nand U10585 (N_10585,N_10257,N_10045);
or U10586 (N_10586,N_10114,N_10383);
xnor U10587 (N_10587,N_10165,N_10449);
or U10588 (N_10588,N_10112,N_10084);
nor U10589 (N_10589,N_10271,N_10491);
or U10590 (N_10590,N_10298,N_10372);
xnor U10591 (N_10591,N_10065,N_10270);
and U10592 (N_10592,N_10484,N_10303);
nor U10593 (N_10593,N_10005,N_10407);
nor U10594 (N_10594,N_10204,N_10001);
xnor U10595 (N_10595,N_10090,N_10201);
nand U10596 (N_10596,N_10117,N_10390);
nand U10597 (N_10597,N_10452,N_10447);
and U10598 (N_10598,N_10134,N_10289);
nand U10599 (N_10599,N_10294,N_10230);
and U10600 (N_10600,N_10365,N_10104);
nor U10601 (N_10601,N_10494,N_10226);
or U10602 (N_10602,N_10126,N_10216);
xor U10603 (N_10603,N_10069,N_10096);
nor U10604 (N_10604,N_10078,N_10229);
or U10605 (N_10605,N_10072,N_10446);
and U10606 (N_10606,N_10401,N_10214);
and U10607 (N_10607,N_10492,N_10091);
or U10608 (N_10608,N_10131,N_10441);
xor U10609 (N_10609,N_10097,N_10087);
and U10610 (N_10610,N_10321,N_10369);
or U10611 (N_10611,N_10403,N_10095);
xor U10612 (N_10612,N_10255,N_10368);
or U10613 (N_10613,N_10411,N_10325);
and U10614 (N_10614,N_10456,N_10273);
or U10615 (N_10615,N_10122,N_10196);
nor U10616 (N_10616,N_10457,N_10423);
nor U10617 (N_10617,N_10269,N_10047);
or U10618 (N_10618,N_10089,N_10203);
or U10619 (N_10619,N_10486,N_10234);
or U10620 (N_10620,N_10267,N_10140);
nor U10621 (N_10621,N_10183,N_10404);
nor U10622 (N_10622,N_10460,N_10110);
or U10623 (N_10623,N_10477,N_10296);
nor U10624 (N_10624,N_10378,N_10288);
or U10625 (N_10625,N_10326,N_10219);
nor U10626 (N_10626,N_10264,N_10012);
or U10627 (N_10627,N_10100,N_10357);
nand U10628 (N_10628,N_10402,N_10262);
xor U10629 (N_10629,N_10360,N_10426);
nand U10630 (N_10630,N_10417,N_10312);
xor U10631 (N_10631,N_10062,N_10060);
nand U10632 (N_10632,N_10323,N_10489);
xnor U10633 (N_10633,N_10156,N_10227);
or U10634 (N_10634,N_10115,N_10220);
xor U10635 (N_10635,N_10418,N_10462);
nand U10636 (N_10636,N_10029,N_10348);
xnor U10637 (N_10637,N_10208,N_10133);
nand U10638 (N_10638,N_10495,N_10245);
xnor U10639 (N_10639,N_10280,N_10341);
or U10640 (N_10640,N_10035,N_10198);
or U10641 (N_10641,N_10200,N_10086);
nand U10642 (N_10642,N_10185,N_10018);
and U10643 (N_10643,N_10304,N_10017);
xor U10644 (N_10644,N_10307,N_10055);
and U10645 (N_10645,N_10152,N_10318);
xnor U10646 (N_10646,N_10222,N_10314);
xor U10647 (N_10647,N_10057,N_10049);
or U10648 (N_10648,N_10237,N_10157);
nand U10649 (N_10649,N_10375,N_10297);
nand U10650 (N_10650,N_10412,N_10434);
nand U10651 (N_10651,N_10437,N_10458);
xnor U10652 (N_10652,N_10265,N_10351);
or U10653 (N_10653,N_10139,N_10033);
nand U10654 (N_10654,N_10362,N_10109);
nor U10655 (N_10655,N_10175,N_10329);
nor U10656 (N_10656,N_10051,N_10440);
or U10657 (N_10657,N_10081,N_10433);
and U10658 (N_10658,N_10146,N_10461);
xnor U10659 (N_10659,N_10163,N_10054);
xnor U10660 (N_10660,N_10339,N_10399);
xor U10661 (N_10661,N_10396,N_10416);
or U10662 (N_10662,N_10176,N_10305);
nand U10663 (N_10663,N_10042,N_10476);
nand U10664 (N_10664,N_10258,N_10427);
xor U10665 (N_10665,N_10025,N_10286);
and U10666 (N_10666,N_10013,N_10448);
nand U10667 (N_10667,N_10118,N_10472);
and U10668 (N_10668,N_10299,N_10002);
and U10669 (N_10669,N_10450,N_10218);
nor U10670 (N_10670,N_10244,N_10147);
or U10671 (N_10671,N_10470,N_10231);
xor U10672 (N_10672,N_10068,N_10359);
nor U10673 (N_10673,N_10083,N_10116);
xor U10674 (N_10674,N_10394,N_10171);
nor U10675 (N_10675,N_10493,N_10228);
and U10676 (N_10676,N_10349,N_10398);
nand U10677 (N_10677,N_10184,N_10182);
nand U10678 (N_10678,N_10092,N_10179);
xnor U10679 (N_10679,N_10287,N_10039);
nor U10680 (N_10680,N_10496,N_10102);
nor U10681 (N_10681,N_10276,N_10308);
xor U10682 (N_10682,N_10088,N_10259);
or U10683 (N_10683,N_10041,N_10187);
nor U10684 (N_10684,N_10291,N_10036);
nor U10685 (N_10685,N_10377,N_10405);
xor U10686 (N_10686,N_10340,N_10022);
nor U10687 (N_10687,N_10410,N_10431);
nand U10688 (N_10688,N_10101,N_10037);
or U10689 (N_10689,N_10111,N_10353);
and U10690 (N_10690,N_10004,N_10044);
and U10691 (N_10691,N_10366,N_10094);
or U10692 (N_10692,N_10364,N_10098);
nand U10693 (N_10693,N_10070,N_10347);
xnor U10694 (N_10694,N_10186,N_10150);
or U10695 (N_10695,N_10248,N_10076);
and U10696 (N_10696,N_10466,N_10178);
xor U10697 (N_10697,N_10274,N_10075);
and U10698 (N_10698,N_10268,N_10195);
xnor U10699 (N_10699,N_10108,N_10436);
xor U10700 (N_10700,N_10302,N_10142);
xor U10701 (N_10701,N_10123,N_10059);
or U10702 (N_10702,N_10174,N_10199);
xnor U10703 (N_10703,N_10473,N_10136);
xor U10704 (N_10704,N_10420,N_10028);
and U10705 (N_10705,N_10138,N_10238);
or U10706 (N_10706,N_10242,N_10293);
nand U10707 (N_10707,N_10333,N_10430);
xor U10708 (N_10708,N_10389,N_10082);
xor U10709 (N_10709,N_10193,N_10246);
and U10710 (N_10710,N_10132,N_10335);
nor U10711 (N_10711,N_10158,N_10056);
nand U10712 (N_10712,N_10105,N_10103);
or U10713 (N_10713,N_10397,N_10145);
nand U10714 (N_10714,N_10282,N_10468);
nor U10715 (N_10715,N_10074,N_10419);
and U10716 (N_10716,N_10413,N_10316);
xor U10717 (N_10717,N_10250,N_10177);
or U10718 (N_10718,N_10487,N_10063);
nor U10719 (N_10719,N_10099,N_10221);
or U10720 (N_10720,N_10254,N_10016);
xor U10721 (N_10721,N_10290,N_10024);
xnor U10722 (N_10722,N_10388,N_10249);
or U10723 (N_10723,N_10067,N_10247);
xnor U10724 (N_10724,N_10251,N_10400);
xor U10725 (N_10725,N_10382,N_10077);
nand U10726 (N_10726,N_10384,N_10135);
nand U10727 (N_10727,N_10125,N_10373);
nor U10728 (N_10728,N_10020,N_10129);
xor U10729 (N_10729,N_10358,N_10272);
nand U10730 (N_10730,N_10315,N_10481);
xor U10731 (N_10731,N_10285,N_10277);
xnor U10732 (N_10732,N_10151,N_10239);
xnor U10733 (N_10733,N_10337,N_10408);
and U10734 (N_10734,N_10310,N_10421);
nand U10735 (N_10735,N_10328,N_10149);
nor U10736 (N_10736,N_10499,N_10026);
nand U10737 (N_10737,N_10172,N_10309);
or U10738 (N_10738,N_10343,N_10009);
and U10739 (N_10739,N_10379,N_10442);
or U10740 (N_10740,N_10206,N_10332);
and U10741 (N_10741,N_10278,N_10483);
nor U10742 (N_10742,N_10371,N_10281);
or U10743 (N_10743,N_10143,N_10038);
xnor U10744 (N_10744,N_10000,N_10261);
or U10745 (N_10745,N_10207,N_10235);
nor U10746 (N_10746,N_10352,N_10052);
xnor U10747 (N_10747,N_10050,N_10160);
nor U10748 (N_10748,N_10439,N_10007);
nand U10749 (N_10749,N_10279,N_10032);
or U10750 (N_10750,N_10068,N_10214);
xnor U10751 (N_10751,N_10415,N_10267);
nor U10752 (N_10752,N_10058,N_10148);
xor U10753 (N_10753,N_10207,N_10274);
nor U10754 (N_10754,N_10122,N_10494);
nor U10755 (N_10755,N_10464,N_10205);
or U10756 (N_10756,N_10265,N_10386);
or U10757 (N_10757,N_10208,N_10228);
nor U10758 (N_10758,N_10302,N_10028);
nand U10759 (N_10759,N_10499,N_10241);
and U10760 (N_10760,N_10200,N_10074);
nor U10761 (N_10761,N_10329,N_10239);
nor U10762 (N_10762,N_10074,N_10111);
and U10763 (N_10763,N_10067,N_10198);
and U10764 (N_10764,N_10033,N_10223);
xnor U10765 (N_10765,N_10469,N_10224);
or U10766 (N_10766,N_10295,N_10308);
nand U10767 (N_10767,N_10058,N_10332);
xnor U10768 (N_10768,N_10497,N_10306);
or U10769 (N_10769,N_10256,N_10214);
or U10770 (N_10770,N_10379,N_10400);
xor U10771 (N_10771,N_10136,N_10345);
xor U10772 (N_10772,N_10386,N_10260);
xnor U10773 (N_10773,N_10239,N_10234);
xnor U10774 (N_10774,N_10362,N_10272);
xor U10775 (N_10775,N_10452,N_10178);
and U10776 (N_10776,N_10254,N_10366);
nor U10777 (N_10777,N_10390,N_10453);
or U10778 (N_10778,N_10083,N_10416);
xor U10779 (N_10779,N_10471,N_10207);
or U10780 (N_10780,N_10054,N_10483);
or U10781 (N_10781,N_10482,N_10378);
xnor U10782 (N_10782,N_10021,N_10043);
xnor U10783 (N_10783,N_10494,N_10240);
nor U10784 (N_10784,N_10398,N_10404);
nor U10785 (N_10785,N_10206,N_10273);
nand U10786 (N_10786,N_10416,N_10284);
xnor U10787 (N_10787,N_10443,N_10220);
or U10788 (N_10788,N_10402,N_10147);
nand U10789 (N_10789,N_10482,N_10072);
nor U10790 (N_10790,N_10329,N_10274);
or U10791 (N_10791,N_10069,N_10073);
nand U10792 (N_10792,N_10155,N_10043);
xor U10793 (N_10793,N_10305,N_10074);
or U10794 (N_10794,N_10433,N_10151);
or U10795 (N_10795,N_10402,N_10412);
nor U10796 (N_10796,N_10484,N_10361);
and U10797 (N_10797,N_10342,N_10010);
nand U10798 (N_10798,N_10148,N_10030);
and U10799 (N_10799,N_10231,N_10038);
or U10800 (N_10800,N_10213,N_10262);
nand U10801 (N_10801,N_10415,N_10168);
and U10802 (N_10802,N_10234,N_10344);
and U10803 (N_10803,N_10235,N_10239);
or U10804 (N_10804,N_10239,N_10396);
nor U10805 (N_10805,N_10348,N_10398);
xnor U10806 (N_10806,N_10082,N_10446);
nor U10807 (N_10807,N_10066,N_10462);
nor U10808 (N_10808,N_10269,N_10460);
nor U10809 (N_10809,N_10288,N_10154);
nand U10810 (N_10810,N_10407,N_10448);
nand U10811 (N_10811,N_10033,N_10327);
xor U10812 (N_10812,N_10332,N_10481);
xnor U10813 (N_10813,N_10275,N_10115);
nor U10814 (N_10814,N_10206,N_10109);
xor U10815 (N_10815,N_10279,N_10294);
nor U10816 (N_10816,N_10263,N_10195);
and U10817 (N_10817,N_10256,N_10359);
and U10818 (N_10818,N_10269,N_10192);
nor U10819 (N_10819,N_10023,N_10149);
nand U10820 (N_10820,N_10260,N_10477);
nor U10821 (N_10821,N_10196,N_10093);
xnor U10822 (N_10822,N_10221,N_10132);
nand U10823 (N_10823,N_10187,N_10199);
nand U10824 (N_10824,N_10064,N_10450);
xnor U10825 (N_10825,N_10232,N_10253);
or U10826 (N_10826,N_10268,N_10366);
or U10827 (N_10827,N_10458,N_10213);
xor U10828 (N_10828,N_10488,N_10305);
and U10829 (N_10829,N_10037,N_10313);
xor U10830 (N_10830,N_10397,N_10456);
and U10831 (N_10831,N_10188,N_10093);
xnor U10832 (N_10832,N_10085,N_10441);
xnor U10833 (N_10833,N_10032,N_10249);
and U10834 (N_10834,N_10340,N_10273);
xor U10835 (N_10835,N_10359,N_10123);
and U10836 (N_10836,N_10094,N_10338);
xor U10837 (N_10837,N_10179,N_10025);
nand U10838 (N_10838,N_10043,N_10038);
xnor U10839 (N_10839,N_10413,N_10064);
or U10840 (N_10840,N_10444,N_10304);
nor U10841 (N_10841,N_10478,N_10377);
or U10842 (N_10842,N_10329,N_10185);
nor U10843 (N_10843,N_10483,N_10153);
xnor U10844 (N_10844,N_10281,N_10314);
nand U10845 (N_10845,N_10465,N_10451);
or U10846 (N_10846,N_10408,N_10024);
and U10847 (N_10847,N_10071,N_10046);
xor U10848 (N_10848,N_10461,N_10496);
nand U10849 (N_10849,N_10018,N_10247);
xnor U10850 (N_10850,N_10244,N_10045);
and U10851 (N_10851,N_10493,N_10270);
and U10852 (N_10852,N_10090,N_10170);
xor U10853 (N_10853,N_10148,N_10010);
or U10854 (N_10854,N_10323,N_10388);
or U10855 (N_10855,N_10375,N_10497);
nor U10856 (N_10856,N_10303,N_10008);
xor U10857 (N_10857,N_10383,N_10477);
nor U10858 (N_10858,N_10146,N_10155);
and U10859 (N_10859,N_10360,N_10450);
nand U10860 (N_10860,N_10406,N_10489);
nor U10861 (N_10861,N_10328,N_10285);
nand U10862 (N_10862,N_10042,N_10283);
xor U10863 (N_10863,N_10440,N_10373);
or U10864 (N_10864,N_10034,N_10278);
and U10865 (N_10865,N_10384,N_10160);
and U10866 (N_10866,N_10004,N_10156);
or U10867 (N_10867,N_10107,N_10086);
nor U10868 (N_10868,N_10213,N_10168);
nor U10869 (N_10869,N_10449,N_10208);
xor U10870 (N_10870,N_10469,N_10119);
or U10871 (N_10871,N_10089,N_10452);
nor U10872 (N_10872,N_10458,N_10092);
and U10873 (N_10873,N_10376,N_10250);
xor U10874 (N_10874,N_10284,N_10461);
and U10875 (N_10875,N_10244,N_10153);
nand U10876 (N_10876,N_10349,N_10337);
nand U10877 (N_10877,N_10400,N_10343);
and U10878 (N_10878,N_10372,N_10264);
nor U10879 (N_10879,N_10089,N_10451);
or U10880 (N_10880,N_10435,N_10427);
xor U10881 (N_10881,N_10457,N_10039);
xor U10882 (N_10882,N_10427,N_10055);
and U10883 (N_10883,N_10325,N_10238);
or U10884 (N_10884,N_10217,N_10367);
and U10885 (N_10885,N_10034,N_10286);
and U10886 (N_10886,N_10013,N_10447);
xnor U10887 (N_10887,N_10033,N_10069);
nand U10888 (N_10888,N_10460,N_10498);
nor U10889 (N_10889,N_10335,N_10163);
xnor U10890 (N_10890,N_10262,N_10366);
xor U10891 (N_10891,N_10027,N_10216);
xor U10892 (N_10892,N_10236,N_10179);
and U10893 (N_10893,N_10462,N_10439);
nand U10894 (N_10894,N_10408,N_10281);
xor U10895 (N_10895,N_10420,N_10152);
or U10896 (N_10896,N_10127,N_10264);
nor U10897 (N_10897,N_10107,N_10066);
or U10898 (N_10898,N_10149,N_10202);
nand U10899 (N_10899,N_10122,N_10174);
or U10900 (N_10900,N_10201,N_10292);
xor U10901 (N_10901,N_10275,N_10059);
and U10902 (N_10902,N_10338,N_10122);
and U10903 (N_10903,N_10496,N_10425);
xor U10904 (N_10904,N_10176,N_10350);
xnor U10905 (N_10905,N_10119,N_10053);
xnor U10906 (N_10906,N_10143,N_10467);
and U10907 (N_10907,N_10331,N_10374);
nand U10908 (N_10908,N_10322,N_10426);
and U10909 (N_10909,N_10191,N_10362);
xnor U10910 (N_10910,N_10153,N_10045);
xnor U10911 (N_10911,N_10004,N_10460);
or U10912 (N_10912,N_10246,N_10160);
nor U10913 (N_10913,N_10060,N_10177);
xor U10914 (N_10914,N_10140,N_10360);
and U10915 (N_10915,N_10139,N_10213);
and U10916 (N_10916,N_10157,N_10472);
xnor U10917 (N_10917,N_10328,N_10128);
or U10918 (N_10918,N_10336,N_10290);
or U10919 (N_10919,N_10155,N_10353);
and U10920 (N_10920,N_10458,N_10017);
or U10921 (N_10921,N_10157,N_10287);
or U10922 (N_10922,N_10363,N_10436);
and U10923 (N_10923,N_10428,N_10113);
xor U10924 (N_10924,N_10003,N_10199);
and U10925 (N_10925,N_10473,N_10410);
xor U10926 (N_10926,N_10254,N_10076);
nor U10927 (N_10927,N_10335,N_10045);
xor U10928 (N_10928,N_10028,N_10355);
and U10929 (N_10929,N_10123,N_10277);
xnor U10930 (N_10930,N_10318,N_10073);
and U10931 (N_10931,N_10026,N_10294);
or U10932 (N_10932,N_10152,N_10483);
and U10933 (N_10933,N_10392,N_10006);
nand U10934 (N_10934,N_10096,N_10427);
xnor U10935 (N_10935,N_10342,N_10233);
nand U10936 (N_10936,N_10475,N_10116);
xnor U10937 (N_10937,N_10268,N_10222);
nand U10938 (N_10938,N_10078,N_10161);
and U10939 (N_10939,N_10272,N_10395);
nor U10940 (N_10940,N_10420,N_10240);
xnor U10941 (N_10941,N_10348,N_10400);
xor U10942 (N_10942,N_10488,N_10071);
or U10943 (N_10943,N_10148,N_10126);
xor U10944 (N_10944,N_10096,N_10267);
xnor U10945 (N_10945,N_10230,N_10095);
nand U10946 (N_10946,N_10037,N_10489);
nand U10947 (N_10947,N_10324,N_10390);
and U10948 (N_10948,N_10008,N_10455);
and U10949 (N_10949,N_10327,N_10336);
or U10950 (N_10950,N_10252,N_10139);
xnor U10951 (N_10951,N_10114,N_10428);
or U10952 (N_10952,N_10476,N_10295);
xor U10953 (N_10953,N_10454,N_10117);
nor U10954 (N_10954,N_10427,N_10016);
xnor U10955 (N_10955,N_10265,N_10025);
nor U10956 (N_10956,N_10301,N_10107);
and U10957 (N_10957,N_10388,N_10035);
xnor U10958 (N_10958,N_10059,N_10497);
xor U10959 (N_10959,N_10000,N_10150);
and U10960 (N_10960,N_10047,N_10481);
nor U10961 (N_10961,N_10367,N_10191);
and U10962 (N_10962,N_10064,N_10063);
nand U10963 (N_10963,N_10221,N_10383);
or U10964 (N_10964,N_10429,N_10219);
nand U10965 (N_10965,N_10402,N_10311);
nand U10966 (N_10966,N_10319,N_10175);
nand U10967 (N_10967,N_10413,N_10380);
nand U10968 (N_10968,N_10015,N_10025);
xnor U10969 (N_10969,N_10320,N_10200);
nor U10970 (N_10970,N_10147,N_10411);
or U10971 (N_10971,N_10157,N_10413);
and U10972 (N_10972,N_10451,N_10247);
xor U10973 (N_10973,N_10027,N_10449);
nor U10974 (N_10974,N_10430,N_10090);
or U10975 (N_10975,N_10075,N_10105);
xnor U10976 (N_10976,N_10399,N_10204);
xor U10977 (N_10977,N_10042,N_10175);
and U10978 (N_10978,N_10216,N_10183);
xnor U10979 (N_10979,N_10226,N_10299);
nand U10980 (N_10980,N_10453,N_10383);
nor U10981 (N_10981,N_10120,N_10401);
and U10982 (N_10982,N_10034,N_10345);
xor U10983 (N_10983,N_10466,N_10056);
nand U10984 (N_10984,N_10190,N_10173);
and U10985 (N_10985,N_10004,N_10002);
or U10986 (N_10986,N_10144,N_10430);
nor U10987 (N_10987,N_10490,N_10151);
nand U10988 (N_10988,N_10360,N_10356);
nor U10989 (N_10989,N_10463,N_10014);
nand U10990 (N_10990,N_10329,N_10368);
nand U10991 (N_10991,N_10336,N_10425);
nand U10992 (N_10992,N_10471,N_10250);
nor U10993 (N_10993,N_10027,N_10270);
nand U10994 (N_10994,N_10108,N_10351);
nor U10995 (N_10995,N_10183,N_10354);
nand U10996 (N_10996,N_10099,N_10107);
and U10997 (N_10997,N_10187,N_10356);
and U10998 (N_10998,N_10447,N_10249);
nor U10999 (N_10999,N_10209,N_10135);
nor U11000 (N_11000,N_10814,N_10820);
nand U11001 (N_11001,N_10960,N_10708);
nor U11002 (N_11002,N_10548,N_10544);
and U11003 (N_11003,N_10679,N_10697);
nor U11004 (N_11004,N_10776,N_10660);
and U11005 (N_11005,N_10609,N_10846);
nor U11006 (N_11006,N_10604,N_10924);
and U11007 (N_11007,N_10718,N_10849);
nand U11008 (N_11008,N_10525,N_10900);
nor U11009 (N_11009,N_10564,N_10978);
nor U11010 (N_11010,N_10657,N_10957);
or U11011 (N_11011,N_10796,N_10508);
xnor U11012 (N_11012,N_10596,N_10744);
xor U11013 (N_11013,N_10944,N_10908);
nor U11014 (N_11014,N_10756,N_10738);
and U11015 (N_11015,N_10551,N_10654);
or U11016 (N_11016,N_10959,N_10536);
nor U11017 (N_11017,N_10748,N_10862);
nor U11018 (N_11018,N_10531,N_10932);
nand U11019 (N_11019,N_10636,N_10671);
xor U11020 (N_11020,N_10802,N_10579);
and U11021 (N_11021,N_10947,N_10894);
nor U11022 (N_11022,N_10887,N_10622);
nor U11023 (N_11023,N_10829,N_10865);
nand U11024 (N_11024,N_10784,N_10889);
and U11025 (N_11025,N_10674,N_10973);
and U11026 (N_11026,N_10639,N_10925);
and U11027 (N_11027,N_10937,N_10746);
or U11028 (N_11028,N_10812,N_10661);
nor U11029 (N_11029,N_10638,N_10730);
or U11030 (N_11030,N_10879,N_10943);
nor U11031 (N_11031,N_10755,N_10935);
xnor U11032 (N_11032,N_10543,N_10619);
nand U11033 (N_11033,N_10790,N_10595);
and U11034 (N_11034,N_10892,N_10689);
nand U11035 (N_11035,N_10620,N_10642);
nand U11036 (N_11036,N_10816,N_10628);
nand U11037 (N_11037,N_10538,N_10761);
nor U11038 (N_11038,N_10580,N_10968);
nand U11039 (N_11039,N_10653,N_10763);
xnor U11040 (N_11040,N_10570,N_10948);
or U11041 (N_11041,N_10860,N_10713);
nand U11042 (N_11042,N_10774,N_10612);
xor U11043 (N_11043,N_10714,N_10866);
nand U11044 (N_11044,N_10882,N_10555);
nand U11045 (N_11045,N_10861,N_10712);
or U11046 (N_11046,N_10810,N_10836);
nand U11047 (N_11047,N_10990,N_10702);
and U11048 (N_11048,N_10557,N_10837);
nor U11049 (N_11049,N_10877,N_10658);
nand U11050 (N_11050,N_10728,N_10747);
and U11051 (N_11051,N_10646,N_10926);
nor U11052 (N_11052,N_10845,N_10807);
nand U11053 (N_11053,N_10872,N_10858);
nor U11054 (N_11054,N_10617,N_10585);
or U11055 (N_11055,N_10535,N_10945);
nor U11056 (N_11056,N_10662,N_10840);
nor U11057 (N_11057,N_10794,N_10791);
or U11058 (N_11058,N_10772,N_10919);
xor U11059 (N_11059,N_10750,N_10667);
or U11060 (N_11060,N_10602,N_10830);
or U11061 (N_11061,N_10923,N_10610);
nor U11062 (N_11062,N_10921,N_10793);
or U11063 (N_11063,N_10690,N_10800);
xor U11064 (N_11064,N_10988,N_10847);
nor U11065 (N_11065,N_10682,N_10513);
and U11066 (N_11066,N_10951,N_10686);
xor U11067 (N_11067,N_10920,N_10561);
or U11068 (N_11068,N_10611,N_10504);
nor U11069 (N_11069,N_10695,N_10854);
and U11070 (N_11070,N_10618,N_10928);
nand U11071 (N_11071,N_10677,N_10905);
nand U11072 (N_11072,N_10896,N_10704);
or U11073 (N_11073,N_10852,N_10914);
nand U11074 (N_11074,N_10627,N_10599);
and U11075 (N_11075,N_10752,N_10521);
nor U11076 (N_11076,N_10833,N_10918);
or U11077 (N_11077,N_10949,N_10640);
xnor U11078 (N_11078,N_10777,N_10716);
nand U11079 (N_11079,N_10859,N_10885);
nand U11080 (N_11080,N_10815,N_10663);
or U11081 (N_11081,N_10700,N_10980);
nand U11082 (N_11082,N_10676,N_10715);
nor U11083 (N_11083,N_10792,N_10855);
nor U11084 (N_11084,N_10766,N_10529);
and U11085 (N_11085,N_10760,N_10933);
or U11086 (N_11086,N_10779,N_10668);
xor U11087 (N_11087,N_10517,N_10764);
nand U11088 (N_11088,N_10641,N_10701);
and U11089 (N_11089,N_10648,N_10939);
or U11090 (N_11090,N_10983,N_10912);
or U11091 (N_11091,N_10853,N_10821);
nor U11092 (N_11092,N_10563,N_10868);
or U11093 (N_11093,N_10706,N_10705);
xor U11094 (N_11094,N_10881,N_10964);
xor U11095 (N_11095,N_10616,N_10975);
nand U11096 (N_11096,N_10606,N_10736);
and U11097 (N_11097,N_10987,N_10664);
and U11098 (N_11098,N_10731,N_10934);
nor U11099 (N_11099,N_10799,N_10871);
and U11100 (N_11100,N_10592,N_10954);
nand U11101 (N_11101,N_10507,N_10514);
nor U11102 (N_11102,N_10675,N_10818);
xnor U11103 (N_11103,N_10647,N_10904);
or U11104 (N_11104,N_10808,N_10603);
nand U11105 (N_11105,N_10553,N_10981);
nand U11106 (N_11106,N_10629,N_10780);
nor U11107 (N_11107,N_10788,N_10897);
nand U11108 (N_11108,N_10518,N_10506);
nand U11109 (N_11109,N_10572,N_10588);
xnor U11110 (N_11110,N_10749,N_10838);
xor U11111 (N_11111,N_10566,N_10797);
nor U11112 (N_11112,N_10630,N_10771);
nor U11113 (N_11113,N_10832,N_10883);
nand U11114 (N_11114,N_10958,N_10888);
and U11115 (N_11115,N_10917,N_10565);
or U11116 (N_11116,N_10541,N_10526);
nor U11117 (N_11117,N_10971,N_10680);
or U11118 (N_11118,N_10965,N_10992);
nand U11119 (N_11119,N_10903,N_10576);
or U11120 (N_11120,N_10844,N_10783);
nor U11121 (N_11121,N_10733,N_10696);
or U11122 (N_11122,N_10737,N_10740);
and U11123 (N_11123,N_10589,N_10765);
nor U11124 (N_11124,N_10922,N_10528);
nand U11125 (N_11125,N_10574,N_10795);
nor U11126 (N_11126,N_10530,N_10607);
nor U11127 (N_11127,N_10575,N_10902);
nor U11128 (N_11128,N_10906,N_10540);
xor U11129 (N_11129,N_10621,N_10512);
or U11130 (N_11130,N_10550,N_10915);
nand U11131 (N_11131,N_10554,N_10880);
nor U11132 (N_11132,N_10962,N_10869);
and U11133 (N_11133,N_10966,N_10938);
and U11134 (N_11134,N_10963,N_10699);
nand U11135 (N_11135,N_10688,N_10825);
nand U11136 (N_11136,N_10527,N_10931);
xor U11137 (N_11137,N_10739,N_10623);
nor U11138 (N_11138,N_10991,N_10505);
nor U11139 (N_11139,N_10831,N_10632);
nor U11140 (N_11140,N_10974,N_10634);
nand U11141 (N_11141,N_10710,N_10930);
nand U11142 (N_11142,N_10758,N_10781);
or U11143 (N_11143,N_10590,N_10631);
and U11144 (N_11144,N_10834,N_10751);
or U11145 (N_11145,N_10510,N_10979);
nor U11146 (N_11146,N_10848,N_10643);
xnor U11147 (N_11147,N_10681,N_10542);
xor U11148 (N_11148,N_10719,N_10722);
xor U11149 (N_11149,N_10562,N_10522);
nand U11150 (N_11150,N_10961,N_10907);
nor U11151 (N_11151,N_10698,N_10594);
or U11152 (N_11152,N_10502,N_10605);
or U11153 (N_11153,N_10711,N_10984);
nand U11154 (N_11154,N_10878,N_10601);
or U11155 (N_11155,N_10672,N_10633);
nand U11156 (N_11156,N_10929,N_10539);
nor U11157 (N_11157,N_10635,N_10941);
and U11158 (N_11158,N_10916,N_10694);
or U11159 (N_11159,N_10656,N_10899);
or U11160 (N_11160,N_10863,N_10598);
and U11161 (N_11161,N_10501,N_10754);
and U11162 (N_11162,N_10996,N_10613);
xor U11163 (N_11163,N_10586,N_10841);
or U11164 (N_11164,N_10851,N_10560);
nand U11165 (N_11165,N_10678,N_10684);
or U11166 (N_11166,N_10725,N_10687);
or U11167 (N_11167,N_10571,N_10952);
and U11168 (N_11168,N_10850,N_10967);
nor U11169 (N_11169,N_10927,N_10946);
or U11170 (N_11170,N_10890,N_10857);
nand U11171 (N_11171,N_10644,N_10614);
nand U11172 (N_11172,N_10950,N_10624);
nor U11173 (N_11173,N_10842,N_10826);
or U11174 (N_11174,N_10913,N_10552);
or U11175 (N_11175,N_10537,N_10666);
nand U11176 (N_11176,N_10515,N_10901);
nor U11177 (N_11177,N_10727,N_10549);
or U11178 (N_11178,N_10545,N_10856);
xnor U11179 (N_11179,N_10985,N_10735);
and U11180 (N_11180,N_10823,N_10651);
xnor U11181 (N_11181,N_10649,N_10723);
nor U11182 (N_11182,N_10685,N_10753);
xnor U11183 (N_11183,N_10782,N_10509);
nand U11184 (N_11184,N_10762,N_10721);
xnor U11185 (N_11185,N_10801,N_10884);
and U11186 (N_11186,N_10745,N_10970);
or U11187 (N_11187,N_10803,N_10546);
nand U11188 (N_11188,N_10956,N_10669);
nand U11189 (N_11189,N_10615,N_10972);
or U11190 (N_11190,N_10843,N_10768);
or U11191 (N_11191,N_10670,N_10626);
or U11192 (N_11192,N_10798,N_10895);
nor U11193 (N_11193,N_10909,N_10720);
or U11194 (N_11194,N_10804,N_10717);
nand U11195 (N_11195,N_10625,N_10875);
nand U11196 (N_11196,N_10742,N_10819);
and U11197 (N_11197,N_10587,N_10982);
xnor U11198 (N_11198,N_10817,N_10910);
nor U11199 (N_11199,N_10683,N_10891);
nor U11200 (N_11200,N_10547,N_10759);
xor U11201 (N_11201,N_10876,N_10995);
xor U11202 (N_11202,N_10608,N_10989);
and U11203 (N_11203,N_10936,N_10828);
or U11204 (N_11204,N_10822,N_10559);
xnor U11205 (N_11205,N_10993,N_10953);
and U11206 (N_11206,N_10581,N_10955);
and U11207 (N_11207,N_10569,N_10556);
xor U11208 (N_11208,N_10809,N_10806);
xnor U11209 (N_11209,N_10593,N_10874);
or U11210 (N_11210,N_10709,N_10597);
nor U11211 (N_11211,N_10976,N_10584);
or U11212 (N_11212,N_10691,N_10940);
xor U11213 (N_11213,N_10864,N_10534);
or U11214 (N_11214,N_10898,N_10650);
and U11215 (N_11215,N_10734,N_10665);
nor U11216 (N_11216,N_10789,N_10523);
nand U11217 (N_11217,N_10773,N_10835);
xor U11218 (N_11218,N_10583,N_10839);
and U11219 (N_11219,N_10533,N_10503);
or U11220 (N_11220,N_10977,N_10786);
nor U11221 (N_11221,N_10692,N_10998);
or U11222 (N_11222,N_10886,N_10591);
or U11223 (N_11223,N_10726,N_10813);
or U11224 (N_11224,N_10693,N_10787);
or U11225 (N_11225,N_10567,N_10811);
and U11226 (N_11226,N_10732,N_10520);
or U11227 (N_11227,N_10673,N_10757);
and U11228 (N_11228,N_10524,N_10600);
xor U11229 (N_11229,N_10893,N_10659);
and U11230 (N_11230,N_10743,N_10655);
nor U11231 (N_11231,N_10767,N_10994);
nand U11232 (N_11232,N_10873,N_10577);
or U11233 (N_11233,N_10769,N_10645);
nand U11234 (N_11234,N_10573,N_10724);
nand U11235 (N_11235,N_10511,N_10911);
or U11236 (N_11236,N_10775,N_10568);
nand U11237 (N_11237,N_10500,N_10805);
and U11238 (N_11238,N_10519,N_10867);
xnor U11239 (N_11239,N_10578,N_10558);
xor U11240 (N_11240,N_10707,N_10741);
and U11241 (N_11241,N_10827,N_10582);
or U11242 (N_11242,N_10870,N_10942);
or U11243 (N_11243,N_10652,N_10997);
or U11244 (N_11244,N_10999,N_10703);
nand U11245 (N_11245,N_10637,N_10516);
xnor U11246 (N_11246,N_10729,N_10770);
nand U11247 (N_11247,N_10986,N_10824);
or U11248 (N_11248,N_10969,N_10778);
xnor U11249 (N_11249,N_10785,N_10532);
nand U11250 (N_11250,N_10605,N_10607);
or U11251 (N_11251,N_10542,N_10501);
xor U11252 (N_11252,N_10979,N_10706);
nor U11253 (N_11253,N_10848,N_10640);
and U11254 (N_11254,N_10912,N_10937);
xor U11255 (N_11255,N_10555,N_10988);
nor U11256 (N_11256,N_10583,N_10853);
xnor U11257 (N_11257,N_10655,N_10542);
nand U11258 (N_11258,N_10787,N_10899);
nand U11259 (N_11259,N_10814,N_10665);
and U11260 (N_11260,N_10769,N_10697);
xor U11261 (N_11261,N_10827,N_10531);
and U11262 (N_11262,N_10892,N_10820);
and U11263 (N_11263,N_10885,N_10824);
nand U11264 (N_11264,N_10692,N_10606);
or U11265 (N_11265,N_10619,N_10944);
or U11266 (N_11266,N_10855,N_10578);
or U11267 (N_11267,N_10887,N_10940);
nand U11268 (N_11268,N_10860,N_10690);
xor U11269 (N_11269,N_10634,N_10530);
and U11270 (N_11270,N_10677,N_10807);
or U11271 (N_11271,N_10802,N_10511);
nor U11272 (N_11272,N_10571,N_10909);
xor U11273 (N_11273,N_10915,N_10866);
or U11274 (N_11274,N_10709,N_10897);
nand U11275 (N_11275,N_10527,N_10558);
and U11276 (N_11276,N_10510,N_10712);
and U11277 (N_11277,N_10730,N_10600);
and U11278 (N_11278,N_10753,N_10522);
nand U11279 (N_11279,N_10632,N_10856);
nor U11280 (N_11280,N_10933,N_10641);
xnor U11281 (N_11281,N_10600,N_10987);
or U11282 (N_11282,N_10836,N_10964);
or U11283 (N_11283,N_10900,N_10769);
or U11284 (N_11284,N_10615,N_10727);
nand U11285 (N_11285,N_10579,N_10667);
and U11286 (N_11286,N_10642,N_10991);
xor U11287 (N_11287,N_10542,N_10995);
nor U11288 (N_11288,N_10567,N_10753);
and U11289 (N_11289,N_10640,N_10941);
nand U11290 (N_11290,N_10939,N_10874);
or U11291 (N_11291,N_10877,N_10705);
and U11292 (N_11292,N_10532,N_10852);
nor U11293 (N_11293,N_10714,N_10673);
or U11294 (N_11294,N_10633,N_10869);
or U11295 (N_11295,N_10533,N_10711);
nor U11296 (N_11296,N_10967,N_10507);
nand U11297 (N_11297,N_10745,N_10660);
nand U11298 (N_11298,N_10928,N_10542);
and U11299 (N_11299,N_10722,N_10856);
or U11300 (N_11300,N_10830,N_10810);
nand U11301 (N_11301,N_10522,N_10729);
nand U11302 (N_11302,N_10948,N_10595);
nor U11303 (N_11303,N_10582,N_10790);
nor U11304 (N_11304,N_10915,N_10543);
and U11305 (N_11305,N_10698,N_10525);
or U11306 (N_11306,N_10999,N_10700);
nor U11307 (N_11307,N_10790,N_10756);
and U11308 (N_11308,N_10872,N_10656);
nor U11309 (N_11309,N_10631,N_10977);
xor U11310 (N_11310,N_10523,N_10742);
or U11311 (N_11311,N_10649,N_10539);
nor U11312 (N_11312,N_10848,N_10994);
xor U11313 (N_11313,N_10541,N_10686);
xor U11314 (N_11314,N_10856,N_10837);
xor U11315 (N_11315,N_10780,N_10910);
and U11316 (N_11316,N_10887,N_10832);
xnor U11317 (N_11317,N_10950,N_10918);
and U11318 (N_11318,N_10919,N_10828);
and U11319 (N_11319,N_10865,N_10569);
or U11320 (N_11320,N_10962,N_10996);
nand U11321 (N_11321,N_10711,N_10935);
xnor U11322 (N_11322,N_10627,N_10514);
or U11323 (N_11323,N_10746,N_10920);
or U11324 (N_11324,N_10538,N_10611);
and U11325 (N_11325,N_10625,N_10690);
xor U11326 (N_11326,N_10960,N_10915);
nor U11327 (N_11327,N_10619,N_10891);
nand U11328 (N_11328,N_10979,N_10974);
nand U11329 (N_11329,N_10535,N_10828);
nand U11330 (N_11330,N_10733,N_10869);
nor U11331 (N_11331,N_10681,N_10921);
nand U11332 (N_11332,N_10858,N_10709);
or U11333 (N_11333,N_10797,N_10749);
nand U11334 (N_11334,N_10611,N_10519);
nand U11335 (N_11335,N_10770,N_10553);
nand U11336 (N_11336,N_10598,N_10792);
and U11337 (N_11337,N_10651,N_10593);
and U11338 (N_11338,N_10601,N_10904);
xor U11339 (N_11339,N_10891,N_10506);
nand U11340 (N_11340,N_10883,N_10530);
xor U11341 (N_11341,N_10916,N_10610);
nand U11342 (N_11342,N_10601,N_10648);
and U11343 (N_11343,N_10682,N_10700);
and U11344 (N_11344,N_10647,N_10714);
nor U11345 (N_11345,N_10857,N_10714);
nor U11346 (N_11346,N_10789,N_10952);
xor U11347 (N_11347,N_10859,N_10661);
and U11348 (N_11348,N_10590,N_10533);
xor U11349 (N_11349,N_10867,N_10601);
and U11350 (N_11350,N_10975,N_10571);
xnor U11351 (N_11351,N_10502,N_10899);
nor U11352 (N_11352,N_10536,N_10754);
or U11353 (N_11353,N_10559,N_10524);
xnor U11354 (N_11354,N_10724,N_10666);
nor U11355 (N_11355,N_10569,N_10880);
nor U11356 (N_11356,N_10934,N_10860);
xnor U11357 (N_11357,N_10621,N_10635);
xor U11358 (N_11358,N_10968,N_10700);
xnor U11359 (N_11359,N_10538,N_10810);
xnor U11360 (N_11360,N_10674,N_10547);
nand U11361 (N_11361,N_10717,N_10737);
or U11362 (N_11362,N_10769,N_10700);
nor U11363 (N_11363,N_10593,N_10886);
and U11364 (N_11364,N_10652,N_10905);
or U11365 (N_11365,N_10546,N_10654);
nand U11366 (N_11366,N_10544,N_10864);
nor U11367 (N_11367,N_10618,N_10700);
and U11368 (N_11368,N_10799,N_10660);
nand U11369 (N_11369,N_10588,N_10867);
nor U11370 (N_11370,N_10785,N_10561);
nor U11371 (N_11371,N_10847,N_10629);
and U11372 (N_11372,N_10588,N_10981);
nor U11373 (N_11373,N_10543,N_10678);
and U11374 (N_11374,N_10561,N_10984);
nand U11375 (N_11375,N_10834,N_10620);
and U11376 (N_11376,N_10582,N_10798);
or U11377 (N_11377,N_10821,N_10797);
nor U11378 (N_11378,N_10691,N_10719);
or U11379 (N_11379,N_10513,N_10642);
and U11380 (N_11380,N_10624,N_10845);
and U11381 (N_11381,N_10792,N_10999);
nand U11382 (N_11382,N_10535,N_10913);
nor U11383 (N_11383,N_10526,N_10834);
xnor U11384 (N_11384,N_10715,N_10878);
xnor U11385 (N_11385,N_10916,N_10988);
or U11386 (N_11386,N_10663,N_10641);
xnor U11387 (N_11387,N_10613,N_10607);
nor U11388 (N_11388,N_10740,N_10507);
xor U11389 (N_11389,N_10629,N_10892);
or U11390 (N_11390,N_10691,N_10835);
or U11391 (N_11391,N_10965,N_10562);
xnor U11392 (N_11392,N_10898,N_10643);
nand U11393 (N_11393,N_10513,N_10591);
nor U11394 (N_11394,N_10893,N_10609);
xnor U11395 (N_11395,N_10986,N_10502);
xnor U11396 (N_11396,N_10813,N_10527);
nand U11397 (N_11397,N_10737,N_10643);
nand U11398 (N_11398,N_10990,N_10785);
and U11399 (N_11399,N_10683,N_10699);
nand U11400 (N_11400,N_10570,N_10800);
nand U11401 (N_11401,N_10802,N_10555);
nand U11402 (N_11402,N_10617,N_10771);
or U11403 (N_11403,N_10728,N_10946);
nand U11404 (N_11404,N_10618,N_10869);
xnor U11405 (N_11405,N_10703,N_10882);
and U11406 (N_11406,N_10820,N_10587);
or U11407 (N_11407,N_10632,N_10592);
xor U11408 (N_11408,N_10986,N_10560);
nor U11409 (N_11409,N_10653,N_10930);
nor U11410 (N_11410,N_10582,N_10507);
xnor U11411 (N_11411,N_10587,N_10835);
and U11412 (N_11412,N_10531,N_10929);
and U11413 (N_11413,N_10693,N_10878);
nand U11414 (N_11414,N_10717,N_10932);
or U11415 (N_11415,N_10820,N_10953);
nor U11416 (N_11416,N_10899,N_10568);
or U11417 (N_11417,N_10852,N_10965);
xor U11418 (N_11418,N_10758,N_10557);
xor U11419 (N_11419,N_10742,N_10536);
xor U11420 (N_11420,N_10560,N_10699);
xnor U11421 (N_11421,N_10751,N_10635);
nand U11422 (N_11422,N_10635,N_10587);
nand U11423 (N_11423,N_10579,N_10809);
nor U11424 (N_11424,N_10963,N_10875);
nor U11425 (N_11425,N_10784,N_10946);
nor U11426 (N_11426,N_10646,N_10698);
xor U11427 (N_11427,N_10718,N_10897);
and U11428 (N_11428,N_10758,N_10874);
nand U11429 (N_11429,N_10809,N_10816);
nor U11430 (N_11430,N_10979,N_10718);
and U11431 (N_11431,N_10549,N_10501);
and U11432 (N_11432,N_10518,N_10901);
xor U11433 (N_11433,N_10650,N_10600);
xor U11434 (N_11434,N_10550,N_10609);
xor U11435 (N_11435,N_10626,N_10584);
nor U11436 (N_11436,N_10639,N_10548);
or U11437 (N_11437,N_10954,N_10911);
and U11438 (N_11438,N_10620,N_10698);
or U11439 (N_11439,N_10530,N_10873);
nor U11440 (N_11440,N_10618,N_10698);
or U11441 (N_11441,N_10898,N_10736);
and U11442 (N_11442,N_10929,N_10882);
nand U11443 (N_11443,N_10945,N_10572);
xnor U11444 (N_11444,N_10568,N_10996);
and U11445 (N_11445,N_10575,N_10785);
nand U11446 (N_11446,N_10510,N_10958);
or U11447 (N_11447,N_10952,N_10502);
nor U11448 (N_11448,N_10810,N_10759);
xor U11449 (N_11449,N_10647,N_10636);
xnor U11450 (N_11450,N_10657,N_10730);
nor U11451 (N_11451,N_10771,N_10977);
xor U11452 (N_11452,N_10541,N_10601);
xnor U11453 (N_11453,N_10812,N_10696);
and U11454 (N_11454,N_10667,N_10628);
nand U11455 (N_11455,N_10574,N_10974);
xor U11456 (N_11456,N_10546,N_10890);
or U11457 (N_11457,N_10728,N_10594);
or U11458 (N_11458,N_10852,N_10750);
nand U11459 (N_11459,N_10519,N_10586);
xor U11460 (N_11460,N_10736,N_10799);
or U11461 (N_11461,N_10502,N_10761);
or U11462 (N_11462,N_10774,N_10788);
and U11463 (N_11463,N_10929,N_10812);
or U11464 (N_11464,N_10841,N_10746);
nor U11465 (N_11465,N_10879,N_10577);
xor U11466 (N_11466,N_10821,N_10872);
nand U11467 (N_11467,N_10828,N_10632);
and U11468 (N_11468,N_10843,N_10632);
and U11469 (N_11469,N_10650,N_10817);
or U11470 (N_11470,N_10777,N_10707);
xnor U11471 (N_11471,N_10978,N_10628);
or U11472 (N_11472,N_10698,N_10729);
or U11473 (N_11473,N_10741,N_10881);
and U11474 (N_11474,N_10930,N_10624);
nand U11475 (N_11475,N_10879,N_10992);
and U11476 (N_11476,N_10583,N_10724);
or U11477 (N_11477,N_10510,N_10936);
xnor U11478 (N_11478,N_10748,N_10506);
xnor U11479 (N_11479,N_10838,N_10643);
or U11480 (N_11480,N_10904,N_10531);
or U11481 (N_11481,N_10742,N_10955);
and U11482 (N_11482,N_10950,N_10607);
and U11483 (N_11483,N_10904,N_10706);
and U11484 (N_11484,N_10626,N_10776);
xnor U11485 (N_11485,N_10645,N_10603);
nor U11486 (N_11486,N_10760,N_10579);
xor U11487 (N_11487,N_10827,N_10960);
and U11488 (N_11488,N_10735,N_10551);
or U11489 (N_11489,N_10695,N_10832);
or U11490 (N_11490,N_10777,N_10811);
and U11491 (N_11491,N_10556,N_10579);
nor U11492 (N_11492,N_10754,N_10549);
nand U11493 (N_11493,N_10601,N_10676);
and U11494 (N_11494,N_10740,N_10716);
and U11495 (N_11495,N_10516,N_10729);
nor U11496 (N_11496,N_10821,N_10542);
xor U11497 (N_11497,N_10589,N_10834);
xor U11498 (N_11498,N_10542,N_10903);
or U11499 (N_11499,N_10610,N_10759);
or U11500 (N_11500,N_11413,N_11231);
or U11501 (N_11501,N_11182,N_11443);
and U11502 (N_11502,N_11077,N_11199);
or U11503 (N_11503,N_11282,N_11125);
xnor U11504 (N_11504,N_11131,N_11300);
or U11505 (N_11505,N_11441,N_11083);
nand U11506 (N_11506,N_11098,N_11190);
or U11507 (N_11507,N_11252,N_11240);
and U11508 (N_11508,N_11337,N_11053);
nor U11509 (N_11509,N_11010,N_11449);
nor U11510 (N_11510,N_11151,N_11273);
nand U11511 (N_11511,N_11408,N_11072);
xor U11512 (N_11512,N_11212,N_11029);
nand U11513 (N_11513,N_11488,N_11444);
nor U11514 (N_11514,N_11426,N_11401);
xnor U11515 (N_11515,N_11019,N_11291);
and U11516 (N_11516,N_11179,N_11299);
nand U11517 (N_11517,N_11255,N_11156);
xor U11518 (N_11518,N_11082,N_11165);
nor U11519 (N_11519,N_11430,N_11411);
xnor U11520 (N_11520,N_11431,N_11372);
and U11521 (N_11521,N_11063,N_11415);
xnor U11522 (N_11522,N_11085,N_11234);
nand U11523 (N_11523,N_11472,N_11219);
nor U11524 (N_11524,N_11475,N_11119);
or U11525 (N_11525,N_11429,N_11128);
and U11526 (N_11526,N_11287,N_11464);
xnor U11527 (N_11527,N_11086,N_11316);
xor U11528 (N_11528,N_11097,N_11324);
or U11529 (N_11529,N_11249,N_11172);
nand U11530 (N_11530,N_11256,N_11008);
and U11531 (N_11531,N_11467,N_11440);
and U11532 (N_11532,N_11268,N_11006);
nand U11533 (N_11533,N_11170,N_11201);
xor U11534 (N_11534,N_11414,N_11496);
and U11535 (N_11535,N_11056,N_11232);
nand U11536 (N_11536,N_11196,N_11129);
or U11537 (N_11537,N_11402,N_11395);
and U11538 (N_11538,N_11452,N_11007);
nand U11539 (N_11539,N_11253,N_11225);
nand U11540 (N_11540,N_11359,N_11205);
xor U11541 (N_11541,N_11152,N_11099);
nand U11542 (N_11542,N_11073,N_11090);
nor U11543 (N_11543,N_11051,N_11117);
nor U11544 (N_11544,N_11378,N_11434);
nand U11545 (N_11545,N_11314,N_11033);
nor U11546 (N_11546,N_11121,N_11484);
or U11547 (N_11547,N_11347,N_11070);
or U11548 (N_11548,N_11294,N_11003);
nand U11549 (N_11549,N_11360,N_11290);
nand U11550 (N_11550,N_11220,N_11318);
nand U11551 (N_11551,N_11242,N_11223);
nand U11552 (N_11552,N_11320,N_11143);
xnor U11553 (N_11553,N_11329,N_11214);
or U11554 (N_11554,N_11343,N_11032);
nor U11555 (N_11555,N_11495,N_11226);
nand U11556 (N_11556,N_11028,N_11306);
nor U11557 (N_11557,N_11215,N_11004);
xor U11558 (N_11558,N_11042,N_11340);
nor U11559 (N_11559,N_11124,N_11177);
nand U11560 (N_11560,N_11130,N_11014);
xor U11561 (N_11561,N_11394,N_11439);
and U11562 (N_11562,N_11396,N_11139);
nand U11563 (N_11563,N_11350,N_11382);
nor U11564 (N_11564,N_11308,N_11147);
xnor U11565 (N_11565,N_11038,N_11067);
nand U11566 (N_11566,N_11096,N_11322);
xor U11567 (N_11567,N_11238,N_11450);
nor U11568 (N_11568,N_11491,N_11262);
and U11569 (N_11569,N_11061,N_11364);
nand U11570 (N_11570,N_11154,N_11188);
nor U11571 (N_11571,N_11257,N_11247);
and U11572 (N_11572,N_11466,N_11417);
or U11573 (N_11573,N_11208,N_11494);
xnor U11574 (N_11574,N_11167,N_11245);
or U11575 (N_11575,N_11492,N_11421);
nor U11576 (N_11576,N_11323,N_11315);
and U11577 (N_11577,N_11277,N_11481);
nand U11578 (N_11578,N_11144,N_11246);
or U11579 (N_11579,N_11134,N_11221);
nand U11580 (N_11580,N_11462,N_11175);
nor U11581 (N_11581,N_11046,N_11305);
and U11582 (N_11582,N_11451,N_11103);
or U11583 (N_11583,N_11206,N_11002);
nand U11584 (N_11584,N_11391,N_11023);
nand U11585 (N_11585,N_11039,N_11260);
nor U11586 (N_11586,N_11250,N_11123);
nand U11587 (N_11587,N_11013,N_11370);
or U11588 (N_11588,N_11222,N_11112);
or U11589 (N_11589,N_11153,N_11357);
or U11590 (N_11590,N_11338,N_11362);
nand U11591 (N_11591,N_11478,N_11163);
and U11592 (N_11592,N_11258,N_11158);
xor U11593 (N_11593,N_11110,N_11118);
and U11594 (N_11594,N_11410,N_11365);
xor U11595 (N_11595,N_11375,N_11381);
and U11596 (N_11596,N_11319,N_11171);
or U11597 (N_11597,N_11024,N_11368);
or U11598 (N_11598,N_11376,N_11000);
nor U11599 (N_11599,N_11034,N_11482);
xnor U11600 (N_11600,N_11457,N_11025);
xor U11601 (N_11601,N_11267,N_11302);
or U11602 (N_11602,N_11180,N_11487);
and U11603 (N_11603,N_11336,N_11239);
nand U11604 (N_11604,N_11204,N_11465);
or U11605 (N_11605,N_11248,N_11122);
or U11606 (N_11606,N_11168,N_11137);
or U11607 (N_11607,N_11266,N_11095);
or U11608 (N_11608,N_11062,N_11344);
xor U11609 (N_11609,N_11427,N_11058);
xor U11610 (N_11610,N_11132,N_11379);
nor U11611 (N_11611,N_11271,N_11387);
and U11612 (N_11612,N_11334,N_11016);
nor U11613 (N_11613,N_11373,N_11052);
and U11614 (N_11614,N_11388,N_11279);
and U11615 (N_11615,N_11263,N_11017);
xnor U11616 (N_11616,N_11176,N_11454);
or U11617 (N_11617,N_11192,N_11209);
nor U11618 (N_11618,N_11397,N_11133);
nor U11619 (N_11619,N_11497,N_11183);
nand U11620 (N_11620,N_11037,N_11020);
or U11621 (N_11621,N_11107,N_11127);
or U11622 (N_11622,N_11331,N_11348);
xnor U11623 (N_11623,N_11217,N_11284);
nand U11624 (N_11624,N_11385,N_11342);
nor U11625 (N_11625,N_11384,N_11297);
or U11626 (N_11626,N_11445,N_11159);
or U11627 (N_11627,N_11393,N_11044);
nor U11628 (N_11628,N_11270,N_11328);
nor U11629 (N_11629,N_11311,N_11489);
xnor U11630 (N_11630,N_11265,N_11114);
or U11631 (N_11631,N_11374,N_11480);
nand U11632 (N_11632,N_11102,N_11354);
and U11633 (N_11633,N_11309,N_11022);
nand U11634 (N_11634,N_11335,N_11295);
and U11635 (N_11635,N_11474,N_11424);
or U11636 (N_11636,N_11218,N_11207);
xor U11637 (N_11637,N_11483,N_11035);
and U11638 (N_11638,N_11050,N_11304);
or U11639 (N_11639,N_11288,N_11150);
and U11640 (N_11640,N_11093,N_11437);
or U11641 (N_11641,N_11195,N_11326);
xnor U11642 (N_11642,N_11422,N_11446);
and U11643 (N_11643,N_11088,N_11135);
xnor U11644 (N_11644,N_11054,N_11198);
nor U11645 (N_11645,N_11109,N_11399);
nor U11646 (N_11646,N_11043,N_11071);
xor U11647 (N_11647,N_11155,N_11169);
xor U11648 (N_11648,N_11210,N_11213);
nor U11649 (N_11649,N_11278,N_11485);
or U11650 (N_11650,N_11100,N_11400);
xor U11651 (N_11651,N_11479,N_11241);
nand U11652 (N_11652,N_11303,N_11420);
xor U11653 (N_11653,N_11161,N_11460);
and U11654 (N_11654,N_11301,N_11065);
nor U11655 (N_11655,N_11386,N_11442);
or U11656 (N_11656,N_11140,N_11490);
nand U11657 (N_11657,N_11283,N_11423);
xnor U11658 (N_11658,N_11499,N_11453);
nand U11659 (N_11659,N_11031,N_11363);
and U11660 (N_11660,N_11371,N_11459);
or U11661 (N_11661,N_11259,N_11406);
and U11662 (N_11662,N_11435,N_11009);
nand U11663 (N_11663,N_11293,N_11055);
and U11664 (N_11664,N_11047,N_11361);
nand U11665 (N_11665,N_11470,N_11191);
and U11666 (N_11666,N_11064,N_11321);
xnor U11667 (N_11667,N_11264,N_11473);
and U11668 (N_11668,N_11261,N_11493);
xnor U11669 (N_11669,N_11157,N_11298);
xnor U11670 (N_11670,N_11230,N_11074);
nand U11671 (N_11671,N_11145,N_11274);
or U11672 (N_11672,N_11419,N_11356);
nand U11673 (N_11673,N_11280,N_11236);
and U11674 (N_11674,N_11228,N_11332);
and U11675 (N_11675,N_11148,N_11200);
xnor U11676 (N_11676,N_11164,N_11469);
or U11677 (N_11677,N_11463,N_11005);
xor U11678 (N_11678,N_11289,N_11233);
nand U11679 (N_11679,N_11281,N_11369);
and U11680 (N_11680,N_11352,N_11447);
nand U11681 (N_11681,N_11015,N_11269);
nor U11682 (N_11682,N_11398,N_11091);
nor U11683 (N_11683,N_11227,N_11078);
nand U11684 (N_11684,N_11377,N_11272);
and U11685 (N_11685,N_11276,N_11011);
and U11686 (N_11686,N_11349,N_11184);
or U11687 (N_11687,N_11229,N_11040);
and U11688 (N_11688,N_11068,N_11194);
nor U11689 (N_11689,N_11346,N_11433);
xnor U11690 (N_11690,N_11407,N_11076);
or U11691 (N_11691,N_11057,N_11313);
or U11692 (N_11692,N_11045,N_11160);
nand U11693 (N_11693,N_11254,N_11136);
or U11694 (N_11694,N_11066,N_11428);
nand U11695 (N_11695,N_11084,N_11089);
or U11696 (N_11696,N_11185,N_11237);
nor U11697 (N_11697,N_11060,N_11243);
nand U11698 (N_11698,N_11235,N_11436);
or U11699 (N_11699,N_11358,N_11366);
and U11700 (N_11700,N_11341,N_11286);
and U11701 (N_11701,N_11432,N_11059);
and U11702 (N_11702,N_11351,N_11456);
nor U11703 (N_11703,N_11081,N_11468);
nor U11704 (N_11704,N_11380,N_11115);
nand U11705 (N_11705,N_11036,N_11126);
or U11706 (N_11706,N_11080,N_11244);
and U11707 (N_11707,N_11404,N_11310);
or U11708 (N_11708,N_11193,N_11189);
or U11709 (N_11709,N_11498,N_11425);
nand U11710 (N_11710,N_11355,N_11146);
nand U11711 (N_11711,N_11187,N_11307);
or U11712 (N_11712,N_11292,N_11075);
and U11713 (N_11713,N_11048,N_11138);
nor U11714 (N_11714,N_11105,N_11416);
xor U11715 (N_11715,N_11116,N_11026);
and U11716 (N_11716,N_11409,N_11027);
and U11717 (N_11717,N_11471,N_11149);
or U11718 (N_11718,N_11461,N_11021);
or U11719 (N_11719,N_11285,N_11216);
nor U11720 (N_11720,N_11173,N_11477);
and U11721 (N_11721,N_11092,N_11012);
nand U11722 (N_11722,N_11383,N_11101);
nand U11723 (N_11723,N_11141,N_11162);
and U11724 (N_11724,N_11486,N_11251);
or U11725 (N_11725,N_11403,N_11390);
or U11726 (N_11726,N_11296,N_11211);
or U11727 (N_11727,N_11069,N_11030);
or U11728 (N_11728,N_11087,N_11018);
xor U11729 (N_11729,N_11094,N_11106);
xor U11730 (N_11730,N_11104,N_11108);
or U11731 (N_11731,N_11476,N_11049);
nand U11732 (N_11732,N_11202,N_11203);
or U11733 (N_11733,N_11275,N_11120);
or U11734 (N_11734,N_11330,N_11186);
xnor U11735 (N_11735,N_11367,N_11166);
and U11736 (N_11736,N_11181,N_11041);
nand U11737 (N_11737,N_11333,N_11001);
nor U11738 (N_11738,N_11448,N_11455);
nand U11739 (N_11739,N_11113,N_11412);
nand U11740 (N_11740,N_11405,N_11142);
and U11741 (N_11741,N_11325,N_11312);
nor U11742 (N_11742,N_11111,N_11389);
nand U11743 (N_11743,N_11197,N_11317);
nor U11744 (N_11744,N_11345,N_11458);
or U11745 (N_11745,N_11327,N_11339);
nand U11746 (N_11746,N_11224,N_11174);
and U11747 (N_11747,N_11079,N_11178);
and U11748 (N_11748,N_11418,N_11353);
and U11749 (N_11749,N_11392,N_11438);
nor U11750 (N_11750,N_11242,N_11439);
xnor U11751 (N_11751,N_11301,N_11047);
nand U11752 (N_11752,N_11304,N_11031);
nand U11753 (N_11753,N_11334,N_11095);
and U11754 (N_11754,N_11244,N_11312);
or U11755 (N_11755,N_11114,N_11450);
xor U11756 (N_11756,N_11130,N_11320);
nand U11757 (N_11757,N_11324,N_11130);
and U11758 (N_11758,N_11242,N_11361);
xnor U11759 (N_11759,N_11008,N_11311);
xnor U11760 (N_11760,N_11316,N_11466);
or U11761 (N_11761,N_11346,N_11133);
nor U11762 (N_11762,N_11496,N_11294);
xnor U11763 (N_11763,N_11432,N_11117);
or U11764 (N_11764,N_11188,N_11305);
or U11765 (N_11765,N_11378,N_11373);
and U11766 (N_11766,N_11287,N_11050);
nand U11767 (N_11767,N_11422,N_11121);
nand U11768 (N_11768,N_11220,N_11489);
or U11769 (N_11769,N_11447,N_11331);
nand U11770 (N_11770,N_11306,N_11006);
and U11771 (N_11771,N_11067,N_11317);
nor U11772 (N_11772,N_11402,N_11008);
xnor U11773 (N_11773,N_11313,N_11007);
nand U11774 (N_11774,N_11031,N_11276);
nand U11775 (N_11775,N_11338,N_11241);
or U11776 (N_11776,N_11423,N_11150);
and U11777 (N_11777,N_11107,N_11288);
and U11778 (N_11778,N_11464,N_11129);
nor U11779 (N_11779,N_11435,N_11268);
or U11780 (N_11780,N_11345,N_11065);
nor U11781 (N_11781,N_11390,N_11274);
nor U11782 (N_11782,N_11338,N_11191);
xor U11783 (N_11783,N_11108,N_11470);
nor U11784 (N_11784,N_11077,N_11094);
or U11785 (N_11785,N_11059,N_11258);
or U11786 (N_11786,N_11033,N_11016);
xnor U11787 (N_11787,N_11200,N_11085);
nand U11788 (N_11788,N_11125,N_11223);
and U11789 (N_11789,N_11181,N_11142);
nor U11790 (N_11790,N_11435,N_11397);
or U11791 (N_11791,N_11242,N_11093);
and U11792 (N_11792,N_11431,N_11025);
xor U11793 (N_11793,N_11132,N_11004);
and U11794 (N_11794,N_11369,N_11490);
nand U11795 (N_11795,N_11321,N_11447);
xnor U11796 (N_11796,N_11142,N_11449);
and U11797 (N_11797,N_11408,N_11105);
xnor U11798 (N_11798,N_11241,N_11170);
xor U11799 (N_11799,N_11311,N_11325);
nor U11800 (N_11800,N_11196,N_11233);
nor U11801 (N_11801,N_11324,N_11406);
nand U11802 (N_11802,N_11101,N_11140);
nor U11803 (N_11803,N_11396,N_11218);
nor U11804 (N_11804,N_11462,N_11130);
nor U11805 (N_11805,N_11398,N_11347);
and U11806 (N_11806,N_11296,N_11074);
or U11807 (N_11807,N_11102,N_11179);
nand U11808 (N_11808,N_11498,N_11028);
and U11809 (N_11809,N_11154,N_11279);
nor U11810 (N_11810,N_11241,N_11156);
and U11811 (N_11811,N_11337,N_11206);
and U11812 (N_11812,N_11105,N_11099);
nor U11813 (N_11813,N_11277,N_11148);
nor U11814 (N_11814,N_11187,N_11381);
and U11815 (N_11815,N_11492,N_11255);
and U11816 (N_11816,N_11349,N_11464);
and U11817 (N_11817,N_11173,N_11175);
nor U11818 (N_11818,N_11145,N_11487);
nor U11819 (N_11819,N_11437,N_11481);
and U11820 (N_11820,N_11495,N_11407);
xnor U11821 (N_11821,N_11002,N_11465);
or U11822 (N_11822,N_11070,N_11256);
xor U11823 (N_11823,N_11245,N_11138);
and U11824 (N_11824,N_11183,N_11108);
xor U11825 (N_11825,N_11255,N_11480);
nand U11826 (N_11826,N_11310,N_11289);
nand U11827 (N_11827,N_11039,N_11366);
or U11828 (N_11828,N_11136,N_11135);
xor U11829 (N_11829,N_11031,N_11253);
nand U11830 (N_11830,N_11084,N_11383);
nor U11831 (N_11831,N_11295,N_11080);
and U11832 (N_11832,N_11386,N_11014);
and U11833 (N_11833,N_11175,N_11193);
or U11834 (N_11834,N_11302,N_11115);
nor U11835 (N_11835,N_11292,N_11363);
and U11836 (N_11836,N_11226,N_11282);
and U11837 (N_11837,N_11285,N_11015);
nand U11838 (N_11838,N_11492,N_11038);
xnor U11839 (N_11839,N_11171,N_11482);
and U11840 (N_11840,N_11009,N_11200);
or U11841 (N_11841,N_11088,N_11175);
and U11842 (N_11842,N_11151,N_11021);
nor U11843 (N_11843,N_11082,N_11094);
xor U11844 (N_11844,N_11424,N_11369);
nor U11845 (N_11845,N_11443,N_11375);
xnor U11846 (N_11846,N_11372,N_11335);
or U11847 (N_11847,N_11489,N_11219);
nor U11848 (N_11848,N_11370,N_11006);
nand U11849 (N_11849,N_11352,N_11410);
nand U11850 (N_11850,N_11354,N_11389);
xor U11851 (N_11851,N_11477,N_11022);
and U11852 (N_11852,N_11061,N_11178);
and U11853 (N_11853,N_11466,N_11184);
and U11854 (N_11854,N_11356,N_11285);
nor U11855 (N_11855,N_11044,N_11145);
nand U11856 (N_11856,N_11043,N_11098);
xor U11857 (N_11857,N_11125,N_11140);
xnor U11858 (N_11858,N_11278,N_11100);
nor U11859 (N_11859,N_11183,N_11285);
nor U11860 (N_11860,N_11227,N_11342);
nor U11861 (N_11861,N_11030,N_11088);
nand U11862 (N_11862,N_11257,N_11250);
or U11863 (N_11863,N_11434,N_11387);
and U11864 (N_11864,N_11015,N_11305);
nand U11865 (N_11865,N_11237,N_11230);
or U11866 (N_11866,N_11140,N_11433);
or U11867 (N_11867,N_11100,N_11187);
xnor U11868 (N_11868,N_11036,N_11236);
nand U11869 (N_11869,N_11335,N_11029);
nand U11870 (N_11870,N_11041,N_11390);
nand U11871 (N_11871,N_11227,N_11176);
or U11872 (N_11872,N_11422,N_11099);
and U11873 (N_11873,N_11108,N_11242);
and U11874 (N_11874,N_11342,N_11180);
and U11875 (N_11875,N_11118,N_11281);
xnor U11876 (N_11876,N_11293,N_11406);
or U11877 (N_11877,N_11479,N_11414);
xor U11878 (N_11878,N_11200,N_11248);
or U11879 (N_11879,N_11065,N_11077);
nor U11880 (N_11880,N_11358,N_11388);
nor U11881 (N_11881,N_11267,N_11310);
nand U11882 (N_11882,N_11391,N_11398);
nor U11883 (N_11883,N_11448,N_11255);
nand U11884 (N_11884,N_11489,N_11454);
and U11885 (N_11885,N_11318,N_11143);
or U11886 (N_11886,N_11081,N_11129);
nand U11887 (N_11887,N_11368,N_11192);
and U11888 (N_11888,N_11234,N_11344);
xnor U11889 (N_11889,N_11173,N_11028);
or U11890 (N_11890,N_11383,N_11440);
xnor U11891 (N_11891,N_11184,N_11268);
nor U11892 (N_11892,N_11476,N_11069);
nor U11893 (N_11893,N_11251,N_11343);
nand U11894 (N_11894,N_11275,N_11309);
nor U11895 (N_11895,N_11201,N_11066);
xor U11896 (N_11896,N_11105,N_11253);
xor U11897 (N_11897,N_11157,N_11079);
xnor U11898 (N_11898,N_11228,N_11174);
nand U11899 (N_11899,N_11436,N_11295);
xor U11900 (N_11900,N_11091,N_11067);
and U11901 (N_11901,N_11013,N_11161);
and U11902 (N_11902,N_11445,N_11348);
and U11903 (N_11903,N_11200,N_11464);
or U11904 (N_11904,N_11058,N_11223);
nor U11905 (N_11905,N_11104,N_11176);
or U11906 (N_11906,N_11170,N_11388);
or U11907 (N_11907,N_11113,N_11112);
nor U11908 (N_11908,N_11193,N_11240);
xor U11909 (N_11909,N_11202,N_11299);
nand U11910 (N_11910,N_11488,N_11450);
nand U11911 (N_11911,N_11450,N_11185);
and U11912 (N_11912,N_11282,N_11097);
or U11913 (N_11913,N_11209,N_11007);
nor U11914 (N_11914,N_11138,N_11094);
xor U11915 (N_11915,N_11003,N_11070);
and U11916 (N_11916,N_11072,N_11080);
or U11917 (N_11917,N_11128,N_11065);
and U11918 (N_11918,N_11348,N_11166);
and U11919 (N_11919,N_11261,N_11365);
nand U11920 (N_11920,N_11325,N_11027);
xor U11921 (N_11921,N_11380,N_11417);
nand U11922 (N_11922,N_11305,N_11428);
or U11923 (N_11923,N_11074,N_11121);
nor U11924 (N_11924,N_11414,N_11083);
or U11925 (N_11925,N_11106,N_11172);
xor U11926 (N_11926,N_11092,N_11044);
and U11927 (N_11927,N_11490,N_11325);
nor U11928 (N_11928,N_11316,N_11246);
or U11929 (N_11929,N_11415,N_11279);
and U11930 (N_11930,N_11482,N_11033);
and U11931 (N_11931,N_11174,N_11153);
xor U11932 (N_11932,N_11334,N_11378);
and U11933 (N_11933,N_11333,N_11261);
xor U11934 (N_11934,N_11400,N_11073);
or U11935 (N_11935,N_11481,N_11463);
and U11936 (N_11936,N_11128,N_11074);
and U11937 (N_11937,N_11108,N_11487);
and U11938 (N_11938,N_11024,N_11121);
or U11939 (N_11939,N_11126,N_11186);
or U11940 (N_11940,N_11056,N_11202);
nor U11941 (N_11941,N_11398,N_11258);
and U11942 (N_11942,N_11307,N_11091);
nand U11943 (N_11943,N_11167,N_11165);
nand U11944 (N_11944,N_11213,N_11007);
nor U11945 (N_11945,N_11274,N_11317);
xnor U11946 (N_11946,N_11245,N_11436);
nand U11947 (N_11947,N_11415,N_11057);
nor U11948 (N_11948,N_11429,N_11332);
and U11949 (N_11949,N_11020,N_11411);
or U11950 (N_11950,N_11481,N_11216);
or U11951 (N_11951,N_11391,N_11264);
xnor U11952 (N_11952,N_11052,N_11172);
xor U11953 (N_11953,N_11228,N_11159);
xnor U11954 (N_11954,N_11241,N_11222);
xnor U11955 (N_11955,N_11416,N_11287);
nor U11956 (N_11956,N_11346,N_11183);
and U11957 (N_11957,N_11283,N_11198);
xnor U11958 (N_11958,N_11189,N_11155);
xor U11959 (N_11959,N_11443,N_11278);
nand U11960 (N_11960,N_11292,N_11255);
xor U11961 (N_11961,N_11078,N_11497);
and U11962 (N_11962,N_11047,N_11206);
nor U11963 (N_11963,N_11390,N_11211);
and U11964 (N_11964,N_11227,N_11424);
or U11965 (N_11965,N_11379,N_11463);
xnor U11966 (N_11966,N_11228,N_11149);
nand U11967 (N_11967,N_11231,N_11303);
nor U11968 (N_11968,N_11036,N_11074);
nand U11969 (N_11969,N_11437,N_11012);
and U11970 (N_11970,N_11075,N_11259);
nand U11971 (N_11971,N_11214,N_11016);
and U11972 (N_11972,N_11246,N_11189);
xor U11973 (N_11973,N_11213,N_11019);
xor U11974 (N_11974,N_11055,N_11359);
and U11975 (N_11975,N_11199,N_11436);
nor U11976 (N_11976,N_11122,N_11135);
or U11977 (N_11977,N_11053,N_11174);
nor U11978 (N_11978,N_11411,N_11170);
and U11979 (N_11979,N_11184,N_11357);
and U11980 (N_11980,N_11376,N_11176);
nand U11981 (N_11981,N_11324,N_11176);
nand U11982 (N_11982,N_11384,N_11043);
and U11983 (N_11983,N_11369,N_11218);
xnor U11984 (N_11984,N_11284,N_11242);
nand U11985 (N_11985,N_11263,N_11130);
nor U11986 (N_11986,N_11490,N_11287);
and U11987 (N_11987,N_11490,N_11303);
and U11988 (N_11988,N_11383,N_11405);
and U11989 (N_11989,N_11294,N_11111);
xor U11990 (N_11990,N_11489,N_11298);
and U11991 (N_11991,N_11260,N_11187);
or U11992 (N_11992,N_11430,N_11190);
or U11993 (N_11993,N_11159,N_11160);
nor U11994 (N_11994,N_11244,N_11220);
nand U11995 (N_11995,N_11052,N_11069);
nand U11996 (N_11996,N_11123,N_11223);
nand U11997 (N_11997,N_11012,N_11412);
xnor U11998 (N_11998,N_11298,N_11240);
and U11999 (N_11999,N_11204,N_11196);
xor U12000 (N_12000,N_11534,N_11978);
nand U12001 (N_12001,N_11602,N_11531);
nand U12002 (N_12002,N_11655,N_11692);
nor U12003 (N_12003,N_11689,N_11881);
and U12004 (N_12004,N_11902,N_11817);
or U12005 (N_12005,N_11972,N_11776);
or U12006 (N_12006,N_11653,N_11539);
and U12007 (N_12007,N_11894,N_11740);
and U12008 (N_12008,N_11821,N_11901);
xor U12009 (N_12009,N_11751,N_11535);
nand U12010 (N_12010,N_11651,N_11828);
nor U12011 (N_12011,N_11861,N_11605);
nand U12012 (N_12012,N_11918,N_11814);
and U12013 (N_12013,N_11779,N_11830);
and U12014 (N_12014,N_11772,N_11594);
nand U12015 (N_12015,N_11648,N_11850);
or U12016 (N_12016,N_11860,N_11573);
nor U12017 (N_12017,N_11611,N_11741);
xnor U12018 (N_12018,N_11796,N_11862);
and U12019 (N_12019,N_11865,N_11792);
nor U12020 (N_12020,N_11701,N_11640);
nor U12021 (N_12021,N_11513,N_11922);
or U12022 (N_12022,N_11987,N_11647);
nand U12023 (N_12023,N_11660,N_11630);
nor U12024 (N_12024,N_11909,N_11744);
xnor U12025 (N_12025,N_11777,N_11937);
and U12026 (N_12026,N_11743,N_11680);
or U12027 (N_12027,N_11912,N_11870);
xnor U12028 (N_12028,N_11957,N_11501);
nand U12029 (N_12029,N_11574,N_11599);
nor U12030 (N_12030,N_11628,N_11613);
nand U12031 (N_12031,N_11643,N_11770);
nor U12032 (N_12032,N_11703,N_11666);
or U12033 (N_12033,N_11866,N_11618);
and U12034 (N_12034,N_11920,N_11664);
or U12035 (N_12035,N_11771,N_11674);
nor U12036 (N_12036,N_11810,N_11632);
and U12037 (N_12037,N_11950,N_11644);
nand U12038 (N_12038,N_11548,N_11963);
or U12039 (N_12039,N_11911,N_11537);
and U12040 (N_12040,N_11614,N_11626);
and U12041 (N_12041,N_11587,N_11526);
and U12042 (N_12042,N_11724,N_11603);
or U12043 (N_12043,N_11543,N_11765);
nor U12044 (N_12044,N_11800,N_11585);
xnor U12045 (N_12045,N_11787,N_11714);
and U12046 (N_12046,N_11519,N_11915);
xor U12047 (N_12047,N_11803,N_11898);
or U12048 (N_12048,N_11849,N_11670);
xor U12049 (N_12049,N_11658,N_11790);
or U12050 (N_12050,N_11693,N_11500);
nand U12051 (N_12051,N_11899,N_11927);
xnor U12052 (N_12052,N_11712,N_11657);
nor U12053 (N_12053,N_11708,N_11782);
nor U12054 (N_12054,N_11876,N_11942);
or U12055 (N_12055,N_11859,N_11729);
and U12056 (N_12056,N_11941,N_11677);
and U12057 (N_12057,N_11928,N_11829);
and U12058 (N_12058,N_11565,N_11515);
and U12059 (N_12059,N_11561,N_11571);
nand U12060 (N_12060,N_11671,N_11590);
nand U12061 (N_12061,N_11930,N_11673);
or U12062 (N_12062,N_11725,N_11697);
nand U12063 (N_12063,N_11516,N_11900);
xor U12064 (N_12064,N_11699,N_11756);
and U12065 (N_12065,N_11806,N_11832);
xor U12066 (N_12066,N_11887,N_11749);
or U12067 (N_12067,N_11775,N_11544);
nor U12068 (N_12068,N_11807,N_11698);
and U12069 (N_12069,N_11781,N_11560);
nor U12070 (N_12070,N_11953,N_11757);
and U12071 (N_12071,N_11669,N_11508);
or U12072 (N_12072,N_11558,N_11654);
nor U12073 (N_12073,N_11623,N_11895);
or U12074 (N_12074,N_11931,N_11527);
nand U12075 (N_12075,N_11837,N_11667);
or U12076 (N_12076,N_11570,N_11562);
xnor U12077 (N_12077,N_11789,N_11715);
and U12078 (N_12078,N_11583,N_11956);
nor U12079 (N_12079,N_11816,N_11877);
and U12080 (N_12080,N_11596,N_11606);
and U12081 (N_12081,N_11636,N_11595);
nor U12082 (N_12082,N_11510,N_11801);
nor U12083 (N_12083,N_11733,N_11704);
and U12084 (N_12084,N_11533,N_11685);
and U12085 (N_12085,N_11718,N_11555);
or U12086 (N_12086,N_11524,N_11608);
and U12087 (N_12087,N_11879,N_11762);
xnor U12088 (N_12088,N_11886,N_11940);
and U12089 (N_12089,N_11855,N_11913);
nand U12090 (N_12090,N_11709,N_11766);
and U12091 (N_12091,N_11853,N_11642);
nor U12092 (N_12092,N_11661,N_11945);
and U12093 (N_12093,N_11995,N_11662);
nor U12094 (N_12094,N_11625,N_11580);
xnor U12095 (N_12095,N_11774,N_11788);
nand U12096 (N_12096,N_11503,N_11577);
nand U12097 (N_12097,N_11758,N_11916);
nand U12098 (N_12098,N_11960,N_11974);
nor U12099 (N_12099,N_11826,N_11554);
nor U12100 (N_12100,N_11885,N_11825);
or U12101 (N_12101,N_11946,N_11967);
xnor U12102 (N_12102,N_11764,N_11778);
and U12103 (N_12103,N_11668,N_11621);
nand U12104 (N_12104,N_11586,N_11867);
or U12105 (N_12105,N_11734,N_11710);
nor U12106 (N_12106,N_11523,N_11903);
nand U12107 (N_12107,N_11889,N_11564);
or U12108 (N_12108,N_11607,N_11917);
and U12109 (N_12109,N_11737,N_11869);
xnor U12110 (N_12110,N_11581,N_11791);
nor U12111 (N_12111,N_11858,N_11906);
xnor U12112 (N_12112,N_11511,N_11933);
or U12113 (N_12113,N_11617,N_11745);
or U12114 (N_12114,N_11522,N_11797);
or U12115 (N_12115,N_11811,N_11955);
and U12116 (N_12116,N_11530,N_11742);
and U12117 (N_12117,N_11904,N_11529);
xnor U12118 (N_12118,N_11846,N_11794);
or U12119 (N_12119,N_11804,N_11897);
nand U12120 (N_12120,N_11923,N_11965);
nand U12121 (N_12121,N_11702,N_11633);
nand U12122 (N_12122,N_11977,N_11629);
xor U12123 (N_12123,N_11656,N_11582);
or U12124 (N_12124,N_11851,N_11649);
nor U12125 (N_12125,N_11553,N_11994);
and U12126 (N_12126,N_11615,N_11549);
and U12127 (N_12127,N_11805,N_11694);
xor U12128 (N_12128,N_11721,N_11507);
nand U12129 (N_12129,N_11739,N_11952);
xnor U12130 (N_12130,N_11732,N_11844);
nor U12131 (N_12131,N_11505,N_11512);
nor U12132 (N_12132,N_11871,N_11888);
nor U12133 (N_12133,N_11892,N_11848);
or U12134 (N_12134,N_11998,N_11600);
or U12135 (N_12135,N_11525,N_11578);
nand U12136 (N_12136,N_11986,N_11641);
or U12137 (N_12137,N_11989,N_11637);
and U12138 (N_12138,N_11569,N_11818);
nand U12139 (N_12139,N_11834,N_11723);
xnor U12140 (N_12140,N_11619,N_11843);
nor U12141 (N_12141,N_11798,N_11682);
nor U12142 (N_12142,N_11552,N_11665);
nor U12143 (N_12143,N_11878,N_11517);
and U12144 (N_12144,N_11722,N_11925);
nand U12145 (N_12145,N_11767,N_11755);
and U12146 (N_12146,N_11890,N_11514);
xnor U12147 (N_12147,N_11983,N_11936);
nor U12148 (N_12148,N_11938,N_11891);
or U12149 (N_12149,N_11992,N_11975);
nor U12150 (N_12150,N_11520,N_11650);
nor U12151 (N_12151,N_11624,N_11842);
or U12152 (N_12152,N_11958,N_11935);
or U12153 (N_12153,N_11783,N_11822);
nor U12154 (N_12154,N_11968,N_11907);
and U12155 (N_12155,N_11696,N_11847);
xnor U12156 (N_12156,N_11663,N_11738);
or U12157 (N_12157,N_11584,N_11563);
nand U12158 (N_12158,N_11827,N_11747);
and U12159 (N_12159,N_11686,N_11597);
nand U12160 (N_12160,N_11924,N_11730);
xor U12161 (N_12161,N_11976,N_11536);
nor U12162 (N_12162,N_11831,N_11717);
or U12163 (N_12163,N_11746,N_11993);
nor U12164 (N_12164,N_11591,N_11979);
and U12165 (N_12165,N_11908,N_11845);
or U12166 (N_12166,N_11609,N_11990);
or U12167 (N_12167,N_11880,N_11559);
nor U12168 (N_12168,N_11864,N_11592);
nor U12169 (N_12169,N_11973,N_11954);
nand U12170 (N_12170,N_11679,N_11612);
nor U12171 (N_12171,N_11620,N_11598);
xor U12172 (N_12172,N_11785,N_11557);
or U12173 (N_12173,N_11688,N_11824);
nor U12174 (N_12174,N_11631,N_11705);
or U12175 (N_12175,N_11991,N_11735);
nand U12176 (N_12176,N_11627,N_11883);
nand U12177 (N_12177,N_11575,N_11921);
or U12178 (N_12178,N_11691,N_11638);
and U12179 (N_12179,N_11932,N_11761);
nor U12180 (N_12180,N_11835,N_11882);
nand U12181 (N_12181,N_11635,N_11506);
or U12182 (N_12182,N_11873,N_11984);
nor U12183 (N_12183,N_11893,N_11874);
nand U12184 (N_12184,N_11634,N_11546);
and U12185 (N_12185,N_11687,N_11645);
nor U12186 (N_12186,N_11566,N_11799);
nor U12187 (N_12187,N_11521,N_11815);
xnor U12188 (N_12188,N_11919,N_11706);
xnor U12189 (N_12189,N_11999,N_11840);
and U12190 (N_12190,N_11616,N_11969);
or U12191 (N_12191,N_11532,N_11572);
and U12192 (N_12192,N_11786,N_11528);
or U12193 (N_12193,N_11753,N_11910);
xnor U12194 (N_12194,N_11759,N_11985);
nand U12195 (N_12195,N_11659,N_11568);
or U12196 (N_12196,N_11711,N_11793);
nand U12197 (N_12197,N_11754,N_11872);
nor U12198 (N_12198,N_11676,N_11646);
xor U12199 (N_12199,N_11833,N_11726);
or U12200 (N_12200,N_11982,N_11716);
nand U12201 (N_12201,N_11678,N_11836);
nand U12202 (N_12202,N_11750,N_11854);
and U12203 (N_12203,N_11707,N_11601);
nand U12204 (N_12204,N_11929,N_11769);
nand U12205 (N_12205,N_11748,N_11545);
nand U12206 (N_12206,N_11784,N_11589);
nor U12207 (N_12207,N_11588,N_11823);
nand U12208 (N_12208,N_11948,N_11857);
nor U12209 (N_12209,N_11763,N_11542);
nand U12210 (N_12210,N_11970,N_11819);
or U12211 (N_12211,N_11947,N_11795);
and U12212 (N_12212,N_11971,N_11802);
nand U12213 (N_12213,N_11820,N_11684);
and U12214 (N_12214,N_11934,N_11719);
and U12215 (N_12215,N_11997,N_11868);
nor U12216 (N_12216,N_11593,N_11622);
or U12217 (N_12217,N_11841,N_11852);
and U12218 (N_12218,N_11905,N_11962);
xnor U12219 (N_12219,N_11856,N_11504);
nor U12220 (N_12220,N_11576,N_11926);
xnor U12221 (N_12221,N_11579,N_11780);
and U12222 (N_12222,N_11809,N_11736);
nand U12223 (N_12223,N_11540,N_11639);
xor U12224 (N_12224,N_11509,N_11713);
xor U12225 (N_12225,N_11556,N_11675);
nor U12226 (N_12226,N_11896,N_11550);
nand U12227 (N_12227,N_11812,N_11700);
and U12228 (N_12228,N_11695,N_11652);
or U12229 (N_12229,N_11551,N_11951);
nor U12230 (N_12230,N_11959,N_11502);
nand U12231 (N_12231,N_11728,N_11914);
or U12232 (N_12232,N_11720,N_11731);
and U12233 (N_12233,N_11839,N_11610);
xor U12234 (N_12234,N_11604,N_11567);
nand U12235 (N_12235,N_11988,N_11813);
xor U12236 (N_12236,N_11727,N_11838);
nor U12237 (N_12237,N_11768,N_11863);
or U12238 (N_12238,N_11541,N_11944);
nor U12239 (N_12239,N_11752,N_11884);
nand U12240 (N_12240,N_11808,N_11943);
nand U12241 (N_12241,N_11980,N_11690);
nand U12242 (N_12242,N_11773,N_11939);
xor U12243 (N_12243,N_11875,N_11547);
xnor U12244 (N_12244,N_11981,N_11538);
nand U12245 (N_12245,N_11760,N_11961);
nand U12246 (N_12246,N_11996,N_11518);
and U12247 (N_12247,N_11681,N_11672);
nor U12248 (N_12248,N_11964,N_11949);
nor U12249 (N_12249,N_11966,N_11683);
xnor U12250 (N_12250,N_11827,N_11784);
or U12251 (N_12251,N_11528,N_11518);
or U12252 (N_12252,N_11729,N_11913);
nand U12253 (N_12253,N_11627,N_11572);
or U12254 (N_12254,N_11906,N_11640);
xnor U12255 (N_12255,N_11586,N_11659);
and U12256 (N_12256,N_11650,N_11697);
nor U12257 (N_12257,N_11565,N_11794);
and U12258 (N_12258,N_11550,N_11820);
nor U12259 (N_12259,N_11948,N_11733);
xor U12260 (N_12260,N_11622,N_11532);
and U12261 (N_12261,N_11599,N_11994);
or U12262 (N_12262,N_11643,N_11601);
nor U12263 (N_12263,N_11921,N_11768);
and U12264 (N_12264,N_11524,N_11940);
and U12265 (N_12265,N_11612,N_11921);
and U12266 (N_12266,N_11878,N_11795);
xor U12267 (N_12267,N_11824,N_11832);
or U12268 (N_12268,N_11789,N_11831);
nor U12269 (N_12269,N_11627,N_11735);
xnor U12270 (N_12270,N_11928,N_11613);
nor U12271 (N_12271,N_11969,N_11953);
xor U12272 (N_12272,N_11633,N_11661);
and U12273 (N_12273,N_11968,N_11624);
and U12274 (N_12274,N_11654,N_11735);
or U12275 (N_12275,N_11562,N_11617);
nor U12276 (N_12276,N_11720,N_11836);
and U12277 (N_12277,N_11785,N_11600);
or U12278 (N_12278,N_11621,N_11704);
xor U12279 (N_12279,N_11860,N_11692);
xor U12280 (N_12280,N_11689,N_11568);
and U12281 (N_12281,N_11893,N_11752);
xnor U12282 (N_12282,N_11982,N_11504);
xor U12283 (N_12283,N_11915,N_11855);
and U12284 (N_12284,N_11668,N_11594);
nand U12285 (N_12285,N_11869,N_11618);
or U12286 (N_12286,N_11783,N_11517);
or U12287 (N_12287,N_11854,N_11681);
nor U12288 (N_12288,N_11560,N_11832);
xor U12289 (N_12289,N_11550,N_11629);
xor U12290 (N_12290,N_11744,N_11951);
nand U12291 (N_12291,N_11608,N_11673);
or U12292 (N_12292,N_11852,N_11929);
xnor U12293 (N_12293,N_11945,N_11834);
or U12294 (N_12294,N_11959,N_11739);
or U12295 (N_12295,N_11944,N_11514);
or U12296 (N_12296,N_11877,N_11697);
or U12297 (N_12297,N_11788,N_11840);
xor U12298 (N_12298,N_11860,N_11745);
nand U12299 (N_12299,N_11931,N_11971);
or U12300 (N_12300,N_11609,N_11974);
xnor U12301 (N_12301,N_11896,N_11723);
nand U12302 (N_12302,N_11743,N_11816);
nand U12303 (N_12303,N_11666,N_11745);
xor U12304 (N_12304,N_11921,N_11766);
or U12305 (N_12305,N_11654,N_11645);
nor U12306 (N_12306,N_11695,N_11931);
nand U12307 (N_12307,N_11779,N_11827);
and U12308 (N_12308,N_11883,N_11643);
nand U12309 (N_12309,N_11872,N_11822);
or U12310 (N_12310,N_11997,N_11772);
xnor U12311 (N_12311,N_11614,N_11710);
nand U12312 (N_12312,N_11975,N_11775);
and U12313 (N_12313,N_11972,N_11855);
or U12314 (N_12314,N_11844,N_11761);
xor U12315 (N_12315,N_11779,N_11782);
xor U12316 (N_12316,N_11734,N_11739);
nor U12317 (N_12317,N_11522,N_11831);
nand U12318 (N_12318,N_11720,N_11937);
nor U12319 (N_12319,N_11681,N_11824);
nand U12320 (N_12320,N_11646,N_11807);
or U12321 (N_12321,N_11737,N_11971);
nand U12322 (N_12322,N_11933,N_11540);
xnor U12323 (N_12323,N_11989,N_11830);
nand U12324 (N_12324,N_11831,N_11545);
and U12325 (N_12325,N_11831,N_11762);
and U12326 (N_12326,N_11974,N_11952);
or U12327 (N_12327,N_11829,N_11675);
xnor U12328 (N_12328,N_11548,N_11887);
or U12329 (N_12329,N_11726,N_11941);
or U12330 (N_12330,N_11586,N_11769);
nand U12331 (N_12331,N_11702,N_11559);
and U12332 (N_12332,N_11799,N_11913);
and U12333 (N_12333,N_11756,N_11762);
or U12334 (N_12334,N_11617,N_11583);
xor U12335 (N_12335,N_11617,N_11802);
nand U12336 (N_12336,N_11888,N_11621);
and U12337 (N_12337,N_11752,N_11640);
xor U12338 (N_12338,N_11939,N_11543);
nor U12339 (N_12339,N_11910,N_11714);
or U12340 (N_12340,N_11676,N_11741);
and U12341 (N_12341,N_11655,N_11827);
and U12342 (N_12342,N_11557,N_11537);
xor U12343 (N_12343,N_11660,N_11896);
or U12344 (N_12344,N_11622,N_11644);
nor U12345 (N_12345,N_11620,N_11523);
nand U12346 (N_12346,N_11677,N_11684);
xnor U12347 (N_12347,N_11968,N_11507);
xnor U12348 (N_12348,N_11633,N_11926);
or U12349 (N_12349,N_11752,N_11947);
and U12350 (N_12350,N_11925,N_11886);
and U12351 (N_12351,N_11728,N_11916);
and U12352 (N_12352,N_11617,N_11986);
xnor U12353 (N_12353,N_11686,N_11553);
or U12354 (N_12354,N_11817,N_11981);
or U12355 (N_12355,N_11838,N_11962);
and U12356 (N_12356,N_11738,N_11759);
xnor U12357 (N_12357,N_11584,N_11684);
nand U12358 (N_12358,N_11638,N_11987);
and U12359 (N_12359,N_11510,N_11530);
xor U12360 (N_12360,N_11998,N_11631);
xor U12361 (N_12361,N_11925,N_11732);
nor U12362 (N_12362,N_11953,N_11663);
or U12363 (N_12363,N_11867,N_11506);
nand U12364 (N_12364,N_11978,N_11646);
nand U12365 (N_12365,N_11953,N_11557);
nand U12366 (N_12366,N_11829,N_11506);
xor U12367 (N_12367,N_11598,N_11758);
and U12368 (N_12368,N_11867,N_11681);
xor U12369 (N_12369,N_11622,N_11549);
nand U12370 (N_12370,N_11975,N_11714);
nor U12371 (N_12371,N_11886,N_11572);
and U12372 (N_12372,N_11678,N_11662);
and U12373 (N_12373,N_11996,N_11813);
or U12374 (N_12374,N_11797,N_11770);
xor U12375 (N_12375,N_11783,N_11613);
and U12376 (N_12376,N_11768,N_11791);
or U12377 (N_12377,N_11604,N_11645);
or U12378 (N_12378,N_11515,N_11578);
and U12379 (N_12379,N_11517,N_11627);
or U12380 (N_12380,N_11904,N_11956);
or U12381 (N_12381,N_11794,N_11795);
nand U12382 (N_12382,N_11643,N_11667);
nor U12383 (N_12383,N_11673,N_11827);
xor U12384 (N_12384,N_11735,N_11561);
and U12385 (N_12385,N_11810,N_11733);
and U12386 (N_12386,N_11995,N_11910);
or U12387 (N_12387,N_11852,N_11993);
nor U12388 (N_12388,N_11986,N_11726);
nand U12389 (N_12389,N_11940,N_11955);
xor U12390 (N_12390,N_11937,N_11502);
nor U12391 (N_12391,N_11635,N_11565);
or U12392 (N_12392,N_11877,N_11808);
or U12393 (N_12393,N_11771,N_11997);
xnor U12394 (N_12394,N_11996,N_11736);
or U12395 (N_12395,N_11596,N_11844);
and U12396 (N_12396,N_11619,N_11805);
nand U12397 (N_12397,N_11771,N_11714);
nand U12398 (N_12398,N_11813,N_11825);
xor U12399 (N_12399,N_11951,N_11656);
nor U12400 (N_12400,N_11785,N_11694);
nand U12401 (N_12401,N_11885,N_11768);
and U12402 (N_12402,N_11522,N_11803);
nand U12403 (N_12403,N_11916,N_11823);
or U12404 (N_12404,N_11851,N_11985);
and U12405 (N_12405,N_11821,N_11598);
nand U12406 (N_12406,N_11711,N_11684);
or U12407 (N_12407,N_11631,N_11649);
nor U12408 (N_12408,N_11926,N_11947);
nand U12409 (N_12409,N_11772,N_11537);
or U12410 (N_12410,N_11799,N_11823);
or U12411 (N_12411,N_11709,N_11876);
nor U12412 (N_12412,N_11813,N_11886);
and U12413 (N_12413,N_11888,N_11803);
nand U12414 (N_12414,N_11961,N_11608);
nor U12415 (N_12415,N_11884,N_11799);
or U12416 (N_12416,N_11630,N_11615);
nor U12417 (N_12417,N_11792,N_11604);
nor U12418 (N_12418,N_11549,N_11656);
or U12419 (N_12419,N_11568,N_11502);
nand U12420 (N_12420,N_11523,N_11780);
and U12421 (N_12421,N_11939,N_11969);
nor U12422 (N_12422,N_11954,N_11747);
nand U12423 (N_12423,N_11512,N_11570);
or U12424 (N_12424,N_11965,N_11664);
or U12425 (N_12425,N_11648,N_11961);
nand U12426 (N_12426,N_11751,N_11937);
nand U12427 (N_12427,N_11883,N_11994);
and U12428 (N_12428,N_11733,N_11652);
or U12429 (N_12429,N_11970,N_11919);
xor U12430 (N_12430,N_11698,N_11696);
nand U12431 (N_12431,N_11642,N_11504);
nor U12432 (N_12432,N_11542,N_11565);
xor U12433 (N_12433,N_11861,N_11501);
nor U12434 (N_12434,N_11687,N_11677);
xor U12435 (N_12435,N_11654,N_11569);
nor U12436 (N_12436,N_11972,N_11518);
or U12437 (N_12437,N_11629,N_11945);
or U12438 (N_12438,N_11999,N_11972);
xnor U12439 (N_12439,N_11597,N_11987);
or U12440 (N_12440,N_11790,N_11594);
nor U12441 (N_12441,N_11709,N_11624);
and U12442 (N_12442,N_11935,N_11598);
or U12443 (N_12443,N_11668,N_11917);
nand U12444 (N_12444,N_11966,N_11656);
nand U12445 (N_12445,N_11548,N_11510);
nand U12446 (N_12446,N_11993,N_11637);
nand U12447 (N_12447,N_11746,N_11675);
nand U12448 (N_12448,N_11763,N_11734);
nor U12449 (N_12449,N_11849,N_11786);
and U12450 (N_12450,N_11678,N_11818);
and U12451 (N_12451,N_11772,N_11961);
nor U12452 (N_12452,N_11699,N_11655);
and U12453 (N_12453,N_11802,N_11676);
xnor U12454 (N_12454,N_11644,N_11884);
nor U12455 (N_12455,N_11515,N_11989);
nand U12456 (N_12456,N_11571,N_11604);
and U12457 (N_12457,N_11742,N_11574);
xnor U12458 (N_12458,N_11934,N_11647);
or U12459 (N_12459,N_11596,N_11531);
and U12460 (N_12460,N_11535,N_11654);
and U12461 (N_12461,N_11800,N_11735);
nand U12462 (N_12462,N_11960,N_11954);
nor U12463 (N_12463,N_11999,N_11681);
nand U12464 (N_12464,N_11749,N_11893);
nor U12465 (N_12465,N_11663,N_11908);
nand U12466 (N_12466,N_11865,N_11821);
and U12467 (N_12467,N_11944,N_11963);
xnor U12468 (N_12468,N_11988,N_11843);
and U12469 (N_12469,N_11693,N_11772);
and U12470 (N_12470,N_11766,N_11654);
and U12471 (N_12471,N_11857,N_11840);
nand U12472 (N_12472,N_11610,N_11712);
or U12473 (N_12473,N_11764,N_11540);
xor U12474 (N_12474,N_11844,N_11873);
nand U12475 (N_12475,N_11735,N_11881);
nor U12476 (N_12476,N_11954,N_11686);
nand U12477 (N_12477,N_11660,N_11934);
xor U12478 (N_12478,N_11701,N_11946);
xnor U12479 (N_12479,N_11684,N_11768);
xor U12480 (N_12480,N_11534,N_11639);
nor U12481 (N_12481,N_11536,N_11682);
nand U12482 (N_12482,N_11802,N_11728);
nand U12483 (N_12483,N_11549,N_11872);
nand U12484 (N_12484,N_11956,N_11969);
nor U12485 (N_12485,N_11924,N_11828);
xnor U12486 (N_12486,N_11803,N_11856);
nand U12487 (N_12487,N_11822,N_11888);
nand U12488 (N_12488,N_11722,N_11708);
and U12489 (N_12489,N_11971,N_11635);
or U12490 (N_12490,N_11620,N_11848);
xor U12491 (N_12491,N_11545,N_11812);
and U12492 (N_12492,N_11773,N_11966);
nor U12493 (N_12493,N_11563,N_11859);
nand U12494 (N_12494,N_11628,N_11869);
nor U12495 (N_12495,N_11551,N_11510);
and U12496 (N_12496,N_11610,N_11765);
xor U12497 (N_12497,N_11993,N_11783);
or U12498 (N_12498,N_11634,N_11858);
nand U12499 (N_12499,N_11519,N_11507);
xnor U12500 (N_12500,N_12172,N_12222);
nor U12501 (N_12501,N_12390,N_12422);
or U12502 (N_12502,N_12384,N_12306);
nor U12503 (N_12503,N_12182,N_12444);
nor U12504 (N_12504,N_12209,N_12161);
nand U12505 (N_12505,N_12063,N_12479);
or U12506 (N_12506,N_12120,N_12369);
nor U12507 (N_12507,N_12437,N_12453);
nor U12508 (N_12508,N_12070,N_12025);
or U12509 (N_12509,N_12155,N_12102);
xor U12510 (N_12510,N_12188,N_12143);
nor U12511 (N_12511,N_12213,N_12321);
or U12512 (N_12512,N_12354,N_12386);
and U12513 (N_12513,N_12225,N_12366);
xnor U12514 (N_12514,N_12158,N_12248);
and U12515 (N_12515,N_12428,N_12331);
or U12516 (N_12516,N_12226,N_12218);
nor U12517 (N_12517,N_12285,N_12455);
or U12518 (N_12518,N_12040,N_12307);
nand U12519 (N_12519,N_12026,N_12094);
xnor U12520 (N_12520,N_12295,N_12006);
nor U12521 (N_12521,N_12169,N_12097);
nand U12522 (N_12522,N_12326,N_12292);
nor U12523 (N_12523,N_12104,N_12033);
nor U12524 (N_12524,N_12170,N_12329);
nor U12525 (N_12525,N_12396,N_12121);
and U12526 (N_12526,N_12137,N_12374);
or U12527 (N_12527,N_12270,N_12375);
or U12528 (N_12528,N_12445,N_12136);
or U12529 (N_12529,N_12122,N_12334);
nand U12530 (N_12530,N_12397,N_12283);
nand U12531 (N_12531,N_12099,N_12024);
and U12532 (N_12532,N_12011,N_12254);
and U12533 (N_12533,N_12176,N_12426);
or U12534 (N_12534,N_12395,N_12340);
xor U12535 (N_12535,N_12410,N_12133);
nor U12536 (N_12536,N_12105,N_12239);
nand U12537 (N_12537,N_12081,N_12309);
nor U12538 (N_12538,N_12262,N_12421);
and U12539 (N_12539,N_12186,N_12019);
xor U12540 (N_12540,N_12048,N_12459);
nor U12541 (N_12541,N_12214,N_12058);
and U12542 (N_12542,N_12150,N_12145);
xor U12543 (N_12543,N_12039,N_12325);
and U12544 (N_12544,N_12371,N_12324);
and U12545 (N_12545,N_12373,N_12287);
and U12546 (N_12546,N_12378,N_12414);
and U12547 (N_12547,N_12101,N_12320);
nand U12548 (N_12548,N_12129,N_12469);
nand U12549 (N_12549,N_12247,N_12191);
nor U12550 (N_12550,N_12093,N_12416);
xor U12551 (N_12551,N_12352,N_12243);
or U12552 (N_12552,N_12002,N_12492);
xnor U12553 (N_12553,N_12330,N_12269);
nand U12554 (N_12554,N_12007,N_12448);
xnor U12555 (N_12555,N_12255,N_12431);
xnor U12556 (N_12556,N_12064,N_12071);
or U12557 (N_12557,N_12030,N_12227);
xor U12558 (N_12558,N_12480,N_12349);
nand U12559 (N_12559,N_12148,N_12245);
or U12560 (N_12560,N_12407,N_12317);
nand U12561 (N_12561,N_12302,N_12343);
xnor U12562 (N_12562,N_12275,N_12013);
and U12563 (N_12563,N_12242,N_12417);
and U12564 (N_12564,N_12429,N_12119);
nor U12565 (N_12565,N_12391,N_12196);
nor U12566 (N_12566,N_12228,N_12299);
or U12567 (N_12567,N_12041,N_12364);
nand U12568 (N_12568,N_12450,N_12207);
and U12569 (N_12569,N_12493,N_12438);
nor U12570 (N_12570,N_12362,N_12481);
xor U12571 (N_12571,N_12156,N_12141);
nand U12572 (N_12572,N_12100,N_12166);
xor U12573 (N_12573,N_12142,N_12047);
nand U12574 (N_12574,N_12003,N_12339);
nor U12575 (N_12575,N_12074,N_12181);
nor U12576 (N_12576,N_12035,N_12229);
and U12577 (N_12577,N_12260,N_12042);
and U12578 (N_12578,N_12452,N_12034);
and U12579 (N_12579,N_12173,N_12050);
xor U12580 (N_12580,N_12418,N_12303);
xnor U12581 (N_12581,N_12276,N_12393);
nor U12582 (N_12582,N_12473,N_12029);
nor U12583 (N_12583,N_12353,N_12211);
nand U12584 (N_12584,N_12338,N_12487);
or U12585 (N_12585,N_12112,N_12079);
nor U12586 (N_12586,N_12062,N_12435);
nor U12587 (N_12587,N_12043,N_12127);
xor U12588 (N_12588,N_12357,N_12082);
and U12589 (N_12589,N_12014,N_12387);
nor U12590 (N_12590,N_12089,N_12441);
nand U12591 (N_12591,N_12277,N_12389);
or U12592 (N_12592,N_12190,N_12356);
nor U12593 (N_12593,N_12092,N_12467);
or U12594 (N_12594,N_12446,N_12210);
or U12595 (N_12595,N_12472,N_12244);
nor U12596 (N_12596,N_12263,N_12365);
xnor U12597 (N_12597,N_12401,N_12151);
nand U12598 (N_12598,N_12208,N_12434);
nand U12599 (N_12599,N_12177,N_12332);
xor U12600 (N_12600,N_12337,N_12004);
xor U12601 (N_12601,N_12425,N_12164);
and U12602 (N_12602,N_12405,N_12404);
and U12603 (N_12603,N_12311,N_12318);
nand U12604 (N_12604,N_12126,N_12335);
nand U12605 (N_12605,N_12061,N_12179);
nand U12606 (N_12606,N_12187,N_12072);
or U12607 (N_12607,N_12496,N_12060);
and U12608 (N_12608,N_12456,N_12235);
or U12609 (N_12609,N_12465,N_12402);
or U12610 (N_12610,N_12403,N_12488);
nor U12611 (N_12611,N_12103,N_12221);
or U12612 (N_12612,N_12195,N_12291);
and U12613 (N_12613,N_12051,N_12268);
or U12614 (N_12614,N_12163,N_12123);
or U12615 (N_12615,N_12084,N_12355);
and U12616 (N_12616,N_12447,N_12001);
nand U12617 (N_12617,N_12153,N_12342);
xor U12618 (N_12618,N_12115,N_12272);
nor U12619 (N_12619,N_12021,N_12341);
xnor U12620 (N_12620,N_12267,N_12288);
or U12621 (N_12621,N_12289,N_12224);
nor U12622 (N_12622,N_12086,N_12394);
nand U12623 (N_12623,N_12206,N_12370);
nand U12624 (N_12624,N_12478,N_12134);
xor U12625 (N_12625,N_12027,N_12462);
and U12626 (N_12626,N_12096,N_12212);
or U12627 (N_12627,N_12385,N_12016);
xnor U12628 (N_12628,N_12471,N_12199);
xor U12629 (N_12629,N_12312,N_12476);
nand U12630 (N_12630,N_12175,N_12189);
and U12631 (N_12631,N_12146,N_12454);
xnor U12632 (N_12632,N_12132,N_12140);
or U12633 (N_12633,N_12485,N_12083);
xor U12634 (N_12634,N_12266,N_12264);
and U12635 (N_12635,N_12216,N_12152);
nand U12636 (N_12636,N_12413,N_12067);
nor U12637 (N_12637,N_12171,N_12457);
and U12638 (N_12638,N_12075,N_12308);
nand U12639 (N_12639,N_12215,N_12439);
and U12640 (N_12640,N_12124,N_12412);
xor U12641 (N_12641,N_12056,N_12497);
and U12642 (N_12642,N_12018,N_12280);
nor U12643 (N_12643,N_12230,N_12408);
nor U12644 (N_12644,N_12109,N_12236);
nor U12645 (N_12645,N_12348,N_12130);
xnor U12646 (N_12646,N_12110,N_12468);
and U12647 (N_12647,N_12284,N_12178);
and U12648 (N_12648,N_12223,N_12198);
xor U12649 (N_12649,N_12194,N_12053);
nand U12650 (N_12650,N_12273,N_12192);
nand U12651 (N_12651,N_12167,N_12427);
xor U12652 (N_12652,N_12162,N_12499);
xor U12653 (N_12653,N_12241,N_12009);
nor U12654 (N_12654,N_12078,N_12159);
or U12655 (N_12655,N_12065,N_12252);
nor U12656 (N_12656,N_12313,N_12157);
nor U12657 (N_12657,N_12464,N_12398);
nand U12658 (N_12658,N_12258,N_12165);
or U12659 (N_12659,N_12279,N_12345);
nor U12660 (N_12660,N_12346,N_12077);
nor U12661 (N_12661,N_12232,N_12293);
nor U12662 (N_12662,N_12117,N_12180);
nor U12663 (N_12663,N_12286,N_12376);
nor U12664 (N_12664,N_12087,N_12409);
and U12665 (N_12665,N_12054,N_12085);
and U12666 (N_12666,N_12234,N_12451);
nor U12667 (N_12667,N_12031,N_12116);
nand U12668 (N_12668,N_12432,N_12361);
and U12669 (N_12669,N_12274,N_12350);
and U12670 (N_12670,N_12367,N_12020);
and U12671 (N_12671,N_12379,N_12098);
or U12672 (N_12672,N_12423,N_12028);
nor U12673 (N_12673,N_12111,N_12015);
or U12674 (N_12674,N_12415,N_12036);
nor U12675 (N_12675,N_12257,N_12183);
nor U12676 (N_12676,N_12106,N_12253);
xnor U12677 (N_12677,N_12149,N_12363);
nor U12678 (N_12678,N_12470,N_12249);
xnor U12679 (N_12679,N_12231,N_12333);
or U12680 (N_12680,N_12200,N_12420);
nor U12681 (N_12681,N_12251,N_12406);
or U12682 (N_12682,N_12113,N_12045);
xor U12683 (N_12683,N_12052,N_12265);
nand U12684 (N_12684,N_12059,N_12336);
nand U12685 (N_12685,N_12197,N_12282);
nand U12686 (N_12686,N_12490,N_12147);
nor U12687 (N_12687,N_12327,N_12237);
nor U12688 (N_12688,N_12203,N_12484);
nor U12689 (N_12689,N_12358,N_12440);
nand U12690 (N_12690,N_12351,N_12238);
or U12691 (N_12691,N_12290,N_12256);
and U12692 (N_12692,N_12217,N_12458);
and U12693 (N_12693,N_12495,N_12037);
nor U12694 (N_12694,N_12125,N_12381);
nor U12695 (N_12695,N_12443,N_12300);
or U12696 (N_12696,N_12298,N_12202);
nand U12697 (N_12697,N_12049,N_12486);
xor U12698 (N_12698,N_12240,N_12250);
or U12699 (N_12699,N_12107,N_12108);
xor U12700 (N_12700,N_12185,N_12310);
nand U12701 (N_12701,N_12090,N_12091);
nor U12702 (N_12702,N_12463,N_12319);
xnor U12703 (N_12703,N_12494,N_12046);
or U12704 (N_12704,N_12205,N_12154);
xor U12705 (N_12705,N_12138,N_12139);
and U12706 (N_12706,N_12305,N_12477);
or U12707 (N_12707,N_12168,N_12430);
xor U12708 (N_12708,N_12032,N_12424);
or U12709 (N_12709,N_12073,N_12360);
or U12710 (N_12710,N_12022,N_12483);
xnor U12711 (N_12711,N_12328,N_12023);
and U12712 (N_12712,N_12436,N_12174);
nand U12713 (N_12713,N_12261,N_12314);
nor U12714 (N_12714,N_12095,N_12220);
nor U12715 (N_12715,N_12377,N_12466);
nand U12716 (N_12716,N_12449,N_12344);
nor U12717 (N_12717,N_12135,N_12038);
nor U12718 (N_12718,N_12301,N_12294);
nor U12719 (N_12719,N_12017,N_12304);
nand U12720 (N_12720,N_12055,N_12012);
nor U12721 (N_12721,N_12233,N_12315);
and U12722 (N_12722,N_12271,N_12411);
nor U12723 (N_12723,N_12316,N_12433);
or U12724 (N_12724,N_12489,N_12296);
or U12725 (N_12725,N_12076,N_12160);
nor U12726 (N_12726,N_12460,N_12057);
and U12727 (N_12727,N_12281,N_12498);
nor U12728 (N_12728,N_12442,N_12114);
xor U12729 (N_12729,N_12144,N_12347);
nand U12730 (N_12730,N_12204,N_12008);
and U12731 (N_12731,N_12044,N_12419);
and U12732 (N_12732,N_12383,N_12010);
nor U12733 (N_12733,N_12259,N_12322);
xor U12734 (N_12734,N_12400,N_12380);
xnor U12735 (N_12735,N_12368,N_12392);
and U12736 (N_12736,N_12201,N_12399);
nor U12737 (N_12737,N_12323,N_12193);
nor U12738 (N_12738,N_12128,N_12382);
or U12739 (N_12739,N_12246,N_12131);
or U12740 (N_12740,N_12474,N_12066);
nand U12741 (N_12741,N_12388,N_12184);
nand U12742 (N_12742,N_12278,N_12080);
xnor U12743 (N_12743,N_12069,N_12475);
nand U12744 (N_12744,N_12359,N_12219);
or U12745 (N_12745,N_12482,N_12491);
and U12746 (N_12746,N_12005,N_12000);
nor U12747 (N_12747,N_12068,N_12461);
nor U12748 (N_12748,N_12297,N_12118);
nand U12749 (N_12749,N_12372,N_12088);
or U12750 (N_12750,N_12382,N_12033);
xor U12751 (N_12751,N_12251,N_12470);
nor U12752 (N_12752,N_12000,N_12235);
xor U12753 (N_12753,N_12236,N_12259);
xnor U12754 (N_12754,N_12289,N_12129);
nor U12755 (N_12755,N_12130,N_12453);
or U12756 (N_12756,N_12162,N_12432);
or U12757 (N_12757,N_12427,N_12416);
nand U12758 (N_12758,N_12140,N_12478);
nand U12759 (N_12759,N_12310,N_12494);
xnor U12760 (N_12760,N_12048,N_12333);
xnor U12761 (N_12761,N_12247,N_12492);
xor U12762 (N_12762,N_12241,N_12095);
nand U12763 (N_12763,N_12121,N_12465);
xor U12764 (N_12764,N_12099,N_12323);
and U12765 (N_12765,N_12112,N_12428);
and U12766 (N_12766,N_12024,N_12179);
or U12767 (N_12767,N_12470,N_12262);
nor U12768 (N_12768,N_12482,N_12019);
nand U12769 (N_12769,N_12379,N_12244);
nor U12770 (N_12770,N_12324,N_12020);
and U12771 (N_12771,N_12041,N_12203);
nor U12772 (N_12772,N_12376,N_12056);
xnor U12773 (N_12773,N_12001,N_12422);
xor U12774 (N_12774,N_12119,N_12087);
nand U12775 (N_12775,N_12353,N_12405);
and U12776 (N_12776,N_12365,N_12145);
xor U12777 (N_12777,N_12368,N_12343);
nand U12778 (N_12778,N_12289,N_12215);
or U12779 (N_12779,N_12108,N_12051);
and U12780 (N_12780,N_12260,N_12359);
xor U12781 (N_12781,N_12487,N_12310);
or U12782 (N_12782,N_12499,N_12265);
and U12783 (N_12783,N_12403,N_12383);
nand U12784 (N_12784,N_12274,N_12445);
nor U12785 (N_12785,N_12354,N_12468);
nand U12786 (N_12786,N_12044,N_12379);
nand U12787 (N_12787,N_12411,N_12048);
xnor U12788 (N_12788,N_12360,N_12469);
and U12789 (N_12789,N_12056,N_12486);
nor U12790 (N_12790,N_12105,N_12295);
nor U12791 (N_12791,N_12111,N_12370);
and U12792 (N_12792,N_12120,N_12233);
nor U12793 (N_12793,N_12316,N_12474);
and U12794 (N_12794,N_12350,N_12422);
or U12795 (N_12795,N_12186,N_12063);
or U12796 (N_12796,N_12498,N_12225);
and U12797 (N_12797,N_12379,N_12096);
or U12798 (N_12798,N_12232,N_12020);
xor U12799 (N_12799,N_12240,N_12180);
or U12800 (N_12800,N_12137,N_12240);
xnor U12801 (N_12801,N_12277,N_12464);
and U12802 (N_12802,N_12037,N_12483);
nor U12803 (N_12803,N_12485,N_12291);
or U12804 (N_12804,N_12462,N_12461);
or U12805 (N_12805,N_12160,N_12064);
or U12806 (N_12806,N_12031,N_12054);
and U12807 (N_12807,N_12378,N_12007);
or U12808 (N_12808,N_12336,N_12274);
xor U12809 (N_12809,N_12213,N_12201);
or U12810 (N_12810,N_12219,N_12211);
nand U12811 (N_12811,N_12233,N_12189);
or U12812 (N_12812,N_12394,N_12345);
xnor U12813 (N_12813,N_12380,N_12134);
nor U12814 (N_12814,N_12139,N_12175);
and U12815 (N_12815,N_12141,N_12001);
xnor U12816 (N_12816,N_12068,N_12271);
nand U12817 (N_12817,N_12295,N_12019);
and U12818 (N_12818,N_12144,N_12446);
nand U12819 (N_12819,N_12130,N_12066);
nand U12820 (N_12820,N_12172,N_12390);
nand U12821 (N_12821,N_12433,N_12095);
nand U12822 (N_12822,N_12466,N_12105);
xnor U12823 (N_12823,N_12216,N_12221);
nand U12824 (N_12824,N_12372,N_12061);
nor U12825 (N_12825,N_12187,N_12016);
nand U12826 (N_12826,N_12007,N_12120);
and U12827 (N_12827,N_12052,N_12122);
or U12828 (N_12828,N_12012,N_12274);
and U12829 (N_12829,N_12168,N_12228);
nor U12830 (N_12830,N_12410,N_12247);
nand U12831 (N_12831,N_12142,N_12131);
xor U12832 (N_12832,N_12002,N_12005);
or U12833 (N_12833,N_12424,N_12094);
xnor U12834 (N_12834,N_12369,N_12351);
nor U12835 (N_12835,N_12172,N_12229);
xor U12836 (N_12836,N_12069,N_12447);
nand U12837 (N_12837,N_12470,N_12146);
or U12838 (N_12838,N_12024,N_12397);
or U12839 (N_12839,N_12392,N_12285);
nor U12840 (N_12840,N_12206,N_12209);
xor U12841 (N_12841,N_12064,N_12377);
nor U12842 (N_12842,N_12299,N_12102);
xnor U12843 (N_12843,N_12314,N_12095);
and U12844 (N_12844,N_12255,N_12236);
nor U12845 (N_12845,N_12012,N_12348);
or U12846 (N_12846,N_12133,N_12225);
nor U12847 (N_12847,N_12396,N_12117);
xnor U12848 (N_12848,N_12378,N_12323);
xor U12849 (N_12849,N_12265,N_12033);
or U12850 (N_12850,N_12185,N_12009);
xor U12851 (N_12851,N_12284,N_12023);
nor U12852 (N_12852,N_12488,N_12189);
and U12853 (N_12853,N_12134,N_12020);
and U12854 (N_12854,N_12475,N_12452);
and U12855 (N_12855,N_12383,N_12022);
and U12856 (N_12856,N_12384,N_12045);
nor U12857 (N_12857,N_12016,N_12493);
xor U12858 (N_12858,N_12454,N_12044);
xor U12859 (N_12859,N_12083,N_12338);
nand U12860 (N_12860,N_12258,N_12242);
xnor U12861 (N_12861,N_12070,N_12052);
nor U12862 (N_12862,N_12377,N_12373);
nor U12863 (N_12863,N_12463,N_12367);
and U12864 (N_12864,N_12264,N_12347);
nand U12865 (N_12865,N_12100,N_12477);
and U12866 (N_12866,N_12396,N_12447);
and U12867 (N_12867,N_12104,N_12102);
or U12868 (N_12868,N_12228,N_12056);
and U12869 (N_12869,N_12477,N_12364);
nand U12870 (N_12870,N_12495,N_12186);
nor U12871 (N_12871,N_12027,N_12496);
nand U12872 (N_12872,N_12383,N_12344);
nand U12873 (N_12873,N_12127,N_12436);
or U12874 (N_12874,N_12180,N_12421);
nor U12875 (N_12875,N_12000,N_12454);
and U12876 (N_12876,N_12063,N_12335);
or U12877 (N_12877,N_12425,N_12166);
xnor U12878 (N_12878,N_12075,N_12167);
nand U12879 (N_12879,N_12077,N_12425);
or U12880 (N_12880,N_12419,N_12073);
nand U12881 (N_12881,N_12107,N_12095);
and U12882 (N_12882,N_12237,N_12374);
and U12883 (N_12883,N_12163,N_12005);
or U12884 (N_12884,N_12089,N_12211);
nand U12885 (N_12885,N_12281,N_12106);
xor U12886 (N_12886,N_12465,N_12113);
or U12887 (N_12887,N_12458,N_12032);
and U12888 (N_12888,N_12380,N_12333);
nor U12889 (N_12889,N_12392,N_12485);
and U12890 (N_12890,N_12161,N_12042);
or U12891 (N_12891,N_12364,N_12066);
nor U12892 (N_12892,N_12172,N_12062);
xor U12893 (N_12893,N_12121,N_12434);
xor U12894 (N_12894,N_12289,N_12198);
nand U12895 (N_12895,N_12275,N_12039);
xnor U12896 (N_12896,N_12123,N_12330);
and U12897 (N_12897,N_12319,N_12227);
and U12898 (N_12898,N_12080,N_12302);
nand U12899 (N_12899,N_12219,N_12138);
nand U12900 (N_12900,N_12075,N_12039);
nor U12901 (N_12901,N_12321,N_12248);
nor U12902 (N_12902,N_12286,N_12272);
and U12903 (N_12903,N_12128,N_12044);
xnor U12904 (N_12904,N_12290,N_12425);
xor U12905 (N_12905,N_12009,N_12308);
nor U12906 (N_12906,N_12187,N_12061);
xnor U12907 (N_12907,N_12286,N_12408);
and U12908 (N_12908,N_12017,N_12174);
nor U12909 (N_12909,N_12347,N_12254);
nand U12910 (N_12910,N_12190,N_12338);
or U12911 (N_12911,N_12104,N_12243);
xor U12912 (N_12912,N_12323,N_12301);
nor U12913 (N_12913,N_12368,N_12081);
or U12914 (N_12914,N_12446,N_12320);
nand U12915 (N_12915,N_12323,N_12249);
nand U12916 (N_12916,N_12266,N_12202);
and U12917 (N_12917,N_12145,N_12045);
nor U12918 (N_12918,N_12350,N_12030);
nand U12919 (N_12919,N_12129,N_12416);
nor U12920 (N_12920,N_12240,N_12457);
xnor U12921 (N_12921,N_12121,N_12021);
xnor U12922 (N_12922,N_12386,N_12180);
or U12923 (N_12923,N_12003,N_12471);
and U12924 (N_12924,N_12185,N_12182);
nand U12925 (N_12925,N_12450,N_12383);
xnor U12926 (N_12926,N_12103,N_12033);
nor U12927 (N_12927,N_12197,N_12373);
xnor U12928 (N_12928,N_12300,N_12190);
and U12929 (N_12929,N_12072,N_12384);
nand U12930 (N_12930,N_12189,N_12481);
and U12931 (N_12931,N_12096,N_12179);
and U12932 (N_12932,N_12183,N_12367);
nor U12933 (N_12933,N_12277,N_12484);
nor U12934 (N_12934,N_12236,N_12287);
xnor U12935 (N_12935,N_12060,N_12495);
nand U12936 (N_12936,N_12449,N_12180);
nor U12937 (N_12937,N_12132,N_12370);
or U12938 (N_12938,N_12188,N_12164);
nand U12939 (N_12939,N_12024,N_12172);
nand U12940 (N_12940,N_12131,N_12439);
xor U12941 (N_12941,N_12346,N_12497);
xor U12942 (N_12942,N_12240,N_12393);
xor U12943 (N_12943,N_12327,N_12443);
xor U12944 (N_12944,N_12469,N_12086);
or U12945 (N_12945,N_12028,N_12080);
nor U12946 (N_12946,N_12134,N_12414);
and U12947 (N_12947,N_12405,N_12157);
and U12948 (N_12948,N_12097,N_12127);
xor U12949 (N_12949,N_12452,N_12317);
nor U12950 (N_12950,N_12241,N_12192);
nor U12951 (N_12951,N_12171,N_12282);
and U12952 (N_12952,N_12468,N_12061);
nand U12953 (N_12953,N_12194,N_12330);
or U12954 (N_12954,N_12156,N_12045);
nor U12955 (N_12955,N_12218,N_12045);
nand U12956 (N_12956,N_12350,N_12194);
nand U12957 (N_12957,N_12220,N_12352);
xnor U12958 (N_12958,N_12476,N_12290);
nand U12959 (N_12959,N_12047,N_12350);
or U12960 (N_12960,N_12104,N_12088);
xnor U12961 (N_12961,N_12135,N_12230);
or U12962 (N_12962,N_12342,N_12395);
xor U12963 (N_12963,N_12307,N_12393);
or U12964 (N_12964,N_12317,N_12293);
xor U12965 (N_12965,N_12204,N_12273);
or U12966 (N_12966,N_12051,N_12229);
nand U12967 (N_12967,N_12225,N_12472);
nand U12968 (N_12968,N_12087,N_12391);
nand U12969 (N_12969,N_12064,N_12422);
nand U12970 (N_12970,N_12065,N_12193);
nor U12971 (N_12971,N_12439,N_12100);
and U12972 (N_12972,N_12400,N_12156);
or U12973 (N_12973,N_12200,N_12431);
xor U12974 (N_12974,N_12046,N_12012);
xor U12975 (N_12975,N_12464,N_12015);
or U12976 (N_12976,N_12227,N_12486);
and U12977 (N_12977,N_12268,N_12460);
and U12978 (N_12978,N_12413,N_12455);
or U12979 (N_12979,N_12465,N_12131);
and U12980 (N_12980,N_12298,N_12204);
nor U12981 (N_12981,N_12388,N_12090);
nand U12982 (N_12982,N_12005,N_12335);
nand U12983 (N_12983,N_12232,N_12075);
xnor U12984 (N_12984,N_12065,N_12118);
xor U12985 (N_12985,N_12271,N_12358);
nand U12986 (N_12986,N_12370,N_12291);
nand U12987 (N_12987,N_12139,N_12415);
xnor U12988 (N_12988,N_12128,N_12076);
nand U12989 (N_12989,N_12027,N_12148);
nand U12990 (N_12990,N_12269,N_12164);
xor U12991 (N_12991,N_12445,N_12002);
or U12992 (N_12992,N_12240,N_12293);
nand U12993 (N_12993,N_12021,N_12493);
and U12994 (N_12994,N_12310,N_12308);
nand U12995 (N_12995,N_12177,N_12088);
and U12996 (N_12996,N_12344,N_12104);
or U12997 (N_12997,N_12106,N_12473);
nor U12998 (N_12998,N_12397,N_12356);
or U12999 (N_12999,N_12107,N_12216);
or U13000 (N_13000,N_12853,N_12712);
or U13001 (N_13001,N_12823,N_12788);
nand U13002 (N_13002,N_12655,N_12854);
and U13003 (N_13003,N_12771,N_12711);
xnor U13004 (N_13004,N_12809,N_12814);
nand U13005 (N_13005,N_12603,N_12919);
nand U13006 (N_13006,N_12954,N_12787);
and U13007 (N_13007,N_12560,N_12967);
and U13008 (N_13008,N_12658,N_12737);
or U13009 (N_13009,N_12745,N_12609);
or U13010 (N_13010,N_12894,N_12836);
or U13011 (N_13011,N_12974,N_12961);
nand U13012 (N_13012,N_12844,N_12707);
or U13013 (N_13013,N_12861,N_12555);
or U13014 (N_13014,N_12671,N_12618);
nand U13015 (N_13015,N_12732,N_12512);
nor U13016 (N_13016,N_12514,N_12834);
and U13017 (N_13017,N_12753,N_12821);
nand U13018 (N_13018,N_12623,N_12940);
xor U13019 (N_13019,N_12587,N_12970);
or U13020 (N_13020,N_12900,N_12932);
or U13021 (N_13021,N_12755,N_12918);
and U13022 (N_13022,N_12741,N_12598);
nand U13023 (N_13023,N_12543,N_12696);
and U13024 (N_13024,N_12622,N_12736);
xor U13025 (N_13025,N_12681,N_12520);
and U13026 (N_13026,N_12518,N_12786);
or U13027 (N_13027,N_12950,N_12629);
nand U13028 (N_13028,N_12626,N_12799);
or U13029 (N_13029,N_12537,N_12693);
or U13030 (N_13030,N_12632,N_12563);
or U13031 (N_13031,N_12766,N_12604);
and U13032 (N_13032,N_12643,N_12890);
nand U13033 (N_13033,N_12503,N_12570);
or U13034 (N_13034,N_12993,N_12927);
and U13035 (N_13035,N_12796,N_12774);
nor U13036 (N_13036,N_12778,N_12558);
and U13037 (N_13037,N_12602,N_12677);
or U13038 (N_13038,N_12931,N_12678);
nand U13039 (N_13039,N_12540,N_12735);
nand U13040 (N_13040,N_12569,N_12656);
nor U13041 (N_13041,N_12627,N_12904);
xnor U13042 (N_13042,N_12977,N_12800);
nand U13043 (N_13043,N_12901,N_12638);
or U13044 (N_13044,N_12783,N_12907);
and U13045 (N_13045,N_12748,N_12840);
xor U13046 (N_13046,N_12532,N_12542);
xor U13047 (N_13047,N_12867,N_12600);
or U13048 (N_13048,N_12651,N_12714);
xnor U13049 (N_13049,N_12946,N_12534);
nor U13050 (N_13050,N_12581,N_12607);
or U13051 (N_13051,N_12945,N_12789);
or U13052 (N_13052,N_12926,N_12841);
and U13053 (N_13053,N_12860,N_12708);
nor U13054 (N_13054,N_12862,N_12885);
and U13055 (N_13055,N_12874,N_12506);
and U13056 (N_13056,N_12527,N_12716);
nor U13057 (N_13057,N_12733,N_12963);
or U13058 (N_13058,N_12815,N_12980);
nand U13059 (N_13059,N_12857,N_12565);
or U13060 (N_13060,N_12688,N_12710);
or U13061 (N_13061,N_12849,N_12759);
or U13062 (N_13062,N_12510,N_12682);
nor U13063 (N_13063,N_12808,N_12972);
xor U13064 (N_13064,N_12728,N_12917);
nand U13065 (N_13065,N_12694,N_12675);
and U13066 (N_13066,N_12553,N_12507);
and U13067 (N_13067,N_12591,N_12513);
nor U13068 (N_13068,N_12526,N_12947);
xor U13069 (N_13069,N_12567,N_12892);
nand U13070 (N_13070,N_12580,N_12976);
or U13071 (N_13071,N_12846,N_12948);
nor U13072 (N_13072,N_12752,N_12538);
nor U13073 (N_13073,N_12848,N_12822);
nor U13074 (N_13074,N_12920,N_12785);
or U13075 (N_13075,N_12646,N_12843);
or U13076 (N_13076,N_12556,N_12606);
nand U13077 (N_13077,N_12636,N_12630);
nor U13078 (N_13078,N_12888,N_12686);
nor U13079 (N_13079,N_12672,N_12751);
nor U13080 (N_13080,N_12650,N_12767);
nand U13081 (N_13081,N_12666,N_12654);
and U13082 (N_13082,N_12747,N_12500);
or U13083 (N_13083,N_12697,N_12943);
or U13084 (N_13084,N_12519,N_12936);
or U13085 (N_13085,N_12583,N_12552);
and U13086 (N_13086,N_12575,N_12589);
nor U13087 (N_13087,N_12812,N_12955);
and U13088 (N_13088,N_12673,N_12517);
nand U13089 (N_13089,N_12839,N_12605);
and U13090 (N_13090,N_12644,N_12760);
nand U13091 (N_13091,N_12897,N_12505);
or U13092 (N_13092,N_12617,N_12908);
or U13093 (N_13093,N_12979,N_12877);
xnor U13094 (N_13094,N_12801,N_12978);
nor U13095 (N_13095,N_12880,N_12964);
or U13096 (N_13096,N_12749,N_12971);
nor U13097 (N_13097,N_12721,N_12842);
or U13098 (N_13098,N_12929,N_12594);
nor U13099 (N_13099,N_12784,N_12795);
or U13100 (N_13100,N_12938,N_12831);
xor U13101 (N_13101,N_12949,N_12962);
xor U13102 (N_13102,N_12889,N_12991);
xor U13103 (N_13103,N_12574,N_12739);
nor U13104 (N_13104,N_12521,N_12935);
or U13105 (N_13105,N_12610,N_12838);
nand U13106 (N_13106,N_12664,N_12983);
or U13107 (N_13107,N_12549,N_12984);
nor U13108 (N_13108,N_12873,N_12941);
nand U13109 (N_13109,N_12699,N_12613);
and U13110 (N_13110,N_12756,N_12529);
or U13111 (N_13111,N_12595,N_12930);
xnor U13112 (N_13112,N_12729,N_12764);
xnor U13113 (N_13113,N_12516,N_12525);
nor U13114 (N_13114,N_12743,N_12813);
or U13115 (N_13115,N_12807,N_12988);
nand U13116 (N_13116,N_12916,N_12817);
or U13117 (N_13117,N_12579,N_12858);
nand U13118 (N_13118,N_12922,N_12535);
xor U13119 (N_13119,N_12875,N_12550);
and U13120 (N_13120,N_12554,N_12968);
xnor U13121 (N_13121,N_12965,N_12830);
nand U13122 (N_13122,N_12829,N_12640);
or U13123 (N_13123,N_12706,N_12902);
xnor U13124 (N_13124,N_12508,N_12698);
nor U13125 (N_13125,N_12794,N_12746);
and U13126 (N_13126,N_12999,N_12937);
and U13127 (N_13127,N_12910,N_12725);
xor U13128 (N_13128,N_12742,N_12744);
nor U13129 (N_13129,N_12523,N_12726);
or U13130 (N_13130,N_12703,N_12661);
nor U13131 (N_13131,N_12960,N_12818);
xor U13132 (N_13132,N_12545,N_12798);
and U13133 (N_13133,N_12966,N_12905);
and U13134 (N_13134,N_12683,N_12832);
xor U13135 (N_13135,N_12691,N_12845);
xor U13136 (N_13136,N_12566,N_12653);
nand U13137 (N_13137,N_12548,N_12701);
and U13138 (N_13138,N_12868,N_12668);
nand U13139 (N_13139,N_12705,N_12913);
or U13140 (N_13140,N_12559,N_12928);
and U13141 (N_13141,N_12670,N_12652);
nor U13142 (N_13142,N_12994,N_12981);
xor U13143 (N_13143,N_12820,N_12722);
xor U13144 (N_13144,N_12776,N_12687);
nand U13145 (N_13145,N_12684,N_12669);
nor U13146 (N_13146,N_12772,N_12806);
or U13147 (N_13147,N_12770,N_12593);
xor U13148 (N_13148,N_12792,N_12588);
or U13149 (N_13149,N_12557,N_12957);
nand U13150 (N_13150,N_12833,N_12871);
nor U13151 (N_13151,N_12649,N_12996);
and U13152 (N_13152,N_12645,N_12522);
or U13153 (N_13153,N_12620,N_12782);
or U13154 (N_13154,N_12989,N_12637);
and U13155 (N_13155,N_12866,N_12738);
nor U13156 (N_13156,N_12590,N_12576);
nor U13157 (N_13157,N_12953,N_12952);
nand U13158 (N_13158,N_12828,N_12956);
nand U13159 (N_13159,N_12859,N_12855);
and U13160 (N_13160,N_12511,N_12660);
xor U13161 (N_13161,N_12524,N_12585);
or U13162 (N_13162,N_12596,N_12856);
xor U13163 (N_13163,N_12723,N_12642);
nor U13164 (N_13164,N_12572,N_12597);
or U13165 (N_13165,N_12612,N_12633);
nor U13166 (N_13166,N_12509,N_12992);
nand U13167 (N_13167,N_12601,N_12758);
and U13168 (N_13168,N_12881,N_12765);
or U13169 (N_13169,N_12539,N_12679);
xor U13170 (N_13170,N_12982,N_12754);
nor U13171 (N_13171,N_12625,N_12912);
xor U13172 (N_13172,N_12939,N_12925);
nand U13173 (N_13173,N_12577,N_12634);
xor U13174 (N_13174,N_12869,N_12884);
xnor U13175 (N_13175,N_12793,N_12731);
and U13176 (N_13176,N_12616,N_12911);
nand U13177 (N_13177,N_12730,N_12611);
nor U13178 (N_13178,N_12803,N_12986);
or U13179 (N_13179,N_12872,N_12680);
nand U13180 (N_13180,N_12504,N_12837);
and U13181 (N_13181,N_12779,N_12958);
nand U13182 (N_13182,N_12985,N_12893);
xnor U13183 (N_13183,N_12921,N_12826);
and U13184 (N_13184,N_12895,N_12657);
and U13185 (N_13185,N_12805,N_12827);
nor U13186 (N_13186,N_12719,N_12891);
nor U13187 (N_13187,N_12761,N_12536);
xnor U13188 (N_13188,N_12791,N_12882);
nor U13189 (N_13189,N_12528,N_12641);
and U13190 (N_13190,N_12899,N_12797);
nand U13191 (N_13191,N_12715,N_12998);
nor U13192 (N_13192,N_12824,N_12777);
nor U13193 (N_13193,N_12663,N_12573);
nand U13194 (N_13194,N_12863,N_12987);
nand U13195 (N_13195,N_12531,N_12690);
nor U13196 (N_13196,N_12924,N_12763);
and U13197 (N_13197,N_12934,N_12773);
and U13198 (N_13198,N_12811,N_12909);
or U13199 (N_13199,N_12933,N_12720);
or U13200 (N_13200,N_12906,N_12944);
or U13201 (N_13201,N_12619,N_12847);
nand U13202 (N_13202,N_12750,N_12997);
nor U13203 (N_13203,N_12802,N_12851);
nand U13204 (N_13204,N_12647,N_12727);
xor U13205 (N_13205,N_12614,N_12975);
xor U13206 (N_13206,N_12586,N_12541);
and U13207 (N_13207,N_12790,N_12969);
and U13208 (N_13208,N_12667,N_12659);
xor U13209 (N_13209,N_12578,N_12810);
nand U13210 (N_13210,N_12886,N_12631);
xnor U13211 (N_13211,N_12870,N_12835);
or U13212 (N_13212,N_12775,N_12724);
or U13213 (N_13213,N_12592,N_12959);
or U13214 (N_13214,N_12819,N_12883);
and U13215 (N_13215,N_12768,N_12571);
nor U13216 (N_13216,N_12898,N_12825);
and U13217 (N_13217,N_12582,N_12702);
xor U13218 (N_13218,N_12816,N_12973);
and U13219 (N_13219,N_12515,N_12689);
xnor U13220 (N_13220,N_12713,N_12757);
or U13221 (N_13221,N_12879,N_12615);
xor U13222 (N_13222,N_12740,N_12662);
xnor U13223 (N_13223,N_12533,N_12568);
nor U13224 (N_13224,N_12564,N_12781);
nor U13225 (N_13225,N_12546,N_12584);
and U13226 (N_13226,N_12608,N_12876);
and U13227 (N_13227,N_12915,N_12709);
nand U13228 (N_13228,N_12864,N_12718);
or U13229 (N_13229,N_12704,N_12562);
and U13230 (N_13230,N_12695,N_12850);
xor U13231 (N_13231,N_12914,N_12635);
and U13232 (N_13232,N_12621,N_12639);
xor U13233 (N_13233,N_12923,N_12674);
nor U13234 (N_13234,N_12551,N_12544);
or U13235 (N_13235,N_12502,N_12734);
and U13236 (N_13236,N_12561,N_12717);
and U13237 (N_13237,N_12990,N_12530);
nand U13238 (N_13238,N_12804,N_12665);
nor U13239 (N_13239,N_12852,N_12995);
or U13240 (N_13240,N_12648,N_12762);
nand U13241 (N_13241,N_12942,N_12887);
nand U13242 (N_13242,N_12951,N_12780);
or U13243 (N_13243,N_12676,N_12903);
and U13244 (N_13244,N_12624,N_12628);
xor U13245 (N_13245,N_12599,N_12547);
nand U13246 (N_13246,N_12685,N_12878);
or U13247 (N_13247,N_12865,N_12692);
nand U13248 (N_13248,N_12769,N_12700);
and U13249 (N_13249,N_12896,N_12501);
and U13250 (N_13250,N_12860,N_12749);
or U13251 (N_13251,N_12717,N_12567);
and U13252 (N_13252,N_12911,N_12774);
and U13253 (N_13253,N_12777,N_12966);
nor U13254 (N_13254,N_12998,N_12789);
nor U13255 (N_13255,N_12893,N_12582);
nor U13256 (N_13256,N_12666,N_12778);
xnor U13257 (N_13257,N_12965,N_12710);
xnor U13258 (N_13258,N_12643,N_12572);
nor U13259 (N_13259,N_12994,N_12703);
nand U13260 (N_13260,N_12843,N_12812);
xnor U13261 (N_13261,N_12613,N_12930);
xnor U13262 (N_13262,N_12699,N_12785);
or U13263 (N_13263,N_12744,N_12866);
nand U13264 (N_13264,N_12812,N_12918);
nand U13265 (N_13265,N_12662,N_12618);
xnor U13266 (N_13266,N_12884,N_12529);
xnor U13267 (N_13267,N_12869,N_12689);
and U13268 (N_13268,N_12768,N_12599);
nor U13269 (N_13269,N_12677,N_12919);
and U13270 (N_13270,N_12981,N_12666);
nand U13271 (N_13271,N_12721,N_12846);
nor U13272 (N_13272,N_12664,N_12563);
or U13273 (N_13273,N_12525,N_12502);
and U13274 (N_13274,N_12632,N_12708);
xnor U13275 (N_13275,N_12801,N_12821);
nor U13276 (N_13276,N_12969,N_12535);
or U13277 (N_13277,N_12822,N_12757);
or U13278 (N_13278,N_12985,N_12972);
and U13279 (N_13279,N_12542,N_12723);
nand U13280 (N_13280,N_12753,N_12731);
or U13281 (N_13281,N_12772,N_12617);
and U13282 (N_13282,N_12784,N_12774);
nand U13283 (N_13283,N_12918,N_12830);
or U13284 (N_13284,N_12716,N_12548);
or U13285 (N_13285,N_12715,N_12681);
or U13286 (N_13286,N_12546,N_12974);
xor U13287 (N_13287,N_12716,N_12595);
nand U13288 (N_13288,N_12739,N_12657);
and U13289 (N_13289,N_12898,N_12522);
xor U13290 (N_13290,N_12889,N_12738);
xnor U13291 (N_13291,N_12897,N_12977);
and U13292 (N_13292,N_12990,N_12710);
nor U13293 (N_13293,N_12696,N_12677);
nand U13294 (N_13294,N_12883,N_12762);
or U13295 (N_13295,N_12500,N_12708);
xor U13296 (N_13296,N_12752,N_12990);
nor U13297 (N_13297,N_12722,N_12695);
nand U13298 (N_13298,N_12503,N_12748);
or U13299 (N_13299,N_12785,N_12542);
and U13300 (N_13300,N_12743,N_12886);
nor U13301 (N_13301,N_12852,N_12922);
or U13302 (N_13302,N_12682,N_12741);
and U13303 (N_13303,N_12654,N_12698);
nor U13304 (N_13304,N_12970,N_12541);
nor U13305 (N_13305,N_12510,N_12715);
xnor U13306 (N_13306,N_12544,N_12895);
nand U13307 (N_13307,N_12803,N_12921);
nor U13308 (N_13308,N_12931,N_12888);
xnor U13309 (N_13309,N_12791,N_12697);
nand U13310 (N_13310,N_12609,N_12583);
nand U13311 (N_13311,N_12972,N_12799);
xnor U13312 (N_13312,N_12647,N_12816);
and U13313 (N_13313,N_12597,N_12746);
or U13314 (N_13314,N_12866,N_12859);
nand U13315 (N_13315,N_12605,N_12595);
nor U13316 (N_13316,N_12982,N_12747);
nand U13317 (N_13317,N_12508,N_12771);
nand U13318 (N_13318,N_12964,N_12704);
nand U13319 (N_13319,N_12936,N_12802);
xor U13320 (N_13320,N_12873,N_12786);
and U13321 (N_13321,N_12807,N_12758);
and U13322 (N_13322,N_12904,N_12748);
nand U13323 (N_13323,N_12526,N_12951);
and U13324 (N_13324,N_12550,N_12607);
nor U13325 (N_13325,N_12767,N_12544);
and U13326 (N_13326,N_12581,N_12540);
nand U13327 (N_13327,N_12666,N_12928);
nand U13328 (N_13328,N_12529,N_12833);
nand U13329 (N_13329,N_12923,N_12715);
nand U13330 (N_13330,N_12816,N_12646);
nor U13331 (N_13331,N_12517,N_12789);
nor U13332 (N_13332,N_12652,N_12921);
and U13333 (N_13333,N_12832,N_12770);
and U13334 (N_13334,N_12534,N_12564);
nor U13335 (N_13335,N_12797,N_12783);
nand U13336 (N_13336,N_12600,N_12741);
and U13337 (N_13337,N_12979,N_12994);
xor U13338 (N_13338,N_12514,N_12504);
nand U13339 (N_13339,N_12563,N_12668);
and U13340 (N_13340,N_12988,N_12883);
and U13341 (N_13341,N_12855,N_12686);
nor U13342 (N_13342,N_12742,N_12864);
and U13343 (N_13343,N_12740,N_12873);
nand U13344 (N_13344,N_12713,N_12777);
nand U13345 (N_13345,N_12612,N_12743);
or U13346 (N_13346,N_12672,N_12557);
xor U13347 (N_13347,N_12814,N_12751);
and U13348 (N_13348,N_12860,N_12509);
nand U13349 (N_13349,N_12691,N_12963);
or U13350 (N_13350,N_12874,N_12714);
nand U13351 (N_13351,N_12618,N_12817);
xor U13352 (N_13352,N_12880,N_12596);
nor U13353 (N_13353,N_12505,N_12833);
and U13354 (N_13354,N_12845,N_12948);
and U13355 (N_13355,N_12973,N_12735);
nand U13356 (N_13356,N_12740,N_12643);
and U13357 (N_13357,N_12761,N_12552);
nor U13358 (N_13358,N_12673,N_12740);
xnor U13359 (N_13359,N_12929,N_12920);
and U13360 (N_13360,N_12797,N_12585);
xor U13361 (N_13361,N_12805,N_12623);
and U13362 (N_13362,N_12934,N_12746);
nor U13363 (N_13363,N_12898,N_12999);
and U13364 (N_13364,N_12753,N_12832);
or U13365 (N_13365,N_12651,N_12908);
and U13366 (N_13366,N_12557,N_12912);
nor U13367 (N_13367,N_12608,N_12699);
and U13368 (N_13368,N_12636,N_12918);
xor U13369 (N_13369,N_12896,N_12970);
nand U13370 (N_13370,N_12509,N_12583);
nor U13371 (N_13371,N_12527,N_12591);
xor U13372 (N_13372,N_12960,N_12648);
and U13373 (N_13373,N_12835,N_12826);
xor U13374 (N_13374,N_12939,N_12902);
xnor U13375 (N_13375,N_12930,N_12983);
nand U13376 (N_13376,N_12624,N_12860);
nor U13377 (N_13377,N_12512,N_12628);
nor U13378 (N_13378,N_12559,N_12790);
nand U13379 (N_13379,N_12717,N_12736);
nor U13380 (N_13380,N_12910,N_12503);
nor U13381 (N_13381,N_12667,N_12618);
xnor U13382 (N_13382,N_12696,N_12877);
nor U13383 (N_13383,N_12849,N_12895);
and U13384 (N_13384,N_12516,N_12532);
xor U13385 (N_13385,N_12553,N_12718);
nor U13386 (N_13386,N_12515,N_12882);
or U13387 (N_13387,N_12910,N_12903);
and U13388 (N_13388,N_12880,N_12845);
xnor U13389 (N_13389,N_12547,N_12626);
nor U13390 (N_13390,N_12842,N_12740);
or U13391 (N_13391,N_12955,N_12698);
and U13392 (N_13392,N_12505,N_12976);
or U13393 (N_13393,N_12651,N_12646);
and U13394 (N_13394,N_12754,N_12623);
nand U13395 (N_13395,N_12641,N_12750);
nor U13396 (N_13396,N_12731,N_12903);
and U13397 (N_13397,N_12926,N_12907);
nand U13398 (N_13398,N_12799,N_12789);
nand U13399 (N_13399,N_12940,N_12876);
nor U13400 (N_13400,N_12598,N_12830);
nor U13401 (N_13401,N_12739,N_12501);
and U13402 (N_13402,N_12501,N_12915);
or U13403 (N_13403,N_12941,N_12683);
or U13404 (N_13404,N_12724,N_12626);
and U13405 (N_13405,N_12774,N_12775);
xnor U13406 (N_13406,N_12632,N_12933);
or U13407 (N_13407,N_12913,N_12813);
nor U13408 (N_13408,N_12554,N_12763);
and U13409 (N_13409,N_12777,N_12644);
xnor U13410 (N_13410,N_12961,N_12683);
nand U13411 (N_13411,N_12532,N_12789);
xor U13412 (N_13412,N_12811,N_12558);
or U13413 (N_13413,N_12968,N_12833);
xnor U13414 (N_13414,N_12516,N_12928);
or U13415 (N_13415,N_12913,N_12653);
and U13416 (N_13416,N_12987,N_12705);
nand U13417 (N_13417,N_12543,N_12980);
nand U13418 (N_13418,N_12606,N_12877);
nand U13419 (N_13419,N_12612,N_12768);
and U13420 (N_13420,N_12647,N_12737);
xor U13421 (N_13421,N_12573,N_12974);
nand U13422 (N_13422,N_12757,N_12965);
xnor U13423 (N_13423,N_12991,N_12984);
and U13424 (N_13424,N_12789,N_12908);
and U13425 (N_13425,N_12534,N_12809);
and U13426 (N_13426,N_12676,N_12608);
or U13427 (N_13427,N_12597,N_12831);
and U13428 (N_13428,N_12676,N_12907);
xnor U13429 (N_13429,N_12907,N_12819);
nand U13430 (N_13430,N_12787,N_12618);
or U13431 (N_13431,N_12905,N_12868);
or U13432 (N_13432,N_12937,N_12784);
nor U13433 (N_13433,N_12825,N_12981);
or U13434 (N_13434,N_12899,N_12922);
and U13435 (N_13435,N_12989,N_12845);
xnor U13436 (N_13436,N_12560,N_12503);
nand U13437 (N_13437,N_12986,N_12634);
nor U13438 (N_13438,N_12731,N_12835);
or U13439 (N_13439,N_12990,N_12951);
or U13440 (N_13440,N_12955,N_12796);
and U13441 (N_13441,N_12837,N_12567);
or U13442 (N_13442,N_12996,N_12692);
or U13443 (N_13443,N_12729,N_12705);
or U13444 (N_13444,N_12938,N_12810);
nand U13445 (N_13445,N_12517,N_12935);
or U13446 (N_13446,N_12762,N_12841);
or U13447 (N_13447,N_12868,N_12800);
or U13448 (N_13448,N_12940,N_12558);
nor U13449 (N_13449,N_12693,N_12690);
and U13450 (N_13450,N_12886,N_12571);
nor U13451 (N_13451,N_12936,N_12987);
or U13452 (N_13452,N_12528,N_12935);
and U13453 (N_13453,N_12790,N_12517);
and U13454 (N_13454,N_12811,N_12769);
nand U13455 (N_13455,N_12539,N_12881);
xnor U13456 (N_13456,N_12993,N_12822);
nand U13457 (N_13457,N_12722,N_12852);
or U13458 (N_13458,N_12606,N_12873);
xor U13459 (N_13459,N_12955,N_12706);
nand U13460 (N_13460,N_12666,N_12883);
xnor U13461 (N_13461,N_12593,N_12825);
or U13462 (N_13462,N_12834,N_12500);
xnor U13463 (N_13463,N_12993,N_12514);
nor U13464 (N_13464,N_12865,N_12770);
xor U13465 (N_13465,N_12674,N_12984);
and U13466 (N_13466,N_12855,N_12674);
and U13467 (N_13467,N_12679,N_12555);
xor U13468 (N_13468,N_12931,N_12835);
nand U13469 (N_13469,N_12904,N_12886);
nor U13470 (N_13470,N_12842,N_12520);
nand U13471 (N_13471,N_12968,N_12591);
nor U13472 (N_13472,N_12783,N_12799);
nor U13473 (N_13473,N_12537,N_12675);
nand U13474 (N_13474,N_12657,N_12735);
xnor U13475 (N_13475,N_12774,N_12760);
xor U13476 (N_13476,N_12807,N_12747);
or U13477 (N_13477,N_12919,N_12935);
nand U13478 (N_13478,N_12521,N_12621);
nand U13479 (N_13479,N_12876,N_12699);
nor U13480 (N_13480,N_12518,N_12694);
and U13481 (N_13481,N_12652,N_12700);
xnor U13482 (N_13482,N_12865,N_12590);
xnor U13483 (N_13483,N_12709,N_12579);
nor U13484 (N_13484,N_12866,N_12553);
nor U13485 (N_13485,N_12580,N_12737);
nor U13486 (N_13486,N_12694,N_12530);
nand U13487 (N_13487,N_12767,N_12768);
xnor U13488 (N_13488,N_12889,N_12602);
nor U13489 (N_13489,N_12677,N_12598);
and U13490 (N_13490,N_12694,N_12707);
nor U13491 (N_13491,N_12920,N_12508);
nor U13492 (N_13492,N_12698,N_12503);
nor U13493 (N_13493,N_12926,N_12520);
nor U13494 (N_13494,N_12937,N_12507);
and U13495 (N_13495,N_12643,N_12863);
or U13496 (N_13496,N_12968,N_12573);
nor U13497 (N_13497,N_12799,N_12945);
xor U13498 (N_13498,N_12774,N_12873);
and U13499 (N_13499,N_12716,N_12665);
nand U13500 (N_13500,N_13051,N_13259);
or U13501 (N_13501,N_13142,N_13186);
nor U13502 (N_13502,N_13412,N_13193);
or U13503 (N_13503,N_13467,N_13289);
xor U13504 (N_13504,N_13099,N_13457);
and U13505 (N_13505,N_13298,N_13162);
and U13506 (N_13506,N_13465,N_13473);
nand U13507 (N_13507,N_13198,N_13338);
or U13508 (N_13508,N_13064,N_13265);
nand U13509 (N_13509,N_13336,N_13464);
nor U13510 (N_13510,N_13287,N_13144);
nand U13511 (N_13511,N_13373,N_13213);
nand U13512 (N_13512,N_13155,N_13368);
nand U13513 (N_13513,N_13078,N_13156);
nor U13514 (N_13514,N_13399,N_13074);
and U13515 (N_13515,N_13366,N_13409);
or U13516 (N_13516,N_13286,N_13341);
nand U13517 (N_13517,N_13154,N_13176);
nand U13518 (N_13518,N_13422,N_13306);
or U13519 (N_13519,N_13216,N_13407);
nand U13520 (N_13520,N_13069,N_13046);
nor U13521 (N_13521,N_13423,N_13278);
nor U13522 (N_13522,N_13451,N_13288);
nand U13523 (N_13523,N_13333,N_13182);
nand U13524 (N_13524,N_13243,N_13017);
or U13525 (N_13525,N_13427,N_13008);
nand U13526 (N_13526,N_13348,N_13299);
nand U13527 (N_13527,N_13215,N_13357);
xor U13528 (N_13528,N_13222,N_13197);
and U13529 (N_13529,N_13461,N_13033);
nand U13530 (N_13530,N_13143,N_13150);
nand U13531 (N_13531,N_13170,N_13443);
nand U13532 (N_13532,N_13095,N_13480);
nand U13533 (N_13533,N_13484,N_13054);
nor U13534 (N_13534,N_13071,N_13383);
and U13535 (N_13535,N_13083,N_13463);
and U13536 (N_13536,N_13019,N_13321);
and U13537 (N_13537,N_13320,N_13126);
xnor U13538 (N_13538,N_13007,N_13195);
nand U13539 (N_13539,N_13135,N_13489);
nor U13540 (N_13540,N_13402,N_13362);
and U13541 (N_13541,N_13108,N_13165);
xor U13542 (N_13542,N_13202,N_13440);
nor U13543 (N_13543,N_13358,N_13158);
or U13544 (N_13544,N_13497,N_13027);
nor U13545 (N_13545,N_13335,N_13055);
nor U13546 (N_13546,N_13456,N_13393);
nor U13547 (N_13547,N_13025,N_13455);
xor U13548 (N_13548,N_13475,N_13248);
and U13549 (N_13549,N_13120,N_13096);
xor U13550 (N_13550,N_13469,N_13075);
or U13551 (N_13551,N_13392,N_13118);
nand U13552 (N_13552,N_13410,N_13325);
or U13553 (N_13553,N_13183,N_13448);
and U13554 (N_13554,N_13491,N_13056);
and U13555 (N_13555,N_13326,N_13225);
nor U13556 (N_13556,N_13136,N_13363);
and U13557 (N_13557,N_13048,N_13230);
nor U13558 (N_13558,N_13349,N_13486);
nand U13559 (N_13559,N_13194,N_13103);
xor U13560 (N_13560,N_13129,N_13240);
and U13561 (N_13561,N_13232,N_13262);
nand U13562 (N_13562,N_13458,N_13107);
and U13563 (N_13563,N_13023,N_13112);
nor U13564 (N_13564,N_13203,N_13449);
xor U13565 (N_13565,N_13192,N_13166);
and U13566 (N_13566,N_13137,N_13400);
nand U13567 (N_13567,N_13324,N_13004);
nor U13568 (N_13568,N_13468,N_13483);
and U13569 (N_13569,N_13346,N_13152);
or U13570 (N_13570,N_13236,N_13452);
or U13571 (N_13571,N_13174,N_13413);
nand U13572 (N_13572,N_13221,N_13115);
or U13573 (N_13573,N_13426,N_13266);
nand U13574 (N_13574,N_13030,N_13429);
nor U13575 (N_13575,N_13050,N_13031);
nor U13576 (N_13576,N_13140,N_13076);
nor U13577 (N_13577,N_13009,N_13488);
nor U13578 (N_13578,N_13442,N_13347);
nand U13579 (N_13579,N_13084,N_13261);
and U13580 (N_13580,N_13001,N_13068);
and U13581 (N_13581,N_13408,N_13220);
or U13582 (N_13582,N_13043,N_13125);
nor U13583 (N_13583,N_13160,N_13376);
xnor U13584 (N_13584,N_13000,N_13028);
nor U13585 (N_13585,N_13119,N_13089);
and U13586 (N_13586,N_13281,N_13411);
nand U13587 (N_13587,N_13284,N_13040);
and U13588 (N_13588,N_13447,N_13179);
xnor U13589 (N_13589,N_13188,N_13312);
or U13590 (N_13590,N_13102,N_13303);
and U13591 (N_13591,N_13344,N_13356);
or U13592 (N_13592,N_13035,N_13481);
nor U13593 (N_13593,N_13010,N_13132);
nor U13594 (N_13594,N_13328,N_13157);
or U13595 (N_13595,N_13257,N_13340);
xnor U13596 (N_13596,N_13477,N_13178);
nand U13597 (N_13597,N_13476,N_13020);
or U13598 (N_13598,N_13351,N_13204);
or U13599 (N_13599,N_13205,N_13384);
nor U13600 (N_13600,N_13238,N_13280);
nand U13601 (N_13601,N_13106,N_13044);
or U13602 (N_13602,N_13191,N_13293);
nor U13603 (N_13603,N_13372,N_13342);
xor U13604 (N_13604,N_13245,N_13370);
and U13605 (N_13605,N_13224,N_13207);
nor U13606 (N_13606,N_13310,N_13304);
nand U13607 (N_13607,N_13271,N_13208);
nand U13608 (N_13608,N_13470,N_13210);
nand U13609 (N_13609,N_13454,N_13403);
nor U13610 (N_13610,N_13450,N_13382);
and U13611 (N_13611,N_13282,N_13290);
nand U13612 (N_13612,N_13005,N_13438);
xor U13613 (N_13613,N_13060,N_13496);
nor U13614 (N_13614,N_13113,N_13459);
nor U13615 (N_13615,N_13141,N_13406);
xor U13616 (N_13616,N_13177,N_13295);
or U13617 (N_13617,N_13337,N_13082);
nand U13618 (N_13618,N_13301,N_13472);
nand U13619 (N_13619,N_13042,N_13153);
or U13620 (N_13620,N_13227,N_13159);
nor U13621 (N_13621,N_13168,N_13432);
xnor U13622 (N_13622,N_13386,N_13087);
or U13623 (N_13623,N_13053,N_13474);
and U13624 (N_13624,N_13223,N_13498);
nand U13625 (N_13625,N_13434,N_13077);
nand U13626 (N_13626,N_13279,N_13499);
xor U13627 (N_13627,N_13199,N_13490);
or U13628 (N_13628,N_13131,N_13441);
nand U13629 (N_13629,N_13385,N_13127);
and U13630 (N_13630,N_13292,N_13479);
or U13631 (N_13631,N_13419,N_13418);
and U13632 (N_13632,N_13369,N_13315);
nand U13633 (N_13633,N_13329,N_13045);
nand U13634 (N_13634,N_13263,N_13163);
nor U13635 (N_13635,N_13181,N_13080);
and U13636 (N_13636,N_13274,N_13218);
or U13637 (N_13637,N_13311,N_13057);
nand U13638 (N_13638,N_13145,N_13308);
or U13639 (N_13639,N_13133,N_13047);
xnor U13640 (N_13640,N_13038,N_13063);
nand U13641 (N_13641,N_13273,N_13388);
or U13642 (N_13642,N_13149,N_13164);
nand U13643 (N_13643,N_13275,N_13002);
xor U13644 (N_13644,N_13254,N_13110);
and U13645 (N_13645,N_13217,N_13122);
and U13646 (N_13646,N_13116,N_13134);
nand U13647 (N_13647,N_13374,N_13021);
nor U13648 (N_13648,N_13396,N_13036);
xor U13649 (N_13649,N_13296,N_13105);
xnor U13650 (N_13650,N_13237,N_13492);
nor U13651 (N_13651,N_13128,N_13466);
nand U13652 (N_13652,N_13146,N_13034);
and U13653 (N_13653,N_13317,N_13073);
nor U13654 (N_13654,N_13173,N_13323);
xnor U13655 (N_13655,N_13277,N_13072);
and U13656 (N_13656,N_13343,N_13052);
xnor U13657 (N_13657,N_13189,N_13209);
nand U13658 (N_13658,N_13026,N_13147);
nand U13659 (N_13659,N_13085,N_13487);
nand U13660 (N_13660,N_13212,N_13255);
and U13661 (N_13661,N_13130,N_13234);
nand U13662 (N_13662,N_13059,N_13401);
or U13663 (N_13663,N_13049,N_13139);
nor U13664 (N_13664,N_13494,N_13390);
nand U13665 (N_13665,N_13439,N_13462);
nand U13666 (N_13666,N_13151,N_13297);
nor U13667 (N_13667,N_13246,N_13196);
and U13668 (N_13668,N_13123,N_13244);
or U13669 (N_13669,N_13252,N_13086);
or U13670 (N_13670,N_13247,N_13214);
nand U13671 (N_13671,N_13493,N_13226);
and U13672 (N_13672,N_13391,N_13322);
nand U13673 (N_13673,N_13319,N_13415);
nand U13674 (N_13674,N_13032,N_13097);
and U13675 (N_13675,N_13309,N_13037);
and U13676 (N_13676,N_13313,N_13375);
or U13677 (N_13677,N_13114,N_13014);
nor U13678 (N_13678,N_13109,N_13478);
or U13679 (N_13679,N_13093,N_13065);
or U13680 (N_13680,N_13219,N_13111);
nand U13681 (N_13681,N_13445,N_13285);
nor U13682 (N_13682,N_13471,N_13003);
or U13683 (N_13683,N_13485,N_13420);
nor U13684 (N_13684,N_13104,N_13229);
nor U13685 (N_13685,N_13314,N_13334);
nand U13686 (N_13686,N_13267,N_13428);
nor U13687 (N_13687,N_13201,N_13062);
and U13688 (N_13688,N_13424,N_13444);
or U13689 (N_13689,N_13161,N_13175);
nor U13690 (N_13690,N_13169,N_13013);
nand U13691 (N_13691,N_13029,N_13332);
nand U13692 (N_13692,N_13389,N_13235);
or U13693 (N_13693,N_13327,N_13241);
nand U13694 (N_13694,N_13416,N_13378);
xor U13695 (N_13695,N_13242,N_13185);
or U13696 (N_13696,N_13421,N_13184);
nor U13697 (N_13697,N_13430,N_13283);
xnor U13698 (N_13698,N_13305,N_13394);
xnor U13699 (N_13699,N_13482,N_13398);
xor U13700 (N_13700,N_13433,N_13361);
nor U13701 (N_13701,N_13015,N_13359);
or U13702 (N_13702,N_13395,N_13016);
nand U13703 (N_13703,N_13291,N_13187);
xnor U13704 (N_13704,N_13354,N_13180);
nor U13705 (N_13705,N_13012,N_13379);
nand U13706 (N_13706,N_13190,N_13387);
nor U13707 (N_13707,N_13171,N_13091);
or U13708 (N_13708,N_13371,N_13039);
nand U13709 (N_13709,N_13100,N_13117);
nor U13710 (N_13710,N_13061,N_13381);
and U13711 (N_13711,N_13058,N_13101);
nand U13712 (N_13712,N_13355,N_13302);
and U13713 (N_13713,N_13253,N_13258);
or U13714 (N_13714,N_13367,N_13024);
and U13715 (N_13715,N_13172,N_13446);
xnor U13716 (N_13716,N_13276,N_13094);
or U13717 (N_13717,N_13272,N_13233);
or U13718 (N_13718,N_13364,N_13404);
nand U13719 (N_13719,N_13353,N_13070);
and U13720 (N_13720,N_13460,N_13331);
xor U13721 (N_13721,N_13350,N_13360);
or U13722 (N_13722,N_13495,N_13066);
nor U13723 (N_13723,N_13436,N_13138);
xor U13724 (N_13724,N_13330,N_13006);
nor U13725 (N_13725,N_13414,N_13079);
nor U13726 (N_13726,N_13377,N_13256);
or U13727 (N_13727,N_13092,N_13417);
nor U13728 (N_13728,N_13380,N_13270);
nor U13729 (N_13729,N_13316,N_13345);
xnor U13730 (N_13730,N_13249,N_13339);
nand U13731 (N_13731,N_13251,N_13431);
nor U13732 (N_13732,N_13405,N_13167);
xnor U13733 (N_13733,N_13365,N_13307);
or U13734 (N_13734,N_13269,N_13011);
nand U13735 (N_13735,N_13318,N_13124);
xor U13736 (N_13736,N_13088,N_13121);
and U13737 (N_13737,N_13260,N_13239);
and U13738 (N_13738,N_13397,N_13200);
xnor U13739 (N_13739,N_13018,N_13300);
nor U13740 (N_13740,N_13148,N_13425);
and U13741 (N_13741,N_13081,N_13228);
nor U13742 (N_13742,N_13268,N_13041);
xnor U13743 (N_13743,N_13352,N_13453);
xor U13744 (N_13744,N_13437,N_13098);
or U13745 (N_13745,N_13206,N_13090);
or U13746 (N_13746,N_13435,N_13022);
or U13747 (N_13747,N_13250,N_13294);
and U13748 (N_13748,N_13211,N_13231);
and U13749 (N_13749,N_13264,N_13067);
and U13750 (N_13750,N_13024,N_13147);
or U13751 (N_13751,N_13274,N_13367);
and U13752 (N_13752,N_13284,N_13045);
xor U13753 (N_13753,N_13373,N_13321);
and U13754 (N_13754,N_13234,N_13133);
or U13755 (N_13755,N_13049,N_13458);
xor U13756 (N_13756,N_13069,N_13133);
nand U13757 (N_13757,N_13498,N_13190);
nand U13758 (N_13758,N_13313,N_13000);
and U13759 (N_13759,N_13224,N_13246);
xnor U13760 (N_13760,N_13008,N_13241);
nor U13761 (N_13761,N_13029,N_13092);
xnor U13762 (N_13762,N_13330,N_13029);
nor U13763 (N_13763,N_13488,N_13381);
or U13764 (N_13764,N_13062,N_13078);
xnor U13765 (N_13765,N_13256,N_13404);
nor U13766 (N_13766,N_13116,N_13426);
and U13767 (N_13767,N_13376,N_13151);
nor U13768 (N_13768,N_13247,N_13153);
xnor U13769 (N_13769,N_13123,N_13049);
nand U13770 (N_13770,N_13203,N_13164);
nor U13771 (N_13771,N_13163,N_13211);
or U13772 (N_13772,N_13337,N_13375);
or U13773 (N_13773,N_13089,N_13314);
nand U13774 (N_13774,N_13342,N_13465);
and U13775 (N_13775,N_13164,N_13391);
xnor U13776 (N_13776,N_13074,N_13076);
nand U13777 (N_13777,N_13155,N_13481);
nor U13778 (N_13778,N_13369,N_13426);
nor U13779 (N_13779,N_13393,N_13088);
and U13780 (N_13780,N_13467,N_13418);
or U13781 (N_13781,N_13097,N_13375);
xor U13782 (N_13782,N_13347,N_13210);
and U13783 (N_13783,N_13144,N_13299);
and U13784 (N_13784,N_13219,N_13472);
and U13785 (N_13785,N_13104,N_13331);
and U13786 (N_13786,N_13411,N_13341);
and U13787 (N_13787,N_13180,N_13261);
or U13788 (N_13788,N_13166,N_13270);
and U13789 (N_13789,N_13317,N_13306);
or U13790 (N_13790,N_13461,N_13451);
nand U13791 (N_13791,N_13345,N_13035);
xor U13792 (N_13792,N_13254,N_13173);
nand U13793 (N_13793,N_13069,N_13296);
nor U13794 (N_13794,N_13039,N_13025);
nand U13795 (N_13795,N_13292,N_13281);
or U13796 (N_13796,N_13263,N_13255);
or U13797 (N_13797,N_13071,N_13102);
and U13798 (N_13798,N_13130,N_13089);
and U13799 (N_13799,N_13331,N_13027);
and U13800 (N_13800,N_13220,N_13469);
xnor U13801 (N_13801,N_13239,N_13295);
nand U13802 (N_13802,N_13068,N_13223);
or U13803 (N_13803,N_13245,N_13420);
or U13804 (N_13804,N_13135,N_13012);
nor U13805 (N_13805,N_13422,N_13116);
nor U13806 (N_13806,N_13462,N_13089);
xnor U13807 (N_13807,N_13347,N_13434);
nand U13808 (N_13808,N_13051,N_13116);
or U13809 (N_13809,N_13353,N_13295);
xor U13810 (N_13810,N_13180,N_13229);
nand U13811 (N_13811,N_13122,N_13220);
nand U13812 (N_13812,N_13344,N_13121);
xor U13813 (N_13813,N_13424,N_13366);
or U13814 (N_13814,N_13490,N_13406);
nand U13815 (N_13815,N_13231,N_13294);
and U13816 (N_13816,N_13404,N_13200);
nor U13817 (N_13817,N_13460,N_13201);
nor U13818 (N_13818,N_13451,N_13298);
nand U13819 (N_13819,N_13193,N_13489);
nor U13820 (N_13820,N_13053,N_13344);
or U13821 (N_13821,N_13202,N_13403);
nor U13822 (N_13822,N_13402,N_13230);
nand U13823 (N_13823,N_13285,N_13474);
xor U13824 (N_13824,N_13324,N_13418);
or U13825 (N_13825,N_13257,N_13275);
nand U13826 (N_13826,N_13327,N_13320);
and U13827 (N_13827,N_13489,N_13401);
and U13828 (N_13828,N_13457,N_13159);
nand U13829 (N_13829,N_13051,N_13351);
nor U13830 (N_13830,N_13329,N_13472);
or U13831 (N_13831,N_13400,N_13262);
or U13832 (N_13832,N_13280,N_13166);
and U13833 (N_13833,N_13359,N_13412);
nand U13834 (N_13834,N_13105,N_13298);
and U13835 (N_13835,N_13490,N_13017);
or U13836 (N_13836,N_13424,N_13298);
xnor U13837 (N_13837,N_13149,N_13174);
xnor U13838 (N_13838,N_13090,N_13212);
xnor U13839 (N_13839,N_13247,N_13178);
nor U13840 (N_13840,N_13094,N_13444);
xnor U13841 (N_13841,N_13145,N_13265);
or U13842 (N_13842,N_13173,N_13118);
nand U13843 (N_13843,N_13063,N_13382);
xnor U13844 (N_13844,N_13249,N_13483);
xnor U13845 (N_13845,N_13043,N_13003);
xnor U13846 (N_13846,N_13379,N_13000);
xnor U13847 (N_13847,N_13357,N_13051);
nand U13848 (N_13848,N_13140,N_13298);
xor U13849 (N_13849,N_13063,N_13089);
and U13850 (N_13850,N_13085,N_13060);
or U13851 (N_13851,N_13437,N_13128);
and U13852 (N_13852,N_13408,N_13458);
nand U13853 (N_13853,N_13137,N_13435);
xnor U13854 (N_13854,N_13267,N_13495);
nor U13855 (N_13855,N_13333,N_13403);
or U13856 (N_13856,N_13026,N_13229);
or U13857 (N_13857,N_13414,N_13472);
or U13858 (N_13858,N_13145,N_13242);
and U13859 (N_13859,N_13028,N_13361);
nand U13860 (N_13860,N_13290,N_13261);
and U13861 (N_13861,N_13144,N_13005);
xor U13862 (N_13862,N_13351,N_13079);
nand U13863 (N_13863,N_13043,N_13014);
xor U13864 (N_13864,N_13134,N_13437);
nand U13865 (N_13865,N_13035,N_13101);
xnor U13866 (N_13866,N_13358,N_13202);
nand U13867 (N_13867,N_13179,N_13212);
nor U13868 (N_13868,N_13160,N_13297);
nor U13869 (N_13869,N_13102,N_13164);
nand U13870 (N_13870,N_13073,N_13479);
or U13871 (N_13871,N_13428,N_13072);
or U13872 (N_13872,N_13021,N_13378);
nand U13873 (N_13873,N_13304,N_13008);
or U13874 (N_13874,N_13097,N_13078);
and U13875 (N_13875,N_13473,N_13264);
nor U13876 (N_13876,N_13417,N_13211);
or U13877 (N_13877,N_13489,N_13247);
xor U13878 (N_13878,N_13414,N_13312);
and U13879 (N_13879,N_13172,N_13352);
nand U13880 (N_13880,N_13482,N_13368);
and U13881 (N_13881,N_13358,N_13339);
and U13882 (N_13882,N_13425,N_13068);
nand U13883 (N_13883,N_13489,N_13079);
or U13884 (N_13884,N_13492,N_13306);
nor U13885 (N_13885,N_13170,N_13400);
nand U13886 (N_13886,N_13226,N_13319);
nor U13887 (N_13887,N_13002,N_13054);
nor U13888 (N_13888,N_13099,N_13089);
or U13889 (N_13889,N_13302,N_13001);
nor U13890 (N_13890,N_13023,N_13092);
nand U13891 (N_13891,N_13370,N_13229);
or U13892 (N_13892,N_13024,N_13463);
nand U13893 (N_13893,N_13058,N_13370);
nor U13894 (N_13894,N_13015,N_13068);
xnor U13895 (N_13895,N_13370,N_13134);
or U13896 (N_13896,N_13040,N_13210);
and U13897 (N_13897,N_13078,N_13205);
and U13898 (N_13898,N_13422,N_13188);
or U13899 (N_13899,N_13138,N_13131);
and U13900 (N_13900,N_13203,N_13190);
or U13901 (N_13901,N_13354,N_13492);
xor U13902 (N_13902,N_13263,N_13259);
xnor U13903 (N_13903,N_13409,N_13313);
nand U13904 (N_13904,N_13314,N_13290);
xnor U13905 (N_13905,N_13092,N_13180);
xor U13906 (N_13906,N_13442,N_13081);
and U13907 (N_13907,N_13224,N_13101);
nand U13908 (N_13908,N_13201,N_13069);
or U13909 (N_13909,N_13350,N_13492);
and U13910 (N_13910,N_13390,N_13057);
xor U13911 (N_13911,N_13098,N_13040);
nand U13912 (N_13912,N_13370,N_13084);
or U13913 (N_13913,N_13070,N_13389);
xor U13914 (N_13914,N_13191,N_13389);
nor U13915 (N_13915,N_13327,N_13138);
nand U13916 (N_13916,N_13159,N_13153);
nor U13917 (N_13917,N_13019,N_13300);
nor U13918 (N_13918,N_13290,N_13486);
or U13919 (N_13919,N_13218,N_13419);
or U13920 (N_13920,N_13367,N_13429);
and U13921 (N_13921,N_13076,N_13447);
nand U13922 (N_13922,N_13043,N_13155);
nor U13923 (N_13923,N_13499,N_13083);
and U13924 (N_13924,N_13191,N_13304);
nand U13925 (N_13925,N_13459,N_13423);
nor U13926 (N_13926,N_13000,N_13155);
or U13927 (N_13927,N_13351,N_13122);
nand U13928 (N_13928,N_13168,N_13009);
xor U13929 (N_13929,N_13166,N_13215);
nor U13930 (N_13930,N_13434,N_13468);
nand U13931 (N_13931,N_13484,N_13083);
or U13932 (N_13932,N_13327,N_13389);
and U13933 (N_13933,N_13019,N_13011);
or U13934 (N_13934,N_13175,N_13258);
nor U13935 (N_13935,N_13359,N_13468);
xnor U13936 (N_13936,N_13175,N_13435);
nand U13937 (N_13937,N_13082,N_13372);
xnor U13938 (N_13938,N_13346,N_13398);
nor U13939 (N_13939,N_13021,N_13138);
or U13940 (N_13940,N_13333,N_13094);
or U13941 (N_13941,N_13410,N_13286);
or U13942 (N_13942,N_13461,N_13407);
or U13943 (N_13943,N_13079,N_13259);
nor U13944 (N_13944,N_13190,N_13188);
and U13945 (N_13945,N_13223,N_13255);
and U13946 (N_13946,N_13447,N_13408);
xor U13947 (N_13947,N_13460,N_13253);
xor U13948 (N_13948,N_13294,N_13077);
nand U13949 (N_13949,N_13002,N_13435);
or U13950 (N_13950,N_13204,N_13096);
nand U13951 (N_13951,N_13173,N_13281);
xor U13952 (N_13952,N_13413,N_13327);
xor U13953 (N_13953,N_13046,N_13380);
xnor U13954 (N_13954,N_13263,N_13148);
or U13955 (N_13955,N_13192,N_13243);
and U13956 (N_13956,N_13299,N_13119);
and U13957 (N_13957,N_13256,N_13248);
and U13958 (N_13958,N_13184,N_13488);
nand U13959 (N_13959,N_13087,N_13165);
nor U13960 (N_13960,N_13330,N_13281);
and U13961 (N_13961,N_13480,N_13224);
nor U13962 (N_13962,N_13299,N_13060);
xnor U13963 (N_13963,N_13245,N_13218);
nand U13964 (N_13964,N_13450,N_13391);
xor U13965 (N_13965,N_13394,N_13380);
and U13966 (N_13966,N_13027,N_13274);
and U13967 (N_13967,N_13094,N_13185);
xnor U13968 (N_13968,N_13406,N_13246);
and U13969 (N_13969,N_13109,N_13195);
nor U13970 (N_13970,N_13092,N_13022);
and U13971 (N_13971,N_13479,N_13371);
or U13972 (N_13972,N_13050,N_13036);
or U13973 (N_13973,N_13440,N_13217);
nand U13974 (N_13974,N_13394,N_13108);
and U13975 (N_13975,N_13329,N_13066);
xor U13976 (N_13976,N_13002,N_13164);
xor U13977 (N_13977,N_13170,N_13153);
nor U13978 (N_13978,N_13365,N_13259);
xor U13979 (N_13979,N_13432,N_13149);
nor U13980 (N_13980,N_13241,N_13103);
or U13981 (N_13981,N_13274,N_13353);
nand U13982 (N_13982,N_13001,N_13449);
or U13983 (N_13983,N_13364,N_13131);
and U13984 (N_13984,N_13248,N_13301);
nand U13985 (N_13985,N_13494,N_13059);
xor U13986 (N_13986,N_13220,N_13219);
or U13987 (N_13987,N_13472,N_13121);
xnor U13988 (N_13988,N_13416,N_13203);
or U13989 (N_13989,N_13482,N_13388);
nand U13990 (N_13990,N_13476,N_13173);
nand U13991 (N_13991,N_13137,N_13058);
or U13992 (N_13992,N_13434,N_13305);
nand U13993 (N_13993,N_13430,N_13052);
and U13994 (N_13994,N_13050,N_13401);
or U13995 (N_13995,N_13427,N_13020);
or U13996 (N_13996,N_13004,N_13189);
xnor U13997 (N_13997,N_13004,N_13425);
nand U13998 (N_13998,N_13045,N_13152);
and U13999 (N_13999,N_13412,N_13361);
or U14000 (N_14000,N_13830,N_13531);
or U14001 (N_14001,N_13690,N_13905);
or U14002 (N_14002,N_13628,N_13934);
xor U14003 (N_14003,N_13778,N_13665);
or U14004 (N_14004,N_13896,N_13655);
or U14005 (N_14005,N_13977,N_13634);
nand U14006 (N_14006,N_13647,N_13715);
or U14007 (N_14007,N_13734,N_13959);
xor U14008 (N_14008,N_13803,N_13857);
xnor U14009 (N_14009,N_13699,N_13917);
nor U14010 (N_14010,N_13923,N_13975);
or U14011 (N_14011,N_13632,N_13595);
nand U14012 (N_14012,N_13853,N_13572);
nand U14013 (N_14013,N_13709,N_13992);
or U14014 (N_14014,N_13805,N_13854);
xor U14015 (N_14015,N_13955,N_13593);
xor U14016 (N_14016,N_13944,N_13991);
xnor U14017 (N_14017,N_13826,N_13693);
xnor U14018 (N_14018,N_13639,N_13621);
or U14019 (N_14019,N_13600,N_13579);
nand U14020 (N_14020,N_13984,N_13653);
nand U14021 (N_14021,N_13766,N_13849);
or U14022 (N_14022,N_13672,N_13696);
or U14023 (N_14023,N_13914,N_13569);
or U14024 (N_14024,N_13719,N_13759);
nand U14025 (N_14025,N_13868,N_13526);
nor U14026 (N_14026,N_13535,N_13506);
or U14027 (N_14027,N_13987,N_13815);
or U14028 (N_14028,N_13701,N_13596);
or U14029 (N_14029,N_13521,N_13687);
xor U14030 (N_14030,N_13666,N_13844);
or U14031 (N_14031,N_13798,N_13697);
xnor U14032 (N_14032,N_13897,N_13786);
nor U14033 (N_14033,N_13771,N_13675);
and U14034 (N_14034,N_13942,N_13883);
and U14035 (N_14035,N_13983,N_13601);
nor U14036 (N_14036,N_13641,N_13587);
xor U14037 (N_14037,N_13500,N_13549);
xor U14038 (N_14038,N_13554,N_13918);
nor U14039 (N_14039,N_13507,N_13631);
or U14040 (N_14040,N_13817,N_13524);
and U14041 (N_14041,N_13866,N_13793);
and U14042 (N_14042,N_13517,N_13941);
xor U14043 (N_14043,N_13671,N_13843);
or U14044 (N_14044,N_13971,N_13643);
or U14045 (N_14045,N_13740,N_13969);
nor U14046 (N_14046,N_13527,N_13910);
xor U14047 (N_14047,N_13575,N_13774);
nand U14048 (N_14048,N_13662,N_13656);
nor U14049 (N_14049,N_13891,N_13860);
xor U14050 (N_14050,N_13960,N_13988);
and U14051 (N_14051,N_13764,N_13967);
or U14052 (N_14052,N_13856,N_13961);
xnor U14053 (N_14053,N_13512,N_13953);
xor U14054 (N_14054,N_13552,N_13795);
nand U14055 (N_14055,N_13839,N_13725);
nor U14056 (N_14056,N_13629,N_13946);
nor U14057 (N_14057,N_13926,N_13543);
nand U14058 (N_14058,N_13576,N_13728);
xnor U14059 (N_14059,N_13878,N_13541);
nand U14060 (N_14060,N_13824,N_13776);
and U14061 (N_14061,N_13516,N_13872);
or U14062 (N_14062,N_13850,N_13851);
or U14063 (N_14063,N_13819,N_13772);
and U14064 (N_14064,N_13838,N_13545);
and U14065 (N_14065,N_13762,N_13695);
or U14066 (N_14066,N_13511,N_13842);
xor U14067 (N_14067,N_13870,N_13752);
or U14068 (N_14068,N_13846,N_13790);
nand U14069 (N_14069,N_13783,N_13540);
or U14070 (N_14070,N_13723,N_13779);
or U14071 (N_14071,N_13927,N_13761);
and U14072 (N_14072,N_13547,N_13722);
xnor U14073 (N_14073,N_13879,N_13586);
or U14074 (N_14074,N_13823,N_13729);
or U14075 (N_14075,N_13726,N_13845);
and U14076 (N_14076,N_13704,N_13997);
xnor U14077 (N_14077,N_13881,N_13518);
or U14078 (N_14078,N_13882,N_13706);
and U14079 (N_14079,N_13788,N_13996);
and U14080 (N_14080,N_13939,N_13974);
xnor U14081 (N_14081,N_13806,N_13737);
nand U14082 (N_14082,N_13710,N_13749);
and U14083 (N_14083,N_13591,N_13683);
and U14084 (N_14084,N_13618,N_13694);
nor U14085 (N_14085,N_13686,N_13711);
and U14086 (N_14086,N_13787,N_13980);
nand U14087 (N_14087,N_13570,N_13863);
and U14088 (N_14088,N_13829,N_13519);
or U14089 (N_14089,N_13898,N_13998);
and U14090 (N_14090,N_13566,N_13963);
nor U14091 (N_14091,N_13670,N_13667);
or U14092 (N_14092,N_13804,N_13911);
or U14093 (N_14093,N_13877,N_13612);
nand U14094 (N_14094,N_13950,N_13724);
and U14095 (N_14095,N_13802,N_13943);
or U14096 (N_14096,N_13584,N_13920);
or U14097 (N_14097,N_13964,N_13677);
or U14098 (N_14098,N_13782,N_13522);
or U14099 (N_14099,N_13907,N_13609);
or U14100 (N_14100,N_13949,N_13604);
and U14101 (N_14101,N_13864,N_13659);
nor U14102 (N_14102,N_13716,N_13718);
xor U14103 (N_14103,N_13550,N_13590);
nor U14104 (N_14104,N_13505,N_13936);
and U14105 (N_14105,N_13698,N_13816);
xnor U14106 (N_14106,N_13742,N_13820);
or U14107 (N_14107,N_13513,N_13906);
or U14108 (N_14108,N_13909,N_13965);
nand U14109 (N_14109,N_13747,N_13525);
nor U14110 (N_14110,N_13504,N_13739);
or U14111 (N_14111,N_13674,N_13865);
nand U14112 (N_14112,N_13578,N_13876);
nand U14113 (N_14113,N_13720,N_13780);
or U14114 (N_14114,N_13688,N_13784);
and U14115 (N_14115,N_13637,N_13733);
or U14116 (N_14116,N_13919,N_13627);
xor U14117 (N_14117,N_13753,N_13777);
and U14118 (N_14118,N_13731,N_13962);
nor U14119 (N_14119,N_13714,N_13937);
nand U14120 (N_14120,N_13903,N_13581);
nand U14121 (N_14121,N_13954,N_13567);
xor U14122 (N_14122,N_13592,N_13822);
nor U14123 (N_14123,N_13808,N_13561);
xor U14124 (N_14124,N_13616,N_13553);
and U14125 (N_14125,N_13681,N_13821);
xnor U14126 (N_14126,N_13833,N_13745);
nand U14127 (N_14127,N_13892,N_13555);
xor U14128 (N_14128,N_13705,N_13855);
xor U14129 (N_14129,N_13649,N_13976);
xnor U14130 (N_14130,N_13945,N_13743);
nor U14131 (N_14131,N_13862,N_13536);
or U14132 (N_14132,N_13573,N_13995);
xor U14133 (N_14133,N_13556,N_13982);
xnor U14134 (N_14134,N_13924,N_13620);
xor U14135 (N_14135,N_13814,N_13800);
and U14136 (N_14136,N_13588,N_13758);
or U14137 (N_14137,N_13712,N_13885);
or U14138 (N_14138,N_13594,N_13861);
nand U14139 (N_14139,N_13895,N_13811);
nand U14140 (N_14140,N_13931,N_13682);
nor U14141 (N_14141,N_13773,N_13608);
or U14142 (N_14142,N_13626,N_13951);
nand U14143 (N_14143,N_13801,N_13617);
or U14144 (N_14144,N_13700,N_13769);
xnor U14145 (N_14145,N_13548,N_13900);
nor U14146 (N_14146,N_13757,N_13669);
and U14147 (N_14147,N_13673,N_13970);
or U14148 (N_14148,N_13832,N_13533);
xor U14149 (N_14149,N_13692,N_13599);
nor U14150 (N_14150,N_13871,N_13538);
nor U14151 (N_14151,N_13929,N_13889);
nand U14152 (N_14152,N_13580,N_13940);
or U14153 (N_14153,N_13508,N_13520);
nor U14154 (N_14154,N_13582,N_13828);
xnor U14155 (N_14155,N_13990,N_13624);
and U14156 (N_14156,N_13933,N_13981);
and U14157 (N_14157,N_13651,N_13558);
nor U14158 (N_14158,N_13565,N_13867);
nor U14159 (N_14159,N_13791,N_13792);
xor U14160 (N_14160,N_13568,N_13614);
and U14161 (N_14161,N_13563,N_13721);
nor U14162 (N_14162,N_13652,N_13703);
and U14163 (N_14163,N_13679,N_13754);
nand U14164 (N_14164,N_13751,N_13661);
nor U14165 (N_14165,N_13585,N_13775);
xor U14166 (N_14166,N_13503,N_13730);
and U14167 (N_14167,N_13858,N_13921);
and U14168 (N_14168,N_13502,N_13736);
and U14169 (N_14169,N_13534,N_13848);
and U14170 (N_14170,N_13571,N_13989);
and U14171 (N_14171,N_13557,N_13765);
xor U14172 (N_14172,N_13886,N_13646);
xnor U14173 (N_14173,N_13630,N_13979);
nand U14174 (N_14174,N_13603,N_13544);
xnor U14175 (N_14175,N_13794,N_13922);
nor U14176 (N_14176,N_13689,N_13741);
and U14177 (N_14177,N_13529,N_13657);
nand U14178 (N_14178,N_13625,N_13873);
nor U14179 (N_14179,N_13606,N_13605);
nand U14180 (N_14180,N_13781,N_13537);
xor U14181 (N_14181,N_13551,N_13515);
nor U14182 (N_14182,N_13812,N_13702);
xor U14183 (N_14183,N_13859,N_13654);
nand U14184 (N_14184,N_13915,N_13648);
xnor U14185 (N_14185,N_13999,N_13642);
and U14186 (N_14186,N_13589,N_13622);
nor U14187 (N_14187,N_13875,N_13887);
nand U14188 (N_14188,N_13899,N_13952);
nor U14189 (N_14189,N_13756,N_13658);
and U14190 (N_14190,N_13660,N_13707);
and U14191 (N_14191,N_13874,N_13528);
nor U14192 (N_14192,N_13501,N_13560);
nor U14193 (N_14193,N_13836,N_13638);
and U14194 (N_14194,N_13746,N_13650);
nand U14195 (N_14195,N_13869,N_13768);
nor U14196 (N_14196,N_13676,N_13912);
and U14197 (N_14197,N_13831,N_13904);
or U14198 (N_14198,N_13750,N_13532);
or U14199 (N_14199,N_13957,N_13744);
and U14200 (N_14200,N_13623,N_13763);
and U14201 (N_14201,N_13938,N_13956);
xor U14202 (N_14202,N_13713,N_13785);
or U14203 (N_14203,N_13925,N_13837);
nand U14204 (N_14204,N_13559,N_13841);
xnor U14205 (N_14205,N_13796,N_13583);
or U14206 (N_14206,N_13748,N_13691);
nand U14207 (N_14207,N_13635,N_13884);
or U14208 (N_14208,N_13901,N_13664);
and U14209 (N_14209,N_13607,N_13644);
and U14210 (N_14210,N_13993,N_13932);
xnor U14211 (N_14211,N_13770,N_13827);
nand U14212 (N_14212,N_13902,N_13678);
xnor U14213 (N_14213,N_13735,N_13523);
or U14214 (N_14214,N_13640,N_13994);
xor U14215 (N_14215,N_13514,N_13893);
or U14216 (N_14216,N_13930,N_13813);
nand U14217 (N_14217,N_13680,N_13546);
nand U14218 (N_14218,N_13966,N_13880);
and U14219 (N_14219,N_13958,N_13789);
xor U14220 (N_14220,N_13530,N_13978);
and U14221 (N_14221,N_13825,N_13986);
nor U14222 (N_14222,N_13968,N_13755);
and U14223 (N_14223,N_13809,N_13913);
nor U14224 (N_14224,N_13539,N_13928);
xor U14225 (N_14225,N_13717,N_13542);
xor U14226 (N_14226,N_13973,N_13810);
xnor U14227 (N_14227,N_13972,N_13611);
xnor U14228 (N_14228,N_13615,N_13847);
xnor U14229 (N_14229,N_13947,N_13835);
and U14230 (N_14230,N_13510,N_13916);
nor U14231 (N_14231,N_13509,N_13797);
xor U14232 (N_14232,N_13807,N_13818);
and U14233 (N_14233,N_13935,N_13613);
nor U14234 (N_14234,N_13834,N_13799);
and U14235 (N_14235,N_13732,N_13767);
xor U14236 (N_14236,N_13852,N_13738);
and U14237 (N_14237,N_13685,N_13663);
or U14238 (N_14238,N_13840,N_13610);
xor U14239 (N_14239,N_13708,N_13597);
xnor U14240 (N_14240,N_13985,N_13684);
nor U14241 (N_14241,N_13602,N_13948);
nand U14242 (N_14242,N_13727,N_13619);
nor U14243 (N_14243,N_13562,N_13888);
nand U14244 (N_14244,N_13598,N_13564);
nand U14245 (N_14245,N_13577,N_13633);
nand U14246 (N_14246,N_13908,N_13668);
and U14247 (N_14247,N_13574,N_13645);
or U14248 (N_14248,N_13636,N_13894);
and U14249 (N_14249,N_13890,N_13760);
or U14250 (N_14250,N_13604,N_13592);
and U14251 (N_14251,N_13556,N_13844);
nor U14252 (N_14252,N_13882,N_13976);
or U14253 (N_14253,N_13859,N_13727);
nand U14254 (N_14254,N_13584,N_13884);
nor U14255 (N_14255,N_13576,N_13951);
xor U14256 (N_14256,N_13827,N_13823);
and U14257 (N_14257,N_13557,N_13758);
nor U14258 (N_14258,N_13969,N_13812);
xnor U14259 (N_14259,N_13770,N_13566);
nor U14260 (N_14260,N_13947,N_13861);
nor U14261 (N_14261,N_13580,N_13784);
and U14262 (N_14262,N_13816,N_13919);
nor U14263 (N_14263,N_13570,N_13780);
xnor U14264 (N_14264,N_13772,N_13986);
nor U14265 (N_14265,N_13949,N_13854);
xor U14266 (N_14266,N_13755,N_13764);
nor U14267 (N_14267,N_13591,N_13563);
xor U14268 (N_14268,N_13560,N_13650);
nand U14269 (N_14269,N_13690,N_13811);
xor U14270 (N_14270,N_13723,N_13972);
xor U14271 (N_14271,N_13587,N_13755);
xor U14272 (N_14272,N_13701,N_13562);
nor U14273 (N_14273,N_13993,N_13669);
or U14274 (N_14274,N_13693,N_13715);
or U14275 (N_14275,N_13764,N_13948);
xnor U14276 (N_14276,N_13893,N_13892);
nor U14277 (N_14277,N_13888,N_13598);
xor U14278 (N_14278,N_13815,N_13640);
and U14279 (N_14279,N_13912,N_13838);
xor U14280 (N_14280,N_13946,N_13885);
or U14281 (N_14281,N_13661,N_13730);
xor U14282 (N_14282,N_13590,N_13945);
and U14283 (N_14283,N_13504,N_13592);
nand U14284 (N_14284,N_13770,N_13974);
xnor U14285 (N_14285,N_13516,N_13623);
nor U14286 (N_14286,N_13522,N_13739);
xnor U14287 (N_14287,N_13959,N_13813);
xor U14288 (N_14288,N_13893,N_13820);
or U14289 (N_14289,N_13546,N_13883);
nand U14290 (N_14290,N_13592,N_13941);
and U14291 (N_14291,N_13951,N_13770);
xnor U14292 (N_14292,N_13909,N_13837);
and U14293 (N_14293,N_13925,N_13737);
nor U14294 (N_14294,N_13823,N_13601);
xnor U14295 (N_14295,N_13655,N_13514);
or U14296 (N_14296,N_13883,N_13559);
nand U14297 (N_14297,N_13654,N_13870);
or U14298 (N_14298,N_13543,N_13548);
or U14299 (N_14299,N_13569,N_13887);
or U14300 (N_14300,N_13716,N_13610);
or U14301 (N_14301,N_13911,N_13873);
nand U14302 (N_14302,N_13569,N_13617);
xor U14303 (N_14303,N_13909,N_13545);
or U14304 (N_14304,N_13546,N_13953);
or U14305 (N_14305,N_13963,N_13873);
xor U14306 (N_14306,N_13822,N_13890);
and U14307 (N_14307,N_13745,N_13703);
and U14308 (N_14308,N_13815,N_13923);
or U14309 (N_14309,N_13980,N_13703);
nor U14310 (N_14310,N_13573,N_13716);
and U14311 (N_14311,N_13533,N_13617);
xnor U14312 (N_14312,N_13964,N_13968);
nand U14313 (N_14313,N_13995,N_13561);
nor U14314 (N_14314,N_13716,N_13710);
nor U14315 (N_14315,N_13623,N_13819);
xor U14316 (N_14316,N_13899,N_13659);
nor U14317 (N_14317,N_13597,N_13923);
nor U14318 (N_14318,N_13592,N_13994);
nand U14319 (N_14319,N_13859,N_13564);
or U14320 (N_14320,N_13866,N_13950);
nor U14321 (N_14321,N_13885,N_13606);
and U14322 (N_14322,N_13876,N_13639);
and U14323 (N_14323,N_13865,N_13609);
xor U14324 (N_14324,N_13874,N_13568);
or U14325 (N_14325,N_13844,N_13631);
or U14326 (N_14326,N_13660,N_13573);
and U14327 (N_14327,N_13715,N_13906);
and U14328 (N_14328,N_13783,N_13560);
and U14329 (N_14329,N_13675,N_13898);
and U14330 (N_14330,N_13656,N_13686);
xnor U14331 (N_14331,N_13693,N_13558);
or U14332 (N_14332,N_13832,N_13535);
nor U14333 (N_14333,N_13886,N_13843);
or U14334 (N_14334,N_13956,N_13833);
and U14335 (N_14335,N_13694,N_13591);
or U14336 (N_14336,N_13600,N_13741);
or U14337 (N_14337,N_13501,N_13870);
xnor U14338 (N_14338,N_13644,N_13699);
or U14339 (N_14339,N_13945,N_13938);
nor U14340 (N_14340,N_13544,N_13680);
or U14341 (N_14341,N_13758,N_13514);
nand U14342 (N_14342,N_13717,N_13731);
and U14343 (N_14343,N_13642,N_13534);
nand U14344 (N_14344,N_13664,N_13619);
and U14345 (N_14345,N_13951,N_13747);
or U14346 (N_14346,N_13521,N_13641);
or U14347 (N_14347,N_13846,N_13801);
nor U14348 (N_14348,N_13625,N_13728);
xor U14349 (N_14349,N_13582,N_13930);
xor U14350 (N_14350,N_13905,N_13831);
nor U14351 (N_14351,N_13983,N_13740);
nand U14352 (N_14352,N_13717,N_13870);
xnor U14353 (N_14353,N_13909,N_13615);
nand U14354 (N_14354,N_13950,N_13845);
xnor U14355 (N_14355,N_13576,N_13899);
and U14356 (N_14356,N_13981,N_13765);
or U14357 (N_14357,N_13779,N_13928);
xor U14358 (N_14358,N_13831,N_13833);
nor U14359 (N_14359,N_13557,N_13787);
xor U14360 (N_14360,N_13813,N_13769);
and U14361 (N_14361,N_13837,N_13689);
xor U14362 (N_14362,N_13639,N_13799);
and U14363 (N_14363,N_13635,N_13737);
xnor U14364 (N_14364,N_13977,N_13924);
nor U14365 (N_14365,N_13668,N_13819);
xor U14366 (N_14366,N_13864,N_13757);
nor U14367 (N_14367,N_13512,N_13547);
nor U14368 (N_14368,N_13663,N_13561);
or U14369 (N_14369,N_13697,N_13550);
and U14370 (N_14370,N_13641,N_13992);
nand U14371 (N_14371,N_13952,N_13696);
and U14372 (N_14372,N_13568,N_13977);
nor U14373 (N_14373,N_13800,N_13576);
and U14374 (N_14374,N_13890,N_13893);
and U14375 (N_14375,N_13618,N_13578);
nand U14376 (N_14376,N_13575,N_13510);
xnor U14377 (N_14377,N_13816,N_13873);
and U14378 (N_14378,N_13540,N_13518);
nor U14379 (N_14379,N_13577,N_13681);
or U14380 (N_14380,N_13658,N_13645);
nand U14381 (N_14381,N_13645,N_13767);
nor U14382 (N_14382,N_13990,N_13780);
and U14383 (N_14383,N_13641,N_13892);
nor U14384 (N_14384,N_13552,N_13775);
nor U14385 (N_14385,N_13951,N_13782);
nor U14386 (N_14386,N_13603,N_13877);
nor U14387 (N_14387,N_13641,N_13888);
nor U14388 (N_14388,N_13747,N_13677);
nand U14389 (N_14389,N_13616,N_13522);
xnor U14390 (N_14390,N_13662,N_13552);
xnor U14391 (N_14391,N_13926,N_13890);
nand U14392 (N_14392,N_13620,N_13713);
and U14393 (N_14393,N_13876,N_13677);
or U14394 (N_14394,N_13861,N_13539);
xor U14395 (N_14395,N_13913,N_13675);
nor U14396 (N_14396,N_13825,N_13864);
and U14397 (N_14397,N_13807,N_13607);
xnor U14398 (N_14398,N_13515,N_13500);
and U14399 (N_14399,N_13561,N_13627);
nand U14400 (N_14400,N_13718,N_13983);
and U14401 (N_14401,N_13858,N_13825);
or U14402 (N_14402,N_13634,N_13655);
xnor U14403 (N_14403,N_13696,N_13572);
or U14404 (N_14404,N_13634,N_13960);
and U14405 (N_14405,N_13837,N_13569);
and U14406 (N_14406,N_13952,N_13995);
nand U14407 (N_14407,N_13773,N_13923);
or U14408 (N_14408,N_13827,N_13637);
and U14409 (N_14409,N_13615,N_13825);
or U14410 (N_14410,N_13856,N_13847);
or U14411 (N_14411,N_13670,N_13930);
and U14412 (N_14412,N_13576,N_13594);
nor U14413 (N_14413,N_13662,N_13801);
nand U14414 (N_14414,N_13641,N_13808);
or U14415 (N_14415,N_13740,N_13857);
and U14416 (N_14416,N_13536,N_13597);
nor U14417 (N_14417,N_13893,N_13803);
xnor U14418 (N_14418,N_13762,N_13685);
nor U14419 (N_14419,N_13622,N_13504);
nand U14420 (N_14420,N_13947,N_13799);
xnor U14421 (N_14421,N_13813,N_13682);
xnor U14422 (N_14422,N_13859,N_13850);
and U14423 (N_14423,N_13503,N_13648);
nor U14424 (N_14424,N_13921,N_13904);
xor U14425 (N_14425,N_13929,N_13907);
xnor U14426 (N_14426,N_13606,N_13786);
nand U14427 (N_14427,N_13917,N_13978);
or U14428 (N_14428,N_13938,N_13988);
nand U14429 (N_14429,N_13901,N_13826);
nor U14430 (N_14430,N_13797,N_13891);
and U14431 (N_14431,N_13693,N_13783);
nor U14432 (N_14432,N_13901,N_13775);
nor U14433 (N_14433,N_13546,N_13716);
nand U14434 (N_14434,N_13645,N_13943);
xnor U14435 (N_14435,N_13779,N_13936);
nand U14436 (N_14436,N_13550,N_13624);
nand U14437 (N_14437,N_13518,N_13977);
nor U14438 (N_14438,N_13667,N_13656);
nand U14439 (N_14439,N_13708,N_13594);
xor U14440 (N_14440,N_13591,N_13819);
and U14441 (N_14441,N_13608,N_13643);
and U14442 (N_14442,N_13979,N_13924);
nand U14443 (N_14443,N_13655,N_13664);
nand U14444 (N_14444,N_13899,N_13632);
nand U14445 (N_14445,N_13716,N_13915);
xnor U14446 (N_14446,N_13671,N_13788);
nor U14447 (N_14447,N_13727,N_13700);
and U14448 (N_14448,N_13568,N_13850);
or U14449 (N_14449,N_13571,N_13898);
xor U14450 (N_14450,N_13503,N_13902);
nor U14451 (N_14451,N_13530,N_13568);
and U14452 (N_14452,N_13500,N_13820);
nand U14453 (N_14453,N_13993,N_13897);
and U14454 (N_14454,N_13662,N_13833);
and U14455 (N_14455,N_13879,N_13652);
or U14456 (N_14456,N_13668,N_13927);
xnor U14457 (N_14457,N_13983,N_13591);
and U14458 (N_14458,N_13767,N_13518);
nand U14459 (N_14459,N_13518,N_13597);
nand U14460 (N_14460,N_13675,N_13684);
xnor U14461 (N_14461,N_13520,N_13929);
and U14462 (N_14462,N_13633,N_13510);
nor U14463 (N_14463,N_13903,N_13583);
and U14464 (N_14464,N_13974,N_13843);
nand U14465 (N_14465,N_13574,N_13862);
nand U14466 (N_14466,N_13695,N_13528);
and U14467 (N_14467,N_13550,N_13545);
nor U14468 (N_14468,N_13567,N_13689);
and U14469 (N_14469,N_13846,N_13859);
xor U14470 (N_14470,N_13648,N_13906);
nand U14471 (N_14471,N_13919,N_13950);
and U14472 (N_14472,N_13867,N_13960);
xor U14473 (N_14473,N_13729,N_13504);
nand U14474 (N_14474,N_13771,N_13536);
xor U14475 (N_14475,N_13813,N_13990);
xnor U14476 (N_14476,N_13962,N_13581);
nand U14477 (N_14477,N_13875,N_13685);
or U14478 (N_14478,N_13773,N_13766);
or U14479 (N_14479,N_13773,N_13565);
nand U14480 (N_14480,N_13948,N_13911);
nand U14481 (N_14481,N_13545,N_13686);
or U14482 (N_14482,N_13997,N_13813);
xnor U14483 (N_14483,N_13503,N_13900);
xor U14484 (N_14484,N_13940,N_13904);
xor U14485 (N_14485,N_13647,N_13609);
nor U14486 (N_14486,N_13544,N_13759);
xor U14487 (N_14487,N_13711,N_13601);
nor U14488 (N_14488,N_13997,N_13798);
nand U14489 (N_14489,N_13581,N_13973);
nand U14490 (N_14490,N_13802,N_13867);
or U14491 (N_14491,N_13845,N_13685);
nor U14492 (N_14492,N_13758,N_13837);
and U14493 (N_14493,N_13548,N_13974);
nand U14494 (N_14494,N_13754,N_13763);
and U14495 (N_14495,N_13923,N_13876);
nor U14496 (N_14496,N_13607,N_13944);
nor U14497 (N_14497,N_13846,N_13643);
or U14498 (N_14498,N_13776,N_13545);
and U14499 (N_14499,N_13575,N_13565);
and U14500 (N_14500,N_14003,N_14244);
and U14501 (N_14501,N_14065,N_14312);
xnor U14502 (N_14502,N_14473,N_14492);
nor U14503 (N_14503,N_14351,N_14225);
or U14504 (N_14504,N_14336,N_14403);
xnor U14505 (N_14505,N_14391,N_14438);
nand U14506 (N_14506,N_14376,N_14317);
and U14507 (N_14507,N_14134,N_14111);
xor U14508 (N_14508,N_14125,N_14216);
and U14509 (N_14509,N_14304,N_14018);
and U14510 (N_14510,N_14254,N_14084);
nand U14511 (N_14511,N_14187,N_14458);
and U14512 (N_14512,N_14296,N_14270);
nand U14513 (N_14513,N_14017,N_14379);
xnor U14514 (N_14514,N_14150,N_14268);
nor U14515 (N_14515,N_14013,N_14373);
nand U14516 (N_14516,N_14449,N_14195);
and U14517 (N_14517,N_14290,N_14162);
xnor U14518 (N_14518,N_14127,N_14407);
nand U14519 (N_14519,N_14217,N_14006);
xor U14520 (N_14520,N_14077,N_14352);
nand U14521 (N_14521,N_14339,N_14277);
nand U14522 (N_14522,N_14165,N_14474);
or U14523 (N_14523,N_14260,N_14020);
and U14524 (N_14524,N_14418,N_14069);
xnor U14525 (N_14525,N_14034,N_14201);
or U14526 (N_14526,N_14309,N_14206);
nand U14527 (N_14527,N_14093,N_14308);
nand U14528 (N_14528,N_14148,N_14412);
nor U14529 (N_14529,N_14116,N_14202);
nand U14530 (N_14530,N_14404,N_14072);
nand U14531 (N_14531,N_14200,N_14487);
or U14532 (N_14532,N_14490,N_14441);
nor U14533 (N_14533,N_14175,N_14040);
xor U14534 (N_14534,N_14298,N_14156);
xnor U14535 (N_14535,N_14051,N_14060);
xor U14536 (N_14536,N_14046,N_14106);
or U14537 (N_14537,N_14497,N_14024);
or U14538 (N_14538,N_14446,N_14213);
and U14539 (N_14539,N_14029,N_14274);
nor U14540 (N_14540,N_14480,N_14154);
nor U14541 (N_14541,N_14266,N_14416);
xnor U14542 (N_14542,N_14253,N_14372);
and U14543 (N_14543,N_14388,N_14121);
nand U14544 (N_14544,N_14435,N_14494);
nand U14545 (N_14545,N_14363,N_14076);
and U14546 (N_14546,N_14251,N_14048);
nand U14547 (N_14547,N_14395,N_14075);
or U14548 (N_14548,N_14205,N_14189);
xnor U14549 (N_14549,N_14219,N_14166);
xor U14550 (N_14550,N_14052,N_14002);
or U14551 (N_14551,N_14207,N_14393);
nand U14552 (N_14552,N_14285,N_14456);
and U14553 (N_14553,N_14311,N_14160);
xor U14554 (N_14554,N_14471,N_14481);
xnor U14555 (N_14555,N_14214,N_14239);
or U14556 (N_14556,N_14280,N_14193);
xnor U14557 (N_14557,N_14316,N_14287);
and U14558 (N_14558,N_14227,N_14089);
or U14559 (N_14559,N_14382,N_14218);
and U14560 (N_14560,N_14347,N_14233);
and U14561 (N_14561,N_14425,N_14235);
and U14562 (N_14562,N_14370,N_14348);
nand U14563 (N_14563,N_14318,N_14356);
and U14564 (N_14564,N_14001,N_14104);
and U14565 (N_14565,N_14050,N_14232);
xor U14566 (N_14566,N_14229,N_14273);
or U14567 (N_14567,N_14240,N_14056);
or U14568 (N_14568,N_14054,N_14291);
nor U14569 (N_14569,N_14431,N_14059);
and U14570 (N_14570,N_14461,N_14468);
xnor U14571 (N_14571,N_14228,N_14132);
and U14572 (N_14572,N_14293,N_14279);
or U14573 (N_14573,N_14381,N_14362);
nand U14574 (N_14574,N_14129,N_14495);
or U14575 (N_14575,N_14000,N_14126);
nand U14576 (N_14576,N_14032,N_14338);
and U14577 (N_14577,N_14271,N_14476);
nor U14578 (N_14578,N_14385,N_14445);
nor U14579 (N_14579,N_14344,N_14022);
nor U14580 (N_14580,N_14158,N_14103);
xor U14581 (N_14581,N_14028,N_14463);
nor U14582 (N_14582,N_14163,N_14210);
or U14583 (N_14583,N_14153,N_14394);
xnor U14584 (N_14584,N_14136,N_14088);
nor U14585 (N_14585,N_14357,N_14030);
xor U14586 (N_14586,N_14236,N_14183);
xor U14587 (N_14587,N_14447,N_14284);
xnor U14588 (N_14588,N_14428,N_14408);
or U14589 (N_14589,N_14499,N_14102);
nor U14590 (N_14590,N_14475,N_14374);
and U14591 (N_14591,N_14122,N_14410);
or U14592 (N_14592,N_14215,N_14267);
and U14593 (N_14593,N_14007,N_14044);
and U14594 (N_14594,N_14263,N_14423);
nand U14595 (N_14595,N_14063,N_14467);
nor U14596 (N_14596,N_14455,N_14442);
and U14597 (N_14597,N_14097,N_14451);
nand U14598 (N_14598,N_14469,N_14249);
nand U14599 (N_14599,N_14432,N_14272);
xor U14600 (N_14600,N_14264,N_14314);
and U14601 (N_14601,N_14367,N_14434);
and U14602 (N_14602,N_14143,N_14101);
xnor U14603 (N_14603,N_14483,N_14406);
or U14604 (N_14604,N_14098,N_14437);
and U14605 (N_14605,N_14064,N_14041);
xor U14606 (N_14606,N_14329,N_14286);
or U14607 (N_14607,N_14074,N_14057);
and U14608 (N_14608,N_14230,N_14283);
nor U14609 (N_14609,N_14333,N_14105);
xor U14610 (N_14610,N_14259,N_14169);
nand U14611 (N_14611,N_14489,N_14026);
and U14612 (N_14612,N_14459,N_14188);
and U14613 (N_14613,N_14349,N_14145);
and U14614 (N_14614,N_14310,N_14377);
nor U14615 (N_14615,N_14096,N_14365);
xnor U14616 (N_14616,N_14371,N_14464);
nor U14617 (N_14617,N_14176,N_14067);
xor U14618 (N_14618,N_14012,N_14439);
or U14619 (N_14619,N_14453,N_14042);
nor U14620 (N_14620,N_14095,N_14341);
nor U14621 (N_14621,N_14212,N_14025);
nor U14622 (N_14622,N_14430,N_14482);
xor U14623 (N_14623,N_14269,N_14429);
nor U14624 (N_14624,N_14004,N_14350);
or U14625 (N_14625,N_14109,N_14378);
nand U14626 (N_14626,N_14295,N_14062);
nor U14627 (N_14627,N_14128,N_14325);
or U14628 (N_14628,N_14384,N_14328);
xnor U14629 (N_14629,N_14208,N_14427);
nand U14630 (N_14630,N_14462,N_14281);
or U14631 (N_14631,N_14409,N_14184);
nand U14632 (N_14632,N_14226,N_14448);
and U14633 (N_14633,N_14426,N_14091);
nand U14634 (N_14634,N_14199,N_14323);
nor U14635 (N_14635,N_14288,N_14300);
and U14636 (N_14636,N_14340,N_14079);
or U14637 (N_14637,N_14436,N_14250);
nand U14638 (N_14638,N_14223,N_14337);
nor U14639 (N_14639,N_14090,N_14016);
xnor U14640 (N_14640,N_14036,N_14100);
xor U14641 (N_14641,N_14297,N_14139);
xnor U14642 (N_14642,N_14112,N_14238);
nor U14643 (N_14643,N_14421,N_14142);
nor U14644 (N_14644,N_14420,N_14019);
or U14645 (N_14645,N_14248,N_14211);
nor U14646 (N_14646,N_14444,N_14010);
nor U14647 (N_14647,N_14324,N_14167);
or U14648 (N_14648,N_14173,N_14196);
and U14649 (N_14649,N_14043,N_14402);
xor U14650 (N_14650,N_14389,N_14400);
nor U14651 (N_14651,N_14155,N_14190);
nand U14652 (N_14652,N_14078,N_14392);
or U14653 (N_14653,N_14247,N_14083);
xor U14654 (N_14654,N_14342,N_14164);
xnor U14655 (N_14655,N_14405,N_14144);
xor U14656 (N_14656,N_14023,N_14231);
nor U14657 (N_14657,N_14086,N_14422);
nor U14658 (N_14658,N_14107,N_14478);
xor U14659 (N_14659,N_14237,N_14417);
or U14660 (N_14660,N_14015,N_14009);
and U14661 (N_14661,N_14488,N_14031);
xnor U14662 (N_14662,N_14361,N_14307);
nand U14663 (N_14663,N_14454,N_14061);
and U14664 (N_14664,N_14011,N_14343);
nand U14665 (N_14665,N_14198,N_14419);
nor U14666 (N_14666,N_14301,N_14209);
nand U14667 (N_14667,N_14053,N_14068);
nor U14668 (N_14668,N_14413,N_14368);
xnor U14669 (N_14669,N_14038,N_14243);
and U14670 (N_14670,N_14037,N_14326);
xnor U14671 (N_14671,N_14354,N_14114);
nor U14672 (N_14672,N_14319,N_14452);
nor U14673 (N_14673,N_14353,N_14070);
nand U14674 (N_14674,N_14222,N_14130);
or U14675 (N_14675,N_14278,N_14181);
or U14676 (N_14676,N_14147,N_14180);
nor U14677 (N_14677,N_14241,N_14203);
nor U14678 (N_14678,N_14360,N_14364);
nand U14679 (N_14679,N_14275,N_14246);
nor U14680 (N_14680,N_14398,N_14411);
xnor U14681 (N_14681,N_14027,N_14123);
nor U14682 (N_14682,N_14282,N_14261);
xor U14683 (N_14683,N_14194,N_14486);
nand U14684 (N_14684,N_14386,N_14185);
nor U14685 (N_14685,N_14322,N_14334);
nand U14686 (N_14686,N_14152,N_14470);
xnor U14687 (N_14687,N_14039,N_14257);
and U14688 (N_14688,N_14465,N_14157);
or U14689 (N_14689,N_14138,N_14440);
xor U14690 (N_14690,N_14120,N_14131);
nor U14691 (N_14691,N_14085,N_14224);
or U14692 (N_14692,N_14177,N_14457);
xor U14693 (N_14693,N_14258,N_14073);
nor U14694 (N_14694,N_14390,N_14256);
or U14695 (N_14695,N_14479,N_14294);
and U14696 (N_14696,N_14276,N_14460);
nor U14697 (N_14697,N_14359,N_14033);
or U14698 (N_14698,N_14047,N_14383);
or U14699 (N_14699,N_14305,N_14265);
xor U14700 (N_14700,N_14055,N_14110);
xnor U14701 (N_14701,N_14182,N_14066);
and U14702 (N_14702,N_14433,N_14321);
and U14703 (N_14703,N_14380,N_14220);
or U14704 (N_14704,N_14133,N_14178);
nor U14705 (N_14705,N_14358,N_14375);
nor U14706 (N_14706,N_14204,N_14192);
and U14707 (N_14707,N_14124,N_14113);
nor U14708 (N_14708,N_14443,N_14117);
nand U14709 (N_14709,N_14399,N_14108);
nor U14710 (N_14710,N_14498,N_14346);
xor U14711 (N_14711,N_14302,N_14306);
xor U14712 (N_14712,N_14387,N_14242);
nand U14713 (N_14713,N_14366,N_14327);
and U14714 (N_14714,N_14466,N_14135);
xor U14715 (N_14715,N_14335,N_14099);
nor U14716 (N_14716,N_14330,N_14484);
nor U14717 (N_14717,N_14146,N_14081);
nand U14718 (N_14718,N_14008,N_14485);
nand U14719 (N_14719,N_14289,N_14424);
nor U14720 (N_14720,N_14186,N_14191);
or U14721 (N_14721,N_14174,N_14472);
xnor U14722 (N_14722,N_14396,N_14049);
nor U14723 (N_14723,N_14369,N_14299);
nand U14724 (N_14724,N_14245,N_14234);
nor U14725 (N_14725,N_14332,N_14303);
and U14726 (N_14726,N_14171,N_14179);
nor U14727 (N_14727,N_14161,N_14094);
or U14728 (N_14728,N_14414,N_14221);
or U14729 (N_14729,N_14045,N_14058);
and U14730 (N_14730,N_14493,N_14315);
nor U14731 (N_14731,N_14172,N_14491);
nand U14732 (N_14732,N_14118,N_14035);
nand U14733 (N_14733,N_14080,N_14496);
nand U14734 (N_14734,N_14255,N_14159);
and U14735 (N_14735,N_14415,N_14005);
nand U14736 (N_14736,N_14071,N_14151);
xnor U14737 (N_14737,N_14014,N_14320);
or U14738 (N_14738,N_14137,N_14450);
nor U14739 (N_14739,N_14331,N_14401);
or U14740 (N_14740,N_14141,N_14292);
and U14741 (N_14741,N_14087,N_14252);
nand U14742 (N_14742,N_14345,N_14170);
xnor U14743 (N_14743,N_14313,N_14082);
nor U14744 (N_14744,N_14197,N_14149);
and U14745 (N_14745,N_14140,N_14355);
xnor U14746 (N_14746,N_14119,N_14262);
xnor U14747 (N_14747,N_14092,N_14477);
xor U14748 (N_14748,N_14397,N_14168);
xnor U14749 (N_14749,N_14021,N_14115);
and U14750 (N_14750,N_14442,N_14397);
or U14751 (N_14751,N_14041,N_14034);
and U14752 (N_14752,N_14007,N_14246);
nor U14753 (N_14753,N_14379,N_14152);
nand U14754 (N_14754,N_14111,N_14124);
nand U14755 (N_14755,N_14197,N_14431);
xor U14756 (N_14756,N_14304,N_14033);
nor U14757 (N_14757,N_14435,N_14398);
and U14758 (N_14758,N_14176,N_14189);
xor U14759 (N_14759,N_14483,N_14318);
or U14760 (N_14760,N_14427,N_14285);
or U14761 (N_14761,N_14059,N_14271);
xor U14762 (N_14762,N_14293,N_14234);
nand U14763 (N_14763,N_14082,N_14183);
and U14764 (N_14764,N_14310,N_14442);
nand U14765 (N_14765,N_14212,N_14391);
xor U14766 (N_14766,N_14481,N_14056);
xnor U14767 (N_14767,N_14346,N_14299);
nand U14768 (N_14768,N_14035,N_14164);
and U14769 (N_14769,N_14117,N_14063);
nand U14770 (N_14770,N_14143,N_14260);
and U14771 (N_14771,N_14112,N_14403);
or U14772 (N_14772,N_14394,N_14194);
nand U14773 (N_14773,N_14107,N_14143);
nor U14774 (N_14774,N_14400,N_14139);
or U14775 (N_14775,N_14055,N_14300);
nand U14776 (N_14776,N_14091,N_14314);
xor U14777 (N_14777,N_14108,N_14345);
and U14778 (N_14778,N_14119,N_14412);
nand U14779 (N_14779,N_14343,N_14055);
and U14780 (N_14780,N_14195,N_14212);
nor U14781 (N_14781,N_14133,N_14281);
and U14782 (N_14782,N_14289,N_14279);
xor U14783 (N_14783,N_14254,N_14055);
xnor U14784 (N_14784,N_14050,N_14230);
and U14785 (N_14785,N_14085,N_14074);
and U14786 (N_14786,N_14358,N_14177);
or U14787 (N_14787,N_14111,N_14177);
and U14788 (N_14788,N_14427,N_14296);
nor U14789 (N_14789,N_14235,N_14056);
nor U14790 (N_14790,N_14080,N_14368);
nand U14791 (N_14791,N_14061,N_14134);
nor U14792 (N_14792,N_14219,N_14107);
nand U14793 (N_14793,N_14109,N_14293);
and U14794 (N_14794,N_14440,N_14192);
xnor U14795 (N_14795,N_14300,N_14301);
or U14796 (N_14796,N_14020,N_14472);
xor U14797 (N_14797,N_14037,N_14491);
nand U14798 (N_14798,N_14412,N_14169);
nor U14799 (N_14799,N_14451,N_14033);
or U14800 (N_14800,N_14354,N_14223);
and U14801 (N_14801,N_14383,N_14104);
or U14802 (N_14802,N_14210,N_14371);
nand U14803 (N_14803,N_14335,N_14488);
nor U14804 (N_14804,N_14139,N_14325);
and U14805 (N_14805,N_14136,N_14399);
nor U14806 (N_14806,N_14161,N_14482);
and U14807 (N_14807,N_14306,N_14147);
xnor U14808 (N_14808,N_14344,N_14295);
or U14809 (N_14809,N_14145,N_14130);
nand U14810 (N_14810,N_14124,N_14350);
and U14811 (N_14811,N_14226,N_14350);
or U14812 (N_14812,N_14041,N_14156);
nor U14813 (N_14813,N_14073,N_14402);
and U14814 (N_14814,N_14387,N_14187);
nand U14815 (N_14815,N_14077,N_14267);
xor U14816 (N_14816,N_14118,N_14227);
xor U14817 (N_14817,N_14396,N_14175);
and U14818 (N_14818,N_14112,N_14225);
or U14819 (N_14819,N_14451,N_14288);
nand U14820 (N_14820,N_14290,N_14204);
xnor U14821 (N_14821,N_14226,N_14487);
or U14822 (N_14822,N_14228,N_14496);
nor U14823 (N_14823,N_14484,N_14307);
and U14824 (N_14824,N_14410,N_14013);
nor U14825 (N_14825,N_14165,N_14463);
nand U14826 (N_14826,N_14372,N_14077);
and U14827 (N_14827,N_14303,N_14334);
or U14828 (N_14828,N_14284,N_14352);
and U14829 (N_14829,N_14039,N_14259);
and U14830 (N_14830,N_14052,N_14443);
xor U14831 (N_14831,N_14394,N_14416);
xor U14832 (N_14832,N_14428,N_14060);
and U14833 (N_14833,N_14133,N_14260);
or U14834 (N_14834,N_14397,N_14491);
xnor U14835 (N_14835,N_14215,N_14349);
or U14836 (N_14836,N_14132,N_14350);
or U14837 (N_14837,N_14055,N_14212);
nand U14838 (N_14838,N_14258,N_14147);
xnor U14839 (N_14839,N_14254,N_14147);
xor U14840 (N_14840,N_14090,N_14027);
and U14841 (N_14841,N_14221,N_14030);
xnor U14842 (N_14842,N_14498,N_14076);
xnor U14843 (N_14843,N_14217,N_14139);
nor U14844 (N_14844,N_14227,N_14228);
nor U14845 (N_14845,N_14434,N_14303);
nor U14846 (N_14846,N_14488,N_14002);
nand U14847 (N_14847,N_14187,N_14012);
nor U14848 (N_14848,N_14024,N_14459);
and U14849 (N_14849,N_14207,N_14037);
and U14850 (N_14850,N_14430,N_14398);
nand U14851 (N_14851,N_14177,N_14336);
nand U14852 (N_14852,N_14094,N_14287);
or U14853 (N_14853,N_14463,N_14313);
xor U14854 (N_14854,N_14004,N_14295);
and U14855 (N_14855,N_14154,N_14229);
nor U14856 (N_14856,N_14471,N_14491);
nor U14857 (N_14857,N_14107,N_14081);
nand U14858 (N_14858,N_14244,N_14088);
or U14859 (N_14859,N_14452,N_14392);
and U14860 (N_14860,N_14095,N_14266);
or U14861 (N_14861,N_14315,N_14287);
xor U14862 (N_14862,N_14019,N_14255);
nor U14863 (N_14863,N_14363,N_14379);
nand U14864 (N_14864,N_14295,N_14177);
or U14865 (N_14865,N_14147,N_14433);
nand U14866 (N_14866,N_14397,N_14000);
and U14867 (N_14867,N_14367,N_14306);
and U14868 (N_14868,N_14158,N_14409);
or U14869 (N_14869,N_14042,N_14090);
nor U14870 (N_14870,N_14346,N_14331);
or U14871 (N_14871,N_14499,N_14357);
nor U14872 (N_14872,N_14470,N_14033);
and U14873 (N_14873,N_14472,N_14008);
nor U14874 (N_14874,N_14258,N_14088);
and U14875 (N_14875,N_14422,N_14226);
nor U14876 (N_14876,N_14371,N_14290);
xor U14877 (N_14877,N_14184,N_14442);
or U14878 (N_14878,N_14409,N_14440);
xor U14879 (N_14879,N_14089,N_14259);
xnor U14880 (N_14880,N_14350,N_14030);
xnor U14881 (N_14881,N_14187,N_14331);
xnor U14882 (N_14882,N_14093,N_14008);
and U14883 (N_14883,N_14268,N_14482);
or U14884 (N_14884,N_14075,N_14490);
and U14885 (N_14885,N_14193,N_14366);
and U14886 (N_14886,N_14362,N_14451);
and U14887 (N_14887,N_14107,N_14188);
xor U14888 (N_14888,N_14085,N_14461);
nor U14889 (N_14889,N_14302,N_14460);
xor U14890 (N_14890,N_14281,N_14220);
nand U14891 (N_14891,N_14162,N_14176);
nor U14892 (N_14892,N_14424,N_14188);
nand U14893 (N_14893,N_14286,N_14157);
nand U14894 (N_14894,N_14148,N_14158);
nor U14895 (N_14895,N_14194,N_14447);
nand U14896 (N_14896,N_14278,N_14330);
and U14897 (N_14897,N_14442,N_14069);
xnor U14898 (N_14898,N_14007,N_14455);
nand U14899 (N_14899,N_14334,N_14247);
nor U14900 (N_14900,N_14180,N_14372);
or U14901 (N_14901,N_14416,N_14048);
or U14902 (N_14902,N_14462,N_14378);
or U14903 (N_14903,N_14354,N_14000);
xor U14904 (N_14904,N_14143,N_14052);
xor U14905 (N_14905,N_14423,N_14123);
or U14906 (N_14906,N_14028,N_14083);
and U14907 (N_14907,N_14432,N_14391);
or U14908 (N_14908,N_14496,N_14480);
and U14909 (N_14909,N_14415,N_14090);
nand U14910 (N_14910,N_14122,N_14236);
xnor U14911 (N_14911,N_14228,N_14239);
or U14912 (N_14912,N_14411,N_14090);
nand U14913 (N_14913,N_14108,N_14298);
xor U14914 (N_14914,N_14319,N_14231);
xor U14915 (N_14915,N_14324,N_14160);
xor U14916 (N_14916,N_14492,N_14163);
nand U14917 (N_14917,N_14010,N_14266);
xnor U14918 (N_14918,N_14172,N_14269);
and U14919 (N_14919,N_14038,N_14170);
xnor U14920 (N_14920,N_14156,N_14169);
and U14921 (N_14921,N_14037,N_14453);
nand U14922 (N_14922,N_14484,N_14281);
or U14923 (N_14923,N_14073,N_14439);
xor U14924 (N_14924,N_14127,N_14257);
and U14925 (N_14925,N_14155,N_14421);
xor U14926 (N_14926,N_14039,N_14262);
and U14927 (N_14927,N_14379,N_14099);
xnor U14928 (N_14928,N_14418,N_14131);
and U14929 (N_14929,N_14406,N_14312);
or U14930 (N_14930,N_14388,N_14184);
nor U14931 (N_14931,N_14002,N_14303);
nand U14932 (N_14932,N_14116,N_14101);
xnor U14933 (N_14933,N_14414,N_14399);
nor U14934 (N_14934,N_14440,N_14268);
nor U14935 (N_14935,N_14368,N_14423);
nand U14936 (N_14936,N_14371,N_14194);
and U14937 (N_14937,N_14068,N_14148);
nand U14938 (N_14938,N_14207,N_14284);
and U14939 (N_14939,N_14253,N_14172);
nor U14940 (N_14940,N_14024,N_14114);
nand U14941 (N_14941,N_14441,N_14321);
or U14942 (N_14942,N_14427,N_14040);
xnor U14943 (N_14943,N_14342,N_14142);
or U14944 (N_14944,N_14378,N_14082);
or U14945 (N_14945,N_14171,N_14365);
nand U14946 (N_14946,N_14274,N_14385);
xor U14947 (N_14947,N_14388,N_14142);
xnor U14948 (N_14948,N_14274,N_14261);
nand U14949 (N_14949,N_14130,N_14327);
xor U14950 (N_14950,N_14246,N_14005);
xnor U14951 (N_14951,N_14342,N_14096);
nor U14952 (N_14952,N_14291,N_14124);
and U14953 (N_14953,N_14233,N_14464);
and U14954 (N_14954,N_14157,N_14178);
or U14955 (N_14955,N_14223,N_14042);
xnor U14956 (N_14956,N_14350,N_14286);
nor U14957 (N_14957,N_14312,N_14170);
nand U14958 (N_14958,N_14194,N_14024);
and U14959 (N_14959,N_14298,N_14222);
or U14960 (N_14960,N_14488,N_14197);
nand U14961 (N_14961,N_14212,N_14127);
xnor U14962 (N_14962,N_14128,N_14361);
nand U14963 (N_14963,N_14147,N_14279);
xnor U14964 (N_14964,N_14464,N_14447);
and U14965 (N_14965,N_14050,N_14123);
nor U14966 (N_14966,N_14492,N_14159);
or U14967 (N_14967,N_14347,N_14292);
and U14968 (N_14968,N_14174,N_14091);
and U14969 (N_14969,N_14106,N_14081);
nor U14970 (N_14970,N_14207,N_14367);
xor U14971 (N_14971,N_14130,N_14268);
or U14972 (N_14972,N_14390,N_14337);
nand U14973 (N_14973,N_14481,N_14090);
nor U14974 (N_14974,N_14033,N_14496);
xnor U14975 (N_14975,N_14395,N_14356);
nand U14976 (N_14976,N_14483,N_14487);
or U14977 (N_14977,N_14224,N_14089);
nor U14978 (N_14978,N_14285,N_14024);
or U14979 (N_14979,N_14381,N_14022);
nand U14980 (N_14980,N_14469,N_14193);
or U14981 (N_14981,N_14249,N_14116);
nor U14982 (N_14982,N_14495,N_14225);
nand U14983 (N_14983,N_14062,N_14229);
nor U14984 (N_14984,N_14272,N_14019);
nand U14985 (N_14985,N_14399,N_14455);
xor U14986 (N_14986,N_14107,N_14137);
or U14987 (N_14987,N_14167,N_14360);
or U14988 (N_14988,N_14280,N_14166);
xnor U14989 (N_14989,N_14380,N_14207);
nand U14990 (N_14990,N_14054,N_14485);
xnor U14991 (N_14991,N_14487,N_14373);
or U14992 (N_14992,N_14352,N_14450);
or U14993 (N_14993,N_14454,N_14286);
xnor U14994 (N_14994,N_14445,N_14425);
xnor U14995 (N_14995,N_14271,N_14371);
nand U14996 (N_14996,N_14007,N_14040);
and U14997 (N_14997,N_14208,N_14150);
nor U14998 (N_14998,N_14110,N_14413);
xnor U14999 (N_14999,N_14024,N_14161);
nor U15000 (N_15000,N_14578,N_14977);
or U15001 (N_15001,N_14633,N_14534);
nor U15002 (N_15002,N_14900,N_14599);
xor U15003 (N_15003,N_14697,N_14753);
xnor U15004 (N_15004,N_14515,N_14645);
xor U15005 (N_15005,N_14615,N_14685);
nor U15006 (N_15006,N_14519,N_14993);
nand U15007 (N_15007,N_14626,N_14548);
and U15008 (N_15008,N_14516,N_14701);
nor U15009 (N_15009,N_14554,N_14544);
nor U15010 (N_15010,N_14862,N_14780);
or U15011 (N_15011,N_14666,N_14819);
nor U15012 (N_15012,N_14600,N_14558);
or U15013 (N_15013,N_14957,N_14939);
xnor U15014 (N_15014,N_14811,N_14816);
nor U15015 (N_15015,N_14768,N_14836);
nand U15016 (N_15016,N_14739,N_14875);
xnor U15017 (N_15017,N_14892,N_14763);
nand U15018 (N_15018,N_14832,N_14770);
or U15019 (N_15019,N_14620,N_14513);
nor U15020 (N_15020,N_14525,N_14536);
xnor U15021 (N_15021,N_14824,N_14781);
and U15022 (N_15022,N_14786,N_14532);
or U15023 (N_15023,N_14775,N_14910);
nor U15024 (N_15024,N_14585,N_14922);
and U15025 (N_15025,N_14876,N_14679);
or U15026 (N_15026,N_14983,N_14877);
nor U15027 (N_15027,N_14627,N_14510);
or U15028 (N_15028,N_14864,N_14800);
and U15029 (N_15029,N_14718,N_14648);
xnor U15030 (N_15030,N_14603,N_14708);
and U15031 (N_15031,N_14611,N_14721);
xor U15032 (N_15032,N_14590,N_14569);
xor U15033 (N_15033,N_14764,N_14767);
nand U15034 (N_15034,N_14621,N_14695);
and U15035 (N_15035,N_14833,N_14867);
xnor U15036 (N_15036,N_14671,N_14973);
and U15037 (N_15037,N_14509,N_14658);
or U15038 (N_15038,N_14559,N_14779);
or U15039 (N_15039,N_14907,N_14637);
nor U15040 (N_15040,N_14562,N_14817);
xnor U15041 (N_15041,N_14681,N_14706);
or U15042 (N_15042,N_14860,N_14809);
nor U15043 (N_15043,N_14804,N_14783);
nand U15044 (N_15044,N_14822,N_14528);
xnor U15045 (N_15045,N_14931,N_14712);
nand U15046 (N_15046,N_14690,N_14674);
nor U15047 (N_15047,N_14890,N_14608);
xnor U15048 (N_15048,N_14547,N_14882);
nand U15049 (N_15049,N_14921,N_14537);
nor U15050 (N_15050,N_14888,N_14623);
and U15051 (N_15051,N_14802,N_14517);
nor U15052 (N_15052,N_14868,N_14514);
and U15053 (N_15053,N_14855,N_14959);
and U15054 (N_15054,N_14814,N_14684);
or U15055 (N_15055,N_14696,N_14619);
nand U15056 (N_15056,N_14917,N_14967);
and U15057 (N_15057,N_14579,N_14932);
nor U15058 (N_15058,N_14575,N_14591);
xor U15059 (N_15059,N_14720,N_14915);
xnor U15060 (N_15060,N_14657,N_14806);
xor U15061 (N_15061,N_14842,N_14796);
or U15062 (N_15062,N_14880,N_14972);
or U15063 (N_15063,N_14595,N_14500);
nand U15064 (N_15064,N_14971,N_14571);
nand U15065 (N_15065,N_14730,N_14556);
nand U15066 (N_15066,N_14873,N_14778);
and U15067 (N_15067,N_14638,N_14747);
nor U15068 (N_15068,N_14676,N_14568);
and U15069 (N_15069,N_14636,N_14731);
xnor U15070 (N_15070,N_14863,N_14606);
and U15071 (N_15071,N_14826,N_14925);
or U15072 (N_15072,N_14656,N_14605);
or U15073 (N_15073,N_14555,N_14808);
and U15074 (N_15074,N_14574,N_14709);
nor U15075 (N_15075,N_14609,N_14991);
xor U15076 (N_15076,N_14791,N_14962);
nand U15077 (N_15077,N_14717,N_14834);
nor U15078 (N_15078,N_14713,N_14845);
and U15079 (N_15079,N_14934,N_14508);
nor U15080 (N_15080,N_14869,N_14761);
nand U15081 (N_15081,N_14948,N_14872);
or U15082 (N_15082,N_14687,N_14805);
or U15083 (N_15083,N_14997,N_14985);
or U15084 (N_15084,N_14693,N_14654);
nor U15085 (N_15085,N_14735,N_14533);
or U15086 (N_15086,N_14522,N_14592);
and U15087 (N_15087,N_14604,N_14602);
and U15088 (N_15088,N_14851,N_14956);
or U15089 (N_15089,N_14572,N_14797);
xor U15090 (N_15090,N_14526,N_14632);
nand U15091 (N_15091,N_14530,N_14771);
nand U15092 (N_15092,N_14901,N_14577);
nor U15093 (N_15093,N_14897,N_14736);
or U15094 (N_15094,N_14879,N_14886);
and U15095 (N_15095,N_14788,N_14689);
and U15096 (N_15096,N_14981,N_14634);
nor U15097 (N_15097,N_14945,N_14918);
nand U15098 (N_15098,N_14738,N_14541);
xor U15099 (N_15099,N_14758,N_14589);
nor U15100 (N_15100,N_14774,N_14828);
nor U15101 (N_15101,N_14520,N_14955);
nor U15102 (N_15102,N_14740,N_14870);
nand U15103 (N_15103,N_14707,N_14573);
nand U15104 (N_15104,N_14649,N_14881);
and U15105 (N_15105,N_14843,N_14839);
and U15106 (N_15106,N_14607,N_14680);
nor U15107 (N_15107,N_14874,N_14821);
and U15108 (N_15108,N_14640,N_14546);
nor U15109 (N_15109,N_14848,N_14567);
or U15110 (N_15110,N_14803,N_14561);
xor U15111 (N_15111,N_14798,N_14705);
or U15112 (N_15112,N_14960,N_14831);
nand U15113 (N_15113,N_14675,N_14686);
nor U15114 (N_15114,N_14952,N_14902);
xnor U15115 (N_15115,N_14540,N_14950);
nand U15116 (N_15116,N_14523,N_14856);
or U15117 (N_15117,N_14930,N_14988);
xnor U15118 (N_15118,N_14969,N_14916);
xnor U15119 (N_15119,N_14908,N_14820);
xor U15120 (N_15120,N_14751,N_14750);
xor U15121 (N_15121,N_14926,N_14813);
xor U15122 (N_15122,N_14777,N_14885);
or U15123 (N_15123,N_14964,N_14992);
xor U15124 (N_15124,N_14723,N_14576);
nor U15125 (N_15125,N_14852,N_14745);
xor U15126 (N_15126,N_14958,N_14672);
nand U15127 (N_15127,N_14664,N_14838);
and U15128 (N_15128,N_14871,N_14641);
xnor U15129 (N_15129,N_14527,N_14728);
or U15130 (N_15130,N_14963,N_14986);
xnor U15131 (N_15131,N_14629,N_14793);
and U15132 (N_15132,N_14665,N_14976);
and U15133 (N_15133,N_14951,N_14953);
or U15134 (N_15134,N_14759,N_14700);
nand U15135 (N_15135,N_14929,N_14812);
nor U15136 (N_15136,N_14789,N_14741);
and U15137 (N_15137,N_14889,N_14743);
and U15138 (N_15138,N_14563,N_14754);
and U15139 (N_15139,N_14724,N_14703);
and U15140 (N_15140,N_14524,N_14699);
xnor U15141 (N_15141,N_14954,N_14841);
nand U15142 (N_15142,N_14887,N_14883);
nand U15143 (N_15143,N_14913,N_14928);
xor U15144 (N_15144,N_14587,N_14504);
or U15145 (N_15145,N_14990,N_14722);
and U15146 (N_15146,N_14702,N_14978);
nor U15147 (N_15147,N_14998,N_14584);
nor U15148 (N_15148,N_14947,N_14949);
nand U15149 (N_15149,N_14503,N_14994);
xnor U15150 (N_15150,N_14807,N_14757);
nand U15151 (N_15151,N_14936,N_14944);
nand U15152 (N_15152,N_14614,N_14861);
xor U15153 (N_15153,N_14529,N_14923);
nor U15154 (N_15154,N_14628,N_14840);
nor U15155 (N_15155,N_14688,N_14975);
and U15156 (N_15156,N_14588,N_14801);
or U15157 (N_15157,N_14586,N_14622);
xnor U15158 (N_15158,N_14711,N_14610);
xor U15159 (N_15159,N_14570,N_14748);
and U15160 (N_15160,N_14765,N_14582);
and U15161 (N_15161,N_14909,N_14837);
nand U15162 (N_15162,N_14726,N_14799);
and U15163 (N_15163,N_14835,N_14815);
xnor U15164 (N_15164,N_14539,N_14650);
xor U15165 (N_15165,N_14933,N_14659);
nor U15166 (N_15166,N_14760,N_14678);
nand U15167 (N_15167,N_14668,N_14551);
xnor U15168 (N_15168,N_14982,N_14827);
nor U15169 (N_15169,N_14938,N_14661);
xnor U15170 (N_15170,N_14894,N_14940);
nor U15171 (N_15171,N_14772,N_14847);
or U15172 (N_15172,N_14552,N_14531);
nand U15173 (N_15173,N_14716,N_14501);
and U15174 (N_15174,N_14698,N_14566);
and U15175 (N_15175,N_14974,N_14598);
or U15176 (N_15176,N_14903,N_14677);
xnor U15177 (N_15177,N_14912,N_14564);
or U15178 (N_15178,N_14752,N_14630);
xor U15179 (N_15179,N_14670,N_14535);
and U15180 (N_15180,N_14792,N_14543);
or U15181 (N_15181,N_14639,N_14596);
and U15182 (N_15182,N_14631,N_14970);
xor U15183 (N_15183,N_14651,N_14612);
and U15184 (N_15184,N_14553,N_14943);
nor U15185 (N_15185,N_14823,N_14647);
or U15186 (N_15186,N_14557,N_14727);
and U15187 (N_15187,N_14904,N_14506);
nand U15188 (N_15188,N_14518,N_14733);
xnor U15189 (N_15189,N_14979,N_14507);
nand U15190 (N_15190,N_14866,N_14853);
nor U15191 (N_15191,N_14941,N_14884);
nand U15192 (N_15192,N_14737,N_14719);
and U15193 (N_15193,N_14818,N_14729);
xnor U15194 (N_15194,N_14660,N_14893);
or U15195 (N_15195,N_14787,N_14987);
nor U15196 (N_15196,N_14635,N_14858);
and U15197 (N_15197,N_14725,N_14996);
nand U15198 (N_15198,N_14502,N_14891);
nor U15199 (N_15199,N_14906,N_14618);
nand U15200 (N_15200,N_14927,N_14776);
nand U15201 (N_15201,N_14646,N_14825);
nand U15202 (N_15202,N_14542,N_14625);
or U15203 (N_15203,N_14505,N_14854);
nand U15204 (N_15204,N_14597,N_14538);
xor U15205 (N_15205,N_14896,N_14755);
and U15206 (N_15206,N_14683,N_14617);
and U15207 (N_15207,N_14662,N_14624);
nor U15208 (N_15208,N_14643,N_14756);
nor U15209 (N_15209,N_14859,N_14914);
and U15210 (N_15210,N_14715,N_14810);
nand U15211 (N_15211,N_14692,N_14694);
nand U15212 (N_15212,N_14911,N_14593);
xor U15213 (N_15213,N_14762,N_14710);
or U15214 (N_15214,N_14663,N_14521);
nand U15215 (N_15215,N_14935,N_14790);
and U15216 (N_15216,N_14580,N_14895);
or U15217 (N_15217,N_14682,N_14924);
nor U15218 (N_15218,N_14920,N_14549);
or U15219 (N_15219,N_14795,N_14644);
or U15220 (N_15220,N_14937,N_14966);
and U15221 (N_15221,N_14989,N_14995);
nand U15222 (N_15222,N_14849,N_14714);
and U15223 (N_15223,N_14905,N_14999);
or U15224 (N_15224,N_14642,N_14667);
or U15225 (N_15225,N_14560,N_14601);
nand U15226 (N_15226,N_14946,N_14773);
nand U15227 (N_15227,N_14766,N_14653);
xnor U15228 (N_15228,N_14769,N_14581);
nand U15229 (N_15229,N_14850,N_14594);
nand U15230 (N_15230,N_14898,N_14732);
xnor U15231 (N_15231,N_14865,N_14512);
and U15232 (N_15232,N_14511,N_14857);
xor U15233 (N_15233,N_14919,N_14744);
nand U15234 (N_15234,N_14942,N_14734);
or U15235 (N_15235,N_14829,N_14673);
nand U15236 (N_15236,N_14583,N_14749);
nor U15237 (N_15237,N_14613,N_14704);
nand U15238 (N_15238,N_14784,N_14961);
xor U15239 (N_15239,N_14655,N_14899);
nand U15240 (N_15240,N_14830,N_14785);
nand U15241 (N_15241,N_14984,N_14878);
nand U15242 (N_15242,N_14782,N_14965);
nand U15243 (N_15243,N_14652,N_14616);
or U15244 (N_15244,N_14746,N_14846);
nor U15245 (N_15245,N_14691,N_14545);
and U15246 (N_15246,N_14794,N_14980);
and U15247 (N_15247,N_14669,N_14968);
nand U15248 (N_15248,N_14565,N_14742);
nand U15249 (N_15249,N_14844,N_14550);
nand U15250 (N_15250,N_14794,N_14923);
or U15251 (N_15251,N_14616,N_14919);
nand U15252 (N_15252,N_14629,N_14761);
xnor U15253 (N_15253,N_14596,N_14795);
nand U15254 (N_15254,N_14901,N_14705);
nand U15255 (N_15255,N_14685,N_14821);
nand U15256 (N_15256,N_14684,N_14900);
or U15257 (N_15257,N_14624,N_14588);
nor U15258 (N_15258,N_14968,N_14853);
nand U15259 (N_15259,N_14954,N_14943);
xnor U15260 (N_15260,N_14618,N_14950);
xnor U15261 (N_15261,N_14895,N_14723);
xnor U15262 (N_15262,N_14659,N_14609);
nor U15263 (N_15263,N_14967,N_14801);
nand U15264 (N_15264,N_14531,N_14605);
xnor U15265 (N_15265,N_14874,N_14871);
nor U15266 (N_15266,N_14739,N_14550);
xnor U15267 (N_15267,N_14870,N_14948);
nor U15268 (N_15268,N_14737,N_14606);
or U15269 (N_15269,N_14788,N_14929);
or U15270 (N_15270,N_14562,N_14741);
nor U15271 (N_15271,N_14857,N_14630);
nand U15272 (N_15272,N_14607,N_14571);
xor U15273 (N_15273,N_14652,N_14828);
nand U15274 (N_15274,N_14561,N_14525);
nand U15275 (N_15275,N_14946,N_14877);
nor U15276 (N_15276,N_14914,N_14976);
xnor U15277 (N_15277,N_14693,N_14964);
or U15278 (N_15278,N_14904,N_14548);
or U15279 (N_15279,N_14674,N_14592);
and U15280 (N_15280,N_14754,N_14591);
xor U15281 (N_15281,N_14722,N_14865);
nand U15282 (N_15282,N_14859,N_14870);
nor U15283 (N_15283,N_14545,N_14670);
nand U15284 (N_15284,N_14746,N_14693);
nand U15285 (N_15285,N_14796,N_14633);
or U15286 (N_15286,N_14901,N_14708);
or U15287 (N_15287,N_14569,N_14829);
xnor U15288 (N_15288,N_14600,N_14564);
and U15289 (N_15289,N_14967,N_14976);
and U15290 (N_15290,N_14631,N_14938);
nor U15291 (N_15291,N_14553,N_14564);
and U15292 (N_15292,N_14932,N_14631);
nand U15293 (N_15293,N_14546,N_14542);
nor U15294 (N_15294,N_14976,N_14699);
xnor U15295 (N_15295,N_14674,N_14668);
xor U15296 (N_15296,N_14827,N_14728);
nor U15297 (N_15297,N_14934,N_14965);
and U15298 (N_15298,N_14568,N_14976);
nand U15299 (N_15299,N_14935,N_14951);
and U15300 (N_15300,N_14706,N_14685);
xnor U15301 (N_15301,N_14702,N_14996);
and U15302 (N_15302,N_14589,N_14759);
or U15303 (N_15303,N_14951,N_14523);
nor U15304 (N_15304,N_14785,N_14995);
xnor U15305 (N_15305,N_14632,N_14905);
or U15306 (N_15306,N_14607,N_14723);
nand U15307 (N_15307,N_14563,N_14762);
nand U15308 (N_15308,N_14697,N_14913);
xor U15309 (N_15309,N_14857,N_14638);
nand U15310 (N_15310,N_14864,N_14669);
and U15311 (N_15311,N_14973,N_14518);
nand U15312 (N_15312,N_14530,N_14619);
xor U15313 (N_15313,N_14887,N_14908);
or U15314 (N_15314,N_14751,N_14819);
and U15315 (N_15315,N_14611,N_14897);
and U15316 (N_15316,N_14723,N_14549);
xor U15317 (N_15317,N_14514,N_14548);
nand U15318 (N_15318,N_14927,N_14645);
and U15319 (N_15319,N_14843,N_14542);
and U15320 (N_15320,N_14901,N_14597);
and U15321 (N_15321,N_14567,N_14575);
or U15322 (N_15322,N_14916,N_14901);
or U15323 (N_15323,N_14769,N_14568);
and U15324 (N_15324,N_14614,N_14505);
nand U15325 (N_15325,N_14705,N_14772);
and U15326 (N_15326,N_14577,N_14963);
xnor U15327 (N_15327,N_14897,N_14655);
xnor U15328 (N_15328,N_14809,N_14824);
or U15329 (N_15329,N_14564,N_14724);
or U15330 (N_15330,N_14633,N_14823);
nand U15331 (N_15331,N_14553,N_14503);
nand U15332 (N_15332,N_14593,N_14855);
nor U15333 (N_15333,N_14793,N_14974);
nand U15334 (N_15334,N_14726,N_14713);
or U15335 (N_15335,N_14646,N_14901);
nand U15336 (N_15336,N_14541,N_14631);
xnor U15337 (N_15337,N_14953,N_14835);
and U15338 (N_15338,N_14624,N_14763);
nand U15339 (N_15339,N_14695,N_14702);
nand U15340 (N_15340,N_14888,N_14737);
nand U15341 (N_15341,N_14835,N_14700);
and U15342 (N_15342,N_14701,N_14533);
or U15343 (N_15343,N_14770,N_14961);
xor U15344 (N_15344,N_14623,N_14603);
nor U15345 (N_15345,N_14847,N_14931);
nand U15346 (N_15346,N_14958,N_14886);
xnor U15347 (N_15347,N_14551,N_14660);
nand U15348 (N_15348,N_14872,N_14949);
or U15349 (N_15349,N_14849,N_14803);
nor U15350 (N_15350,N_14541,N_14886);
and U15351 (N_15351,N_14552,N_14561);
nor U15352 (N_15352,N_14565,N_14923);
or U15353 (N_15353,N_14927,N_14875);
or U15354 (N_15354,N_14979,N_14794);
nand U15355 (N_15355,N_14798,N_14805);
nand U15356 (N_15356,N_14940,N_14998);
and U15357 (N_15357,N_14787,N_14984);
or U15358 (N_15358,N_14657,N_14819);
nor U15359 (N_15359,N_14559,N_14540);
nor U15360 (N_15360,N_14964,N_14620);
and U15361 (N_15361,N_14696,N_14707);
or U15362 (N_15362,N_14761,N_14860);
or U15363 (N_15363,N_14526,N_14705);
or U15364 (N_15364,N_14523,N_14878);
nor U15365 (N_15365,N_14579,N_14833);
xnor U15366 (N_15366,N_14845,N_14875);
nand U15367 (N_15367,N_14771,N_14772);
nand U15368 (N_15368,N_14999,N_14560);
or U15369 (N_15369,N_14785,N_14754);
or U15370 (N_15370,N_14729,N_14821);
and U15371 (N_15371,N_14505,N_14557);
and U15372 (N_15372,N_14665,N_14725);
and U15373 (N_15373,N_14797,N_14732);
xnor U15374 (N_15374,N_14556,N_14593);
nor U15375 (N_15375,N_14746,N_14582);
nand U15376 (N_15376,N_14953,N_14719);
nor U15377 (N_15377,N_14563,N_14901);
nand U15378 (N_15378,N_14772,N_14544);
xor U15379 (N_15379,N_14566,N_14660);
and U15380 (N_15380,N_14536,N_14896);
nand U15381 (N_15381,N_14796,N_14573);
nor U15382 (N_15382,N_14542,N_14512);
and U15383 (N_15383,N_14525,N_14601);
nand U15384 (N_15384,N_14743,N_14913);
nand U15385 (N_15385,N_14555,N_14877);
xnor U15386 (N_15386,N_14978,N_14760);
nor U15387 (N_15387,N_14571,N_14806);
nand U15388 (N_15388,N_14802,N_14820);
xnor U15389 (N_15389,N_14598,N_14683);
or U15390 (N_15390,N_14942,N_14860);
nor U15391 (N_15391,N_14662,N_14807);
nor U15392 (N_15392,N_14669,N_14678);
xor U15393 (N_15393,N_14898,N_14806);
or U15394 (N_15394,N_14991,N_14935);
or U15395 (N_15395,N_14833,N_14742);
or U15396 (N_15396,N_14581,N_14685);
or U15397 (N_15397,N_14796,N_14724);
and U15398 (N_15398,N_14744,N_14712);
xor U15399 (N_15399,N_14748,N_14701);
and U15400 (N_15400,N_14840,N_14674);
and U15401 (N_15401,N_14549,N_14645);
or U15402 (N_15402,N_14890,N_14772);
xnor U15403 (N_15403,N_14640,N_14619);
or U15404 (N_15404,N_14797,N_14716);
or U15405 (N_15405,N_14560,N_14818);
xnor U15406 (N_15406,N_14796,N_14758);
and U15407 (N_15407,N_14781,N_14624);
or U15408 (N_15408,N_14606,N_14944);
nor U15409 (N_15409,N_14733,N_14932);
nor U15410 (N_15410,N_14810,N_14760);
xor U15411 (N_15411,N_14721,N_14686);
nand U15412 (N_15412,N_14943,N_14795);
xnor U15413 (N_15413,N_14951,N_14604);
and U15414 (N_15414,N_14596,N_14832);
nand U15415 (N_15415,N_14813,N_14539);
or U15416 (N_15416,N_14832,N_14644);
or U15417 (N_15417,N_14930,N_14821);
and U15418 (N_15418,N_14897,N_14550);
and U15419 (N_15419,N_14850,N_14683);
nand U15420 (N_15420,N_14845,N_14628);
or U15421 (N_15421,N_14767,N_14827);
and U15422 (N_15422,N_14951,N_14680);
or U15423 (N_15423,N_14984,N_14888);
nand U15424 (N_15424,N_14583,N_14703);
or U15425 (N_15425,N_14769,N_14976);
or U15426 (N_15426,N_14998,N_14793);
nand U15427 (N_15427,N_14646,N_14876);
nand U15428 (N_15428,N_14732,N_14851);
xnor U15429 (N_15429,N_14580,N_14900);
nor U15430 (N_15430,N_14864,N_14950);
xnor U15431 (N_15431,N_14752,N_14928);
nor U15432 (N_15432,N_14819,N_14983);
or U15433 (N_15433,N_14781,N_14744);
nor U15434 (N_15434,N_14617,N_14918);
or U15435 (N_15435,N_14777,N_14688);
nand U15436 (N_15436,N_14871,N_14662);
and U15437 (N_15437,N_14984,N_14791);
nand U15438 (N_15438,N_14635,N_14785);
or U15439 (N_15439,N_14742,N_14696);
nor U15440 (N_15440,N_14895,N_14526);
or U15441 (N_15441,N_14913,N_14717);
and U15442 (N_15442,N_14997,N_14821);
xnor U15443 (N_15443,N_14810,N_14603);
xnor U15444 (N_15444,N_14804,N_14714);
xnor U15445 (N_15445,N_14701,N_14534);
and U15446 (N_15446,N_14897,N_14927);
or U15447 (N_15447,N_14512,N_14828);
and U15448 (N_15448,N_14784,N_14836);
or U15449 (N_15449,N_14947,N_14545);
and U15450 (N_15450,N_14753,N_14620);
or U15451 (N_15451,N_14578,N_14657);
nand U15452 (N_15452,N_14591,N_14881);
or U15453 (N_15453,N_14598,N_14919);
and U15454 (N_15454,N_14855,N_14933);
nor U15455 (N_15455,N_14556,N_14666);
nand U15456 (N_15456,N_14930,N_14919);
nor U15457 (N_15457,N_14639,N_14845);
and U15458 (N_15458,N_14864,N_14820);
nand U15459 (N_15459,N_14688,N_14698);
nand U15460 (N_15460,N_14813,N_14718);
or U15461 (N_15461,N_14764,N_14712);
nor U15462 (N_15462,N_14590,N_14700);
and U15463 (N_15463,N_14718,N_14762);
xnor U15464 (N_15464,N_14810,N_14563);
xnor U15465 (N_15465,N_14983,N_14894);
and U15466 (N_15466,N_14957,N_14594);
and U15467 (N_15467,N_14754,N_14668);
xor U15468 (N_15468,N_14904,N_14686);
and U15469 (N_15469,N_14875,N_14761);
and U15470 (N_15470,N_14971,N_14843);
xor U15471 (N_15471,N_14727,N_14769);
nor U15472 (N_15472,N_14952,N_14719);
xnor U15473 (N_15473,N_14732,N_14605);
nor U15474 (N_15474,N_14574,N_14597);
and U15475 (N_15475,N_14851,N_14601);
nand U15476 (N_15476,N_14803,N_14810);
nand U15477 (N_15477,N_14836,N_14799);
and U15478 (N_15478,N_14547,N_14952);
nor U15479 (N_15479,N_14657,N_14502);
nand U15480 (N_15480,N_14819,N_14772);
nor U15481 (N_15481,N_14620,N_14507);
nor U15482 (N_15482,N_14941,N_14624);
xnor U15483 (N_15483,N_14614,N_14901);
and U15484 (N_15484,N_14937,N_14628);
and U15485 (N_15485,N_14620,N_14849);
xor U15486 (N_15486,N_14975,N_14910);
nor U15487 (N_15487,N_14806,N_14919);
xor U15488 (N_15488,N_14772,N_14859);
or U15489 (N_15489,N_14737,N_14980);
or U15490 (N_15490,N_14655,N_14682);
nand U15491 (N_15491,N_14821,N_14537);
nor U15492 (N_15492,N_14838,N_14688);
and U15493 (N_15493,N_14654,N_14581);
xnor U15494 (N_15494,N_14921,N_14713);
and U15495 (N_15495,N_14849,N_14955);
xor U15496 (N_15496,N_14951,N_14750);
xor U15497 (N_15497,N_14816,N_14880);
nand U15498 (N_15498,N_14552,N_14873);
nor U15499 (N_15499,N_14521,N_14585);
and U15500 (N_15500,N_15249,N_15018);
nand U15501 (N_15501,N_15009,N_15488);
nor U15502 (N_15502,N_15479,N_15276);
nor U15503 (N_15503,N_15057,N_15355);
or U15504 (N_15504,N_15275,N_15152);
xnor U15505 (N_15505,N_15281,N_15243);
xor U15506 (N_15506,N_15215,N_15196);
or U15507 (N_15507,N_15201,N_15138);
or U15508 (N_15508,N_15239,N_15484);
or U15509 (N_15509,N_15208,N_15042);
nand U15510 (N_15510,N_15133,N_15336);
nand U15511 (N_15511,N_15012,N_15106);
and U15512 (N_15512,N_15376,N_15418);
nor U15513 (N_15513,N_15467,N_15000);
nor U15514 (N_15514,N_15121,N_15309);
or U15515 (N_15515,N_15314,N_15225);
and U15516 (N_15516,N_15465,N_15036);
nor U15517 (N_15517,N_15037,N_15011);
nor U15518 (N_15518,N_15289,N_15401);
or U15519 (N_15519,N_15450,N_15179);
or U15520 (N_15520,N_15245,N_15293);
nor U15521 (N_15521,N_15282,N_15188);
nand U15522 (N_15522,N_15260,N_15415);
and U15523 (N_15523,N_15395,N_15206);
nor U15524 (N_15524,N_15257,N_15204);
nor U15525 (N_15525,N_15217,N_15186);
xnor U15526 (N_15526,N_15396,N_15246);
nand U15527 (N_15527,N_15406,N_15124);
nand U15528 (N_15528,N_15177,N_15081);
nor U15529 (N_15529,N_15040,N_15344);
xor U15530 (N_15530,N_15187,N_15471);
nand U15531 (N_15531,N_15420,N_15279);
xor U15532 (N_15532,N_15075,N_15034);
and U15533 (N_15533,N_15097,N_15176);
nor U15534 (N_15534,N_15297,N_15445);
xor U15535 (N_15535,N_15024,N_15178);
or U15536 (N_15536,N_15154,N_15033);
or U15537 (N_15537,N_15308,N_15094);
or U15538 (N_15538,N_15291,N_15301);
nand U15539 (N_15539,N_15014,N_15359);
xor U15540 (N_15540,N_15356,N_15302);
xnor U15541 (N_15541,N_15425,N_15227);
nor U15542 (N_15542,N_15161,N_15270);
nand U15543 (N_15543,N_15210,N_15140);
nor U15544 (N_15544,N_15258,N_15262);
xor U15545 (N_15545,N_15168,N_15323);
xnor U15546 (N_15546,N_15459,N_15429);
nor U15547 (N_15547,N_15424,N_15170);
and U15548 (N_15548,N_15159,N_15393);
nand U15549 (N_15549,N_15489,N_15167);
and U15550 (N_15550,N_15280,N_15101);
or U15551 (N_15551,N_15151,N_15329);
and U15552 (N_15552,N_15253,N_15416);
or U15553 (N_15553,N_15076,N_15205);
or U15554 (N_15554,N_15322,N_15470);
and U15555 (N_15555,N_15242,N_15050);
or U15556 (N_15556,N_15362,N_15345);
nor U15557 (N_15557,N_15383,N_15238);
xor U15558 (N_15558,N_15126,N_15248);
nor U15559 (N_15559,N_15122,N_15043);
nor U15560 (N_15560,N_15372,N_15147);
or U15561 (N_15561,N_15026,N_15377);
or U15562 (N_15562,N_15473,N_15093);
or U15563 (N_15563,N_15194,N_15234);
nor U15564 (N_15564,N_15296,N_15495);
nor U15565 (N_15565,N_15137,N_15364);
nor U15566 (N_15566,N_15305,N_15386);
nand U15567 (N_15567,N_15221,N_15318);
nand U15568 (N_15568,N_15353,N_15062);
nor U15569 (N_15569,N_15265,N_15095);
and U15570 (N_15570,N_15430,N_15369);
xor U15571 (N_15571,N_15405,N_15378);
nand U15572 (N_15572,N_15190,N_15426);
xor U15573 (N_15573,N_15013,N_15385);
nand U15574 (N_15574,N_15273,N_15340);
xnor U15575 (N_15575,N_15368,N_15320);
nor U15576 (N_15576,N_15351,N_15358);
xnor U15577 (N_15577,N_15398,N_15422);
and U15578 (N_15578,N_15255,N_15472);
nand U15579 (N_15579,N_15145,N_15163);
xnor U15580 (N_15580,N_15001,N_15419);
nand U15581 (N_15581,N_15123,N_15046);
nor U15582 (N_15582,N_15494,N_15021);
xnor U15583 (N_15583,N_15141,N_15496);
or U15584 (N_15584,N_15115,N_15028);
xnor U15585 (N_15585,N_15328,N_15098);
nor U15586 (N_15586,N_15113,N_15071);
nor U15587 (N_15587,N_15016,N_15118);
and U15588 (N_15588,N_15454,N_15051);
xor U15589 (N_15589,N_15338,N_15226);
nand U15590 (N_15590,N_15212,N_15108);
and U15591 (N_15591,N_15294,N_15413);
and U15592 (N_15592,N_15144,N_15209);
or U15593 (N_15593,N_15149,N_15084);
and U15594 (N_15594,N_15184,N_15300);
or U15595 (N_15595,N_15035,N_15223);
nand U15596 (N_15596,N_15200,N_15380);
or U15597 (N_15597,N_15499,N_15290);
xnor U15598 (N_15598,N_15409,N_15441);
or U15599 (N_15599,N_15072,N_15131);
nand U15600 (N_15600,N_15049,N_15211);
xnor U15601 (N_15601,N_15158,N_15236);
and U15602 (N_15602,N_15174,N_15082);
xor U15603 (N_15603,N_15363,N_15327);
xor U15604 (N_15604,N_15411,N_15460);
and U15605 (N_15605,N_15218,N_15224);
xnor U15606 (N_15606,N_15132,N_15397);
and U15607 (N_15607,N_15483,N_15102);
nor U15608 (N_15608,N_15352,N_15462);
nand U15609 (N_15609,N_15134,N_15143);
and U15610 (N_15610,N_15475,N_15304);
nand U15611 (N_15611,N_15442,N_15354);
or U15612 (N_15612,N_15423,N_15182);
and U15613 (N_15613,N_15172,N_15216);
and U15614 (N_15614,N_15349,N_15259);
nor U15615 (N_15615,N_15185,N_15490);
nor U15616 (N_15616,N_15414,N_15180);
nor U15617 (N_15617,N_15015,N_15432);
and U15618 (N_15618,N_15402,N_15031);
nand U15619 (N_15619,N_15434,N_15162);
and U15620 (N_15620,N_15023,N_15100);
nor U15621 (N_15621,N_15065,N_15464);
nor U15622 (N_15622,N_15346,N_15319);
nand U15623 (N_15623,N_15417,N_15153);
nor U15624 (N_15624,N_15099,N_15456);
or U15625 (N_15625,N_15271,N_15285);
nor U15626 (N_15626,N_15148,N_15222);
or U15627 (N_15627,N_15466,N_15444);
or U15628 (N_15628,N_15335,N_15019);
nor U15629 (N_15629,N_15437,N_15128);
nor U15630 (N_15630,N_15191,N_15261);
and U15631 (N_15631,N_15142,N_15321);
nand U15632 (N_15632,N_15135,N_15292);
and U15633 (N_15633,N_15017,N_15427);
or U15634 (N_15634,N_15350,N_15111);
xnor U15635 (N_15635,N_15474,N_15244);
nand U15636 (N_15636,N_15348,N_15008);
nor U15637 (N_15637,N_15461,N_15087);
nand U15638 (N_15638,N_15375,N_15139);
nand U15639 (N_15639,N_15384,N_15054);
nand U15640 (N_15640,N_15056,N_15400);
nand U15641 (N_15641,N_15478,N_15029);
and U15642 (N_15642,N_15298,N_15315);
or U15643 (N_15643,N_15286,N_15130);
nor U15644 (N_15644,N_15371,N_15195);
nor U15645 (N_15645,N_15391,N_15250);
xnor U15646 (N_15646,N_15252,N_15090);
and U15647 (N_15647,N_15127,N_15404);
or U15648 (N_15648,N_15433,N_15160);
xnor U15649 (N_15649,N_15078,N_15272);
nor U15650 (N_15650,N_15324,N_15455);
and U15651 (N_15651,N_15005,N_15480);
or U15652 (N_15652,N_15337,N_15256);
or U15653 (N_15653,N_15477,N_15197);
or U15654 (N_15654,N_15183,N_15379);
nand U15655 (N_15655,N_15171,N_15213);
and U15656 (N_15656,N_15096,N_15310);
nor U15657 (N_15657,N_15498,N_15267);
xnor U15658 (N_15658,N_15476,N_15447);
nand U15659 (N_15659,N_15408,N_15365);
or U15660 (N_15660,N_15347,N_15463);
nand U15661 (N_15661,N_15333,N_15313);
or U15662 (N_15662,N_15482,N_15073);
xor U15663 (N_15663,N_15357,N_15435);
and U15664 (N_15664,N_15045,N_15164);
nand U15665 (N_15665,N_15436,N_15020);
nand U15666 (N_15666,N_15278,N_15287);
nor U15667 (N_15667,N_15083,N_15214);
nor U15668 (N_15668,N_15058,N_15193);
xor U15669 (N_15669,N_15374,N_15146);
nor U15670 (N_15670,N_15388,N_15104);
nand U15671 (N_15671,N_15202,N_15030);
xor U15672 (N_15672,N_15006,N_15264);
or U15673 (N_15673,N_15230,N_15175);
xor U15674 (N_15674,N_15064,N_15361);
and U15675 (N_15675,N_15306,N_15277);
and U15676 (N_15676,N_15370,N_15317);
or U15677 (N_15677,N_15284,N_15063);
and U15678 (N_15678,N_15247,N_15325);
nor U15679 (N_15679,N_15241,N_15399);
nand U15680 (N_15680,N_15240,N_15382);
nand U15681 (N_15681,N_15440,N_15055);
nor U15682 (N_15682,N_15039,N_15449);
nand U15683 (N_15683,N_15032,N_15228);
or U15684 (N_15684,N_15068,N_15198);
xnor U15685 (N_15685,N_15091,N_15189);
nor U15686 (N_15686,N_15231,N_15166);
and U15687 (N_15687,N_15157,N_15403);
nor U15688 (N_15688,N_15468,N_15390);
and U15689 (N_15689,N_15199,N_15116);
nor U15690 (N_15690,N_15085,N_15169);
and U15691 (N_15691,N_15077,N_15458);
and U15692 (N_15692,N_15394,N_15129);
or U15693 (N_15693,N_15112,N_15339);
or U15694 (N_15694,N_15469,N_15343);
and U15695 (N_15695,N_15366,N_15497);
or U15696 (N_15696,N_15254,N_15446);
or U15697 (N_15697,N_15004,N_15079);
and U15698 (N_15698,N_15181,N_15453);
xor U15699 (N_15699,N_15010,N_15220);
and U15700 (N_15700,N_15047,N_15105);
and U15701 (N_15701,N_15038,N_15451);
xnor U15702 (N_15702,N_15114,N_15491);
and U15703 (N_15703,N_15070,N_15235);
xor U15704 (N_15704,N_15269,N_15412);
and U15705 (N_15705,N_15207,N_15438);
and U15706 (N_15706,N_15002,N_15295);
or U15707 (N_15707,N_15069,N_15237);
xnor U15708 (N_15708,N_15203,N_15150);
xor U15709 (N_15709,N_15263,N_15229);
nand U15710 (N_15710,N_15092,N_15251);
nor U15711 (N_15711,N_15155,N_15332);
and U15712 (N_15712,N_15312,N_15331);
and U15713 (N_15713,N_15311,N_15316);
nor U15714 (N_15714,N_15274,N_15088);
and U15715 (N_15715,N_15080,N_15431);
and U15716 (N_15716,N_15299,N_15059);
xnor U15717 (N_15717,N_15410,N_15120);
and U15718 (N_15718,N_15443,N_15367);
or U15719 (N_15719,N_15334,N_15044);
and U15720 (N_15720,N_15330,N_15117);
and U15721 (N_15721,N_15428,N_15452);
xnor U15722 (N_15722,N_15041,N_15389);
and U15723 (N_15723,N_15448,N_15439);
and U15724 (N_15724,N_15003,N_15481);
or U15725 (N_15725,N_15341,N_15342);
nand U15726 (N_15726,N_15283,N_15407);
or U15727 (N_15727,N_15074,N_15486);
and U15728 (N_15728,N_15067,N_15303);
nand U15729 (N_15729,N_15119,N_15136);
or U15730 (N_15730,N_15027,N_15232);
xnor U15731 (N_15731,N_15061,N_15156);
nor U15732 (N_15732,N_15219,N_15485);
nor U15733 (N_15733,N_15052,N_15487);
xnor U15734 (N_15734,N_15066,N_15268);
xnor U15735 (N_15735,N_15421,N_15103);
nor U15736 (N_15736,N_15007,N_15025);
nor U15737 (N_15737,N_15060,N_15125);
nand U15738 (N_15738,N_15307,N_15048);
nor U15739 (N_15739,N_15089,N_15381);
nor U15740 (N_15740,N_15493,N_15109);
or U15741 (N_15741,N_15266,N_15233);
nor U15742 (N_15742,N_15165,N_15022);
xor U15743 (N_15743,N_15107,N_15086);
or U15744 (N_15744,N_15387,N_15288);
nand U15745 (N_15745,N_15492,N_15173);
nor U15746 (N_15746,N_15326,N_15192);
and U15747 (N_15747,N_15053,N_15360);
or U15748 (N_15748,N_15457,N_15373);
or U15749 (N_15749,N_15110,N_15392);
or U15750 (N_15750,N_15409,N_15394);
and U15751 (N_15751,N_15443,N_15436);
xnor U15752 (N_15752,N_15281,N_15069);
and U15753 (N_15753,N_15018,N_15314);
nand U15754 (N_15754,N_15497,N_15013);
nor U15755 (N_15755,N_15003,N_15420);
nand U15756 (N_15756,N_15320,N_15287);
nand U15757 (N_15757,N_15254,N_15216);
and U15758 (N_15758,N_15402,N_15214);
nand U15759 (N_15759,N_15463,N_15301);
nor U15760 (N_15760,N_15307,N_15364);
nand U15761 (N_15761,N_15023,N_15226);
xnor U15762 (N_15762,N_15058,N_15252);
nand U15763 (N_15763,N_15394,N_15422);
and U15764 (N_15764,N_15418,N_15018);
nand U15765 (N_15765,N_15405,N_15376);
xnor U15766 (N_15766,N_15260,N_15035);
nor U15767 (N_15767,N_15281,N_15276);
nand U15768 (N_15768,N_15481,N_15305);
xor U15769 (N_15769,N_15256,N_15303);
xnor U15770 (N_15770,N_15005,N_15396);
or U15771 (N_15771,N_15347,N_15187);
nand U15772 (N_15772,N_15289,N_15113);
and U15773 (N_15773,N_15496,N_15194);
or U15774 (N_15774,N_15129,N_15419);
and U15775 (N_15775,N_15147,N_15141);
nor U15776 (N_15776,N_15121,N_15097);
or U15777 (N_15777,N_15321,N_15104);
or U15778 (N_15778,N_15169,N_15325);
nor U15779 (N_15779,N_15254,N_15057);
nand U15780 (N_15780,N_15317,N_15112);
and U15781 (N_15781,N_15030,N_15219);
nor U15782 (N_15782,N_15347,N_15138);
nor U15783 (N_15783,N_15332,N_15450);
nor U15784 (N_15784,N_15393,N_15278);
and U15785 (N_15785,N_15244,N_15487);
nor U15786 (N_15786,N_15342,N_15151);
nand U15787 (N_15787,N_15258,N_15364);
nor U15788 (N_15788,N_15075,N_15458);
nor U15789 (N_15789,N_15034,N_15250);
nor U15790 (N_15790,N_15483,N_15112);
and U15791 (N_15791,N_15016,N_15389);
or U15792 (N_15792,N_15433,N_15223);
xor U15793 (N_15793,N_15127,N_15315);
xor U15794 (N_15794,N_15482,N_15263);
xnor U15795 (N_15795,N_15329,N_15178);
nor U15796 (N_15796,N_15037,N_15118);
xor U15797 (N_15797,N_15487,N_15208);
nand U15798 (N_15798,N_15029,N_15073);
nor U15799 (N_15799,N_15329,N_15063);
nand U15800 (N_15800,N_15051,N_15212);
nand U15801 (N_15801,N_15045,N_15086);
xnor U15802 (N_15802,N_15190,N_15367);
or U15803 (N_15803,N_15293,N_15027);
or U15804 (N_15804,N_15366,N_15161);
and U15805 (N_15805,N_15380,N_15094);
and U15806 (N_15806,N_15061,N_15377);
xor U15807 (N_15807,N_15382,N_15171);
nor U15808 (N_15808,N_15403,N_15089);
nand U15809 (N_15809,N_15108,N_15231);
xor U15810 (N_15810,N_15043,N_15356);
or U15811 (N_15811,N_15111,N_15241);
nor U15812 (N_15812,N_15155,N_15038);
or U15813 (N_15813,N_15183,N_15263);
and U15814 (N_15814,N_15354,N_15101);
nand U15815 (N_15815,N_15399,N_15210);
or U15816 (N_15816,N_15284,N_15408);
or U15817 (N_15817,N_15316,N_15111);
nand U15818 (N_15818,N_15392,N_15464);
and U15819 (N_15819,N_15257,N_15402);
xnor U15820 (N_15820,N_15155,N_15218);
nand U15821 (N_15821,N_15374,N_15430);
and U15822 (N_15822,N_15447,N_15282);
nand U15823 (N_15823,N_15080,N_15122);
and U15824 (N_15824,N_15198,N_15360);
or U15825 (N_15825,N_15447,N_15431);
and U15826 (N_15826,N_15052,N_15047);
xor U15827 (N_15827,N_15125,N_15161);
or U15828 (N_15828,N_15340,N_15000);
xnor U15829 (N_15829,N_15380,N_15382);
nor U15830 (N_15830,N_15105,N_15021);
or U15831 (N_15831,N_15143,N_15073);
and U15832 (N_15832,N_15008,N_15411);
or U15833 (N_15833,N_15461,N_15033);
xnor U15834 (N_15834,N_15309,N_15246);
or U15835 (N_15835,N_15094,N_15317);
nand U15836 (N_15836,N_15148,N_15427);
nand U15837 (N_15837,N_15235,N_15403);
or U15838 (N_15838,N_15466,N_15146);
nor U15839 (N_15839,N_15388,N_15048);
nand U15840 (N_15840,N_15388,N_15316);
and U15841 (N_15841,N_15429,N_15229);
and U15842 (N_15842,N_15158,N_15329);
xnor U15843 (N_15843,N_15383,N_15100);
nor U15844 (N_15844,N_15094,N_15086);
and U15845 (N_15845,N_15378,N_15400);
or U15846 (N_15846,N_15263,N_15035);
and U15847 (N_15847,N_15023,N_15025);
and U15848 (N_15848,N_15306,N_15085);
xor U15849 (N_15849,N_15055,N_15108);
nand U15850 (N_15850,N_15039,N_15152);
and U15851 (N_15851,N_15253,N_15163);
or U15852 (N_15852,N_15197,N_15493);
or U15853 (N_15853,N_15377,N_15163);
and U15854 (N_15854,N_15117,N_15140);
nand U15855 (N_15855,N_15228,N_15327);
nand U15856 (N_15856,N_15319,N_15071);
and U15857 (N_15857,N_15170,N_15198);
nor U15858 (N_15858,N_15451,N_15239);
nand U15859 (N_15859,N_15035,N_15018);
and U15860 (N_15860,N_15223,N_15105);
or U15861 (N_15861,N_15257,N_15040);
nand U15862 (N_15862,N_15360,N_15088);
xnor U15863 (N_15863,N_15483,N_15387);
or U15864 (N_15864,N_15349,N_15019);
and U15865 (N_15865,N_15479,N_15135);
and U15866 (N_15866,N_15207,N_15378);
nand U15867 (N_15867,N_15228,N_15356);
or U15868 (N_15868,N_15098,N_15055);
or U15869 (N_15869,N_15142,N_15165);
and U15870 (N_15870,N_15385,N_15374);
or U15871 (N_15871,N_15479,N_15271);
and U15872 (N_15872,N_15141,N_15211);
or U15873 (N_15873,N_15368,N_15139);
or U15874 (N_15874,N_15091,N_15188);
and U15875 (N_15875,N_15129,N_15259);
nor U15876 (N_15876,N_15365,N_15299);
xnor U15877 (N_15877,N_15191,N_15243);
and U15878 (N_15878,N_15306,N_15075);
or U15879 (N_15879,N_15125,N_15388);
nand U15880 (N_15880,N_15321,N_15337);
nor U15881 (N_15881,N_15480,N_15308);
or U15882 (N_15882,N_15307,N_15176);
xnor U15883 (N_15883,N_15308,N_15111);
or U15884 (N_15884,N_15165,N_15039);
nand U15885 (N_15885,N_15184,N_15239);
xnor U15886 (N_15886,N_15369,N_15209);
or U15887 (N_15887,N_15410,N_15192);
or U15888 (N_15888,N_15440,N_15459);
or U15889 (N_15889,N_15028,N_15110);
nor U15890 (N_15890,N_15098,N_15292);
or U15891 (N_15891,N_15472,N_15424);
nor U15892 (N_15892,N_15278,N_15342);
nor U15893 (N_15893,N_15284,N_15020);
and U15894 (N_15894,N_15286,N_15037);
nand U15895 (N_15895,N_15429,N_15148);
or U15896 (N_15896,N_15415,N_15023);
nor U15897 (N_15897,N_15496,N_15246);
and U15898 (N_15898,N_15328,N_15202);
xor U15899 (N_15899,N_15433,N_15203);
nand U15900 (N_15900,N_15200,N_15096);
xnor U15901 (N_15901,N_15092,N_15429);
nand U15902 (N_15902,N_15038,N_15337);
nand U15903 (N_15903,N_15129,N_15140);
nor U15904 (N_15904,N_15260,N_15257);
and U15905 (N_15905,N_15480,N_15090);
or U15906 (N_15906,N_15355,N_15185);
xnor U15907 (N_15907,N_15190,N_15152);
xnor U15908 (N_15908,N_15009,N_15096);
and U15909 (N_15909,N_15105,N_15446);
or U15910 (N_15910,N_15452,N_15271);
nand U15911 (N_15911,N_15462,N_15145);
or U15912 (N_15912,N_15012,N_15198);
and U15913 (N_15913,N_15434,N_15157);
nand U15914 (N_15914,N_15156,N_15233);
or U15915 (N_15915,N_15001,N_15403);
xor U15916 (N_15916,N_15444,N_15021);
or U15917 (N_15917,N_15232,N_15191);
or U15918 (N_15918,N_15409,N_15312);
nor U15919 (N_15919,N_15164,N_15287);
and U15920 (N_15920,N_15253,N_15475);
nor U15921 (N_15921,N_15316,N_15079);
or U15922 (N_15922,N_15349,N_15230);
and U15923 (N_15923,N_15057,N_15451);
nor U15924 (N_15924,N_15053,N_15406);
nand U15925 (N_15925,N_15445,N_15155);
xnor U15926 (N_15926,N_15433,N_15122);
xnor U15927 (N_15927,N_15499,N_15257);
or U15928 (N_15928,N_15409,N_15135);
and U15929 (N_15929,N_15404,N_15106);
and U15930 (N_15930,N_15356,N_15079);
nor U15931 (N_15931,N_15206,N_15455);
or U15932 (N_15932,N_15429,N_15050);
xnor U15933 (N_15933,N_15201,N_15392);
and U15934 (N_15934,N_15406,N_15334);
xnor U15935 (N_15935,N_15231,N_15317);
or U15936 (N_15936,N_15039,N_15304);
and U15937 (N_15937,N_15001,N_15154);
or U15938 (N_15938,N_15204,N_15212);
nor U15939 (N_15939,N_15111,N_15383);
or U15940 (N_15940,N_15151,N_15254);
and U15941 (N_15941,N_15034,N_15145);
and U15942 (N_15942,N_15377,N_15336);
nor U15943 (N_15943,N_15412,N_15210);
or U15944 (N_15944,N_15004,N_15284);
xnor U15945 (N_15945,N_15082,N_15172);
nand U15946 (N_15946,N_15080,N_15400);
nor U15947 (N_15947,N_15088,N_15285);
nor U15948 (N_15948,N_15055,N_15423);
nor U15949 (N_15949,N_15377,N_15207);
nand U15950 (N_15950,N_15164,N_15335);
nand U15951 (N_15951,N_15390,N_15180);
xnor U15952 (N_15952,N_15349,N_15417);
xnor U15953 (N_15953,N_15075,N_15149);
nand U15954 (N_15954,N_15162,N_15330);
nor U15955 (N_15955,N_15050,N_15399);
and U15956 (N_15956,N_15038,N_15272);
or U15957 (N_15957,N_15084,N_15408);
xor U15958 (N_15958,N_15495,N_15027);
or U15959 (N_15959,N_15420,N_15303);
and U15960 (N_15960,N_15344,N_15386);
nand U15961 (N_15961,N_15408,N_15305);
nor U15962 (N_15962,N_15248,N_15141);
or U15963 (N_15963,N_15177,N_15028);
nor U15964 (N_15964,N_15022,N_15284);
nor U15965 (N_15965,N_15343,N_15195);
nor U15966 (N_15966,N_15119,N_15384);
nor U15967 (N_15967,N_15437,N_15226);
xor U15968 (N_15968,N_15150,N_15494);
nand U15969 (N_15969,N_15120,N_15169);
xnor U15970 (N_15970,N_15328,N_15480);
nand U15971 (N_15971,N_15296,N_15470);
nor U15972 (N_15972,N_15307,N_15284);
xor U15973 (N_15973,N_15338,N_15358);
and U15974 (N_15974,N_15034,N_15185);
nor U15975 (N_15975,N_15224,N_15482);
and U15976 (N_15976,N_15406,N_15057);
xnor U15977 (N_15977,N_15175,N_15344);
nand U15978 (N_15978,N_15463,N_15304);
xor U15979 (N_15979,N_15485,N_15302);
nand U15980 (N_15980,N_15132,N_15471);
or U15981 (N_15981,N_15370,N_15334);
xor U15982 (N_15982,N_15495,N_15070);
xnor U15983 (N_15983,N_15100,N_15052);
and U15984 (N_15984,N_15439,N_15145);
nor U15985 (N_15985,N_15249,N_15180);
nand U15986 (N_15986,N_15116,N_15235);
xnor U15987 (N_15987,N_15261,N_15055);
or U15988 (N_15988,N_15037,N_15030);
and U15989 (N_15989,N_15414,N_15436);
nor U15990 (N_15990,N_15085,N_15019);
xor U15991 (N_15991,N_15185,N_15007);
or U15992 (N_15992,N_15463,N_15092);
nor U15993 (N_15993,N_15391,N_15149);
nand U15994 (N_15994,N_15174,N_15301);
and U15995 (N_15995,N_15035,N_15137);
and U15996 (N_15996,N_15464,N_15282);
nor U15997 (N_15997,N_15317,N_15326);
xor U15998 (N_15998,N_15400,N_15245);
nor U15999 (N_15999,N_15012,N_15400);
and U16000 (N_16000,N_15914,N_15981);
nand U16001 (N_16001,N_15931,N_15696);
nor U16002 (N_16002,N_15978,N_15602);
nand U16003 (N_16003,N_15884,N_15895);
or U16004 (N_16004,N_15578,N_15718);
and U16005 (N_16005,N_15804,N_15891);
nor U16006 (N_16006,N_15692,N_15947);
nand U16007 (N_16007,N_15669,N_15663);
nor U16008 (N_16008,N_15882,N_15883);
xnor U16009 (N_16009,N_15561,N_15666);
nand U16010 (N_16010,N_15705,N_15542);
or U16011 (N_16011,N_15592,N_15509);
nor U16012 (N_16012,N_15852,N_15969);
xnor U16013 (N_16013,N_15965,N_15876);
nand U16014 (N_16014,N_15620,N_15778);
and U16015 (N_16015,N_15880,N_15904);
nor U16016 (N_16016,N_15789,N_15552);
or U16017 (N_16017,N_15942,N_15512);
and U16018 (N_16018,N_15672,N_15707);
nand U16019 (N_16019,N_15694,N_15656);
nand U16020 (N_16020,N_15511,N_15745);
or U16021 (N_16021,N_15953,N_15861);
xor U16022 (N_16022,N_15689,N_15564);
xnor U16023 (N_16023,N_15715,N_15554);
xor U16024 (N_16024,N_15830,N_15783);
nor U16025 (N_16025,N_15649,N_15526);
nand U16026 (N_16026,N_15684,N_15950);
nor U16027 (N_16027,N_15614,N_15651);
xnor U16028 (N_16028,N_15836,N_15762);
and U16029 (N_16029,N_15648,N_15647);
or U16030 (N_16030,N_15779,N_15749);
nand U16031 (N_16031,N_15945,N_15726);
xor U16032 (N_16032,N_15626,N_15844);
nor U16033 (N_16033,N_15834,N_15679);
xnor U16034 (N_16034,N_15577,N_15551);
nor U16035 (N_16035,N_15941,N_15784);
and U16036 (N_16036,N_15714,N_15719);
and U16037 (N_16037,N_15706,N_15608);
nand U16038 (N_16038,N_15553,N_15898);
nand U16039 (N_16039,N_15801,N_15951);
xnor U16040 (N_16040,N_15522,N_15536);
and U16041 (N_16041,N_15655,N_15916);
nor U16042 (N_16042,N_15865,N_15675);
nor U16043 (N_16043,N_15510,N_15806);
nand U16044 (N_16044,N_15514,N_15579);
or U16045 (N_16045,N_15671,N_15757);
nor U16046 (N_16046,N_15567,N_15917);
xnor U16047 (N_16047,N_15535,N_15847);
and U16048 (N_16048,N_15767,N_15559);
xnor U16049 (N_16049,N_15868,N_15973);
xnor U16050 (N_16050,N_15777,N_15831);
xnor U16051 (N_16051,N_15869,N_15710);
nand U16052 (N_16052,N_15576,N_15530);
xor U16053 (N_16053,N_15629,N_15738);
or U16054 (N_16054,N_15957,N_15949);
or U16055 (N_16055,N_15731,N_15538);
nor U16056 (N_16056,N_15725,N_15885);
nor U16057 (N_16057,N_15505,N_15913);
nand U16058 (N_16058,N_15839,N_15761);
and U16059 (N_16059,N_15922,N_15964);
nand U16060 (N_16060,N_15952,N_15636);
or U16061 (N_16061,N_15759,N_15686);
xor U16062 (N_16062,N_15665,N_15618);
or U16063 (N_16063,N_15585,N_15624);
nor U16064 (N_16064,N_15772,N_15703);
xor U16065 (N_16065,N_15859,N_15607);
and U16066 (N_16066,N_15874,N_15890);
nor U16067 (N_16067,N_15766,N_15625);
and U16068 (N_16068,N_15506,N_15754);
and U16069 (N_16069,N_15743,N_15637);
xnor U16070 (N_16070,N_15790,N_15643);
or U16071 (N_16071,N_15701,N_15652);
and U16072 (N_16072,N_15589,N_15716);
or U16073 (N_16073,N_15840,N_15853);
or U16074 (N_16074,N_15741,N_15590);
or U16075 (N_16075,N_15617,N_15797);
nand U16076 (N_16076,N_15593,N_15528);
or U16077 (N_16077,N_15548,N_15764);
or U16078 (N_16078,N_15918,N_15730);
and U16079 (N_16079,N_15619,N_15842);
xnor U16080 (N_16080,N_15824,N_15845);
nor U16081 (N_16081,N_15713,N_15920);
nor U16082 (N_16082,N_15747,N_15843);
xor U16083 (N_16083,N_15668,N_15992);
and U16084 (N_16084,N_15570,N_15879);
and U16085 (N_16085,N_15755,N_15888);
or U16086 (N_16086,N_15724,N_15803);
and U16087 (N_16087,N_15968,N_15582);
nand U16088 (N_16088,N_15785,N_15569);
nor U16089 (N_16089,N_15930,N_15688);
xor U16090 (N_16090,N_15899,N_15580);
or U16091 (N_16091,N_15555,N_15984);
nor U16092 (N_16092,N_15955,N_15566);
xor U16093 (N_16093,N_15596,N_15776);
and U16094 (N_16094,N_15996,N_15939);
or U16095 (N_16095,N_15961,N_15556);
and U16096 (N_16096,N_15682,N_15502);
nand U16097 (N_16097,N_15954,N_15588);
and U16098 (N_16098,N_15826,N_15537);
xor U16099 (N_16099,N_15604,N_15662);
and U16100 (N_16100,N_15832,N_15809);
or U16101 (N_16101,N_15781,N_15991);
nand U16102 (N_16102,N_15758,N_15854);
nor U16103 (N_16103,N_15721,N_15644);
nor U16104 (N_16104,N_15972,N_15595);
nor U16105 (N_16105,N_15583,N_15775);
or U16106 (N_16106,N_15900,N_15780);
nand U16107 (N_16107,N_15658,N_15875);
and U16108 (N_16108,N_15574,N_15709);
xor U16109 (N_16109,N_15599,N_15886);
or U16110 (N_16110,N_15612,N_15999);
nor U16111 (N_16111,N_15587,N_15722);
xor U16112 (N_16112,N_15687,N_15615);
and U16113 (N_16113,N_15998,N_15810);
nand U16114 (N_16114,N_15560,N_15912);
xnor U16115 (N_16115,N_15820,N_15774);
nor U16116 (N_16116,N_15645,N_15937);
and U16117 (N_16117,N_15929,N_15763);
nor U16118 (N_16118,N_15500,N_15848);
xnor U16119 (N_16119,N_15905,N_15678);
nand U16120 (N_16120,N_15565,N_15788);
nor U16121 (N_16121,N_15704,N_15562);
and U16122 (N_16122,N_15685,N_15990);
nor U16123 (N_16123,N_15518,N_15867);
or U16124 (N_16124,N_15690,N_15674);
nand U16125 (N_16125,N_15639,N_15603);
and U16126 (N_16126,N_15911,N_15616);
and U16127 (N_16127,N_15925,N_15986);
and U16128 (N_16128,N_15708,N_15539);
nor U16129 (N_16129,N_15717,N_15581);
or U16130 (N_16130,N_15927,N_15727);
and U16131 (N_16131,N_15621,N_15933);
or U16132 (N_16132,N_15627,N_15878);
nor U16133 (N_16133,N_15997,N_15700);
or U16134 (N_16134,N_15513,N_15959);
nand U16135 (N_16135,N_15752,N_15841);
nand U16136 (N_16136,N_15558,N_15507);
and U16137 (N_16137,N_15563,N_15963);
nor U16138 (N_16138,N_15516,N_15871);
or U16139 (N_16139,N_15676,N_15837);
nand U16140 (N_16140,N_15910,N_15795);
nor U16141 (N_16141,N_15728,N_15736);
and U16142 (N_16142,N_15938,N_15835);
nand U16143 (N_16143,N_15693,N_15936);
nand U16144 (N_16144,N_15846,N_15800);
nor U16145 (N_16145,N_15681,N_15695);
nor U16146 (N_16146,N_15822,N_15744);
and U16147 (N_16147,N_15975,N_15943);
nand U16148 (N_16148,N_15597,N_15753);
xor U16149 (N_16149,N_15851,N_15944);
nand U16150 (N_16150,N_15971,N_15811);
and U16151 (N_16151,N_15907,N_15680);
or U16152 (N_16152,N_15823,N_15683);
nand U16153 (N_16153,N_15515,N_15571);
xnor U16154 (N_16154,N_15849,N_15995);
nor U16155 (N_16155,N_15988,N_15598);
xor U16156 (N_16156,N_15979,N_15773);
xnor U16157 (N_16157,N_15549,N_15534);
or U16158 (N_16158,N_15786,N_15729);
and U16159 (N_16159,N_15926,N_15934);
and U16160 (N_16160,N_15746,N_15863);
nor U16161 (N_16161,N_15635,N_15812);
or U16162 (N_16162,N_15921,N_15768);
nor U16163 (N_16163,N_15631,N_15909);
nand U16164 (N_16164,N_15740,N_15805);
and U16165 (N_16165,N_15575,N_15993);
nor U16166 (N_16166,N_15628,N_15808);
or U16167 (N_16167,N_15546,N_15935);
and U16168 (N_16168,N_15985,N_15814);
xnor U16169 (N_16169,N_15545,N_15734);
and U16170 (N_16170,N_15833,N_15923);
or U16171 (N_16171,N_15543,N_15894);
nor U16172 (N_16172,N_15723,N_15769);
nand U16173 (N_16173,N_15521,N_15928);
or U16174 (N_16174,N_15661,N_15544);
nor U16175 (N_16175,N_15702,N_15994);
or U16176 (N_16176,N_15557,N_15653);
and U16177 (N_16177,N_15903,N_15670);
and U16178 (N_16178,N_15525,N_15873);
nor U16179 (N_16179,N_15802,N_15858);
and U16180 (N_16180,N_15791,N_15524);
xor U16181 (N_16181,N_15813,N_15782);
xnor U16182 (N_16182,N_15742,N_15611);
nand U16183 (N_16183,N_15760,N_15646);
xor U16184 (N_16184,N_15642,N_15605);
and U16185 (N_16185,N_15908,N_15664);
or U16186 (N_16186,N_15815,N_15568);
nor U16187 (N_16187,N_15829,N_15987);
nor U16188 (N_16188,N_15792,N_15896);
or U16189 (N_16189,N_15889,N_15756);
xor U16190 (N_16190,N_15613,N_15657);
or U16191 (N_16191,N_15531,N_15677);
nand U16192 (N_16192,N_15850,N_15881);
nor U16193 (N_16193,N_15584,N_15946);
and U16194 (N_16194,N_15817,N_15892);
or U16195 (N_16195,N_15520,N_15739);
and U16196 (N_16196,N_15962,N_15591);
nand U16197 (N_16197,N_15902,N_15819);
xor U16198 (N_16198,N_15956,N_15667);
or U16199 (N_16199,N_15504,N_15586);
and U16200 (N_16200,N_15632,N_15601);
nand U16201 (N_16201,N_15540,N_15600);
nor U16202 (N_16202,N_15573,N_15825);
nor U16203 (N_16203,N_15733,N_15983);
nor U16204 (N_16204,N_15866,N_15924);
nor U16205 (N_16205,N_15654,N_15609);
xor U16206 (N_16206,N_15796,N_15901);
nand U16207 (N_16207,N_15640,N_15610);
nand U16208 (N_16208,N_15720,N_15659);
nor U16209 (N_16209,N_15860,N_15622);
nand U16210 (N_16210,N_15862,N_15980);
xnor U16211 (N_16211,N_15966,N_15735);
nor U16212 (N_16212,N_15807,N_15989);
nor U16213 (N_16213,N_15711,N_15906);
nor U16214 (N_16214,N_15751,N_15897);
or U16215 (N_16215,N_15960,N_15732);
nor U16216 (N_16216,N_15697,N_15572);
xnor U16217 (N_16217,N_15523,N_15529);
or U16218 (N_16218,N_15793,N_15550);
or U16219 (N_16219,N_15787,N_15750);
xor U16220 (N_16220,N_15877,N_15623);
and U16221 (N_16221,N_15818,N_15919);
nand U16222 (N_16222,N_15638,N_15517);
or U16223 (N_16223,N_15606,N_15932);
nand U16224 (N_16224,N_15857,N_15872);
or U16225 (N_16225,N_15650,N_15864);
nand U16226 (N_16226,N_15856,N_15519);
nor U16227 (N_16227,N_15893,N_15828);
and U16228 (N_16228,N_15976,N_15771);
or U16229 (N_16229,N_15977,N_15737);
nand U16230 (N_16230,N_15855,N_15533);
nor U16231 (N_16231,N_15508,N_15970);
or U16232 (N_16232,N_15633,N_15915);
and U16233 (N_16233,N_15541,N_15948);
or U16234 (N_16234,N_15887,N_15958);
and U16235 (N_16235,N_15673,N_15660);
or U16236 (N_16236,N_15940,N_15748);
nand U16237 (N_16237,N_15634,N_15982);
and U16238 (N_16238,N_15827,N_15974);
and U16239 (N_16239,N_15794,N_15698);
xnor U16240 (N_16240,N_15967,N_15799);
and U16241 (N_16241,N_15816,N_15798);
and U16242 (N_16242,N_15821,N_15594);
and U16243 (N_16243,N_15641,N_15691);
nand U16244 (N_16244,N_15527,N_15699);
and U16245 (N_16245,N_15630,N_15532);
nor U16246 (N_16246,N_15501,N_15547);
nand U16247 (N_16247,N_15712,N_15765);
and U16248 (N_16248,N_15770,N_15870);
nor U16249 (N_16249,N_15838,N_15503);
nand U16250 (N_16250,N_15881,N_15583);
xor U16251 (N_16251,N_15625,N_15993);
and U16252 (N_16252,N_15952,N_15909);
and U16253 (N_16253,N_15634,N_15939);
or U16254 (N_16254,N_15604,N_15574);
nor U16255 (N_16255,N_15811,N_15792);
xnor U16256 (N_16256,N_15997,N_15691);
nor U16257 (N_16257,N_15788,N_15889);
nand U16258 (N_16258,N_15919,N_15986);
nand U16259 (N_16259,N_15840,N_15882);
nor U16260 (N_16260,N_15520,N_15600);
or U16261 (N_16261,N_15512,N_15785);
or U16262 (N_16262,N_15701,N_15864);
nand U16263 (N_16263,N_15888,N_15611);
nor U16264 (N_16264,N_15541,N_15503);
nand U16265 (N_16265,N_15858,N_15748);
nand U16266 (N_16266,N_15653,N_15548);
and U16267 (N_16267,N_15755,N_15608);
and U16268 (N_16268,N_15869,N_15583);
xnor U16269 (N_16269,N_15636,N_15711);
and U16270 (N_16270,N_15510,N_15652);
nand U16271 (N_16271,N_15901,N_15511);
xor U16272 (N_16272,N_15551,N_15648);
xor U16273 (N_16273,N_15877,N_15756);
or U16274 (N_16274,N_15535,N_15680);
nor U16275 (N_16275,N_15500,N_15532);
nand U16276 (N_16276,N_15935,N_15635);
or U16277 (N_16277,N_15799,N_15559);
or U16278 (N_16278,N_15676,N_15715);
and U16279 (N_16279,N_15908,N_15543);
and U16280 (N_16280,N_15845,N_15552);
or U16281 (N_16281,N_15899,N_15657);
nand U16282 (N_16282,N_15867,N_15830);
nor U16283 (N_16283,N_15855,N_15993);
and U16284 (N_16284,N_15738,N_15574);
or U16285 (N_16285,N_15558,N_15736);
or U16286 (N_16286,N_15785,N_15756);
or U16287 (N_16287,N_15640,N_15906);
and U16288 (N_16288,N_15830,N_15939);
or U16289 (N_16289,N_15504,N_15934);
and U16290 (N_16290,N_15589,N_15551);
and U16291 (N_16291,N_15535,N_15677);
and U16292 (N_16292,N_15807,N_15937);
and U16293 (N_16293,N_15899,N_15984);
xnor U16294 (N_16294,N_15946,N_15860);
and U16295 (N_16295,N_15770,N_15906);
nor U16296 (N_16296,N_15752,N_15706);
or U16297 (N_16297,N_15587,N_15565);
and U16298 (N_16298,N_15989,N_15575);
and U16299 (N_16299,N_15536,N_15876);
nand U16300 (N_16300,N_15683,N_15850);
xnor U16301 (N_16301,N_15592,N_15887);
and U16302 (N_16302,N_15821,N_15866);
nor U16303 (N_16303,N_15995,N_15574);
xor U16304 (N_16304,N_15984,N_15565);
xnor U16305 (N_16305,N_15620,N_15920);
and U16306 (N_16306,N_15908,N_15643);
and U16307 (N_16307,N_15746,N_15798);
xnor U16308 (N_16308,N_15929,N_15576);
nor U16309 (N_16309,N_15645,N_15958);
and U16310 (N_16310,N_15812,N_15628);
nor U16311 (N_16311,N_15620,N_15878);
nand U16312 (N_16312,N_15514,N_15947);
or U16313 (N_16313,N_15706,N_15921);
xor U16314 (N_16314,N_15970,N_15993);
and U16315 (N_16315,N_15759,N_15810);
and U16316 (N_16316,N_15627,N_15750);
or U16317 (N_16317,N_15548,N_15655);
or U16318 (N_16318,N_15818,N_15547);
and U16319 (N_16319,N_15728,N_15899);
or U16320 (N_16320,N_15860,N_15701);
xor U16321 (N_16321,N_15962,N_15898);
and U16322 (N_16322,N_15910,N_15889);
nor U16323 (N_16323,N_15640,N_15871);
nor U16324 (N_16324,N_15701,N_15904);
nand U16325 (N_16325,N_15805,N_15964);
or U16326 (N_16326,N_15993,N_15850);
nor U16327 (N_16327,N_15766,N_15945);
and U16328 (N_16328,N_15520,N_15678);
nor U16329 (N_16329,N_15686,N_15651);
nor U16330 (N_16330,N_15678,N_15597);
or U16331 (N_16331,N_15985,N_15974);
nor U16332 (N_16332,N_15782,N_15735);
or U16333 (N_16333,N_15904,N_15627);
or U16334 (N_16334,N_15590,N_15902);
nor U16335 (N_16335,N_15641,N_15808);
nor U16336 (N_16336,N_15533,N_15986);
or U16337 (N_16337,N_15935,N_15748);
xnor U16338 (N_16338,N_15986,N_15659);
nor U16339 (N_16339,N_15997,N_15905);
and U16340 (N_16340,N_15651,N_15802);
xor U16341 (N_16341,N_15753,N_15586);
nand U16342 (N_16342,N_15789,N_15734);
and U16343 (N_16343,N_15617,N_15958);
or U16344 (N_16344,N_15696,N_15748);
xor U16345 (N_16345,N_15560,N_15837);
and U16346 (N_16346,N_15663,N_15613);
xor U16347 (N_16347,N_15552,N_15811);
or U16348 (N_16348,N_15502,N_15596);
xnor U16349 (N_16349,N_15868,N_15624);
xor U16350 (N_16350,N_15558,N_15602);
nand U16351 (N_16351,N_15638,N_15987);
xnor U16352 (N_16352,N_15689,N_15719);
or U16353 (N_16353,N_15802,N_15915);
and U16354 (N_16354,N_15709,N_15935);
or U16355 (N_16355,N_15858,N_15558);
xor U16356 (N_16356,N_15846,N_15753);
nand U16357 (N_16357,N_15593,N_15579);
or U16358 (N_16358,N_15700,N_15622);
nand U16359 (N_16359,N_15516,N_15913);
xnor U16360 (N_16360,N_15836,N_15608);
nand U16361 (N_16361,N_15684,N_15928);
nand U16362 (N_16362,N_15903,N_15809);
nor U16363 (N_16363,N_15546,N_15693);
nand U16364 (N_16364,N_15967,N_15609);
nor U16365 (N_16365,N_15950,N_15693);
xor U16366 (N_16366,N_15862,N_15847);
and U16367 (N_16367,N_15749,N_15665);
and U16368 (N_16368,N_15500,N_15527);
nor U16369 (N_16369,N_15934,N_15824);
nor U16370 (N_16370,N_15582,N_15571);
or U16371 (N_16371,N_15755,N_15763);
and U16372 (N_16372,N_15944,N_15707);
and U16373 (N_16373,N_15510,N_15638);
nand U16374 (N_16374,N_15853,N_15923);
or U16375 (N_16375,N_15520,N_15911);
nor U16376 (N_16376,N_15580,N_15594);
and U16377 (N_16377,N_15659,N_15908);
nor U16378 (N_16378,N_15959,N_15803);
or U16379 (N_16379,N_15860,N_15663);
or U16380 (N_16380,N_15560,N_15784);
and U16381 (N_16381,N_15920,N_15818);
or U16382 (N_16382,N_15825,N_15720);
nand U16383 (N_16383,N_15729,N_15860);
xor U16384 (N_16384,N_15627,N_15910);
or U16385 (N_16385,N_15949,N_15705);
nor U16386 (N_16386,N_15942,N_15659);
and U16387 (N_16387,N_15815,N_15894);
nor U16388 (N_16388,N_15948,N_15530);
xnor U16389 (N_16389,N_15856,N_15760);
xor U16390 (N_16390,N_15721,N_15787);
nand U16391 (N_16391,N_15672,N_15660);
nand U16392 (N_16392,N_15895,N_15862);
and U16393 (N_16393,N_15590,N_15838);
or U16394 (N_16394,N_15818,N_15878);
nor U16395 (N_16395,N_15934,N_15564);
and U16396 (N_16396,N_15566,N_15517);
xor U16397 (N_16397,N_15585,N_15635);
nand U16398 (N_16398,N_15772,N_15808);
and U16399 (N_16399,N_15993,N_15965);
nand U16400 (N_16400,N_15838,N_15622);
or U16401 (N_16401,N_15537,N_15942);
nand U16402 (N_16402,N_15856,N_15776);
nor U16403 (N_16403,N_15713,N_15864);
xor U16404 (N_16404,N_15627,N_15531);
nor U16405 (N_16405,N_15539,N_15835);
xor U16406 (N_16406,N_15717,N_15751);
nor U16407 (N_16407,N_15924,N_15625);
or U16408 (N_16408,N_15928,N_15784);
or U16409 (N_16409,N_15988,N_15835);
xor U16410 (N_16410,N_15669,N_15975);
or U16411 (N_16411,N_15856,N_15653);
xnor U16412 (N_16412,N_15679,N_15950);
and U16413 (N_16413,N_15600,N_15623);
and U16414 (N_16414,N_15854,N_15512);
nand U16415 (N_16415,N_15649,N_15746);
or U16416 (N_16416,N_15636,N_15751);
xor U16417 (N_16417,N_15667,N_15525);
nand U16418 (N_16418,N_15613,N_15822);
or U16419 (N_16419,N_15683,N_15913);
or U16420 (N_16420,N_15502,N_15626);
nand U16421 (N_16421,N_15918,N_15812);
nand U16422 (N_16422,N_15995,N_15873);
and U16423 (N_16423,N_15988,N_15875);
xor U16424 (N_16424,N_15723,N_15896);
xor U16425 (N_16425,N_15917,N_15557);
nand U16426 (N_16426,N_15730,N_15952);
xnor U16427 (N_16427,N_15598,N_15628);
xor U16428 (N_16428,N_15911,N_15906);
and U16429 (N_16429,N_15614,N_15504);
or U16430 (N_16430,N_15783,N_15607);
xor U16431 (N_16431,N_15580,N_15726);
nor U16432 (N_16432,N_15819,N_15942);
xor U16433 (N_16433,N_15848,N_15653);
or U16434 (N_16434,N_15937,N_15675);
xnor U16435 (N_16435,N_15852,N_15714);
and U16436 (N_16436,N_15510,N_15759);
xnor U16437 (N_16437,N_15818,N_15967);
xnor U16438 (N_16438,N_15614,N_15653);
or U16439 (N_16439,N_15887,N_15627);
and U16440 (N_16440,N_15635,N_15656);
nand U16441 (N_16441,N_15926,N_15559);
and U16442 (N_16442,N_15725,N_15938);
or U16443 (N_16443,N_15543,N_15619);
nand U16444 (N_16444,N_15707,N_15990);
xnor U16445 (N_16445,N_15711,N_15684);
or U16446 (N_16446,N_15841,N_15543);
nand U16447 (N_16447,N_15593,N_15825);
and U16448 (N_16448,N_15861,N_15696);
xor U16449 (N_16449,N_15773,N_15516);
nand U16450 (N_16450,N_15707,N_15681);
xor U16451 (N_16451,N_15947,N_15879);
xor U16452 (N_16452,N_15849,N_15601);
nand U16453 (N_16453,N_15848,N_15870);
or U16454 (N_16454,N_15739,N_15551);
and U16455 (N_16455,N_15687,N_15848);
xnor U16456 (N_16456,N_15959,N_15724);
or U16457 (N_16457,N_15833,N_15625);
nand U16458 (N_16458,N_15572,N_15633);
nand U16459 (N_16459,N_15881,N_15898);
xnor U16460 (N_16460,N_15931,N_15798);
nor U16461 (N_16461,N_15593,N_15962);
or U16462 (N_16462,N_15721,N_15890);
and U16463 (N_16463,N_15770,N_15659);
nor U16464 (N_16464,N_15892,N_15681);
xor U16465 (N_16465,N_15658,N_15610);
and U16466 (N_16466,N_15652,N_15532);
nand U16467 (N_16467,N_15861,N_15967);
xnor U16468 (N_16468,N_15890,N_15853);
and U16469 (N_16469,N_15869,N_15640);
nor U16470 (N_16470,N_15600,N_15777);
xnor U16471 (N_16471,N_15875,N_15780);
xnor U16472 (N_16472,N_15723,N_15502);
nor U16473 (N_16473,N_15509,N_15811);
xnor U16474 (N_16474,N_15616,N_15896);
or U16475 (N_16475,N_15928,N_15956);
nand U16476 (N_16476,N_15602,N_15844);
nor U16477 (N_16477,N_15962,N_15740);
and U16478 (N_16478,N_15557,N_15676);
xor U16479 (N_16479,N_15719,N_15618);
nor U16480 (N_16480,N_15811,N_15675);
xor U16481 (N_16481,N_15834,N_15975);
xnor U16482 (N_16482,N_15854,N_15887);
nand U16483 (N_16483,N_15784,N_15717);
xor U16484 (N_16484,N_15540,N_15616);
and U16485 (N_16485,N_15804,N_15545);
xnor U16486 (N_16486,N_15584,N_15698);
xnor U16487 (N_16487,N_15579,N_15685);
or U16488 (N_16488,N_15963,N_15869);
nor U16489 (N_16489,N_15776,N_15965);
nor U16490 (N_16490,N_15823,N_15897);
xnor U16491 (N_16491,N_15630,N_15958);
nand U16492 (N_16492,N_15851,N_15961);
nor U16493 (N_16493,N_15894,N_15737);
or U16494 (N_16494,N_15778,N_15993);
or U16495 (N_16495,N_15799,N_15669);
nand U16496 (N_16496,N_15729,N_15904);
and U16497 (N_16497,N_15521,N_15706);
nand U16498 (N_16498,N_15579,N_15984);
or U16499 (N_16499,N_15689,N_15908);
and U16500 (N_16500,N_16013,N_16137);
and U16501 (N_16501,N_16381,N_16136);
xor U16502 (N_16502,N_16435,N_16220);
nand U16503 (N_16503,N_16192,N_16116);
xnor U16504 (N_16504,N_16465,N_16335);
nor U16505 (N_16505,N_16436,N_16401);
xnor U16506 (N_16506,N_16411,N_16457);
or U16507 (N_16507,N_16298,N_16160);
nand U16508 (N_16508,N_16458,N_16405);
xor U16509 (N_16509,N_16170,N_16200);
and U16510 (N_16510,N_16259,N_16452);
and U16511 (N_16511,N_16224,N_16043);
xnor U16512 (N_16512,N_16319,N_16470);
nand U16513 (N_16513,N_16450,N_16423);
nand U16514 (N_16514,N_16364,N_16242);
or U16515 (N_16515,N_16366,N_16288);
nand U16516 (N_16516,N_16246,N_16026);
or U16517 (N_16517,N_16362,N_16353);
xnor U16518 (N_16518,N_16077,N_16199);
nor U16519 (N_16519,N_16069,N_16083);
and U16520 (N_16520,N_16023,N_16201);
or U16521 (N_16521,N_16451,N_16312);
xor U16522 (N_16522,N_16165,N_16301);
xnor U16523 (N_16523,N_16219,N_16463);
or U16524 (N_16524,N_16359,N_16247);
nor U16525 (N_16525,N_16037,N_16406);
or U16526 (N_16526,N_16210,N_16253);
xnor U16527 (N_16527,N_16391,N_16328);
xor U16528 (N_16528,N_16268,N_16261);
and U16529 (N_16529,N_16025,N_16325);
xnor U16530 (N_16530,N_16140,N_16213);
xor U16531 (N_16531,N_16475,N_16095);
xnor U16532 (N_16532,N_16074,N_16087);
and U16533 (N_16533,N_16464,N_16340);
nand U16534 (N_16534,N_16015,N_16299);
xnor U16535 (N_16535,N_16115,N_16058);
or U16536 (N_16536,N_16202,N_16208);
nand U16537 (N_16537,N_16339,N_16008);
xnor U16538 (N_16538,N_16035,N_16172);
nor U16539 (N_16539,N_16356,N_16499);
or U16540 (N_16540,N_16343,N_16168);
nand U16541 (N_16541,N_16047,N_16085);
and U16542 (N_16542,N_16098,N_16324);
or U16543 (N_16543,N_16379,N_16412);
and U16544 (N_16544,N_16046,N_16417);
or U16545 (N_16545,N_16012,N_16321);
nand U16546 (N_16546,N_16029,N_16307);
nand U16547 (N_16547,N_16142,N_16016);
nand U16548 (N_16548,N_16327,N_16304);
or U16549 (N_16549,N_16461,N_16432);
and U16550 (N_16550,N_16385,N_16131);
nor U16551 (N_16551,N_16326,N_16150);
xnor U16552 (N_16552,N_16103,N_16292);
nand U16553 (N_16553,N_16119,N_16146);
or U16554 (N_16554,N_16196,N_16471);
nand U16555 (N_16555,N_16264,N_16084);
or U16556 (N_16556,N_16444,N_16446);
xor U16557 (N_16557,N_16212,N_16110);
and U16558 (N_16558,N_16291,N_16493);
and U16559 (N_16559,N_16260,N_16222);
nor U16560 (N_16560,N_16061,N_16177);
xnor U16561 (N_16561,N_16473,N_16185);
and U16562 (N_16562,N_16141,N_16266);
or U16563 (N_16563,N_16236,N_16104);
xnor U16564 (N_16564,N_16494,N_16333);
nor U16565 (N_16565,N_16322,N_16138);
xnor U16566 (N_16566,N_16289,N_16243);
or U16567 (N_16567,N_16389,N_16062);
and U16568 (N_16568,N_16102,N_16252);
xnor U16569 (N_16569,N_16409,N_16360);
nor U16570 (N_16570,N_16193,N_16229);
or U16571 (N_16571,N_16075,N_16109);
nor U16572 (N_16572,N_16216,N_16375);
or U16573 (N_16573,N_16245,N_16332);
or U16574 (N_16574,N_16238,N_16280);
nand U16575 (N_16575,N_16021,N_16189);
or U16576 (N_16576,N_16030,N_16349);
nor U16577 (N_16577,N_16005,N_16311);
xor U16578 (N_16578,N_16420,N_16014);
or U16579 (N_16579,N_16313,N_16392);
nand U16580 (N_16580,N_16300,N_16348);
nor U16581 (N_16581,N_16318,N_16113);
xor U16582 (N_16582,N_16002,N_16370);
nand U16583 (N_16583,N_16302,N_16265);
nand U16584 (N_16584,N_16225,N_16135);
or U16585 (N_16585,N_16000,N_16134);
and U16586 (N_16586,N_16357,N_16020);
nand U16587 (N_16587,N_16305,N_16296);
nor U16588 (N_16588,N_16351,N_16433);
or U16589 (N_16589,N_16235,N_16211);
xor U16590 (N_16590,N_16445,N_16231);
xnor U16591 (N_16591,N_16408,N_16334);
nand U16592 (N_16592,N_16485,N_16459);
or U16593 (N_16593,N_16257,N_16094);
xnor U16594 (N_16594,N_16010,N_16162);
nor U16595 (N_16595,N_16440,N_16341);
and U16596 (N_16596,N_16228,N_16278);
nand U16597 (N_16597,N_16143,N_16218);
or U16598 (N_16598,N_16100,N_16107);
nand U16599 (N_16599,N_16466,N_16164);
nand U16600 (N_16600,N_16276,N_16378);
nand U16601 (N_16601,N_16114,N_16315);
xor U16602 (N_16602,N_16358,N_16082);
or U16603 (N_16603,N_16441,N_16028);
or U16604 (N_16604,N_16101,N_16293);
and U16605 (N_16605,N_16443,N_16111);
nor U16606 (N_16606,N_16376,N_16407);
xor U16607 (N_16607,N_16284,N_16112);
nor U16608 (N_16608,N_16181,N_16352);
xnor U16609 (N_16609,N_16024,N_16019);
nor U16610 (N_16610,N_16064,N_16174);
xnor U16611 (N_16611,N_16422,N_16044);
and U16612 (N_16612,N_16428,N_16286);
and U16613 (N_16613,N_16039,N_16051);
xor U16614 (N_16614,N_16027,N_16067);
or U16615 (N_16615,N_16171,N_16402);
xnor U16616 (N_16616,N_16057,N_16003);
nand U16617 (N_16617,N_16032,N_16240);
nand U16618 (N_16618,N_16303,N_16486);
xnor U16619 (N_16619,N_16400,N_16195);
nor U16620 (N_16620,N_16159,N_16294);
xor U16621 (N_16621,N_16049,N_16209);
or U16622 (N_16622,N_16413,N_16439);
xor U16623 (N_16623,N_16017,N_16447);
or U16624 (N_16624,N_16380,N_16271);
xnor U16625 (N_16625,N_16279,N_16410);
nor U16626 (N_16626,N_16425,N_16456);
and U16627 (N_16627,N_16022,N_16495);
and U16628 (N_16628,N_16151,N_16490);
nor U16629 (N_16629,N_16125,N_16053);
or U16630 (N_16630,N_16317,N_16217);
nand U16631 (N_16631,N_16093,N_16108);
xnor U16632 (N_16632,N_16206,N_16234);
and U16633 (N_16633,N_16283,N_16155);
nand U16634 (N_16634,N_16052,N_16316);
xnor U16635 (N_16635,N_16045,N_16190);
nand U16636 (N_16636,N_16144,N_16361);
or U16637 (N_16637,N_16281,N_16059);
and U16638 (N_16638,N_16184,N_16398);
and U16639 (N_16639,N_16429,N_16065);
or U16640 (N_16640,N_16418,N_16282);
and U16641 (N_16641,N_16481,N_16421);
and U16642 (N_16642,N_16258,N_16214);
nor U16643 (N_16643,N_16187,N_16484);
nand U16644 (N_16644,N_16118,N_16106);
and U16645 (N_16645,N_16197,N_16419);
or U16646 (N_16646,N_16078,N_16180);
xnor U16647 (N_16647,N_16384,N_16152);
or U16648 (N_16648,N_16018,N_16403);
nor U16649 (N_16649,N_16011,N_16467);
nor U16650 (N_16650,N_16272,N_16230);
nor U16651 (N_16651,N_16176,N_16431);
xnor U16652 (N_16652,N_16454,N_16215);
or U16653 (N_16653,N_16329,N_16068);
nor U16654 (N_16654,N_16350,N_16223);
nand U16655 (N_16655,N_16416,N_16123);
xor U16656 (N_16656,N_16121,N_16394);
or U16657 (N_16657,N_16241,N_16092);
nor U16658 (N_16658,N_16161,N_16221);
nor U16659 (N_16659,N_16158,N_16255);
and U16660 (N_16660,N_16397,N_16060);
nand U16661 (N_16661,N_16396,N_16479);
nor U16662 (N_16662,N_16331,N_16076);
xor U16663 (N_16663,N_16133,N_16497);
nand U16664 (N_16664,N_16460,N_16194);
and U16665 (N_16665,N_16117,N_16033);
and U16666 (N_16666,N_16472,N_16041);
and U16667 (N_16667,N_16330,N_16167);
xnor U16668 (N_16668,N_16346,N_16145);
and U16669 (N_16669,N_16034,N_16239);
nor U16670 (N_16670,N_16338,N_16274);
nand U16671 (N_16671,N_16128,N_16480);
and U16672 (N_16672,N_16437,N_16369);
and U16673 (N_16673,N_16081,N_16275);
or U16674 (N_16674,N_16295,N_16476);
nand U16675 (N_16675,N_16426,N_16404);
nor U16676 (N_16676,N_16250,N_16469);
and U16677 (N_16677,N_16427,N_16249);
nor U16678 (N_16678,N_16182,N_16129);
nand U16679 (N_16679,N_16132,N_16173);
nand U16680 (N_16680,N_16154,N_16448);
nand U16681 (N_16681,N_16166,N_16001);
or U16682 (N_16682,N_16383,N_16483);
nor U16683 (N_16683,N_16310,N_16468);
nor U16684 (N_16684,N_16347,N_16097);
nor U16685 (N_16685,N_16153,N_16478);
nor U16686 (N_16686,N_16090,N_16449);
nor U16687 (N_16687,N_16474,N_16323);
nand U16688 (N_16688,N_16367,N_16424);
xnor U16689 (N_16689,N_16256,N_16462);
and U16690 (N_16690,N_16254,N_16186);
or U16691 (N_16691,N_16105,N_16377);
nor U16692 (N_16692,N_16147,N_16120);
or U16693 (N_16693,N_16482,N_16089);
or U16694 (N_16694,N_16270,N_16226);
or U16695 (N_16695,N_16086,N_16169);
xor U16696 (N_16696,N_16127,N_16442);
xor U16697 (N_16697,N_16354,N_16487);
or U16698 (N_16698,N_16066,N_16390);
and U16699 (N_16699,N_16232,N_16007);
nor U16700 (N_16700,N_16496,N_16345);
xor U16701 (N_16701,N_16368,N_16244);
nand U16702 (N_16702,N_16096,N_16175);
nor U16703 (N_16703,N_16056,N_16363);
nor U16704 (N_16704,N_16099,N_16183);
xnor U16705 (N_16705,N_16262,N_16477);
or U16706 (N_16706,N_16157,N_16124);
nand U16707 (N_16707,N_16205,N_16438);
xnor U16708 (N_16708,N_16399,N_16309);
or U16709 (N_16709,N_16163,N_16371);
or U16710 (N_16710,N_16009,N_16285);
xnor U16711 (N_16711,N_16387,N_16048);
nand U16712 (N_16712,N_16372,N_16453);
xnor U16713 (N_16713,N_16308,N_16336);
or U16714 (N_16714,N_16126,N_16297);
or U16715 (N_16715,N_16373,N_16073);
nand U16716 (N_16716,N_16038,N_16355);
xor U16717 (N_16717,N_16203,N_16050);
xnor U16718 (N_16718,N_16227,N_16042);
xor U16719 (N_16719,N_16344,N_16178);
and U16720 (N_16720,N_16040,N_16365);
and U16721 (N_16721,N_16139,N_16036);
or U16722 (N_16722,N_16263,N_16148);
xor U16723 (N_16723,N_16149,N_16251);
nand U16724 (N_16724,N_16415,N_16337);
or U16725 (N_16725,N_16492,N_16430);
xnor U16726 (N_16726,N_16179,N_16054);
and U16727 (N_16727,N_16388,N_16072);
or U16728 (N_16728,N_16374,N_16489);
nor U16729 (N_16729,N_16314,N_16055);
nor U16730 (N_16730,N_16004,N_16063);
or U16731 (N_16731,N_16277,N_16191);
or U16732 (N_16732,N_16267,N_16006);
and U16733 (N_16733,N_16070,N_16342);
xnor U16734 (N_16734,N_16269,N_16130);
and U16735 (N_16735,N_16395,N_16290);
and U16736 (N_16736,N_16491,N_16088);
nand U16737 (N_16737,N_16204,N_16188);
or U16738 (N_16738,N_16207,N_16455);
or U16739 (N_16739,N_16306,N_16287);
nand U16740 (N_16740,N_16248,N_16273);
xnor U16741 (N_16741,N_16031,N_16393);
nor U16742 (N_16742,N_16237,N_16198);
nand U16743 (N_16743,N_16156,N_16071);
nand U16744 (N_16744,N_16233,N_16386);
or U16745 (N_16745,N_16080,N_16498);
nand U16746 (N_16746,N_16079,N_16091);
or U16747 (N_16747,N_16382,N_16488);
or U16748 (N_16748,N_16414,N_16122);
xor U16749 (N_16749,N_16320,N_16434);
or U16750 (N_16750,N_16311,N_16455);
and U16751 (N_16751,N_16144,N_16262);
and U16752 (N_16752,N_16376,N_16104);
xnor U16753 (N_16753,N_16116,N_16224);
nor U16754 (N_16754,N_16358,N_16433);
nand U16755 (N_16755,N_16055,N_16385);
nand U16756 (N_16756,N_16409,N_16167);
nor U16757 (N_16757,N_16070,N_16389);
xnor U16758 (N_16758,N_16064,N_16225);
or U16759 (N_16759,N_16451,N_16064);
nor U16760 (N_16760,N_16287,N_16107);
nand U16761 (N_16761,N_16064,N_16324);
or U16762 (N_16762,N_16166,N_16173);
and U16763 (N_16763,N_16386,N_16390);
xnor U16764 (N_16764,N_16257,N_16303);
nor U16765 (N_16765,N_16311,N_16007);
and U16766 (N_16766,N_16387,N_16194);
nor U16767 (N_16767,N_16497,N_16410);
and U16768 (N_16768,N_16319,N_16127);
or U16769 (N_16769,N_16336,N_16366);
nand U16770 (N_16770,N_16128,N_16036);
xor U16771 (N_16771,N_16008,N_16312);
or U16772 (N_16772,N_16048,N_16378);
nand U16773 (N_16773,N_16041,N_16034);
and U16774 (N_16774,N_16164,N_16373);
and U16775 (N_16775,N_16409,N_16159);
nor U16776 (N_16776,N_16194,N_16394);
or U16777 (N_16777,N_16328,N_16127);
or U16778 (N_16778,N_16022,N_16426);
xor U16779 (N_16779,N_16254,N_16470);
and U16780 (N_16780,N_16233,N_16356);
or U16781 (N_16781,N_16031,N_16456);
or U16782 (N_16782,N_16327,N_16421);
and U16783 (N_16783,N_16217,N_16319);
nor U16784 (N_16784,N_16377,N_16450);
and U16785 (N_16785,N_16227,N_16340);
nor U16786 (N_16786,N_16466,N_16135);
or U16787 (N_16787,N_16363,N_16220);
or U16788 (N_16788,N_16380,N_16075);
nand U16789 (N_16789,N_16133,N_16143);
and U16790 (N_16790,N_16209,N_16018);
or U16791 (N_16791,N_16277,N_16207);
nand U16792 (N_16792,N_16426,N_16493);
nor U16793 (N_16793,N_16015,N_16474);
nor U16794 (N_16794,N_16029,N_16222);
xnor U16795 (N_16795,N_16353,N_16366);
nor U16796 (N_16796,N_16197,N_16129);
xnor U16797 (N_16797,N_16352,N_16300);
xor U16798 (N_16798,N_16031,N_16200);
nor U16799 (N_16799,N_16073,N_16259);
or U16800 (N_16800,N_16070,N_16487);
xnor U16801 (N_16801,N_16357,N_16350);
nor U16802 (N_16802,N_16153,N_16241);
and U16803 (N_16803,N_16259,N_16359);
nand U16804 (N_16804,N_16403,N_16233);
xor U16805 (N_16805,N_16225,N_16161);
nor U16806 (N_16806,N_16270,N_16199);
nor U16807 (N_16807,N_16310,N_16107);
xor U16808 (N_16808,N_16165,N_16095);
xnor U16809 (N_16809,N_16450,N_16030);
or U16810 (N_16810,N_16167,N_16194);
xor U16811 (N_16811,N_16241,N_16057);
or U16812 (N_16812,N_16489,N_16026);
or U16813 (N_16813,N_16121,N_16271);
xor U16814 (N_16814,N_16426,N_16125);
nor U16815 (N_16815,N_16480,N_16335);
nor U16816 (N_16816,N_16431,N_16345);
or U16817 (N_16817,N_16087,N_16112);
or U16818 (N_16818,N_16034,N_16119);
nand U16819 (N_16819,N_16368,N_16343);
nand U16820 (N_16820,N_16317,N_16273);
xnor U16821 (N_16821,N_16406,N_16151);
nand U16822 (N_16822,N_16264,N_16255);
xor U16823 (N_16823,N_16010,N_16073);
nand U16824 (N_16824,N_16253,N_16376);
or U16825 (N_16825,N_16119,N_16408);
or U16826 (N_16826,N_16203,N_16459);
or U16827 (N_16827,N_16079,N_16228);
nor U16828 (N_16828,N_16146,N_16406);
nor U16829 (N_16829,N_16436,N_16097);
or U16830 (N_16830,N_16487,N_16452);
and U16831 (N_16831,N_16291,N_16301);
nand U16832 (N_16832,N_16344,N_16055);
and U16833 (N_16833,N_16378,N_16175);
and U16834 (N_16834,N_16491,N_16272);
and U16835 (N_16835,N_16186,N_16388);
nor U16836 (N_16836,N_16252,N_16417);
xnor U16837 (N_16837,N_16038,N_16139);
or U16838 (N_16838,N_16294,N_16289);
nor U16839 (N_16839,N_16234,N_16177);
and U16840 (N_16840,N_16376,N_16348);
xor U16841 (N_16841,N_16363,N_16235);
nor U16842 (N_16842,N_16033,N_16384);
nor U16843 (N_16843,N_16166,N_16287);
and U16844 (N_16844,N_16474,N_16426);
nand U16845 (N_16845,N_16049,N_16456);
and U16846 (N_16846,N_16323,N_16430);
and U16847 (N_16847,N_16298,N_16462);
or U16848 (N_16848,N_16320,N_16390);
and U16849 (N_16849,N_16151,N_16265);
nor U16850 (N_16850,N_16395,N_16089);
and U16851 (N_16851,N_16285,N_16494);
or U16852 (N_16852,N_16466,N_16429);
nor U16853 (N_16853,N_16194,N_16039);
nor U16854 (N_16854,N_16357,N_16424);
xnor U16855 (N_16855,N_16444,N_16096);
and U16856 (N_16856,N_16305,N_16239);
nor U16857 (N_16857,N_16113,N_16172);
and U16858 (N_16858,N_16441,N_16354);
and U16859 (N_16859,N_16229,N_16296);
or U16860 (N_16860,N_16187,N_16352);
nor U16861 (N_16861,N_16332,N_16155);
nor U16862 (N_16862,N_16463,N_16310);
nor U16863 (N_16863,N_16464,N_16395);
nor U16864 (N_16864,N_16452,N_16149);
nor U16865 (N_16865,N_16261,N_16355);
xor U16866 (N_16866,N_16308,N_16384);
nand U16867 (N_16867,N_16244,N_16128);
and U16868 (N_16868,N_16071,N_16293);
nor U16869 (N_16869,N_16184,N_16207);
xor U16870 (N_16870,N_16251,N_16371);
xnor U16871 (N_16871,N_16335,N_16372);
nand U16872 (N_16872,N_16156,N_16232);
nand U16873 (N_16873,N_16299,N_16428);
nand U16874 (N_16874,N_16384,N_16402);
or U16875 (N_16875,N_16056,N_16173);
xor U16876 (N_16876,N_16182,N_16251);
nand U16877 (N_16877,N_16363,N_16038);
nor U16878 (N_16878,N_16020,N_16390);
and U16879 (N_16879,N_16183,N_16217);
nand U16880 (N_16880,N_16309,N_16408);
xnor U16881 (N_16881,N_16192,N_16152);
nand U16882 (N_16882,N_16039,N_16408);
and U16883 (N_16883,N_16003,N_16384);
or U16884 (N_16884,N_16327,N_16466);
xnor U16885 (N_16885,N_16347,N_16330);
nand U16886 (N_16886,N_16085,N_16204);
xor U16887 (N_16887,N_16320,N_16450);
xor U16888 (N_16888,N_16199,N_16249);
and U16889 (N_16889,N_16025,N_16485);
nor U16890 (N_16890,N_16233,N_16254);
nor U16891 (N_16891,N_16324,N_16489);
or U16892 (N_16892,N_16450,N_16184);
or U16893 (N_16893,N_16102,N_16390);
or U16894 (N_16894,N_16124,N_16402);
nor U16895 (N_16895,N_16114,N_16142);
nand U16896 (N_16896,N_16059,N_16426);
and U16897 (N_16897,N_16074,N_16027);
or U16898 (N_16898,N_16290,N_16115);
and U16899 (N_16899,N_16459,N_16314);
or U16900 (N_16900,N_16373,N_16480);
or U16901 (N_16901,N_16274,N_16031);
and U16902 (N_16902,N_16388,N_16333);
or U16903 (N_16903,N_16444,N_16276);
or U16904 (N_16904,N_16243,N_16385);
nor U16905 (N_16905,N_16090,N_16187);
nor U16906 (N_16906,N_16291,N_16368);
nand U16907 (N_16907,N_16312,N_16112);
xnor U16908 (N_16908,N_16072,N_16363);
nor U16909 (N_16909,N_16037,N_16284);
nor U16910 (N_16910,N_16438,N_16096);
or U16911 (N_16911,N_16273,N_16265);
nand U16912 (N_16912,N_16223,N_16111);
or U16913 (N_16913,N_16303,N_16110);
xor U16914 (N_16914,N_16287,N_16311);
or U16915 (N_16915,N_16327,N_16019);
or U16916 (N_16916,N_16283,N_16431);
nor U16917 (N_16917,N_16448,N_16073);
and U16918 (N_16918,N_16351,N_16446);
xnor U16919 (N_16919,N_16217,N_16134);
nor U16920 (N_16920,N_16268,N_16057);
nand U16921 (N_16921,N_16332,N_16055);
nor U16922 (N_16922,N_16014,N_16210);
xnor U16923 (N_16923,N_16211,N_16167);
and U16924 (N_16924,N_16108,N_16002);
xor U16925 (N_16925,N_16044,N_16276);
nand U16926 (N_16926,N_16413,N_16328);
xor U16927 (N_16927,N_16146,N_16390);
xor U16928 (N_16928,N_16344,N_16112);
or U16929 (N_16929,N_16328,N_16064);
xor U16930 (N_16930,N_16441,N_16333);
nand U16931 (N_16931,N_16191,N_16252);
nor U16932 (N_16932,N_16212,N_16224);
nor U16933 (N_16933,N_16495,N_16362);
and U16934 (N_16934,N_16289,N_16339);
or U16935 (N_16935,N_16008,N_16278);
and U16936 (N_16936,N_16451,N_16162);
and U16937 (N_16937,N_16115,N_16096);
or U16938 (N_16938,N_16036,N_16190);
and U16939 (N_16939,N_16473,N_16372);
nor U16940 (N_16940,N_16334,N_16400);
and U16941 (N_16941,N_16464,N_16030);
nand U16942 (N_16942,N_16403,N_16357);
and U16943 (N_16943,N_16497,N_16335);
nand U16944 (N_16944,N_16372,N_16443);
xor U16945 (N_16945,N_16130,N_16381);
or U16946 (N_16946,N_16135,N_16232);
and U16947 (N_16947,N_16448,N_16338);
nand U16948 (N_16948,N_16218,N_16123);
xor U16949 (N_16949,N_16440,N_16382);
and U16950 (N_16950,N_16271,N_16310);
xnor U16951 (N_16951,N_16289,N_16114);
nor U16952 (N_16952,N_16243,N_16150);
or U16953 (N_16953,N_16479,N_16401);
nor U16954 (N_16954,N_16170,N_16160);
nor U16955 (N_16955,N_16211,N_16128);
nand U16956 (N_16956,N_16239,N_16359);
nor U16957 (N_16957,N_16390,N_16117);
and U16958 (N_16958,N_16424,N_16229);
xor U16959 (N_16959,N_16339,N_16314);
xnor U16960 (N_16960,N_16001,N_16185);
and U16961 (N_16961,N_16448,N_16104);
xnor U16962 (N_16962,N_16273,N_16151);
and U16963 (N_16963,N_16175,N_16009);
and U16964 (N_16964,N_16285,N_16183);
or U16965 (N_16965,N_16489,N_16184);
nand U16966 (N_16966,N_16378,N_16009);
or U16967 (N_16967,N_16178,N_16006);
xor U16968 (N_16968,N_16167,N_16075);
and U16969 (N_16969,N_16297,N_16405);
nand U16970 (N_16970,N_16323,N_16259);
or U16971 (N_16971,N_16285,N_16140);
or U16972 (N_16972,N_16438,N_16118);
nand U16973 (N_16973,N_16290,N_16074);
and U16974 (N_16974,N_16135,N_16370);
xor U16975 (N_16975,N_16257,N_16231);
nor U16976 (N_16976,N_16180,N_16198);
nand U16977 (N_16977,N_16484,N_16252);
or U16978 (N_16978,N_16442,N_16496);
nor U16979 (N_16979,N_16339,N_16349);
or U16980 (N_16980,N_16267,N_16090);
nor U16981 (N_16981,N_16308,N_16443);
nor U16982 (N_16982,N_16304,N_16451);
xnor U16983 (N_16983,N_16229,N_16045);
nor U16984 (N_16984,N_16005,N_16474);
xor U16985 (N_16985,N_16038,N_16193);
xor U16986 (N_16986,N_16003,N_16496);
and U16987 (N_16987,N_16017,N_16133);
nand U16988 (N_16988,N_16213,N_16160);
nand U16989 (N_16989,N_16299,N_16159);
nand U16990 (N_16990,N_16448,N_16429);
and U16991 (N_16991,N_16230,N_16068);
nand U16992 (N_16992,N_16417,N_16228);
xnor U16993 (N_16993,N_16112,N_16232);
and U16994 (N_16994,N_16496,N_16402);
and U16995 (N_16995,N_16222,N_16078);
nor U16996 (N_16996,N_16432,N_16345);
or U16997 (N_16997,N_16257,N_16193);
nand U16998 (N_16998,N_16052,N_16420);
nor U16999 (N_16999,N_16007,N_16238);
xnor U17000 (N_17000,N_16962,N_16522);
xor U17001 (N_17001,N_16756,N_16630);
nor U17002 (N_17002,N_16923,N_16767);
or U17003 (N_17003,N_16573,N_16623);
nand U17004 (N_17004,N_16832,N_16880);
nand U17005 (N_17005,N_16904,N_16699);
nor U17006 (N_17006,N_16902,N_16976);
and U17007 (N_17007,N_16993,N_16857);
and U17008 (N_17008,N_16824,N_16546);
nor U17009 (N_17009,N_16787,N_16636);
or U17010 (N_17010,N_16728,N_16854);
nand U17011 (N_17011,N_16607,N_16778);
xnor U17012 (N_17012,N_16761,N_16618);
or U17013 (N_17013,N_16763,N_16501);
xor U17014 (N_17014,N_16863,N_16974);
nand U17015 (N_17015,N_16706,N_16885);
nand U17016 (N_17016,N_16870,N_16614);
xnor U17017 (N_17017,N_16658,N_16650);
and U17018 (N_17018,N_16820,N_16861);
nand U17019 (N_17019,N_16814,N_16887);
nor U17020 (N_17020,N_16825,N_16682);
and U17021 (N_17021,N_16506,N_16505);
nor U17022 (N_17022,N_16987,N_16813);
or U17023 (N_17023,N_16540,N_16687);
nand U17024 (N_17024,N_16674,N_16587);
nand U17025 (N_17025,N_16991,N_16586);
and U17026 (N_17026,N_16806,N_16879);
or U17027 (N_17027,N_16542,N_16717);
nand U17028 (N_17028,N_16627,N_16664);
or U17029 (N_17029,N_16519,N_16979);
xor U17030 (N_17030,N_16708,N_16898);
nor U17031 (N_17031,N_16510,N_16855);
and U17032 (N_17032,N_16570,N_16713);
and U17033 (N_17033,N_16560,N_16942);
nor U17034 (N_17034,N_16828,N_16966);
xor U17035 (N_17035,N_16792,N_16817);
xnor U17036 (N_17036,N_16638,N_16982);
or U17037 (N_17037,N_16804,N_16836);
nor U17038 (N_17038,N_16666,N_16949);
nor U17039 (N_17039,N_16507,N_16574);
and U17040 (N_17040,N_16801,N_16597);
or U17041 (N_17041,N_16919,N_16697);
and U17042 (N_17042,N_16973,N_16661);
and U17043 (N_17043,N_16803,N_16534);
xnor U17044 (N_17044,N_16943,N_16707);
and U17045 (N_17045,N_16997,N_16797);
nand U17046 (N_17046,N_16716,N_16785);
nand U17047 (N_17047,N_16826,N_16755);
and U17048 (N_17048,N_16891,N_16884);
xor U17049 (N_17049,N_16670,N_16984);
nand U17050 (N_17050,N_16823,N_16729);
nor U17051 (N_17051,N_16509,N_16970);
xor U17052 (N_17052,N_16833,N_16951);
nand U17053 (N_17053,N_16912,N_16642);
nand U17054 (N_17054,N_16894,N_16635);
nand U17055 (N_17055,N_16536,N_16892);
and U17056 (N_17056,N_16740,N_16705);
or U17057 (N_17057,N_16646,N_16754);
and U17058 (N_17058,N_16901,N_16503);
and U17059 (N_17059,N_16888,N_16606);
and U17060 (N_17060,N_16511,N_16788);
nand U17061 (N_17061,N_16599,N_16882);
and U17062 (N_17062,N_16559,N_16521);
nand U17063 (N_17063,N_16848,N_16620);
nor U17064 (N_17064,N_16750,N_16669);
nand U17065 (N_17065,N_16977,N_16652);
nor U17066 (N_17066,N_16684,N_16629);
and U17067 (N_17067,N_16628,N_16959);
nor U17068 (N_17068,N_16624,N_16742);
nor U17069 (N_17069,N_16512,N_16758);
nand U17070 (N_17070,N_16701,N_16960);
nor U17071 (N_17071,N_16749,N_16853);
xnor U17072 (N_17072,N_16517,N_16622);
nor U17073 (N_17073,N_16829,N_16938);
nor U17074 (N_17074,N_16548,N_16551);
or U17075 (N_17075,N_16715,N_16500);
and U17076 (N_17076,N_16897,N_16565);
xnor U17077 (N_17077,N_16995,N_16948);
nor U17078 (N_17078,N_16641,N_16547);
xor U17079 (N_17079,N_16648,N_16865);
nand U17080 (N_17080,N_16694,N_16588);
nor U17081 (N_17081,N_16846,N_16910);
nor U17082 (N_17082,N_16769,N_16777);
nor U17083 (N_17083,N_16562,N_16860);
nand U17084 (N_17084,N_16924,N_16837);
xnor U17085 (N_17085,N_16578,N_16703);
nand U17086 (N_17086,N_16616,N_16655);
nor U17087 (N_17087,N_16608,N_16602);
nor U17088 (N_17088,N_16572,N_16558);
nand U17089 (N_17089,N_16665,N_16795);
nor U17090 (N_17090,N_16604,N_16866);
and U17091 (N_17091,N_16957,N_16662);
or U17092 (N_17092,N_16890,N_16986);
or U17093 (N_17093,N_16821,N_16981);
nand U17094 (N_17094,N_16771,N_16998);
nand U17095 (N_17095,N_16834,N_16903);
nor U17096 (N_17096,N_16685,N_16719);
or U17097 (N_17097,N_16816,N_16739);
nand U17098 (N_17098,N_16581,N_16794);
xor U17099 (N_17099,N_16946,N_16690);
and U17100 (N_17100,N_16594,N_16613);
nand U17101 (N_17101,N_16675,N_16759);
nand U17102 (N_17102,N_16876,N_16667);
and U17103 (N_17103,N_16555,N_16789);
and U17104 (N_17104,N_16809,N_16626);
nand U17105 (N_17105,N_16818,N_16733);
nor U17106 (N_17106,N_16858,N_16935);
nor U17107 (N_17107,N_16576,N_16812);
and U17108 (N_17108,N_16781,N_16563);
or U17109 (N_17109,N_16680,N_16566);
nor U17110 (N_17110,N_16933,N_16671);
nand U17111 (N_17111,N_16593,N_16695);
nor U17112 (N_17112,N_16856,N_16569);
xor U17113 (N_17113,N_16550,N_16696);
and U17114 (N_17114,N_16954,N_16950);
and U17115 (N_17115,N_16969,N_16502);
and U17116 (N_17116,N_16735,N_16520);
nor U17117 (N_17117,N_16612,N_16805);
nor U17118 (N_17118,N_16908,N_16598);
nor U17119 (N_17119,N_16643,N_16516);
nor U17120 (N_17120,N_16723,N_16538);
xor U17121 (N_17121,N_16862,N_16796);
nand U17122 (N_17122,N_16741,N_16744);
or U17123 (N_17123,N_16878,N_16544);
and U17124 (N_17124,N_16975,N_16609);
or U17125 (N_17125,N_16752,N_16615);
xor U17126 (N_17126,N_16838,N_16929);
xnor U17127 (N_17127,N_16914,N_16819);
xnor U17128 (N_17128,N_16831,N_16965);
or U17129 (N_17129,N_16808,N_16779);
nand U17130 (N_17130,N_16790,N_16745);
and U17131 (N_17131,N_16964,N_16896);
nand U17132 (N_17132,N_16656,N_16724);
and U17133 (N_17133,N_16945,N_16786);
and U17134 (N_17134,N_16541,N_16840);
nor U17135 (N_17135,N_16844,N_16681);
nor U17136 (N_17136,N_16589,N_16722);
xnor U17137 (N_17137,N_16686,N_16867);
xor U17138 (N_17138,N_16782,N_16532);
xor U17139 (N_17139,N_16508,N_16757);
nand U17140 (N_17140,N_16872,N_16654);
xnor U17141 (N_17141,N_16531,N_16647);
or U17142 (N_17142,N_16692,N_16784);
or U17143 (N_17143,N_16637,N_16514);
and U17144 (N_17144,N_16601,N_16704);
or U17145 (N_17145,N_16610,N_16845);
xor U17146 (N_17146,N_16753,N_16800);
and U17147 (N_17147,N_16734,N_16631);
or U17148 (N_17148,N_16523,N_16543);
and U17149 (N_17149,N_16649,N_16900);
or U17150 (N_17150,N_16727,N_16659);
nor U17151 (N_17151,N_16525,N_16726);
nor U17152 (N_17152,N_16822,N_16811);
nand U17153 (N_17153,N_16625,N_16683);
xor U17154 (N_17154,N_16721,N_16596);
or U17155 (N_17155,N_16944,N_16875);
and U17156 (N_17156,N_16537,N_16841);
nand U17157 (N_17157,N_16881,N_16592);
and U17158 (N_17158,N_16852,N_16772);
xor U17159 (N_17159,N_16830,N_16720);
xor U17160 (N_17160,N_16958,N_16760);
or U17161 (N_17161,N_16774,N_16994);
or U17162 (N_17162,N_16568,N_16961);
or U17163 (N_17163,N_16968,N_16850);
and U17164 (N_17164,N_16590,N_16766);
nor U17165 (N_17165,N_16839,N_16718);
nor U17166 (N_17166,N_16515,N_16645);
and U17167 (N_17167,N_16835,N_16693);
nand U17168 (N_17168,N_16571,N_16732);
nor U17169 (N_17169,N_16899,N_16776);
xor U17170 (N_17170,N_16895,N_16600);
nor U17171 (N_17171,N_16921,N_16714);
or U17172 (N_17172,N_16561,N_16913);
nand U17173 (N_17173,N_16634,N_16504);
or U17174 (N_17174,N_16632,N_16639);
xnor U17175 (N_17175,N_16877,N_16621);
or U17176 (N_17176,N_16827,N_16925);
xor U17177 (N_17177,N_16930,N_16751);
or U17178 (N_17178,N_16668,N_16556);
nand U17179 (N_17179,N_16762,N_16851);
nor U17180 (N_17180,N_16513,N_16842);
and U17181 (N_17181,N_16584,N_16564);
nor U17182 (N_17182,N_16985,N_16990);
xnor U17183 (N_17183,N_16527,N_16941);
nand U17184 (N_17184,N_16815,N_16545);
or U17185 (N_17185,N_16864,N_16747);
and U17186 (N_17186,N_16660,N_16528);
and U17187 (N_17187,N_16712,N_16605);
or U17188 (N_17188,N_16736,N_16883);
nand U17189 (N_17189,N_16579,N_16983);
nor U17190 (N_17190,N_16698,N_16529);
nor U17191 (N_17191,N_16730,N_16911);
nor U17192 (N_17192,N_16677,N_16928);
nand U17193 (N_17193,N_16988,N_16768);
nor U17194 (N_17194,N_16678,N_16927);
nor U17195 (N_17195,N_16915,N_16886);
xnor U17196 (N_17196,N_16971,N_16780);
nor U17197 (N_17197,N_16802,N_16651);
nand U17198 (N_17198,N_16535,N_16676);
and U17199 (N_17199,N_16688,N_16530);
nor U17200 (N_17200,N_16582,N_16583);
nand U17201 (N_17201,N_16849,N_16999);
or U17202 (N_17202,N_16764,N_16552);
or U17203 (N_17203,N_16868,N_16533);
or U17204 (N_17204,N_16710,N_16807);
nand U17205 (N_17205,N_16917,N_16871);
or U17206 (N_17206,N_16595,N_16799);
nand U17207 (N_17207,N_16737,N_16619);
or U17208 (N_17208,N_16567,N_16526);
or U17209 (N_17209,N_16518,N_16711);
or U17210 (N_17210,N_16553,N_16770);
or U17211 (N_17211,N_16731,N_16775);
nor U17212 (N_17212,N_16793,N_16554);
and U17213 (N_17213,N_16798,N_16738);
nor U17214 (N_17214,N_16689,N_16748);
nor U17215 (N_17215,N_16743,N_16557);
xnor U17216 (N_17216,N_16773,N_16972);
xnor U17217 (N_17217,N_16869,N_16905);
and U17218 (N_17218,N_16934,N_16765);
and U17219 (N_17219,N_16936,N_16746);
nand U17220 (N_17220,N_16810,N_16918);
or U17221 (N_17221,N_16963,N_16580);
xnor U17222 (N_17222,N_16611,N_16932);
xnor U17223 (N_17223,N_16644,N_16916);
and U17224 (N_17224,N_16926,N_16955);
nor U17225 (N_17225,N_16992,N_16653);
xor U17226 (N_17226,N_16524,N_16937);
and U17227 (N_17227,N_16980,N_16591);
nand U17228 (N_17228,N_16920,N_16939);
or U17229 (N_17229,N_16657,N_16603);
nor U17230 (N_17230,N_16922,N_16978);
xor U17231 (N_17231,N_16539,N_16967);
xor U17232 (N_17232,N_16577,N_16952);
nor U17233 (N_17233,N_16931,N_16549);
and U17234 (N_17234,N_16673,N_16947);
nand U17235 (N_17235,N_16843,N_16893);
xor U17236 (N_17236,N_16907,N_16889);
nand U17237 (N_17237,N_16585,N_16640);
xnor U17238 (N_17238,N_16874,N_16791);
xnor U17239 (N_17239,N_16691,N_16663);
xor U17240 (N_17240,N_16847,N_16989);
xnor U17241 (N_17241,N_16725,N_16859);
xnor U17242 (N_17242,N_16906,N_16633);
or U17243 (N_17243,N_16956,N_16996);
xor U17244 (N_17244,N_16940,N_16617);
xnor U17245 (N_17245,N_16953,N_16672);
nor U17246 (N_17246,N_16873,N_16700);
xnor U17247 (N_17247,N_16702,N_16909);
nand U17248 (N_17248,N_16575,N_16679);
or U17249 (N_17249,N_16709,N_16783);
and U17250 (N_17250,N_16571,N_16601);
or U17251 (N_17251,N_16540,N_16813);
and U17252 (N_17252,N_16918,N_16646);
nand U17253 (N_17253,N_16725,N_16950);
nand U17254 (N_17254,N_16717,N_16944);
or U17255 (N_17255,N_16985,N_16562);
xor U17256 (N_17256,N_16631,N_16639);
nand U17257 (N_17257,N_16822,N_16971);
or U17258 (N_17258,N_16612,N_16966);
nand U17259 (N_17259,N_16815,N_16871);
xnor U17260 (N_17260,N_16626,N_16621);
or U17261 (N_17261,N_16999,N_16795);
and U17262 (N_17262,N_16998,N_16812);
xor U17263 (N_17263,N_16702,N_16860);
or U17264 (N_17264,N_16742,N_16939);
and U17265 (N_17265,N_16616,N_16618);
and U17266 (N_17266,N_16817,N_16934);
xor U17267 (N_17267,N_16963,N_16899);
or U17268 (N_17268,N_16971,N_16594);
nor U17269 (N_17269,N_16715,N_16514);
and U17270 (N_17270,N_16653,N_16722);
and U17271 (N_17271,N_16507,N_16627);
or U17272 (N_17272,N_16759,N_16990);
and U17273 (N_17273,N_16777,N_16655);
xnor U17274 (N_17274,N_16796,N_16693);
nand U17275 (N_17275,N_16890,N_16785);
or U17276 (N_17276,N_16600,N_16820);
nor U17277 (N_17277,N_16829,N_16682);
or U17278 (N_17278,N_16894,N_16700);
nor U17279 (N_17279,N_16538,N_16664);
and U17280 (N_17280,N_16702,N_16840);
or U17281 (N_17281,N_16752,N_16662);
and U17282 (N_17282,N_16994,N_16550);
xnor U17283 (N_17283,N_16642,N_16581);
or U17284 (N_17284,N_16724,N_16629);
and U17285 (N_17285,N_16716,N_16533);
or U17286 (N_17286,N_16943,N_16907);
nand U17287 (N_17287,N_16599,N_16696);
nor U17288 (N_17288,N_16644,N_16827);
nor U17289 (N_17289,N_16945,N_16648);
and U17290 (N_17290,N_16507,N_16774);
or U17291 (N_17291,N_16676,N_16995);
or U17292 (N_17292,N_16960,N_16974);
nor U17293 (N_17293,N_16759,N_16894);
or U17294 (N_17294,N_16707,N_16941);
xor U17295 (N_17295,N_16505,N_16541);
or U17296 (N_17296,N_16701,N_16605);
nand U17297 (N_17297,N_16909,N_16949);
nor U17298 (N_17298,N_16766,N_16890);
xnor U17299 (N_17299,N_16789,N_16544);
nand U17300 (N_17300,N_16584,N_16646);
nor U17301 (N_17301,N_16856,N_16521);
and U17302 (N_17302,N_16716,N_16976);
and U17303 (N_17303,N_16695,N_16591);
nand U17304 (N_17304,N_16971,N_16641);
nor U17305 (N_17305,N_16719,N_16778);
or U17306 (N_17306,N_16604,N_16964);
nor U17307 (N_17307,N_16837,N_16621);
or U17308 (N_17308,N_16677,N_16705);
nand U17309 (N_17309,N_16822,N_16528);
and U17310 (N_17310,N_16633,N_16688);
nor U17311 (N_17311,N_16548,N_16879);
or U17312 (N_17312,N_16787,N_16760);
nor U17313 (N_17313,N_16718,N_16628);
and U17314 (N_17314,N_16937,N_16856);
nand U17315 (N_17315,N_16697,N_16666);
and U17316 (N_17316,N_16572,N_16681);
nor U17317 (N_17317,N_16820,N_16565);
or U17318 (N_17318,N_16851,N_16857);
or U17319 (N_17319,N_16598,N_16754);
nand U17320 (N_17320,N_16953,N_16521);
and U17321 (N_17321,N_16987,N_16525);
xnor U17322 (N_17322,N_16676,N_16670);
nand U17323 (N_17323,N_16535,N_16910);
xnor U17324 (N_17324,N_16537,N_16898);
nor U17325 (N_17325,N_16764,N_16915);
nand U17326 (N_17326,N_16796,N_16568);
or U17327 (N_17327,N_16775,N_16924);
or U17328 (N_17328,N_16868,N_16590);
nor U17329 (N_17329,N_16696,N_16606);
nor U17330 (N_17330,N_16571,N_16604);
xor U17331 (N_17331,N_16576,N_16807);
nand U17332 (N_17332,N_16937,N_16994);
xnor U17333 (N_17333,N_16868,N_16975);
and U17334 (N_17334,N_16885,N_16987);
or U17335 (N_17335,N_16703,N_16551);
or U17336 (N_17336,N_16776,N_16821);
nor U17337 (N_17337,N_16925,N_16831);
and U17338 (N_17338,N_16587,N_16816);
xnor U17339 (N_17339,N_16943,N_16575);
and U17340 (N_17340,N_16968,N_16993);
nand U17341 (N_17341,N_16713,N_16919);
or U17342 (N_17342,N_16563,N_16913);
nand U17343 (N_17343,N_16548,N_16560);
nor U17344 (N_17344,N_16821,N_16720);
or U17345 (N_17345,N_16691,N_16929);
nor U17346 (N_17346,N_16723,N_16574);
or U17347 (N_17347,N_16998,N_16880);
xor U17348 (N_17348,N_16949,N_16663);
nor U17349 (N_17349,N_16589,N_16574);
and U17350 (N_17350,N_16953,N_16802);
xnor U17351 (N_17351,N_16598,N_16619);
nor U17352 (N_17352,N_16849,N_16588);
or U17353 (N_17353,N_16759,N_16927);
nor U17354 (N_17354,N_16844,N_16962);
nand U17355 (N_17355,N_16531,N_16894);
xor U17356 (N_17356,N_16655,N_16780);
or U17357 (N_17357,N_16917,N_16845);
nand U17358 (N_17358,N_16926,N_16625);
xnor U17359 (N_17359,N_16616,N_16657);
or U17360 (N_17360,N_16751,N_16970);
nor U17361 (N_17361,N_16682,N_16576);
and U17362 (N_17362,N_16998,N_16617);
or U17363 (N_17363,N_16718,N_16556);
and U17364 (N_17364,N_16813,N_16546);
xor U17365 (N_17365,N_16900,N_16685);
or U17366 (N_17366,N_16767,N_16753);
and U17367 (N_17367,N_16992,N_16785);
xor U17368 (N_17368,N_16525,N_16757);
and U17369 (N_17369,N_16581,N_16635);
and U17370 (N_17370,N_16740,N_16676);
nand U17371 (N_17371,N_16949,N_16568);
nor U17372 (N_17372,N_16711,N_16856);
nand U17373 (N_17373,N_16623,N_16943);
xnor U17374 (N_17374,N_16686,N_16518);
xnor U17375 (N_17375,N_16741,N_16594);
xnor U17376 (N_17376,N_16844,N_16785);
or U17377 (N_17377,N_16989,N_16747);
and U17378 (N_17378,N_16595,N_16748);
and U17379 (N_17379,N_16562,N_16725);
nand U17380 (N_17380,N_16940,N_16828);
xor U17381 (N_17381,N_16730,N_16529);
nor U17382 (N_17382,N_16990,N_16589);
nand U17383 (N_17383,N_16833,N_16764);
and U17384 (N_17384,N_16502,N_16790);
and U17385 (N_17385,N_16768,N_16736);
nor U17386 (N_17386,N_16734,N_16836);
and U17387 (N_17387,N_16772,N_16978);
xor U17388 (N_17388,N_16517,N_16522);
and U17389 (N_17389,N_16877,N_16710);
and U17390 (N_17390,N_16870,N_16752);
nor U17391 (N_17391,N_16830,N_16962);
or U17392 (N_17392,N_16757,N_16561);
nand U17393 (N_17393,N_16502,N_16710);
or U17394 (N_17394,N_16942,N_16569);
and U17395 (N_17395,N_16864,N_16644);
nor U17396 (N_17396,N_16611,N_16684);
and U17397 (N_17397,N_16546,N_16701);
xor U17398 (N_17398,N_16505,N_16745);
or U17399 (N_17399,N_16887,N_16883);
or U17400 (N_17400,N_16660,N_16669);
and U17401 (N_17401,N_16881,N_16924);
nor U17402 (N_17402,N_16525,N_16686);
nor U17403 (N_17403,N_16662,N_16825);
nand U17404 (N_17404,N_16626,N_16713);
xor U17405 (N_17405,N_16829,N_16797);
or U17406 (N_17406,N_16850,N_16566);
or U17407 (N_17407,N_16905,N_16871);
and U17408 (N_17408,N_16954,N_16506);
nand U17409 (N_17409,N_16705,N_16633);
nand U17410 (N_17410,N_16665,N_16805);
nand U17411 (N_17411,N_16527,N_16550);
xor U17412 (N_17412,N_16810,N_16870);
xor U17413 (N_17413,N_16520,N_16785);
or U17414 (N_17414,N_16839,N_16607);
nand U17415 (N_17415,N_16598,N_16947);
nor U17416 (N_17416,N_16889,N_16839);
or U17417 (N_17417,N_16697,N_16859);
nand U17418 (N_17418,N_16780,N_16528);
nand U17419 (N_17419,N_16650,N_16874);
and U17420 (N_17420,N_16813,N_16956);
and U17421 (N_17421,N_16875,N_16835);
and U17422 (N_17422,N_16887,N_16930);
nand U17423 (N_17423,N_16615,N_16932);
and U17424 (N_17424,N_16946,N_16506);
or U17425 (N_17425,N_16654,N_16944);
and U17426 (N_17426,N_16859,N_16686);
nor U17427 (N_17427,N_16771,N_16874);
and U17428 (N_17428,N_16880,N_16633);
and U17429 (N_17429,N_16809,N_16673);
nor U17430 (N_17430,N_16719,N_16979);
or U17431 (N_17431,N_16833,N_16986);
and U17432 (N_17432,N_16758,N_16682);
and U17433 (N_17433,N_16835,N_16983);
nor U17434 (N_17434,N_16787,N_16909);
nor U17435 (N_17435,N_16614,N_16625);
nand U17436 (N_17436,N_16517,N_16857);
or U17437 (N_17437,N_16888,N_16557);
and U17438 (N_17438,N_16699,N_16622);
nand U17439 (N_17439,N_16906,N_16689);
nor U17440 (N_17440,N_16543,N_16801);
nor U17441 (N_17441,N_16794,N_16658);
nand U17442 (N_17442,N_16589,N_16741);
xor U17443 (N_17443,N_16702,N_16981);
and U17444 (N_17444,N_16602,N_16546);
nor U17445 (N_17445,N_16511,N_16738);
nand U17446 (N_17446,N_16855,N_16973);
nand U17447 (N_17447,N_16566,N_16761);
nor U17448 (N_17448,N_16677,N_16947);
or U17449 (N_17449,N_16582,N_16717);
xor U17450 (N_17450,N_16818,N_16545);
nand U17451 (N_17451,N_16974,N_16676);
nand U17452 (N_17452,N_16505,N_16863);
or U17453 (N_17453,N_16979,N_16981);
and U17454 (N_17454,N_16711,N_16951);
nand U17455 (N_17455,N_16894,N_16822);
xor U17456 (N_17456,N_16891,N_16663);
and U17457 (N_17457,N_16920,N_16634);
xor U17458 (N_17458,N_16906,N_16772);
nand U17459 (N_17459,N_16726,N_16733);
nand U17460 (N_17460,N_16968,N_16683);
or U17461 (N_17461,N_16561,N_16634);
and U17462 (N_17462,N_16680,N_16835);
and U17463 (N_17463,N_16826,N_16778);
and U17464 (N_17464,N_16510,N_16538);
nor U17465 (N_17465,N_16891,N_16621);
or U17466 (N_17466,N_16854,N_16568);
nand U17467 (N_17467,N_16845,N_16647);
xor U17468 (N_17468,N_16989,N_16990);
and U17469 (N_17469,N_16703,N_16840);
xor U17470 (N_17470,N_16922,N_16798);
and U17471 (N_17471,N_16569,N_16543);
nand U17472 (N_17472,N_16940,N_16542);
xnor U17473 (N_17473,N_16646,N_16693);
or U17474 (N_17474,N_16700,N_16893);
and U17475 (N_17475,N_16652,N_16938);
nand U17476 (N_17476,N_16939,N_16804);
xnor U17477 (N_17477,N_16972,N_16883);
nor U17478 (N_17478,N_16937,N_16823);
and U17479 (N_17479,N_16511,N_16730);
and U17480 (N_17480,N_16997,N_16738);
and U17481 (N_17481,N_16931,N_16570);
xnor U17482 (N_17482,N_16995,N_16561);
or U17483 (N_17483,N_16904,N_16768);
or U17484 (N_17484,N_16685,N_16786);
xnor U17485 (N_17485,N_16879,N_16927);
and U17486 (N_17486,N_16875,N_16547);
and U17487 (N_17487,N_16777,N_16861);
or U17488 (N_17488,N_16548,N_16835);
xnor U17489 (N_17489,N_16524,N_16688);
nand U17490 (N_17490,N_16575,N_16652);
nor U17491 (N_17491,N_16574,N_16841);
or U17492 (N_17492,N_16531,N_16874);
xnor U17493 (N_17493,N_16539,N_16685);
or U17494 (N_17494,N_16920,N_16531);
xnor U17495 (N_17495,N_16772,N_16697);
and U17496 (N_17496,N_16509,N_16694);
and U17497 (N_17497,N_16555,N_16871);
nand U17498 (N_17498,N_16671,N_16543);
or U17499 (N_17499,N_16517,N_16815);
nor U17500 (N_17500,N_17165,N_17248);
nor U17501 (N_17501,N_17445,N_17250);
nand U17502 (N_17502,N_17437,N_17149);
nor U17503 (N_17503,N_17369,N_17223);
xnor U17504 (N_17504,N_17345,N_17358);
or U17505 (N_17505,N_17498,N_17129);
and U17506 (N_17506,N_17231,N_17068);
nand U17507 (N_17507,N_17191,N_17113);
and U17508 (N_17508,N_17044,N_17254);
xor U17509 (N_17509,N_17204,N_17153);
xor U17510 (N_17510,N_17399,N_17132);
nand U17511 (N_17511,N_17105,N_17266);
nand U17512 (N_17512,N_17481,N_17324);
xnor U17513 (N_17513,N_17354,N_17385);
or U17514 (N_17514,N_17241,N_17334);
or U17515 (N_17515,N_17446,N_17147);
nand U17516 (N_17516,N_17283,N_17387);
and U17517 (N_17517,N_17102,N_17476);
nor U17518 (N_17518,N_17257,N_17066);
and U17519 (N_17519,N_17171,N_17252);
and U17520 (N_17520,N_17449,N_17470);
nor U17521 (N_17521,N_17074,N_17025);
and U17522 (N_17522,N_17421,N_17318);
or U17523 (N_17523,N_17383,N_17403);
xnor U17524 (N_17524,N_17036,N_17062);
or U17525 (N_17525,N_17145,N_17349);
or U17526 (N_17526,N_17336,N_17377);
nand U17527 (N_17527,N_17039,N_17396);
nor U17528 (N_17528,N_17016,N_17169);
nand U17529 (N_17529,N_17031,N_17010);
or U17530 (N_17530,N_17404,N_17320);
and U17531 (N_17531,N_17144,N_17456);
and U17532 (N_17532,N_17014,N_17269);
nor U17533 (N_17533,N_17157,N_17143);
and U17534 (N_17534,N_17209,N_17285);
nor U17535 (N_17535,N_17356,N_17221);
or U17536 (N_17536,N_17214,N_17020);
nand U17537 (N_17537,N_17187,N_17493);
and U17538 (N_17538,N_17071,N_17392);
xnor U17539 (N_17539,N_17482,N_17466);
nor U17540 (N_17540,N_17263,N_17409);
xor U17541 (N_17541,N_17402,N_17453);
xnor U17542 (N_17542,N_17452,N_17448);
and U17543 (N_17543,N_17242,N_17131);
nor U17544 (N_17544,N_17339,N_17175);
nand U17545 (N_17545,N_17299,N_17003);
xor U17546 (N_17546,N_17056,N_17229);
nand U17547 (N_17547,N_17027,N_17217);
and U17548 (N_17548,N_17183,N_17467);
xor U17549 (N_17549,N_17009,N_17367);
or U17550 (N_17550,N_17422,N_17152);
and U17551 (N_17551,N_17479,N_17473);
or U17552 (N_17552,N_17045,N_17284);
or U17553 (N_17553,N_17150,N_17096);
xor U17554 (N_17554,N_17206,N_17117);
and U17555 (N_17555,N_17465,N_17220);
or U17556 (N_17556,N_17451,N_17215);
or U17557 (N_17557,N_17281,N_17464);
or U17558 (N_17558,N_17468,N_17355);
or U17559 (N_17559,N_17291,N_17041);
or U17560 (N_17560,N_17368,N_17256);
xnor U17561 (N_17561,N_17099,N_17158);
nand U17562 (N_17562,N_17076,N_17378);
or U17563 (N_17563,N_17161,N_17490);
or U17564 (N_17564,N_17443,N_17048);
xor U17565 (N_17565,N_17127,N_17001);
and U17566 (N_17566,N_17251,N_17277);
and U17567 (N_17567,N_17111,N_17006);
nor U17568 (N_17568,N_17059,N_17416);
xnor U17569 (N_17569,N_17365,N_17093);
or U17570 (N_17570,N_17271,N_17095);
or U17571 (N_17571,N_17239,N_17330);
and U17572 (N_17572,N_17112,N_17103);
and U17573 (N_17573,N_17347,N_17015);
xnor U17574 (N_17574,N_17125,N_17176);
and U17575 (N_17575,N_17091,N_17194);
and U17576 (N_17576,N_17188,N_17341);
xor U17577 (N_17577,N_17382,N_17186);
or U17578 (N_17578,N_17434,N_17494);
or U17579 (N_17579,N_17134,N_17070);
nand U17580 (N_17580,N_17380,N_17342);
nor U17581 (N_17581,N_17160,N_17499);
nand U17582 (N_17582,N_17412,N_17234);
xnor U17583 (N_17583,N_17233,N_17197);
or U17584 (N_17584,N_17037,N_17474);
nand U17585 (N_17585,N_17357,N_17272);
xnor U17586 (N_17586,N_17433,N_17237);
and U17587 (N_17587,N_17088,N_17371);
or U17588 (N_17588,N_17447,N_17323);
or U17589 (N_17589,N_17072,N_17028);
nor U17590 (N_17590,N_17350,N_17172);
nor U17591 (N_17591,N_17075,N_17236);
nand U17592 (N_17592,N_17340,N_17436);
and U17593 (N_17593,N_17026,N_17331);
or U17594 (N_17594,N_17139,N_17244);
or U17595 (N_17595,N_17430,N_17114);
or U17596 (N_17596,N_17492,N_17258);
and U17597 (N_17597,N_17115,N_17487);
nand U17598 (N_17598,N_17261,N_17000);
xnor U17599 (N_17599,N_17282,N_17007);
or U17600 (N_17600,N_17270,N_17109);
nor U17601 (N_17601,N_17363,N_17346);
or U17602 (N_17602,N_17118,N_17344);
xor U17603 (N_17603,N_17373,N_17084);
or U17604 (N_17604,N_17080,N_17213);
xor U17605 (N_17605,N_17138,N_17064);
and U17606 (N_17606,N_17401,N_17338);
and U17607 (N_17607,N_17394,N_17240);
nand U17608 (N_17608,N_17224,N_17264);
xor U17609 (N_17609,N_17246,N_17051);
nor U17610 (N_17610,N_17086,N_17055);
and U17611 (N_17611,N_17216,N_17301);
xor U17612 (N_17612,N_17019,N_17413);
nor U17613 (N_17613,N_17124,N_17418);
nand U17614 (N_17614,N_17410,N_17222);
nand U17615 (N_17615,N_17312,N_17292);
or U17616 (N_17616,N_17079,N_17126);
nand U17617 (N_17617,N_17249,N_17419);
nand U17618 (N_17618,N_17211,N_17397);
xor U17619 (N_17619,N_17218,N_17107);
nand U17620 (N_17620,N_17495,N_17173);
or U17621 (N_17621,N_17278,N_17327);
or U17622 (N_17622,N_17463,N_17438);
nor U17623 (N_17623,N_17203,N_17322);
and U17624 (N_17624,N_17276,N_17290);
nand U17625 (N_17625,N_17415,N_17302);
nor U17626 (N_17626,N_17198,N_17018);
and U17627 (N_17627,N_17423,N_17130);
nor U17628 (N_17628,N_17428,N_17458);
and U17629 (N_17629,N_17489,N_17308);
nor U17630 (N_17630,N_17178,N_17067);
nor U17631 (N_17631,N_17304,N_17179);
nor U17632 (N_17632,N_17348,N_17008);
nor U17633 (N_17633,N_17405,N_17119);
nand U17634 (N_17634,N_17230,N_17444);
nand U17635 (N_17635,N_17073,N_17366);
nand U17636 (N_17636,N_17496,N_17329);
nor U17637 (N_17637,N_17200,N_17390);
nor U17638 (N_17638,N_17477,N_17395);
and U17639 (N_17639,N_17455,N_17136);
or U17640 (N_17640,N_17488,N_17253);
nand U17641 (N_17641,N_17441,N_17189);
and U17642 (N_17642,N_17030,N_17040);
and U17643 (N_17643,N_17137,N_17004);
nand U17644 (N_17644,N_17435,N_17052);
nand U17645 (N_17645,N_17287,N_17310);
or U17646 (N_17646,N_17021,N_17328);
and U17647 (N_17647,N_17303,N_17128);
or U17648 (N_17648,N_17012,N_17089);
nor U17649 (N_17649,N_17332,N_17227);
nand U17650 (N_17650,N_17199,N_17309);
and U17651 (N_17651,N_17120,N_17225);
xor U17652 (N_17652,N_17315,N_17391);
or U17653 (N_17653,N_17190,N_17351);
or U17654 (N_17654,N_17212,N_17029);
nand U17655 (N_17655,N_17011,N_17123);
xnor U17656 (N_17656,N_17289,N_17226);
nand U17657 (N_17657,N_17381,N_17427);
nor U17658 (N_17658,N_17353,N_17142);
xnor U17659 (N_17659,N_17462,N_17060);
or U17660 (N_17660,N_17228,N_17432);
nand U17661 (N_17661,N_17255,N_17243);
nor U17662 (N_17662,N_17259,N_17085);
and U17663 (N_17663,N_17219,N_17090);
and U17664 (N_17664,N_17431,N_17375);
nand U17665 (N_17665,N_17326,N_17185);
nand U17666 (N_17666,N_17440,N_17042);
nand U17667 (N_17667,N_17267,N_17038);
nor U17668 (N_17668,N_17374,N_17092);
or U17669 (N_17669,N_17098,N_17260);
and U17670 (N_17670,N_17081,N_17457);
xor U17671 (N_17671,N_17192,N_17155);
and U17672 (N_17672,N_17484,N_17022);
or U17673 (N_17673,N_17141,N_17472);
nand U17674 (N_17674,N_17478,N_17279);
nor U17675 (N_17675,N_17486,N_17298);
xor U17676 (N_17676,N_17097,N_17317);
and U17677 (N_17677,N_17497,N_17002);
or U17678 (N_17678,N_17400,N_17359);
nand U17679 (N_17679,N_17110,N_17491);
or U17680 (N_17680,N_17388,N_17274);
nor U17681 (N_17681,N_17170,N_17094);
xnor U17682 (N_17682,N_17406,N_17485);
or U17683 (N_17683,N_17047,N_17471);
nand U17684 (N_17684,N_17288,N_17439);
nand U17685 (N_17685,N_17083,N_17362);
or U17686 (N_17686,N_17193,N_17265);
or U17687 (N_17687,N_17293,N_17337);
nand U17688 (N_17688,N_17311,N_17316);
nor U17689 (N_17689,N_17177,N_17133);
or U17690 (N_17690,N_17370,N_17148);
xor U17691 (N_17691,N_17034,N_17164);
or U17692 (N_17692,N_17425,N_17013);
and U17693 (N_17693,N_17201,N_17386);
nor U17694 (N_17694,N_17364,N_17376);
nand U17695 (N_17695,N_17389,N_17426);
nand U17696 (N_17696,N_17154,N_17411);
xnor U17697 (N_17697,N_17166,N_17063);
or U17698 (N_17698,N_17294,N_17163);
nor U17699 (N_17699,N_17077,N_17162);
nor U17700 (N_17700,N_17296,N_17280);
nand U17701 (N_17701,N_17054,N_17033);
nand U17702 (N_17702,N_17005,N_17460);
nand U17703 (N_17703,N_17297,N_17069);
xor U17704 (N_17704,N_17101,N_17407);
xnor U17705 (N_17705,N_17450,N_17268);
and U17706 (N_17706,N_17417,N_17235);
or U17707 (N_17707,N_17307,N_17273);
or U17708 (N_17708,N_17319,N_17087);
xnor U17709 (N_17709,N_17049,N_17106);
and U17710 (N_17710,N_17343,N_17174);
or U17711 (N_17711,N_17061,N_17205);
nor U17712 (N_17712,N_17275,N_17286);
xor U17713 (N_17713,N_17306,N_17459);
xor U17714 (N_17714,N_17195,N_17454);
or U17715 (N_17715,N_17181,N_17082);
and U17716 (N_17716,N_17408,N_17180);
and U17717 (N_17717,N_17295,N_17167);
nand U17718 (N_17718,N_17325,N_17140);
or U17719 (N_17719,N_17361,N_17352);
xor U17720 (N_17720,N_17116,N_17065);
xor U17721 (N_17721,N_17483,N_17053);
nor U17722 (N_17722,N_17058,N_17121);
and U17723 (N_17723,N_17196,N_17057);
nor U17724 (N_17724,N_17314,N_17414);
and U17725 (N_17725,N_17469,N_17429);
or U17726 (N_17726,N_17156,N_17108);
nand U17727 (N_17727,N_17262,N_17043);
nor U17728 (N_17728,N_17393,N_17305);
and U17729 (N_17729,N_17104,N_17151);
nand U17730 (N_17730,N_17184,N_17122);
and U17731 (N_17731,N_17238,N_17379);
and U17732 (N_17732,N_17360,N_17135);
and U17733 (N_17733,N_17461,N_17046);
nor U17734 (N_17734,N_17480,N_17313);
nand U17735 (N_17735,N_17168,N_17424);
nand U17736 (N_17736,N_17100,N_17078);
or U17737 (N_17737,N_17398,N_17202);
and U17738 (N_17738,N_17159,N_17024);
nor U17739 (N_17739,N_17335,N_17321);
xor U17740 (N_17740,N_17247,N_17208);
or U17741 (N_17741,N_17333,N_17210);
xnor U17742 (N_17742,N_17035,N_17420);
nand U17743 (N_17743,N_17245,N_17182);
and U17744 (N_17744,N_17442,N_17207);
xnor U17745 (N_17745,N_17017,N_17232);
and U17746 (N_17746,N_17023,N_17384);
nand U17747 (N_17747,N_17300,N_17475);
or U17748 (N_17748,N_17050,N_17146);
xnor U17749 (N_17749,N_17032,N_17372);
nor U17750 (N_17750,N_17460,N_17452);
nor U17751 (N_17751,N_17065,N_17256);
or U17752 (N_17752,N_17156,N_17360);
nor U17753 (N_17753,N_17018,N_17461);
nand U17754 (N_17754,N_17442,N_17390);
or U17755 (N_17755,N_17279,N_17170);
or U17756 (N_17756,N_17298,N_17150);
nand U17757 (N_17757,N_17218,N_17083);
or U17758 (N_17758,N_17204,N_17341);
nand U17759 (N_17759,N_17001,N_17442);
nand U17760 (N_17760,N_17155,N_17157);
xor U17761 (N_17761,N_17461,N_17219);
and U17762 (N_17762,N_17290,N_17429);
nor U17763 (N_17763,N_17281,N_17080);
nand U17764 (N_17764,N_17102,N_17323);
nor U17765 (N_17765,N_17007,N_17177);
nand U17766 (N_17766,N_17271,N_17468);
xnor U17767 (N_17767,N_17047,N_17168);
and U17768 (N_17768,N_17135,N_17023);
nand U17769 (N_17769,N_17242,N_17477);
xor U17770 (N_17770,N_17097,N_17268);
and U17771 (N_17771,N_17216,N_17396);
nand U17772 (N_17772,N_17403,N_17374);
and U17773 (N_17773,N_17117,N_17264);
or U17774 (N_17774,N_17376,N_17100);
nor U17775 (N_17775,N_17233,N_17328);
xor U17776 (N_17776,N_17450,N_17252);
nor U17777 (N_17777,N_17036,N_17222);
or U17778 (N_17778,N_17487,N_17040);
nor U17779 (N_17779,N_17244,N_17217);
nor U17780 (N_17780,N_17026,N_17402);
nor U17781 (N_17781,N_17225,N_17270);
or U17782 (N_17782,N_17215,N_17494);
nand U17783 (N_17783,N_17291,N_17206);
xor U17784 (N_17784,N_17113,N_17344);
nor U17785 (N_17785,N_17081,N_17298);
nor U17786 (N_17786,N_17346,N_17155);
and U17787 (N_17787,N_17259,N_17412);
nand U17788 (N_17788,N_17134,N_17288);
and U17789 (N_17789,N_17185,N_17172);
nor U17790 (N_17790,N_17017,N_17256);
or U17791 (N_17791,N_17121,N_17129);
nand U17792 (N_17792,N_17139,N_17181);
nor U17793 (N_17793,N_17014,N_17071);
nand U17794 (N_17794,N_17358,N_17011);
and U17795 (N_17795,N_17443,N_17365);
xnor U17796 (N_17796,N_17429,N_17326);
or U17797 (N_17797,N_17131,N_17155);
and U17798 (N_17798,N_17015,N_17081);
or U17799 (N_17799,N_17112,N_17400);
nand U17800 (N_17800,N_17458,N_17362);
or U17801 (N_17801,N_17158,N_17423);
nand U17802 (N_17802,N_17089,N_17273);
nand U17803 (N_17803,N_17198,N_17315);
and U17804 (N_17804,N_17280,N_17259);
and U17805 (N_17805,N_17431,N_17448);
xor U17806 (N_17806,N_17174,N_17433);
and U17807 (N_17807,N_17282,N_17081);
and U17808 (N_17808,N_17052,N_17026);
xor U17809 (N_17809,N_17308,N_17451);
and U17810 (N_17810,N_17003,N_17183);
xnor U17811 (N_17811,N_17152,N_17475);
nand U17812 (N_17812,N_17048,N_17416);
xor U17813 (N_17813,N_17009,N_17424);
and U17814 (N_17814,N_17111,N_17101);
and U17815 (N_17815,N_17117,N_17225);
and U17816 (N_17816,N_17100,N_17152);
or U17817 (N_17817,N_17389,N_17371);
nor U17818 (N_17818,N_17431,N_17230);
or U17819 (N_17819,N_17418,N_17121);
nor U17820 (N_17820,N_17373,N_17079);
nor U17821 (N_17821,N_17389,N_17381);
nand U17822 (N_17822,N_17096,N_17048);
nand U17823 (N_17823,N_17181,N_17085);
nor U17824 (N_17824,N_17428,N_17317);
or U17825 (N_17825,N_17317,N_17379);
or U17826 (N_17826,N_17400,N_17269);
xor U17827 (N_17827,N_17266,N_17319);
nor U17828 (N_17828,N_17403,N_17129);
nor U17829 (N_17829,N_17232,N_17495);
xnor U17830 (N_17830,N_17462,N_17242);
or U17831 (N_17831,N_17003,N_17042);
or U17832 (N_17832,N_17323,N_17058);
xor U17833 (N_17833,N_17159,N_17384);
nand U17834 (N_17834,N_17415,N_17355);
nor U17835 (N_17835,N_17045,N_17059);
xnor U17836 (N_17836,N_17341,N_17302);
and U17837 (N_17837,N_17369,N_17316);
or U17838 (N_17838,N_17158,N_17061);
or U17839 (N_17839,N_17491,N_17118);
nand U17840 (N_17840,N_17216,N_17403);
and U17841 (N_17841,N_17258,N_17330);
and U17842 (N_17842,N_17446,N_17251);
nand U17843 (N_17843,N_17421,N_17331);
nor U17844 (N_17844,N_17250,N_17049);
xnor U17845 (N_17845,N_17018,N_17459);
nor U17846 (N_17846,N_17039,N_17411);
or U17847 (N_17847,N_17274,N_17169);
xnor U17848 (N_17848,N_17296,N_17214);
nand U17849 (N_17849,N_17469,N_17377);
or U17850 (N_17850,N_17195,N_17220);
nand U17851 (N_17851,N_17261,N_17401);
nor U17852 (N_17852,N_17147,N_17032);
nor U17853 (N_17853,N_17032,N_17382);
and U17854 (N_17854,N_17284,N_17446);
and U17855 (N_17855,N_17212,N_17396);
xnor U17856 (N_17856,N_17347,N_17221);
nor U17857 (N_17857,N_17183,N_17371);
nand U17858 (N_17858,N_17088,N_17188);
nor U17859 (N_17859,N_17352,N_17334);
nand U17860 (N_17860,N_17488,N_17197);
xnor U17861 (N_17861,N_17095,N_17187);
and U17862 (N_17862,N_17072,N_17261);
nor U17863 (N_17863,N_17200,N_17455);
xnor U17864 (N_17864,N_17391,N_17009);
nand U17865 (N_17865,N_17199,N_17153);
nor U17866 (N_17866,N_17364,N_17077);
nand U17867 (N_17867,N_17268,N_17159);
or U17868 (N_17868,N_17003,N_17498);
nor U17869 (N_17869,N_17456,N_17432);
xor U17870 (N_17870,N_17499,N_17099);
and U17871 (N_17871,N_17331,N_17335);
or U17872 (N_17872,N_17380,N_17434);
xnor U17873 (N_17873,N_17001,N_17469);
or U17874 (N_17874,N_17295,N_17144);
nand U17875 (N_17875,N_17252,N_17040);
nor U17876 (N_17876,N_17212,N_17342);
nand U17877 (N_17877,N_17285,N_17203);
nand U17878 (N_17878,N_17015,N_17011);
or U17879 (N_17879,N_17178,N_17169);
and U17880 (N_17880,N_17008,N_17408);
and U17881 (N_17881,N_17071,N_17216);
nand U17882 (N_17882,N_17474,N_17267);
and U17883 (N_17883,N_17130,N_17175);
nor U17884 (N_17884,N_17114,N_17263);
nand U17885 (N_17885,N_17434,N_17159);
xor U17886 (N_17886,N_17182,N_17447);
xnor U17887 (N_17887,N_17399,N_17356);
xnor U17888 (N_17888,N_17025,N_17249);
xor U17889 (N_17889,N_17300,N_17031);
nand U17890 (N_17890,N_17480,N_17349);
xor U17891 (N_17891,N_17267,N_17183);
xnor U17892 (N_17892,N_17079,N_17199);
nor U17893 (N_17893,N_17180,N_17429);
or U17894 (N_17894,N_17009,N_17086);
nor U17895 (N_17895,N_17018,N_17477);
or U17896 (N_17896,N_17041,N_17312);
and U17897 (N_17897,N_17441,N_17113);
xor U17898 (N_17898,N_17046,N_17218);
nand U17899 (N_17899,N_17385,N_17132);
or U17900 (N_17900,N_17268,N_17195);
or U17901 (N_17901,N_17295,N_17177);
and U17902 (N_17902,N_17412,N_17303);
or U17903 (N_17903,N_17239,N_17456);
xnor U17904 (N_17904,N_17466,N_17234);
nand U17905 (N_17905,N_17358,N_17402);
nand U17906 (N_17906,N_17072,N_17427);
nor U17907 (N_17907,N_17000,N_17129);
nand U17908 (N_17908,N_17149,N_17061);
and U17909 (N_17909,N_17103,N_17077);
nand U17910 (N_17910,N_17245,N_17352);
or U17911 (N_17911,N_17040,N_17242);
xnor U17912 (N_17912,N_17395,N_17183);
nor U17913 (N_17913,N_17495,N_17143);
or U17914 (N_17914,N_17485,N_17438);
xor U17915 (N_17915,N_17091,N_17414);
nand U17916 (N_17916,N_17021,N_17199);
and U17917 (N_17917,N_17431,N_17470);
xor U17918 (N_17918,N_17453,N_17220);
nand U17919 (N_17919,N_17423,N_17001);
nor U17920 (N_17920,N_17122,N_17076);
nor U17921 (N_17921,N_17452,N_17073);
nor U17922 (N_17922,N_17212,N_17000);
nor U17923 (N_17923,N_17481,N_17359);
xor U17924 (N_17924,N_17022,N_17367);
and U17925 (N_17925,N_17241,N_17158);
xnor U17926 (N_17926,N_17113,N_17437);
and U17927 (N_17927,N_17460,N_17337);
and U17928 (N_17928,N_17040,N_17026);
and U17929 (N_17929,N_17158,N_17049);
and U17930 (N_17930,N_17425,N_17239);
nor U17931 (N_17931,N_17001,N_17198);
and U17932 (N_17932,N_17405,N_17447);
nand U17933 (N_17933,N_17243,N_17485);
nand U17934 (N_17934,N_17277,N_17354);
nand U17935 (N_17935,N_17296,N_17169);
xor U17936 (N_17936,N_17233,N_17100);
and U17937 (N_17937,N_17122,N_17313);
or U17938 (N_17938,N_17258,N_17118);
nand U17939 (N_17939,N_17162,N_17331);
or U17940 (N_17940,N_17353,N_17497);
nor U17941 (N_17941,N_17098,N_17348);
nand U17942 (N_17942,N_17137,N_17442);
xor U17943 (N_17943,N_17270,N_17436);
nor U17944 (N_17944,N_17132,N_17128);
nor U17945 (N_17945,N_17483,N_17357);
nand U17946 (N_17946,N_17433,N_17296);
xor U17947 (N_17947,N_17026,N_17165);
nand U17948 (N_17948,N_17404,N_17418);
or U17949 (N_17949,N_17193,N_17328);
nor U17950 (N_17950,N_17112,N_17461);
or U17951 (N_17951,N_17407,N_17368);
and U17952 (N_17952,N_17318,N_17353);
nand U17953 (N_17953,N_17392,N_17015);
and U17954 (N_17954,N_17083,N_17053);
nand U17955 (N_17955,N_17112,N_17425);
nand U17956 (N_17956,N_17385,N_17487);
nor U17957 (N_17957,N_17211,N_17014);
xnor U17958 (N_17958,N_17488,N_17001);
nor U17959 (N_17959,N_17319,N_17130);
nor U17960 (N_17960,N_17234,N_17111);
xor U17961 (N_17961,N_17363,N_17081);
nor U17962 (N_17962,N_17092,N_17024);
nor U17963 (N_17963,N_17401,N_17352);
xor U17964 (N_17964,N_17048,N_17298);
nand U17965 (N_17965,N_17492,N_17374);
nand U17966 (N_17966,N_17392,N_17452);
nor U17967 (N_17967,N_17002,N_17320);
and U17968 (N_17968,N_17383,N_17206);
xnor U17969 (N_17969,N_17388,N_17257);
nand U17970 (N_17970,N_17467,N_17465);
xor U17971 (N_17971,N_17453,N_17097);
nand U17972 (N_17972,N_17140,N_17320);
nor U17973 (N_17973,N_17258,N_17432);
and U17974 (N_17974,N_17317,N_17033);
nand U17975 (N_17975,N_17314,N_17228);
nand U17976 (N_17976,N_17039,N_17306);
xnor U17977 (N_17977,N_17158,N_17374);
nor U17978 (N_17978,N_17013,N_17075);
and U17979 (N_17979,N_17317,N_17467);
xnor U17980 (N_17980,N_17467,N_17361);
nor U17981 (N_17981,N_17432,N_17156);
or U17982 (N_17982,N_17343,N_17405);
xor U17983 (N_17983,N_17419,N_17414);
xnor U17984 (N_17984,N_17099,N_17224);
and U17985 (N_17985,N_17338,N_17111);
nand U17986 (N_17986,N_17438,N_17393);
and U17987 (N_17987,N_17482,N_17467);
or U17988 (N_17988,N_17110,N_17494);
xor U17989 (N_17989,N_17300,N_17255);
nand U17990 (N_17990,N_17358,N_17165);
xnor U17991 (N_17991,N_17266,N_17001);
and U17992 (N_17992,N_17036,N_17076);
or U17993 (N_17993,N_17073,N_17470);
and U17994 (N_17994,N_17087,N_17476);
nor U17995 (N_17995,N_17341,N_17271);
nand U17996 (N_17996,N_17498,N_17278);
xor U17997 (N_17997,N_17491,N_17141);
xnor U17998 (N_17998,N_17242,N_17043);
nand U17999 (N_17999,N_17252,N_17200);
xnor U18000 (N_18000,N_17648,N_17515);
and U18001 (N_18001,N_17812,N_17641);
xnor U18002 (N_18002,N_17665,N_17957);
nor U18003 (N_18003,N_17654,N_17704);
or U18004 (N_18004,N_17593,N_17973);
xnor U18005 (N_18005,N_17892,N_17840);
nor U18006 (N_18006,N_17747,N_17563);
nor U18007 (N_18007,N_17612,N_17874);
or U18008 (N_18008,N_17666,N_17581);
nor U18009 (N_18009,N_17530,N_17958);
or U18010 (N_18010,N_17989,N_17520);
xor U18011 (N_18011,N_17643,N_17824);
xor U18012 (N_18012,N_17998,N_17568);
nor U18013 (N_18013,N_17866,N_17614);
or U18014 (N_18014,N_17619,N_17608);
or U18015 (N_18015,N_17625,N_17725);
nor U18016 (N_18016,N_17726,N_17735);
xnor U18017 (N_18017,N_17942,N_17660);
or U18018 (N_18018,N_17599,N_17683);
nor U18019 (N_18019,N_17750,N_17711);
and U18020 (N_18020,N_17823,N_17566);
nand U18021 (N_18021,N_17668,N_17736);
or U18022 (N_18022,N_17926,N_17871);
and U18023 (N_18023,N_17854,N_17542);
or U18024 (N_18024,N_17756,N_17510);
or U18025 (N_18025,N_17831,N_17797);
and U18026 (N_18026,N_17632,N_17502);
nand U18027 (N_18027,N_17946,N_17544);
and U18028 (N_18028,N_17754,N_17771);
xor U18029 (N_18029,N_17876,N_17557);
and U18030 (N_18030,N_17540,N_17622);
and U18031 (N_18031,N_17597,N_17609);
or U18032 (N_18032,N_17877,N_17807);
xnor U18033 (N_18033,N_17847,N_17737);
and U18034 (N_18034,N_17706,N_17729);
xnor U18035 (N_18035,N_17816,N_17999);
xnor U18036 (N_18036,N_17887,N_17921);
nor U18037 (N_18037,N_17522,N_17805);
nor U18038 (N_18038,N_17923,N_17821);
xor U18039 (N_18039,N_17889,N_17913);
or U18040 (N_18040,N_17903,N_17995);
and U18041 (N_18041,N_17664,N_17762);
and U18042 (N_18042,N_17810,N_17611);
or U18043 (N_18043,N_17959,N_17940);
and U18044 (N_18044,N_17616,N_17601);
nor U18045 (N_18045,N_17780,N_17813);
xnor U18046 (N_18046,N_17865,N_17948);
xnor U18047 (N_18047,N_17842,N_17993);
nand U18048 (N_18048,N_17784,N_17728);
nand U18049 (N_18049,N_17789,N_17734);
xnor U18050 (N_18050,N_17899,N_17945);
nor U18051 (N_18051,N_17752,N_17634);
xor U18052 (N_18052,N_17550,N_17523);
and U18053 (N_18053,N_17629,N_17739);
nand U18054 (N_18054,N_17577,N_17983);
nand U18055 (N_18055,N_17639,N_17825);
xor U18056 (N_18056,N_17873,N_17799);
xnor U18057 (N_18057,N_17981,N_17875);
nand U18058 (N_18058,N_17576,N_17732);
xnor U18059 (N_18059,N_17588,N_17953);
or U18060 (N_18060,N_17621,N_17943);
and U18061 (N_18061,N_17819,N_17602);
nand U18062 (N_18062,N_17642,N_17675);
or U18063 (N_18063,N_17992,N_17843);
and U18064 (N_18064,N_17846,N_17720);
nand U18065 (N_18065,N_17553,N_17900);
and U18066 (N_18066,N_17930,N_17518);
or U18067 (N_18067,N_17950,N_17638);
nand U18068 (N_18068,N_17769,N_17558);
and U18069 (N_18069,N_17982,N_17669);
or U18070 (N_18070,N_17538,N_17570);
nor U18071 (N_18071,N_17681,N_17988);
nor U18072 (N_18072,N_17727,N_17861);
and U18073 (N_18073,N_17549,N_17644);
xnor U18074 (N_18074,N_17961,N_17759);
xor U18075 (N_18075,N_17698,N_17994);
xnor U18076 (N_18076,N_17569,N_17925);
nand U18077 (N_18077,N_17891,N_17582);
and U18078 (N_18078,N_17917,N_17796);
or U18079 (N_18079,N_17909,N_17653);
and U18080 (N_18080,N_17979,N_17897);
or U18081 (N_18081,N_17938,N_17922);
nor U18082 (N_18082,N_17817,N_17844);
or U18083 (N_18083,N_17541,N_17676);
xor U18084 (N_18084,N_17578,N_17751);
nor U18085 (N_18085,N_17963,N_17630);
nor U18086 (N_18086,N_17969,N_17650);
xnor U18087 (N_18087,N_17802,N_17867);
xnor U18088 (N_18088,N_17770,N_17699);
nand U18089 (N_18089,N_17811,N_17855);
and U18090 (N_18090,N_17775,N_17710);
xnor U18091 (N_18091,N_17803,N_17667);
and U18092 (N_18092,N_17859,N_17898);
or U18093 (N_18093,N_17589,N_17693);
nand U18094 (N_18094,N_17934,N_17841);
and U18095 (N_18095,N_17907,N_17894);
xnor U18096 (N_18096,N_17856,N_17908);
and U18097 (N_18097,N_17765,N_17977);
nand U18098 (N_18098,N_17850,N_17543);
nor U18099 (N_18099,N_17504,N_17635);
nor U18100 (N_18100,N_17809,N_17741);
xnor U18101 (N_18101,N_17500,N_17748);
xor U18102 (N_18102,N_17529,N_17554);
nand U18103 (N_18103,N_17968,N_17620);
nor U18104 (N_18104,N_17610,N_17919);
or U18105 (N_18105,N_17997,N_17966);
or U18106 (N_18106,N_17857,N_17848);
and U18107 (N_18107,N_17572,N_17545);
nand U18108 (N_18108,N_17673,N_17924);
nor U18109 (N_18109,N_17503,N_17932);
nor U18110 (N_18110,N_17656,N_17839);
nor U18111 (N_18111,N_17837,N_17767);
or U18112 (N_18112,N_17531,N_17584);
and U18113 (N_18113,N_17559,N_17936);
nand U18114 (N_18114,N_17818,N_17768);
nor U18115 (N_18115,N_17604,N_17742);
or U18116 (N_18116,N_17896,N_17575);
and U18117 (N_18117,N_17657,N_17760);
xor U18118 (N_18118,N_17978,N_17971);
nand U18119 (N_18119,N_17594,N_17501);
or U18120 (N_18120,N_17905,N_17590);
or U18121 (N_18121,N_17680,N_17783);
xnor U18122 (N_18122,N_17690,N_17514);
or U18123 (N_18123,N_17893,N_17670);
or U18124 (N_18124,N_17547,N_17580);
and U18125 (N_18125,N_17562,N_17902);
nor U18126 (N_18126,N_17852,N_17869);
and U18127 (N_18127,N_17679,N_17822);
and U18128 (N_18128,N_17967,N_17505);
xor U18129 (N_18129,N_17546,N_17965);
xnor U18130 (N_18130,N_17561,N_17651);
or U18131 (N_18131,N_17827,N_17890);
or U18132 (N_18132,N_17860,N_17798);
or U18133 (N_18133,N_17782,N_17512);
xnor U18134 (N_18134,N_17738,N_17764);
or U18135 (N_18135,N_17603,N_17949);
nand U18136 (N_18136,N_17915,N_17606);
nand U18137 (N_18137,N_17627,N_17591);
and U18138 (N_18138,N_17956,N_17773);
and U18139 (N_18139,N_17636,N_17596);
nand U18140 (N_18140,N_17689,N_17788);
xnor U18141 (N_18141,N_17774,N_17740);
and U18142 (N_18142,N_17933,N_17864);
nor U18143 (N_18143,N_17571,N_17659);
and U18144 (N_18144,N_17672,N_17592);
nand U18145 (N_18145,N_17806,N_17834);
nand U18146 (N_18146,N_17777,N_17613);
nand U18147 (N_18147,N_17920,N_17781);
and U18148 (N_18148,N_17787,N_17631);
nand U18149 (N_18149,N_17637,N_17785);
nand U18150 (N_18150,N_17708,N_17928);
nand U18151 (N_18151,N_17586,N_17695);
and U18152 (N_18152,N_17692,N_17962);
xnor U18153 (N_18153,N_17972,N_17939);
and U18154 (N_18154,N_17628,N_17794);
nor U18155 (N_18155,N_17990,N_17617);
or U18156 (N_18156,N_17743,N_17687);
and U18157 (N_18157,N_17886,N_17996);
and U18158 (N_18158,N_17832,N_17885);
xnor U18159 (N_18159,N_17686,N_17713);
and U18160 (N_18160,N_17655,N_17772);
and U18161 (N_18161,N_17513,N_17539);
or U18162 (N_18162,N_17560,N_17829);
nor U18163 (N_18163,N_17941,N_17684);
nor U18164 (N_18164,N_17790,N_17955);
and U18165 (N_18165,N_17835,N_17793);
xor U18166 (N_18166,N_17511,N_17649);
nor U18167 (N_18167,N_17718,N_17814);
or U18168 (N_18168,N_17532,N_17691);
nand U18169 (N_18169,N_17838,N_17707);
or U18170 (N_18170,N_17524,N_17791);
nor U18171 (N_18171,N_17951,N_17600);
xnor U18172 (N_18172,N_17984,N_17929);
nor U18173 (N_18173,N_17694,N_17779);
and U18174 (N_18174,N_17533,N_17652);
and U18175 (N_18175,N_17828,N_17862);
nor U18176 (N_18176,N_17858,N_17986);
nor U18177 (N_18177,N_17960,N_17753);
xor U18178 (N_18178,N_17548,N_17552);
nor U18179 (N_18179,N_17991,N_17755);
nor U18180 (N_18180,N_17700,N_17509);
or U18181 (N_18181,N_17724,N_17723);
or U18182 (N_18182,N_17536,N_17815);
and U18183 (N_18183,N_17671,N_17944);
or U18184 (N_18184,N_17870,N_17678);
and U18185 (N_18185,N_17906,N_17574);
and U18186 (N_18186,N_17749,N_17633);
nor U18187 (N_18187,N_17914,N_17974);
nand U18188 (N_18188,N_17826,N_17702);
nand U18189 (N_18189,N_17911,N_17647);
nand U18190 (N_18190,N_17895,N_17882);
nor U18191 (N_18191,N_17964,N_17795);
and U18192 (N_18192,N_17927,N_17808);
and U18193 (N_18193,N_17525,N_17935);
or U18194 (N_18194,N_17674,N_17853);
nand U18195 (N_18195,N_17585,N_17663);
or U18196 (N_18196,N_17658,N_17712);
and U18197 (N_18197,N_17598,N_17766);
nor U18198 (N_18198,N_17758,N_17607);
or U18199 (N_18199,N_17918,N_17975);
nand U18200 (N_18200,N_17804,N_17987);
or U18201 (N_18201,N_17904,N_17879);
xor U18202 (N_18202,N_17763,N_17952);
xor U18203 (N_18203,N_17980,N_17851);
nor U18204 (N_18204,N_17624,N_17761);
and U18205 (N_18205,N_17517,N_17746);
nand U18206 (N_18206,N_17573,N_17565);
nand U18207 (N_18207,N_17868,N_17567);
nor U18208 (N_18208,N_17880,N_17506);
nor U18209 (N_18209,N_17709,N_17733);
nand U18210 (N_18210,N_17801,N_17626);
or U18211 (N_18211,N_17836,N_17744);
xor U18212 (N_18212,N_17776,N_17595);
nor U18213 (N_18213,N_17719,N_17715);
nand U18214 (N_18214,N_17845,N_17537);
and U18215 (N_18215,N_17730,N_17833);
and U18216 (N_18216,N_17976,N_17646);
or U18217 (N_18217,N_17551,N_17535);
and U18218 (N_18218,N_17910,N_17507);
and U18219 (N_18219,N_17714,N_17745);
and U18220 (N_18220,N_17697,N_17526);
nand U18221 (N_18221,N_17872,N_17661);
nor U18222 (N_18222,N_17605,N_17519);
xnor U18223 (N_18223,N_17881,N_17640);
or U18224 (N_18224,N_17701,N_17716);
and U18225 (N_18225,N_17849,N_17792);
nor U18226 (N_18226,N_17662,N_17618);
and U18227 (N_18227,N_17587,N_17623);
xor U18228 (N_18228,N_17778,N_17579);
or U18229 (N_18229,N_17731,N_17888);
or U18230 (N_18230,N_17688,N_17527);
or U18231 (N_18231,N_17677,N_17528);
xor U18232 (N_18232,N_17721,N_17985);
nor U18233 (N_18233,N_17534,N_17705);
or U18234 (N_18234,N_17970,N_17583);
or U18235 (N_18235,N_17916,N_17820);
nor U18236 (N_18236,N_17564,N_17863);
or U18237 (N_18237,N_17757,N_17830);
nor U18238 (N_18238,N_17555,N_17786);
xor U18239 (N_18239,N_17800,N_17954);
and U18240 (N_18240,N_17722,N_17521);
and U18241 (N_18241,N_17947,N_17703);
or U18242 (N_18242,N_17556,N_17615);
nor U18243 (N_18243,N_17901,N_17937);
nand U18244 (N_18244,N_17878,N_17645);
xnor U18245 (N_18245,N_17685,N_17912);
xor U18246 (N_18246,N_17508,N_17516);
nor U18247 (N_18247,N_17682,N_17696);
nor U18248 (N_18248,N_17884,N_17931);
and U18249 (N_18249,N_17883,N_17717);
xnor U18250 (N_18250,N_17756,N_17897);
nor U18251 (N_18251,N_17952,N_17973);
nor U18252 (N_18252,N_17988,N_17733);
nor U18253 (N_18253,N_17955,N_17960);
xnor U18254 (N_18254,N_17916,N_17834);
xnor U18255 (N_18255,N_17940,N_17983);
xor U18256 (N_18256,N_17527,N_17736);
and U18257 (N_18257,N_17952,N_17592);
nand U18258 (N_18258,N_17524,N_17619);
xnor U18259 (N_18259,N_17728,N_17527);
or U18260 (N_18260,N_17934,N_17602);
or U18261 (N_18261,N_17751,N_17730);
and U18262 (N_18262,N_17627,N_17756);
or U18263 (N_18263,N_17915,N_17785);
nand U18264 (N_18264,N_17876,N_17788);
xor U18265 (N_18265,N_17942,N_17876);
xor U18266 (N_18266,N_17856,N_17528);
nor U18267 (N_18267,N_17839,N_17614);
and U18268 (N_18268,N_17795,N_17576);
xor U18269 (N_18269,N_17903,N_17771);
nor U18270 (N_18270,N_17774,N_17552);
and U18271 (N_18271,N_17986,N_17627);
and U18272 (N_18272,N_17839,N_17770);
xnor U18273 (N_18273,N_17979,N_17779);
and U18274 (N_18274,N_17724,N_17719);
or U18275 (N_18275,N_17874,N_17929);
or U18276 (N_18276,N_17633,N_17556);
nor U18277 (N_18277,N_17749,N_17908);
nand U18278 (N_18278,N_17801,N_17691);
xor U18279 (N_18279,N_17595,N_17693);
nor U18280 (N_18280,N_17722,N_17828);
or U18281 (N_18281,N_17990,N_17945);
nand U18282 (N_18282,N_17679,N_17835);
nand U18283 (N_18283,N_17925,N_17575);
nor U18284 (N_18284,N_17597,N_17708);
and U18285 (N_18285,N_17876,N_17994);
and U18286 (N_18286,N_17837,N_17720);
nand U18287 (N_18287,N_17698,N_17600);
nor U18288 (N_18288,N_17588,N_17592);
and U18289 (N_18289,N_17622,N_17848);
or U18290 (N_18290,N_17953,N_17880);
xnor U18291 (N_18291,N_17735,N_17511);
xnor U18292 (N_18292,N_17619,N_17865);
and U18293 (N_18293,N_17747,N_17537);
nand U18294 (N_18294,N_17513,N_17934);
xor U18295 (N_18295,N_17880,N_17820);
nand U18296 (N_18296,N_17921,N_17557);
nand U18297 (N_18297,N_17669,N_17851);
nand U18298 (N_18298,N_17747,N_17976);
and U18299 (N_18299,N_17729,N_17771);
xnor U18300 (N_18300,N_17984,N_17753);
xnor U18301 (N_18301,N_17504,N_17623);
nand U18302 (N_18302,N_17883,N_17746);
xnor U18303 (N_18303,N_17854,N_17948);
xor U18304 (N_18304,N_17645,N_17684);
nor U18305 (N_18305,N_17527,N_17656);
nor U18306 (N_18306,N_17699,N_17990);
or U18307 (N_18307,N_17979,N_17752);
or U18308 (N_18308,N_17538,N_17751);
nor U18309 (N_18309,N_17689,N_17822);
or U18310 (N_18310,N_17663,N_17635);
xnor U18311 (N_18311,N_17838,N_17560);
nand U18312 (N_18312,N_17880,N_17968);
xnor U18313 (N_18313,N_17763,N_17652);
nor U18314 (N_18314,N_17926,N_17766);
and U18315 (N_18315,N_17515,N_17958);
xnor U18316 (N_18316,N_17884,N_17689);
and U18317 (N_18317,N_17719,N_17646);
or U18318 (N_18318,N_17618,N_17968);
nand U18319 (N_18319,N_17788,N_17795);
xnor U18320 (N_18320,N_17766,N_17579);
and U18321 (N_18321,N_17572,N_17913);
and U18322 (N_18322,N_17983,N_17731);
and U18323 (N_18323,N_17694,N_17775);
or U18324 (N_18324,N_17537,N_17906);
or U18325 (N_18325,N_17771,N_17862);
and U18326 (N_18326,N_17700,N_17699);
or U18327 (N_18327,N_17951,N_17556);
nor U18328 (N_18328,N_17636,N_17527);
nor U18329 (N_18329,N_17749,N_17607);
nor U18330 (N_18330,N_17835,N_17821);
nand U18331 (N_18331,N_17805,N_17936);
nor U18332 (N_18332,N_17862,N_17574);
nand U18333 (N_18333,N_17675,N_17974);
or U18334 (N_18334,N_17681,N_17670);
nor U18335 (N_18335,N_17804,N_17950);
nor U18336 (N_18336,N_17582,N_17637);
nand U18337 (N_18337,N_17658,N_17839);
nor U18338 (N_18338,N_17652,N_17532);
nand U18339 (N_18339,N_17992,N_17663);
or U18340 (N_18340,N_17737,N_17655);
nand U18341 (N_18341,N_17571,N_17790);
nand U18342 (N_18342,N_17510,N_17524);
and U18343 (N_18343,N_17673,N_17747);
xnor U18344 (N_18344,N_17688,N_17514);
or U18345 (N_18345,N_17838,N_17730);
nand U18346 (N_18346,N_17519,N_17741);
and U18347 (N_18347,N_17944,N_17971);
or U18348 (N_18348,N_17649,N_17967);
nand U18349 (N_18349,N_17922,N_17695);
and U18350 (N_18350,N_17766,N_17767);
nand U18351 (N_18351,N_17756,N_17548);
nor U18352 (N_18352,N_17514,N_17852);
xnor U18353 (N_18353,N_17743,N_17634);
nand U18354 (N_18354,N_17546,N_17751);
xnor U18355 (N_18355,N_17878,N_17750);
xnor U18356 (N_18356,N_17547,N_17625);
or U18357 (N_18357,N_17572,N_17685);
xnor U18358 (N_18358,N_17932,N_17929);
xor U18359 (N_18359,N_17871,N_17824);
nand U18360 (N_18360,N_17797,N_17878);
xnor U18361 (N_18361,N_17646,N_17886);
nand U18362 (N_18362,N_17760,N_17510);
and U18363 (N_18363,N_17903,N_17767);
or U18364 (N_18364,N_17845,N_17789);
nor U18365 (N_18365,N_17930,N_17520);
and U18366 (N_18366,N_17854,N_17502);
and U18367 (N_18367,N_17689,N_17514);
nor U18368 (N_18368,N_17599,N_17866);
xor U18369 (N_18369,N_17535,N_17911);
nor U18370 (N_18370,N_17960,N_17630);
nor U18371 (N_18371,N_17827,N_17657);
xnor U18372 (N_18372,N_17853,N_17549);
or U18373 (N_18373,N_17532,N_17620);
or U18374 (N_18374,N_17563,N_17741);
nand U18375 (N_18375,N_17611,N_17528);
nand U18376 (N_18376,N_17584,N_17603);
xor U18377 (N_18377,N_17585,N_17771);
nand U18378 (N_18378,N_17906,N_17568);
nor U18379 (N_18379,N_17640,N_17966);
xor U18380 (N_18380,N_17706,N_17957);
or U18381 (N_18381,N_17708,N_17546);
or U18382 (N_18382,N_17524,N_17978);
and U18383 (N_18383,N_17746,N_17693);
xnor U18384 (N_18384,N_17931,N_17833);
or U18385 (N_18385,N_17884,N_17703);
nor U18386 (N_18386,N_17828,N_17532);
and U18387 (N_18387,N_17902,N_17647);
nor U18388 (N_18388,N_17562,N_17555);
nand U18389 (N_18389,N_17997,N_17782);
nor U18390 (N_18390,N_17606,N_17645);
or U18391 (N_18391,N_17586,N_17507);
and U18392 (N_18392,N_17726,N_17721);
xor U18393 (N_18393,N_17935,N_17899);
nor U18394 (N_18394,N_17856,N_17890);
xor U18395 (N_18395,N_17795,N_17782);
xor U18396 (N_18396,N_17808,N_17975);
nand U18397 (N_18397,N_17881,N_17600);
or U18398 (N_18398,N_17918,N_17939);
or U18399 (N_18399,N_17534,N_17709);
nor U18400 (N_18400,N_17720,N_17672);
and U18401 (N_18401,N_17515,N_17998);
nand U18402 (N_18402,N_17807,N_17968);
nand U18403 (N_18403,N_17773,N_17822);
and U18404 (N_18404,N_17664,N_17689);
and U18405 (N_18405,N_17927,N_17705);
or U18406 (N_18406,N_17698,N_17647);
xor U18407 (N_18407,N_17716,N_17967);
nor U18408 (N_18408,N_17527,N_17977);
or U18409 (N_18409,N_17658,N_17552);
xnor U18410 (N_18410,N_17740,N_17629);
or U18411 (N_18411,N_17541,N_17557);
nor U18412 (N_18412,N_17532,N_17862);
nor U18413 (N_18413,N_17857,N_17992);
nand U18414 (N_18414,N_17822,N_17687);
and U18415 (N_18415,N_17504,N_17894);
nor U18416 (N_18416,N_17797,N_17894);
nor U18417 (N_18417,N_17606,N_17506);
and U18418 (N_18418,N_17658,N_17661);
nand U18419 (N_18419,N_17945,N_17649);
nand U18420 (N_18420,N_17535,N_17778);
or U18421 (N_18421,N_17862,N_17685);
and U18422 (N_18422,N_17582,N_17813);
xnor U18423 (N_18423,N_17640,N_17526);
or U18424 (N_18424,N_17860,N_17724);
xnor U18425 (N_18425,N_17777,N_17884);
and U18426 (N_18426,N_17877,N_17860);
and U18427 (N_18427,N_17631,N_17869);
nand U18428 (N_18428,N_17774,N_17558);
xor U18429 (N_18429,N_17521,N_17958);
nand U18430 (N_18430,N_17574,N_17814);
xor U18431 (N_18431,N_17673,N_17614);
nand U18432 (N_18432,N_17947,N_17841);
nor U18433 (N_18433,N_17586,N_17520);
and U18434 (N_18434,N_17819,N_17581);
nor U18435 (N_18435,N_17697,N_17708);
or U18436 (N_18436,N_17550,N_17729);
nand U18437 (N_18437,N_17524,N_17859);
nand U18438 (N_18438,N_17549,N_17890);
xor U18439 (N_18439,N_17742,N_17992);
and U18440 (N_18440,N_17652,N_17576);
nand U18441 (N_18441,N_17756,N_17672);
nand U18442 (N_18442,N_17696,N_17949);
xor U18443 (N_18443,N_17856,N_17602);
nand U18444 (N_18444,N_17694,N_17525);
and U18445 (N_18445,N_17885,N_17664);
or U18446 (N_18446,N_17971,N_17902);
or U18447 (N_18447,N_17859,N_17661);
nor U18448 (N_18448,N_17965,N_17771);
nand U18449 (N_18449,N_17833,N_17746);
nor U18450 (N_18450,N_17602,N_17527);
or U18451 (N_18451,N_17593,N_17644);
and U18452 (N_18452,N_17522,N_17776);
xor U18453 (N_18453,N_17853,N_17705);
xor U18454 (N_18454,N_17819,N_17806);
xor U18455 (N_18455,N_17727,N_17562);
and U18456 (N_18456,N_17840,N_17588);
nand U18457 (N_18457,N_17517,N_17956);
nand U18458 (N_18458,N_17906,N_17580);
xnor U18459 (N_18459,N_17630,N_17823);
nor U18460 (N_18460,N_17747,N_17756);
xnor U18461 (N_18461,N_17551,N_17874);
nand U18462 (N_18462,N_17833,N_17547);
or U18463 (N_18463,N_17829,N_17901);
and U18464 (N_18464,N_17749,N_17587);
xnor U18465 (N_18465,N_17686,N_17716);
and U18466 (N_18466,N_17720,N_17627);
and U18467 (N_18467,N_17984,N_17875);
nand U18468 (N_18468,N_17654,N_17737);
nor U18469 (N_18469,N_17645,N_17881);
and U18470 (N_18470,N_17882,N_17762);
nand U18471 (N_18471,N_17703,N_17970);
and U18472 (N_18472,N_17908,N_17888);
or U18473 (N_18473,N_17550,N_17925);
xnor U18474 (N_18474,N_17537,N_17700);
xor U18475 (N_18475,N_17650,N_17507);
nor U18476 (N_18476,N_17897,N_17993);
and U18477 (N_18477,N_17565,N_17767);
or U18478 (N_18478,N_17921,N_17531);
nand U18479 (N_18479,N_17943,N_17859);
and U18480 (N_18480,N_17922,N_17581);
nor U18481 (N_18481,N_17540,N_17676);
and U18482 (N_18482,N_17829,N_17723);
xnor U18483 (N_18483,N_17722,N_17896);
or U18484 (N_18484,N_17983,N_17784);
nand U18485 (N_18485,N_17733,N_17792);
and U18486 (N_18486,N_17500,N_17546);
nand U18487 (N_18487,N_17532,N_17953);
xnor U18488 (N_18488,N_17626,N_17568);
xnor U18489 (N_18489,N_17986,N_17637);
or U18490 (N_18490,N_17712,N_17962);
nand U18491 (N_18491,N_17617,N_17915);
nor U18492 (N_18492,N_17964,N_17946);
xnor U18493 (N_18493,N_17693,N_17562);
xnor U18494 (N_18494,N_17625,N_17846);
nor U18495 (N_18495,N_17686,N_17814);
nor U18496 (N_18496,N_17751,N_17821);
and U18497 (N_18497,N_17570,N_17752);
nand U18498 (N_18498,N_17563,N_17525);
nor U18499 (N_18499,N_17648,N_17895);
nand U18500 (N_18500,N_18237,N_18490);
nand U18501 (N_18501,N_18431,N_18119);
nor U18502 (N_18502,N_18198,N_18308);
nand U18503 (N_18503,N_18451,N_18444);
nand U18504 (N_18504,N_18225,N_18343);
and U18505 (N_18505,N_18337,N_18371);
nor U18506 (N_18506,N_18322,N_18229);
nor U18507 (N_18507,N_18392,N_18019);
nor U18508 (N_18508,N_18064,N_18273);
xnor U18509 (N_18509,N_18005,N_18338);
and U18510 (N_18510,N_18321,N_18289);
xor U18511 (N_18511,N_18235,N_18405);
and U18512 (N_18512,N_18452,N_18004);
xnor U18513 (N_18513,N_18102,N_18044);
and U18514 (N_18514,N_18200,N_18447);
nand U18515 (N_18515,N_18034,N_18189);
or U18516 (N_18516,N_18012,N_18038);
and U18517 (N_18517,N_18448,N_18382);
nand U18518 (N_18518,N_18181,N_18021);
nor U18519 (N_18519,N_18245,N_18194);
or U18520 (N_18520,N_18336,N_18088);
nor U18521 (N_18521,N_18416,N_18261);
nand U18522 (N_18522,N_18456,N_18369);
xnor U18523 (N_18523,N_18109,N_18412);
nand U18524 (N_18524,N_18413,N_18330);
nand U18525 (N_18525,N_18182,N_18464);
and U18526 (N_18526,N_18140,N_18354);
and U18527 (N_18527,N_18108,N_18049);
nand U18528 (N_18528,N_18065,N_18357);
and U18529 (N_18529,N_18305,N_18248);
nand U18530 (N_18530,N_18139,N_18481);
nor U18531 (N_18531,N_18009,N_18161);
xor U18532 (N_18532,N_18095,N_18016);
or U18533 (N_18533,N_18487,N_18185);
nor U18534 (N_18534,N_18436,N_18247);
nor U18535 (N_18535,N_18014,N_18302);
or U18536 (N_18536,N_18318,N_18278);
xor U18537 (N_18537,N_18097,N_18409);
and U18538 (N_18538,N_18350,N_18145);
nor U18539 (N_18539,N_18141,N_18192);
or U18540 (N_18540,N_18489,N_18255);
xnor U18541 (N_18541,N_18491,N_18332);
nand U18542 (N_18542,N_18231,N_18495);
nor U18543 (N_18543,N_18290,N_18121);
nor U18544 (N_18544,N_18258,N_18018);
nand U18545 (N_18545,N_18297,N_18317);
and U18546 (N_18546,N_18351,N_18226);
nand U18547 (N_18547,N_18313,N_18461);
and U18548 (N_18548,N_18328,N_18374);
nand U18549 (N_18549,N_18144,N_18050);
and U18550 (N_18550,N_18202,N_18315);
nor U18551 (N_18551,N_18234,N_18474);
and U18552 (N_18552,N_18363,N_18284);
or U18553 (N_18553,N_18469,N_18041);
or U18554 (N_18554,N_18162,N_18341);
and U18555 (N_18555,N_18285,N_18378);
nor U18556 (N_18556,N_18213,N_18372);
and U18557 (N_18557,N_18045,N_18152);
xnor U18558 (N_18558,N_18184,N_18172);
nand U18559 (N_18559,N_18439,N_18087);
nand U18560 (N_18560,N_18477,N_18023);
nor U18561 (N_18561,N_18218,N_18327);
nand U18562 (N_18562,N_18134,N_18274);
or U18563 (N_18563,N_18260,N_18057);
and U18564 (N_18564,N_18206,N_18124);
nor U18565 (N_18565,N_18101,N_18026);
and U18566 (N_18566,N_18320,N_18323);
xor U18567 (N_18567,N_18298,N_18210);
xnor U18568 (N_18568,N_18475,N_18453);
nand U18569 (N_18569,N_18483,N_18053);
xor U18570 (N_18570,N_18003,N_18471);
nand U18571 (N_18571,N_18190,N_18393);
xnor U18572 (N_18572,N_18163,N_18132);
and U18573 (N_18573,N_18485,N_18345);
nor U18574 (N_18574,N_18060,N_18061);
or U18575 (N_18575,N_18007,N_18178);
nand U18576 (N_18576,N_18253,N_18227);
nor U18577 (N_18577,N_18107,N_18277);
nor U18578 (N_18578,N_18169,N_18187);
xor U18579 (N_18579,N_18484,N_18129);
xor U18580 (N_18580,N_18280,N_18271);
nor U18581 (N_18581,N_18286,N_18265);
nor U18582 (N_18582,N_18083,N_18070);
nor U18583 (N_18583,N_18063,N_18168);
or U18584 (N_18584,N_18348,N_18389);
and U18585 (N_18585,N_18000,N_18296);
nand U18586 (N_18586,N_18333,N_18457);
xnor U18587 (N_18587,N_18092,N_18171);
and U18588 (N_18588,N_18463,N_18113);
or U18589 (N_18589,N_18243,N_18156);
or U18590 (N_18590,N_18052,N_18074);
or U18591 (N_18591,N_18137,N_18306);
and U18592 (N_18592,N_18496,N_18059);
nand U18593 (N_18593,N_18266,N_18268);
nand U18594 (N_18594,N_18086,N_18035);
nor U18595 (N_18595,N_18391,N_18138);
xor U18596 (N_18596,N_18498,N_18460);
nor U18597 (N_18597,N_18326,N_18440);
xnor U18598 (N_18598,N_18173,N_18186);
or U18599 (N_18599,N_18397,N_18224);
and U18600 (N_18600,N_18404,N_18370);
or U18601 (N_18601,N_18269,N_18188);
or U18602 (N_18602,N_18179,N_18478);
nand U18603 (N_18603,N_18426,N_18155);
and U18604 (N_18604,N_18311,N_18325);
or U18605 (N_18605,N_18380,N_18017);
xnor U18606 (N_18606,N_18242,N_18233);
xor U18607 (N_18607,N_18028,N_18191);
xnor U18608 (N_18608,N_18068,N_18470);
nor U18609 (N_18609,N_18090,N_18013);
nor U18610 (N_18610,N_18153,N_18100);
or U18611 (N_18611,N_18089,N_18419);
or U18612 (N_18612,N_18459,N_18301);
nor U18613 (N_18613,N_18054,N_18116);
or U18614 (N_18614,N_18223,N_18197);
and U18615 (N_18615,N_18373,N_18408);
xnor U18616 (N_18616,N_18443,N_18069);
nor U18617 (N_18617,N_18340,N_18428);
nand U18618 (N_18618,N_18263,N_18388);
nand U18619 (N_18619,N_18473,N_18098);
nor U18620 (N_18620,N_18251,N_18445);
or U18621 (N_18621,N_18011,N_18072);
and U18622 (N_18622,N_18025,N_18376);
nor U18623 (N_18623,N_18434,N_18259);
nor U18624 (N_18624,N_18055,N_18379);
nand U18625 (N_18625,N_18300,N_18293);
nand U18626 (N_18626,N_18110,N_18492);
xnor U18627 (N_18627,N_18177,N_18292);
xnor U18628 (N_18628,N_18022,N_18236);
xnor U18629 (N_18629,N_18240,N_18291);
xnor U18630 (N_18630,N_18486,N_18176);
or U18631 (N_18631,N_18066,N_18433);
and U18632 (N_18632,N_18353,N_18203);
and U18633 (N_18633,N_18062,N_18359);
xor U18634 (N_18634,N_18067,N_18476);
nor U18635 (N_18635,N_18335,N_18358);
xor U18636 (N_18636,N_18073,N_18159);
and U18637 (N_18637,N_18395,N_18215);
xnor U18638 (N_18638,N_18417,N_18400);
nor U18639 (N_18639,N_18123,N_18015);
nand U18640 (N_18640,N_18199,N_18114);
nand U18641 (N_18641,N_18377,N_18221);
and U18642 (N_18642,N_18076,N_18310);
and U18643 (N_18643,N_18466,N_18331);
xor U18644 (N_18644,N_18410,N_18080);
or U18645 (N_18645,N_18275,N_18314);
and U18646 (N_18646,N_18126,N_18180);
or U18647 (N_18647,N_18104,N_18299);
or U18648 (N_18648,N_18122,N_18128);
nor U18649 (N_18649,N_18030,N_18105);
nor U18650 (N_18650,N_18027,N_18112);
nor U18651 (N_18651,N_18307,N_18216);
nor U18652 (N_18652,N_18131,N_18304);
xor U18653 (N_18653,N_18324,N_18430);
nor U18654 (N_18654,N_18394,N_18099);
xor U18655 (N_18655,N_18143,N_18127);
nor U18656 (N_18656,N_18056,N_18250);
nor U18657 (N_18657,N_18407,N_18406);
nand U18658 (N_18658,N_18033,N_18111);
xor U18659 (N_18659,N_18157,N_18077);
or U18660 (N_18660,N_18402,N_18149);
nand U18661 (N_18661,N_18091,N_18207);
or U18662 (N_18662,N_18421,N_18232);
or U18663 (N_18663,N_18272,N_18195);
or U18664 (N_18664,N_18120,N_18096);
nor U18665 (N_18665,N_18058,N_18465);
xnor U18666 (N_18666,N_18165,N_18219);
nor U18667 (N_18667,N_18267,N_18287);
and U18668 (N_18668,N_18422,N_18047);
nor U18669 (N_18669,N_18252,N_18093);
xor U18670 (N_18670,N_18349,N_18454);
or U18671 (N_18671,N_18442,N_18346);
xnor U18672 (N_18672,N_18164,N_18036);
and U18673 (N_18673,N_18010,N_18174);
and U18674 (N_18674,N_18201,N_18204);
nand U18675 (N_18675,N_18365,N_18130);
xnor U18676 (N_18676,N_18002,N_18048);
nand U18677 (N_18677,N_18295,N_18029);
xnor U18678 (N_18678,N_18220,N_18079);
or U18679 (N_18679,N_18387,N_18118);
or U18680 (N_18680,N_18270,N_18472);
and U18681 (N_18681,N_18228,N_18467);
or U18682 (N_18682,N_18386,N_18212);
xor U18683 (N_18683,N_18368,N_18264);
xor U18684 (N_18684,N_18411,N_18241);
xnor U18685 (N_18685,N_18425,N_18039);
and U18686 (N_18686,N_18214,N_18024);
nand U18687 (N_18687,N_18367,N_18479);
or U18688 (N_18688,N_18071,N_18106);
xnor U18689 (N_18689,N_18020,N_18344);
nand U18690 (N_18690,N_18366,N_18037);
xor U18691 (N_18691,N_18384,N_18441);
or U18692 (N_18692,N_18329,N_18257);
and U18693 (N_18693,N_18450,N_18493);
xnor U18694 (N_18694,N_18103,N_18084);
nand U18695 (N_18695,N_18424,N_18455);
nand U18696 (N_18696,N_18146,N_18167);
xor U18697 (N_18697,N_18468,N_18362);
xor U18698 (N_18698,N_18051,N_18316);
nand U18699 (N_18699,N_18193,N_18446);
nand U18700 (N_18700,N_18148,N_18282);
nand U18701 (N_18701,N_18081,N_18211);
nor U18702 (N_18702,N_18082,N_18438);
nor U18703 (N_18703,N_18488,N_18166);
nor U18704 (N_18704,N_18401,N_18078);
nor U18705 (N_18705,N_18383,N_18217);
and U18706 (N_18706,N_18175,N_18319);
and U18707 (N_18707,N_18254,N_18435);
or U18708 (N_18708,N_18244,N_18281);
xnor U18709 (N_18709,N_18352,N_18334);
and U18710 (N_18710,N_18385,N_18239);
xor U18711 (N_18711,N_18437,N_18117);
or U18712 (N_18712,N_18427,N_18482);
and U18713 (N_18713,N_18339,N_18356);
nor U18714 (N_18714,N_18283,N_18494);
nand U18715 (N_18715,N_18480,N_18396);
xor U18716 (N_18716,N_18256,N_18381);
and U18717 (N_18717,N_18364,N_18135);
nand U18718 (N_18718,N_18403,N_18458);
and U18719 (N_18719,N_18085,N_18208);
and U18720 (N_18720,N_18133,N_18040);
nand U18721 (N_18721,N_18249,N_18042);
nand U18722 (N_18722,N_18312,N_18262);
nor U18723 (N_18723,N_18399,N_18046);
and U18724 (N_18724,N_18375,N_18418);
xnor U18725 (N_18725,N_18230,N_18288);
xor U18726 (N_18726,N_18361,N_18449);
nor U18727 (N_18727,N_18158,N_18294);
nand U18728 (N_18728,N_18355,N_18420);
nor U18729 (N_18729,N_18390,N_18183);
nand U18730 (N_18730,N_18423,N_18136);
or U18731 (N_18731,N_18160,N_18032);
nor U18732 (N_18732,N_18222,N_18147);
nand U18733 (N_18733,N_18415,N_18043);
xnor U18734 (N_18734,N_18309,N_18196);
xor U18735 (N_18735,N_18205,N_18347);
and U18736 (N_18736,N_18150,N_18125);
and U18737 (N_18737,N_18462,N_18154);
and U18738 (N_18738,N_18432,N_18303);
or U18739 (N_18739,N_18414,N_18170);
nor U18740 (N_18740,N_18429,N_18497);
xor U18741 (N_18741,N_18142,N_18360);
nor U18742 (N_18742,N_18209,N_18238);
or U18743 (N_18743,N_18001,N_18115);
nand U18744 (N_18744,N_18276,N_18075);
nand U18745 (N_18745,N_18342,N_18246);
nor U18746 (N_18746,N_18279,N_18398);
nor U18747 (N_18747,N_18006,N_18094);
or U18748 (N_18748,N_18008,N_18031);
nor U18749 (N_18749,N_18151,N_18499);
or U18750 (N_18750,N_18257,N_18484);
and U18751 (N_18751,N_18290,N_18336);
nor U18752 (N_18752,N_18433,N_18469);
nor U18753 (N_18753,N_18341,N_18426);
xor U18754 (N_18754,N_18356,N_18004);
nand U18755 (N_18755,N_18305,N_18234);
xor U18756 (N_18756,N_18155,N_18251);
xor U18757 (N_18757,N_18015,N_18045);
and U18758 (N_18758,N_18036,N_18167);
nor U18759 (N_18759,N_18221,N_18129);
or U18760 (N_18760,N_18155,N_18196);
nand U18761 (N_18761,N_18104,N_18429);
xor U18762 (N_18762,N_18161,N_18008);
and U18763 (N_18763,N_18460,N_18165);
xor U18764 (N_18764,N_18076,N_18279);
or U18765 (N_18765,N_18228,N_18194);
or U18766 (N_18766,N_18263,N_18094);
and U18767 (N_18767,N_18184,N_18205);
or U18768 (N_18768,N_18393,N_18289);
nand U18769 (N_18769,N_18082,N_18256);
and U18770 (N_18770,N_18303,N_18205);
nor U18771 (N_18771,N_18295,N_18007);
and U18772 (N_18772,N_18021,N_18018);
nand U18773 (N_18773,N_18386,N_18322);
xnor U18774 (N_18774,N_18058,N_18332);
nand U18775 (N_18775,N_18064,N_18380);
and U18776 (N_18776,N_18399,N_18121);
nand U18777 (N_18777,N_18273,N_18302);
nand U18778 (N_18778,N_18247,N_18352);
and U18779 (N_18779,N_18203,N_18105);
and U18780 (N_18780,N_18332,N_18255);
and U18781 (N_18781,N_18449,N_18350);
nand U18782 (N_18782,N_18429,N_18138);
xnor U18783 (N_18783,N_18168,N_18302);
xor U18784 (N_18784,N_18412,N_18275);
nor U18785 (N_18785,N_18319,N_18017);
nor U18786 (N_18786,N_18296,N_18351);
and U18787 (N_18787,N_18377,N_18099);
xnor U18788 (N_18788,N_18346,N_18145);
nand U18789 (N_18789,N_18458,N_18045);
xnor U18790 (N_18790,N_18169,N_18355);
and U18791 (N_18791,N_18478,N_18163);
nand U18792 (N_18792,N_18332,N_18463);
nor U18793 (N_18793,N_18389,N_18360);
nor U18794 (N_18794,N_18151,N_18289);
or U18795 (N_18795,N_18465,N_18008);
and U18796 (N_18796,N_18456,N_18160);
and U18797 (N_18797,N_18214,N_18291);
xor U18798 (N_18798,N_18009,N_18457);
and U18799 (N_18799,N_18409,N_18095);
nand U18800 (N_18800,N_18135,N_18165);
xnor U18801 (N_18801,N_18426,N_18374);
xnor U18802 (N_18802,N_18214,N_18183);
and U18803 (N_18803,N_18463,N_18080);
xnor U18804 (N_18804,N_18114,N_18150);
or U18805 (N_18805,N_18291,N_18135);
or U18806 (N_18806,N_18391,N_18290);
nand U18807 (N_18807,N_18446,N_18189);
and U18808 (N_18808,N_18140,N_18385);
and U18809 (N_18809,N_18239,N_18211);
or U18810 (N_18810,N_18203,N_18004);
and U18811 (N_18811,N_18282,N_18194);
and U18812 (N_18812,N_18218,N_18234);
nor U18813 (N_18813,N_18456,N_18146);
and U18814 (N_18814,N_18387,N_18478);
and U18815 (N_18815,N_18392,N_18043);
nand U18816 (N_18816,N_18445,N_18442);
or U18817 (N_18817,N_18137,N_18468);
nand U18818 (N_18818,N_18257,N_18212);
nand U18819 (N_18819,N_18124,N_18035);
nand U18820 (N_18820,N_18285,N_18124);
nand U18821 (N_18821,N_18087,N_18285);
and U18822 (N_18822,N_18499,N_18414);
nor U18823 (N_18823,N_18302,N_18158);
and U18824 (N_18824,N_18133,N_18465);
nand U18825 (N_18825,N_18090,N_18348);
or U18826 (N_18826,N_18436,N_18242);
nor U18827 (N_18827,N_18223,N_18290);
and U18828 (N_18828,N_18361,N_18282);
and U18829 (N_18829,N_18424,N_18304);
or U18830 (N_18830,N_18132,N_18223);
nand U18831 (N_18831,N_18280,N_18458);
xor U18832 (N_18832,N_18207,N_18441);
and U18833 (N_18833,N_18046,N_18364);
xor U18834 (N_18834,N_18083,N_18490);
nand U18835 (N_18835,N_18236,N_18086);
or U18836 (N_18836,N_18242,N_18134);
xnor U18837 (N_18837,N_18287,N_18233);
nor U18838 (N_18838,N_18078,N_18133);
and U18839 (N_18839,N_18476,N_18447);
xnor U18840 (N_18840,N_18475,N_18096);
nor U18841 (N_18841,N_18170,N_18268);
nor U18842 (N_18842,N_18256,N_18361);
and U18843 (N_18843,N_18338,N_18059);
or U18844 (N_18844,N_18114,N_18090);
nand U18845 (N_18845,N_18363,N_18092);
or U18846 (N_18846,N_18304,N_18323);
or U18847 (N_18847,N_18111,N_18005);
and U18848 (N_18848,N_18007,N_18000);
nor U18849 (N_18849,N_18249,N_18013);
nand U18850 (N_18850,N_18470,N_18309);
and U18851 (N_18851,N_18216,N_18303);
nor U18852 (N_18852,N_18210,N_18194);
and U18853 (N_18853,N_18486,N_18032);
nand U18854 (N_18854,N_18430,N_18283);
nand U18855 (N_18855,N_18432,N_18149);
xnor U18856 (N_18856,N_18368,N_18350);
and U18857 (N_18857,N_18429,N_18309);
or U18858 (N_18858,N_18318,N_18047);
nor U18859 (N_18859,N_18228,N_18117);
and U18860 (N_18860,N_18070,N_18414);
and U18861 (N_18861,N_18372,N_18105);
xnor U18862 (N_18862,N_18482,N_18135);
nand U18863 (N_18863,N_18045,N_18277);
nand U18864 (N_18864,N_18342,N_18251);
or U18865 (N_18865,N_18397,N_18019);
xnor U18866 (N_18866,N_18213,N_18352);
nand U18867 (N_18867,N_18112,N_18201);
nor U18868 (N_18868,N_18196,N_18207);
nand U18869 (N_18869,N_18484,N_18335);
and U18870 (N_18870,N_18257,N_18292);
nand U18871 (N_18871,N_18294,N_18153);
xor U18872 (N_18872,N_18384,N_18108);
nor U18873 (N_18873,N_18096,N_18372);
xor U18874 (N_18874,N_18166,N_18308);
or U18875 (N_18875,N_18197,N_18337);
nand U18876 (N_18876,N_18348,N_18192);
xnor U18877 (N_18877,N_18094,N_18372);
nor U18878 (N_18878,N_18494,N_18416);
nor U18879 (N_18879,N_18020,N_18229);
xor U18880 (N_18880,N_18341,N_18183);
and U18881 (N_18881,N_18117,N_18111);
xnor U18882 (N_18882,N_18056,N_18241);
or U18883 (N_18883,N_18361,N_18220);
xor U18884 (N_18884,N_18407,N_18193);
and U18885 (N_18885,N_18319,N_18145);
xnor U18886 (N_18886,N_18104,N_18001);
xnor U18887 (N_18887,N_18288,N_18068);
and U18888 (N_18888,N_18009,N_18382);
or U18889 (N_18889,N_18402,N_18342);
and U18890 (N_18890,N_18240,N_18081);
xnor U18891 (N_18891,N_18487,N_18404);
xor U18892 (N_18892,N_18176,N_18493);
and U18893 (N_18893,N_18292,N_18416);
nor U18894 (N_18894,N_18275,N_18045);
xor U18895 (N_18895,N_18325,N_18083);
nor U18896 (N_18896,N_18260,N_18233);
nor U18897 (N_18897,N_18411,N_18413);
xor U18898 (N_18898,N_18492,N_18227);
xor U18899 (N_18899,N_18218,N_18045);
xnor U18900 (N_18900,N_18113,N_18334);
or U18901 (N_18901,N_18458,N_18106);
or U18902 (N_18902,N_18097,N_18116);
nand U18903 (N_18903,N_18122,N_18131);
nand U18904 (N_18904,N_18203,N_18346);
and U18905 (N_18905,N_18379,N_18098);
or U18906 (N_18906,N_18429,N_18310);
xor U18907 (N_18907,N_18091,N_18039);
nand U18908 (N_18908,N_18274,N_18366);
nor U18909 (N_18909,N_18350,N_18107);
xnor U18910 (N_18910,N_18446,N_18439);
or U18911 (N_18911,N_18028,N_18409);
nor U18912 (N_18912,N_18476,N_18008);
xnor U18913 (N_18913,N_18048,N_18355);
nor U18914 (N_18914,N_18040,N_18268);
or U18915 (N_18915,N_18294,N_18473);
xor U18916 (N_18916,N_18460,N_18274);
nor U18917 (N_18917,N_18307,N_18050);
and U18918 (N_18918,N_18451,N_18058);
nand U18919 (N_18919,N_18088,N_18355);
xor U18920 (N_18920,N_18085,N_18393);
and U18921 (N_18921,N_18017,N_18420);
nor U18922 (N_18922,N_18112,N_18069);
and U18923 (N_18923,N_18419,N_18288);
or U18924 (N_18924,N_18162,N_18325);
and U18925 (N_18925,N_18324,N_18493);
and U18926 (N_18926,N_18433,N_18435);
nand U18927 (N_18927,N_18396,N_18030);
or U18928 (N_18928,N_18493,N_18414);
nand U18929 (N_18929,N_18461,N_18071);
nor U18930 (N_18930,N_18457,N_18080);
xor U18931 (N_18931,N_18072,N_18356);
xnor U18932 (N_18932,N_18172,N_18119);
xnor U18933 (N_18933,N_18220,N_18386);
or U18934 (N_18934,N_18066,N_18431);
nor U18935 (N_18935,N_18303,N_18029);
nor U18936 (N_18936,N_18348,N_18405);
and U18937 (N_18937,N_18396,N_18131);
nor U18938 (N_18938,N_18476,N_18261);
and U18939 (N_18939,N_18347,N_18074);
nand U18940 (N_18940,N_18100,N_18276);
nor U18941 (N_18941,N_18488,N_18037);
xor U18942 (N_18942,N_18426,N_18278);
nand U18943 (N_18943,N_18114,N_18161);
nor U18944 (N_18944,N_18139,N_18476);
nor U18945 (N_18945,N_18405,N_18464);
nor U18946 (N_18946,N_18255,N_18306);
and U18947 (N_18947,N_18209,N_18433);
or U18948 (N_18948,N_18194,N_18376);
nand U18949 (N_18949,N_18287,N_18262);
xnor U18950 (N_18950,N_18293,N_18375);
or U18951 (N_18951,N_18135,N_18417);
and U18952 (N_18952,N_18002,N_18127);
and U18953 (N_18953,N_18075,N_18100);
nor U18954 (N_18954,N_18245,N_18498);
xnor U18955 (N_18955,N_18126,N_18415);
nand U18956 (N_18956,N_18391,N_18110);
and U18957 (N_18957,N_18211,N_18364);
and U18958 (N_18958,N_18397,N_18060);
nor U18959 (N_18959,N_18293,N_18382);
and U18960 (N_18960,N_18069,N_18166);
nand U18961 (N_18961,N_18464,N_18371);
and U18962 (N_18962,N_18368,N_18241);
nor U18963 (N_18963,N_18097,N_18126);
nand U18964 (N_18964,N_18094,N_18127);
xnor U18965 (N_18965,N_18200,N_18179);
and U18966 (N_18966,N_18387,N_18127);
nand U18967 (N_18967,N_18151,N_18309);
and U18968 (N_18968,N_18379,N_18456);
xnor U18969 (N_18969,N_18264,N_18346);
or U18970 (N_18970,N_18445,N_18001);
and U18971 (N_18971,N_18176,N_18041);
or U18972 (N_18972,N_18057,N_18420);
xnor U18973 (N_18973,N_18191,N_18097);
or U18974 (N_18974,N_18280,N_18338);
or U18975 (N_18975,N_18130,N_18406);
nand U18976 (N_18976,N_18235,N_18201);
and U18977 (N_18977,N_18094,N_18441);
nand U18978 (N_18978,N_18228,N_18242);
nand U18979 (N_18979,N_18383,N_18094);
nor U18980 (N_18980,N_18112,N_18071);
nor U18981 (N_18981,N_18220,N_18311);
and U18982 (N_18982,N_18323,N_18486);
nor U18983 (N_18983,N_18492,N_18459);
nor U18984 (N_18984,N_18085,N_18185);
xor U18985 (N_18985,N_18086,N_18246);
nor U18986 (N_18986,N_18192,N_18108);
nand U18987 (N_18987,N_18049,N_18350);
or U18988 (N_18988,N_18341,N_18179);
xor U18989 (N_18989,N_18282,N_18000);
xnor U18990 (N_18990,N_18043,N_18130);
or U18991 (N_18991,N_18267,N_18431);
and U18992 (N_18992,N_18138,N_18021);
and U18993 (N_18993,N_18458,N_18372);
and U18994 (N_18994,N_18042,N_18227);
and U18995 (N_18995,N_18195,N_18388);
or U18996 (N_18996,N_18487,N_18118);
nand U18997 (N_18997,N_18419,N_18055);
nand U18998 (N_18998,N_18436,N_18354);
and U18999 (N_18999,N_18376,N_18288);
nor U19000 (N_19000,N_18570,N_18903);
and U19001 (N_19001,N_18658,N_18676);
or U19002 (N_19002,N_18759,N_18739);
and U19003 (N_19003,N_18673,N_18945);
nand U19004 (N_19004,N_18687,N_18718);
or U19005 (N_19005,N_18794,N_18523);
nand U19006 (N_19006,N_18603,N_18848);
nor U19007 (N_19007,N_18926,N_18619);
nor U19008 (N_19008,N_18934,N_18521);
nand U19009 (N_19009,N_18669,N_18777);
nor U19010 (N_19010,N_18768,N_18968);
xnor U19011 (N_19011,N_18646,N_18559);
nor U19012 (N_19012,N_18510,N_18636);
nor U19013 (N_19013,N_18839,N_18917);
xnor U19014 (N_19014,N_18890,N_18784);
or U19015 (N_19015,N_18617,N_18858);
nand U19016 (N_19016,N_18554,N_18626);
nand U19017 (N_19017,N_18754,N_18850);
or U19018 (N_19018,N_18702,N_18597);
nor U19019 (N_19019,N_18745,N_18614);
or U19020 (N_19020,N_18908,N_18911);
and U19021 (N_19021,N_18827,N_18751);
or U19022 (N_19022,N_18688,N_18772);
nor U19023 (N_19023,N_18633,N_18954);
nand U19024 (N_19024,N_18502,N_18585);
nor U19025 (N_19025,N_18514,N_18834);
xor U19026 (N_19026,N_18984,N_18760);
nor U19027 (N_19027,N_18837,N_18844);
nor U19028 (N_19028,N_18861,N_18667);
nor U19029 (N_19029,N_18698,N_18990);
xnor U19030 (N_19030,N_18790,N_18821);
or U19031 (N_19031,N_18788,N_18887);
xnor U19032 (N_19032,N_18690,N_18769);
xnor U19033 (N_19033,N_18573,N_18994);
and U19034 (N_19034,N_18993,N_18539);
nor U19035 (N_19035,N_18775,N_18668);
nand U19036 (N_19036,N_18774,N_18895);
nand U19037 (N_19037,N_18660,N_18662);
or U19038 (N_19038,N_18548,N_18755);
and U19039 (N_19039,N_18828,N_18561);
and U19040 (N_19040,N_18734,N_18558);
xor U19041 (N_19041,N_18936,N_18714);
xnor U19042 (N_19042,N_18823,N_18518);
nand U19043 (N_19043,N_18746,N_18520);
or U19044 (N_19044,N_18829,N_18683);
and U19045 (N_19045,N_18655,N_18628);
and U19046 (N_19046,N_18991,N_18500);
or U19047 (N_19047,N_18808,N_18873);
nand U19048 (N_19048,N_18569,N_18512);
nor U19049 (N_19049,N_18878,N_18699);
or U19050 (N_19050,N_18577,N_18505);
nand U19051 (N_19051,N_18813,N_18762);
and U19052 (N_19052,N_18963,N_18931);
xnor U19053 (N_19053,N_18842,N_18966);
or U19054 (N_19054,N_18770,N_18845);
and U19055 (N_19055,N_18904,N_18782);
and U19056 (N_19056,N_18924,N_18923);
nand U19057 (N_19057,N_18789,N_18757);
xnor U19058 (N_19058,N_18773,N_18553);
xnor U19059 (N_19059,N_18781,N_18863);
or U19060 (N_19060,N_18637,N_18961);
nor U19061 (N_19061,N_18889,N_18802);
and U19062 (N_19062,N_18712,N_18592);
or U19063 (N_19063,N_18600,N_18817);
nand U19064 (N_19064,N_18747,N_18519);
and U19065 (N_19065,N_18910,N_18675);
or U19066 (N_19066,N_18749,N_18820);
nand U19067 (N_19067,N_18651,N_18616);
xnor U19068 (N_19068,N_18508,N_18664);
nand U19069 (N_19069,N_18639,N_18935);
or U19070 (N_19070,N_18711,N_18741);
or U19071 (N_19071,N_18752,N_18882);
and U19072 (N_19072,N_18709,N_18960);
xor U19073 (N_19073,N_18522,N_18672);
nor U19074 (N_19074,N_18976,N_18846);
xor U19075 (N_19075,N_18684,N_18606);
and U19076 (N_19076,N_18691,N_18909);
nand U19077 (N_19077,N_18981,N_18927);
or U19078 (N_19078,N_18796,N_18942);
nand U19079 (N_19079,N_18835,N_18611);
nor U19080 (N_19080,N_18725,N_18517);
or U19081 (N_19081,N_18511,N_18851);
and U19082 (N_19082,N_18750,N_18605);
or U19083 (N_19083,N_18753,N_18995);
xnor U19084 (N_19084,N_18534,N_18946);
nor U19085 (N_19085,N_18891,N_18696);
or U19086 (N_19086,N_18663,N_18645);
nor U19087 (N_19087,N_18647,N_18971);
nor U19088 (N_19088,N_18596,N_18677);
nand U19089 (N_19089,N_18792,N_18630);
or U19090 (N_19090,N_18533,N_18849);
and U19091 (N_19091,N_18886,N_18893);
xor U19092 (N_19092,N_18581,N_18560);
or U19093 (N_19093,N_18503,N_18965);
xor U19094 (N_19094,N_18610,N_18949);
and U19095 (N_19095,N_18665,N_18885);
nand U19096 (N_19096,N_18700,N_18959);
nor U19097 (N_19097,N_18756,N_18557);
nand U19098 (N_19098,N_18550,N_18578);
nor U19099 (N_19099,N_18972,N_18874);
nor U19100 (N_19100,N_18701,N_18912);
xnor U19101 (N_19101,N_18804,N_18621);
nand U19102 (N_19102,N_18726,N_18525);
nor U19103 (N_19103,N_18962,N_18722);
nor U19104 (N_19104,N_18836,N_18881);
nand U19105 (N_19105,N_18728,N_18634);
nand U19106 (N_19106,N_18919,N_18830);
nor U19107 (N_19107,N_18738,N_18812);
xor U19108 (N_19108,N_18778,N_18806);
or U19109 (N_19109,N_18902,N_18871);
xnor U19110 (N_19110,N_18916,N_18670);
nand U19111 (N_19111,N_18674,N_18776);
and U19112 (N_19112,N_18705,N_18707);
and U19113 (N_19113,N_18780,N_18579);
and U19114 (N_19114,N_18609,N_18855);
and U19115 (N_19115,N_18689,N_18652);
nor U19116 (N_19116,N_18763,N_18513);
nand U19117 (N_19117,N_18930,N_18783);
nor U19118 (N_19118,N_18627,N_18974);
xor U19119 (N_19119,N_18801,N_18799);
nand U19120 (N_19120,N_18985,N_18642);
nand U19121 (N_19121,N_18719,N_18786);
and U19122 (N_19122,N_18529,N_18818);
or U19123 (N_19123,N_18536,N_18716);
nor U19124 (N_19124,N_18809,N_18922);
nor U19125 (N_19125,N_18532,N_18531);
nor U19126 (N_19126,N_18681,N_18859);
xor U19127 (N_19127,N_18545,N_18825);
or U19128 (N_19128,N_18814,N_18815);
nand U19129 (N_19129,N_18939,N_18625);
nand U19130 (N_19130,N_18501,N_18840);
or U19131 (N_19131,N_18727,N_18593);
xnor U19132 (N_19132,N_18692,N_18929);
or U19133 (N_19133,N_18787,N_18898);
nor U19134 (N_19134,N_18831,N_18740);
nand U19135 (N_19135,N_18506,N_18552);
nand U19136 (N_19136,N_18706,N_18979);
or U19137 (N_19137,N_18811,N_18970);
nand U19138 (N_19138,N_18847,N_18944);
or U19139 (N_19139,N_18955,N_18967);
nor U19140 (N_19140,N_18798,N_18743);
or U19141 (N_19141,N_18805,N_18989);
or U19142 (N_19142,N_18551,N_18631);
or U19143 (N_19143,N_18657,N_18595);
or U19144 (N_19144,N_18576,N_18527);
or U19145 (N_19145,N_18999,N_18791);
xnor U19146 (N_19146,N_18925,N_18638);
nor U19147 (N_19147,N_18950,N_18643);
and U19148 (N_19148,N_18897,N_18973);
and U19149 (N_19149,N_18869,N_18562);
nor U19150 (N_19150,N_18682,N_18824);
or U19151 (N_19151,N_18862,N_18988);
nand U19152 (N_19152,N_18879,N_18964);
nand U19153 (N_19153,N_18736,N_18733);
and U19154 (N_19154,N_18986,N_18983);
or U19155 (N_19155,N_18819,N_18530);
nor U19156 (N_19156,N_18838,N_18724);
or U19157 (N_19157,N_18516,N_18807);
and U19158 (N_19158,N_18771,N_18507);
xnor U19159 (N_19159,N_18678,N_18666);
nand U19160 (N_19160,N_18659,N_18883);
nor U19161 (N_19161,N_18880,N_18629);
nand U19162 (N_19162,N_18918,N_18661);
xnor U19163 (N_19163,N_18795,N_18915);
nand U19164 (N_19164,N_18737,N_18731);
and U19165 (N_19165,N_18713,N_18860);
nor U19166 (N_19166,N_18721,N_18998);
nor U19167 (N_19167,N_18624,N_18537);
nor U19168 (N_19168,N_18932,N_18940);
or U19169 (N_19169,N_18694,N_18648);
and U19170 (N_19170,N_18956,N_18875);
and U19171 (N_19171,N_18572,N_18833);
nor U19172 (N_19172,N_18598,N_18622);
nor U19173 (N_19173,N_18566,N_18555);
nor U19174 (N_19174,N_18717,N_18586);
nor U19175 (N_19175,N_18816,N_18793);
nor U19176 (N_19176,N_18549,N_18623);
and U19177 (N_19177,N_18876,N_18649);
and U19178 (N_19178,N_18564,N_18635);
nand U19179 (N_19179,N_18947,N_18715);
and U19180 (N_19180,N_18618,N_18867);
or U19181 (N_19181,N_18703,N_18571);
nand U19182 (N_19182,N_18748,N_18951);
and U19183 (N_19183,N_18574,N_18866);
nand U19184 (N_19184,N_18894,N_18899);
and U19185 (N_19185,N_18900,N_18987);
xor U19186 (N_19186,N_18547,N_18853);
or U19187 (N_19187,N_18582,N_18896);
or U19188 (N_19188,N_18868,N_18544);
nor U19189 (N_19189,N_18535,N_18854);
nand U19190 (N_19190,N_18546,N_18526);
or U19191 (N_19191,N_18615,N_18953);
or U19192 (N_19192,N_18832,N_18613);
nand U19193 (N_19193,N_18892,N_18686);
xor U19194 (N_19194,N_18941,N_18913);
or U19195 (N_19195,N_18803,N_18921);
and U19196 (N_19196,N_18608,N_18653);
nand U19197 (N_19197,N_18997,N_18800);
nor U19198 (N_19198,N_18524,N_18758);
nor U19199 (N_19199,N_18540,N_18865);
nand U19200 (N_19200,N_18541,N_18650);
or U19201 (N_19201,N_18556,N_18693);
xor U19202 (N_19202,N_18607,N_18980);
and U19203 (N_19203,N_18841,N_18958);
or U19204 (N_19204,N_18978,N_18785);
and U19205 (N_19205,N_18977,N_18723);
xor U19206 (N_19206,N_18565,N_18744);
nand U19207 (N_19207,N_18620,N_18644);
or U19208 (N_19208,N_18822,N_18568);
or U19209 (N_19209,N_18599,N_18509);
or U19210 (N_19210,N_18870,N_18843);
or U19211 (N_19211,N_18735,N_18679);
xnor U19212 (N_19212,N_18612,N_18604);
and U19213 (N_19213,N_18938,N_18656);
nand U19214 (N_19214,N_18587,N_18697);
xor U19215 (N_19215,N_18641,N_18937);
and U19216 (N_19216,N_18905,N_18907);
or U19217 (N_19217,N_18543,N_18856);
or U19218 (N_19218,N_18906,N_18720);
nand U19219 (N_19219,N_18730,N_18928);
nand U19220 (N_19220,N_18680,N_18996);
and U19221 (N_19221,N_18761,N_18589);
nand U19222 (N_19222,N_18542,N_18584);
and U19223 (N_19223,N_18708,N_18901);
xnor U19224 (N_19224,N_18884,N_18704);
and U19225 (N_19225,N_18975,N_18583);
xor U19226 (N_19226,N_18797,N_18538);
or U19227 (N_19227,N_18588,N_18969);
nand U19228 (N_19228,N_18732,N_18695);
nor U19229 (N_19229,N_18567,N_18729);
nor U19230 (N_19230,N_18515,N_18575);
nand U19231 (N_19231,N_18810,N_18563);
nor U19232 (N_19232,N_18779,N_18654);
xor U19233 (N_19233,N_18957,N_18590);
nand U19234 (N_19234,N_18952,N_18888);
and U19235 (N_19235,N_18852,N_18765);
and U19236 (N_19236,N_18742,N_18948);
and U19237 (N_19237,N_18504,N_18864);
nor U19238 (N_19238,N_18943,N_18764);
or U19239 (N_19239,N_18982,N_18671);
and U19240 (N_19240,N_18601,N_18591);
and U19241 (N_19241,N_18602,N_18933);
nand U19242 (N_19242,N_18528,N_18992);
xnor U19243 (N_19243,N_18920,N_18872);
and U19244 (N_19244,N_18877,N_18594);
and U19245 (N_19245,N_18640,N_18710);
or U19246 (N_19246,N_18580,N_18632);
or U19247 (N_19247,N_18767,N_18685);
nor U19248 (N_19248,N_18914,N_18766);
xor U19249 (N_19249,N_18857,N_18826);
nor U19250 (N_19250,N_18704,N_18879);
xor U19251 (N_19251,N_18846,N_18552);
and U19252 (N_19252,N_18979,N_18775);
xnor U19253 (N_19253,N_18738,N_18589);
xnor U19254 (N_19254,N_18669,N_18893);
xnor U19255 (N_19255,N_18921,N_18766);
xnor U19256 (N_19256,N_18661,N_18549);
nand U19257 (N_19257,N_18592,N_18697);
nand U19258 (N_19258,N_18731,N_18925);
nand U19259 (N_19259,N_18810,N_18839);
nor U19260 (N_19260,N_18816,N_18857);
or U19261 (N_19261,N_18510,N_18524);
nand U19262 (N_19262,N_18656,N_18752);
xor U19263 (N_19263,N_18513,N_18727);
xnor U19264 (N_19264,N_18575,N_18583);
and U19265 (N_19265,N_18708,N_18534);
nor U19266 (N_19266,N_18630,N_18769);
nor U19267 (N_19267,N_18969,N_18930);
nor U19268 (N_19268,N_18513,N_18834);
nor U19269 (N_19269,N_18605,N_18782);
and U19270 (N_19270,N_18847,N_18918);
nor U19271 (N_19271,N_18533,N_18575);
xor U19272 (N_19272,N_18609,N_18997);
nand U19273 (N_19273,N_18876,N_18758);
nand U19274 (N_19274,N_18800,N_18777);
and U19275 (N_19275,N_18754,N_18897);
or U19276 (N_19276,N_18508,N_18670);
nor U19277 (N_19277,N_18607,N_18764);
nand U19278 (N_19278,N_18603,N_18633);
nor U19279 (N_19279,N_18523,N_18857);
or U19280 (N_19280,N_18589,N_18780);
nor U19281 (N_19281,N_18804,N_18697);
nand U19282 (N_19282,N_18755,N_18689);
nor U19283 (N_19283,N_18876,N_18644);
nand U19284 (N_19284,N_18651,N_18583);
nor U19285 (N_19285,N_18898,N_18903);
nor U19286 (N_19286,N_18612,N_18742);
nand U19287 (N_19287,N_18674,N_18562);
or U19288 (N_19288,N_18686,N_18572);
or U19289 (N_19289,N_18757,N_18949);
or U19290 (N_19290,N_18846,N_18657);
or U19291 (N_19291,N_18873,N_18738);
nor U19292 (N_19292,N_18831,N_18793);
and U19293 (N_19293,N_18836,N_18878);
nand U19294 (N_19294,N_18620,N_18559);
or U19295 (N_19295,N_18916,N_18771);
xor U19296 (N_19296,N_18996,N_18923);
xnor U19297 (N_19297,N_18534,N_18689);
xor U19298 (N_19298,N_18997,N_18908);
nand U19299 (N_19299,N_18640,N_18960);
and U19300 (N_19300,N_18833,N_18927);
nand U19301 (N_19301,N_18796,N_18683);
nor U19302 (N_19302,N_18684,N_18659);
xnor U19303 (N_19303,N_18601,N_18769);
or U19304 (N_19304,N_18753,N_18847);
nor U19305 (N_19305,N_18977,N_18927);
and U19306 (N_19306,N_18707,N_18976);
or U19307 (N_19307,N_18624,N_18802);
and U19308 (N_19308,N_18850,N_18864);
nand U19309 (N_19309,N_18747,N_18638);
or U19310 (N_19310,N_18620,N_18970);
nor U19311 (N_19311,N_18983,N_18872);
xnor U19312 (N_19312,N_18947,N_18957);
or U19313 (N_19313,N_18881,N_18738);
nor U19314 (N_19314,N_18717,N_18875);
nor U19315 (N_19315,N_18616,N_18768);
nor U19316 (N_19316,N_18584,N_18823);
and U19317 (N_19317,N_18608,N_18685);
and U19318 (N_19318,N_18613,N_18711);
or U19319 (N_19319,N_18531,N_18655);
or U19320 (N_19320,N_18565,N_18794);
and U19321 (N_19321,N_18621,N_18818);
xor U19322 (N_19322,N_18700,N_18680);
or U19323 (N_19323,N_18877,N_18809);
xor U19324 (N_19324,N_18980,N_18582);
and U19325 (N_19325,N_18605,N_18570);
nand U19326 (N_19326,N_18543,N_18678);
nand U19327 (N_19327,N_18703,N_18652);
xnor U19328 (N_19328,N_18969,N_18825);
nor U19329 (N_19329,N_18953,N_18532);
nand U19330 (N_19330,N_18854,N_18563);
xor U19331 (N_19331,N_18638,N_18876);
and U19332 (N_19332,N_18953,N_18515);
nand U19333 (N_19333,N_18530,N_18896);
nor U19334 (N_19334,N_18750,N_18660);
nor U19335 (N_19335,N_18733,N_18937);
nor U19336 (N_19336,N_18704,N_18745);
or U19337 (N_19337,N_18943,N_18961);
nand U19338 (N_19338,N_18761,N_18550);
or U19339 (N_19339,N_18890,N_18847);
or U19340 (N_19340,N_18753,N_18749);
nor U19341 (N_19341,N_18800,N_18760);
nor U19342 (N_19342,N_18759,N_18937);
or U19343 (N_19343,N_18667,N_18808);
nand U19344 (N_19344,N_18836,N_18884);
nand U19345 (N_19345,N_18572,N_18828);
nor U19346 (N_19346,N_18690,N_18907);
and U19347 (N_19347,N_18677,N_18997);
or U19348 (N_19348,N_18857,N_18988);
and U19349 (N_19349,N_18677,N_18615);
or U19350 (N_19350,N_18860,N_18874);
nand U19351 (N_19351,N_18592,N_18774);
nor U19352 (N_19352,N_18760,N_18564);
nor U19353 (N_19353,N_18761,N_18908);
nor U19354 (N_19354,N_18735,N_18619);
or U19355 (N_19355,N_18530,N_18771);
nor U19356 (N_19356,N_18650,N_18969);
and U19357 (N_19357,N_18725,N_18542);
or U19358 (N_19358,N_18649,N_18858);
xor U19359 (N_19359,N_18621,N_18603);
or U19360 (N_19360,N_18591,N_18538);
nand U19361 (N_19361,N_18954,N_18923);
xnor U19362 (N_19362,N_18962,N_18842);
xnor U19363 (N_19363,N_18896,N_18845);
and U19364 (N_19364,N_18931,N_18661);
nand U19365 (N_19365,N_18736,N_18791);
or U19366 (N_19366,N_18812,N_18684);
or U19367 (N_19367,N_18742,N_18731);
xor U19368 (N_19368,N_18836,N_18574);
or U19369 (N_19369,N_18984,N_18859);
and U19370 (N_19370,N_18634,N_18981);
nand U19371 (N_19371,N_18703,N_18751);
or U19372 (N_19372,N_18867,N_18557);
nor U19373 (N_19373,N_18501,N_18649);
nand U19374 (N_19374,N_18827,N_18506);
and U19375 (N_19375,N_18710,N_18839);
nand U19376 (N_19376,N_18777,N_18822);
nor U19377 (N_19377,N_18966,N_18717);
nor U19378 (N_19378,N_18549,N_18630);
xnor U19379 (N_19379,N_18776,N_18783);
xor U19380 (N_19380,N_18631,N_18698);
or U19381 (N_19381,N_18591,N_18791);
xor U19382 (N_19382,N_18720,N_18735);
xor U19383 (N_19383,N_18526,N_18776);
and U19384 (N_19384,N_18602,N_18831);
xnor U19385 (N_19385,N_18925,N_18817);
nand U19386 (N_19386,N_18840,N_18875);
xor U19387 (N_19387,N_18758,N_18657);
or U19388 (N_19388,N_18886,N_18641);
xnor U19389 (N_19389,N_18542,N_18793);
nor U19390 (N_19390,N_18647,N_18947);
or U19391 (N_19391,N_18512,N_18731);
or U19392 (N_19392,N_18954,N_18660);
xor U19393 (N_19393,N_18616,N_18902);
nor U19394 (N_19394,N_18924,N_18593);
xnor U19395 (N_19395,N_18774,N_18731);
nand U19396 (N_19396,N_18877,N_18989);
nand U19397 (N_19397,N_18902,N_18874);
nand U19398 (N_19398,N_18524,N_18856);
nand U19399 (N_19399,N_18529,N_18686);
and U19400 (N_19400,N_18848,N_18663);
and U19401 (N_19401,N_18613,N_18626);
nand U19402 (N_19402,N_18501,N_18894);
or U19403 (N_19403,N_18715,N_18887);
xor U19404 (N_19404,N_18640,N_18954);
nand U19405 (N_19405,N_18791,N_18664);
or U19406 (N_19406,N_18502,N_18740);
and U19407 (N_19407,N_18721,N_18755);
or U19408 (N_19408,N_18693,N_18651);
xnor U19409 (N_19409,N_18810,N_18726);
nand U19410 (N_19410,N_18558,N_18908);
nor U19411 (N_19411,N_18957,N_18806);
nor U19412 (N_19412,N_18710,N_18767);
and U19413 (N_19413,N_18828,N_18577);
and U19414 (N_19414,N_18654,N_18787);
nor U19415 (N_19415,N_18533,N_18800);
and U19416 (N_19416,N_18797,N_18854);
xor U19417 (N_19417,N_18680,N_18922);
nand U19418 (N_19418,N_18872,N_18529);
or U19419 (N_19419,N_18957,N_18856);
xor U19420 (N_19420,N_18737,N_18565);
or U19421 (N_19421,N_18709,N_18799);
or U19422 (N_19422,N_18703,N_18679);
nor U19423 (N_19423,N_18929,N_18537);
or U19424 (N_19424,N_18886,N_18860);
nand U19425 (N_19425,N_18514,N_18548);
xnor U19426 (N_19426,N_18587,N_18643);
nand U19427 (N_19427,N_18940,N_18963);
nor U19428 (N_19428,N_18893,N_18726);
or U19429 (N_19429,N_18998,N_18577);
xor U19430 (N_19430,N_18927,N_18784);
nand U19431 (N_19431,N_18920,N_18595);
nor U19432 (N_19432,N_18672,N_18891);
or U19433 (N_19433,N_18749,N_18748);
xor U19434 (N_19434,N_18539,N_18905);
or U19435 (N_19435,N_18611,N_18870);
and U19436 (N_19436,N_18516,N_18562);
and U19437 (N_19437,N_18741,N_18560);
and U19438 (N_19438,N_18807,N_18964);
or U19439 (N_19439,N_18851,N_18748);
xnor U19440 (N_19440,N_18726,N_18932);
and U19441 (N_19441,N_18882,N_18948);
xor U19442 (N_19442,N_18659,N_18763);
nand U19443 (N_19443,N_18879,N_18644);
and U19444 (N_19444,N_18954,N_18937);
nand U19445 (N_19445,N_18984,N_18968);
nor U19446 (N_19446,N_18969,N_18713);
and U19447 (N_19447,N_18923,N_18913);
nor U19448 (N_19448,N_18790,N_18689);
nor U19449 (N_19449,N_18645,N_18799);
and U19450 (N_19450,N_18964,N_18968);
xnor U19451 (N_19451,N_18942,N_18739);
nand U19452 (N_19452,N_18918,N_18872);
and U19453 (N_19453,N_18669,N_18577);
nand U19454 (N_19454,N_18639,N_18930);
or U19455 (N_19455,N_18718,N_18684);
nand U19456 (N_19456,N_18501,N_18565);
xnor U19457 (N_19457,N_18815,N_18548);
and U19458 (N_19458,N_18552,N_18577);
or U19459 (N_19459,N_18882,N_18804);
nand U19460 (N_19460,N_18785,N_18611);
nand U19461 (N_19461,N_18543,N_18619);
nor U19462 (N_19462,N_18577,N_18698);
and U19463 (N_19463,N_18569,N_18898);
nand U19464 (N_19464,N_18698,N_18614);
and U19465 (N_19465,N_18730,N_18877);
xor U19466 (N_19466,N_18554,N_18576);
nand U19467 (N_19467,N_18580,N_18748);
and U19468 (N_19468,N_18798,N_18756);
xor U19469 (N_19469,N_18716,N_18638);
and U19470 (N_19470,N_18594,N_18671);
nor U19471 (N_19471,N_18810,N_18701);
nor U19472 (N_19472,N_18612,N_18653);
nand U19473 (N_19473,N_18838,N_18808);
nand U19474 (N_19474,N_18761,N_18548);
nor U19475 (N_19475,N_18884,N_18986);
nor U19476 (N_19476,N_18770,N_18609);
and U19477 (N_19477,N_18688,N_18857);
nor U19478 (N_19478,N_18627,N_18664);
nor U19479 (N_19479,N_18952,N_18772);
and U19480 (N_19480,N_18700,N_18541);
or U19481 (N_19481,N_18853,N_18888);
nor U19482 (N_19482,N_18934,N_18847);
and U19483 (N_19483,N_18937,N_18516);
nand U19484 (N_19484,N_18529,N_18858);
nand U19485 (N_19485,N_18979,N_18810);
xnor U19486 (N_19486,N_18642,N_18608);
xor U19487 (N_19487,N_18899,N_18977);
nand U19488 (N_19488,N_18909,N_18969);
and U19489 (N_19489,N_18644,N_18862);
nor U19490 (N_19490,N_18607,N_18720);
nand U19491 (N_19491,N_18962,N_18938);
or U19492 (N_19492,N_18879,N_18759);
nor U19493 (N_19493,N_18627,N_18959);
or U19494 (N_19494,N_18792,N_18991);
xor U19495 (N_19495,N_18903,N_18983);
nand U19496 (N_19496,N_18762,N_18520);
xor U19497 (N_19497,N_18757,N_18739);
nor U19498 (N_19498,N_18990,N_18792);
nand U19499 (N_19499,N_18879,N_18750);
or U19500 (N_19500,N_19084,N_19232);
or U19501 (N_19501,N_19105,N_19327);
and U19502 (N_19502,N_19140,N_19284);
and U19503 (N_19503,N_19425,N_19361);
xnor U19504 (N_19504,N_19355,N_19283);
and U19505 (N_19505,N_19391,N_19173);
nor U19506 (N_19506,N_19144,N_19466);
xor U19507 (N_19507,N_19346,N_19223);
xor U19508 (N_19508,N_19026,N_19274);
nand U19509 (N_19509,N_19062,N_19297);
or U19510 (N_19510,N_19047,N_19158);
nor U19511 (N_19511,N_19028,N_19354);
nor U19512 (N_19512,N_19418,N_19392);
xnor U19513 (N_19513,N_19176,N_19243);
and U19514 (N_19514,N_19395,N_19076);
or U19515 (N_19515,N_19489,N_19290);
and U19516 (N_19516,N_19427,N_19317);
and U19517 (N_19517,N_19277,N_19436);
nor U19518 (N_19518,N_19342,N_19226);
or U19519 (N_19519,N_19396,N_19068);
xor U19520 (N_19520,N_19204,N_19357);
nand U19521 (N_19521,N_19155,N_19293);
nor U19522 (N_19522,N_19167,N_19270);
nand U19523 (N_19523,N_19246,N_19302);
and U19524 (N_19524,N_19213,N_19292);
xor U19525 (N_19525,N_19258,N_19424);
nand U19526 (N_19526,N_19151,N_19136);
nand U19527 (N_19527,N_19032,N_19216);
nand U19528 (N_19528,N_19483,N_19325);
xor U19529 (N_19529,N_19043,N_19334);
nor U19530 (N_19530,N_19397,N_19042);
xnor U19531 (N_19531,N_19078,N_19372);
nor U19532 (N_19532,N_19021,N_19016);
nor U19533 (N_19533,N_19240,N_19338);
nor U19534 (N_19534,N_19071,N_19400);
or U19535 (N_19535,N_19492,N_19348);
xnor U19536 (N_19536,N_19091,N_19141);
or U19537 (N_19537,N_19005,N_19153);
and U19538 (N_19538,N_19253,N_19012);
nor U19539 (N_19539,N_19107,N_19434);
or U19540 (N_19540,N_19380,N_19299);
nand U19541 (N_19541,N_19499,N_19428);
xor U19542 (N_19542,N_19145,N_19367);
nor U19543 (N_19543,N_19377,N_19426);
or U19544 (N_19544,N_19175,N_19234);
nand U19545 (N_19545,N_19461,N_19497);
or U19546 (N_19546,N_19450,N_19134);
and U19547 (N_19547,N_19237,N_19099);
nand U19548 (N_19548,N_19018,N_19316);
or U19549 (N_19549,N_19331,N_19387);
nor U19550 (N_19550,N_19459,N_19255);
xor U19551 (N_19551,N_19041,N_19094);
nor U19552 (N_19552,N_19329,N_19291);
xnor U19553 (N_19553,N_19196,N_19064);
xnor U19554 (N_19554,N_19287,N_19369);
xnor U19555 (N_19555,N_19356,N_19447);
nor U19556 (N_19556,N_19161,N_19476);
xor U19557 (N_19557,N_19166,N_19206);
nand U19558 (N_19558,N_19444,N_19343);
and U19559 (N_19559,N_19079,N_19315);
nand U19560 (N_19560,N_19264,N_19421);
nor U19561 (N_19561,N_19414,N_19104);
xnor U19562 (N_19562,N_19265,N_19138);
nand U19563 (N_19563,N_19469,N_19229);
or U19564 (N_19564,N_19239,N_19388);
or U19565 (N_19565,N_19422,N_19326);
xor U19566 (N_19566,N_19247,N_19275);
xor U19567 (N_19567,N_19089,N_19164);
nor U19568 (N_19568,N_19221,N_19106);
nor U19569 (N_19569,N_19464,N_19238);
nand U19570 (N_19570,N_19061,N_19478);
or U19571 (N_19571,N_19095,N_19301);
xor U19572 (N_19572,N_19199,N_19098);
and U19573 (N_19573,N_19405,N_19220);
or U19574 (N_19574,N_19114,N_19092);
or U19575 (N_19575,N_19252,N_19403);
nand U19576 (N_19576,N_19118,N_19117);
or U19577 (N_19577,N_19137,N_19431);
and U19578 (N_19578,N_19188,N_19437);
or U19579 (N_19579,N_19055,N_19126);
xnor U19580 (N_19580,N_19458,N_19452);
nand U19581 (N_19581,N_19182,N_19318);
nor U19582 (N_19582,N_19360,N_19177);
and U19583 (N_19583,N_19472,N_19310);
nor U19584 (N_19584,N_19011,N_19113);
nand U19585 (N_19585,N_19410,N_19097);
nor U19586 (N_19586,N_19203,N_19143);
or U19587 (N_19587,N_19149,N_19251);
xnor U19588 (N_19588,N_19050,N_19462);
or U19589 (N_19589,N_19244,N_19368);
or U19590 (N_19590,N_19314,N_19451);
nand U19591 (N_19591,N_19259,N_19474);
nand U19592 (N_19592,N_19040,N_19096);
xor U19593 (N_19593,N_19051,N_19004);
xor U19594 (N_19594,N_19101,N_19069);
and U19595 (N_19595,N_19415,N_19350);
and U19596 (N_19596,N_19193,N_19341);
nand U19597 (N_19597,N_19086,N_19228);
xnor U19598 (N_19598,N_19448,N_19139);
and U19599 (N_19599,N_19323,N_19121);
or U19600 (N_19600,N_19305,N_19148);
and U19601 (N_19601,N_19194,N_19183);
xnor U19602 (N_19602,N_19067,N_19457);
and U19603 (N_19603,N_19273,N_19147);
xor U19604 (N_19604,N_19411,N_19172);
xor U19605 (N_19605,N_19195,N_19300);
nor U19606 (N_19606,N_19419,N_19322);
or U19607 (N_19607,N_19029,N_19242);
or U19608 (N_19608,N_19103,N_19201);
nor U19609 (N_19609,N_19218,N_19465);
or U19610 (N_19610,N_19420,N_19442);
and U19611 (N_19611,N_19260,N_19192);
xor U19612 (N_19612,N_19481,N_19333);
and U19613 (N_19613,N_19030,N_19313);
nand U19614 (N_19614,N_19120,N_19109);
nor U19615 (N_19615,N_19031,N_19335);
nor U19616 (N_19616,N_19351,N_19445);
nand U19617 (N_19617,N_19254,N_19198);
and U19618 (N_19618,N_19007,N_19054);
nor U19619 (N_19619,N_19443,N_19053);
nand U19620 (N_19620,N_19046,N_19233);
or U19621 (N_19621,N_19495,N_19044);
nand U19622 (N_19622,N_19152,N_19268);
or U19623 (N_19623,N_19404,N_19150);
xor U19624 (N_19624,N_19430,N_19477);
nor U19625 (N_19625,N_19340,N_19449);
or U19626 (N_19626,N_19025,N_19321);
or U19627 (N_19627,N_19438,N_19065);
nor U19628 (N_19628,N_19319,N_19278);
xor U19629 (N_19629,N_19132,N_19460);
or U19630 (N_19630,N_19473,N_19470);
xnor U19631 (N_19631,N_19169,N_19487);
nor U19632 (N_19632,N_19189,N_19123);
or U19633 (N_19633,N_19394,N_19439);
or U19634 (N_19634,N_19399,N_19231);
or U19635 (N_19635,N_19250,N_19288);
nor U19636 (N_19636,N_19467,N_19225);
and U19637 (N_19637,N_19130,N_19453);
nor U19638 (N_19638,N_19142,N_19115);
or U19639 (N_19639,N_19498,N_19215);
nand U19640 (N_19640,N_19056,N_19363);
nand U19641 (N_19641,N_19073,N_19339);
nor U19642 (N_19642,N_19208,N_19324);
nand U19643 (N_19643,N_19306,N_19129);
and U19644 (N_19644,N_19190,N_19257);
nor U19645 (N_19645,N_19365,N_19261);
and U19646 (N_19646,N_19217,N_19441);
nor U19647 (N_19647,N_19312,N_19127);
xor U19648 (N_19648,N_19010,N_19308);
and U19649 (N_19649,N_19307,N_19022);
xor U19650 (N_19650,N_19282,N_19154);
nor U19651 (N_19651,N_19162,N_19384);
or U19652 (N_19652,N_19320,N_19235);
nand U19653 (N_19653,N_19200,N_19370);
and U19654 (N_19654,N_19432,N_19416);
nand U19655 (N_19655,N_19386,N_19295);
and U19656 (N_19656,N_19186,N_19330);
xor U19657 (N_19657,N_19376,N_19146);
and U19658 (N_19658,N_19000,N_19456);
xor U19659 (N_19659,N_19245,N_19379);
nor U19660 (N_19660,N_19048,N_19383);
nor U19661 (N_19661,N_19468,N_19358);
nor U19662 (N_19662,N_19389,N_19075);
nand U19663 (N_19663,N_19087,N_19085);
and U19664 (N_19664,N_19219,N_19174);
or U19665 (N_19665,N_19423,N_19241);
and U19666 (N_19666,N_19493,N_19222);
nand U19667 (N_19667,N_19006,N_19057);
and U19668 (N_19668,N_19034,N_19165);
nor U19669 (N_19669,N_19205,N_19074);
nand U19670 (N_19670,N_19267,N_19353);
or U19671 (N_19671,N_19197,N_19266);
and U19672 (N_19672,N_19125,N_19133);
and U19673 (N_19673,N_19393,N_19408);
xnor U19674 (N_19674,N_19036,N_19170);
nand U19675 (N_19675,N_19072,N_19433);
nand U19676 (N_19676,N_19224,N_19381);
nand U19677 (N_19677,N_19180,N_19080);
nand U19678 (N_19678,N_19328,N_19289);
nand U19679 (N_19679,N_19116,N_19280);
and U19680 (N_19680,N_19406,N_19463);
nor U19681 (N_19681,N_19382,N_19081);
nor U19682 (N_19682,N_19185,N_19093);
or U19683 (N_19683,N_19332,N_19008);
xor U19684 (N_19684,N_19063,N_19210);
xnor U19685 (N_19685,N_19269,N_19013);
xnor U19686 (N_19686,N_19413,N_19017);
xor U19687 (N_19687,N_19045,N_19248);
or U19688 (N_19688,N_19088,N_19263);
nand U19689 (N_19689,N_19187,N_19385);
and U19690 (N_19690,N_19168,N_19336);
nand U19691 (N_19691,N_19286,N_19037);
or U19692 (N_19692,N_19060,N_19440);
nor U19693 (N_19693,N_19412,N_19362);
or U19694 (N_19694,N_19344,N_19119);
nor U19695 (N_19695,N_19271,N_19135);
and U19696 (N_19696,N_19131,N_19407);
xnor U19697 (N_19697,N_19214,N_19202);
or U19698 (N_19698,N_19446,N_19490);
nor U19699 (N_19699,N_19352,N_19178);
and U19700 (N_19700,N_19390,N_19309);
xor U19701 (N_19701,N_19038,N_19409);
and U19702 (N_19702,N_19304,N_19077);
nand U19703 (N_19703,N_19294,N_19157);
nor U19704 (N_19704,N_19491,N_19480);
or U19705 (N_19705,N_19272,N_19475);
or U19706 (N_19706,N_19279,N_19015);
or U19707 (N_19707,N_19285,N_19375);
and U19708 (N_19708,N_19179,N_19281);
nand U19709 (N_19709,N_19366,N_19378);
nand U19710 (N_19710,N_19002,N_19471);
nor U19711 (N_19711,N_19303,N_19052);
nor U19712 (N_19712,N_19102,N_19184);
nor U19713 (N_19713,N_19371,N_19488);
or U19714 (N_19714,N_19494,N_19211);
xnor U19715 (N_19715,N_19337,N_19454);
or U19716 (N_19716,N_19359,N_19160);
xor U19717 (N_19717,N_19209,N_19111);
nor U19718 (N_19718,N_19023,N_19256);
or U19719 (N_19719,N_19128,N_19455);
and U19720 (N_19720,N_19311,N_19124);
and U19721 (N_19721,N_19066,N_19398);
or U19722 (N_19722,N_19207,N_19401);
nor U19723 (N_19723,N_19014,N_19003);
or U19724 (N_19724,N_19296,N_19236);
nand U19725 (N_19725,N_19298,N_19171);
xnor U19726 (N_19726,N_19227,N_19496);
and U19727 (N_19727,N_19108,N_19249);
or U19728 (N_19728,N_19484,N_19181);
nor U19729 (N_19729,N_19435,N_19345);
and U19730 (N_19730,N_19009,N_19122);
or U19731 (N_19731,N_19024,N_19349);
and U19732 (N_19732,N_19001,N_19486);
or U19733 (N_19733,N_19374,N_19027);
nor U19734 (N_19734,N_19479,N_19059);
nand U19735 (N_19735,N_19019,N_19020);
or U19736 (N_19736,N_19230,N_19191);
xor U19737 (N_19737,N_19364,N_19485);
or U19738 (N_19738,N_19156,N_19070);
nor U19739 (N_19739,N_19049,N_19212);
and U19740 (N_19740,N_19112,N_19039);
xnor U19741 (N_19741,N_19163,N_19110);
and U19742 (N_19742,N_19090,N_19347);
or U19743 (N_19743,N_19429,N_19035);
and U19744 (N_19744,N_19402,N_19417);
or U19745 (N_19745,N_19082,N_19159);
nand U19746 (N_19746,N_19262,N_19058);
xor U19747 (N_19747,N_19083,N_19482);
nand U19748 (N_19748,N_19276,N_19100);
nor U19749 (N_19749,N_19373,N_19033);
and U19750 (N_19750,N_19086,N_19159);
nor U19751 (N_19751,N_19496,N_19035);
xnor U19752 (N_19752,N_19259,N_19492);
nand U19753 (N_19753,N_19304,N_19357);
or U19754 (N_19754,N_19094,N_19164);
nor U19755 (N_19755,N_19399,N_19487);
and U19756 (N_19756,N_19285,N_19201);
or U19757 (N_19757,N_19418,N_19299);
or U19758 (N_19758,N_19121,N_19436);
and U19759 (N_19759,N_19441,N_19198);
xor U19760 (N_19760,N_19435,N_19017);
nand U19761 (N_19761,N_19488,N_19406);
and U19762 (N_19762,N_19348,N_19356);
nor U19763 (N_19763,N_19003,N_19345);
nand U19764 (N_19764,N_19494,N_19303);
nor U19765 (N_19765,N_19042,N_19494);
nor U19766 (N_19766,N_19388,N_19292);
xor U19767 (N_19767,N_19482,N_19186);
xnor U19768 (N_19768,N_19051,N_19421);
and U19769 (N_19769,N_19437,N_19349);
nor U19770 (N_19770,N_19393,N_19128);
or U19771 (N_19771,N_19150,N_19011);
and U19772 (N_19772,N_19336,N_19034);
or U19773 (N_19773,N_19465,N_19485);
or U19774 (N_19774,N_19085,N_19388);
and U19775 (N_19775,N_19075,N_19405);
xor U19776 (N_19776,N_19349,N_19330);
or U19777 (N_19777,N_19167,N_19319);
and U19778 (N_19778,N_19305,N_19133);
and U19779 (N_19779,N_19437,N_19096);
nand U19780 (N_19780,N_19147,N_19302);
nor U19781 (N_19781,N_19207,N_19054);
xnor U19782 (N_19782,N_19047,N_19353);
nand U19783 (N_19783,N_19386,N_19463);
or U19784 (N_19784,N_19293,N_19435);
or U19785 (N_19785,N_19333,N_19494);
nand U19786 (N_19786,N_19127,N_19474);
xor U19787 (N_19787,N_19367,N_19426);
nand U19788 (N_19788,N_19104,N_19086);
nor U19789 (N_19789,N_19038,N_19262);
nor U19790 (N_19790,N_19080,N_19078);
and U19791 (N_19791,N_19325,N_19242);
nor U19792 (N_19792,N_19030,N_19467);
nor U19793 (N_19793,N_19317,N_19026);
xor U19794 (N_19794,N_19481,N_19316);
xor U19795 (N_19795,N_19086,N_19129);
and U19796 (N_19796,N_19484,N_19173);
xor U19797 (N_19797,N_19493,N_19170);
nor U19798 (N_19798,N_19464,N_19388);
or U19799 (N_19799,N_19044,N_19319);
nor U19800 (N_19800,N_19134,N_19057);
nor U19801 (N_19801,N_19121,N_19453);
nand U19802 (N_19802,N_19254,N_19390);
or U19803 (N_19803,N_19046,N_19487);
nor U19804 (N_19804,N_19494,N_19149);
nor U19805 (N_19805,N_19477,N_19259);
and U19806 (N_19806,N_19110,N_19194);
nand U19807 (N_19807,N_19436,N_19320);
or U19808 (N_19808,N_19256,N_19372);
and U19809 (N_19809,N_19483,N_19191);
and U19810 (N_19810,N_19139,N_19385);
nor U19811 (N_19811,N_19161,N_19138);
and U19812 (N_19812,N_19392,N_19422);
nand U19813 (N_19813,N_19221,N_19008);
xor U19814 (N_19814,N_19244,N_19300);
xor U19815 (N_19815,N_19021,N_19039);
and U19816 (N_19816,N_19391,N_19079);
nor U19817 (N_19817,N_19125,N_19496);
and U19818 (N_19818,N_19170,N_19024);
nand U19819 (N_19819,N_19006,N_19167);
nand U19820 (N_19820,N_19053,N_19056);
and U19821 (N_19821,N_19103,N_19099);
and U19822 (N_19822,N_19409,N_19007);
or U19823 (N_19823,N_19021,N_19022);
and U19824 (N_19824,N_19007,N_19074);
xor U19825 (N_19825,N_19436,N_19308);
xnor U19826 (N_19826,N_19094,N_19165);
and U19827 (N_19827,N_19244,N_19076);
and U19828 (N_19828,N_19002,N_19441);
nor U19829 (N_19829,N_19292,N_19168);
nor U19830 (N_19830,N_19486,N_19487);
nor U19831 (N_19831,N_19056,N_19384);
or U19832 (N_19832,N_19041,N_19004);
and U19833 (N_19833,N_19197,N_19243);
and U19834 (N_19834,N_19357,N_19459);
nor U19835 (N_19835,N_19098,N_19001);
or U19836 (N_19836,N_19238,N_19186);
nor U19837 (N_19837,N_19060,N_19093);
and U19838 (N_19838,N_19256,N_19285);
or U19839 (N_19839,N_19029,N_19472);
or U19840 (N_19840,N_19488,N_19023);
xnor U19841 (N_19841,N_19283,N_19161);
or U19842 (N_19842,N_19062,N_19440);
or U19843 (N_19843,N_19125,N_19393);
nand U19844 (N_19844,N_19309,N_19488);
nand U19845 (N_19845,N_19096,N_19016);
nor U19846 (N_19846,N_19099,N_19409);
and U19847 (N_19847,N_19358,N_19002);
xnor U19848 (N_19848,N_19368,N_19216);
nor U19849 (N_19849,N_19105,N_19485);
or U19850 (N_19850,N_19252,N_19011);
nand U19851 (N_19851,N_19299,N_19347);
or U19852 (N_19852,N_19344,N_19128);
or U19853 (N_19853,N_19488,N_19448);
and U19854 (N_19854,N_19498,N_19092);
nand U19855 (N_19855,N_19385,N_19275);
nand U19856 (N_19856,N_19174,N_19460);
nor U19857 (N_19857,N_19294,N_19436);
and U19858 (N_19858,N_19155,N_19489);
or U19859 (N_19859,N_19456,N_19418);
or U19860 (N_19860,N_19135,N_19140);
nor U19861 (N_19861,N_19125,N_19293);
xor U19862 (N_19862,N_19137,N_19471);
nand U19863 (N_19863,N_19470,N_19282);
xnor U19864 (N_19864,N_19001,N_19000);
xnor U19865 (N_19865,N_19033,N_19008);
xnor U19866 (N_19866,N_19179,N_19069);
xor U19867 (N_19867,N_19089,N_19050);
and U19868 (N_19868,N_19210,N_19104);
or U19869 (N_19869,N_19411,N_19465);
nand U19870 (N_19870,N_19435,N_19108);
and U19871 (N_19871,N_19220,N_19242);
and U19872 (N_19872,N_19374,N_19330);
xor U19873 (N_19873,N_19487,N_19083);
and U19874 (N_19874,N_19157,N_19322);
xor U19875 (N_19875,N_19390,N_19289);
nor U19876 (N_19876,N_19175,N_19143);
nand U19877 (N_19877,N_19400,N_19390);
nand U19878 (N_19878,N_19129,N_19047);
nor U19879 (N_19879,N_19403,N_19170);
nor U19880 (N_19880,N_19212,N_19328);
xnor U19881 (N_19881,N_19293,N_19224);
and U19882 (N_19882,N_19411,N_19451);
nand U19883 (N_19883,N_19285,N_19302);
nand U19884 (N_19884,N_19110,N_19391);
or U19885 (N_19885,N_19123,N_19495);
xnor U19886 (N_19886,N_19319,N_19353);
xnor U19887 (N_19887,N_19446,N_19081);
or U19888 (N_19888,N_19089,N_19470);
and U19889 (N_19889,N_19189,N_19231);
nor U19890 (N_19890,N_19063,N_19471);
xnor U19891 (N_19891,N_19199,N_19112);
and U19892 (N_19892,N_19005,N_19165);
nand U19893 (N_19893,N_19010,N_19316);
or U19894 (N_19894,N_19334,N_19308);
nand U19895 (N_19895,N_19063,N_19427);
nor U19896 (N_19896,N_19270,N_19170);
xor U19897 (N_19897,N_19491,N_19172);
and U19898 (N_19898,N_19278,N_19078);
or U19899 (N_19899,N_19452,N_19379);
and U19900 (N_19900,N_19396,N_19387);
and U19901 (N_19901,N_19133,N_19037);
xnor U19902 (N_19902,N_19173,N_19275);
xnor U19903 (N_19903,N_19491,N_19210);
or U19904 (N_19904,N_19029,N_19085);
and U19905 (N_19905,N_19318,N_19368);
nor U19906 (N_19906,N_19213,N_19034);
nand U19907 (N_19907,N_19182,N_19476);
nand U19908 (N_19908,N_19258,N_19389);
nand U19909 (N_19909,N_19470,N_19173);
or U19910 (N_19910,N_19211,N_19479);
or U19911 (N_19911,N_19182,N_19152);
nand U19912 (N_19912,N_19489,N_19042);
or U19913 (N_19913,N_19039,N_19007);
nor U19914 (N_19914,N_19286,N_19340);
and U19915 (N_19915,N_19420,N_19113);
or U19916 (N_19916,N_19321,N_19121);
nor U19917 (N_19917,N_19386,N_19043);
xnor U19918 (N_19918,N_19150,N_19494);
or U19919 (N_19919,N_19024,N_19106);
xnor U19920 (N_19920,N_19317,N_19121);
xnor U19921 (N_19921,N_19448,N_19032);
nand U19922 (N_19922,N_19262,N_19012);
nor U19923 (N_19923,N_19158,N_19251);
xnor U19924 (N_19924,N_19457,N_19146);
and U19925 (N_19925,N_19217,N_19103);
or U19926 (N_19926,N_19024,N_19185);
xnor U19927 (N_19927,N_19393,N_19207);
or U19928 (N_19928,N_19192,N_19040);
and U19929 (N_19929,N_19463,N_19034);
and U19930 (N_19930,N_19477,N_19489);
nand U19931 (N_19931,N_19281,N_19250);
or U19932 (N_19932,N_19078,N_19335);
or U19933 (N_19933,N_19185,N_19265);
and U19934 (N_19934,N_19182,N_19418);
xnor U19935 (N_19935,N_19161,N_19353);
nor U19936 (N_19936,N_19013,N_19455);
xor U19937 (N_19937,N_19279,N_19397);
nor U19938 (N_19938,N_19168,N_19388);
and U19939 (N_19939,N_19163,N_19023);
nand U19940 (N_19940,N_19204,N_19396);
nand U19941 (N_19941,N_19182,N_19433);
nor U19942 (N_19942,N_19491,N_19085);
nand U19943 (N_19943,N_19049,N_19108);
or U19944 (N_19944,N_19112,N_19473);
and U19945 (N_19945,N_19289,N_19270);
xor U19946 (N_19946,N_19312,N_19059);
nor U19947 (N_19947,N_19237,N_19312);
and U19948 (N_19948,N_19198,N_19360);
nand U19949 (N_19949,N_19408,N_19061);
and U19950 (N_19950,N_19144,N_19254);
nor U19951 (N_19951,N_19456,N_19169);
nand U19952 (N_19952,N_19062,N_19363);
and U19953 (N_19953,N_19076,N_19092);
xor U19954 (N_19954,N_19436,N_19499);
and U19955 (N_19955,N_19487,N_19066);
nor U19956 (N_19956,N_19318,N_19063);
or U19957 (N_19957,N_19337,N_19120);
xor U19958 (N_19958,N_19438,N_19022);
xor U19959 (N_19959,N_19472,N_19374);
and U19960 (N_19960,N_19312,N_19378);
and U19961 (N_19961,N_19305,N_19292);
or U19962 (N_19962,N_19489,N_19370);
nor U19963 (N_19963,N_19376,N_19474);
and U19964 (N_19964,N_19046,N_19214);
xnor U19965 (N_19965,N_19266,N_19344);
xor U19966 (N_19966,N_19143,N_19099);
xor U19967 (N_19967,N_19435,N_19256);
xor U19968 (N_19968,N_19316,N_19286);
xor U19969 (N_19969,N_19210,N_19258);
or U19970 (N_19970,N_19168,N_19374);
and U19971 (N_19971,N_19474,N_19268);
nand U19972 (N_19972,N_19053,N_19160);
nand U19973 (N_19973,N_19151,N_19094);
nor U19974 (N_19974,N_19193,N_19410);
xor U19975 (N_19975,N_19334,N_19327);
and U19976 (N_19976,N_19043,N_19300);
or U19977 (N_19977,N_19163,N_19387);
xnor U19978 (N_19978,N_19196,N_19204);
nor U19979 (N_19979,N_19039,N_19048);
nand U19980 (N_19980,N_19305,N_19345);
nor U19981 (N_19981,N_19062,N_19082);
xor U19982 (N_19982,N_19320,N_19146);
xnor U19983 (N_19983,N_19340,N_19199);
nor U19984 (N_19984,N_19268,N_19222);
and U19985 (N_19985,N_19144,N_19330);
and U19986 (N_19986,N_19465,N_19155);
or U19987 (N_19987,N_19445,N_19344);
or U19988 (N_19988,N_19485,N_19090);
xor U19989 (N_19989,N_19108,N_19310);
or U19990 (N_19990,N_19276,N_19012);
or U19991 (N_19991,N_19432,N_19332);
or U19992 (N_19992,N_19149,N_19209);
nor U19993 (N_19993,N_19421,N_19087);
or U19994 (N_19994,N_19246,N_19336);
nand U19995 (N_19995,N_19472,N_19031);
or U19996 (N_19996,N_19351,N_19030);
and U19997 (N_19997,N_19307,N_19477);
nand U19998 (N_19998,N_19131,N_19037);
or U19999 (N_19999,N_19406,N_19440);
nand U20000 (N_20000,N_19921,N_19580);
nor U20001 (N_20001,N_19682,N_19694);
nand U20002 (N_20002,N_19613,N_19625);
xor U20003 (N_20003,N_19742,N_19574);
xor U20004 (N_20004,N_19610,N_19700);
nand U20005 (N_20005,N_19729,N_19759);
xor U20006 (N_20006,N_19588,N_19507);
nand U20007 (N_20007,N_19644,N_19581);
nand U20008 (N_20008,N_19643,N_19904);
nor U20009 (N_20009,N_19524,N_19878);
and U20010 (N_20010,N_19826,N_19672);
nand U20011 (N_20011,N_19774,N_19534);
nor U20012 (N_20012,N_19519,N_19992);
and U20013 (N_20013,N_19881,N_19535);
and U20014 (N_20014,N_19989,N_19693);
xor U20015 (N_20015,N_19523,N_19640);
or U20016 (N_20016,N_19834,N_19666);
or U20017 (N_20017,N_19938,N_19577);
nor U20018 (N_20018,N_19950,N_19751);
or U20019 (N_20019,N_19932,N_19976);
or U20020 (N_20020,N_19839,N_19600);
or U20021 (N_20021,N_19718,N_19847);
and U20022 (N_20022,N_19968,N_19850);
nand U20023 (N_20023,N_19629,N_19608);
nor U20024 (N_20024,N_19863,N_19925);
nand U20025 (N_20025,N_19645,N_19614);
and U20026 (N_20026,N_19884,N_19598);
and U20027 (N_20027,N_19855,N_19870);
or U20028 (N_20028,N_19628,N_19750);
nor U20029 (N_20029,N_19697,N_19810);
nand U20030 (N_20030,N_19698,N_19674);
and U20031 (N_20031,N_19997,N_19501);
nand U20032 (N_20032,N_19823,N_19967);
and U20033 (N_20033,N_19898,N_19673);
nand U20034 (N_20034,N_19707,N_19833);
and U20035 (N_20035,N_19579,N_19536);
nand U20036 (N_20036,N_19931,N_19618);
and U20037 (N_20037,N_19787,N_19566);
nor U20038 (N_20038,N_19948,N_19830);
or U20039 (N_20039,N_19602,N_19745);
xnor U20040 (N_20040,N_19746,N_19765);
and U20041 (N_20041,N_19680,N_19930);
and U20042 (N_20042,N_19763,N_19906);
and U20043 (N_20043,N_19996,N_19973);
or U20044 (N_20044,N_19514,N_19775);
nor U20045 (N_20045,N_19633,N_19892);
nor U20046 (N_20046,N_19962,N_19540);
and U20047 (N_20047,N_19651,N_19798);
or U20048 (N_20048,N_19549,N_19741);
nor U20049 (N_20049,N_19738,N_19840);
xor U20050 (N_20050,N_19846,N_19905);
and U20051 (N_20051,N_19772,N_19727);
nand U20052 (N_20052,N_19963,N_19732);
xnor U20053 (N_20053,N_19800,N_19734);
or U20054 (N_20054,N_19955,N_19939);
nand U20055 (N_20055,N_19736,N_19791);
nor U20056 (N_20056,N_19546,N_19530);
nor U20057 (N_20057,N_19564,N_19928);
xnor U20058 (N_20058,N_19735,N_19893);
xor U20059 (N_20059,N_19764,N_19533);
nand U20060 (N_20060,N_19794,N_19652);
nand U20061 (N_20061,N_19615,N_19896);
xnor U20062 (N_20062,N_19943,N_19937);
xnor U20063 (N_20063,N_19910,N_19824);
or U20064 (N_20064,N_19946,N_19703);
or U20065 (N_20065,N_19553,N_19808);
nor U20066 (N_20066,N_19785,N_19724);
or U20067 (N_20067,N_19781,N_19872);
nand U20068 (N_20068,N_19515,N_19873);
and U20069 (N_20069,N_19619,N_19758);
nand U20070 (N_20070,N_19941,N_19563);
xnor U20071 (N_20071,N_19934,N_19686);
nor U20072 (N_20072,N_19720,N_19717);
and U20073 (N_20073,N_19565,N_19874);
nor U20074 (N_20074,N_19531,N_19578);
or U20075 (N_20075,N_19829,N_19517);
nor U20076 (N_20076,N_19502,N_19656);
or U20077 (N_20077,N_19913,N_19803);
or U20078 (N_20078,N_19689,N_19518);
and U20079 (N_20079,N_19795,N_19940);
or U20080 (N_20080,N_19719,N_19599);
xor U20081 (N_20081,N_19877,N_19634);
nand U20082 (N_20082,N_19716,N_19711);
xnor U20083 (N_20083,N_19883,N_19835);
xor U20084 (N_20084,N_19594,N_19662);
and U20085 (N_20085,N_19899,N_19880);
or U20086 (N_20086,N_19709,N_19544);
or U20087 (N_20087,N_19504,N_19854);
or U20088 (N_20088,N_19861,N_19609);
xnor U20089 (N_20089,N_19942,N_19661);
nor U20090 (N_20090,N_19953,N_19918);
and U20091 (N_20091,N_19550,N_19744);
or U20092 (N_20092,N_19993,N_19538);
xor U20093 (N_20093,N_19516,N_19596);
or U20094 (N_20094,N_19995,N_19837);
nand U20095 (N_20095,N_19677,N_19797);
nor U20096 (N_20096,N_19556,N_19985);
or U20097 (N_20097,N_19575,N_19623);
and U20098 (N_20098,N_19617,N_19852);
nand U20099 (N_20099,N_19903,N_19585);
xnor U20100 (N_20100,N_19919,N_19676);
or U20101 (N_20101,N_19601,N_19739);
nand U20102 (N_20102,N_19767,N_19650);
and U20103 (N_20103,N_19554,N_19994);
nor U20104 (N_20104,N_19622,N_19859);
xor U20105 (N_20105,N_19844,N_19926);
and U20106 (N_20106,N_19635,N_19589);
and U20107 (N_20107,N_19522,N_19821);
nand U20108 (N_20108,N_19513,N_19587);
nand U20109 (N_20109,N_19804,N_19667);
nor U20110 (N_20110,N_19762,N_19604);
xnor U20111 (N_20111,N_19627,N_19961);
or U20112 (N_20112,N_19848,N_19512);
or U20113 (N_20113,N_19782,N_19867);
and U20114 (N_20114,N_19780,N_19971);
and U20115 (N_20115,N_19702,N_19648);
xor U20116 (N_20116,N_19528,N_19678);
and U20117 (N_20117,N_19778,N_19715);
or U20118 (N_20118,N_19789,N_19664);
xor U20119 (N_20119,N_19658,N_19974);
or U20120 (N_20120,N_19525,N_19561);
and U20121 (N_20121,N_19815,N_19558);
and U20122 (N_20122,N_19977,N_19595);
xnor U20123 (N_20123,N_19783,N_19721);
nor U20124 (N_20124,N_19593,N_19584);
and U20125 (N_20125,N_19510,N_19777);
nand U20126 (N_20126,N_19935,N_19799);
nor U20127 (N_20127,N_19814,N_19802);
nor U20128 (N_20128,N_19722,N_19966);
and U20129 (N_20129,N_19914,N_19969);
nand U20130 (N_20130,N_19527,N_19590);
and U20131 (N_20131,N_19813,N_19889);
and U20132 (N_20132,N_19675,N_19944);
xor U20133 (N_20133,N_19954,N_19555);
and U20134 (N_20134,N_19760,N_19624);
nor U20135 (N_20135,N_19552,N_19822);
nor U20136 (N_20136,N_19503,N_19696);
and U20137 (N_20137,N_19856,N_19568);
or U20138 (N_20138,N_19621,N_19509);
xor U20139 (N_20139,N_19894,N_19607);
xor U20140 (N_20140,N_19838,N_19790);
and U20141 (N_20141,N_19888,N_19690);
nand U20142 (N_20142,N_19999,N_19740);
or U20143 (N_20143,N_19979,N_19957);
xor U20144 (N_20144,N_19557,N_19987);
xnor U20145 (N_20145,N_19978,N_19537);
nor U20146 (N_20146,N_19816,N_19529);
nand U20147 (N_20147,N_19630,N_19573);
nand U20148 (N_20148,N_19638,N_19920);
xor U20149 (N_20149,N_19520,N_19982);
and U20150 (N_20150,N_19949,N_19890);
xnor U20151 (N_20151,N_19769,N_19965);
and U20152 (N_20152,N_19924,N_19761);
and U20153 (N_20153,N_19917,N_19646);
xnor U20154 (N_20154,N_19655,N_19901);
nor U20155 (N_20155,N_19879,N_19909);
or U20156 (N_20156,N_19701,N_19688);
xnor U20157 (N_20157,N_19842,N_19784);
or U20158 (N_20158,N_19811,N_19508);
and U20159 (N_20159,N_19947,N_19768);
and U20160 (N_20160,N_19752,N_19548);
and U20161 (N_20161,N_19730,N_19773);
or U20162 (N_20162,N_19659,N_19684);
nor U20163 (N_20163,N_19706,N_19642);
or U20164 (N_20164,N_19869,N_19860);
nor U20165 (N_20165,N_19572,N_19828);
xor U20166 (N_20166,N_19704,N_19737);
or U20167 (N_20167,N_19731,N_19970);
xnor U20168 (N_20168,N_19505,N_19900);
and U20169 (N_20169,N_19858,N_19866);
xnor U20170 (N_20170,N_19851,N_19923);
nand U20171 (N_20171,N_19886,N_19521);
nand U20172 (N_20172,N_19868,N_19776);
or U20173 (N_20173,N_19660,N_19766);
xor U20174 (N_20174,N_19733,N_19639);
and U20175 (N_20175,N_19984,N_19543);
nand U20176 (N_20176,N_19862,N_19567);
or U20177 (N_20177,N_19857,N_19951);
or U20178 (N_20178,N_19705,N_19532);
xnor U20179 (N_20179,N_19849,N_19807);
or U20180 (N_20180,N_19668,N_19649);
and U20181 (N_20181,N_19865,N_19959);
xor U20182 (N_20182,N_19753,N_19831);
or U20183 (N_20183,N_19853,N_19685);
xor U20184 (N_20184,N_19818,N_19990);
xor U20185 (N_20185,N_19713,N_19771);
or U20186 (N_20186,N_19972,N_19864);
and U20187 (N_20187,N_19841,N_19796);
nor U20188 (N_20188,N_19755,N_19571);
nand U20189 (N_20189,N_19551,N_19945);
nand U20190 (N_20190,N_19933,N_19506);
nor U20191 (N_20191,N_19562,N_19975);
nand U20192 (N_20192,N_19569,N_19812);
or U20193 (N_20193,N_19541,N_19631);
nand U20194 (N_20194,N_19936,N_19952);
nor U20195 (N_20195,N_19699,N_19606);
nand U20196 (N_20196,N_19788,N_19809);
xor U20197 (N_20197,N_19981,N_19725);
or U20198 (N_20198,N_19681,N_19980);
xor U20199 (N_20199,N_19756,N_19641);
nand U20200 (N_20200,N_19902,N_19582);
or U20201 (N_20201,N_19597,N_19805);
xnor U20202 (N_20202,N_19747,N_19960);
xor U20203 (N_20203,N_19882,N_19875);
nand U20204 (N_20204,N_19576,N_19793);
xnor U20205 (N_20205,N_19620,N_19691);
nor U20206 (N_20206,N_19876,N_19526);
nand U20207 (N_20207,N_19647,N_19632);
or U20208 (N_20208,N_19726,N_19922);
nand U20209 (N_20209,N_19583,N_19636);
nand U20210 (N_20210,N_19912,N_19511);
or U20211 (N_20211,N_19885,N_19806);
and U20212 (N_20212,N_19670,N_19908);
or U20213 (N_20213,N_19836,N_19687);
nand U20214 (N_20214,N_19657,N_19605);
and U20215 (N_20215,N_19907,N_19916);
nor U20216 (N_20216,N_19845,N_19714);
nor U20217 (N_20217,N_19637,N_19539);
and U20218 (N_20218,N_19871,N_19786);
nand U20219 (N_20219,N_19710,N_19895);
nor U20220 (N_20220,N_19983,N_19779);
nand U20221 (N_20221,N_19591,N_19559);
nand U20222 (N_20222,N_19542,N_19956);
nor U20223 (N_20223,N_19665,N_19728);
and U20224 (N_20224,N_19692,N_19891);
nand U20225 (N_20225,N_19825,N_19911);
and U20226 (N_20226,N_19832,N_19998);
nor U20227 (N_20227,N_19723,N_19757);
and U20228 (N_20228,N_19683,N_19801);
nand U20229 (N_20229,N_19749,N_19929);
nand U20230 (N_20230,N_19663,N_19560);
or U20231 (N_20231,N_19586,N_19991);
nand U20232 (N_20232,N_19827,N_19770);
xnor U20233 (N_20233,N_19915,N_19669);
nand U20234 (N_20234,N_19592,N_19708);
xnor U20235 (N_20235,N_19653,N_19695);
nor U20236 (N_20236,N_19626,N_19988);
nor U20237 (N_20237,N_19612,N_19817);
xor U20238 (N_20238,N_19671,N_19819);
nand U20239 (N_20239,N_19820,N_19611);
and U20240 (N_20240,N_19743,N_19843);
xnor U20241 (N_20241,N_19792,N_19748);
xor U20242 (N_20242,N_19958,N_19712);
or U20243 (N_20243,N_19679,N_19754);
xor U20244 (N_20244,N_19986,N_19570);
nor U20245 (N_20245,N_19616,N_19897);
xnor U20246 (N_20246,N_19887,N_19545);
and U20247 (N_20247,N_19927,N_19603);
or U20248 (N_20248,N_19654,N_19964);
or U20249 (N_20249,N_19547,N_19500);
nand U20250 (N_20250,N_19914,N_19978);
nor U20251 (N_20251,N_19873,N_19947);
and U20252 (N_20252,N_19934,N_19609);
and U20253 (N_20253,N_19760,N_19918);
nor U20254 (N_20254,N_19632,N_19579);
and U20255 (N_20255,N_19863,N_19972);
nor U20256 (N_20256,N_19686,N_19972);
xor U20257 (N_20257,N_19541,N_19854);
xnor U20258 (N_20258,N_19636,N_19685);
xor U20259 (N_20259,N_19598,N_19713);
and U20260 (N_20260,N_19677,N_19770);
nand U20261 (N_20261,N_19518,N_19884);
nor U20262 (N_20262,N_19743,N_19989);
nand U20263 (N_20263,N_19812,N_19772);
xor U20264 (N_20264,N_19952,N_19614);
xnor U20265 (N_20265,N_19805,N_19534);
nand U20266 (N_20266,N_19782,N_19633);
and U20267 (N_20267,N_19571,N_19808);
or U20268 (N_20268,N_19781,N_19624);
and U20269 (N_20269,N_19643,N_19804);
nor U20270 (N_20270,N_19639,N_19738);
or U20271 (N_20271,N_19935,N_19990);
xnor U20272 (N_20272,N_19959,N_19937);
xor U20273 (N_20273,N_19918,N_19735);
and U20274 (N_20274,N_19799,N_19740);
nor U20275 (N_20275,N_19832,N_19811);
and U20276 (N_20276,N_19550,N_19573);
xnor U20277 (N_20277,N_19745,N_19633);
nand U20278 (N_20278,N_19596,N_19897);
or U20279 (N_20279,N_19878,N_19922);
xor U20280 (N_20280,N_19541,N_19600);
xor U20281 (N_20281,N_19793,N_19950);
xor U20282 (N_20282,N_19595,N_19708);
nor U20283 (N_20283,N_19771,N_19862);
xnor U20284 (N_20284,N_19508,N_19785);
nand U20285 (N_20285,N_19946,N_19870);
or U20286 (N_20286,N_19828,N_19519);
or U20287 (N_20287,N_19876,N_19901);
xnor U20288 (N_20288,N_19609,N_19802);
and U20289 (N_20289,N_19531,N_19961);
or U20290 (N_20290,N_19553,N_19961);
nor U20291 (N_20291,N_19652,N_19757);
and U20292 (N_20292,N_19779,N_19722);
or U20293 (N_20293,N_19551,N_19858);
nor U20294 (N_20294,N_19924,N_19845);
nand U20295 (N_20295,N_19708,N_19905);
or U20296 (N_20296,N_19837,N_19721);
and U20297 (N_20297,N_19883,N_19599);
and U20298 (N_20298,N_19500,N_19920);
and U20299 (N_20299,N_19966,N_19565);
nor U20300 (N_20300,N_19657,N_19802);
and U20301 (N_20301,N_19711,N_19878);
xnor U20302 (N_20302,N_19747,N_19804);
xor U20303 (N_20303,N_19690,N_19531);
nand U20304 (N_20304,N_19536,N_19535);
or U20305 (N_20305,N_19759,N_19850);
xor U20306 (N_20306,N_19758,N_19637);
xnor U20307 (N_20307,N_19548,N_19713);
and U20308 (N_20308,N_19867,N_19675);
nand U20309 (N_20309,N_19865,N_19947);
nand U20310 (N_20310,N_19534,N_19710);
and U20311 (N_20311,N_19637,N_19942);
and U20312 (N_20312,N_19614,N_19595);
and U20313 (N_20313,N_19925,N_19689);
nand U20314 (N_20314,N_19769,N_19827);
or U20315 (N_20315,N_19727,N_19687);
and U20316 (N_20316,N_19509,N_19681);
nor U20317 (N_20317,N_19833,N_19966);
and U20318 (N_20318,N_19779,N_19780);
xor U20319 (N_20319,N_19661,N_19508);
or U20320 (N_20320,N_19760,N_19554);
or U20321 (N_20321,N_19863,N_19677);
nor U20322 (N_20322,N_19696,N_19569);
nand U20323 (N_20323,N_19704,N_19528);
xnor U20324 (N_20324,N_19561,N_19537);
or U20325 (N_20325,N_19909,N_19586);
or U20326 (N_20326,N_19922,N_19690);
nor U20327 (N_20327,N_19603,N_19954);
and U20328 (N_20328,N_19662,N_19844);
xor U20329 (N_20329,N_19762,N_19848);
or U20330 (N_20330,N_19509,N_19688);
and U20331 (N_20331,N_19752,N_19845);
nor U20332 (N_20332,N_19546,N_19793);
and U20333 (N_20333,N_19552,N_19652);
nor U20334 (N_20334,N_19751,N_19629);
and U20335 (N_20335,N_19914,N_19825);
and U20336 (N_20336,N_19563,N_19967);
and U20337 (N_20337,N_19889,N_19896);
nand U20338 (N_20338,N_19744,N_19527);
nor U20339 (N_20339,N_19810,N_19657);
or U20340 (N_20340,N_19570,N_19715);
nor U20341 (N_20341,N_19812,N_19976);
xor U20342 (N_20342,N_19743,N_19927);
nor U20343 (N_20343,N_19899,N_19705);
nand U20344 (N_20344,N_19807,N_19605);
or U20345 (N_20345,N_19739,N_19808);
nor U20346 (N_20346,N_19727,N_19942);
xnor U20347 (N_20347,N_19603,N_19884);
and U20348 (N_20348,N_19823,N_19507);
nand U20349 (N_20349,N_19809,N_19683);
or U20350 (N_20350,N_19901,N_19895);
nor U20351 (N_20351,N_19787,N_19632);
xnor U20352 (N_20352,N_19753,N_19593);
nand U20353 (N_20353,N_19629,N_19528);
nand U20354 (N_20354,N_19734,N_19727);
nor U20355 (N_20355,N_19538,N_19596);
or U20356 (N_20356,N_19819,N_19640);
or U20357 (N_20357,N_19745,N_19845);
or U20358 (N_20358,N_19535,N_19798);
and U20359 (N_20359,N_19795,N_19843);
and U20360 (N_20360,N_19607,N_19754);
nand U20361 (N_20361,N_19702,N_19503);
and U20362 (N_20362,N_19833,N_19577);
xor U20363 (N_20363,N_19558,N_19835);
nor U20364 (N_20364,N_19825,N_19554);
and U20365 (N_20365,N_19686,N_19616);
nand U20366 (N_20366,N_19929,N_19676);
xor U20367 (N_20367,N_19548,N_19639);
and U20368 (N_20368,N_19622,N_19647);
nand U20369 (N_20369,N_19655,N_19873);
xnor U20370 (N_20370,N_19602,N_19673);
nor U20371 (N_20371,N_19992,N_19550);
or U20372 (N_20372,N_19757,N_19738);
nor U20373 (N_20373,N_19584,N_19994);
or U20374 (N_20374,N_19932,N_19660);
xnor U20375 (N_20375,N_19709,N_19814);
or U20376 (N_20376,N_19538,N_19700);
nand U20377 (N_20377,N_19752,N_19549);
nand U20378 (N_20378,N_19858,N_19910);
and U20379 (N_20379,N_19668,N_19841);
nor U20380 (N_20380,N_19909,N_19804);
nor U20381 (N_20381,N_19617,N_19803);
or U20382 (N_20382,N_19595,N_19761);
xor U20383 (N_20383,N_19965,N_19542);
nand U20384 (N_20384,N_19540,N_19568);
or U20385 (N_20385,N_19978,N_19915);
nor U20386 (N_20386,N_19788,N_19760);
xor U20387 (N_20387,N_19632,N_19580);
nor U20388 (N_20388,N_19791,N_19504);
xor U20389 (N_20389,N_19669,N_19646);
or U20390 (N_20390,N_19764,N_19571);
xor U20391 (N_20391,N_19764,N_19705);
or U20392 (N_20392,N_19962,N_19821);
nor U20393 (N_20393,N_19992,N_19754);
or U20394 (N_20394,N_19889,N_19807);
xor U20395 (N_20395,N_19764,N_19546);
nor U20396 (N_20396,N_19559,N_19976);
and U20397 (N_20397,N_19803,N_19873);
nor U20398 (N_20398,N_19751,N_19768);
xnor U20399 (N_20399,N_19982,N_19989);
nand U20400 (N_20400,N_19536,N_19547);
and U20401 (N_20401,N_19755,N_19861);
or U20402 (N_20402,N_19775,N_19969);
and U20403 (N_20403,N_19835,N_19796);
nor U20404 (N_20404,N_19692,N_19903);
nand U20405 (N_20405,N_19631,N_19734);
nand U20406 (N_20406,N_19692,N_19748);
xnor U20407 (N_20407,N_19586,N_19911);
nor U20408 (N_20408,N_19709,N_19736);
nor U20409 (N_20409,N_19642,N_19995);
nand U20410 (N_20410,N_19785,N_19964);
nor U20411 (N_20411,N_19757,N_19688);
or U20412 (N_20412,N_19569,N_19994);
and U20413 (N_20413,N_19674,N_19978);
and U20414 (N_20414,N_19881,N_19742);
nor U20415 (N_20415,N_19781,N_19635);
xor U20416 (N_20416,N_19762,N_19889);
and U20417 (N_20417,N_19675,N_19880);
xor U20418 (N_20418,N_19685,N_19890);
xnor U20419 (N_20419,N_19729,N_19632);
or U20420 (N_20420,N_19927,N_19800);
xor U20421 (N_20421,N_19837,N_19974);
nand U20422 (N_20422,N_19952,N_19872);
xor U20423 (N_20423,N_19898,N_19574);
xor U20424 (N_20424,N_19699,N_19907);
xor U20425 (N_20425,N_19709,N_19515);
nand U20426 (N_20426,N_19559,N_19713);
or U20427 (N_20427,N_19686,N_19834);
nor U20428 (N_20428,N_19858,N_19783);
or U20429 (N_20429,N_19516,N_19861);
nor U20430 (N_20430,N_19819,N_19972);
xnor U20431 (N_20431,N_19668,N_19672);
nand U20432 (N_20432,N_19910,N_19646);
nor U20433 (N_20433,N_19958,N_19999);
nand U20434 (N_20434,N_19975,N_19570);
nand U20435 (N_20435,N_19851,N_19675);
and U20436 (N_20436,N_19646,N_19512);
xnor U20437 (N_20437,N_19591,N_19712);
or U20438 (N_20438,N_19780,N_19838);
or U20439 (N_20439,N_19517,N_19846);
or U20440 (N_20440,N_19508,N_19606);
nor U20441 (N_20441,N_19543,N_19909);
nor U20442 (N_20442,N_19708,N_19594);
nand U20443 (N_20443,N_19564,N_19996);
nand U20444 (N_20444,N_19727,N_19704);
and U20445 (N_20445,N_19880,N_19808);
nand U20446 (N_20446,N_19874,N_19767);
xor U20447 (N_20447,N_19878,N_19706);
and U20448 (N_20448,N_19626,N_19517);
and U20449 (N_20449,N_19763,N_19540);
and U20450 (N_20450,N_19902,N_19719);
nor U20451 (N_20451,N_19611,N_19711);
or U20452 (N_20452,N_19559,N_19630);
nor U20453 (N_20453,N_19668,N_19582);
or U20454 (N_20454,N_19777,N_19582);
and U20455 (N_20455,N_19595,N_19747);
and U20456 (N_20456,N_19792,N_19969);
or U20457 (N_20457,N_19527,N_19936);
nand U20458 (N_20458,N_19965,N_19986);
xnor U20459 (N_20459,N_19731,N_19626);
nor U20460 (N_20460,N_19802,N_19989);
or U20461 (N_20461,N_19511,N_19909);
or U20462 (N_20462,N_19592,N_19580);
xor U20463 (N_20463,N_19953,N_19999);
nor U20464 (N_20464,N_19614,N_19600);
and U20465 (N_20465,N_19827,N_19686);
and U20466 (N_20466,N_19682,N_19502);
or U20467 (N_20467,N_19815,N_19871);
or U20468 (N_20468,N_19949,N_19595);
or U20469 (N_20469,N_19789,N_19666);
and U20470 (N_20470,N_19978,N_19755);
nor U20471 (N_20471,N_19793,N_19672);
xnor U20472 (N_20472,N_19595,N_19607);
or U20473 (N_20473,N_19771,N_19988);
and U20474 (N_20474,N_19869,N_19852);
nand U20475 (N_20475,N_19763,N_19689);
nand U20476 (N_20476,N_19545,N_19896);
and U20477 (N_20477,N_19546,N_19758);
or U20478 (N_20478,N_19793,N_19956);
xor U20479 (N_20479,N_19697,N_19658);
xor U20480 (N_20480,N_19740,N_19861);
nand U20481 (N_20481,N_19987,N_19522);
nand U20482 (N_20482,N_19662,N_19751);
and U20483 (N_20483,N_19896,N_19587);
xnor U20484 (N_20484,N_19829,N_19993);
xor U20485 (N_20485,N_19962,N_19819);
nor U20486 (N_20486,N_19610,N_19671);
or U20487 (N_20487,N_19841,N_19956);
xnor U20488 (N_20488,N_19824,N_19570);
or U20489 (N_20489,N_19503,N_19547);
xor U20490 (N_20490,N_19941,N_19681);
nand U20491 (N_20491,N_19740,N_19769);
xor U20492 (N_20492,N_19666,N_19758);
or U20493 (N_20493,N_19522,N_19806);
and U20494 (N_20494,N_19709,N_19779);
nand U20495 (N_20495,N_19582,N_19745);
nor U20496 (N_20496,N_19633,N_19922);
and U20497 (N_20497,N_19701,N_19617);
or U20498 (N_20498,N_19942,N_19579);
xor U20499 (N_20499,N_19855,N_19816);
xnor U20500 (N_20500,N_20477,N_20103);
nand U20501 (N_20501,N_20450,N_20136);
or U20502 (N_20502,N_20098,N_20027);
nand U20503 (N_20503,N_20161,N_20411);
nor U20504 (N_20504,N_20359,N_20169);
and U20505 (N_20505,N_20300,N_20171);
nand U20506 (N_20506,N_20280,N_20270);
nor U20507 (N_20507,N_20099,N_20260);
or U20508 (N_20508,N_20019,N_20256);
nand U20509 (N_20509,N_20251,N_20250);
nand U20510 (N_20510,N_20034,N_20229);
nor U20511 (N_20511,N_20274,N_20425);
nor U20512 (N_20512,N_20129,N_20088);
xor U20513 (N_20513,N_20339,N_20015);
nor U20514 (N_20514,N_20388,N_20165);
or U20515 (N_20515,N_20228,N_20493);
nand U20516 (N_20516,N_20231,N_20266);
nor U20517 (N_20517,N_20175,N_20148);
nor U20518 (N_20518,N_20041,N_20211);
xor U20519 (N_20519,N_20361,N_20018);
nand U20520 (N_20520,N_20310,N_20456);
nor U20521 (N_20521,N_20417,N_20068);
nor U20522 (N_20522,N_20268,N_20030);
nor U20523 (N_20523,N_20439,N_20091);
or U20524 (N_20524,N_20010,N_20090);
and U20525 (N_20525,N_20447,N_20024);
and U20526 (N_20526,N_20055,N_20047);
xnor U20527 (N_20527,N_20150,N_20200);
or U20528 (N_20528,N_20466,N_20126);
nor U20529 (N_20529,N_20470,N_20420);
and U20530 (N_20530,N_20037,N_20213);
nand U20531 (N_20531,N_20315,N_20014);
xor U20532 (N_20532,N_20166,N_20180);
nand U20533 (N_20533,N_20288,N_20051);
and U20534 (N_20534,N_20155,N_20490);
nor U20535 (N_20535,N_20192,N_20414);
nor U20536 (N_20536,N_20040,N_20328);
nor U20537 (N_20537,N_20065,N_20341);
xnor U20538 (N_20538,N_20354,N_20246);
and U20539 (N_20539,N_20120,N_20327);
nand U20540 (N_20540,N_20061,N_20198);
and U20541 (N_20541,N_20272,N_20356);
xnor U20542 (N_20542,N_20436,N_20471);
nor U20543 (N_20543,N_20386,N_20381);
or U20544 (N_20544,N_20087,N_20431);
and U20545 (N_20545,N_20304,N_20483);
and U20546 (N_20546,N_20033,N_20344);
nor U20547 (N_20547,N_20162,N_20348);
and U20548 (N_20548,N_20465,N_20476);
nor U20549 (N_20549,N_20028,N_20285);
xor U20550 (N_20550,N_20102,N_20371);
or U20551 (N_20551,N_20006,N_20408);
xor U20552 (N_20552,N_20392,N_20404);
nand U20553 (N_20553,N_20253,N_20212);
and U20554 (N_20554,N_20054,N_20009);
nor U20555 (N_20555,N_20105,N_20400);
xnor U20556 (N_20556,N_20275,N_20096);
xor U20557 (N_20557,N_20311,N_20022);
nand U20558 (N_20558,N_20355,N_20457);
nor U20559 (N_20559,N_20294,N_20295);
xnor U20560 (N_20560,N_20316,N_20084);
nor U20561 (N_20561,N_20445,N_20340);
xnor U20562 (N_20562,N_20230,N_20458);
xor U20563 (N_20563,N_20049,N_20403);
or U20564 (N_20564,N_20263,N_20209);
nor U20565 (N_20565,N_20062,N_20043);
nand U20566 (N_20566,N_20397,N_20455);
and U20567 (N_20567,N_20303,N_20244);
or U20568 (N_20568,N_20208,N_20410);
xnor U20569 (N_20569,N_20261,N_20132);
nand U20570 (N_20570,N_20170,N_20324);
or U20571 (N_20571,N_20100,N_20462);
and U20572 (N_20572,N_20469,N_20013);
xnor U20573 (N_20573,N_20191,N_20226);
xor U20574 (N_20574,N_20196,N_20485);
and U20575 (N_20575,N_20207,N_20215);
nor U20576 (N_20576,N_20484,N_20265);
nor U20577 (N_20577,N_20038,N_20432);
nor U20578 (N_20578,N_20117,N_20202);
nor U20579 (N_20579,N_20454,N_20326);
xor U20580 (N_20580,N_20337,N_20141);
and U20581 (N_20581,N_20112,N_20488);
or U20582 (N_20582,N_20017,N_20314);
or U20583 (N_20583,N_20377,N_20107);
xor U20584 (N_20584,N_20056,N_20044);
or U20585 (N_20585,N_20448,N_20080);
nor U20586 (N_20586,N_20104,N_20463);
xor U20587 (N_20587,N_20159,N_20323);
and U20588 (N_20588,N_20384,N_20429);
and U20589 (N_20589,N_20093,N_20154);
xnor U20590 (N_20590,N_20183,N_20446);
nor U20591 (N_20591,N_20139,N_20168);
or U20592 (N_20592,N_20347,N_20216);
or U20593 (N_20593,N_20157,N_20428);
and U20594 (N_20594,N_20186,N_20110);
nor U20595 (N_20595,N_20444,N_20077);
xnor U20596 (N_20596,N_20299,N_20172);
nand U20597 (N_20597,N_20057,N_20050);
and U20598 (N_20598,N_20421,N_20357);
nor U20599 (N_20599,N_20293,N_20188);
xnor U20600 (N_20600,N_20368,N_20369);
nand U20601 (N_20601,N_20343,N_20245);
nand U20602 (N_20602,N_20453,N_20438);
nor U20603 (N_20603,N_20257,N_20320);
nand U20604 (N_20604,N_20284,N_20273);
nand U20605 (N_20605,N_20002,N_20423);
nand U20606 (N_20606,N_20309,N_20204);
nor U20607 (N_20607,N_20407,N_20427);
nor U20608 (N_20608,N_20474,N_20193);
nor U20609 (N_20609,N_20335,N_20351);
and U20610 (N_20610,N_20406,N_20482);
or U20611 (N_20611,N_20382,N_20296);
and U20612 (N_20612,N_20277,N_20243);
nor U20613 (N_20613,N_20353,N_20074);
nor U20614 (N_20614,N_20064,N_20233);
and U20615 (N_20615,N_20185,N_20005);
and U20616 (N_20616,N_20402,N_20021);
nor U20617 (N_20617,N_20116,N_20012);
or U20618 (N_20618,N_20391,N_20398);
and U20619 (N_20619,N_20362,N_20127);
and U20620 (N_20620,N_20366,N_20210);
and U20621 (N_20621,N_20472,N_20237);
nor U20622 (N_20622,N_20312,N_20473);
nor U20623 (N_20623,N_20415,N_20241);
nand U20624 (N_20624,N_20158,N_20345);
nand U20625 (N_20625,N_20152,N_20329);
xor U20626 (N_20626,N_20167,N_20094);
nand U20627 (N_20627,N_20205,N_20184);
or U20628 (N_20628,N_20258,N_20111);
and U20629 (N_20629,N_20060,N_20292);
and U20630 (N_20630,N_20058,N_20222);
and U20631 (N_20631,N_20481,N_20071);
and U20632 (N_20632,N_20045,N_20433);
xnor U20633 (N_20633,N_20011,N_20332);
nor U20634 (N_20634,N_20114,N_20480);
nor U20635 (N_20635,N_20350,N_20418);
or U20636 (N_20636,N_20199,N_20026);
or U20637 (N_20637,N_20160,N_20372);
xor U20638 (N_20638,N_20413,N_20264);
nand U20639 (N_20639,N_20016,N_20422);
nand U20640 (N_20640,N_20187,N_20365);
or U20641 (N_20641,N_20426,N_20236);
xor U20642 (N_20642,N_20254,N_20346);
or U20643 (N_20643,N_20048,N_20489);
nand U20644 (N_20644,N_20467,N_20118);
and U20645 (N_20645,N_20281,N_20240);
and U20646 (N_20646,N_20452,N_20036);
nor U20647 (N_20647,N_20029,N_20072);
or U20648 (N_20648,N_20302,N_20238);
xor U20649 (N_20649,N_20321,N_20135);
nor U20650 (N_20650,N_20478,N_20227);
nand U20651 (N_20651,N_20079,N_20374);
or U20652 (N_20652,N_20387,N_20095);
nand U20653 (N_20653,N_20283,N_20106);
and U20654 (N_20654,N_20066,N_20499);
and U20655 (N_20655,N_20308,N_20318);
and U20656 (N_20656,N_20442,N_20086);
or U20657 (N_20657,N_20247,N_20435);
nand U20658 (N_20658,N_20333,N_20130);
xor U20659 (N_20659,N_20430,N_20486);
xor U20660 (N_20660,N_20075,N_20214);
or U20661 (N_20661,N_20195,N_20449);
or U20662 (N_20662,N_20437,N_20182);
xor U20663 (N_20663,N_20405,N_20298);
nand U20664 (N_20664,N_20317,N_20242);
nor U20665 (N_20665,N_20078,N_20031);
nor U20666 (N_20666,N_20225,N_20234);
nor U20667 (N_20667,N_20137,N_20451);
and U20668 (N_20668,N_20443,N_20142);
nand U20669 (N_20669,N_20069,N_20239);
nand U20670 (N_20670,N_20330,N_20495);
or U20671 (N_20671,N_20334,N_20460);
and U20672 (N_20672,N_20046,N_20390);
nand U20673 (N_20673,N_20143,N_20101);
nor U20674 (N_20674,N_20032,N_20279);
or U20675 (N_20675,N_20306,N_20189);
nand U20676 (N_20676,N_20115,N_20434);
or U20677 (N_20677,N_20349,N_20221);
nor U20678 (N_20678,N_20395,N_20206);
nand U20679 (N_20679,N_20367,N_20140);
or U20680 (N_20680,N_20151,N_20201);
nand U20681 (N_20681,N_20352,N_20370);
nor U20682 (N_20682,N_20396,N_20394);
nor U20683 (N_20683,N_20385,N_20059);
and U20684 (N_20684,N_20203,N_20393);
and U20685 (N_20685,N_20149,N_20085);
and U20686 (N_20686,N_20378,N_20389);
xor U20687 (N_20687,N_20262,N_20379);
nor U20688 (N_20688,N_20305,N_20479);
nand U20689 (N_20689,N_20419,N_20290);
or U20690 (N_20690,N_20138,N_20287);
or U20691 (N_20691,N_20178,N_20122);
nand U20692 (N_20692,N_20125,N_20089);
or U20693 (N_20693,N_20163,N_20492);
or U20694 (N_20694,N_20383,N_20409);
xnor U20695 (N_20695,N_20124,N_20399);
or U20696 (N_20696,N_20267,N_20291);
nor U20697 (N_20697,N_20363,N_20174);
or U20698 (N_20698,N_20301,N_20487);
or U20699 (N_20699,N_20235,N_20416);
xnor U20700 (N_20700,N_20176,N_20042);
xnor U20701 (N_20701,N_20373,N_20271);
or U20702 (N_20702,N_20092,N_20109);
nor U20703 (N_20703,N_20255,N_20123);
or U20704 (N_20704,N_20082,N_20156);
and U20705 (N_20705,N_20494,N_20322);
or U20706 (N_20706,N_20083,N_20121);
xnor U20707 (N_20707,N_20146,N_20338);
or U20708 (N_20708,N_20220,N_20496);
xor U20709 (N_20709,N_20342,N_20219);
or U20710 (N_20710,N_20181,N_20025);
nor U20711 (N_20711,N_20217,N_20003);
xnor U20712 (N_20712,N_20197,N_20440);
nor U20713 (N_20713,N_20259,N_20194);
nor U20714 (N_20714,N_20459,N_20461);
or U20715 (N_20715,N_20424,N_20375);
xor U20716 (N_20716,N_20224,N_20076);
xnor U20717 (N_20717,N_20053,N_20008);
nor U20718 (N_20718,N_20313,N_20131);
or U20719 (N_20719,N_20498,N_20286);
nor U20720 (N_20720,N_20052,N_20358);
nand U20721 (N_20721,N_20007,N_20232);
xnor U20722 (N_20722,N_20113,N_20468);
nand U20723 (N_20723,N_20223,N_20278);
and U20724 (N_20724,N_20081,N_20153);
or U20725 (N_20725,N_20000,N_20020);
nand U20726 (N_20726,N_20289,N_20401);
nand U20727 (N_20727,N_20412,N_20164);
nand U20728 (N_20728,N_20475,N_20179);
xor U20729 (N_20729,N_20147,N_20380);
and U20730 (N_20730,N_20108,N_20360);
xnor U20731 (N_20731,N_20190,N_20023);
xor U20732 (N_20732,N_20269,N_20464);
or U20733 (N_20733,N_20177,N_20144);
nand U20734 (N_20734,N_20249,N_20491);
nor U20735 (N_20735,N_20070,N_20119);
and U20736 (N_20736,N_20276,N_20001);
and U20737 (N_20737,N_20039,N_20297);
or U20738 (N_20738,N_20376,N_20325);
nand U20739 (N_20739,N_20441,N_20035);
nand U20740 (N_20740,N_20173,N_20145);
and U20741 (N_20741,N_20004,N_20336);
nor U20742 (N_20742,N_20134,N_20307);
nor U20743 (N_20743,N_20248,N_20497);
nand U20744 (N_20744,N_20252,N_20133);
and U20745 (N_20745,N_20282,N_20128);
or U20746 (N_20746,N_20073,N_20364);
xor U20747 (N_20747,N_20319,N_20218);
nor U20748 (N_20748,N_20331,N_20097);
nand U20749 (N_20749,N_20067,N_20063);
nor U20750 (N_20750,N_20125,N_20186);
xor U20751 (N_20751,N_20199,N_20268);
xor U20752 (N_20752,N_20406,N_20088);
nand U20753 (N_20753,N_20230,N_20143);
and U20754 (N_20754,N_20022,N_20225);
or U20755 (N_20755,N_20450,N_20343);
xnor U20756 (N_20756,N_20111,N_20164);
xnor U20757 (N_20757,N_20123,N_20192);
or U20758 (N_20758,N_20369,N_20442);
or U20759 (N_20759,N_20019,N_20421);
and U20760 (N_20760,N_20331,N_20069);
xor U20761 (N_20761,N_20225,N_20431);
and U20762 (N_20762,N_20206,N_20239);
nand U20763 (N_20763,N_20033,N_20232);
xor U20764 (N_20764,N_20151,N_20103);
nand U20765 (N_20765,N_20436,N_20237);
nand U20766 (N_20766,N_20001,N_20124);
nand U20767 (N_20767,N_20181,N_20428);
nand U20768 (N_20768,N_20002,N_20474);
and U20769 (N_20769,N_20096,N_20427);
and U20770 (N_20770,N_20178,N_20143);
and U20771 (N_20771,N_20497,N_20361);
xor U20772 (N_20772,N_20081,N_20050);
nand U20773 (N_20773,N_20476,N_20234);
nand U20774 (N_20774,N_20063,N_20274);
or U20775 (N_20775,N_20071,N_20060);
xnor U20776 (N_20776,N_20484,N_20427);
xnor U20777 (N_20777,N_20157,N_20006);
xor U20778 (N_20778,N_20138,N_20396);
xnor U20779 (N_20779,N_20245,N_20321);
nand U20780 (N_20780,N_20478,N_20365);
nand U20781 (N_20781,N_20139,N_20343);
nor U20782 (N_20782,N_20140,N_20078);
and U20783 (N_20783,N_20061,N_20340);
nand U20784 (N_20784,N_20065,N_20129);
or U20785 (N_20785,N_20479,N_20065);
nand U20786 (N_20786,N_20039,N_20227);
or U20787 (N_20787,N_20016,N_20025);
xor U20788 (N_20788,N_20261,N_20293);
or U20789 (N_20789,N_20366,N_20228);
nand U20790 (N_20790,N_20091,N_20376);
xor U20791 (N_20791,N_20232,N_20213);
nor U20792 (N_20792,N_20379,N_20010);
xor U20793 (N_20793,N_20105,N_20068);
nor U20794 (N_20794,N_20184,N_20385);
xnor U20795 (N_20795,N_20471,N_20357);
nor U20796 (N_20796,N_20294,N_20418);
nor U20797 (N_20797,N_20377,N_20125);
and U20798 (N_20798,N_20419,N_20098);
and U20799 (N_20799,N_20192,N_20034);
nor U20800 (N_20800,N_20084,N_20427);
xor U20801 (N_20801,N_20116,N_20287);
nand U20802 (N_20802,N_20160,N_20177);
or U20803 (N_20803,N_20240,N_20086);
and U20804 (N_20804,N_20341,N_20276);
or U20805 (N_20805,N_20317,N_20267);
and U20806 (N_20806,N_20310,N_20485);
or U20807 (N_20807,N_20109,N_20292);
or U20808 (N_20808,N_20172,N_20276);
nand U20809 (N_20809,N_20440,N_20231);
nand U20810 (N_20810,N_20079,N_20029);
xnor U20811 (N_20811,N_20026,N_20296);
nand U20812 (N_20812,N_20013,N_20254);
or U20813 (N_20813,N_20315,N_20295);
or U20814 (N_20814,N_20452,N_20022);
and U20815 (N_20815,N_20441,N_20157);
xnor U20816 (N_20816,N_20476,N_20472);
and U20817 (N_20817,N_20268,N_20379);
or U20818 (N_20818,N_20385,N_20357);
and U20819 (N_20819,N_20264,N_20247);
and U20820 (N_20820,N_20090,N_20320);
or U20821 (N_20821,N_20091,N_20401);
nor U20822 (N_20822,N_20015,N_20169);
or U20823 (N_20823,N_20185,N_20172);
xnor U20824 (N_20824,N_20281,N_20366);
nand U20825 (N_20825,N_20147,N_20106);
nor U20826 (N_20826,N_20277,N_20137);
nand U20827 (N_20827,N_20252,N_20161);
or U20828 (N_20828,N_20204,N_20287);
nand U20829 (N_20829,N_20411,N_20197);
nor U20830 (N_20830,N_20361,N_20458);
nor U20831 (N_20831,N_20059,N_20271);
xor U20832 (N_20832,N_20395,N_20089);
nor U20833 (N_20833,N_20136,N_20485);
nor U20834 (N_20834,N_20382,N_20236);
nor U20835 (N_20835,N_20265,N_20337);
nor U20836 (N_20836,N_20261,N_20031);
and U20837 (N_20837,N_20123,N_20493);
nor U20838 (N_20838,N_20272,N_20040);
nor U20839 (N_20839,N_20235,N_20128);
nand U20840 (N_20840,N_20047,N_20264);
and U20841 (N_20841,N_20411,N_20242);
nor U20842 (N_20842,N_20211,N_20399);
nand U20843 (N_20843,N_20340,N_20234);
nand U20844 (N_20844,N_20257,N_20029);
xnor U20845 (N_20845,N_20258,N_20315);
xor U20846 (N_20846,N_20030,N_20062);
nand U20847 (N_20847,N_20279,N_20162);
and U20848 (N_20848,N_20360,N_20363);
nand U20849 (N_20849,N_20060,N_20019);
nand U20850 (N_20850,N_20383,N_20163);
and U20851 (N_20851,N_20456,N_20063);
nor U20852 (N_20852,N_20443,N_20209);
and U20853 (N_20853,N_20331,N_20266);
nor U20854 (N_20854,N_20323,N_20230);
and U20855 (N_20855,N_20387,N_20267);
and U20856 (N_20856,N_20465,N_20067);
and U20857 (N_20857,N_20019,N_20414);
xnor U20858 (N_20858,N_20094,N_20316);
xnor U20859 (N_20859,N_20160,N_20313);
xor U20860 (N_20860,N_20419,N_20354);
nand U20861 (N_20861,N_20317,N_20233);
xnor U20862 (N_20862,N_20164,N_20229);
or U20863 (N_20863,N_20280,N_20364);
xnor U20864 (N_20864,N_20442,N_20465);
nor U20865 (N_20865,N_20323,N_20300);
nand U20866 (N_20866,N_20354,N_20010);
or U20867 (N_20867,N_20450,N_20459);
nand U20868 (N_20868,N_20127,N_20327);
or U20869 (N_20869,N_20381,N_20224);
and U20870 (N_20870,N_20441,N_20069);
nor U20871 (N_20871,N_20480,N_20494);
nor U20872 (N_20872,N_20087,N_20209);
and U20873 (N_20873,N_20198,N_20482);
and U20874 (N_20874,N_20022,N_20413);
xnor U20875 (N_20875,N_20238,N_20336);
and U20876 (N_20876,N_20028,N_20277);
or U20877 (N_20877,N_20230,N_20049);
nor U20878 (N_20878,N_20428,N_20407);
xor U20879 (N_20879,N_20183,N_20044);
or U20880 (N_20880,N_20330,N_20174);
and U20881 (N_20881,N_20379,N_20215);
xor U20882 (N_20882,N_20347,N_20145);
and U20883 (N_20883,N_20002,N_20069);
or U20884 (N_20884,N_20398,N_20203);
and U20885 (N_20885,N_20123,N_20294);
nor U20886 (N_20886,N_20455,N_20052);
nand U20887 (N_20887,N_20262,N_20254);
xnor U20888 (N_20888,N_20382,N_20287);
nor U20889 (N_20889,N_20166,N_20157);
xor U20890 (N_20890,N_20225,N_20253);
nor U20891 (N_20891,N_20159,N_20376);
nor U20892 (N_20892,N_20130,N_20312);
nor U20893 (N_20893,N_20187,N_20244);
or U20894 (N_20894,N_20216,N_20212);
or U20895 (N_20895,N_20085,N_20182);
nor U20896 (N_20896,N_20441,N_20027);
nand U20897 (N_20897,N_20372,N_20432);
or U20898 (N_20898,N_20334,N_20432);
nand U20899 (N_20899,N_20458,N_20100);
nand U20900 (N_20900,N_20231,N_20235);
or U20901 (N_20901,N_20471,N_20120);
and U20902 (N_20902,N_20339,N_20072);
xnor U20903 (N_20903,N_20255,N_20088);
nor U20904 (N_20904,N_20433,N_20082);
and U20905 (N_20905,N_20030,N_20184);
xor U20906 (N_20906,N_20163,N_20222);
xnor U20907 (N_20907,N_20353,N_20061);
nor U20908 (N_20908,N_20390,N_20250);
and U20909 (N_20909,N_20151,N_20086);
nand U20910 (N_20910,N_20202,N_20285);
nor U20911 (N_20911,N_20064,N_20112);
nor U20912 (N_20912,N_20341,N_20029);
nand U20913 (N_20913,N_20181,N_20118);
xnor U20914 (N_20914,N_20346,N_20400);
and U20915 (N_20915,N_20407,N_20337);
and U20916 (N_20916,N_20345,N_20010);
and U20917 (N_20917,N_20210,N_20422);
nor U20918 (N_20918,N_20414,N_20201);
nor U20919 (N_20919,N_20215,N_20002);
or U20920 (N_20920,N_20119,N_20254);
or U20921 (N_20921,N_20278,N_20220);
nand U20922 (N_20922,N_20004,N_20322);
xor U20923 (N_20923,N_20434,N_20028);
nor U20924 (N_20924,N_20007,N_20357);
and U20925 (N_20925,N_20412,N_20459);
nand U20926 (N_20926,N_20152,N_20122);
xor U20927 (N_20927,N_20224,N_20092);
nor U20928 (N_20928,N_20314,N_20293);
and U20929 (N_20929,N_20195,N_20490);
or U20930 (N_20930,N_20001,N_20245);
and U20931 (N_20931,N_20131,N_20008);
or U20932 (N_20932,N_20237,N_20438);
or U20933 (N_20933,N_20017,N_20460);
and U20934 (N_20934,N_20252,N_20002);
nand U20935 (N_20935,N_20361,N_20146);
or U20936 (N_20936,N_20242,N_20346);
or U20937 (N_20937,N_20311,N_20374);
xnor U20938 (N_20938,N_20167,N_20002);
nor U20939 (N_20939,N_20189,N_20068);
xnor U20940 (N_20940,N_20040,N_20226);
nand U20941 (N_20941,N_20388,N_20346);
and U20942 (N_20942,N_20137,N_20211);
and U20943 (N_20943,N_20084,N_20226);
or U20944 (N_20944,N_20204,N_20457);
and U20945 (N_20945,N_20281,N_20393);
or U20946 (N_20946,N_20052,N_20344);
and U20947 (N_20947,N_20214,N_20307);
and U20948 (N_20948,N_20321,N_20265);
nor U20949 (N_20949,N_20277,N_20407);
and U20950 (N_20950,N_20327,N_20354);
nor U20951 (N_20951,N_20308,N_20384);
nand U20952 (N_20952,N_20017,N_20212);
xor U20953 (N_20953,N_20037,N_20175);
nor U20954 (N_20954,N_20289,N_20457);
xnor U20955 (N_20955,N_20333,N_20093);
xor U20956 (N_20956,N_20415,N_20148);
and U20957 (N_20957,N_20324,N_20106);
nor U20958 (N_20958,N_20432,N_20395);
and U20959 (N_20959,N_20399,N_20063);
or U20960 (N_20960,N_20106,N_20395);
or U20961 (N_20961,N_20265,N_20240);
and U20962 (N_20962,N_20232,N_20316);
nor U20963 (N_20963,N_20274,N_20247);
nand U20964 (N_20964,N_20213,N_20401);
nor U20965 (N_20965,N_20296,N_20073);
nor U20966 (N_20966,N_20157,N_20125);
nor U20967 (N_20967,N_20344,N_20214);
nor U20968 (N_20968,N_20391,N_20056);
nor U20969 (N_20969,N_20350,N_20142);
or U20970 (N_20970,N_20338,N_20409);
and U20971 (N_20971,N_20221,N_20323);
and U20972 (N_20972,N_20076,N_20015);
or U20973 (N_20973,N_20251,N_20087);
or U20974 (N_20974,N_20457,N_20132);
xor U20975 (N_20975,N_20449,N_20215);
and U20976 (N_20976,N_20359,N_20143);
nand U20977 (N_20977,N_20396,N_20190);
or U20978 (N_20978,N_20242,N_20078);
nor U20979 (N_20979,N_20232,N_20445);
nor U20980 (N_20980,N_20420,N_20144);
xnor U20981 (N_20981,N_20481,N_20459);
or U20982 (N_20982,N_20025,N_20395);
nand U20983 (N_20983,N_20158,N_20429);
xor U20984 (N_20984,N_20251,N_20434);
nor U20985 (N_20985,N_20395,N_20348);
xnor U20986 (N_20986,N_20202,N_20020);
and U20987 (N_20987,N_20172,N_20261);
or U20988 (N_20988,N_20357,N_20396);
xnor U20989 (N_20989,N_20364,N_20358);
nand U20990 (N_20990,N_20421,N_20112);
nand U20991 (N_20991,N_20078,N_20302);
nor U20992 (N_20992,N_20138,N_20393);
nand U20993 (N_20993,N_20354,N_20323);
nor U20994 (N_20994,N_20467,N_20152);
and U20995 (N_20995,N_20415,N_20188);
or U20996 (N_20996,N_20375,N_20341);
nor U20997 (N_20997,N_20317,N_20147);
nand U20998 (N_20998,N_20388,N_20183);
and U20999 (N_20999,N_20261,N_20327);
nor U21000 (N_21000,N_20783,N_20866);
and U21001 (N_21001,N_20694,N_20935);
or U21002 (N_21002,N_20707,N_20683);
xnor U21003 (N_21003,N_20727,N_20562);
nand U21004 (N_21004,N_20863,N_20893);
or U21005 (N_21005,N_20854,N_20734);
xor U21006 (N_21006,N_20872,N_20641);
xor U21007 (N_21007,N_20503,N_20899);
or U21008 (N_21008,N_20965,N_20617);
nand U21009 (N_21009,N_20542,N_20767);
xnor U21010 (N_21010,N_20826,N_20917);
nor U21011 (N_21011,N_20753,N_20650);
xnor U21012 (N_21012,N_20981,N_20631);
and U21013 (N_21013,N_20787,N_20565);
xor U21014 (N_21014,N_20797,N_20953);
or U21015 (N_21015,N_20582,N_20968);
xor U21016 (N_21016,N_20585,N_20554);
nand U21017 (N_21017,N_20771,N_20776);
nor U21018 (N_21018,N_20894,N_20875);
xnor U21019 (N_21019,N_20836,N_20931);
nor U21020 (N_21020,N_20583,N_20505);
nand U21021 (N_21021,N_20906,N_20999);
and U21022 (N_21022,N_20918,N_20985);
or U21023 (N_21023,N_20561,N_20969);
or U21024 (N_21024,N_20880,N_20937);
nor U21025 (N_21025,N_20611,N_20785);
and U21026 (N_21026,N_20544,N_20890);
or U21027 (N_21027,N_20603,N_20667);
xor U21028 (N_21028,N_20512,N_20747);
nand U21029 (N_21029,N_20764,N_20812);
nor U21030 (N_21030,N_20710,N_20573);
xnor U21031 (N_21031,N_20830,N_20598);
nand U21032 (N_21032,N_20672,N_20994);
xnor U21033 (N_21033,N_20853,N_20577);
nand U21034 (N_21034,N_20892,N_20639);
xor U21035 (N_21035,N_20809,N_20526);
xor U21036 (N_21036,N_20599,N_20926);
nand U21037 (N_21037,N_20795,N_20742);
nand U21038 (N_21038,N_20916,N_20986);
or U21039 (N_21039,N_20665,N_20769);
xnor U21040 (N_21040,N_20557,N_20861);
or U21041 (N_21041,N_20592,N_20622);
nor U21042 (N_21042,N_20704,N_20886);
xor U21043 (N_21043,N_20946,N_20515);
and U21044 (N_21044,N_20539,N_20612);
and U21045 (N_21045,N_20756,N_20609);
or U21046 (N_21046,N_20685,N_20740);
or U21047 (N_21047,N_20647,N_20675);
xnor U21048 (N_21048,N_20658,N_20676);
or U21049 (N_21049,N_20898,N_20807);
or U21050 (N_21050,N_20668,N_20649);
xor U21051 (N_21051,N_20950,N_20849);
nand U21052 (N_21052,N_20614,N_20746);
xnor U21053 (N_21053,N_20816,N_20957);
nand U21054 (N_21054,N_20663,N_20600);
nor U21055 (N_21055,N_20885,N_20750);
nor U21056 (N_21056,N_20975,N_20788);
nor U21057 (N_21057,N_20961,N_20778);
nor U21058 (N_21058,N_20835,N_20703);
or U21059 (N_21059,N_20630,N_20628);
nor U21060 (N_21060,N_20948,N_20934);
xnor U21061 (N_21061,N_20971,N_20654);
or U21062 (N_21062,N_20633,N_20869);
xnor U21063 (N_21063,N_20643,N_20989);
nor U21064 (N_21064,N_20721,N_20709);
xnor U21065 (N_21065,N_20855,N_20621);
xnor U21066 (N_21066,N_20824,N_20902);
and U21067 (N_21067,N_20843,N_20519);
or U21068 (N_21068,N_20550,N_20524);
and U21069 (N_21069,N_20729,N_20716);
xnor U21070 (N_21070,N_20578,N_20731);
or U21071 (N_21071,N_20605,N_20556);
or U21072 (N_21072,N_20547,N_20574);
xnor U21073 (N_21073,N_20817,N_20960);
or U21074 (N_21074,N_20543,N_20674);
or U21075 (N_21075,N_20932,N_20990);
nand U21076 (N_21076,N_20827,N_20511);
or U21077 (N_21077,N_20768,N_20838);
nor U21078 (N_21078,N_20638,N_20848);
nand U21079 (N_21079,N_20933,N_20798);
and U21080 (N_21080,N_20586,N_20927);
xor U21081 (N_21081,N_20558,N_20888);
xor U21082 (N_21082,N_20770,N_20864);
xor U21083 (N_21083,N_20992,N_20741);
nor U21084 (N_21084,N_20858,N_20745);
nand U21085 (N_21085,N_20692,N_20518);
xor U21086 (N_21086,N_20867,N_20613);
nor U21087 (N_21087,N_20711,N_20684);
xnor U21088 (N_21088,N_20878,N_20514);
and U21089 (N_21089,N_20792,N_20737);
nand U21090 (N_21090,N_20588,N_20587);
or U21091 (N_21091,N_20720,N_20998);
and U21092 (N_21092,N_20686,N_20806);
nor U21093 (N_21093,N_20620,N_20677);
and U21094 (N_21094,N_20559,N_20528);
or U21095 (N_21095,N_20952,N_20755);
nor U21096 (N_21096,N_20629,N_20713);
nor U21097 (N_21097,N_20996,N_20831);
nand U21098 (N_21098,N_20634,N_20506);
or U21099 (N_21099,N_20736,N_20991);
xnor U21100 (N_21100,N_20666,N_20604);
xor U21101 (N_21101,N_20819,N_20532);
nor U21102 (N_21102,N_20718,N_20618);
nand U21103 (N_21103,N_20627,N_20794);
or U21104 (N_21104,N_20936,N_20921);
nand U21105 (N_21105,N_20680,N_20735);
and U21106 (N_21106,N_20758,N_20607);
or U21107 (N_21107,N_20963,N_20567);
xor U21108 (N_21108,N_20661,N_20615);
nor U21109 (N_21109,N_20874,N_20842);
nor U21110 (N_21110,N_20801,N_20723);
xnor U21111 (N_21111,N_20944,N_20743);
xor U21112 (N_21112,N_20608,N_20689);
nand U21113 (N_21113,N_20681,N_20571);
and U21114 (N_21114,N_20911,N_20651);
xor U21115 (N_21115,N_20988,N_20974);
xor U21116 (N_21116,N_20870,N_20943);
or U21117 (N_21117,N_20715,N_20509);
nand U21118 (N_21118,N_20763,N_20871);
xnor U21119 (N_21119,N_20859,N_20576);
and U21120 (N_21120,N_20945,N_20891);
xnor U21121 (N_21121,N_20796,N_20669);
nand U21122 (N_21122,N_20821,N_20865);
nor U21123 (N_21123,N_20976,N_20572);
and U21124 (N_21124,N_20897,N_20517);
or U21125 (N_21125,N_20939,N_20876);
and U21126 (N_21126,N_20593,N_20664);
xor U21127 (N_21127,N_20800,N_20982);
or U21128 (N_21128,N_20706,N_20850);
xnor U21129 (N_21129,N_20722,N_20920);
and U21130 (N_21130,N_20712,N_20564);
nor U21131 (N_21131,N_20860,N_20852);
and U21132 (N_21132,N_20697,N_20760);
or U21133 (N_21133,N_20749,N_20534);
nand U21134 (N_21134,N_20823,N_20695);
and U21135 (N_21135,N_20648,N_20657);
xnor U21136 (N_21136,N_20903,N_20616);
nor U21137 (N_21137,N_20958,N_20780);
or U21138 (N_21138,N_20705,N_20752);
or U21139 (N_21139,N_20546,N_20868);
nor U21140 (N_21140,N_20732,N_20540);
or U21141 (N_21141,N_20688,N_20660);
and U21142 (N_21142,N_20580,N_20766);
xor U21143 (N_21143,N_20761,N_20653);
nor U21144 (N_21144,N_20837,N_20527);
nand U21145 (N_21145,N_20635,N_20825);
nand U21146 (N_21146,N_20726,N_20698);
xor U21147 (N_21147,N_20938,N_20765);
xor U21148 (N_21148,N_20645,N_20815);
nand U21149 (N_21149,N_20700,N_20533);
nor U21150 (N_21150,N_20808,N_20995);
or U21151 (N_21151,N_20791,N_20956);
and U21152 (N_21152,N_20719,N_20507);
or U21153 (N_21153,N_20775,N_20520);
xor U21154 (N_21154,N_20530,N_20966);
nor U21155 (N_21155,N_20671,N_20714);
and U21156 (N_21156,N_20959,N_20951);
or U21157 (N_21157,N_20513,N_20909);
xor U21158 (N_21158,N_20922,N_20904);
nand U21159 (N_21159,N_20896,N_20717);
nor U21160 (N_21160,N_20744,N_20846);
nand U21161 (N_21161,N_20662,N_20883);
xor U21162 (N_21162,N_20644,N_20606);
nor U21163 (N_21163,N_20560,N_20820);
nor U21164 (N_21164,N_20673,N_20579);
nand U21165 (N_21165,N_20594,N_20678);
and U21166 (N_21166,N_20925,N_20905);
or U21167 (N_21167,N_20708,N_20522);
nor U21168 (N_21168,N_20529,N_20738);
xor U21169 (N_21169,N_20774,N_20777);
nand U21170 (N_21170,N_20730,N_20551);
nor U21171 (N_21171,N_20851,N_20637);
or U21172 (N_21172,N_20923,N_20987);
and U21173 (N_21173,N_20632,N_20782);
or U21174 (N_21174,N_20977,N_20814);
nor U21175 (N_21175,N_20829,N_20954);
xor U21176 (N_21176,N_20679,N_20873);
nor U21177 (N_21177,N_20523,N_20907);
nor U21178 (N_21178,N_20822,N_20724);
nor U21179 (N_21179,N_20504,N_20701);
nand U21180 (N_21180,N_20832,N_20748);
nand U21181 (N_21181,N_20979,N_20919);
nand U21182 (N_21182,N_20924,N_20793);
and U21183 (N_21183,N_20623,N_20563);
nand U21184 (N_21184,N_20828,N_20862);
xnor U21185 (N_21185,N_20589,N_20844);
or U21186 (N_21186,N_20656,N_20652);
xor U21187 (N_21187,N_20789,N_20941);
and U21188 (N_21188,N_20913,N_20912);
xor U21189 (N_21189,N_20610,N_20591);
and U21190 (N_21190,N_20659,N_20940);
or U21191 (N_21191,N_20553,N_20900);
or U21192 (N_21192,N_20799,N_20502);
and U21193 (N_21193,N_20877,N_20696);
nor U21194 (N_21194,N_20786,N_20699);
and U21195 (N_21195,N_20915,N_20790);
xor U21196 (N_21196,N_20624,N_20847);
nor U21197 (N_21197,N_20839,N_20549);
nand U21198 (N_21198,N_20702,N_20619);
nand U21199 (N_21199,N_20537,N_20569);
xor U21200 (N_21200,N_20626,N_20640);
nand U21201 (N_21201,N_20772,N_20857);
nor U21202 (N_21202,N_20687,N_20818);
or U21203 (N_21203,N_20584,N_20840);
nand U21204 (N_21204,N_20601,N_20779);
or U21205 (N_21205,N_20942,N_20541);
or U21206 (N_21206,N_20682,N_20501);
xnor U21207 (N_21207,N_20983,N_20725);
nand U21208 (N_21208,N_20972,N_20762);
nor U21209 (N_21209,N_20552,N_20895);
xnor U21210 (N_21210,N_20575,N_20910);
nand U21211 (N_21211,N_20970,N_20930);
xor U21212 (N_21212,N_20646,N_20636);
nor U21213 (N_21213,N_20879,N_20984);
nand U21214 (N_21214,N_20548,N_20805);
nand U21215 (N_21215,N_20536,N_20690);
nand U21216 (N_21216,N_20884,N_20516);
or U21217 (N_21217,N_20545,N_20803);
or U21218 (N_21218,N_20882,N_20811);
and U21219 (N_21219,N_20568,N_20595);
and U21220 (N_21220,N_20508,N_20914);
nor U21221 (N_21221,N_20773,N_20590);
or U21222 (N_21222,N_20881,N_20784);
nor U21223 (N_21223,N_20655,N_20833);
nor U21224 (N_21224,N_20670,N_20993);
and U21225 (N_21225,N_20997,N_20510);
nor U21226 (N_21226,N_20555,N_20521);
or U21227 (N_21227,N_20693,N_20691);
nand U21228 (N_21228,N_20802,N_20602);
nor U21229 (N_21229,N_20804,N_20973);
nand U21230 (N_21230,N_20813,N_20566);
nand U21231 (N_21231,N_20889,N_20733);
nand U21232 (N_21232,N_20845,N_20908);
nor U21233 (N_21233,N_20570,N_20967);
nand U21234 (N_21234,N_20581,N_20759);
and U21235 (N_21235,N_20538,N_20901);
or U21236 (N_21236,N_20596,N_20955);
nand U21237 (N_21237,N_20856,N_20928);
or U21238 (N_21238,N_20531,N_20841);
nand U21239 (N_21239,N_20625,N_20947);
and U21240 (N_21240,N_20781,N_20739);
or U21241 (N_21241,N_20535,N_20929);
nand U21242 (N_21242,N_20597,N_20949);
nor U21243 (N_21243,N_20980,N_20728);
xnor U21244 (N_21244,N_20962,N_20810);
nor U21245 (N_21245,N_20887,N_20642);
or U21246 (N_21246,N_20757,N_20500);
and U21247 (N_21247,N_20754,N_20978);
xor U21248 (N_21248,N_20834,N_20964);
nand U21249 (N_21249,N_20751,N_20525);
nor U21250 (N_21250,N_20628,N_20551);
or U21251 (N_21251,N_20922,N_20923);
xnor U21252 (N_21252,N_20905,N_20612);
or U21253 (N_21253,N_20915,N_20745);
nand U21254 (N_21254,N_20636,N_20609);
nor U21255 (N_21255,N_20965,N_20924);
and U21256 (N_21256,N_20692,N_20577);
or U21257 (N_21257,N_20884,N_20749);
nand U21258 (N_21258,N_20792,N_20875);
nand U21259 (N_21259,N_20584,N_20623);
xor U21260 (N_21260,N_20848,N_20551);
or U21261 (N_21261,N_20851,N_20978);
xor U21262 (N_21262,N_20841,N_20778);
or U21263 (N_21263,N_20814,N_20809);
nand U21264 (N_21264,N_20737,N_20526);
or U21265 (N_21265,N_20673,N_20963);
nand U21266 (N_21266,N_20957,N_20970);
and U21267 (N_21267,N_20931,N_20667);
xor U21268 (N_21268,N_20930,N_20816);
xnor U21269 (N_21269,N_20895,N_20862);
nand U21270 (N_21270,N_20918,N_20681);
nand U21271 (N_21271,N_20945,N_20883);
or U21272 (N_21272,N_20946,N_20676);
nand U21273 (N_21273,N_20833,N_20606);
nor U21274 (N_21274,N_20900,N_20712);
and U21275 (N_21275,N_20742,N_20561);
or U21276 (N_21276,N_20638,N_20874);
nand U21277 (N_21277,N_20501,N_20878);
and U21278 (N_21278,N_20532,N_20713);
nor U21279 (N_21279,N_20928,N_20689);
nor U21280 (N_21280,N_20939,N_20864);
and U21281 (N_21281,N_20766,N_20557);
or U21282 (N_21282,N_20686,N_20556);
nand U21283 (N_21283,N_20877,N_20513);
nor U21284 (N_21284,N_20664,N_20967);
xor U21285 (N_21285,N_20853,N_20854);
xor U21286 (N_21286,N_20654,N_20536);
and U21287 (N_21287,N_20857,N_20875);
and U21288 (N_21288,N_20974,N_20684);
xor U21289 (N_21289,N_20546,N_20958);
nand U21290 (N_21290,N_20870,N_20957);
nor U21291 (N_21291,N_20646,N_20519);
xnor U21292 (N_21292,N_20806,N_20525);
nand U21293 (N_21293,N_20882,N_20960);
nand U21294 (N_21294,N_20620,N_20659);
and U21295 (N_21295,N_20885,N_20987);
xor U21296 (N_21296,N_20943,N_20836);
nand U21297 (N_21297,N_20721,N_20859);
xnor U21298 (N_21298,N_20838,N_20770);
and U21299 (N_21299,N_20672,N_20872);
xnor U21300 (N_21300,N_20678,N_20610);
nor U21301 (N_21301,N_20673,N_20853);
and U21302 (N_21302,N_20905,N_20916);
or U21303 (N_21303,N_20675,N_20504);
xor U21304 (N_21304,N_20918,N_20995);
nand U21305 (N_21305,N_20934,N_20821);
and U21306 (N_21306,N_20903,N_20799);
or U21307 (N_21307,N_20666,N_20557);
nand U21308 (N_21308,N_20933,N_20940);
or U21309 (N_21309,N_20987,N_20837);
and U21310 (N_21310,N_20620,N_20711);
nor U21311 (N_21311,N_20989,N_20968);
and U21312 (N_21312,N_20636,N_20712);
xnor U21313 (N_21313,N_20927,N_20886);
nand U21314 (N_21314,N_20749,N_20909);
xnor U21315 (N_21315,N_20846,N_20743);
nor U21316 (N_21316,N_20715,N_20668);
nor U21317 (N_21317,N_20553,N_20795);
nand U21318 (N_21318,N_20901,N_20917);
nand U21319 (N_21319,N_20702,N_20560);
and U21320 (N_21320,N_20613,N_20562);
nand U21321 (N_21321,N_20752,N_20882);
xor U21322 (N_21322,N_20886,N_20767);
xnor U21323 (N_21323,N_20937,N_20668);
or U21324 (N_21324,N_20872,N_20808);
and U21325 (N_21325,N_20996,N_20722);
and U21326 (N_21326,N_20868,N_20750);
nand U21327 (N_21327,N_20981,N_20968);
and U21328 (N_21328,N_20560,N_20735);
and U21329 (N_21329,N_20504,N_20848);
xor U21330 (N_21330,N_20540,N_20871);
xor U21331 (N_21331,N_20775,N_20646);
xor U21332 (N_21332,N_20963,N_20783);
or U21333 (N_21333,N_20532,N_20607);
nand U21334 (N_21334,N_20572,N_20540);
or U21335 (N_21335,N_20604,N_20945);
and U21336 (N_21336,N_20729,N_20932);
xor U21337 (N_21337,N_20655,N_20964);
and U21338 (N_21338,N_20836,N_20819);
and U21339 (N_21339,N_20964,N_20863);
and U21340 (N_21340,N_20887,N_20942);
nor U21341 (N_21341,N_20764,N_20721);
xnor U21342 (N_21342,N_20769,N_20813);
nor U21343 (N_21343,N_20996,N_20948);
xor U21344 (N_21344,N_20914,N_20680);
and U21345 (N_21345,N_20552,N_20979);
nand U21346 (N_21346,N_20859,N_20564);
and U21347 (N_21347,N_20760,N_20938);
nand U21348 (N_21348,N_20656,N_20586);
or U21349 (N_21349,N_20967,N_20893);
nand U21350 (N_21350,N_20527,N_20992);
nand U21351 (N_21351,N_20715,N_20535);
nand U21352 (N_21352,N_20921,N_20883);
nand U21353 (N_21353,N_20611,N_20679);
xnor U21354 (N_21354,N_20821,N_20509);
and U21355 (N_21355,N_20962,N_20639);
xnor U21356 (N_21356,N_20735,N_20966);
nor U21357 (N_21357,N_20520,N_20720);
nand U21358 (N_21358,N_20579,N_20819);
and U21359 (N_21359,N_20765,N_20729);
nor U21360 (N_21360,N_20859,N_20756);
xor U21361 (N_21361,N_20583,N_20596);
and U21362 (N_21362,N_20864,N_20851);
nand U21363 (N_21363,N_20581,N_20664);
or U21364 (N_21364,N_20865,N_20739);
or U21365 (N_21365,N_20629,N_20741);
xnor U21366 (N_21366,N_20851,N_20867);
and U21367 (N_21367,N_20703,N_20614);
or U21368 (N_21368,N_20844,N_20732);
nand U21369 (N_21369,N_20803,N_20753);
nor U21370 (N_21370,N_20633,N_20903);
and U21371 (N_21371,N_20699,N_20666);
or U21372 (N_21372,N_20786,N_20611);
nor U21373 (N_21373,N_20881,N_20846);
or U21374 (N_21374,N_20935,N_20846);
xor U21375 (N_21375,N_20775,N_20619);
xor U21376 (N_21376,N_20799,N_20781);
xor U21377 (N_21377,N_20958,N_20837);
and U21378 (N_21378,N_20931,N_20898);
nand U21379 (N_21379,N_20970,N_20650);
nor U21380 (N_21380,N_20626,N_20504);
and U21381 (N_21381,N_20560,N_20917);
nand U21382 (N_21382,N_20959,N_20613);
xnor U21383 (N_21383,N_20814,N_20584);
nor U21384 (N_21384,N_20876,N_20975);
nor U21385 (N_21385,N_20715,N_20664);
nand U21386 (N_21386,N_20626,N_20576);
or U21387 (N_21387,N_20751,N_20651);
nor U21388 (N_21388,N_20950,N_20915);
nor U21389 (N_21389,N_20909,N_20792);
nand U21390 (N_21390,N_20929,N_20845);
nor U21391 (N_21391,N_20572,N_20608);
nor U21392 (N_21392,N_20815,N_20914);
and U21393 (N_21393,N_20655,N_20887);
nand U21394 (N_21394,N_20593,N_20665);
nand U21395 (N_21395,N_20695,N_20528);
nand U21396 (N_21396,N_20541,N_20976);
and U21397 (N_21397,N_20709,N_20649);
nand U21398 (N_21398,N_20987,N_20776);
nor U21399 (N_21399,N_20989,N_20613);
xnor U21400 (N_21400,N_20562,N_20808);
or U21401 (N_21401,N_20766,N_20728);
or U21402 (N_21402,N_20598,N_20963);
nor U21403 (N_21403,N_20805,N_20712);
or U21404 (N_21404,N_20980,N_20889);
xor U21405 (N_21405,N_20759,N_20647);
and U21406 (N_21406,N_20888,N_20857);
nor U21407 (N_21407,N_20618,N_20908);
nand U21408 (N_21408,N_20705,N_20952);
or U21409 (N_21409,N_20723,N_20774);
nor U21410 (N_21410,N_20556,N_20912);
or U21411 (N_21411,N_20644,N_20812);
or U21412 (N_21412,N_20925,N_20961);
and U21413 (N_21413,N_20986,N_20742);
xnor U21414 (N_21414,N_20883,N_20869);
or U21415 (N_21415,N_20893,N_20998);
nor U21416 (N_21416,N_20562,N_20523);
nand U21417 (N_21417,N_20894,N_20735);
or U21418 (N_21418,N_20666,N_20705);
or U21419 (N_21419,N_20843,N_20518);
nor U21420 (N_21420,N_20783,N_20637);
or U21421 (N_21421,N_20817,N_20581);
and U21422 (N_21422,N_20928,N_20579);
nor U21423 (N_21423,N_20698,N_20552);
xor U21424 (N_21424,N_20598,N_20927);
nand U21425 (N_21425,N_20864,N_20807);
and U21426 (N_21426,N_20516,N_20737);
nor U21427 (N_21427,N_20619,N_20960);
nor U21428 (N_21428,N_20791,N_20670);
nor U21429 (N_21429,N_20653,N_20855);
or U21430 (N_21430,N_20892,N_20878);
and U21431 (N_21431,N_20613,N_20726);
nor U21432 (N_21432,N_20862,N_20674);
xor U21433 (N_21433,N_20964,N_20841);
nor U21434 (N_21434,N_20643,N_20959);
xor U21435 (N_21435,N_20926,N_20760);
nand U21436 (N_21436,N_20842,N_20509);
xor U21437 (N_21437,N_20645,N_20710);
and U21438 (N_21438,N_20620,N_20993);
and U21439 (N_21439,N_20735,N_20564);
and U21440 (N_21440,N_20584,N_20632);
nor U21441 (N_21441,N_20928,N_20576);
nor U21442 (N_21442,N_20960,N_20703);
and U21443 (N_21443,N_20546,N_20826);
nor U21444 (N_21444,N_20814,N_20756);
and U21445 (N_21445,N_20741,N_20954);
nand U21446 (N_21446,N_20990,N_20998);
nor U21447 (N_21447,N_20945,N_20575);
nand U21448 (N_21448,N_20544,N_20760);
nor U21449 (N_21449,N_20721,N_20733);
and U21450 (N_21450,N_20839,N_20837);
xnor U21451 (N_21451,N_20916,N_20751);
nand U21452 (N_21452,N_20745,N_20668);
nand U21453 (N_21453,N_20677,N_20671);
and U21454 (N_21454,N_20656,N_20549);
xnor U21455 (N_21455,N_20916,N_20712);
and U21456 (N_21456,N_20731,N_20505);
xnor U21457 (N_21457,N_20698,N_20607);
and U21458 (N_21458,N_20918,N_20714);
and U21459 (N_21459,N_20726,N_20930);
nor U21460 (N_21460,N_20653,N_20582);
xnor U21461 (N_21461,N_20985,N_20949);
nand U21462 (N_21462,N_20948,N_20541);
or U21463 (N_21463,N_20783,N_20640);
or U21464 (N_21464,N_20729,N_20820);
and U21465 (N_21465,N_20640,N_20674);
or U21466 (N_21466,N_20510,N_20632);
and U21467 (N_21467,N_20729,N_20870);
and U21468 (N_21468,N_20529,N_20568);
nand U21469 (N_21469,N_20988,N_20659);
nand U21470 (N_21470,N_20902,N_20961);
or U21471 (N_21471,N_20712,N_20953);
nor U21472 (N_21472,N_20849,N_20964);
or U21473 (N_21473,N_20831,N_20544);
nand U21474 (N_21474,N_20892,N_20605);
or U21475 (N_21475,N_20625,N_20527);
xnor U21476 (N_21476,N_20974,N_20556);
xnor U21477 (N_21477,N_20637,N_20770);
xor U21478 (N_21478,N_20616,N_20837);
or U21479 (N_21479,N_20649,N_20730);
nand U21480 (N_21480,N_20534,N_20836);
nand U21481 (N_21481,N_20561,N_20569);
nand U21482 (N_21482,N_20665,N_20639);
or U21483 (N_21483,N_20555,N_20854);
xor U21484 (N_21484,N_20559,N_20677);
nor U21485 (N_21485,N_20683,N_20564);
and U21486 (N_21486,N_20592,N_20652);
xnor U21487 (N_21487,N_20502,N_20797);
and U21488 (N_21488,N_20859,N_20916);
or U21489 (N_21489,N_20858,N_20971);
or U21490 (N_21490,N_20731,N_20532);
nand U21491 (N_21491,N_20563,N_20718);
nor U21492 (N_21492,N_20848,N_20734);
xnor U21493 (N_21493,N_20932,N_20903);
xnor U21494 (N_21494,N_20833,N_20942);
and U21495 (N_21495,N_20702,N_20943);
xor U21496 (N_21496,N_20821,N_20959);
xor U21497 (N_21497,N_20945,N_20802);
nand U21498 (N_21498,N_20721,N_20857);
nor U21499 (N_21499,N_20920,N_20650);
xnor U21500 (N_21500,N_21335,N_21084);
xnor U21501 (N_21501,N_21019,N_21179);
nor U21502 (N_21502,N_21227,N_21059);
nor U21503 (N_21503,N_21085,N_21418);
xnor U21504 (N_21504,N_21425,N_21138);
xnor U21505 (N_21505,N_21254,N_21024);
nor U21506 (N_21506,N_21011,N_21265);
nand U21507 (N_21507,N_21332,N_21397);
xnor U21508 (N_21508,N_21268,N_21412);
nand U21509 (N_21509,N_21384,N_21442);
nand U21510 (N_21510,N_21487,N_21427);
or U21511 (N_21511,N_21454,N_21220);
or U21512 (N_21512,N_21329,N_21074);
nand U21513 (N_21513,N_21090,N_21020);
or U21514 (N_21514,N_21103,N_21344);
nor U21515 (N_21515,N_21197,N_21486);
and U21516 (N_21516,N_21353,N_21471);
xnor U21517 (N_21517,N_21290,N_21099);
xnor U21518 (N_21518,N_21441,N_21255);
xor U21519 (N_21519,N_21192,N_21079);
and U21520 (N_21520,N_21194,N_21027);
or U21521 (N_21521,N_21330,N_21060);
nand U21522 (N_21522,N_21392,N_21328);
or U21523 (N_21523,N_21434,N_21191);
xor U21524 (N_21524,N_21070,N_21023);
and U21525 (N_21525,N_21346,N_21495);
or U21526 (N_21526,N_21012,N_21081);
and U21527 (N_21527,N_21480,N_21307);
nor U21528 (N_21528,N_21008,N_21014);
nor U21529 (N_21529,N_21243,N_21363);
nand U21530 (N_21530,N_21201,N_21280);
nand U21531 (N_21531,N_21342,N_21388);
nand U21532 (N_21532,N_21244,N_21127);
xor U21533 (N_21533,N_21285,N_21190);
xor U21534 (N_21534,N_21176,N_21082);
nor U21535 (N_21535,N_21301,N_21206);
and U21536 (N_21536,N_21018,N_21222);
or U21537 (N_21537,N_21132,N_21025);
xor U21538 (N_21538,N_21391,N_21241);
nor U21539 (N_21539,N_21338,N_21393);
xor U21540 (N_21540,N_21459,N_21266);
xnor U21541 (N_21541,N_21137,N_21310);
nand U21542 (N_21542,N_21144,N_21210);
xor U21543 (N_21543,N_21112,N_21433);
and U21544 (N_21544,N_21386,N_21360);
or U21545 (N_21545,N_21325,N_21369);
xnor U21546 (N_21546,N_21409,N_21350);
nor U21547 (N_21547,N_21272,N_21147);
or U21548 (N_21548,N_21064,N_21443);
nand U21549 (N_21549,N_21479,N_21234);
and U21550 (N_21550,N_21087,N_21106);
xnor U21551 (N_21551,N_21080,N_21041);
and U21552 (N_21552,N_21093,N_21499);
or U21553 (N_21553,N_21037,N_21130);
and U21554 (N_21554,N_21049,N_21073);
or U21555 (N_21555,N_21256,N_21490);
or U21556 (N_21556,N_21086,N_21058);
and U21557 (N_21557,N_21390,N_21348);
xnor U21558 (N_21558,N_21212,N_21071);
or U21559 (N_21559,N_21383,N_21422);
or U21560 (N_21560,N_21199,N_21380);
nor U21561 (N_21561,N_21170,N_21450);
xnor U21562 (N_21562,N_21236,N_21213);
or U21563 (N_21563,N_21108,N_21322);
xnor U21564 (N_21564,N_21373,N_21336);
nor U21565 (N_21565,N_21264,N_21215);
or U21566 (N_21566,N_21477,N_21410);
and U21567 (N_21567,N_21283,N_21052);
or U21568 (N_21568,N_21200,N_21318);
nor U21569 (N_21569,N_21096,N_21028);
and U21570 (N_21570,N_21345,N_21046);
and U21571 (N_21571,N_21035,N_21382);
nand U21572 (N_21572,N_21149,N_21146);
and U21573 (N_21573,N_21022,N_21276);
nor U21574 (N_21574,N_21033,N_21327);
and U21575 (N_21575,N_21333,N_21180);
or U21576 (N_21576,N_21467,N_21349);
or U21577 (N_21577,N_21361,N_21447);
nand U21578 (N_21578,N_21293,N_21164);
or U21579 (N_21579,N_21061,N_21140);
and U21580 (N_21580,N_21182,N_21155);
and U21581 (N_21581,N_21337,N_21026);
or U21582 (N_21582,N_21262,N_21048);
xnor U21583 (N_21583,N_21102,N_21436);
xnor U21584 (N_21584,N_21284,N_21303);
or U21585 (N_21585,N_21143,N_21439);
nor U21586 (N_21586,N_21015,N_21152);
and U21587 (N_21587,N_21016,N_21317);
nor U21588 (N_21588,N_21472,N_21407);
nand U21589 (N_21589,N_21187,N_21211);
nand U21590 (N_21590,N_21116,N_21121);
and U21591 (N_21591,N_21316,N_21141);
and U21592 (N_21592,N_21413,N_21160);
nand U21593 (N_21593,N_21150,N_21078);
nand U21594 (N_21594,N_21068,N_21324);
nor U21595 (N_21595,N_21168,N_21151);
or U21596 (N_21596,N_21072,N_21420);
nand U21597 (N_21597,N_21107,N_21063);
nand U21598 (N_21598,N_21057,N_21435);
nand U21599 (N_21599,N_21295,N_21431);
or U21600 (N_21600,N_21229,N_21000);
nor U21601 (N_21601,N_21381,N_21083);
xnor U21602 (N_21602,N_21288,N_21437);
xor U21603 (N_21603,N_21257,N_21379);
nor U21604 (N_21604,N_21476,N_21173);
xnor U21605 (N_21605,N_21470,N_21294);
nand U21606 (N_21606,N_21251,N_21453);
nand U21607 (N_21607,N_21319,N_21448);
nor U21608 (N_21608,N_21242,N_21183);
and U21609 (N_21609,N_21461,N_21389);
or U21610 (N_21610,N_21189,N_21050);
nand U21611 (N_21611,N_21167,N_21445);
nand U21612 (N_21612,N_21204,N_21094);
nand U21613 (N_21613,N_21414,N_21358);
or U21614 (N_21614,N_21387,N_21408);
xor U21615 (N_21615,N_21278,N_21494);
nor U21616 (N_21616,N_21374,N_21030);
or U21617 (N_21617,N_21209,N_21091);
xor U21618 (N_21618,N_21029,N_21223);
nor U21619 (N_21619,N_21009,N_21088);
xnor U21620 (N_21620,N_21031,N_21498);
xor U21621 (N_21621,N_21075,N_21034);
nand U21622 (N_21622,N_21017,N_21343);
nand U21623 (N_21623,N_21111,N_21249);
and U21624 (N_21624,N_21003,N_21119);
nand U21625 (N_21625,N_21292,N_21286);
and U21626 (N_21626,N_21247,N_21115);
nand U21627 (N_21627,N_21488,N_21421);
xnor U21628 (N_21628,N_21069,N_21039);
and U21629 (N_21629,N_21440,N_21474);
nor U21630 (N_21630,N_21216,N_21297);
xor U21631 (N_21631,N_21145,N_21411);
and U21632 (N_21632,N_21245,N_21100);
xor U21633 (N_21633,N_21267,N_21153);
nor U21634 (N_21634,N_21238,N_21148);
or U21635 (N_21635,N_21481,N_21444);
nor U21636 (N_21636,N_21493,N_21298);
nor U21637 (N_21637,N_21277,N_21271);
or U21638 (N_21638,N_21331,N_21371);
or U21639 (N_21639,N_21218,N_21237);
xnor U21640 (N_21640,N_21469,N_21460);
nand U21641 (N_21641,N_21497,N_21010);
and U21642 (N_21642,N_21341,N_21366);
or U21643 (N_21643,N_21178,N_21214);
and U21644 (N_21644,N_21118,N_21438);
or U21645 (N_21645,N_21205,N_21308);
nor U21646 (N_21646,N_21203,N_21423);
xnor U21647 (N_21647,N_21171,N_21123);
nand U21648 (N_21648,N_21161,N_21250);
nand U21649 (N_21649,N_21181,N_21306);
and U21650 (N_21650,N_21177,N_21491);
and U21651 (N_21651,N_21246,N_21230);
nand U21652 (N_21652,N_21260,N_21136);
and U21653 (N_21653,N_21275,N_21133);
xor U21654 (N_21654,N_21394,N_21452);
nor U21655 (N_21655,N_21456,N_21312);
and U21656 (N_21656,N_21475,N_21056);
nor U21657 (N_21657,N_21021,N_21231);
or U21658 (N_21658,N_21270,N_21261);
and U21659 (N_21659,N_21117,N_21359);
xnor U21660 (N_21660,N_21128,N_21269);
or U21661 (N_21661,N_21375,N_21184);
or U21662 (N_21662,N_21279,N_21125);
nand U21663 (N_21663,N_21134,N_21273);
or U21664 (N_21664,N_21097,N_21196);
nor U21665 (N_21665,N_21291,N_21482);
xor U21666 (N_21666,N_21355,N_21114);
nor U21667 (N_21667,N_21304,N_21352);
or U21668 (N_21668,N_21315,N_21326);
and U21669 (N_21669,N_21398,N_21385);
nor U21670 (N_21670,N_21370,N_21208);
and U21671 (N_21671,N_21362,N_21378);
and U21672 (N_21672,N_21428,N_21154);
or U21673 (N_21673,N_21289,N_21005);
and U21674 (N_21674,N_21235,N_21406);
or U21675 (N_21675,N_21110,N_21104);
nor U21676 (N_21676,N_21468,N_21400);
nand U21677 (N_21677,N_21483,N_21228);
or U21678 (N_21678,N_21013,N_21162);
or U21679 (N_21679,N_21044,N_21376);
xor U21680 (N_21680,N_21492,N_21430);
or U21681 (N_21681,N_21287,N_21354);
xor U21682 (N_21682,N_21051,N_21157);
nor U21683 (N_21683,N_21496,N_21321);
nor U21684 (N_21684,N_21159,N_21062);
and U21685 (N_21685,N_21124,N_21174);
and U21686 (N_21686,N_21240,N_21139);
xnor U21687 (N_21687,N_21426,N_21122);
nand U21688 (N_21688,N_21109,N_21156);
and U21689 (N_21689,N_21403,N_21263);
nand U21690 (N_21690,N_21217,N_21357);
xnor U21691 (N_21691,N_21040,N_21458);
and U21692 (N_21692,N_21038,N_21252);
nand U21693 (N_21693,N_21478,N_21006);
and U21694 (N_21694,N_21175,N_21462);
xnor U21695 (N_21695,N_21198,N_21351);
nand U21696 (N_21696,N_21053,N_21202);
xnor U21697 (N_21697,N_21395,N_21457);
xnor U21698 (N_21698,N_21339,N_21232);
and U21699 (N_21699,N_21004,N_21424);
or U21700 (N_21700,N_21314,N_21042);
nand U21701 (N_21701,N_21195,N_21101);
nand U21702 (N_21702,N_21258,N_21484);
and U21703 (N_21703,N_21186,N_21185);
or U21704 (N_21704,N_21113,N_21045);
and U21705 (N_21705,N_21429,N_21092);
nor U21706 (N_21706,N_21007,N_21451);
and U21707 (N_21707,N_21415,N_21281);
nand U21708 (N_21708,N_21226,N_21404);
or U21709 (N_21709,N_21002,N_21449);
xor U21710 (N_21710,N_21169,N_21105);
or U21711 (N_21711,N_21055,N_21432);
xor U21712 (N_21712,N_21098,N_21402);
nand U21713 (N_21713,N_21067,N_21282);
nand U21714 (N_21714,N_21163,N_21259);
nor U21715 (N_21715,N_21473,N_21465);
nor U21716 (N_21716,N_21323,N_21464);
nor U21717 (N_21717,N_21221,N_21248);
nor U21718 (N_21718,N_21077,N_21399);
nand U21719 (N_21719,N_21233,N_21207);
and U21720 (N_21720,N_21367,N_21043);
or U21721 (N_21721,N_21309,N_21446);
or U21722 (N_21722,N_21166,N_21334);
or U21723 (N_21723,N_21047,N_21417);
and U21724 (N_21724,N_21054,N_21225);
and U21725 (N_21725,N_21347,N_21300);
or U21726 (N_21726,N_21142,N_21340);
nand U21727 (N_21727,N_21401,N_21356);
or U21728 (N_21728,N_21364,N_21466);
nand U21729 (N_21729,N_21274,N_21126);
nand U21730 (N_21730,N_21135,N_21032);
nand U21731 (N_21731,N_21158,N_21419);
nor U21732 (N_21732,N_21489,N_21095);
and U21733 (N_21733,N_21485,N_21188);
nand U21734 (N_21734,N_21313,N_21396);
nor U21735 (N_21735,N_21165,N_21172);
nand U21736 (N_21736,N_21120,N_21076);
xnor U21737 (N_21737,N_21368,N_21455);
xor U21738 (N_21738,N_21036,N_21296);
nand U21739 (N_21739,N_21129,N_21305);
nand U21740 (N_21740,N_21219,N_21463);
nor U21741 (N_21741,N_21299,N_21193);
nor U21742 (N_21742,N_21416,N_21372);
nor U21743 (N_21743,N_21065,N_21302);
or U21744 (N_21744,N_21089,N_21131);
or U21745 (N_21745,N_21001,N_21224);
nand U21746 (N_21746,N_21066,N_21253);
or U21747 (N_21747,N_21405,N_21311);
nor U21748 (N_21748,N_21377,N_21239);
nor U21749 (N_21749,N_21365,N_21320);
nor U21750 (N_21750,N_21455,N_21171);
or U21751 (N_21751,N_21412,N_21139);
or U21752 (N_21752,N_21185,N_21198);
or U21753 (N_21753,N_21311,N_21161);
or U21754 (N_21754,N_21298,N_21305);
and U21755 (N_21755,N_21037,N_21265);
nand U21756 (N_21756,N_21198,N_21202);
nand U21757 (N_21757,N_21014,N_21034);
or U21758 (N_21758,N_21283,N_21477);
nand U21759 (N_21759,N_21162,N_21393);
nor U21760 (N_21760,N_21353,N_21456);
nand U21761 (N_21761,N_21441,N_21155);
or U21762 (N_21762,N_21181,N_21365);
and U21763 (N_21763,N_21182,N_21039);
xnor U21764 (N_21764,N_21083,N_21234);
or U21765 (N_21765,N_21356,N_21063);
and U21766 (N_21766,N_21269,N_21334);
nor U21767 (N_21767,N_21433,N_21457);
nor U21768 (N_21768,N_21109,N_21136);
nor U21769 (N_21769,N_21413,N_21148);
or U21770 (N_21770,N_21400,N_21218);
and U21771 (N_21771,N_21050,N_21445);
and U21772 (N_21772,N_21440,N_21003);
nand U21773 (N_21773,N_21117,N_21139);
nor U21774 (N_21774,N_21415,N_21199);
or U21775 (N_21775,N_21360,N_21480);
xor U21776 (N_21776,N_21482,N_21344);
and U21777 (N_21777,N_21440,N_21336);
or U21778 (N_21778,N_21315,N_21317);
xnor U21779 (N_21779,N_21152,N_21201);
xnor U21780 (N_21780,N_21191,N_21292);
and U21781 (N_21781,N_21337,N_21418);
xor U21782 (N_21782,N_21262,N_21127);
or U21783 (N_21783,N_21272,N_21416);
nand U21784 (N_21784,N_21214,N_21062);
xor U21785 (N_21785,N_21276,N_21136);
and U21786 (N_21786,N_21491,N_21007);
nor U21787 (N_21787,N_21120,N_21147);
nor U21788 (N_21788,N_21343,N_21131);
nor U21789 (N_21789,N_21154,N_21370);
or U21790 (N_21790,N_21461,N_21190);
nand U21791 (N_21791,N_21141,N_21063);
and U21792 (N_21792,N_21356,N_21391);
or U21793 (N_21793,N_21260,N_21023);
xor U21794 (N_21794,N_21410,N_21498);
nand U21795 (N_21795,N_21032,N_21294);
and U21796 (N_21796,N_21055,N_21206);
and U21797 (N_21797,N_21335,N_21354);
nor U21798 (N_21798,N_21422,N_21077);
and U21799 (N_21799,N_21351,N_21156);
or U21800 (N_21800,N_21440,N_21319);
or U21801 (N_21801,N_21286,N_21272);
or U21802 (N_21802,N_21027,N_21428);
nor U21803 (N_21803,N_21198,N_21262);
and U21804 (N_21804,N_21042,N_21259);
nor U21805 (N_21805,N_21058,N_21141);
and U21806 (N_21806,N_21274,N_21016);
xnor U21807 (N_21807,N_21123,N_21305);
or U21808 (N_21808,N_21459,N_21235);
nor U21809 (N_21809,N_21009,N_21368);
or U21810 (N_21810,N_21295,N_21237);
or U21811 (N_21811,N_21037,N_21193);
nor U21812 (N_21812,N_21012,N_21265);
nor U21813 (N_21813,N_21109,N_21201);
or U21814 (N_21814,N_21025,N_21431);
and U21815 (N_21815,N_21408,N_21495);
and U21816 (N_21816,N_21273,N_21192);
xnor U21817 (N_21817,N_21340,N_21041);
xnor U21818 (N_21818,N_21398,N_21000);
nand U21819 (N_21819,N_21212,N_21325);
xnor U21820 (N_21820,N_21073,N_21207);
nor U21821 (N_21821,N_21195,N_21042);
or U21822 (N_21822,N_21186,N_21241);
and U21823 (N_21823,N_21436,N_21169);
nor U21824 (N_21824,N_21248,N_21063);
and U21825 (N_21825,N_21328,N_21259);
nor U21826 (N_21826,N_21227,N_21330);
nor U21827 (N_21827,N_21258,N_21454);
and U21828 (N_21828,N_21216,N_21488);
and U21829 (N_21829,N_21057,N_21252);
nand U21830 (N_21830,N_21222,N_21281);
xnor U21831 (N_21831,N_21127,N_21229);
nor U21832 (N_21832,N_21473,N_21341);
and U21833 (N_21833,N_21479,N_21121);
or U21834 (N_21834,N_21406,N_21490);
or U21835 (N_21835,N_21481,N_21136);
xor U21836 (N_21836,N_21327,N_21039);
nand U21837 (N_21837,N_21132,N_21075);
xor U21838 (N_21838,N_21212,N_21365);
nand U21839 (N_21839,N_21435,N_21430);
nand U21840 (N_21840,N_21471,N_21031);
and U21841 (N_21841,N_21267,N_21291);
and U21842 (N_21842,N_21255,N_21435);
xnor U21843 (N_21843,N_21082,N_21085);
xor U21844 (N_21844,N_21426,N_21108);
xnor U21845 (N_21845,N_21182,N_21185);
nor U21846 (N_21846,N_21325,N_21189);
or U21847 (N_21847,N_21198,N_21071);
xor U21848 (N_21848,N_21304,N_21006);
and U21849 (N_21849,N_21188,N_21408);
and U21850 (N_21850,N_21181,N_21489);
nand U21851 (N_21851,N_21311,N_21341);
nand U21852 (N_21852,N_21334,N_21311);
nand U21853 (N_21853,N_21169,N_21012);
nor U21854 (N_21854,N_21468,N_21293);
xnor U21855 (N_21855,N_21185,N_21201);
and U21856 (N_21856,N_21434,N_21377);
and U21857 (N_21857,N_21071,N_21199);
xnor U21858 (N_21858,N_21438,N_21073);
or U21859 (N_21859,N_21438,N_21478);
nor U21860 (N_21860,N_21384,N_21317);
and U21861 (N_21861,N_21214,N_21405);
nand U21862 (N_21862,N_21133,N_21376);
or U21863 (N_21863,N_21458,N_21382);
and U21864 (N_21864,N_21186,N_21242);
nor U21865 (N_21865,N_21343,N_21051);
nor U21866 (N_21866,N_21346,N_21063);
and U21867 (N_21867,N_21409,N_21096);
nand U21868 (N_21868,N_21320,N_21254);
and U21869 (N_21869,N_21377,N_21309);
xnor U21870 (N_21870,N_21382,N_21111);
nor U21871 (N_21871,N_21181,N_21427);
nand U21872 (N_21872,N_21312,N_21213);
or U21873 (N_21873,N_21121,N_21263);
nor U21874 (N_21874,N_21145,N_21292);
and U21875 (N_21875,N_21166,N_21103);
nor U21876 (N_21876,N_21450,N_21481);
nor U21877 (N_21877,N_21370,N_21190);
or U21878 (N_21878,N_21206,N_21125);
and U21879 (N_21879,N_21249,N_21474);
xnor U21880 (N_21880,N_21321,N_21247);
or U21881 (N_21881,N_21000,N_21135);
nand U21882 (N_21882,N_21205,N_21038);
nor U21883 (N_21883,N_21123,N_21426);
and U21884 (N_21884,N_21018,N_21113);
xnor U21885 (N_21885,N_21209,N_21181);
nor U21886 (N_21886,N_21080,N_21157);
xor U21887 (N_21887,N_21002,N_21020);
xor U21888 (N_21888,N_21480,N_21493);
and U21889 (N_21889,N_21324,N_21106);
nand U21890 (N_21890,N_21261,N_21142);
nand U21891 (N_21891,N_21322,N_21193);
nand U21892 (N_21892,N_21190,N_21051);
xor U21893 (N_21893,N_21215,N_21048);
and U21894 (N_21894,N_21373,N_21444);
or U21895 (N_21895,N_21056,N_21371);
or U21896 (N_21896,N_21410,N_21012);
or U21897 (N_21897,N_21049,N_21039);
nand U21898 (N_21898,N_21397,N_21041);
or U21899 (N_21899,N_21319,N_21240);
nor U21900 (N_21900,N_21033,N_21281);
xnor U21901 (N_21901,N_21268,N_21111);
nor U21902 (N_21902,N_21166,N_21211);
nand U21903 (N_21903,N_21043,N_21140);
nand U21904 (N_21904,N_21392,N_21314);
xnor U21905 (N_21905,N_21479,N_21487);
nand U21906 (N_21906,N_21140,N_21251);
nand U21907 (N_21907,N_21388,N_21239);
nor U21908 (N_21908,N_21225,N_21289);
or U21909 (N_21909,N_21242,N_21165);
nor U21910 (N_21910,N_21278,N_21035);
xor U21911 (N_21911,N_21459,N_21378);
nor U21912 (N_21912,N_21311,N_21395);
and U21913 (N_21913,N_21414,N_21123);
nand U21914 (N_21914,N_21268,N_21238);
nand U21915 (N_21915,N_21009,N_21148);
xor U21916 (N_21916,N_21463,N_21133);
or U21917 (N_21917,N_21440,N_21404);
nor U21918 (N_21918,N_21045,N_21413);
nand U21919 (N_21919,N_21315,N_21290);
or U21920 (N_21920,N_21346,N_21463);
nor U21921 (N_21921,N_21114,N_21077);
xnor U21922 (N_21922,N_21454,N_21027);
and U21923 (N_21923,N_21035,N_21293);
nor U21924 (N_21924,N_21218,N_21111);
and U21925 (N_21925,N_21251,N_21273);
or U21926 (N_21926,N_21066,N_21257);
xnor U21927 (N_21927,N_21098,N_21474);
xor U21928 (N_21928,N_21165,N_21178);
nor U21929 (N_21929,N_21075,N_21193);
nand U21930 (N_21930,N_21213,N_21233);
nand U21931 (N_21931,N_21288,N_21123);
and U21932 (N_21932,N_21173,N_21085);
xor U21933 (N_21933,N_21138,N_21161);
xnor U21934 (N_21934,N_21163,N_21119);
nor U21935 (N_21935,N_21016,N_21197);
xnor U21936 (N_21936,N_21099,N_21043);
and U21937 (N_21937,N_21286,N_21444);
xnor U21938 (N_21938,N_21238,N_21255);
nand U21939 (N_21939,N_21201,N_21475);
xnor U21940 (N_21940,N_21081,N_21160);
and U21941 (N_21941,N_21128,N_21188);
xnor U21942 (N_21942,N_21288,N_21380);
nand U21943 (N_21943,N_21030,N_21490);
and U21944 (N_21944,N_21384,N_21020);
and U21945 (N_21945,N_21046,N_21315);
or U21946 (N_21946,N_21137,N_21430);
or U21947 (N_21947,N_21435,N_21463);
or U21948 (N_21948,N_21143,N_21011);
or U21949 (N_21949,N_21194,N_21196);
or U21950 (N_21950,N_21307,N_21453);
nor U21951 (N_21951,N_21058,N_21215);
and U21952 (N_21952,N_21108,N_21096);
or U21953 (N_21953,N_21178,N_21021);
or U21954 (N_21954,N_21203,N_21279);
xor U21955 (N_21955,N_21113,N_21151);
nand U21956 (N_21956,N_21071,N_21413);
nand U21957 (N_21957,N_21133,N_21014);
and U21958 (N_21958,N_21172,N_21076);
nand U21959 (N_21959,N_21008,N_21362);
and U21960 (N_21960,N_21351,N_21105);
and U21961 (N_21961,N_21195,N_21245);
or U21962 (N_21962,N_21375,N_21239);
nand U21963 (N_21963,N_21121,N_21161);
or U21964 (N_21964,N_21442,N_21175);
xnor U21965 (N_21965,N_21220,N_21421);
nand U21966 (N_21966,N_21255,N_21068);
nor U21967 (N_21967,N_21027,N_21038);
or U21968 (N_21968,N_21424,N_21123);
and U21969 (N_21969,N_21125,N_21275);
nand U21970 (N_21970,N_21468,N_21366);
nand U21971 (N_21971,N_21021,N_21206);
nand U21972 (N_21972,N_21207,N_21397);
and U21973 (N_21973,N_21332,N_21053);
nand U21974 (N_21974,N_21329,N_21009);
nor U21975 (N_21975,N_21046,N_21252);
or U21976 (N_21976,N_21485,N_21155);
nor U21977 (N_21977,N_21032,N_21374);
nand U21978 (N_21978,N_21048,N_21354);
or U21979 (N_21979,N_21210,N_21476);
nand U21980 (N_21980,N_21003,N_21207);
nor U21981 (N_21981,N_21028,N_21030);
or U21982 (N_21982,N_21334,N_21036);
xnor U21983 (N_21983,N_21289,N_21477);
xor U21984 (N_21984,N_21424,N_21270);
or U21985 (N_21985,N_21233,N_21419);
xnor U21986 (N_21986,N_21349,N_21194);
xor U21987 (N_21987,N_21356,N_21484);
nand U21988 (N_21988,N_21138,N_21490);
and U21989 (N_21989,N_21176,N_21077);
xor U21990 (N_21990,N_21201,N_21265);
xnor U21991 (N_21991,N_21129,N_21428);
nand U21992 (N_21992,N_21275,N_21410);
xor U21993 (N_21993,N_21328,N_21450);
or U21994 (N_21994,N_21205,N_21365);
or U21995 (N_21995,N_21293,N_21445);
or U21996 (N_21996,N_21211,N_21067);
nand U21997 (N_21997,N_21168,N_21031);
nand U21998 (N_21998,N_21443,N_21135);
and U21999 (N_21999,N_21163,N_21465);
or U22000 (N_22000,N_21500,N_21646);
or U22001 (N_22001,N_21655,N_21997);
or U22002 (N_22002,N_21845,N_21984);
nor U22003 (N_22003,N_21697,N_21912);
nor U22004 (N_22004,N_21641,N_21792);
nor U22005 (N_22005,N_21994,N_21680);
nor U22006 (N_22006,N_21864,N_21897);
xnor U22007 (N_22007,N_21919,N_21873);
or U22008 (N_22008,N_21776,N_21558);
and U22009 (N_22009,N_21800,N_21632);
xor U22010 (N_22010,N_21764,N_21742);
nand U22011 (N_22011,N_21916,N_21532);
nand U22012 (N_22012,N_21913,N_21585);
and U22013 (N_22013,N_21566,N_21967);
and U22014 (N_22014,N_21601,N_21708);
or U22015 (N_22015,N_21778,N_21723);
nor U22016 (N_22016,N_21827,N_21594);
or U22017 (N_22017,N_21810,N_21672);
nor U22018 (N_22018,N_21665,N_21877);
or U22019 (N_22019,N_21957,N_21750);
nor U22020 (N_22020,N_21917,N_21628);
nand U22021 (N_22021,N_21699,N_21989);
or U22022 (N_22022,N_21551,N_21821);
nand U22023 (N_22023,N_21749,N_21979);
nand U22024 (N_22024,N_21974,N_21740);
or U22025 (N_22025,N_21744,N_21662);
or U22026 (N_22026,N_21563,N_21931);
and U22027 (N_22027,N_21935,N_21629);
nand U22028 (N_22028,N_21714,N_21861);
nor U22029 (N_22029,N_21613,N_21542);
and U22030 (N_22030,N_21941,N_21829);
nand U22031 (N_22031,N_21622,N_21738);
nand U22032 (N_22032,N_21717,N_21898);
xnor U22033 (N_22033,N_21549,N_21734);
or U22034 (N_22034,N_21607,N_21603);
and U22035 (N_22035,N_21999,N_21674);
nand U22036 (N_22036,N_21652,N_21884);
xnor U22037 (N_22037,N_21722,N_21506);
and U22038 (N_22038,N_21528,N_21546);
and U22039 (N_22039,N_21619,N_21715);
or U22040 (N_22040,N_21857,N_21520);
xnor U22041 (N_22041,N_21611,N_21733);
nand U22042 (N_22042,N_21523,N_21605);
and U22043 (N_22043,N_21961,N_21820);
nor U22044 (N_22044,N_21896,N_21779);
nand U22045 (N_22045,N_21858,N_21683);
nor U22046 (N_22046,N_21872,N_21704);
nor U22047 (N_22047,N_21530,N_21850);
and U22048 (N_22048,N_21595,N_21955);
nor U22049 (N_22049,N_21584,N_21654);
nand U22050 (N_22050,N_21910,N_21502);
nor U22051 (N_22051,N_21799,N_21525);
nor U22052 (N_22052,N_21944,N_21824);
and U22053 (N_22053,N_21653,N_21940);
and U22054 (N_22054,N_21785,N_21587);
xor U22055 (N_22055,N_21787,N_21658);
nor U22056 (N_22056,N_21564,N_21735);
nand U22057 (N_22057,N_21968,N_21664);
nand U22058 (N_22058,N_21817,N_21995);
nor U22059 (N_22059,N_21681,N_21721);
or U22060 (N_22060,N_21814,N_21772);
nor U22061 (N_22061,N_21720,N_21909);
xnor U22062 (N_22062,N_21640,N_21795);
xor U22063 (N_22063,N_21951,N_21656);
nand U22064 (N_22064,N_21696,N_21895);
xor U22065 (N_22065,N_21539,N_21701);
nand U22066 (N_22066,N_21887,N_21643);
nand U22067 (N_22067,N_21712,N_21908);
xor U22068 (N_22068,N_21907,N_21876);
nand U22069 (N_22069,N_21782,N_21899);
and U22070 (N_22070,N_21579,N_21561);
nor U22071 (N_22071,N_21920,N_21928);
and U22072 (N_22072,N_21922,N_21947);
nor U22073 (N_22073,N_21702,N_21926);
nand U22074 (N_22074,N_21602,N_21838);
nor U22075 (N_22075,N_21834,N_21988);
and U22076 (N_22076,N_21837,N_21959);
nor U22077 (N_22077,N_21797,N_21668);
or U22078 (N_22078,N_21582,N_21518);
and U22079 (N_22079,N_21533,N_21589);
and U22080 (N_22080,N_21577,N_21915);
xnor U22081 (N_22081,N_21854,N_21962);
nand U22082 (N_22082,N_21842,N_21692);
xor U22083 (N_22083,N_21706,N_21610);
nor U22084 (N_22084,N_21883,N_21774);
and U22085 (N_22085,N_21902,N_21833);
xnor U22086 (N_22086,N_21626,N_21557);
nor U22087 (N_22087,N_21759,N_21853);
xnor U22088 (N_22088,N_21686,N_21828);
nand U22089 (N_22089,N_21536,N_21752);
or U22090 (N_22090,N_21676,N_21921);
nand U22091 (N_22091,N_21559,N_21870);
and U22092 (N_22092,N_21685,N_21630);
or U22093 (N_22093,N_21569,N_21574);
or U22094 (N_22094,N_21946,N_21773);
xnor U22095 (N_22095,N_21540,N_21892);
nor U22096 (N_22096,N_21960,N_21952);
nor U22097 (N_22097,N_21573,N_21783);
nand U22098 (N_22098,N_21729,N_21554);
xnor U22099 (N_22099,N_21975,N_21571);
nand U22100 (N_22100,N_21648,N_21608);
and U22101 (N_22101,N_21966,N_21621);
nand U22102 (N_22102,N_21846,N_21874);
nand U22103 (N_22103,N_21728,N_21812);
or U22104 (N_22104,N_21945,N_21700);
nand U22105 (N_22105,N_21512,N_21516);
and U22106 (N_22106,N_21517,N_21860);
or U22107 (N_22107,N_21878,N_21624);
nand U22108 (N_22108,N_21831,N_21791);
and U22109 (N_22109,N_21599,N_21875);
or U22110 (N_22110,N_21847,N_21793);
or U22111 (N_22111,N_21666,N_21780);
and U22112 (N_22112,N_21527,N_21597);
nand U22113 (N_22113,N_21889,N_21986);
xor U22114 (N_22114,N_21971,N_21775);
nand U22115 (N_22115,N_21830,N_21990);
or U22116 (N_22116,N_21637,N_21852);
nand U22117 (N_22117,N_21803,N_21954);
xor U22118 (N_22118,N_21544,N_21511);
nor U22119 (N_22119,N_21514,N_21911);
or U22120 (N_22120,N_21970,N_21906);
xor U22121 (N_22121,N_21679,N_21562);
and U22122 (N_22122,N_21725,N_21609);
nor U22123 (N_22123,N_21871,N_21900);
and U22124 (N_22124,N_21855,N_21890);
or U22125 (N_22125,N_21592,N_21885);
xnor U22126 (N_22126,N_21600,N_21736);
nand U22127 (N_22127,N_21541,N_21796);
nand U22128 (N_22128,N_21805,N_21649);
and U22129 (N_22129,N_21713,N_21659);
nand U22130 (N_22130,N_21743,N_21567);
nand U22131 (N_22131,N_21925,N_21768);
and U22132 (N_22132,N_21711,N_21556);
nor U22133 (N_22133,N_21623,N_21880);
xor U22134 (N_22134,N_21816,N_21976);
and U22135 (N_22135,N_21586,N_21578);
or U22136 (N_22136,N_21784,N_21770);
or U22137 (N_22137,N_21719,N_21948);
or U22138 (N_22138,N_21843,N_21741);
nor U22139 (N_22139,N_21588,N_21893);
nand U22140 (N_22140,N_21977,N_21918);
or U22141 (N_22141,N_21591,N_21865);
nand U22142 (N_22142,N_21753,N_21548);
nor U22143 (N_22143,N_21866,N_21832);
and U22144 (N_22144,N_21636,N_21509);
xor U22145 (N_22145,N_21781,N_21767);
or U22146 (N_22146,N_21851,N_21901);
nand U22147 (N_22147,N_21580,N_21639);
or U22148 (N_22148,N_21671,N_21507);
or U22149 (N_22149,N_21848,N_21663);
nor U22150 (N_22150,N_21745,N_21691);
xor U22151 (N_22151,N_21612,N_21929);
nor U22152 (N_22152,N_21727,N_21937);
or U22153 (N_22153,N_21992,N_21942);
or U22154 (N_22154,N_21927,N_21684);
and U22155 (N_22155,N_21547,N_21615);
nor U22156 (N_22156,N_21933,N_21703);
and U22157 (N_22157,N_21938,N_21604);
nand U22158 (N_22158,N_21936,N_21746);
xnor U22159 (N_22159,N_21726,N_21981);
and U22160 (N_22160,N_21905,N_21755);
or U22161 (N_22161,N_21560,N_21983);
nand U22162 (N_22162,N_21709,N_21510);
and U22163 (N_22163,N_21661,N_21529);
nand U22164 (N_22164,N_21677,N_21756);
nor U22165 (N_22165,N_21669,N_21982);
nor U22166 (N_22166,N_21969,N_21730);
nor U22167 (N_22167,N_21798,N_21757);
and U22168 (N_22168,N_21687,N_21835);
nor U22169 (N_22169,N_21863,N_21627);
nor U22170 (N_22170,N_21972,N_21934);
nand U22171 (N_22171,N_21524,N_21930);
nand U22172 (N_22172,N_21732,N_21859);
nand U22173 (N_22173,N_21923,N_21570);
nor U22174 (N_22174,N_21645,N_21786);
xor U22175 (N_22175,N_21963,N_21675);
nor U22176 (N_22176,N_21631,N_21788);
nand U22177 (N_22177,N_21739,N_21822);
xor U22178 (N_22178,N_21537,N_21769);
nand U22179 (N_22179,N_21904,N_21598);
xor U22180 (N_22180,N_21705,N_21534);
and U22181 (N_22181,N_21503,N_21504);
nand U22182 (N_22182,N_21932,N_21590);
xnor U22183 (N_22183,N_21678,N_21731);
or U22184 (N_22184,N_21813,N_21924);
or U22185 (N_22185,N_21939,N_21616);
or U22186 (N_22186,N_21758,N_21695);
nor U22187 (N_22187,N_21823,N_21862);
or U22188 (N_22188,N_21555,N_21760);
or U22189 (N_22189,N_21765,N_21638);
nand U22190 (N_22190,N_21707,N_21886);
or U22191 (N_22191,N_21766,N_21980);
xnor U22192 (N_22192,N_21614,N_21596);
xnor U22193 (N_22193,N_21737,N_21505);
nor U22194 (N_22194,N_21515,N_21818);
nor U22195 (N_22195,N_21794,N_21841);
nand U22196 (N_22196,N_21763,N_21958);
nor U22197 (N_22197,N_21943,N_21531);
or U22198 (N_22198,N_21964,N_21844);
nand U22199 (N_22199,N_21762,N_21519);
and U22200 (N_22200,N_21545,N_21693);
nand U22201 (N_22201,N_21815,N_21635);
nand U22202 (N_22202,N_21633,N_21513);
or U22203 (N_22203,N_21973,N_21868);
nor U22204 (N_22204,N_21583,N_21650);
and U22205 (N_22205,N_21985,N_21568);
nor U22206 (N_22206,N_21790,N_21550);
nor U22207 (N_22207,N_21840,N_21751);
and U22208 (N_22208,N_21538,N_21956);
nor U22209 (N_22209,N_21552,N_21521);
nand U22210 (N_22210,N_21949,N_21606);
or U22211 (N_22211,N_21657,N_21993);
or U22212 (N_22212,N_21903,N_21526);
nand U22213 (N_22213,N_21647,N_21882);
xor U22214 (N_22214,N_21618,N_21651);
or U22215 (N_22215,N_21716,N_21501);
nand U22216 (N_22216,N_21522,N_21879);
or U22217 (N_22217,N_21535,N_21804);
nand U22218 (N_22218,N_21710,N_21617);
nand U22219 (N_22219,N_21978,N_21572);
and U22220 (N_22220,N_21688,N_21670);
and U22221 (N_22221,N_21543,N_21620);
xnor U22222 (N_22222,N_21553,N_21811);
nor U22223 (N_22223,N_21826,N_21953);
nand U22224 (N_22224,N_21718,N_21698);
or U22225 (N_22225,N_21806,N_21682);
nor U22226 (N_22226,N_21777,N_21801);
or U22227 (N_22227,N_21667,N_21819);
and U22228 (N_22228,N_21856,N_21565);
xor U22229 (N_22229,N_21576,N_21724);
nand U22230 (N_22230,N_21771,N_21575);
and U22231 (N_22231,N_21642,N_21748);
nand U22232 (N_22232,N_21881,N_21789);
nor U22233 (N_22233,N_21914,N_21809);
nand U22234 (N_22234,N_21987,N_21625);
and U22235 (N_22235,N_21965,N_21849);
xnor U22236 (N_22236,N_21998,N_21808);
xnor U22237 (N_22237,N_21690,N_21694);
or U22238 (N_22238,N_21754,N_21747);
nor U22239 (N_22239,N_21996,N_21894);
nand U22240 (N_22240,N_21634,N_21839);
and U22241 (N_22241,N_21673,N_21689);
nor U22242 (N_22242,N_21888,N_21581);
nand U22243 (N_22243,N_21508,N_21644);
and U22244 (N_22244,N_21807,N_21869);
or U22245 (N_22245,N_21802,N_21825);
xor U22246 (N_22246,N_21950,N_21593);
xnor U22247 (N_22247,N_21891,N_21867);
or U22248 (N_22248,N_21761,N_21836);
nor U22249 (N_22249,N_21660,N_21991);
xor U22250 (N_22250,N_21508,N_21626);
and U22251 (N_22251,N_21858,N_21646);
nor U22252 (N_22252,N_21947,N_21629);
and U22253 (N_22253,N_21680,N_21579);
nor U22254 (N_22254,N_21565,N_21794);
and U22255 (N_22255,N_21593,N_21547);
and U22256 (N_22256,N_21804,N_21706);
or U22257 (N_22257,N_21958,N_21542);
and U22258 (N_22258,N_21873,N_21752);
and U22259 (N_22259,N_21672,N_21643);
and U22260 (N_22260,N_21521,N_21635);
xnor U22261 (N_22261,N_21868,N_21702);
nand U22262 (N_22262,N_21901,N_21897);
xor U22263 (N_22263,N_21752,N_21622);
and U22264 (N_22264,N_21555,N_21857);
nor U22265 (N_22265,N_21828,N_21991);
or U22266 (N_22266,N_21577,N_21510);
xnor U22267 (N_22267,N_21533,N_21603);
nor U22268 (N_22268,N_21961,N_21957);
nand U22269 (N_22269,N_21607,N_21847);
nand U22270 (N_22270,N_21932,N_21957);
and U22271 (N_22271,N_21726,N_21649);
nor U22272 (N_22272,N_21596,N_21919);
nor U22273 (N_22273,N_21720,N_21770);
nand U22274 (N_22274,N_21501,N_21568);
nor U22275 (N_22275,N_21764,N_21823);
nor U22276 (N_22276,N_21599,N_21926);
nand U22277 (N_22277,N_21701,N_21644);
or U22278 (N_22278,N_21998,N_21682);
xnor U22279 (N_22279,N_21536,N_21788);
xor U22280 (N_22280,N_21675,N_21624);
or U22281 (N_22281,N_21789,N_21610);
nor U22282 (N_22282,N_21980,N_21747);
nor U22283 (N_22283,N_21943,N_21787);
and U22284 (N_22284,N_21849,N_21988);
xor U22285 (N_22285,N_21945,N_21507);
or U22286 (N_22286,N_21963,N_21757);
nor U22287 (N_22287,N_21886,N_21749);
xnor U22288 (N_22288,N_21827,N_21943);
nor U22289 (N_22289,N_21796,N_21758);
or U22290 (N_22290,N_21689,N_21792);
nor U22291 (N_22291,N_21978,N_21996);
and U22292 (N_22292,N_21548,N_21714);
xor U22293 (N_22293,N_21510,N_21641);
and U22294 (N_22294,N_21756,N_21940);
nor U22295 (N_22295,N_21565,N_21881);
xor U22296 (N_22296,N_21559,N_21889);
xnor U22297 (N_22297,N_21896,N_21839);
nor U22298 (N_22298,N_21857,N_21708);
nand U22299 (N_22299,N_21713,N_21716);
nand U22300 (N_22300,N_21569,N_21911);
nand U22301 (N_22301,N_21594,N_21595);
and U22302 (N_22302,N_21508,N_21639);
nand U22303 (N_22303,N_21962,N_21807);
nor U22304 (N_22304,N_21917,N_21554);
and U22305 (N_22305,N_21784,N_21767);
or U22306 (N_22306,N_21726,N_21587);
nor U22307 (N_22307,N_21510,N_21597);
nor U22308 (N_22308,N_21859,N_21878);
xnor U22309 (N_22309,N_21623,N_21503);
nor U22310 (N_22310,N_21941,N_21820);
nand U22311 (N_22311,N_21669,N_21636);
nor U22312 (N_22312,N_21666,N_21557);
or U22313 (N_22313,N_21557,N_21740);
nor U22314 (N_22314,N_21746,N_21622);
or U22315 (N_22315,N_21711,N_21910);
xor U22316 (N_22316,N_21524,N_21662);
xor U22317 (N_22317,N_21944,N_21677);
xor U22318 (N_22318,N_21632,N_21705);
xor U22319 (N_22319,N_21582,N_21519);
xor U22320 (N_22320,N_21840,N_21896);
nand U22321 (N_22321,N_21701,N_21819);
xor U22322 (N_22322,N_21527,N_21888);
nand U22323 (N_22323,N_21981,N_21880);
and U22324 (N_22324,N_21552,N_21700);
and U22325 (N_22325,N_21839,N_21908);
and U22326 (N_22326,N_21849,N_21984);
nor U22327 (N_22327,N_21838,N_21595);
nor U22328 (N_22328,N_21523,N_21722);
nand U22329 (N_22329,N_21758,N_21894);
and U22330 (N_22330,N_21757,N_21516);
or U22331 (N_22331,N_21602,N_21939);
xor U22332 (N_22332,N_21722,N_21611);
and U22333 (N_22333,N_21632,N_21587);
and U22334 (N_22334,N_21887,N_21766);
xor U22335 (N_22335,N_21948,N_21724);
xnor U22336 (N_22336,N_21648,N_21855);
and U22337 (N_22337,N_21583,N_21564);
xnor U22338 (N_22338,N_21502,N_21744);
nand U22339 (N_22339,N_21814,N_21735);
nor U22340 (N_22340,N_21983,N_21865);
nor U22341 (N_22341,N_21676,N_21739);
and U22342 (N_22342,N_21586,N_21980);
xor U22343 (N_22343,N_21931,N_21701);
nand U22344 (N_22344,N_21731,N_21998);
or U22345 (N_22345,N_21651,N_21993);
or U22346 (N_22346,N_21998,N_21653);
nor U22347 (N_22347,N_21842,N_21959);
or U22348 (N_22348,N_21519,N_21754);
and U22349 (N_22349,N_21972,N_21929);
or U22350 (N_22350,N_21632,N_21510);
nor U22351 (N_22351,N_21660,N_21745);
xnor U22352 (N_22352,N_21713,N_21617);
or U22353 (N_22353,N_21697,N_21585);
nor U22354 (N_22354,N_21874,N_21955);
or U22355 (N_22355,N_21503,N_21533);
and U22356 (N_22356,N_21518,N_21926);
nor U22357 (N_22357,N_21924,N_21919);
nand U22358 (N_22358,N_21808,N_21755);
nor U22359 (N_22359,N_21926,N_21758);
and U22360 (N_22360,N_21619,N_21606);
xnor U22361 (N_22361,N_21846,N_21864);
or U22362 (N_22362,N_21739,N_21966);
and U22363 (N_22363,N_21611,N_21684);
or U22364 (N_22364,N_21875,N_21831);
nor U22365 (N_22365,N_21577,N_21901);
and U22366 (N_22366,N_21879,N_21876);
nor U22367 (N_22367,N_21501,N_21768);
or U22368 (N_22368,N_21611,N_21726);
or U22369 (N_22369,N_21923,N_21833);
nand U22370 (N_22370,N_21733,N_21538);
or U22371 (N_22371,N_21685,N_21637);
and U22372 (N_22372,N_21623,N_21818);
or U22373 (N_22373,N_21909,N_21896);
and U22374 (N_22374,N_21701,N_21867);
nand U22375 (N_22375,N_21805,N_21610);
xnor U22376 (N_22376,N_21777,N_21882);
and U22377 (N_22377,N_21933,N_21784);
and U22378 (N_22378,N_21630,N_21701);
nor U22379 (N_22379,N_21852,N_21901);
xor U22380 (N_22380,N_21680,N_21521);
nor U22381 (N_22381,N_21918,N_21894);
nor U22382 (N_22382,N_21815,N_21734);
xnor U22383 (N_22383,N_21601,N_21609);
or U22384 (N_22384,N_21595,N_21522);
or U22385 (N_22385,N_21955,N_21902);
nand U22386 (N_22386,N_21791,N_21661);
or U22387 (N_22387,N_21517,N_21633);
or U22388 (N_22388,N_21507,N_21726);
nor U22389 (N_22389,N_21650,N_21805);
or U22390 (N_22390,N_21658,N_21544);
xnor U22391 (N_22391,N_21815,N_21824);
xnor U22392 (N_22392,N_21786,N_21830);
nand U22393 (N_22393,N_21807,N_21821);
or U22394 (N_22394,N_21631,N_21626);
nand U22395 (N_22395,N_21802,N_21877);
nand U22396 (N_22396,N_21879,N_21791);
xor U22397 (N_22397,N_21819,N_21517);
nand U22398 (N_22398,N_21871,N_21745);
or U22399 (N_22399,N_21755,N_21691);
or U22400 (N_22400,N_21955,N_21916);
and U22401 (N_22401,N_21630,N_21505);
xor U22402 (N_22402,N_21880,N_21515);
nor U22403 (N_22403,N_21990,N_21975);
or U22404 (N_22404,N_21826,N_21512);
nor U22405 (N_22405,N_21725,N_21556);
nor U22406 (N_22406,N_21842,N_21697);
or U22407 (N_22407,N_21564,N_21568);
or U22408 (N_22408,N_21961,N_21789);
nand U22409 (N_22409,N_21619,N_21694);
nor U22410 (N_22410,N_21968,N_21685);
nor U22411 (N_22411,N_21844,N_21697);
and U22412 (N_22412,N_21547,N_21893);
nand U22413 (N_22413,N_21902,N_21840);
nand U22414 (N_22414,N_21507,N_21915);
nand U22415 (N_22415,N_21707,N_21772);
xor U22416 (N_22416,N_21500,N_21768);
xnor U22417 (N_22417,N_21875,N_21924);
nor U22418 (N_22418,N_21511,N_21912);
or U22419 (N_22419,N_21574,N_21586);
nand U22420 (N_22420,N_21568,N_21982);
and U22421 (N_22421,N_21668,N_21809);
or U22422 (N_22422,N_21530,N_21848);
or U22423 (N_22423,N_21965,N_21644);
or U22424 (N_22424,N_21773,N_21742);
xnor U22425 (N_22425,N_21781,N_21507);
and U22426 (N_22426,N_21834,N_21518);
nor U22427 (N_22427,N_21874,N_21867);
and U22428 (N_22428,N_21676,N_21705);
and U22429 (N_22429,N_21928,N_21900);
nor U22430 (N_22430,N_21771,N_21577);
and U22431 (N_22431,N_21536,N_21572);
or U22432 (N_22432,N_21998,N_21897);
and U22433 (N_22433,N_21600,N_21585);
nand U22434 (N_22434,N_21699,N_21883);
or U22435 (N_22435,N_21987,N_21778);
nand U22436 (N_22436,N_21737,N_21664);
xor U22437 (N_22437,N_21827,N_21704);
or U22438 (N_22438,N_21933,N_21794);
nand U22439 (N_22439,N_21609,N_21829);
nand U22440 (N_22440,N_21862,N_21898);
nor U22441 (N_22441,N_21794,N_21905);
xnor U22442 (N_22442,N_21989,N_21625);
nand U22443 (N_22443,N_21997,N_21892);
xor U22444 (N_22444,N_21944,N_21562);
xnor U22445 (N_22445,N_21931,N_21999);
xnor U22446 (N_22446,N_21704,N_21748);
nor U22447 (N_22447,N_21823,N_21706);
and U22448 (N_22448,N_21572,N_21595);
nand U22449 (N_22449,N_21696,N_21502);
and U22450 (N_22450,N_21955,N_21935);
and U22451 (N_22451,N_21942,N_21622);
nor U22452 (N_22452,N_21703,N_21853);
xor U22453 (N_22453,N_21687,N_21536);
xor U22454 (N_22454,N_21910,N_21556);
or U22455 (N_22455,N_21513,N_21580);
nand U22456 (N_22456,N_21877,N_21830);
xor U22457 (N_22457,N_21676,N_21835);
xnor U22458 (N_22458,N_21707,N_21765);
xor U22459 (N_22459,N_21579,N_21910);
nand U22460 (N_22460,N_21738,N_21632);
or U22461 (N_22461,N_21567,N_21579);
nor U22462 (N_22462,N_21810,N_21669);
xor U22463 (N_22463,N_21717,N_21951);
and U22464 (N_22464,N_21846,N_21948);
xnor U22465 (N_22465,N_21810,N_21553);
or U22466 (N_22466,N_21954,N_21722);
and U22467 (N_22467,N_21669,N_21834);
nand U22468 (N_22468,N_21815,N_21518);
or U22469 (N_22469,N_21565,N_21527);
nor U22470 (N_22470,N_21659,N_21751);
or U22471 (N_22471,N_21850,N_21734);
or U22472 (N_22472,N_21648,N_21585);
or U22473 (N_22473,N_21950,N_21571);
and U22474 (N_22474,N_21543,N_21529);
and U22475 (N_22475,N_21952,N_21771);
nor U22476 (N_22476,N_21521,N_21582);
or U22477 (N_22477,N_21851,N_21619);
xor U22478 (N_22478,N_21673,N_21814);
xor U22479 (N_22479,N_21748,N_21590);
xnor U22480 (N_22480,N_21503,N_21927);
and U22481 (N_22481,N_21502,N_21550);
or U22482 (N_22482,N_21915,N_21713);
xnor U22483 (N_22483,N_21532,N_21755);
nor U22484 (N_22484,N_21900,N_21930);
or U22485 (N_22485,N_21913,N_21680);
and U22486 (N_22486,N_21616,N_21933);
or U22487 (N_22487,N_21572,N_21680);
nor U22488 (N_22488,N_21759,N_21869);
nand U22489 (N_22489,N_21575,N_21789);
and U22490 (N_22490,N_21785,N_21741);
nor U22491 (N_22491,N_21726,N_21887);
nor U22492 (N_22492,N_21714,N_21889);
nand U22493 (N_22493,N_21875,N_21762);
nor U22494 (N_22494,N_21602,N_21764);
nor U22495 (N_22495,N_21954,N_21967);
nand U22496 (N_22496,N_21501,N_21681);
or U22497 (N_22497,N_21863,N_21818);
nor U22498 (N_22498,N_21995,N_21806);
nor U22499 (N_22499,N_21602,N_21903);
nand U22500 (N_22500,N_22453,N_22041);
and U22501 (N_22501,N_22447,N_22217);
and U22502 (N_22502,N_22036,N_22305);
xnor U22503 (N_22503,N_22261,N_22027);
xnor U22504 (N_22504,N_22039,N_22426);
nor U22505 (N_22505,N_22363,N_22270);
nand U22506 (N_22506,N_22365,N_22196);
and U22507 (N_22507,N_22372,N_22263);
and U22508 (N_22508,N_22090,N_22244);
nand U22509 (N_22509,N_22064,N_22197);
and U22510 (N_22510,N_22351,N_22257);
xor U22511 (N_22511,N_22369,N_22038);
and U22512 (N_22512,N_22304,N_22419);
nor U22513 (N_22513,N_22017,N_22336);
and U22514 (N_22514,N_22403,N_22104);
xnor U22515 (N_22515,N_22326,N_22170);
nand U22516 (N_22516,N_22012,N_22292);
nand U22517 (N_22517,N_22226,N_22433);
or U22518 (N_22518,N_22281,N_22457);
nor U22519 (N_22519,N_22271,N_22138);
or U22520 (N_22520,N_22449,N_22398);
nor U22521 (N_22521,N_22025,N_22044);
nand U22522 (N_22522,N_22497,N_22330);
xnor U22523 (N_22523,N_22215,N_22240);
nand U22524 (N_22524,N_22420,N_22030);
nor U22525 (N_22525,N_22461,N_22362);
or U22526 (N_22526,N_22052,N_22317);
and U22527 (N_22527,N_22357,N_22278);
or U22528 (N_22528,N_22496,N_22258);
xnor U22529 (N_22529,N_22190,N_22051);
nor U22530 (N_22530,N_22004,N_22061);
nor U22531 (N_22531,N_22283,N_22349);
or U22532 (N_22532,N_22286,N_22432);
or U22533 (N_22533,N_22247,N_22152);
xnor U22534 (N_22534,N_22473,N_22075);
xor U22535 (N_22535,N_22467,N_22415);
and U22536 (N_22536,N_22289,N_22183);
and U22537 (N_22537,N_22153,N_22301);
nand U22538 (N_22538,N_22213,N_22356);
nor U22539 (N_22539,N_22414,N_22282);
nor U22540 (N_22540,N_22484,N_22311);
and U22541 (N_22541,N_22423,N_22245);
nand U22542 (N_22542,N_22162,N_22057);
nand U22543 (N_22543,N_22337,N_22216);
xnor U22544 (N_22544,N_22042,N_22268);
and U22545 (N_22545,N_22462,N_22296);
nand U22546 (N_22546,N_22425,N_22407);
and U22547 (N_22547,N_22063,N_22413);
nand U22548 (N_22548,N_22358,N_22237);
or U22549 (N_22549,N_22127,N_22018);
and U22550 (N_22550,N_22177,N_22010);
nand U22551 (N_22551,N_22024,N_22359);
and U22552 (N_22552,N_22174,N_22302);
or U22553 (N_22553,N_22463,N_22115);
and U22554 (N_22554,N_22055,N_22441);
nor U22555 (N_22555,N_22102,N_22070);
or U22556 (N_22556,N_22435,N_22404);
nand U22557 (N_22557,N_22318,N_22327);
nand U22558 (N_22558,N_22384,N_22109);
nand U22559 (N_22559,N_22002,N_22037);
nand U22560 (N_22560,N_22067,N_22122);
nand U22561 (N_22561,N_22130,N_22011);
xor U22562 (N_22562,N_22253,N_22401);
or U22563 (N_22563,N_22287,N_22186);
nand U22564 (N_22564,N_22192,N_22243);
or U22565 (N_22565,N_22066,N_22139);
and U22566 (N_22566,N_22267,N_22176);
or U22567 (N_22567,N_22150,N_22074);
nor U22568 (N_22568,N_22344,N_22440);
or U22569 (N_22569,N_22393,N_22182);
or U22570 (N_22570,N_22254,N_22079);
nor U22571 (N_22571,N_22342,N_22092);
nand U22572 (N_22572,N_22009,N_22133);
nand U22573 (N_22573,N_22233,N_22123);
nor U22574 (N_22574,N_22339,N_22083);
or U22575 (N_22575,N_22489,N_22178);
and U22576 (N_22576,N_22208,N_22137);
xor U22577 (N_22577,N_22439,N_22181);
nor U22578 (N_22578,N_22347,N_22128);
or U22579 (N_22579,N_22495,N_22389);
and U22580 (N_22580,N_22029,N_22147);
nand U22581 (N_22581,N_22350,N_22218);
nand U22582 (N_22582,N_22214,N_22341);
nor U22583 (N_22583,N_22144,N_22246);
nor U22584 (N_22584,N_22205,N_22101);
nor U22585 (N_22585,N_22402,N_22200);
and U22586 (N_22586,N_22396,N_22360);
or U22587 (N_22587,N_22048,N_22418);
xnor U22588 (N_22588,N_22154,N_22234);
or U22589 (N_22589,N_22265,N_22417);
or U22590 (N_22590,N_22185,N_22000);
nor U22591 (N_22591,N_22272,N_22368);
nor U22592 (N_22592,N_22284,N_22448);
nand U22593 (N_22593,N_22442,N_22405);
or U22594 (N_22594,N_22071,N_22392);
or U22595 (N_22595,N_22498,N_22468);
and U22596 (N_22596,N_22033,N_22175);
or U22597 (N_22597,N_22231,N_22077);
nand U22598 (N_22598,N_22209,N_22391);
xor U22599 (N_22599,N_22266,N_22285);
nor U22600 (N_22600,N_22416,N_22187);
xor U22601 (N_22601,N_22431,N_22082);
and U22602 (N_22602,N_22219,N_22161);
xor U22603 (N_22603,N_22164,N_22295);
and U22604 (N_22604,N_22494,N_22100);
xor U22605 (N_22605,N_22276,N_22471);
nand U22606 (N_22606,N_22179,N_22103);
nand U22607 (N_22607,N_22236,N_22450);
nand U22608 (N_22608,N_22492,N_22483);
nand U22609 (N_22609,N_22470,N_22015);
nor U22610 (N_22610,N_22238,N_22445);
and U22611 (N_22611,N_22166,N_22195);
xnor U22612 (N_22612,N_22202,N_22212);
nor U22613 (N_22613,N_22141,N_22379);
nand U22614 (N_22614,N_22062,N_22228);
nor U22615 (N_22615,N_22001,N_22499);
or U22616 (N_22616,N_22366,N_22280);
and U22617 (N_22617,N_22068,N_22333);
nand U22618 (N_22618,N_22400,N_22045);
xor U22619 (N_22619,N_22399,N_22163);
xnor U22620 (N_22620,N_22008,N_22262);
or U22621 (N_22621,N_22408,N_22348);
or U22622 (N_22622,N_22198,N_22095);
or U22623 (N_22623,N_22383,N_22054);
xor U22624 (N_22624,N_22140,N_22136);
and U22625 (N_22625,N_22475,N_22387);
and U22626 (N_22626,N_22151,N_22260);
nand U22627 (N_22627,N_22110,N_22478);
nand U22628 (N_22628,N_22412,N_22020);
nand U22629 (N_22629,N_22080,N_22006);
and U22630 (N_22630,N_22375,N_22376);
and U22631 (N_22631,N_22021,N_22129);
nor U22632 (N_22632,N_22394,N_22224);
nand U22633 (N_22633,N_22316,N_22466);
nand U22634 (N_22634,N_22211,N_22108);
xnor U22635 (N_22635,N_22487,N_22331);
xnor U22636 (N_22636,N_22003,N_22374);
nand U22637 (N_22637,N_22474,N_22320);
and U22638 (N_22638,N_22235,N_22116);
and U22639 (N_22639,N_22220,N_22364);
or U22640 (N_22640,N_22321,N_22355);
nand U22641 (N_22641,N_22091,N_22410);
or U22642 (N_22642,N_22146,N_22105);
xor U22643 (N_22643,N_22345,N_22016);
nand U22644 (N_22644,N_22315,N_22455);
and U22645 (N_22645,N_22274,N_22112);
xnor U22646 (N_22646,N_22319,N_22210);
or U22647 (N_22647,N_22193,N_22157);
nor U22648 (N_22648,N_22132,N_22451);
and U22649 (N_22649,N_22159,N_22490);
nand U22650 (N_22650,N_22291,N_22436);
nor U22651 (N_22651,N_22397,N_22421);
and U22652 (N_22652,N_22134,N_22242);
nor U22653 (N_22653,N_22297,N_22120);
and U22654 (N_22654,N_22354,N_22361);
xnor U22655 (N_22655,N_22443,N_22032);
nand U22656 (N_22656,N_22332,N_22329);
and U22657 (N_22657,N_22371,N_22382);
nand U22658 (N_22658,N_22458,N_22346);
and U22659 (N_22659,N_22126,N_22013);
nand U22660 (N_22660,N_22078,N_22251);
nand U22661 (N_22661,N_22023,N_22098);
and U22662 (N_22662,N_22111,N_22125);
nor U22663 (N_22663,N_22249,N_22294);
or U22664 (N_22664,N_22084,N_22485);
or U22665 (N_22665,N_22491,N_22460);
or U22666 (N_22666,N_22093,N_22022);
xnor U22667 (N_22667,N_22203,N_22241);
and U22668 (N_22668,N_22239,N_22121);
nand U22669 (N_22669,N_22299,N_22381);
xnor U22670 (N_22670,N_22380,N_22476);
or U22671 (N_22671,N_22264,N_22480);
nand U22672 (N_22672,N_22060,N_22288);
or U22673 (N_22673,N_22142,N_22043);
nor U22674 (N_22674,N_22259,N_22169);
nand U22675 (N_22675,N_22388,N_22118);
or U22676 (N_22676,N_22145,N_22135);
nor U22677 (N_22677,N_22089,N_22386);
nor U22678 (N_22678,N_22300,N_22156);
and U22679 (N_22679,N_22189,N_22230);
or U22680 (N_22680,N_22081,N_22221);
or U22681 (N_22681,N_22312,N_22201);
or U22682 (N_22682,N_22028,N_22073);
nand U22683 (N_22683,N_22303,N_22390);
or U22684 (N_22684,N_22086,N_22378);
and U22685 (N_22685,N_22155,N_22464);
and U22686 (N_22686,N_22085,N_22308);
nor U22687 (N_22687,N_22456,N_22422);
and U22688 (N_22688,N_22465,N_22310);
nor U22689 (N_22689,N_22325,N_22005);
or U22690 (N_22690,N_22059,N_22222);
and U22691 (N_22691,N_22056,N_22395);
nand U22692 (N_22692,N_22046,N_22385);
nor U22693 (N_22693,N_22184,N_22314);
xor U22694 (N_22694,N_22477,N_22409);
xor U22695 (N_22695,N_22481,N_22148);
or U22696 (N_22696,N_22087,N_22065);
xor U22697 (N_22697,N_22293,N_22309);
or U22698 (N_22698,N_22223,N_22275);
or U22699 (N_22699,N_22113,N_22072);
and U22700 (N_22700,N_22107,N_22097);
and U22701 (N_22701,N_22227,N_22047);
or U22702 (N_22702,N_22049,N_22279);
xnor U22703 (N_22703,N_22277,N_22406);
nand U22704 (N_22704,N_22007,N_22437);
xnor U22705 (N_22705,N_22199,N_22096);
xor U22706 (N_22706,N_22273,N_22167);
or U22707 (N_22707,N_22119,N_22207);
or U22708 (N_22708,N_22035,N_22014);
and U22709 (N_22709,N_22307,N_22088);
or U22710 (N_22710,N_22324,N_22250);
or U22711 (N_22711,N_22173,N_22313);
nor U22712 (N_22712,N_22143,N_22069);
xnor U22713 (N_22713,N_22298,N_22444);
xnor U22714 (N_22714,N_22031,N_22290);
and U22715 (N_22715,N_22367,N_22114);
nor U22716 (N_22716,N_22335,N_22053);
xnor U22717 (N_22717,N_22430,N_22323);
xnor U22718 (N_22718,N_22117,N_22131);
or U22719 (N_22719,N_22434,N_22165);
and U22720 (N_22720,N_22191,N_22438);
xor U22721 (N_22721,N_22269,N_22172);
and U22722 (N_22722,N_22482,N_22411);
nor U22723 (N_22723,N_22171,N_22019);
xor U22724 (N_22724,N_22188,N_22076);
and U22725 (N_22725,N_22424,N_22454);
and U22726 (N_22726,N_22429,N_22168);
or U22727 (N_22727,N_22428,N_22058);
or U22728 (N_22728,N_22486,N_22232);
nand U22729 (N_22729,N_22334,N_22459);
nand U22730 (N_22730,N_22452,N_22050);
nor U22731 (N_22731,N_22488,N_22328);
and U22732 (N_22732,N_22343,N_22149);
or U22733 (N_22733,N_22352,N_22040);
nor U22734 (N_22734,N_22353,N_22340);
and U22735 (N_22735,N_22180,N_22469);
nor U22736 (N_22736,N_22493,N_22370);
nor U22737 (N_22737,N_22446,N_22248);
xnor U22738 (N_22738,N_22472,N_22206);
or U22739 (N_22739,N_22225,N_22373);
nor U22740 (N_22740,N_22094,N_22479);
nor U22741 (N_22741,N_22158,N_22229);
xor U22742 (N_22742,N_22306,N_22204);
and U22743 (N_22743,N_22338,N_22427);
xnor U22744 (N_22744,N_22160,N_22034);
nor U22745 (N_22745,N_22124,N_22194);
nand U22746 (N_22746,N_22377,N_22322);
and U22747 (N_22747,N_22252,N_22255);
or U22748 (N_22748,N_22099,N_22106);
or U22749 (N_22749,N_22256,N_22026);
and U22750 (N_22750,N_22447,N_22177);
and U22751 (N_22751,N_22457,N_22458);
nand U22752 (N_22752,N_22059,N_22241);
nor U22753 (N_22753,N_22331,N_22485);
xor U22754 (N_22754,N_22246,N_22182);
nand U22755 (N_22755,N_22146,N_22087);
nor U22756 (N_22756,N_22168,N_22490);
nor U22757 (N_22757,N_22099,N_22072);
nand U22758 (N_22758,N_22425,N_22370);
xor U22759 (N_22759,N_22489,N_22000);
xor U22760 (N_22760,N_22055,N_22313);
xnor U22761 (N_22761,N_22279,N_22343);
nor U22762 (N_22762,N_22335,N_22327);
or U22763 (N_22763,N_22388,N_22328);
or U22764 (N_22764,N_22281,N_22393);
xor U22765 (N_22765,N_22000,N_22441);
xor U22766 (N_22766,N_22338,N_22191);
or U22767 (N_22767,N_22051,N_22339);
nor U22768 (N_22768,N_22086,N_22194);
nor U22769 (N_22769,N_22319,N_22105);
nand U22770 (N_22770,N_22466,N_22255);
or U22771 (N_22771,N_22408,N_22163);
nor U22772 (N_22772,N_22197,N_22182);
or U22773 (N_22773,N_22310,N_22233);
and U22774 (N_22774,N_22447,N_22070);
xor U22775 (N_22775,N_22057,N_22286);
or U22776 (N_22776,N_22149,N_22427);
nand U22777 (N_22777,N_22324,N_22260);
nand U22778 (N_22778,N_22414,N_22399);
nand U22779 (N_22779,N_22457,N_22210);
xnor U22780 (N_22780,N_22408,N_22256);
or U22781 (N_22781,N_22121,N_22411);
nor U22782 (N_22782,N_22009,N_22291);
and U22783 (N_22783,N_22279,N_22453);
nor U22784 (N_22784,N_22478,N_22042);
nand U22785 (N_22785,N_22492,N_22417);
or U22786 (N_22786,N_22204,N_22344);
and U22787 (N_22787,N_22154,N_22268);
xor U22788 (N_22788,N_22441,N_22122);
and U22789 (N_22789,N_22003,N_22407);
or U22790 (N_22790,N_22289,N_22122);
nor U22791 (N_22791,N_22030,N_22388);
or U22792 (N_22792,N_22160,N_22319);
nor U22793 (N_22793,N_22029,N_22174);
nor U22794 (N_22794,N_22428,N_22145);
nor U22795 (N_22795,N_22314,N_22122);
nor U22796 (N_22796,N_22490,N_22477);
nand U22797 (N_22797,N_22150,N_22487);
xor U22798 (N_22798,N_22338,N_22388);
xor U22799 (N_22799,N_22475,N_22175);
or U22800 (N_22800,N_22162,N_22329);
nor U22801 (N_22801,N_22064,N_22321);
nand U22802 (N_22802,N_22336,N_22060);
and U22803 (N_22803,N_22335,N_22185);
and U22804 (N_22804,N_22187,N_22158);
nand U22805 (N_22805,N_22178,N_22078);
nor U22806 (N_22806,N_22460,N_22058);
nor U22807 (N_22807,N_22071,N_22106);
and U22808 (N_22808,N_22464,N_22066);
and U22809 (N_22809,N_22321,N_22381);
or U22810 (N_22810,N_22358,N_22329);
or U22811 (N_22811,N_22235,N_22328);
xnor U22812 (N_22812,N_22268,N_22490);
nor U22813 (N_22813,N_22199,N_22321);
nand U22814 (N_22814,N_22214,N_22038);
or U22815 (N_22815,N_22164,N_22052);
or U22816 (N_22816,N_22423,N_22148);
and U22817 (N_22817,N_22362,N_22169);
or U22818 (N_22818,N_22064,N_22180);
or U22819 (N_22819,N_22436,N_22385);
nand U22820 (N_22820,N_22112,N_22031);
nor U22821 (N_22821,N_22449,N_22040);
nor U22822 (N_22822,N_22071,N_22240);
and U22823 (N_22823,N_22142,N_22488);
or U22824 (N_22824,N_22434,N_22448);
nand U22825 (N_22825,N_22387,N_22312);
nor U22826 (N_22826,N_22136,N_22061);
nand U22827 (N_22827,N_22126,N_22355);
nor U22828 (N_22828,N_22494,N_22404);
nand U22829 (N_22829,N_22304,N_22238);
or U22830 (N_22830,N_22208,N_22183);
xor U22831 (N_22831,N_22368,N_22242);
xnor U22832 (N_22832,N_22081,N_22379);
xor U22833 (N_22833,N_22243,N_22392);
or U22834 (N_22834,N_22211,N_22135);
nor U22835 (N_22835,N_22034,N_22436);
nor U22836 (N_22836,N_22385,N_22253);
and U22837 (N_22837,N_22031,N_22421);
xnor U22838 (N_22838,N_22277,N_22481);
or U22839 (N_22839,N_22036,N_22078);
nor U22840 (N_22840,N_22238,N_22213);
and U22841 (N_22841,N_22389,N_22485);
or U22842 (N_22842,N_22091,N_22292);
xnor U22843 (N_22843,N_22224,N_22201);
nand U22844 (N_22844,N_22007,N_22170);
or U22845 (N_22845,N_22035,N_22365);
xnor U22846 (N_22846,N_22482,N_22095);
nor U22847 (N_22847,N_22053,N_22466);
or U22848 (N_22848,N_22215,N_22042);
nor U22849 (N_22849,N_22360,N_22466);
xor U22850 (N_22850,N_22481,N_22082);
nor U22851 (N_22851,N_22065,N_22305);
or U22852 (N_22852,N_22382,N_22236);
nor U22853 (N_22853,N_22067,N_22214);
or U22854 (N_22854,N_22478,N_22010);
nand U22855 (N_22855,N_22226,N_22332);
and U22856 (N_22856,N_22095,N_22085);
or U22857 (N_22857,N_22027,N_22039);
xor U22858 (N_22858,N_22146,N_22280);
xnor U22859 (N_22859,N_22401,N_22057);
nor U22860 (N_22860,N_22314,N_22483);
nor U22861 (N_22861,N_22228,N_22054);
nand U22862 (N_22862,N_22197,N_22013);
or U22863 (N_22863,N_22039,N_22068);
nand U22864 (N_22864,N_22282,N_22025);
nor U22865 (N_22865,N_22112,N_22451);
or U22866 (N_22866,N_22164,N_22350);
xor U22867 (N_22867,N_22382,N_22191);
nor U22868 (N_22868,N_22051,N_22013);
xnor U22869 (N_22869,N_22082,N_22340);
or U22870 (N_22870,N_22055,N_22489);
xnor U22871 (N_22871,N_22010,N_22492);
nor U22872 (N_22872,N_22184,N_22027);
and U22873 (N_22873,N_22140,N_22424);
nand U22874 (N_22874,N_22302,N_22204);
or U22875 (N_22875,N_22308,N_22267);
and U22876 (N_22876,N_22126,N_22271);
and U22877 (N_22877,N_22444,N_22241);
or U22878 (N_22878,N_22175,N_22435);
nand U22879 (N_22879,N_22042,N_22476);
or U22880 (N_22880,N_22141,N_22036);
nor U22881 (N_22881,N_22274,N_22336);
or U22882 (N_22882,N_22065,N_22169);
nand U22883 (N_22883,N_22446,N_22487);
xnor U22884 (N_22884,N_22109,N_22041);
nand U22885 (N_22885,N_22342,N_22335);
xnor U22886 (N_22886,N_22325,N_22271);
nand U22887 (N_22887,N_22389,N_22207);
or U22888 (N_22888,N_22203,N_22127);
nand U22889 (N_22889,N_22212,N_22397);
and U22890 (N_22890,N_22476,N_22132);
and U22891 (N_22891,N_22302,N_22449);
nor U22892 (N_22892,N_22291,N_22303);
xor U22893 (N_22893,N_22057,N_22426);
nor U22894 (N_22894,N_22298,N_22306);
nor U22895 (N_22895,N_22227,N_22424);
nand U22896 (N_22896,N_22465,N_22116);
nor U22897 (N_22897,N_22347,N_22293);
or U22898 (N_22898,N_22130,N_22014);
nor U22899 (N_22899,N_22081,N_22020);
nor U22900 (N_22900,N_22414,N_22093);
nor U22901 (N_22901,N_22088,N_22240);
or U22902 (N_22902,N_22208,N_22159);
nor U22903 (N_22903,N_22138,N_22306);
xnor U22904 (N_22904,N_22083,N_22208);
xnor U22905 (N_22905,N_22488,N_22189);
xor U22906 (N_22906,N_22343,N_22454);
nor U22907 (N_22907,N_22049,N_22412);
nand U22908 (N_22908,N_22071,N_22284);
nor U22909 (N_22909,N_22119,N_22382);
xnor U22910 (N_22910,N_22218,N_22065);
nor U22911 (N_22911,N_22402,N_22323);
nand U22912 (N_22912,N_22188,N_22207);
or U22913 (N_22913,N_22344,N_22323);
or U22914 (N_22914,N_22365,N_22140);
and U22915 (N_22915,N_22174,N_22244);
nor U22916 (N_22916,N_22396,N_22326);
nand U22917 (N_22917,N_22381,N_22049);
nand U22918 (N_22918,N_22222,N_22154);
xnor U22919 (N_22919,N_22070,N_22010);
nand U22920 (N_22920,N_22407,N_22362);
nor U22921 (N_22921,N_22466,N_22224);
nor U22922 (N_22922,N_22399,N_22405);
nor U22923 (N_22923,N_22431,N_22418);
nor U22924 (N_22924,N_22343,N_22119);
xnor U22925 (N_22925,N_22406,N_22297);
and U22926 (N_22926,N_22345,N_22066);
nand U22927 (N_22927,N_22366,N_22277);
and U22928 (N_22928,N_22374,N_22407);
nor U22929 (N_22929,N_22432,N_22272);
xor U22930 (N_22930,N_22408,N_22005);
xnor U22931 (N_22931,N_22348,N_22480);
xor U22932 (N_22932,N_22113,N_22041);
and U22933 (N_22933,N_22223,N_22016);
and U22934 (N_22934,N_22351,N_22371);
xnor U22935 (N_22935,N_22154,N_22315);
xnor U22936 (N_22936,N_22367,N_22428);
nor U22937 (N_22937,N_22496,N_22472);
and U22938 (N_22938,N_22159,N_22328);
and U22939 (N_22939,N_22287,N_22020);
or U22940 (N_22940,N_22221,N_22258);
or U22941 (N_22941,N_22418,N_22408);
nand U22942 (N_22942,N_22227,N_22003);
xnor U22943 (N_22943,N_22058,N_22370);
or U22944 (N_22944,N_22244,N_22268);
and U22945 (N_22945,N_22257,N_22168);
nand U22946 (N_22946,N_22174,N_22436);
nand U22947 (N_22947,N_22171,N_22203);
and U22948 (N_22948,N_22468,N_22119);
and U22949 (N_22949,N_22439,N_22497);
nor U22950 (N_22950,N_22340,N_22027);
or U22951 (N_22951,N_22482,N_22371);
and U22952 (N_22952,N_22103,N_22493);
nand U22953 (N_22953,N_22075,N_22175);
nor U22954 (N_22954,N_22267,N_22285);
or U22955 (N_22955,N_22364,N_22238);
nor U22956 (N_22956,N_22408,N_22071);
or U22957 (N_22957,N_22412,N_22212);
nand U22958 (N_22958,N_22306,N_22389);
or U22959 (N_22959,N_22074,N_22366);
and U22960 (N_22960,N_22018,N_22335);
and U22961 (N_22961,N_22258,N_22499);
nand U22962 (N_22962,N_22471,N_22312);
and U22963 (N_22963,N_22151,N_22001);
and U22964 (N_22964,N_22162,N_22209);
xnor U22965 (N_22965,N_22457,N_22238);
xnor U22966 (N_22966,N_22364,N_22015);
and U22967 (N_22967,N_22382,N_22387);
nand U22968 (N_22968,N_22465,N_22488);
or U22969 (N_22969,N_22097,N_22148);
or U22970 (N_22970,N_22147,N_22184);
nor U22971 (N_22971,N_22233,N_22449);
and U22972 (N_22972,N_22260,N_22309);
xor U22973 (N_22973,N_22494,N_22058);
and U22974 (N_22974,N_22149,N_22411);
nand U22975 (N_22975,N_22226,N_22370);
xor U22976 (N_22976,N_22048,N_22155);
and U22977 (N_22977,N_22402,N_22015);
nor U22978 (N_22978,N_22354,N_22151);
xor U22979 (N_22979,N_22195,N_22304);
xnor U22980 (N_22980,N_22109,N_22286);
xnor U22981 (N_22981,N_22033,N_22078);
or U22982 (N_22982,N_22016,N_22161);
or U22983 (N_22983,N_22380,N_22117);
or U22984 (N_22984,N_22187,N_22307);
nand U22985 (N_22985,N_22040,N_22264);
and U22986 (N_22986,N_22362,N_22221);
xor U22987 (N_22987,N_22418,N_22333);
xnor U22988 (N_22988,N_22308,N_22230);
xor U22989 (N_22989,N_22250,N_22039);
xor U22990 (N_22990,N_22267,N_22213);
or U22991 (N_22991,N_22265,N_22331);
nand U22992 (N_22992,N_22114,N_22164);
or U22993 (N_22993,N_22092,N_22032);
xor U22994 (N_22994,N_22075,N_22205);
and U22995 (N_22995,N_22099,N_22324);
or U22996 (N_22996,N_22429,N_22079);
nand U22997 (N_22997,N_22148,N_22295);
or U22998 (N_22998,N_22010,N_22027);
or U22999 (N_22999,N_22148,N_22229);
and U23000 (N_23000,N_22591,N_22952);
or U23001 (N_23001,N_22698,N_22526);
xnor U23002 (N_23002,N_22899,N_22917);
nor U23003 (N_23003,N_22503,N_22836);
nor U23004 (N_23004,N_22864,N_22753);
and U23005 (N_23005,N_22657,N_22598);
xor U23006 (N_23006,N_22746,N_22908);
or U23007 (N_23007,N_22937,N_22841);
and U23008 (N_23008,N_22826,N_22688);
nor U23009 (N_23009,N_22985,N_22564);
and U23010 (N_23010,N_22946,N_22811);
xor U23011 (N_23011,N_22606,N_22837);
nand U23012 (N_23012,N_22786,N_22510);
nor U23013 (N_23013,N_22918,N_22911);
nor U23014 (N_23014,N_22672,N_22938);
or U23015 (N_23015,N_22709,N_22764);
nand U23016 (N_23016,N_22782,N_22724);
nand U23017 (N_23017,N_22798,N_22717);
nand U23018 (N_23018,N_22643,N_22880);
xnor U23019 (N_23019,N_22663,N_22758);
or U23020 (N_23020,N_22857,N_22973);
xnor U23021 (N_23021,N_22642,N_22860);
xnor U23022 (N_23022,N_22733,N_22781);
xnor U23023 (N_23023,N_22674,N_22518);
and U23024 (N_23024,N_22892,N_22677);
or U23025 (N_23025,N_22656,N_22673);
nand U23026 (N_23026,N_22921,N_22705);
nand U23027 (N_23027,N_22589,N_22844);
nor U23028 (N_23028,N_22902,N_22873);
or U23029 (N_23029,N_22605,N_22727);
xor U23030 (N_23030,N_22759,N_22633);
and U23031 (N_23031,N_22795,N_22628);
or U23032 (N_23032,N_22504,N_22616);
nor U23033 (N_23033,N_22517,N_22829);
nand U23034 (N_23034,N_22772,N_22687);
or U23035 (N_23035,N_22919,N_22925);
nor U23036 (N_23036,N_22914,N_22878);
and U23037 (N_23037,N_22960,N_22586);
xnor U23038 (N_23038,N_22726,N_22872);
or U23039 (N_23039,N_22942,N_22541);
nor U23040 (N_23040,N_22755,N_22824);
nor U23041 (N_23041,N_22689,N_22557);
and U23042 (N_23042,N_22777,N_22978);
nand U23043 (N_23043,N_22723,N_22654);
or U23044 (N_23044,N_22794,N_22940);
xor U23045 (N_23045,N_22515,N_22767);
xnor U23046 (N_23046,N_22729,N_22570);
nand U23047 (N_23047,N_22868,N_22757);
nand U23048 (N_23048,N_22981,N_22632);
or U23049 (N_23049,N_22585,N_22553);
nand U23050 (N_23050,N_22832,N_22820);
xnor U23051 (N_23051,N_22704,N_22538);
nand U23052 (N_23052,N_22732,N_22527);
xor U23053 (N_23053,N_22924,N_22810);
or U23054 (N_23054,N_22660,N_22690);
xor U23055 (N_23055,N_22506,N_22863);
and U23056 (N_23056,N_22613,N_22813);
nand U23057 (N_23057,N_22608,N_22650);
and U23058 (N_23058,N_22742,N_22520);
xnor U23059 (N_23059,N_22610,N_22659);
nand U23060 (N_23060,N_22516,N_22664);
or U23061 (N_23061,N_22971,N_22619);
nand U23062 (N_23062,N_22821,N_22966);
or U23063 (N_23063,N_22988,N_22554);
and U23064 (N_23064,N_22913,N_22947);
nor U23065 (N_23065,N_22686,N_22684);
and U23066 (N_23066,N_22648,N_22840);
and U23067 (N_23067,N_22768,N_22621);
nand U23068 (N_23068,N_22876,N_22900);
xor U23069 (N_23069,N_22696,N_22790);
xor U23070 (N_23070,N_22855,N_22627);
nor U23071 (N_23071,N_22850,N_22641);
nor U23072 (N_23072,N_22569,N_22852);
nor U23073 (N_23073,N_22734,N_22539);
and U23074 (N_23074,N_22970,N_22572);
nor U23075 (N_23075,N_22640,N_22653);
or U23076 (N_23076,N_22895,N_22760);
nor U23077 (N_23077,N_22675,N_22521);
nor U23078 (N_23078,N_22853,N_22883);
or U23079 (N_23079,N_22563,N_22962);
and U23080 (N_23080,N_22611,N_22901);
xor U23081 (N_23081,N_22828,N_22949);
and U23082 (N_23082,N_22814,N_22602);
nor U23083 (N_23083,N_22825,N_22915);
xnor U23084 (N_23084,N_22927,N_22576);
and U23085 (N_23085,N_22617,N_22730);
nor U23086 (N_23086,N_22514,N_22839);
or U23087 (N_23087,N_22969,N_22509);
and U23088 (N_23088,N_22630,N_22751);
and U23089 (N_23089,N_22972,N_22953);
xor U23090 (N_23090,N_22568,N_22754);
nand U23091 (N_23091,N_22738,N_22625);
and U23092 (N_23092,N_22920,N_22791);
xor U23093 (N_23093,N_22702,N_22594);
xor U23094 (N_23094,N_22649,N_22870);
xnor U23095 (N_23095,N_22776,N_22739);
nor U23096 (N_23096,N_22590,N_22596);
or U23097 (N_23097,N_22858,N_22647);
and U23098 (N_23098,N_22773,N_22834);
and U23099 (N_23099,N_22959,N_22551);
xor U23100 (N_23100,N_22979,N_22561);
and U23101 (N_23101,N_22999,N_22588);
nand U23102 (N_23102,N_22540,N_22546);
or U23103 (N_23103,N_22519,N_22685);
and U23104 (N_23104,N_22965,N_22620);
nand U23105 (N_23105,N_22667,N_22603);
xor U23106 (N_23106,N_22968,N_22866);
nor U23107 (N_23107,N_22885,N_22762);
xor U23108 (N_23108,N_22618,N_22725);
xor U23109 (N_23109,N_22804,N_22882);
xnor U23110 (N_23110,N_22793,N_22592);
nand U23111 (N_23111,N_22771,N_22827);
xor U23112 (N_23112,N_22678,N_22903);
or U23113 (N_23113,N_22671,N_22547);
and U23114 (N_23114,N_22565,N_22955);
nand U23115 (N_23115,N_22907,N_22713);
and U23116 (N_23116,N_22706,N_22898);
xnor U23117 (N_23117,N_22893,N_22976);
nor U23118 (N_23118,N_22577,N_22805);
nand U23119 (N_23119,N_22512,N_22812);
nor U23120 (N_23120,N_22566,N_22708);
or U23121 (N_23121,N_22692,N_22502);
nor U23122 (N_23122,N_22580,N_22635);
nand U23123 (N_23123,N_22575,N_22756);
nor U23124 (N_23124,N_22823,N_22644);
xnor U23125 (N_23125,N_22948,N_22770);
xor U23126 (N_23126,N_22500,N_22939);
xnor U23127 (N_23127,N_22682,N_22714);
or U23128 (N_23128,N_22865,N_22797);
nor U23129 (N_23129,N_22958,N_22549);
xor U23130 (N_23130,N_22763,N_22721);
xnor U23131 (N_23131,N_22928,N_22604);
or U23132 (N_23132,N_22703,N_22501);
or U23133 (N_23133,N_22909,N_22505);
xor U23134 (N_23134,N_22728,N_22681);
xor U23135 (N_23135,N_22508,N_22612);
nand U23136 (N_23136,N_22694,N_22548);
and U23137 (N_23137,N_22623,N_22996);
and U23138 (N_23138,N_22854,N_22974);
nand U23139 (N_23139,N_22740,N_22666);
nand U23140 (N_23140,N_22774,N_22951);
nand U23141 (N_23141,N_22887,N_22513);
xor U23142 (N_23142,N_22808,N_22997);
and U23143 (N_23143,N_22904,N_22993);
nor U23144 (N_23144,N_22990,N_22780);
nor U23145 (N_23145,N_22987,N_22769);
nor U23146 (N_23146,N_22761,N_22775);
or U23147 (N_23147,N_22809,N_22819);
xnor U23148 (N_23148,N_22542,N_22711);
nor U23149 (N_23149,N_22789,N_22545);
nor U23150 (N_23150,N_22982,N_22856);
and U23151 (N_23151,N_22579,N_22897);
nor U23152 (N_23152,N_22584,N_22802);
nand U23153 (N_23153,N_22567,N_22524);
nand U23154 (N_23154,N_22954,N_22595);
or U23155 (N_23155,N_22670,N_22910);
or U23156 (N_23156,N_22994,N_22783);
or U23157 (N_23157,N_22835,N_22923);
or U23158 (N_23158,N_22637,N_22930);
xnor U23159 (N_23159,N_22846,N_22535);
nand U23160 (N_23160,N_22735,N_22983);
nor U23161 (N_23161,N_22697,N_22523);
nand U23162 (N_23162,N_22583,N_22668);
nand U23163 (N_23163,N_22977,N_22749);
nor U23164 (N_23164,N_22693,N_22905);
nand U23165 (N_23165,N_22935,N_22862);
nand U23166 (N_23166,N_22533,N_22599);
xnor U23167 (N_23167,N_22933,N_22944);
nand U23168 (N_23168,N_22556,N_22741);
or U23169 (N_23169,N_22869,N_22587);
nand U23170 (N_23170,N_22701,N_22943);
and U23171 (N_23171,N_22552,N_22646);
nor U23172 (N_23172,N_22838,N_22867);
or U23173 (N_23173,N_22531,N_22799);
nor U23174 (N_23174,N_22787,N_22691);
or U23175 (N_23175,N_22629,N_22800);
and U23176 (N_23176,N_22831,N_22558);
nor U23177 (N_23177,N_22661,N_22597);
nand U23178 (N_23178,N_22712,N_22743);
or U23179 (N_23179,N_22879,N_22778);
or U23180 (N_23180,N_22984,N_22680);
xor U23181 (N_23181,N_22581,N_22747);
nor U23182 (N_23182,N_22766,N_22859);
and U23183 (N_23183,N_22655,N_22784);
xor U23184 (N_23184,N_22536,N_22932);
nor U23185 (N_23185,N_22716,N_22975);
or U23186 (N_23186,N_22529,N_22651);
xor U23187 (N_23187,N_22624,N_22639);
xor U23188 (N_23188,N_22731,N_22950);
or U23189 (N_23189,N_22736,N_22956);
nand U23190 (N_23190,N_22638,N_22998);
nand U23191 (N_23191,N_22607,N_22816);
nand U23192 (N_23192,N_22967,N_22522);
and U23193 (N_23193,N_22995,N_22582);
xor U23194 (N_23194,N_22645,N_22626);
xnor U23195 (N_23195,N_22964,N_22788);
nor U23196 (N_23196,N_22992,N_22622);
and U23197 (N_23197,N_22765,N_22719);
and U23198 (N_23198,N_22871,N_22722);
nor U23199 (N_23199,N_22600,N_22888);
xor U23200 (N_23200,N_22785,N_22843);
xnor U23201 (N_23201,N_22614,N_22571);
nand U23202 (N_23202,N_22941,N_22851);
or U23203 (N_23203,N_22573,N_22574);
nor U23204 (N_23204,N_22931,N_22822);
nor U23205 (N_23205,N_22662,N_22815);
nand U23206 (N_23206,N_22779,N_22896);
nor U23207 (N_23207,N_22679,N_22601);
nand U23208 (N_23208,N_22874,N_22926);
nor U23209 (N_23209,N_22525,N_22560);
nor U23210 (N_23210,N_22665,N_22683);
nand U23211 (N_23211,N_22912,N_22631);
or U23212 (N_23212,N_22796,N_22986);
or U23213 (N_23213,N_22916,N_22877);
and U23214 (N_23214,N_22894,N_22818);
nand U23215 (N_23215,N_22700,N_22745);
xor U23216 (N_23216,N_22980,N_22750);
and U23217 (N_23217,N_22669,N_22737);
nor U23218 (N_23218,N_22884,N_22578);
nor U23219 (N_23219,N_22890,N_22530);
nor U23220 (N_23220,N_22562,N_22652);
and U23221 (N_23221,N_22550,N_22861);
or U23222 (N_23222,N_22676,N_22936);
or U23223 (N_23223,N_22801,N_22989);
and U23224 (N_23224,N_22961,N_22830);
nand U23225 (N_23225,N_22991,N_22922);
and U23226 (N_23226,N_22636,N_22792);
xor U23227 (N_23227,N_22609,N_22833);
xnor U23228 (N_23228,N_22555,N_22845);
xnor U23229 (N_23229,N_22615,N_22534);
and U23230 (N_23230,N_22803,N_22710);
nor U23231 (N_23231,N_22543,N_22817);
nand U23232 (N_23232,N_22891,N_22695);
nand U23233 (N_23233,N_22889,N_22634);
or U23234 (N_23234,N_22507,N_22963);
nand U23235 (N_23235,N_22559,N_22906);
nand U23236 (N_23236,N_22886,N_22707);
and U23237 (N_23237,N_22847,N_22806);
or U23238 (N_23238,N_22532,N_22544);
or U23239 (N_23239,N_22699,N_22849);
or U23240 (N_23240,N_22528,N_22848);
nor U23241 (N_23241,N_22945,N_22718);
xor U23242 (N_23242,N_22744,N_22875);
or U23243 (N_23243,N_22537,N_22752);
or U23244 (N_23244,N_22511,N_22842);
nor U23245 (N_23245,N_22929,N_22720);
xor U23246 (N_23246,N_22881,N_22934);
or U23247 (N_23247,N_22658,N_22957);
and U23248 (N_23248,N_22593,N_22715);
and U23249 (N_23249,N_22807,N_22748);
nor U23250 (N_23250,N_22671,N_22641);
and U23251 (N_23251,N_22606,N_22588);
or U23252 (N_23252,N_22799,N_22970);
and U23253 (N_23253,N_22795,N_22836);
and U23254 (N_23254,N_22758,N_22970);
nor U23255 (N_23255,N_22850,N_22831);
or U23256 (N_23256,N_22879,N_22771);
or U23257 (N_23257,N_22651,N_22885);
and U23258 (N_23258,N_22656,N_22712);
and U23259 (N_23259,N_22741,N_22801);
nor U23260 (N_23260,N_22607,N_22757);
or U23261 (N_23261,N_22632,N_22658);
xnor U23262 (N_23262,N_22749,N_22898);
xor U23263 (N_23263,N_22558,N_22705);
nor U23264 (N_23264,N_22817,N_22841);
xor U23265 (N_23265,N_22865,N_22718);
xnor U23266 (N_23266,N_22579,N_22916);
xnor U23267 (N_23267,N_22531,N_22947);
xnor U23268 (N_23268,N_22710,N_22816);
nor U23269 (N_23269,N_22699,N_22835);
and U23270 (N_23270,N_22528,N_22792);
nor U23271 (N_23271,N_22892,N_22861);
and U23272 (N_23272,N_22928,N_22925);
or U23273 (N_23273,N_22556,N_22576);
or U23274 (N_23274,N_22811,N_22858);
or U23275 (N_23275,N_22714,N_22767);
nor U23276 (N_23276,N_22890,N_22702);
and U23277 (N_23277,N_22605,N_22958);
xor U23278 (N_23278,N_22916,N_22911);
and U23279 (N_23279,N_22936,N_22618);
or U23280 (N_23280,N_22546,N_22883);
and U23281 (N_23281,N_22549,N_22623);
xor U23282 (N_23282,N_22532,N_22789);
nand U23283 (N_23283,N_22956,N_22893);
and U23284 (N_23284,N_22573,N_22796);
nor U23285 (N_23285,N_22858,N_22805);
or U23286 (N_23286,N_22680,N_22837);
nand U23287 (N_23287,N_22622,N_22720);
nand U23288 (N_23288,N_22751,N_22927);
xnor U23289 (N_23289,N_22722,N_22979);
or U23290 (N_23290,N_22598,N_22837);
xor U23291 (N_23291,N_22896,N_22773);
and U23292 (N_23292,N_22940,N_22913);
or U23293 (N_23293,N_22633,N_22583);
and U23294 (N_23294,N_22769,N_22723);
nor U23295 (N_23295,N_22510,N_22645);
and U23296 (N_23296,N_22702,N_22969);
nor U23297 (N_23297,N_22970,N_22718);
xor U23298 (N_23298,N_22546,N_22500);
nor U23299 (N_23299,N_22812,N_22615);
nor U23300 (N_23300,N_22636,N_22863);
or U23301 (N_23301,N_22965,N_22700);
nor U23302 (N_23302,N_22649,N_22681);
nor U23303 (N_23303,N_22589,N_22594);
or U23304 (N_23304,N_22915,N_22820);
and U23305 (N_23305,N_22871,N_22857);
and U23306 (N_23306,N_22716,N_22837);
and U23307 (N_23307,N_22531,N_22542);
and U23308 (N_23308,N_22922,N_22683);
xnor U23309 (N_23309,N_22532,N_22793);
or U23310 (N_23310,N_22763,N_22626);
nand U23311 (N_23311,N_22607,N_22976);
and U23312 (N_23312,N_22532,N_22765);
nor U23313 (N_23313,N_22850,N_22695);
nand U23314 (N_23314,N_22583,N_22701);
and U23315 (N_23315,N_22620,N_22920);
and U23316 (N_23316,N_22631,N_22925);
or U23317 (N_23317,N_22692,N_22534);
xnor U23318 (N_23318,N_22994,N_22755);
and U23319 (N_23319,N_22921,N_22781);
or U23320 (N_23320,N_22976,N_22772);
xor U23321 (N_23321,N_22581,N_22955);
or U23322 (N_23322,N_22909,N_22674);
xnor U23323 (N_23323,N_22929,N_22971);
and U23324 (N_23324,N_22567,N_22844);
and U23325 (N_23325,N_22923,N_22749);
and U23326 (N_23326,N_22682,N_22672);
nor U23327 (N_23327,N_22604,N_22590);
nand U23328 (N_23328,N_22504,N_22969);
or U23329 (N_23329,N_22719,N_22588);
or U23330 (N_23330,N_22667,N_22997);
nor U23331 (N_23331,N_22678,N_22913);
nor U23332 (N_23332,N_22944,N_22655);
nor U23333 (N_23333,N_22553,N_22948);
xor U23334 (N_23334,N_22661,N_22890);
nand U23335 (N_23335,N_22639,N_22881);
or U23336 (N_23336,N_22816,N_22723);
nand U23337 (N_23337,N_22951,N_22957);
nand U23338 (N_23338,N_22714,N_22616);
nand U23339 (N_23339,N_22618,N_22908);
nor U23340 (N_23340,N_22980,N_22850);
nor U23341 (N_23341,N_22972,N_22561);
xor U23342 (N_23342,N_22819,N_22783);
nand U23343 (N_23343,N_22706,N_22609);
and U23344 (N_23344,N_22717,N_22771);
xnor U23345 (N_23345,N_22544,N_22969);
or U23346 (N_23346,N_22588,N_22697);
nor U23347 (N_23347,N_22833,N_22931);
nor U23348 (N_23348,N_22660,N_22546);
xor U23349 (N_23349,N_22802,N_22998);
nor U23350 (N_23350,N_22517,N_22708);
nor U23351 (N_23351,N_22511,N_22813);
and U23352 (N_23352,N_22785,N_22909);
and U23353 (N_23353,N_22850,N_22856);
nand U23354 (N_23354,N_22671,N_22840);
nand U23355 (N_23355,N_22596,N_22866);
or U23356 (N_23356,N_22664,N_22633);
and U23357 (N_23357,N_22782,N_22620);
nand U23358 (N_23358,N_22560,N_22955);
and U23359 (N_23359,N_22897,N_22626);
xnor U23360 (N_23360,N_22660,N_22963);
and U23361 (N_23361,N_22907,N_22845);
and U23362 (N_23362,N_22692,N_22568);
nand U23363 (N_23363,N_22862,N_22954);
or U23364 (N_23364,N_22841,N_22806);
xnor U23365 (N_23365,N_22729,N_22703);
xnor U23366 (N_23366,N_22585,N_22944);
nor U23367 (N_23367,N_22584,N_22936);
or U23368 (N_23368,N_22599,N_22725);
xnor U23369 (N_23369,N_22684,N_22943);
and U23370 (N_23370,N_22550,N_22687);
xnor U23371 (N_23371,N_22940,N_22861);
nor U23372 (N_23372,N_22891,N_22502);
nand U23373 (N_23373,N_22875,N_22719);
or U23374 (N_23374,N_22706,N_22552);
xor U23375 (N_23375,N_22758,N_22971);
or U23376 (N_23376,N_22589,N_22906);
or U23377 (N_23377,N_22517,N_22971);
or U23378 (N_23378,N_22674,N_22948);
or U23379 (N_23379,N_22893,N_22667);
nor U23380 (N_23380,N_22917,N_22768);
nor U23381 (N_23381,N_22958,N_22529);
xnor U23382 (N_23382,N_22633,N_22778);
or U23383 (N_23383,N_22919,N_22861);
nand U23384 (N_23384,N_22644,N_22515);
and U23385 (N_23385,N_22855,N_22570);
or U23386 (N_23386,N_22941,N_22674);
xnor U23387 (N_23387,N_22614,N_22911);
and U23388 (N_23388,N_22722,N_22703);
nor U23389 (N_23389,N_22596,N_22715);
nor U23390 (N_23390,N_22757,N_22829);
xnor U23391 (N_23391,N_22662,N_22598);
and U23392 (N_23392,N_22569,N_22823);
nand U23393 (N_23393,N_22537,N_22576);
or U23394 (N_23394,N_22861,N_22634);
nor U23395 (N_23395,N_22525,N_22558);
and U23396 (N_23396,N_22870,N_22608);
and U23397 (N_23397,N_22517,N_22751);
nor U23398 (N_23398,N_22919,N_22621);
nor U23399 (N_23399,N_22682,N_22546);
nor U23400 (N_23400,N_22883,N_22862);
or U23401 (N_23401,N_22596,N_22687);
nor U23402 (N_23402,N_22757,N_22748);
nand U23403 (N_23403,N_22976,N_22915);
xnor U23404 (N_23404,N_22991,N_22726);
or U23405 (N_23405,N_22650,N_22603);
nor U23406 (N_23406,N_22644,N_22939);
or U23407 (N_23407,N_22983,N_22558);
nand U23408 (N_23408,N_22808,N_22769);
xor U23409 (N_23409,N_22746,N_22593);
xor U23410 (N_23410,N_22949,N_22521);
xnor U23411 (N_23411,N_22669,N_22821);
nand U23412 (N_23412,N_22806,N_22660);
or U23413 (N_23413,N_22656,N_22911);
xor U23414 (N_23414,N_22779,N_22725);
xnor U23415 (N_23415,N_22891,N_22869);
nor U23416 (N_23416,N_22747,N_22927);
nor U23417 (N_23417,N_22813,N_22915);
nor U23418 (N_23418,N_22913,N_22723);
xnor U23419 (N_23419,N_22728,N_22692);
and U23420 (N_23420,N_22779,N_22535);
or U23421 (N_23421,N_22717,N_22897);
nand U23422 (N_23422,N_22548,N_22946);
or U23423 (N_23423,N_22600,N_22784);
nor U23424 (N_23424,N_22623,N_22692);
or U23425 (N_23425,N_22698,N_22512);
nor U23426 (N_23426,N_22868,N_22632);
nor U23427 (N_23427,N_22959,N_22967);
xor U23428 (N_23428,N_22918,N_22736);
nand U23429 (N_23429,N_22768,N_22859);
nor U23430 (N_23430,N_22883,N_22742);
or U23431 (N_23431,N_22654,N_22756);
nor U23432 (N_23432,N_22698,N_22565);
xor U23433 (N_23433,N_22812,N_22670);
and U23434 (N_23434,N_22915,N_22749);
xor U23435 (N_23435,N_22890,N_22536);
xnor U23436 (N_23436,N_22564,N_22861);
nand U23437 (N_23437,N_22566,N_22647);
nor U23438 (N_23438,N_22891,N_22613);
or U23439 (N_23439,N_22698,N_22929);
xor U23440 (N_23440,N_22674,N_22646);
or U23441 (N_23441,N_22810,N_22580);
xor U23442 (N_23442,N_22572,N_22997);
or U23443 (N_23443,N_22744,N_22977);
and U23444 (N_23444,N_22838,N_22786);
nor U23445 (N_23445,N_22638,N_22641);
nor U23446 (N_23446,N_22927,N_22874);
xnor U23447 (N_23447,N_22703,N_22857);
or U23448 (N_23448,N_22729,N_22585);
and U23449 (N_23449,N_22979,N_22541);
or U23450 (N_23450,N_22691,N_22515);
nor U23451 (N_23451,N_22872,N_22582);
or U23452 (N_23452,N_22953,N_22649);
or U23453 (N_23453,N_22792,N_22937);
xnor U23454 (N_23454,N_22805,N_22589);
nor U23455 (N_23455,N_22907,N_22865);
and U23456 (N_23456,N_22584,N_22812);
or U23457 (N_23457,N_22511,N_22841);
or U23458 (N_23458,N_22734,N_22861);
nor U23459 (N_23459,N_22763,N_22526);
and U23460 (N_23460,N_22532,N_22762);
and U23461 (N_23461,N_22719,N_22526);
nand U23462 (N_23462,N_22963,N_22590);
xnor U23463 (N_23463,N_22564,N_22682);
or U23464 (N_23464,N_22570,N_22586);
or U23465 (N_23465,N_22784,N_22910);
nor U23466 (N_23466,N_22710,N_22831);
nand U23467 (N_23467,N_22508,N_22808);
or U23468 (N_23468,N_22649,N_22666);
nand U23469 (N_23469,N_22637,N_22724);
or U23470 (N_23470,N_22977,N_22584);
xor U23471 (N_23471,N_22573,N_22657);
nor U23472 (N_23472,N_22630,N_22993);
and U23473 (N_23473,N_22528,N_22935);
and U23474 (N_23474,N_22988,N_22634);
nor U23475 (N_23475,N_22713,N_22892);
and U23476 (N_23476,N_22962,N_22761);
and U23477 (N_23477,N_22530,N_22901);
xor U23478 (N_23478,N_22908,N_22763);
nor U23479 (N_23479,N_22744,N_22832);
and U23480 (N_23480,N_22723,N_22852);
and U23481 (N_23481,N_22839,N_22699);
nand U23482 (N_23482,N_22881,N_22930);
nand U23483 (N_23483,N_22959,N_22994);
xnor U23484 (N_23484,N_22954,N_22833);
and U23485 (N_23485,N_22636,N_22997);
or U23486 (N_23486,N_22985,N_22951);
nor U23487 (N_23487,N_22876,N_22668);
nor U23488 (N_23488,N_22803,N_22744);
and U23489 (N_23489,N_22534,N_22532);
nor U23490 (N_23490,N_22864,N_22877);
nand U23491 (N_23491,N_22508,N_22754);
or U23492 (N_23492,N_22951,N_22791);
or U23493 (N_23493,N_22984,N_22891);
xor U23494 (N_23494,N_22991,N_22815);
nand U23495 (N_23495,N_22661,N_22861);
xor U23496 (N_23496,N_22947,N_22868);
or U23497 (N_23497,N_22933,N_22755);
nor U23498 (N_23498,N_22549,N_22901);
nor U23499 (N_23499,N_22798,N_22904);
nand U23500 (N_23500,N_23430,N_23249);
nand U23501 (N_23501,N_23149,N_23028);
or U23502 (N_23502,N_23373,N_23263);
and U23503 (N_23503,N_23122,N_23157);
or U23504 (N_23504,N_23154,N_23477);
or U23505 (N_23505,N_23248,N_23493);
and U23506 (N_23506,N_23050,N_23343);
nor U23507 (N_23507,N_23364,N_23062);
or U23508 (N_23508,N_23135,N_23034);
nand U23509 (N_23509,N_23499,N_23195);
xor U23510 (N_23510,N_23369,N_23346);
and U23511 (N_23511,N_23087,N_23338);
nor U23512 (N_23512,N_23146,N_23102);
xnor U23513 (N_23513,N_23459,N_23478);
and U23514 (N_23514,N_23242,N_23189);
xnor U23515 (N_23515,N_23185,N_23236);
nand U23516 (N_23516,N_23496,N_23255);
xor U23517 (N_23517,N_23440,N_23424);
or U23518 (N_23518,N_23183,N_23417);
xor U23519 (N_23519,N_23309,N_23112);
nand U23520 (N_23520,N_23426,N_23040);
nor U23521 (N_23521,N_23386,N_23179);
xnor U23522 (N_23522,N_23095,N_23490);
or U23523 (N_23523,N_23344,N_23193);
nand U23524 (N_23524,N_23103,N_23350);
and U23525 (N_23525,N_23181,N_23258);
nor U23526 (N_23526,N_23170,N_23205);
nor U23527 (N_23527,N_23360,N_23412);
and U23528 (N_23528,N_23024,N_23140);
or U23529 (N_23529,N_23152,N_23158);
or U23530 (N_23530,N_23167,N_23042);
and U23531 (N_23531,N_23268,N_23199);
nor U23532 (N_23532,N_23401,N_23053);
and U23533 (N_23533,N_23056,N_23172);
and U23534 (N_23534,N_23296,N_23041);
and U23535 (N_23535,N_23367,N_23267);
nand U23536 (N_23536,N_23194,N_23022);
or U23537 (N_23537,N_23332,N_23191);
or U23538 (N_23538,N_23409,N_23282);
or U23539 (N_23539,N_23120,N_23388);
or U23540 (N_23540,N_23304,N_23432);
and U23541 (N_23541,N_23488,N_23302);
or U23542 (N_23542,N_23331,N_23037);
xnor U23543 (N_23543,N_23380,N_23245);
nand U23544 (N_23544,N_23252,N_23210);
nor U23545 (N_23545,N_23074,N_23368);
nand U23546 (N_23546,N_23222,N_23330);
or U23547 (N_23547,N_23136,N_23025);
nor U23548 (N_23548,N_23353,N_23305);
xor U23549 (N_23549,N_23144,N_23241);
nor U23550 (N_23550,N_23235,N_23107);
nand U23551 (N_23551,N_23009,N_23212);
or U23552 (N_23552,N_23481,N_23049);
or U23553 (N_23553,N_23473,N_23291);
nor U23554 (N_23554,N_23370,N_23137);
or U23555 (N_23555,N_23035,N_23202);
xor U23556 (N_23556,N_23200,N_23403);
nand U23557 (N_23557,N_23465,N_23308);
nand U23558 (N_23558,N_23196,N_23339);
xnor U23559 (N_23559,N_23247,N_23182);
and U23560 (N_23560,N_23351,N_23164);
nor U23561 (N_23561,N_23471,N_23410);
nor U23562 (N_23562,N_23358,N_23067);
nor U23563 (N_23563,N_23010,N_23390);
nor U23564 (N_23564,N_23138,N_23127);
and U23565 (N_23565,N_23150,N_23059);
nor U23566 (N_23566,N_23392,N_23450);
nor U23567 (N_23567,N_23257,N_23318);
nor U23568 (N_23568,N_23008,N_23007);
nand U23569 (N_23569,N_23280,N_23111);
xnor U23570 (N_23570,N_23303,N_23231);
nand U23571 (N_23571,N_23246,N_23314);
nand U23572 (N_23572,N_23307,N_23029);
and U23573 (N_23573,N_23153,N_23229);
nor U23574 (N_23574,N_23123,N_23480);
xnor U23575 (N_23575,N_23352,N_23214);
xnor U23576 (N_23576,N_23470,N_23461);
nand U23577 (N_23577,N_23209,N_23463);
nor U23578 (N_23578,N_23130,N_23462);
or U23579 (N_23579,N_23436,N_23016);
xor U23580 (N_23580,N_23383,N_23043);
nand U23581 (N_23581,N_23211,N_23064);
nor U23582 (N_23582,N_23115,N_23237);
nor U23583 (N_23583,N_23047,N_23306);
and U23584 (N_23584,N_23491,N_23418);
and U23585 (N_23585,N_23293,N_23001);
or U23586 (N_23586,N_23228,N_23190);
xor U23587 (N_23587,N_23097,N_23279);
nand U23588 (N_23588,N_23243,N_23080);
nor U23589 (N_23589,N_23166,N_23327);
nand U23590 (N_23590,N_23299,N_23260);
nor U23591 (N_23591,N_23208,N_23396);
nand U23592 (N_23592,N_23232,N_23437);
xor U23593 (N_23593,N_23377,N_23084);
or U23594 (N_23594,N_23495,N_23227);
and U23595 (N_23595,N_23326,N_23472);
and U23596 (N_23596,N_23448,N_23278);
nor U23597 (N_23597,N_23175,N_23233);
xor U23598 (N_23598,N_23316,N_23163);
and U23599 (N_23599,N_23474,N_23482);
or U23600 (N_23600,N_23375,N_23178);
xnor U23601 (N_23601,N_23186,N_23323);
nor U23602 (N_23602,N_23265,N_23328);
or U23603 (N_23603,N_23230,N_23468);
nor U23604 (N_23604,N_23438,N_23169);
nand U23605 (N_23605,N_23366,N_23203);
xnor U23606 (N_23606,N_23239,N_23384);
nand U23607 (N_23607,N_23286,N_23421);
or U23608 (N_23608,N_23483,N_23301);
nor U23609 (N_23609,N_23151,N_23272);
or U23610 (N_23610,N_23479,N_23070);
nand U23611 (N_23611,N_23441,N_23033);
nand U23612 (N_23612,N_23294,N_23487);
or U23613 (N_23613,N_23273,N_23439);
and U23614 (N_23614,N_23031,N_23073);
nor U23615 (N_23615,N_23363,N_23069);
and U23616 (N_23616,N_23192,N_23362);
or U23617 (N_23617,N_23443,N_23391);
and U23618 (N_23618,N_23124,N_23032);
or U23619 (N_23619,N_23093,N_23334);
nor U23620 (N_23620,N_23134,N_23374);
or U23621 (N_23621,N_23141,N_23213);
nand U23622 (N_23622,N_23177,N_23006);
nand U23623 (N_23623,N_23425,N_23125);
xnor U23624 (N_23624,N_23184,N_23337);
or U23625 (N_23625,N_23261,N_23058);
or U23626 (N_23626,N_23288,N_23311);
nand U23627 (N_23627,N_23420,N_23066);
or U23628 (N_23628,N_23054,N_23398);
nand U23629 (N_23629,N_23250,N_23456);
nand U23630 (N_23630,N_23096,N_23492);
xor U23631 (N_23631,N_23206,N_23297);
xnor U23632 (N_23632,N_23086,N_23004);
nand U23633 (N_23633,N_23027,N_23379);
and U23634 (N_23634,N_23416,N_23313);
xnor U23635 (N_23635,N_23218,N_23023);
nor U23636 (N_23636,N_23197,N_23395);
or U23637 (N_23637,N_23110,N_23251);
or U23638 (N_23638,N_23065,N_23238);
and U23639 (N_23639,N_23108,N_23295);
xor U23640 (N_23640,N_23335,N_23497);
or U23641 (N_23641,N_23460,N_23106);
or U23642 (N_23642,N_23216,N_23381);
xnor U23643 (N_23643,N_23148,N_23240);
or U23644 (N_23644,N_23378,N_23394);
and U23645 (N_23645,N_23142,N_23429);
nand U23646 (N_23646,N_23341,N_23442);
and U23647 (N_23647,N_23092,N_23259);
or U23648 (N_23648,N_23319,N_23133);
nand U23649 (N_23649,N_23117,N_23168);
and U23650 (N_23650,N_23419,N_23101);
xor U23651 (N_23651,N_23405,N_23081);
nor U23652 (N_23652,N_23285,N_23089);
and U23653 (N_23653,N_23264,N_23310);
or U23654 (N_23654,N_23464,N_23447);
or U23655 (N_23655,N_23382,N_23005);
and U23656 (N_23656,N_23345,N_23026);
or U23657 (N_23657,N_23290,N_23276);
and U23658 (N_23658,N_23423,N_23165);
nand U23659 (N_23659,N_23322,N_23173);
or U23660 (N_23660,N_23090,N_23176);
or U23661 (N_23661,N_23467,N_23044);
nor U23662 (N_23662,N_23454,N_23253);
nand U23663 (N_23663,N_23348,N_23099);
xnor U23664 (N_23664,N_23171,N_23275);
nand U23665 (N_23665,N_23393,N_23466);
or U23666 (N_23666,N_23220,N_23427);
xnor U23667 (N_23667,N_23281,N_23453);
xor U23668 (N_23668,N_23078,N_23098);
xor U23669 (N_23669,N_23128,N_23320);
xnor U23670 (N_23670,N_23160,N_23215);
and U23671 (N_23671,N_23428,N_23372);
nor U23672 (N_23672,N_23071,N_23019);
nand U23673 (N_23673,N_23361,N_23063);
xnor U23674 (N_23674,N_23365,N_23055);
nand U23675 (N_23675,N_23011,N_23036);
nand U23676 (N_23676,N_23399,N_23254);
nand U23677 (N_23677,N_23486,N_23413);
nor U23678 (N_23678,N_23020,N_23325);
and U23679 (N_23679,N_23408,N_23289);
nand U23680 (N_23680,N_23476,N_23109);
or U23681 (N_23681,N_23445,N_23444);
nand U23682 (N_23682,N_23003,N_23126);
and U23683 (N_23683,N_23132,N_23030);
nand U23684 (N_23684,N_23226,N_23449);
xnor U23685 (N_23685,N_23376,N_23162);
nand U23686 (N_23686,N_23347,N_23406);
and U23687 (N_23687,N_23431,N_23079);
nand U23688 (N_23688,N_23129,N_23455);
nor U23689 (N_23689,N_23155,N_23002);
or U23690 (N_23690,N_23411,N_23298);
or U23691 (N_23691,N_23052,N_23113);
nor U23692 (N_23692,N_23244,N_23000);
nor U23693 (N_23693,N_23397,N_23224);
or U23694 (N_23694,N_23085,N_23180);
xnor U23695 (N_23695,N_23434,N_23475);
xor U23696 (N_23696,N_23270,N_23038);
and U23697 (N_23697,N_23105,N_23371);
nand U23698 (N_23698,N_23271,N_23159);
or U23699 (N_23699,N_23094,N_23415);
nand U23700 (N_23700,N_23225,N_23355);
nand U23701 (N_23701,N_23156,N_23342);
xor U23702 (N_23702,N_23404,N_23458);
nand U23703 (N_23703,N_23389,N_23435);
and U23704 (N_23704,N_23207,N_23048);
and U23705 (N_23705,N_23329,N_23407);
and U23706 (N_23706,N_23015,N_23201);
and U23707 (N_23707,N_23118,N_23217);
nand U23708 (N_23708,N_23221,N_23300);
nor U23709 (N_23709,N_23324,N_23385);
or U23710 (N_23710,N_23072,N_23457);
or U23711 (N_23711,N_23114,N_23356);
or U23712 (N_23712,N_23139,N_23400);
nor U23713 (N_23713,N_23121,N_23187);
or U23714 (N_23714,N_23104,N_23317);
or U23715 (N_23715,N_23336,N_23269);
and U23716 (N_23716,N_23489,N_23340);
xnor U23717 (N_23717,N_23451,N_23387);
and U23718 (N_23718,N_23131,N_23077);
nand U23719 (N_23719,N_23161,N_23145);
or U23720 (N_23720,N_23469,N_23083);
xnor U23721 (N_23721,N_23147,N_23452);
xor U23722 (N_23722,N_23060,N_23292);
nor U23723 (N_23723,N_23357,N_23116);
or U23724 (N_23724,N_23312,N_23076);
nor U23725 (N_23725,N_23446,N_23349);
or U23726 (N_23726,N_23354,N_23422);
or U23727 (N_23727,N_23321,N_23198);
and U23728 (N_23728,N_23219,N_23283);
or U23729 (N_23729,N_23277,N_23287);
xnor U23730 (N_23730,N_23274,N_23262);
and U23731 (N_23731,N_23014,N_23333);
or U23732 (N_23732,N_23256,N_23484);
xor U23733 (N_23733,N_23045,N_23039);
nand U23734 (N_23734,N_23012,N_23119);
nand U23735 (N_23735,N_23498,N_23091);
and U23736 (N_23736,N_23013,N_23204);
and U23737 (N_23737,N_23068,N_23433);
xnor U23738 (N_23738,N_23266,N_23174);
nand U23739 (N_23739,N_23082,N_23057);
or U23740 (N_23740,N_23234,N_23018);
xor U23741 (N_23741,N_23143,N_23051);
nand U23742 (N_23742,N_23315,N_23075);
xnor U23743 (N_23743,N_23061,N_23223);
xnor U23744 (N_23744,N_23402,N_23188);
or U23745 (N_23745,N_23414,N_23284);
xor U23746 (N_23746,N_23100,N_23359);
nand U23747 (N_23747,N_23485,N_23088);
xor U23748 (N_23748,N_23017,N_23046);
nand U23749 (N_23749,N_23494,N_23021);
xnor U23750 (N_23750,N_23480,N_23462);
or U23751 (N_23751,N_23193,N_23148);
and U23752 (N_23752,N_23071,N_23480);
nand U23753 (N_23753,N_23238,N_23223);
nor U23754 (N_23754,N_23404,N_23343);
and U23755 (N_23755,N_23047,N_23271);
nor U23756 (N_23756,N_23000,N_23449);
nor U23757 (N_23757,N_23180,N_23220);
xnor U23758 (N_23758,N_23129,N_23317);
nor U23759 (N_23759,N_23452,N_23287);
nand U23760 (N_23760,N_23154,N_23049);
or U23761 (N_23761,N_23354,N_23460);
xnor U23762 (N_23762,N_23106,N_23124);
nor U23763 (N_23763,N_23134,N_23226);
xnor U23764 (N_23764,N_23156,N_23363);
nor U23765 (N_23765,N_23281,N_23320);
xnor U23766 (N_23766,N_23056,N_23424);
xnor U23767 (N_23767,N_23383,N_23483);
xnor U23768 (N_23768,N_23338,N_23107);
xnor U23769 (N_23769,N_23384,N_23021);
or U23770 (N_23770,N_23291,N_23368);
and U23771 (N_23771,N_23238,N_23452);
nand U23772 (N_23772,N_23113,N_23018);
nor U23773 (N_23773,N_23415,N_23104);
and U23774 (N_23774,N_23341,N_23287);
xor U23775 (N_23775,N_23054,N_23324);
xnor U23776 (N_23776,N_23446,N_23016);
and U23777 (N_23777,N_23130,N_23461);
and U23778 (N_23778,N_23314,N_23363);
and U23779 (N_23779,N_23422,N_23032);
nor U23780 (N_23780,N_23223,N_23196);
xnor U23781 (N_23781,N_23213,N_23043);
nor U23782 (N_23782,N_23282,N_23477);
nor U23783 (N_23783,N_23127,N_23080);
nor U23784 (N_23784,N_23411,N_23409);
xor U23785 (N_23785,N_23133,N_23175);
or U23786 (N_23786,N_23259,N_23192);
nand U23787 (N_23787,N_23051,N_23206);
nor U23788 (N_23788,N_23187,N_23137);
or U23789 (N_23789,N_23407,N_23145);
xnor U23790 (N_23790,N_23131,N_23135);
nor U23791 (N_23791,N_23143,N_23028);
or U23792 (N_23792,N_23392,N_23240);
and U23793 (N_23793,N_23046,N_23296);
nor U23794 (N_23794,N_23472,N_23061);
xnor U23795 (N_23795,N_23454,N_23331);
and U23796 (N_23796,N_23280,N_23254);
xnor U23797 (N_23797,N_23320,N_23296);
or U23798 (N_23798,N_23010,N_23017);
and U23799 (N_23799,N_23404,N_23214);
and U23800 (N_23800,N_23375,N_23167);
or U23801 (N_23801,N_23126,N_23109);
nand U23802 (N_23802,N_23425,N_23135);
nor U23803 (N_23803,N_23069,N_23054);
nand U23804 (N_23804,N_23303,N_23326);
xnor U23805 (N_23805,N_23450,N_23321);
and U23806 (N_23806,N_23423,N_23371);
and U23807 (N_23807,N_23003,N_23477);
xnor U23808 (N_23808,N_23078,N_23300);
xor U23809 (N_23809,N_23245,N_23329);
and U23810 (N_23810,N_23442,N_23488);
or U23811 (N_23811,N_23479,N_23172);
nor U23812 (N_23812,N_23172,N_23168);
nor U23813 (N_23813,N_23214,N_23485);
or U23814 (N_23814,N_23016,N_23115);
or U23815 (N_23815,N_23083,N_23153);
nand U23816 (N_23816,N_23305,N_23004);
or U23817 (N_23817,N_23428,N_23371);
xnor U23818 (N_23818,N_23245,N_23056);
and U23819 (N_23819,N_23213,N_23242);
or U23820 (N_23820,N_23186,N_23464);
and U23821 (N_23821,N_23268,N_23349);
xnor U23822 (N_23822,N_23405,N_23479);
or U23823 (N_23823,N_23171,N_23492);
nor U23824 (N_23824,N_23102,N_23144);
nor U23825 (N_23825,N_23369,N_23110);
nor U23826 (N_23826,N_23313,N_23187);
nor U23827 (N_23827,N_23289,N_23456);
or U23828 (N_23828,N_23240,N_23471);
xnor U23829 (N_23829,N_23474,N_23260);
nand U23830 (N_23830,N_23341,N_23060);
or U23831 (N_23831,N_23418,N_23373);
xor U23832 (N_23832,N_23233,N_23055);
xor U23833 (N_23833,N_23289,N_23190);
nand U23834 (N_23834,N_23143,N_23429);
or U23835 (N_23835,N_23474,N_23173);
and U23836 (N_23836,N_23100,N_23300);
nor U23837 (N_23837,N_23329,N_23185);
or U23838 (N_23838,N_23022,N_23347);
or U23839 (N_23839,N_23026,N_23226);
and U23840 (N_23840,N_23151,N_23442);
xnor U23841 (N_23841,N_23423,N_23381);
nand U23842 (N_23842,N_23073,N_23481);
xnor U23843 (N_23843,N_23275,N_23472);
xnor U23844 (N_23844,N_23227,N_23458);
nand U23845 (N_23845,N_23349,N_23391);
or U23846 (N_23846,N_23483,N_23423);
nand U23847 (N_23847,N_23426,N_23176);
nor U23848 (N_23848,N_23214,N_23296);
nand U23849 (N_23849,N_23033,N_23056);
and U23850 (N_23850,N_23308,N_23162);
nand U23851 (N_23851,N_23216,N_23103);
or U23852 (N_23852,N_23445,N_23462);
nor U23853 (N_23853,N_23088,N_23151);
or U23854 (N_23854,N_23314,N_23431);
or U23855 (N_23855,N_23132,N_23190);
nand U23856 (N_23856,N_23011,N_23325);
nor U23857 (N_23857,N_23236,N_23336);
nand U23858 (N_23858,N_23152,N_23004);
xor U23859 (N_23859,N_23051,N_23261);
xnor U23860 (N_23860,N_23365,N_23334);
xnor U23861 (N_23861,N_23413,N_23435);
xnor U23862 (N_23862,N_23049,N_23020);
nand U23863 (N_23863,N_23119,N_23406);
and U23864 (N_23864,N_23476,N_23087);
or U23865 (N_23865,N_23353,N_23040);
xnor U23866 (N_23866,N_23316,N_23283);
nor U23867 (N_23867,N_23056,N_23423);
xnor U23868 (N_23868,N_23110,N_23114);
nand U23869 (N_23869,N_23121,N_23197);
or U23870 (N_23870,N_23181,N_23082);
nor U23871 (N_23871,N_23232,N_23416);
nand U23872 (N_23872,N_23123,N_23439);
and U23873 (N_23873,N_23381,N_23087);
xnor U23874 (N_23874,N_23408,N_23039);
and U23875 (N_23875,N_23432,N_23175);
nand U23876 (N_23876,N_23102,N_23352);
nand U23877 (N_23877,N_23486,N_23159);
nor U23878 (N_23878,N_23481,N_23227);
and U23879 (N_23879,N_23291,N_23084);
nor U23880 (N_23880,N_23129,N_23251);
nand U23881 (N_23881,N_23097,N_23017);
nor U23882 (N_23882,N_23007,N_23268);
xnor U23883 (N_23883,N_23088,N_23313);
or U23884 (N_23884,N_23211,N_23306);
nor U23885 (N_23885,N_23068,N_23150);
nor U23886 (N_23886,N_23270,N_23437);
nor U23887 (N_23887,N_23441,N_23204);
or U23888 (N_23888,N_23499,N_23455);
nand U23889 (N_23889,N_23023,N_23012);
nor U23890 (N_23890,N_23085,N_23342);
xor U23891 (N_23891,N_23491,N_23213);
or U23892 (N_23892,N_23139,N_23348);
nand U23893 (N_23893,N_23376,N_23451);
nand U23894 (N_23894,N_23471,N_23124);
nand U23895 (N_23895,N_23212,N_23483);
nor U23896 (N_23896,N_23374,N_23066);
nor U23897 (N_23897,N_23031,N_23344);
and U23898 (N_23898,N_23323,N_23264);
and U23899 (N_23899,N_23002,N_23394);
and U23900 (N_23900,N_23359,N_23477);
nand U23901 (N_23901,N_23363,N_23407);
nand U23902 (N_23902,N_23358,N_23379);
and U23903 (N_23903,N_23487,N_23000);
nor U23904 (N_23904,N_23023,N_23429);
and U23905 (N_23905,N_23034,N_23249);
or U23906 (N_23906,N_23359,N_23488);
or U23907 (N_23907,N_23162,N_23433);
nand U23908 (N_23908,N_23063,N_23295);
or U23909 (N_23909,N_23170,N_23180);
and U23910 (N_23910,N_23324,N_23486);
nand U23911 (N_23911,N_23037,N_23334);
and U23912 (N_23912,N_23318,N_23192);
xnor U23913 (N_23913,N_23352,N_23407);
nor U23914 (N_23914,N_23073,N_23122);
or U23915 (N_23915,N_23256,N_23081);
and U23916 (N_23916,N_23311,N_23032);
and U23917 (N_23917,N_23262,N_23225);
xnor U23918 (N_23918,N_23255,N_23314);
nand U23919 (N_23919,N_23400,N_23234);
nand U23920 (N_23920,N_23032,N_23158);
xor U23921 (N_23921,N_23183,N_23102);
or U23922 (N_23922,N_23232,N_23410);
nor U23923 (N_23923,N_23232,N_23438);
or U23924 (N_23924,N_23343,N_23163);
nand U23925 (N_23925,N_23023,N_23482);
nor U23926 (N_23926,N_23178,N_23457);
nand U23927 (N_23927,N_23423,N_23387);
nand U23928 (N_23928,N_23467,N_23491);
xor U23929 (N_23929,N_23221,N_23195);
nand U23930 (N_23930,N_23446,N_23199);
and U23931 (N_23931,N_23452,N_23023);
nor U23932 (N_23932,N_23396,N_23210);
nor U23933 (N_23933,N_23385,N_23152);
and U23934 (N_23934,N_23394,N_23190);
or U23935 (N_23935,N_23223,N_23052);
nor U23936 (N_23936,N_23060,N_23330);
nor U23937 (N_23937,N_23153,N_23432);
xor U23938 (N_23938,N_23401,N_23216);
xnor U23939 (N_23939,N_23209,N_23061);
nand U23940 (N_23940,N_23271,N_23473);
nand U23941 (N_23941,N_23199,N_23065);
or U23942 (N_23942,N_23430,N_23422);
nor U23943 (N_23943,N_23121,N_23327);
and U23944 (N_23944,N_23309,N_23487);
nor U23945 (N_23945,N_23332,N_23022);
nor U23946 (N_23946,N_23165,N_23485);
xor U23947 (N_23947,N_23268,N_23232);
nor U23948 (N_23948,N_23149,N_23005);
nor U23949 (N_23949,N_23468,N_23421);
nand U23950 (N_23950,N_23198,N_23257);
nand U23951 (N_23951,N_23037,N_23433);
and U23952 (N_23952,N_23204,N_23489);
nor U23953 (N_23953,N_23097,N_23026);
or U23954 (N_23954,N_23132,N_23169);
and U23955 (N_23955,N_23129,N_23163);
nor U23956 (N_23956,N_23484,N_23262);
nor U23957 (N_23957,N_23280,N_23377);
and U23958 (N_23958,N_23103,N_23136);
nor U23959 (N_23959,N_23021,N_23123);
and U23960 (N_23960,N_23269,N_23113);
xnor U23961 (N_23961,N_23115,N_23132);
or U23962 (N_23962,N_23445,N_23077);
and U23963 (N_23963,N_23186,N_23056);
nand U23964 (N_23964,N_23429,N_23438);
and U23965 (N_23965,N_23436,N_23026);
nor U23966 (N_23966,N_23168,N_23002);
nor U23967 (N_23967,N_23399,N_23014);
and U23968 (N_23968,N_23329,N_23018);
nand U23969 (N_23969,N_23496,N_23442);
nand U23970 (N_23970,N_23476,N_23092);
xor U23971 (N_23971,N_23208,N_23483);
nand U23972 (N_23972,N_23360,N_23391);
or U23973 (N_23973,N_23474,N_23211);
xor U23974 (N_23974,N_23127,N_23269);
nand U23975 (N_23975,N_23158,N_23236);
and U23976 (N_23976,N_23208,N_23273);
xor U23977 (N_23977,N_23094,N_23159);
and U23978 (N_23978,N_23220,N_23431);
or U23979 (N_23979,N_23063,N_23226);
xor U23980 (N_23980,N_23128,N_23258);
xnor U23981 (N_23981,N_23335,N_23212);
nand U23982 (N_23982,N_23258,N_23247);
or U23983 (N_23983,N_23120,N_23219);
or U23984 (N_23984,N_23229,N_23206);
xnor U23985 (N_23985,N_23364,N_23157);
and U23986 (N_23986,N_23418,N_23393);
or U23987 (N_23987,N_23395,N_23314);
nor U23988 (N_23988,N_23424,N_23375);
or U23989 (N_23989,N_23063,N_23079);
and U23990 (N_23990,N_23227,N_23073);
nor U23991 (N_23991,N_23232,N_23486);
and U23992 (N_23992,N_23420,N_23430);
or U23993 (N_23993,N_23444,N_23324);
xnor U23994 (N_23994,N_23387,N_23021);
xnor U23995 (N_23995,N_23371,N_23198);
and U23996 (N_23996,N_23318,N_23412);
nand U23997 (N_23997,N_23455,N_23433);
nor U23998 (N_23998,N_23229,N_23361);
xor U23999 (N_23999,N_23209,N_23464);
xor U24000 (N_24000,N_23662,N_23715);
nor U24001 (N_24001,N_23733,N_23777);
nand U24002 (N_24002,N_23543,N_23632);
xnor U24003 (N_24003,N_23775,N_23619);
or U24004 (N_24004,N_23982,N_23660);
and U24005 (N_24005,N_23669,N_23554);
nand U24006 (N_24006,N_23714,N_23833);
xnor U24007 (N_24007,N_23676,N_23559);
and U24008 (N_24008,N_23712,N_23514);
and U24009 (N_24009,N_23963,N_23689);
nand U24010 (N_24010,N_23779,N_23788);
nand U24011 (N_24011,N_23601,N_23919);
or U24012 (N_24012,N_23888,N_23599);
nand U24013 (N_24013,N_23500,N_23872);
and U24014 (N_24014,N_23761,N_23708);
xor U24015 (N_24015,N_23868,N_23939);
nor U24016 (N_24016,N_23925,N_23892);
nor U24017 (N_24017,N_23659,N_23582);
nor U24018 (N_24018,N_23757,N_23956);
xnor U24019 (N_24019,N_23501,N_23597);
or U24020 (N_24020,N_23807,N_23780);
nand U24021 (N_24021,N_23821,N_23759);
or U24022 (N_24022,N_23600,N_23851);
and U24023 (N_24023,N_23640,N_23639);
or U24024 (N_24024,N_23911,N_23756);
and U24025 (N_24025,N_23558,N_23881);
nor U24026 (N_24026,N_23535,N_23952);
nand U24027 (N_24027,N_23739,N_23529);
nand U24028 (N_24028,N_23837,N_23670);
xnor U24029 (N_24029,N_23920,N_23753);
xor U24030 (N_24030,N_23754,N_23655);
or U24031 (N_24031,N_23867,N_23572);
and U24032 (N_24032,N_23584,N_23637);
nand U24033 (N_24033,N_23947,N_23506);
and U24034 (N_24034,N_23738,N_23511);
and U24035 (N_24035,N_23841,N_23913);
nand U24036 (N_24036,N_23850,N_23521);
nand U24037 (N_24037,N_23745,N_23786);
xnor U24038 (N_24038,N_23908,N_23583);
and U24039 (N_24039,N_23541,N_23969);
and U24040 (N_24040,N_23813,N_23718);
and U24041 (N_24041,N_23871,N_23997);
and U24042 (N_24042,N_23800,N_23980);
nand U24043 (N_24043,N_23575,N_23882);
xor U24044 (N_24044,N_23773,N_23527);
nand U24045 (N_24045,N_23590,N_23612);
xnor U24046 (N_24046,N_23723,N_23649);
nor U24047 (N_24047,N_23697,N_23658);
nand U24048 (N_24048,N_23799,N_23949);
or U24049 (N_24049,N_23565,N_23921);
nand U24050 (N_24050,N_23776,N_23507);
xor U24051 (N_24051,N_23940,N_23705);
nor U24052 (N_24052,N_23825,N_23700);
and U24053 (N_24053,N_23695,N_23974);
xnor U24054 (N_24054,N_23645,N_23822);
nand U24055 (N_24055,N_23585,N_23664);
nor U24056 (N_24056,N_23861,N_23968);
nor U24057 (N_24057,N_23663,N_23741);
or U24058 (N_24058,N_23542,N_23883);
nor U24059 (N_24059,N_23654,N_23806);
nor U24060 (N_24060,N_23534,N_23557);
or U24061 (N_24061,N_23692,N_23631);
or U24062 (N_24062,N_23680,N_23914);
nand U24063 (N_24063,N_23604,N_23886);
nand U24064 (N_24064,N_23876,N_23657);
xor U24065 (N_24065,N_23628,N_23931);
xnor U24066 (N_24066,N_23652,N_23834);
or U24067 (N_24067,N_23711,N_23504);
or U24068 (N_24068,N_23661,N_23853);
nor U24069 (N_24069,N_23537,N_23643);
nand U24070 (N_24070,N_23991,N_23869);
nor U24071 (N_24071,N_23512,N_23625);
nand U24072 (N_24072,N_23993,N_23984);
nand U24073 (N_24073,N_23677,N_23577);
and U24074 (N_24074,N_23764,N_23587);
or U24075 (N_24075,N_23904,N_23889);
and U24076 (N_24076,N_23546,N_23835);
and U24077 (N_24077,N_23912,N_23752);
xnor U24078 (N_24078,N_23722,N_23790);
or U24079 (N_24079,N_23636,N_23578);
and U24080 (N_24080,N_23877,N_23962);
or U24081 (N_24081,N_23609,N_23593);
nand U24082 (N_24082,N_23784,N_23648);
nand U24083 (N_24083,N_23950,N_23610);
nand U24084 (N_24084,N_23944,N_23580);
xor U24085 (N_24085,N_23573,N_23895);
xor U24086 (N_24086,N_23890,N_23618);
and U24087 (N_24087,N_23792,N_23884);
nor U24088 (N_24088,N_23977,N_23897);
and U24089 (N_24089,N_23688,N_23617);
nor U24090 (N_24090,N_23513,N_23772);
and U24091 (N_24091,N_23734,N_23709);
nor U24092 (N_24092,N_23793,N_23523);
nand U24093 (N_24093,N_23975,N_23864);
nor U24094 (N_24094,N_23763,N_23650);
xor U24095 (N_24095,N_23926,N_23830);
nand U24096 (N_24096,N_23568,N_23614);
nor U24097 (N_24097,N_23874,N_23994);
xor U24098 (N_24098,N_23902,N_23638);
or U24099 (N_24099,N_23938,N_23725);
nand U24100 (N_24100,N_23603,N_23970);
and U24101 (N_24101,N_23951,N_23816);
or U24102 (N_24102,N_23880,N_23783);
nor U24103 (N_24103,N_23934,N_23943);
or U24104 (N_24104,N_23698,N_23948);
nor U24105 (N_24105,N_23656,N_23553);
nand U24106 (N_24106,N_23690,N_23887);
and U24107 (N_24107,N_23544,N_23740);
nand U24108 (N_24108,N_23804,N_23987);
nand U24109 (N_24109,N_23675,N_23995);
nor U24110 (N_24110,N_23898,N_23576);
xnor U24111 (N_24111,N_23860,N_23909);
or U24112 (N_24112,N_23906,N_23815);
and U24113 (N_24113,N_23955,N_23960);
xor U24114 (N_24114,N_23602,N_23567);
or U24115 (N_24115,N_23893,N_23809);
nor U24116 (N_24116,N_23642,N_23966);
xnor U24117 (N_24117,N_23717,N_23781);
nor U24118 (N_24118,N_23937,N_23929);
and U24119 (N_24119,N_23928,N_23569);
nand U24120 (N_24120,N_23641,N_23540);
and U24121 (N_24121,N_23996,N_23891);
or U24122 (N_24122,N_23682,N_23620);
and U24123 (N_24123,N_23588,N_23684);
nand U24124 (N_24124,N_23586,N_23563);
or U24125 (N_24125,N_23516,N_23693);
xor U24126 (N_24126,N_23976,N_23769);
nor U24127 (N_24127,N_23958,N_23515);
and U24128 (N_24128,N_23536,N_23899);
nor U24129 (N_24129,N_23802,N_23770);
xor U24130 (N_24130,N_23613,N_23621);
nor U24131 (N_24131,N_23696,N_23986);
nor U24132 (N_24132,N_23903,N_23627);
nor U24133 (N_24133,N_23701,N_23848);
or U24134 (N_24134,N_23924,N_23524);
nand U24135 (N_24135,N_23812,N_23870);
and U24136 (N_24136,N_23596,N_23798);
nand U24137 (N_24137,N_23724,N_23981);
or U24138 (N_24138,N_23917,N_23967);
and U24139 (N_24139,N_23828,N_23915);
xor U24140 (N_24140,N_23644,N_23748);
or U24141 (N_24141,N_23983,N_23607);
or U24142 (N_24142,N_23999,N_23556);
nor U24143 (N_24143,N_23747,N_23589);
xor U24144 (N_24144,N_23707,N_23771);
or U24145 (N_24145,N_23526,N_23824);
and U24146 (N_24146,N_23846,N_23819);
and U24147 (N_24147,N_23930,N_23918);
nand U24148 (N_24148,N_23594,N_23598);
and U24149 (N_24149,N_23672,N_23907);
xnor U24150 (N_24150,N_23579,N_23787);
or U24151 (N_24151,N_23863,N_23760);
or U24152 (N_24152,N_23901,N_23791);
nor U24153 (N_24153,N_23510,N_23946);
nand U24154 (N_24154,N_23750,N_23570);
nor U24155 (N_24155,N_23778,N_23520);
nand U24156 (N_24156,N_23623,N_23726);
nand U24157 (N_24157,N_23564,N_23933);
nand U24158 (N_24158,N_23615,N_23865);
or U24159 (N_24159,N_23562,N_23720);
xnor U24160 (N_24160,N_23730,N_23852);
and U24161 (N_24161,N_23716,N_23935);
or U24162 (N_24162,N_23885,N_23998);
or U24163 (N_24163,N_23679,N_23875);
or U24164 (N_24164,N_23561,N_23704);
or U24165 (N_24165,N_23719,N_23518);
xnor U24166 (N_24166,N_23762,N_23817);
or U24167 (N_24167,N_23606,N_23550);
or U24168 (N_24168,N_23910,N_23818);
and U24169 (N_24169,N_23706,N_23988);
nand U24170 (N_24170,N_23651,N_23808);
nor U24171 (N_24171,N_23743,N_23774);
nor U24172 (N_24172,N_23849,N_23635);
nand U24173 (N_24173,N_23517,N_23985);
nand U24174 (N_24174,N_23646,N_23765);
nand U24175 (N_24175,N_23687,N_23845);
nor U24176 (N_24176,N_23932,N_23878);
nand U24177 (N_24177,N_23629,N_23927);
or U24178 (N_24178,N_23710,N_23923);
or U24179 (N_24179,N_23810,N_23566);
or U24180 (N_24180,N_23595,N_23560);
xnor U24181 (N_24181,N_23842,N_23826);
or U24182 (N_24182,N_23694,N_23971);
and U24183 (N_24183,N_23840,N_23525);
or U24184 (N_24184,N_23746,N_23855);
xor U24185 (N_24185,N_23794,N_23916);
nand U24186 (N_24186,N_23736,N_23814);
and U24187 (N_24187,N_23699,N_23766);
and U24188 (N_24188,N_23796,N_23805);
and U24189 (N_24189,N_23729,N_23789);
or U24190 (N_24190,N_23608,N_23686);
xor U24191 (N_24191,N_23626,N_23528);
xor U24192 (N_24192,N_23989,N_23811);
or U24193 (N_24193,N_23674,N_23879);
or U24194 (N_24194,N_23744,N_23633);
nor U24195 (N_24195,N_23979,N_23768);
or U24196 (N_24196,N_23647,N_23862);
or U24197 (N_24197,N_23571,N_23592);
nor U24198 (N_24198,N_23803,N_23728);
and U24199 (N_24199,N_23555,N_23547);
xnor U24200 (N_24200,N_23847,N_23503);
and U24201 (N_24201,N_23702,N_23782);
nand U24202 (N_24202,N_23732,N_23795);
or U24203 (N_24203,N_23591,N_23936);
and U24204 (N_24204,N_23703,N_23973);
xnor U24205 (N_24205,N_23894,N_23866);
nor U24206 (N_24206,N_23519,N_23843);
nand U24207 (N_24207,N_23549,N_23678);
nand U24208 (N_24208,N_23727,N_23751);
or U24209 (N_24209,N_23505,N_23942);
nor U24210 (N_24210,N_23538,N_23823);
nand U24211 (N_24211,N_23616,N_23767);
nand U24212 (N_24212,N_23530,N_23838);
nand U24213 (N_24213,N_23539,N_23836);
nand U24214 (N_24214,N_23990,N_23856);
nor U24215 (N_24215,N_23522,N_23737);
nor U24216 (N_24216,N_23839,N_23622);
xor U24217 (N_24217,N_23574,N_23905);
nor U24218 (N_24218,N_23953,N_23666);
nand U24219 (N_24219,N_23755,N_23611);
and U24220 (N_24220,N_23531,N_23961);
and U24221 (N_24221,N_23832,N_23954);
or U24222 (N_24222,N_23873,N_23665);
nor U24223 (N_24223,N_23785,N_23992);
nand U24224 (N_24224,N_23581,N_23683);
or U24225 (N_24225,N_23713,N_23854);
or U24226 (N_24226,N_23858,N_23900);
nor U24227 (N_24227,N_23758,N_23671);
nand U24228 (N_24228,N_23630,N_23829);
xnor U24229 (N_24229,N_23673,N_23502);
xnor U24230 (N_24230,N_23957,N_23972);
nor U24231 (N_24231,N_23667,N_23721);
nand U24232 (N_24232,N_23681,N_23742);
or U24233 (N_24233,N_23797,N_23533);
nand U24234 (N_24234,N_23653,N_23634);
or U24235 (N_24235,N_23941,N_23545);
and U24236 (N_24236,N_23844,N_23959);
and U24237 (N_24237,N_23945,N_23978);
xor U24238 (N_24238,N_23691,N_23831);
nand U24239 (N_24239,N_23749,N_23685);
xor U24240 (N_24240,N_23820,N_23509);
and U24241 (N_24241,N_23605,N_23857);
nor U24242 (N_24242,N_23552,N_23922);
nand U24243 (N_24243,N_23548,N_23731);
and U24244 (N_24244,N_23508,N_23668);
and U24245 (N_24245,N_23532,N_23965);
or U24246 (N_24246,N_23801,N_23859);
or U24247 (N_24247,N_23827,N_23735);
and U24248 (N_24248,N_23624,N_23551);
nor U24249 (N_24249,N_23964,N_23896);
xnor U24250 (N_24250,N_23583,N_23769);
nand U24251 (N_24251,N_23764,N_23771);
nand U24252 (N_24252,N_23520,N_23960);
and U24253 (N_24253,N_23937,N_23977);
nor U24254 (N_24254,N_23770,N_23696);
and U24255 (N_24255,N_23637,N_23634);
or U24256 (N_24256,N_23501,N_23578);
nand U24257 (N_24257,N_23678,N_23587);
xnor U24258 (N_24258,N_23874,N_23701);
xor U24259 (N_24259,N_23669,N_23545);
xor U24260 (N_24260,N_23805,N_23607);
nor U24261 (N_24261,N_23521,N_23979);
nor U24262 (N_24262,N_23579,N_23562);
and U24263 (N_24263,N_23805,N_23716);
nor U24264 (N_24264,N_23646,N_23795);
nand U24265 (N_24265,N_23752,N_23544);
nor U24266 (N_24266,N_23654,N_23644);
or U24267 (N_24267,N_23764,N_23757);
xnor U24268 (N_24268,N_23835,N_23654);
nor U24269 (N_24269,N_23859,N_23917);
or U24270 (N_24270,N_23729,N_23893);
nand U24271 (N_24271,N_23770,N_23646);
nor U24272 (N_24272,N_23693,N_23737);
xor U24273 (N_24273,N_23816,N_23665);
and U24274 (N_24274,N_23664,N_23858);
or U24275 (N_24275,N_23545,N_23633);
and U24276 (N_24276,N_23913,N_23564);
nor U24277 (N_24277,N_23542,N_23529);
or U24278 (N_24278,N_23553,N_23597);
xor U24279 (N_24279,N_23568,N_23748);
nor U24280 (N_24280,N_23822,N_23958);
nor U24281 (N_24281,N_23871,N_23718);
or U24282 (N_24282,N_23868,N_23816);
xnor U24283 (N_24283,N_23759,N_23576);
and U24284 (N_24284,N_23601,N_23554);
nand U24285 (N_24285,N_23917,N_23896);
or U24286 (N_24286,N_23608,N_23844);
or U24287 (N_24287,N_23826,N_23629);
nand U24288 (N_24288,N_23917,N_23561);
nand U24289 (N_24289,N_23946,N_23847);
or U24290 (N_24290,N_23552,N_23675);
nand U24291 (N_24291,N_23613,N_23845);
xnor U24292 (N_24292,N_23896,N_23774);
nor U24293 (N_24293,N_23730,N_23876);
or U24294 (N_24294,N_23537,N_23707);
and U24295 (N_24295,N_23933,N_23531);
xor U24296 (N_24296,N_23661,N_23909);
nand U24297 (N_24297,N_23787,N_23564);
nor U24298 (N_24298,N_23999,N_23598);
or U24299 (N_24299,N_23991,N_23829);
and U24300 (N_24300,N_23704,N_23592);
xnor U24301 (N_24301,N_23711,N_23913);
nor U24302 (N_24302,N_23906,N_23793);
xnor U24303 (N_24303,N_23734,N_23950);
xnor U24304 (N_24304,N_23820,N_23537);
and U24305 (N_24305,N_23987,N_23781);
xor U24306 (N_24306,N_23642,N_23644);
nand U24307 (N_24307,N_23800,N_23505);
and U24308 (N_24308,N_23804,N_23551);
and U24309 (N_24309,N_23753,N_23659);
nand U24310 (N_24310,N_23528,N_23760);
nand U24311 (N_24311,N_23903,N_23758);
and U24312 (N_24312,N_23930,N_23913);
or U24313 (N_24313,N_23923,N_23680);
and U24314 (N_24314,N_23621,N_23909);
xor U24315 (N_24315,N_23632,N_23882);
xnor U24316 (N_24316,N_23723,N_23526);
or U24317 (N_24317,N_23611,N_23588);
xor U24318 (N_24318,N_23686,N_23784);
or U24319 (N_24319,N_23636,N_23568);
xnor U24320 (N_24320,N_23970,N_23733);
nand U24321 (N_24321,N_23517,N_23732);
or U24322 (N_24322,N_23778,N_23869);
nor U24323 (N_24323,N_23780,N_23676);
and U24324 (N_24324,N_23683,N_23884);
or U24325 (N_24325,N_23915,N_23618);
and U24326 (N_24326,N_23693,N_23748);
or U24327 (N_24327,N_23853,N_23707);
xnor U24328 (N_24328,N_23696,N_23851);
and U24329 (N_24329,N_23839,N_23812);
or U24330 (N_24330,N_23589,N_23786);
nand U24331 (N_24331,N_23722,N_23779);
or U24332 (N_24332,N_23630,N_23618);
and U24333 (N_24333,N_23982,N_23955);
nand U24334 (N_24334,N_23630,N_23727);
xnor U24335 (N_24335,N_23831,N_23829);
or U24336 (N_24336,N_23906,N_23634);
nor U24337 (N_24337,N_23827,N_23885);
or U24338 (N_24338,N_23715,N_23897);
and U24339 (N_24339,N_23850,N_23585);
nor U24340 (N_24340,N_23670,N_23785);
xor U24341 (N_24341,N_23658,N_23882);
or U24342 (N_24342,N_23577,N_23531);
nor U24343 (N_24343,N_23604,N_23613);
xor U24344 (N_24344,N_23728,N_23562);
xor U24345 (N_24345,N_23696,N_23755);
or U24346 (N_24346,N_23894,N_23654);
xnor U24347 (N_24347,N_23716,N_23871);
xor U24348 (N_24348,N_23922,N_23878);
xor U24349 (N_24349,N_23638,N_23605);
nand U24350 (N_24350,N_23585,N_23676);
nand U24351 (N_24351,N_23620,N_23929);
or U24352 (N_24352,N_23644,N_23820);
nand U24353 (N_24353,N_23665,N_23751);
or U24354 (N_24354,N_23897,N_23530);
xor U24355 (N_24355,N_23959,N_23784);
or U24356 (N_24356,N_23999,N_23578);
xor U24357 (N_24357,N_23677,N_23765);
and U24358 (N_24358,N_23703,N_23821);
or U24359 (N_24359,N_23881,N_23644);
and U24360 (N_24360,N_23624,N_23919);
xnor U24361 (N_24361,N_23562,N_23649);
nor U24362 (N_24362,N_23776,N_23753);
nor U24363 (N_24363,N_23504,N_23693);
nand U24364 (N_24364,N_23862,N_23522);
or U24365 (N_24365,N_23879,N_23615);
and U24366 (N_24366,N_23971,N_23608);
or U24367 (N_24367,N_23886,N_23540);
and U24368 (N_24368,N_23712,N_23611);
nand U24369 (N_24369,N_23519,N_23955);
nand U24370 (N_24370,N_23850,N_23736);
or U24371 (N_24371,N_23741,N_23810);
xor U24372 (N_24372,N_23661,N_23523);
nor U24373 (N_24373,N_23790,N_23842);
nor U24374 (N_24374,N_23555,N_23503);
nor U24375 (N_24375,N_23771,N_23967);
nor U24376 (N_24376,N_23528,N_23810);
nand U24377 (N_24377,N_23842,N_23800);
and U24378 (N_24378,N_23813,N_23693);
nor U24379 (N_24379,N_23790,N_23822);
xor U24380 (N_24380,N_23751,N_23708);
xor U24381 (N_24381,N_23690,N_23617);
nand U24382 (N_24382,N_23519,N_23526);
nor U24383 (N_24383,N_23884,N_23652);
or U24384 (N_24384,N_23820,N_23640);
nor U24385 (N_24385,N_23573,N_23649);
nand U24386 (N_24386,N_23978,N_23859);
nor U24387 (N_24387,N_23724,N_23528);
nor U24388 (N_24388,N_23572,N_23953);
or U24389 (N_24389,N_23511,N_23757);
and U24390 (N_24390,N_23944,N_23841);
nor U24391 (N_24391,N_23741,N_23559);
nor U24392 (N_24392,N_23625,N_23983);
nand U24393 (N_24393,N_23746,N_23665);
or U24394 (N_24394,N_23611,N_23634);
xor U24395 (N_24395,N_23819,N_23872);
nand U24396 (N_24396,N_23575,N_23994);
and U24397 (N_24397,N_23868,N_23554);
nand U24398 (N_24398,N_23571,N_23945);
xnor U24399 (N_24399,N_23987,N_23532);
nor U24400 (N_24400,N_23621,N_23567);
nand U24401 (N_24401,N_23941,N_23550);
or U24402 (N_24402,N_23806,N_23996);
and U24403 (N_24403,N_23945,N_23918);
xor U24404 (N_24404,N_23598,N_23559);
or U24405 (N_24405,N_23539,N_23733);
xor U24406 (N_24406,N_23758,N_23736);
and U24407 (N_24407,N_23721,N_23772);
or U24408 (N_24408,N_23642,N_23993);
nor U24409 (N_24409,N_23874,N_23628);
nor U24410 (N_24410,N_23534,N_23758);
nand U24411 (N_24411,N_23997,N_23998);
nor U24412 (N_24412,N_23756,N_23688);
and U24413 (N_24413,N_23536,N_23814);
nand U24414 (N_24414,N_23791,N_23555);
nand U24415 (N_24415,N_23595,N_23862);
nand U24416 (N_24416,N_23693,N_23604);
nand U24417 (N_24417,N_23811,N_23501);
nand U24418 (N_24418,N_23790,N_23980);
nand U24419 (N_24419,N_23905,N_23754);
xor U24420 (N_24420,N_23726,N_23743);
or U24421 (N_24421,N_23512,N_23724);
or U24422 (N_24422,N_23690,N_23686);
or U24423 (N_24423,N_23949,N_23579);
and U24424 (N_24424,N_23863,N_23574);
and U24425 (N_24425,N_23929,N_23792);
or U24426 (N_24426,N_23852,N_23779);
nor U24427 (N_24427,N_23512,N_23521);
nand U24428 (N_24428,N_23962,N_23504);
nor U24429 (N_24429,N_23910,N_23595);
or U24430 (N_24430,N_23965,N_23546);
xor U24431 (N_24431,N_23723,N_23918);
or U24432 (N_24432,N_23908,N_23657);
nand U24433 (N_24433,N_23775,N_23893);
xor U24434 (N_24434,N_23602,N_23639);
nand U24435 (N_24435,N_23506,N_23777);
nor U24436 (N_24436,N_23882,N_23579);
nor U24437 (N_24437,N_23823,N_23785);
or U24438 (N_24438,N_23694,N_23599);
or U24439 (N_24439,N_23770,N_23901);
nor U24440 (N_24440,N_23843,N_23827);
xor U24441 (N_24441,N_23767,N_23738);
xnor U24442 (N_24442,N_23910,N_23932);
and U24443 (N_24443,N_23519,N_23865);
nand U24444 (N_24444,N_23770,N_23924);
and U24445 (N_24445,N_23813,N_23655);
nor U24446 (N_24446,N_23820,N_23985);
and U24447 (N_24447,N_23771,N_23969);
xor U24448 (N_24448,N_23582,N_23856);
or U24449 (N_24449,N_23582,N_23566);
nor U24450 (N_24450,N_23508,N_23874);
nand U24451 (N_24451,N_23710,N_23579);
nand U24452 (N_24452,N_23852,N_23753);
nor U24453 (N_24453,N_23770,N_23891);
nand U24454 (N_24454,N_23956,N_23595);
xnor U24455 (N_24455,N_23862,N_23753);
or U24456 (N_24456,N_23526,N_23985);
nor U24457 (N_24457,N_23946,N_23773);
nor U24458 (N_24458,N_23521,N_23544);
or U24459 (N_24459,N_23603,N_23741);
nand U24460 (N_24460,N_23803,N_23731);
nand U24461 (N_24461,N_23913,N_23657);
nand U24462 (N_24462,N_23807,N_23643);
and U24463 (N_24463,N_23648,N_23575);
and U24464 (N_24464,N_23607,N_23928);
and U24465 (N_24465,N_23851,N_23619);
xor U24466 (N_24466,N_23589,N_23738);
and U24467 (N_24467,N_23734,N_23841);
nand U24468 (N_24468,N_23505,N_23920);
nand U24469 (N_24469,N_23679,N_23825);
xnor U24470 (N_24470,N_23663,N_23925);
nand U24471 (N_24471,N_23630,N_23652);
or U24472 (N_24472,N_23921,N_23527);
xnor U24473 (N_24473,N_23576,N_23856);
or U24474 (N_24474,N_23960,N_23673);
or U24475 (N_24475,N_23761,N_23962);
xnor U24476 (N_24476,N_23589,N_23769);
and U24477 (N_24477,N_23519,N_23746);
nand U24478 (N_24478,N_23699,N_23808);
or U24479 (N_24479,N_23675,N_23743);
nor U24480 (N_24480,N_23647,N_23503);
and U24481 (N_24481,N_23781,N_23821);
nand U24482 (N_24482,N_23991,N_23645);
nand U24483 (N_24483,N_23732,N_23534);
nor U24484 (N_24484,N_23578,N_23721);
nor U24485 (N_24485,N_23616,N_23588);
or U24486 (N_24486,N_23887,N_23847);
nand U24487 (N_24487,N_23927,N_23985);
or U24488 (N_24488,N_23577,N_23782);
nor U24489 (N_24489,N_23981,N_23945);
and U24490 (N_24490,N_23834,N_23520);
or U24491 (N_24491,N_23905,N_23556);
or U24492 (N_24492,N_23945,N_23645);
and U24493 (N_24493,N_23983,N_23588);
xnor U24494 (N_24494,N_23776,N_23511);
and U24495 (N_24495,N_23597,N_23637);
nand U24496 (N_24496,N_23981,N_23903);
or U24497 (N_24497,N_23602,N_23780);
xnor U24498 (N_24498,N_23600,N_23935);
xnor U24499 (N_24499,N_23754,N_23508);
or U24500 (N_24500,N_24171,N_24096);
or U24501 (N_24501,N_24234,N_24183);
nor U24502 (N_24502,N_24446,N_24182);
and U24503 (N_24503,N_24105,N_24447);
nor U24504 (N_24504,N_24225,N_24391);
and U24505 (N_24505,N_24005,N_24073);
nor U24506 (N_24506,N_24455,N_24349);
and U24507 (N_24507,N_24168,N_24437);
xor U24508 (N_24508,N_24232,N_24064);
nor U24509 (N_24509,N_24336,N_24240);
or U24510 (N_24510,N_24373,N_24244);
nand U24511 (N_24511,N_24486,N_24128);
or U24512 (N_24512,N_24425,N_24457);
and U24513 (N_24513,N_24039,N_24332);
nor U24514 (N_24514,N_24320,N_24024);
xnor U24515 (N_24515,N_24499,N_24348);
nand U24516 (N_24516,N_24169,N_24101);
xnor U24517 (N_24517,N_24372,N_24357);
nor U24518 (N_24518,N_24103,N_24401);
or U24519 (N_24519,N_24159,N_24152);
nand U24520 (N_24520,N_24335,N_24377);
nand U24521 (N_24521,N_24384,N_24160);
xor U24522 (N_24522,N_24371,N_24076);
nor U24523 (N_24523,N_24082,N_24350);
and U24524 (N_24524,N_24338,N_24172);
xor U24525 (N_24525,N_24154,N_24125);
xnor U24526 (N_24526,N_24390,N_24104);
nor U24527 (N_24527,N_24421,N_24268);
nor U24528 (N_24528,N_24204,N_24286);
and U24529 (N_24529,N_24111,N_24032);
and U24530 (N_24530,N_24131,N_24462);
nor U24531 (N_24531,N_24296,N_24444);
xor U24532 (N_24532,N_24334,N_24046);
and U24533 (N_24533,N_24189,N_24069);
xnor U24534 (N_24534,N_24496,N_24321);
nand U24535 (N_24535,N_24009,N_24043);
nor U24536 (N_24536,N_24048,N_24044);
xor U24537 (N_24537,N_24195,N_24379);
nand U24538 (N_24538,N_24074,N_24161);
nand U24539 (N_24539,N_24235,N_24414);
nor U24540 (N_24540,N_24280,N_24084);
and U24541 (N_24541,N_24156,N_24275);
nand U24542 (N_24542,N_24419,N_24192);
xor U24543 (N_24543,N_24187,N_24461);
or U24544 (N_24544,N_24456,N_24113);
or U24545 (N_24545,N_24214,N_24435);
nor U24546 (N_24546,N_24000,N_24155);
nand U24547 (N_24547,N_24114,N_24071);
nand U24548 (N_24548,N_24163,N_24400);
and U24549 (N_24549,N_24130,N_24300);
or U24550 (N_24550,N_24067,N_24145);
nand U24551 (N_24551,N_24418,N_24259);
and U24552 (N_24552,N_24339,N_24215);
or U24553 (N_24553,N_24281,N_24452);
and U24554 (N_24554,N_24135,N_24248);
and U24555 (N_24555,N_24303,N_24309);
nand U24556 (N_24556,N_24451,N_24245);
nand U24557 (N_24557,N_24424,N_24494);
nand U24558 (N_24558,N_24072,N_24266);
nand U24559 (N_24559,N_24075,N_24293);
nor U24560 (N_24560,N_24238,N_24016);
nand U24561 (N_24561,N_24138,N_24242);
or U24562 (N_24562,N_24106,N_24146);
nand U24563 (N_24563,N_24207,N_24487);
and U24564 (N_24564,N_24036,N_24180);
nand U24565 (N_24565,N_24026,N_24480);
xnor U24566 (N_24566,N_24177,N_24190);
or U24567 (N_24567,N_24299,N_24206);
nand U24568 (N_24568,N_24329,N_24353);
xnor U24569 (N_24569,N_24136,N_24053);
xnor U24570 (N_24570,N_24020,N_24313);
and U24571 (N_24571,N_24098,N_24038);
nand U24572 (N_24572,N_24316,N_24010);
nand U24573 (N_24573,N_24448,N_24258);
nand U24574 (N_24574,N_24228,N_24041);
xor U24575 (N_24575,N_24194,N_24360);
xnor U24576 (N_24576,N_24137,N_24199);
nand U24577 (N_24577,N_24202,N_24277);
and U24578 (N_24578,N_24148,N_24263);
nand U24579 (N_24579,N_24273,N_24237);
or U24580 (N_24580,N_24364,N_24388);
nand U24581 (N_24581,N_24328,N_24359);
or U24582 (N_24582,N_24251,N_24308);
and U24583 (N_24583,N_24100,N_24068);
and U24584 (N_24584,N_24031,N_24422);
or U24585 (N_24585,N_24257,N_24165);
and U24586 (N_24586,N_24395,N_24438);
or U24587 (N_24587,N_24093,N_24434);
nand U24588 (N_24588,N_24287,N_24013);
nand U24589 (N_24589,N_24459,N_24256);
nand U24590 (N_24590,N_24035,N_24077);
xor U24591 (N_24591,N_24483,N_24181);
xnor U24592 (N_24592,N_24198,N_24343);
nand U24593 (N_24593,N_24250,N_24099);
nand U24594 (N_24594,N_24352,N_24340);
and U24595 (N_24595,N_24231,N_24465);
and U24596 (N_24596,N_24209,N_24272);
xnor U24597 (N_24597,N_24021,N_24471);
nor U24598 (N_24598,N_24479,N_24179);
and U24599 (N_24599,N_24003,N_24351);
nand U24600 (N_24600,N_24089,N_24166);
xor U24601 (N_24601,N_24178,N_24366);
nor U24602 (N_24602,N_24430,N_24212);
or U24603 (N_24603,N_24324,N_24023);
nand U24604 (N_24604,N_24413,N_24055);
nor U24605 (N_24605,N_24243,N_24126);
nand U24606 (N_24606,N_24033,N_24274);
nand U24607 (N_24607,N_24185,N_24008);
xnor U24608 (N_24608,N_24197,N_24110);
nor U24609 (N_24609,N_24330,N_24186);
nand U24610 (N_24610,N_24019,N_24367);
and U24611 (N_24611,N_24375,N_24188);
or U24612 (N_24612,N_24354,N_24314);
nand U24613 (N_24613,N_24025,N_24174);
or U24614 (N_24614,N_24355,N_24470);
nor U24615 (N_24615,N_24345,N_24417);
xor U24616 (N_24616,N_24311,N_24376);
or U24617 (N_24617,N_24060,N_24405);
and U24618 (N_24618,N_24004,N_24489);
nand U24619 (N_24619,N_24219,N_24034);
xnor U24620 (N_24620,N_24065,N_24102);
xor U24621 (N_24621,N_24498,N_24382);
or U24622 (N_24622,N_24392,N_24014);
xor U24623 (N_24623,N_24306,N_24066);
or U24624 (N_24624,N_24001,N_24247);
nand U24625 (N_24625,N_24488,N_24403);
and U24626 (N_24626,N_24307,N_24327);
xor U24627 (N_24627,N_24426,N_24233);
nor U24628 (N_24628,N_24346,N_24433);
xnor U24629 (N_24629,N_24191,N_24216);
xor U24630 (N_24630,N_24284,N_24117);
and U24631 (N_24631,N_24201,N_24173);
nor U24632 (N_24632,N_24411,N_24460);
and U24633 (N_24633,N_24222,N_24112);
nor U24634 (N_24634,N_24213,N_24265);
nor U24635 (N_24635,N_24302,N_24141);
or U24636 (N_24636,N_24319,N_24081);
nor U24637 (N_24637,N_24029,N_24368);
xor U24638 (N_24638,N_24449,N_24078);
and U24639 (N_24639,N_24092,N_24333);
nor U24640 (N_24640,N_24261,N_24227);
nor U24641 (N_24641,N_24211,N_24383);
and U24642 (N_24642,N_24151,N_24436);
or U24643 (N_24643,N_24458,N_24429);
nor U24644 (N_24644,N_24223,N_24022);
xnor U24645 (N_24645,N_24057,N_24045);
nor U24646 (N_24646,N_24396,N_24279);
nor U24647 (N_24647,N_24415,N_24200);
or U24648 (N_24648,N_24063,N_24331);
or U24649 (N_24649,N_24080,N_24472);
and U24650 (N_24650,N_24475,N_24205);
nand U24651 (N_24651,N_24290,N_24495);
or U24652 (N_24652,N_24040,N_24030);
or U24653 (N_24653,N_24049,N_24252);
nor U24654 (N_24654,N_24469,N_24132);
nand U24655 (N_24655,N_24002,N_24229);
nor U24656 (N_24656,N_24399,N_24468);
xor U24657 (N_24657,N_24441,N_24369);
or U24658 (N_24658,N_24253,N_24176);
and U24659 (N_24659,N_24050,N_24362);
xnor U24660 (N_24660,N_24407,N_24109);
nor U24661 (N_24661,N_24341,N_24006);
or U24662 (N_24662,N_24018,N_24255);
xor U24663 (N_24663,N_24322,N_24028);
or U24664 (N_24664,N_24086,N_24363);
and U24665 (N_24665,N_24342,N_24164);
nor U24666 (N_24666,N_24094,N_24184);
xor U24667 (N_24667,N_24254,N_24052);
or U24668 (N_24668,N_24464,N_24267);
xor U24669 (N_24669,N_24440,N_24149);
and U24670 (N_24670,N_24467,N_24431);
and U24671 (N_24671,N_24393,N_24482);
and U24672 (N_24672,N_24450,N_24276);
xnor U24673 (N_24673,N_24133,N_24143);
xor U24674 (N_24674,N_24122,N_24397);
or U24675 (N_24675,N_24047,N_24158);
xnor U24676 (N_24676,N_24404,N_24042);
nor U24677 (N_24677,N_24297,N_24007);
nor U24678 (N_24678,N_24056,N_24466);
nand U24679 (N_24679,N_24153,N_24298);
or U24680 (N_24680,N_24017,N_24325);
xor U24681 (N_24681,N_24289,N_24485);
xor U24682 (N_24682,N_24090,N_24217);
nor U24683 (N_24683,N_24108,N_24323);
nand U24684 (N_24684,N_24374,N_24490);
xnor U24685 (N_24685,N_24295,N_24241);
or U24686 (N_24686,N_24292,N_24385);
and U24687 (N_24687,N_24365,N_24304);
and U24688 (N_24688,N_24142,N_24107);
and U24689 (N_24689,N_24134,N_24123);
or U24690 (N_24690,N_24398,N_24270);
xnor U24691 (N_24691,N_24370,N_24051);
nand U24692 (N_24692,N_24428,N_24079);
or U24693 (N_24693,N_24140,N_24484);
nor U24694 (N_24694,N_24406,N_24260);
nand U24695 (N_24695,N_24453,N_24119);
and U24696 (N_24696,N_24116,N_24118);
or U24697 (N_24697,N_24129,N_24271);
xnor U24698 (N_24698,N_24283,N_24492);
and U24699 (N_24699,N_24423,N_24095);
xnor U24700 (N_24700,N_24262,N_24127);
and U24701 (N_24701,N_24054,N_24378);
or U24702 (N_24702,N_24193,N_24124);
and U24703 (N_24703,N_24410,N_24394);
and U24704 (N_24704,N_24058,N_24224);
nor U24705 (N_24705,N_24062,N_24474);
and U24706 (N_24706,N_24445,N_24203);
nand U24707 (N_24707,N_24285,N_24463);
and U24708 (N_24708,N_24120,N_24037);
and U24709 (N_24709,N_24015,N_24477);
nand U24710 (N_24710,N_24220,N_24432);
xnor U24711 (N_24711,N_24121,N_24150);
or U24712 (N_24712,N_24497,N_24115);
nor U24713 (N_24713,N_24097,N_24409);
xnor U24714 (N_24714,N_24358,N_24381);
and U24715 (N_24715,N_24061,N_24088);
xnor U24716 (N_24716,N_24337,N_24291);
or U24717 (N_24717,N_24312,N_24236);
xnor U24718 (N_24718,N_24210,N_24175);
or U24719 (N_24719,N_24196,N_24442);
and U24720 (N_24720,N_24139,N_24361);
or U24721 (N_24721,N_24218,N_24157);
nand U24722 (N_24722,N_24239,N_24305);
and U24723 (N_24723,N_24294,N_24315);
nor U24724 (N_24724,N_24027,N_24389);
xor U24725 (N_24725,N_24481,N_24326);
xnor U24726 (N_24726,N_24221,N_24420);
or U24727 (N_24727,N_24012,N_24167);
nor U24728 (N_24728,N_24478,N_24170);
or U24729 (N_24729,N_24226,N_24246);
nand U24730 (N_24730,N_24347,N_24147);
nor U24731 (N_24731,N_24318,N_24083);
and U24732 (N_24732,N_24408,N_24317);
xnor U24733 (N_24733,N_24380,N_24230);
nand U24734 (N_24734,N_24091,N_24344);
or U24735 (N_24735,N_24473,N_24386);
or U24736 (N_24736,N_24491,N_24387);
xnor U24737 (N_24737,N_24310,N_24269);
xnor U24738 (N_24738,N_24454,N_24144);
and U24739 (N_24739,N_24412,N_24162);
or U24740 (N_24740,N_24264,N_24070);
nor U24741 (N_24741,N_24208,N_24282);
and U24742 (N_24742,N_24439,N_24493);
and U24743 (N_24743,N_24085,N_24301);
or U24744 (N_24744,N_24476,N_24443);
nand U24745 (N_24745,N_24416,N_24288);
nand U24746 (N_24746,N_24011,N_24402);
xnor U24747 (N_24747,N_24356,N_24278);
xor U24748 (N_24748,N_24087,N_24059);
xnor U24749 (N_24749,N_24427,N_24249);
nor U24750 (N_24750,N_24059,N_24377);
or U24751 (N_24751,N_24398,N_24250);
nor U24752 (N_24752,N_24309,N_24282);
and U24753 (N_24753,N_24159,N_24093);
xnor U24754 (N_24754,N_24163,N_24342);
or U24755 (N_24755,N_24215,N_24463);
nand U24756 (N_24756,N_24472,N_24377);
or U24757 (N_24757,N_24017,N_24151);
nor U24758 (N_24758,N_24393,N_24465);
and U24759 (N_24759,N_24265,N_24434);
nand U24760 (N_24760,N_24057,N_24425);
xnor U24761 (N_24761,N_24331,N_24186);
nor U24762 (N_24762,N_24178,N_24218);
and U24763 (N_24763,N_24196,N_24331);
or U24764 (N_24764,N_24300,N_24235);
nor U24765 (N_24765,N_24060,N_24435);
nor U24766 (N_24766,N_24201,N_24153);
or U24767 (N_24767,N_24259,N_24197);
or U24768 (N_24768,N_24233,N_24328);
nor U24769 (N_24769,N_24193,N_24474);
nor U24770 (N_24770,N_24412,N_24387);
or U24771 (N_24771,N_24124,N_24416);
and U24772 (N_24772,N_24275,N_24164);
nor U24773 (N_24773,N_24491,N_24179);
nand U24774 (N_24774,N_24400,N_24264);
nor U24775 (N_24775,N_24388,N_24307);
nor U24776 (N_24776,N_24355,N_24026);
and U24777 (N_24777,N_24450,N_24201);
nand U24778 (N_24778,N_24123,N_24014);
nor U24779 (N_24779,N_24209,N_24070);
nand U24780 (N_24780,N_24397,N_24181);
nor U24781 (N_24781,N_24071,N_24115);
nor U24782 (N_24782,N_24336,N_24074);
and U24783 (N_24783,N_24186,N_24160);
and U24784 (N_24784,N_24358,N_24407);
xnor U24785 (N_24785,N_24014,N_24425);
or U24786 (N_24786,N_24348,N_24130);
xor U24787 (N_24787,N_24065,N_24048);
and U24788 (N_24788,N_24316,N_24225);
and U24789 (N_24789,N_24435,N_24109);
and U24790 (N_24790,N_24313,N_24153);
or U24791 (N_24791,N_24388,N_24101);
nand U24792 (N_24792,N_24267,N_24444);
xor U24793 (N_24793,N_24496,N_24361);
or U24794 (N_24794,N_24484,N_24185);
and U24795 (N_24795,N_24413,N_24421);
and U24796 (N_24796,N_24064,N_24434);
and U24797 (N_24797,N_24389,N_24230);
or U24798 (N_24798,N_24008,N_24336);
nand U24799 (N_24799,N_24304,N_24419);
nor U24800 (N_24800,N_24206,N_24189);
and U24801 (N_24801,N_24455,N_24212);
nor U24802 (N_24802,N_24032,N_24227);
xnor U24803 (N_24803,N_24482,N_24146);
nor U24804 (N_24804,N_24085,N_24441);
nand U24805 (N_24805,N_24339,N_24369);
and U24806 (N_24806,N_24481,N_24459);
and U24807 (N_24807,N_24002,N_24324);
or U24808 (N_24808,N_24011,N_24466);
xnor U24809 (N_24809,N_24387,N_24401);
and U24810 (N_24810,N_24242,N_24199);
xnor U24811 (N_24811,N_24360,N_24286);
xor U24812 (N_24812,N_24338,N_24424);
xor U24813 (N_24813,N_24357,N_24110);
and U24814 (N_24814,N_24009,N_24003);
xnor U24815 (N_24815,N_24409,N_24157);
nand U24816 (N_24816,N_24387,N_24310);
and U24817 (N_24817,N_24105,N_24359);
or U24818 (N_24818,N_24361,N_24196);
and U24819 (N_24819,N_24261,N_24223);
or U24820 (N_24820,N_24147,N_24002);
and U24821 (N_24821,N_24171,N_24090);
or U24822 (N_24822,N_24424,N_24276);
xor U24823 (N_24823,N_24127,N_24490);
xor U24824 (N_24824,N_24040,N_24055);
or U24825 (N_24825,N_24130,N_24265);
nor U24826 (N_24826,N_24446,N_24275);
nand U24827 (N_24827,N_24053,N_24184);
xnor U24828 (N_24828,N_24094,N_24409);
xor U24829 (N_24829,N_24086,N_24059);
and U24830 (N_24830,N_24434,N_24016);
nor U24831 (N_24831,N_24223,N_24449);
xor U24832 (N_24832,N_24381,N_24236);
nand U24833 (N_24833,N_24124,N_24047);
nor U24834 (N_24834,N_24435,N_24428);
nor U24835 (N_24835,N_24448,N_24151);
nor U24836 (N_24836,N_24156,N_24233);
nand U24837 (N_24837,N_24295,N_24104);
and U24838 (N_24838,N_24319,N_24470);
or U24839 (N_24839,N_24034,N_24426);
nor U24840 (N_24840,N_24118,N_24430);
or U24841 (N_24841,N_24295,N_24461);
nor U24842 (N_24842,N_24280,N_24133);
or U24843 (N_24843,N_24230,N_24241);
nand U24844 (N_24844,N_24312,N_24478);
xnor U24845 (N_24845,N_24038,N_24071);
or U24846 (N_24846,N_24496,N_24059);
and U24847 (N_24847,N_24014,N_24085);
nor U24848 (N_24848,N_24169,N_24042);
nand U24849 (N_24849,N_24025,N_24030);
nand U24850 (N_24850,N_24469,N_24420);
nand U24851 (N_24851,N_24166,N_24422);
xnor U24852 (N_24852,N_24158,N_24028);
nand U24853 (N_24853,N_24097,N_24378);
nor U24854 (N_24854,N_24004,N_24412);
nand U24855 (N_24855,N_24333,N_24180);
nor U24856 (N_24856,N_24470,N_24298);
xor U24857 (N_24857,N_24012,N_24351);
or U24858 (N_24858,N_24492,N_24202);
xnor U24859 (N_24859,N_24214,N_24154);
or U24860 (N_24860,N_24419,N_24229);
and U24861 (N_24861,N_24274,N_24175);
or U24862 (N_24862,N_24499,N_24254);
nand U24863 (N_24863,N_24148,N_24100);
and U24864 (N_24864,N_24286,N_24018);
xnor U24865 (N_24865,N_24168,N_24197);
nor U24866 (N_24866,N_24420,N_24267);
and U24867 (N_24867,N_24044,N_24083);
xor U24868 (N_24868,N_24368,N_24351);
or U24869 (N_24869,N_24265,N_24472);
xor U24870 (N_24870,N_24476,N_24072);
or U24871 (N_24871,N_24054,N_24243);
nand U24872 (N_24872,N_24072,N_24315);
xor U24873 (N_24873,N_24456,N_24191);
nor U24874 (N_24874,N_24313,N_24451);
and U24875 (N_24875,N_24377,N_24364);
and U24876 (N_24876,N_24314,N_24376);
nor U24877 (N_24877,N_24498,N_24455);
nor U24878 (N_24878,N_24237,N_24178);
xnor U24879 (N_24879,N_24293,N_24462);
nand U24880 (N_24880,N_24051,N_24365);
and U24881 (N_24881,N_24039,N_24481);
or U24882 (N_24882,N_24334,N_24028);
nor U24883 (N_24883,N_24119,N_24040);
and U24884 (N_24884,N_24024,N_24180);
nor U24885 (N_24885,N_24137,N_24186);
xnor U24886 (N_24886,N_24341,N_24362);
xnor U24887 (N_24887,N_24002,N_24409);
nor U24888 (N_24888,N_24472,N_24091);
xor U24889 (N_24889,N_24100,N_24375);
nand U24890 (N_24890,N_24290,N_24320);
nand U24891 (N_24891,N_24348,N_24092);
or U24892 (N_24892,N_24270,N_24339);
or U24893 (N_24893,N_24398,N_24389);
nand U24894 (N_24894,N_24264,N_24363);
xnor U24895 (N_24895,N_24073,N_24422);
xnor U24896 (N_24896,N_24040,N_24197);
nor U24897 (N_24897,N_24162,N_24327);
and U24898 (N_24898,N_24479,N_24375);
or U24899 (N_24899,N_24068,N_24345);
nand U24900 (N_24900,N_24083,N_24441);
xnor U24901 (N_24901,N_24407,N_24287);
nand U24902 (N_24902,N_24240,N_24236);
xnor U24903 (N_24903,N_24053,N_24066);
nand U24904 (N_24904,N_24498,N_24221);
or U24905 (N_24905,N_24004,N_24224);
nor U24906 (N_24906,N_24153,N_24177);
and U24907 (N_24907,N_24471,N_24058);
nand U24908 (N_24908,N_24161,N_24387);
nor U24909 (N_24909,N_24210,N_24472);
and U24910 (N_24910,N_24210,N_24409);
and U24911 (N_24911,N_24457,N_24025);
nor U24912 (N_24912,N_24313,N_24007);
nor U24913 (N_24913,N_24049,N_24275);
and U24914 (N_24914,N_24043,N_24139);
xnor U24915 (N_24915,N_24010,N_24322);
xor U24916 (N_24916,N_24277,N_24050);
and U24917 (N_24917,N_24272,N_24205);
nor U24918 (N_24918,N_24224,N_24285);
or U24919 (N_24919,N_24144,N_24178);
nor U24920 (N_24920,N_24483,N_24242);
or U24921 (N_24921,N_24174,N_24240);
or U24922 (N_24922,N_24212,N_24271);
and U24923 (N_24923,N_24091,N_24467);
and U24924 (N_24924,N_24000,N_24132);
nor U24925 (N_24925,N_24401,N_24282);
and U24926 (N_24926,N_24447,N_24436);
nor U24927 (N_24927,N_24249,N_24012);
nor U24928 (N_24928,N_24279,N_24381);
nand U24929 (N_24929,N_24449,N_24308);
or U24930 (N_24930,N_24281,N_24249);
and U24931 (N_24931,N_24204,N_24068);
nand U24932 (N_24932,N_24351,N_24204);
xor U24933 (N_24933,N_24108,N_24256);
or U24934 (N_24934,N_24076,N_24485);
or U24935 (N_24935,N_24047,N_24462);
nand U24936 (N_24936,N_24224,N_24399);
or U24937 (N_24937,N_24436,N_24027);
or U24938 (N_24938,N_24498,N_24057);
nor U24939 (N_24939,N_24177,N_24342);
xnor U24940 (N_24940,N_24061,N_24331);
or U24941 (N_24941,N_24028,N_24432);
and U24942 (N_24942,N_24154,N_24063);
or U24943 (N_24943,N_24414,N_24363);
nand U24944 (N_24944,N_24206,N_24030);
and U24945 (N_24945,N_24033,N_24237);
nand U24946 (N_24946,N_24424,N_24250);
and U24947 (N_24947,N_24146,N_24484);
nor U24948 (N_24948,N_24092,N_24057);
nor U24949 (N_24949,N_24434,N_24068);
nor U24950 (N_24950,N_24271,N_24390);
and U24951 (N_24951,N_24335,N_24228);
nor U24952 (N_24952,N_24198,N_24285);
and U24953 (N_24953,N_24375,N_24260);
nand U24954 (N_24954,N_24281,N_24079);
and U24955 (N_24955,N_24156,N_24050);
nor U24956 (N_24956,N_24070,N_24301);
nor U24957 (N_24957,N_24373,N_24428);
or U24958 (N_24958,N_24450,N_24251);
and U24959 (N_24959,N_24032,N_24095);
or U24960 (N_24960,N_24207,N_24471);
and U24961 (N_24961,N_24359,N_24278);
nand U24962 (N_24962,N_24353,N_24125);
xnor U24963 (N_24963,N_24252,N_24137);
nand U24964 (N_24964,N_24018,N_24212);
nand U24965 (N_24965,N_24135,N_24110);
or U24966 (N_24966,N_24108,N_24291);
xor U24967 (N_24967,N_24373,N_24408);
nor U24968 (N_24968,N_24186,N_24282);
and U24969 (N_24969,N_24256,N_24027);
nand U24970 (N_24970,N_24337,N_24418);
nand U24971 (N_24971,N_24315,N_24203);
or U24972 (N_24972,N_24339,N_24022);
or U24973 (N_24973,N_24022,N_24318);
and U24974 (N_24974,N_24128,N_24115);
nand U24975 (N_24975,N_24084,N_24164);
nor U24976 (N_24976,N_24296,N_24358);
or U24977 (N_24977,N_24360,N_24312);
or U24978 (N_24978,N_24179,N_24010);
nor U24979 (N_24979,N_24063,N_24210);
or U24980 (N_24980,N_24410,N_24095);
nand U24981 (N_24981,N_24497,N_24060);
nor U24982 (N_24982,N_24171,N_24150);
nor U24983 (N_24983,N_24357,N_24077);
nor U24984 (N_24984,N_24274,N_24134);
or U24985 (N_24985,N_24396,N_24468);
nor U24986 (N_24986,N_24231,N_24209);
and U24987 (N_24987,N_24156,N_24299);
nor U24988 (N_24988,N_24276,N_24174);
nor U24989 (N_24989,N_24446,N_24044);
nor U24990 (N_24990,N_24007,N_24289);
nand U24991 (N_24991,N_24447,N_24217);
nand U24992 (N_24992,N_24078,N_24362);
nor U24993 (N_24993,N_24162,N_24181);
nor U24994 (N_24994,N_24250,N_24039);
xnor U24995 (N_24995,N_24067,N_24326);
xor U24996 (N_24996,N_24484,N_24025);
and U24997 (N_24997,N_24497,N_24091);
and U24998 (N_24998,N_24033,N_24295);
xnor U24999 (N_24999,N_24095,N_24252);
nand U25000 (N_25000,N_24886,N_24777);
xnor U25001 (N_25001,N_24993,N_24916);
nor U25002 (N_25002,N_24589,N_24878);
or U25003 (N_25003,N_24781,N_24674);
xnor U25004 (N_25004,N_24784,N_24561);
nand U25005 (N_25005,N_24556,N_24707);
and U25006 (N_25006,N_24900,N_24542);
xor U25007 (N_25007,N_24939,N_24554);
xor U25008 (N_25008,N_24563,N_24823);
nand U25009 (N_25009,N_24789,N_24779);
xnor U25010 (N_25010,N_24955,N_24545);
nor U25011 (N_25011,N_24767,N_24866);
nor U25012 (N_25012,N_24942,N_24530);
and U25013 (N_25013,N_24731,N_24967);
and U25014 (N_25014,N_24816,N_24696);
xnor U25015 (N_25015,N_24758,N_24596);
and U25016 (N_25016,N_24843,N_24629);
xor U25017 (N_25017,N_24990,N_24863);
or U25018 (N_25018,N_24951,N_24883);
and U25019 (N_25019,N_24714,N_24922);
or U25020 (N_25020,N_24943,N_24601);
or U25021 (N_25021,N_24756,N_24931);
or U25022 (N_25022,N_24928,N_24812);
nor U25023 (N_25023,N_24617,N_24595);
nor U25024 (N_25024,N_24902,N_24745);
xnor U25025 (N_25025,N_24853,N_24628);
and U25026 (N_25026,N_24988,N_24734);
nand U25027 (N_25027,N_24665,N_24537);
and U25028 (N_25028,N_24568,N_24898);
xor U25029 (N_25029,N_24792,N_24847);
nand U25030 (N_25030,N_24606,N_24856);
nand U25031 (N_25031,N_24526,N_24814);
or U25032 (N_25032,N_24936,N_24641);
xnor U25033 (N_25033,N_24509,N_24581);
nor U25034 (N_25034,N_24803,N_24919);
nor U25035 (N_25035,N_24840,N_24875);
nor U25036 (N_25036,N_24819,N_24887);
and U25037 (N_25037,N_24656,N_24712);
nand U25038 (N_25038,N_24686,N_24682);
xnor U25039 (N_25039,N_24820,N_24986);
or U25040 (N_25040,N_24753,N_24760);
xor U25041 (N_25041,N_24549,N_24927);
xnor U25042 (N_25042,N_24857,N_24764);
nor U25043 (N_25043,N_24889,N_24982);
or U25044 (N_25044,N_24852,N_24829);
nor U25045 (N_25045,N_24685,N_24564);
and U25046 (N_25046,N_24858,N_24653);
and U25047 (N_25047,N_24867,N_24778);
nand U25048 (N_25048,N_24799,N_24703);
nor U25049 (N_25049,N_24985,N_24839);
and U25050 (N_25050,N_24648,N_24626);
or U25051 (N_25051,N_24968,N_24773);
xnor U25052 (N_25052,N_24582,N_24870);
nor U25053 (N_25053,N_24972,N_24520);
nand U25054 (N_25054,N_24695,N_24506);
nand U25055 (N_25055,N_24925,N_24527);
nor U25056 (N_25056,N_24590,N_24908);
and U25057 (N_25057,N_24701,N_24638);
nor U25058 (N_25058,N_24871,N_24678);
nor U25059 (N_25059,N_24669,N_24736);
nand U25060 (N_25060,N_24947,N_24591);
or U25061 (N_25061,N_24598,N_24924);
xor U25062 (N_25062,N_24605,N_24964);
and U25063 (N_25063,N_24969,N_24644);
and U25064 (N_25064,N_24739,N_24607);
xnor U25065 (N_25065,N_24907,N_24504);
nor U25066 (N_25066,N_24539,N_24592);
xor U25067 (N_25067,N_24802,N_24865);
nor U25068 (N_25068,N_24921,N_24555);
xor U25069 (N_25069,N_24827,N_24622);
nand U25070 (N_25070,N_24965,N_24643);
xor U25071 (N_25071,N_24891,N_24660);
or U25072 (N_25072,N_24973,N_24721);
and U25073 (N_25073,N_24646,N_24516);
xnor U25074 (N_25074,N_24511,N_24888);
xnor U25075 (N_25075,N_24818,N_24904);
nor U25076 (N_25076,N_24838,N_24998);
or U25077 (N_25077,N_24882,N_24810);
or U25078 (N_25078,N_24880,N_24740);
nand U25079 (N_25079,N_24979,N_24984);
or U25080 (N_25080,N_24860,N_24726);
or U25081 (N_25081,N_24541,N_24672);
nor U25082 (N_25082,N_24748,N_24710);
or U25083 (N_25083,N_24661,N_24876);
xor U25084 (N_25084,N_24742,N_24879);
nor U25085 (N_25085,N_24873,N_24536);
xor U25086 (N_25086,N_24649,N_24835);
and U25087 (N_25087,N_24851,N_24558);
and U25088 (N_25088,N_24794,N_24708);
and U25089 (N_25089,N_24978,N_24691);
or U25090 (N_25090,N_24671,N_24687);
nand U25091 (N_25091,N_24930,N_24914);
xor U25092 (N_25092,N_24747,N_24750);
and U25093 (N_25093,N_24722,N_24694);
nor U25094 (N_25094,N_24632,N_24732);
or U25095 (N_25095,N_24983,N_24651);
nand U25096 (N_25096,N_24533,N_24776);
or U25097 (N_25097,N_24627,N_24946);
or U25098 (N_25098,N_24807,N_24974);
or U25099 (N_25099,N_24593,N_24510);
nand U25100 (N_25100,N_24508,N_24705);
nand U25101 (N_25101,N_24738,N_24833);
and U25102 (N_25102,N_24692,N_24825);
xnor U25103 (N_25103,N_24597,N_24676);
and U25104 (N_25104,N_24585,N_24521);
or U25105 (N_25105,N_24956,N_24751);
xnor U25106 (N_25106,N_24728,N_24937);
or U25107 (N_25107,N_24514,N_24911);
nand U25108 (N_25108,N_24980,N_24841);
or U25109 (N_25109,N_24614,N_24602);
and U25110 (N_25110,N_24971,N_24884);
and U25111 (N_25111,N_24952,N_24583);
nand U25112 (N_25112,N_24567,N_24757);
nor U25113 (N_25113,N_24633,N_24821);
xnor U25114 (N_25114,N_24795,N_24892);
nor U25115 (N_25115,N_24670,N_24501);
nand U25116 (N_25116,N_24548,N_24899);
xnor U25117 (N_25117,N_24553,N_24640);
or U25118 (N_25118,N_24940,N_24618);
nand U25119 (N_25119,N_24890,N_24689);
nor U25120 (N_25120,N_24552,N_24645);
nand U25121 (N_25121,N_24797,N_24538);
nor U25122 (N_25122,N_24845,N_24918);
xor U25123 (N_25123,N_24735,N_24953);
or U25124 (N_25124,N_24636,N_24805);
nor U25125 (N_25125,N_24609,N_24631);
nor U25126 (N_25126,N_24733,N_24948);
xor U25127 (N_25127,N_24588,N_24775);
and U25128 (N_25128,N_24711,N_24994);
nor U25129 (N_25129,N_24662,N_24547);
nor U25130 (N_25130,N_24848,N_24611);
or U25131 (N_25131,N_24949,N_24769);
and U25132 (N_25132,N_24737,N_24862);
nor U25133 (N_25133,N_24809,N_24824);
or U25134 (N_25134,N_24771,N_24713);
nand U25135 (N_25135,N_24715,N_24724);
nand U25136 (N_25136,N_24718,N_24950);
or U25137 (N_25137,N_24761,N_24762);
and U25138 (N_25138,N_24657,N_24546);
nor U25139 (N_25139,N_24906,N_24650);
or U25140 (N_25140,N_24855,N_24594);
or U25141 (N_25141,N_24868,N_24954);
xnor U25142 (N_25142,N_24704,N_24575);
nor U25143 (N_25143,N_24741,N_24804);
xor U25144 (N_25144,N_24752,N_24897);
nand U25145 (N_25145,N_24620,N_24569);
xnor U25146 (N_25146,N_24634,N_24859);
or U25147 (N_25147,N_24828,N_24912);
or U25148 (N_25148,N_24793,N_24673);
or U25149 (N_25149,N_24850,N_24987);
nand U25150 (N_25150,N_24920,N_24540);
xnor U25151 (N_25151,N_24608,N_24668);
nand U25152 (N_25152,N_24624,N_24679);
nand U25153 (N_25153,N_24615,N_24832);
nor U25154 (N_25154,N_24677,N_24528);
and U25155 (N_25155,N_24621,N_24500);
nor U25156 (N_25156,N_24997,N_24522);
nand U25157 (N_25157,N_24959,N_24610);
nor U25158 (N_25158,N_24532,N_24861);
nand U25159 (N_25159,N_24765,N_24977);
xnor U25160 (N_25160,N_24958,N_24702);
nor U25161 (N_25161,N_24562,N_24523);
and U25162 (N_25162,N_24512,N_24680);
and U25163 (N_25163,N_24642,N_24637);
and U25164 (N_25164,N_24697,N_24603);
and U25165 (N_25165,N_24658,N_24749);
and U25166 (N_25166,N_24580,N_24565);
nand U25167 (N_25167,N_24559,N_24616);
nand U25168 (N_25168,N_24830,N_24913);
and U25169 (N_25169,N_24699,N_24744);
and U25170 (N_25170,N_24652,N_24881);
and U25171 (N_25171,N_24566,N_24577);
nor U25172 (N_25172,N_24507,N_24935);
and U25173 (N_25173,N_24957,N_24966);
or U25174 (N_25174,N_24944,N_24550);
xor U25175 (N_25175,N_24877,N_24534);
and U25176 (N_25176,N_24716,N_24801);
xnor U25177 (N_25177,N_24806,N_24574);
nand U25178 (N_25178,N_24782,N_24630);
or U25179 (N_25179,N_24725,N_24837);
and U25180 (N_25180,N_24926,N_24570);
or U25181 (N_25181,N_24654,N_24573);
and U25182 (N_25182,N_24667,N_24992);
and U25183 (N_25183,N_24743,N_24639);
nor U25184 (N_25184,N_24834,N_24791);
or U25185 (N_25185,N_24976,N_24675);
or U25186 (N_25186,N_24576,N_24901);
xor U25187 (N_25187,N_24783,N_24766);
nand U25188 (N_25188,N_24720,N_24960);
and U25189 (N_25189,N_24655,N_24836);
nor U25190 (N_25190,N_24513,N_24730);
and U25191 (N_25191,N_24719,N_24529);
and U25192 (N_25192,N_24941,N_24619);
xor U25193 (N_25193,N_24915,N_24842);
xnor U25194 (N_25194,N_24932,N_24826);
and U25195 (N_25195,N_24613,N_24663);
nand U25196 (N_25196,N_24989,N_24535);
or U25197 (N_25197,N_24854,N_24917);
nor U25198 (N_25198,N_24659,N_24578);
and U25199 (N_25199,N_24893,N_24808);
or U25200 (N_25200,N_24869,N_24923);
or U25201 (N_25201,N_24698,N_24505);
nor U25202 (N_25202,N_24683,N_24772);
and U25203 (N_25203,N_24962,N_24933);
nand U25204 (N_25204,N_24587,N_24625);
or U25205 (N_25205,N_24584,N_24961);
nand U25206 (N_25206,N_24770,N_24690);
or U25207 (N_25207,N_24813,N_24785);
and U25208 (N_25208,N_24991,N_24709);
and U25209 (N_25209,N_24945,N_24786);
or U25210 (N_25210,N_24503,N_24934);
nor U25211 (N_25211,N_24684,N_24717);
and U25212 (N_25212,N_24763,N_24963);
or U25213 (N_25213,N_24600,N_24754);
or U25214 (N_25214,N_24688,N_24896);
xor U25215 (N_25215,N_24790,N_24664);
and U25216 (N_25216,N_24905,N_24727);
xnor U25217 (N_25217,N_24515,N_24759);
or U25218 (N_25218,N_24604,N_24844);
nand U25219 (N_25219,N_24551,N_24681);
xnor U25220 (N_25220,N_24910,N_24846);
nor U25221 (N_25221,N_24519,N_24502);
or U25222 (N_25222,N_24822,N_24815);
and U25223 (N_25223,N_24755,N_24938);
or U25224 (N_25224,N_24723,N_24872);
or U25225 (N_25225,N_24929,N_24864);
or U25226 (N_25226,N_24996,N_24811);
nor U25227 (N_25227,N_24531,N_24524);
nor U25228 (N_25228,N_24995,N_24557);
or U25229 (N_25229,N_24612,N_24903);
or U25230 (N_25230,N_24975,N_24543);
or U25231 (N_25231,N_24849,N_24831);
nand U25232 (N_25232,N_24798,N_24746);
xnor U25233 (N_25233,N_24700,N_24788);
nor U25234 (N_25234,N_24666,N_24729);
nand U25235 (N_25235,N_24599,N_24774);
nand U25236 (N_25236,N_24572,N_24800);
nor U25237 (N_25237,N_24571,N_24525);
xor U25238 (N_25238,N_24693,N_24895);
or U25239 (N_25239,N_24909,N_24885);
nand U25240 (N_25240,N_24517,N_24874);
nand U25241 (N_25241,N_24817,N_24635);
and U25242 (N_25242,N_24518,N_24787);
and U25243 (N_25243,N_24623,N_24970);
xor U25244 (N_25244,N_24999,N_24981);
or U25245 (N_25245,N_24586,N_24796);
and U25246 (N_25246,N_24768,N_24780);
and U25247 (N_25247,N_24894,N_24560);
xnor U25248 (N_25248,N_24647,N_24544);
nand U25249 (N_25249,N_24579,N_24706);
nand U25250 (N_25250,N_24915,N_24745);
nand U25251 (N_25251,N_24681,N_24925);
and U25252 (N_25252,N_24742,N_24829);
nand U25253 (N_25253,N_24668,N_24642);
xnor U25254 (N_25254,N_24942,N_24605);
nor U25255 (N_25255,N_24985,N_24958);
nor U25256 (N_25256,N_24617,N_24833);
nor U25257 (N_25257,N_24641,N_24996);
and U25258 (N_25258,N_24957,N_24984);
and U25259 (N_25259,N_24671,N_24956);
and U25260 (N_25260,N_24703,N_24792);
xnor U25261 (N_25261,N_24980,N_24872);
or U25262 (N_25262,N_24791,N_24698);
xnor U25263 (N_25263,N_24957,N_24702);
or U25264 (N_25264,N_24509,N_24897);
nand U25265 (N_25265,N_24982,N_24906);
or U25266 (N_25266,N_24816,N_24632);
nand U25267 (N_25267,N_24946,N_24933);
xnor U25268 (N_25268,N_24816,N_24515);
nor U25269 (N_25269,N_24835,N_24939);
or U25270 (N_25270,N_24812,N_24878);
nor U25271 (N_25271,N_24604,N_24611);
nand U25272 (N_25272,N_24850,N_24957);
nor U25273 (N_25273,N_24733,N_24506);
nor U25274 (N_25274,N_24724,N_24684);
or U25275 (N_25275,N_24626,N_24986);
and U25276 (N_25276,N_24649,N_24549);
nand U25277 (N_25277,N_24507,N_24833);
xor U25278 (N_25278,N_24948,N_24944);
nor U25279 (N_25279,N_24613,N_24784);
nor U25280 (N_25280,N_24525,N_24897);
and U25281 (N_25281,N_24768,N_24562);
xnor U25282 (N_25282,N_24617,N_24607);
and U25283 (N_25283,N_24936,N_24930);
xnor U25284 (N_25284,N_24962,N_24593);
nor U25285 (N_25285,N_24723,N_24649);
nor U25286 (N_25286,N_24628,N_24515);
and U25287 (N_25287,N_24506,N_24711);
nor U25288 (N_25288,N_24524,N_24745);
xor U25289 (N_25289,N_24880,N_24998);
nand U25290 (N_25290,N_24845,N_24533);
xnor U25291 (N_25291,N_24990,N_24875);
xnor U25292 (N_25292,N_24704,N_24845);
xor U25293 (N_25293,N_24697,N_24898);
or U25294 (N_25294,N_24527,N_24766);
and U25295 (N_25295,N_24731,N_24691);
xor U25296 (N_25296,N_24765,N_24827);
nand U25297 (N_25297,N_24875,N_24785);
nand U25298 (N_25298,N_24523,N_24992);
nor U25299 (N_25299,N_24913,N_24574);
nor U25300 (N_25300,N_24581,N_24779);
xnor U25301 (N_25301,N_24770,N_24568);
and U25302 (N_25302,N_24586,N_24926);
or U25303 (N_25303,N_24530,N_24889);
or U25304 (N_25304,N_24559,N_24544);
nand U25305 (N_25305,N_24883,N_24692);
or U25306 (N_25306,N_24689,N_24942);
xor U25307 (N_25307,N_24503,N_24555);
and U25308 (N_25308,N_24725,N_24984);
nand U25309 (N_25309,N_24643,N_24549);
xor U25310 (N_25310,N_24969,N_24539);
nor U25311 (N_25311,N_24709,N_24867);
nor U25312 (N_25312,N_24540,N_24562);
xor U25313 (N_25313,N_24997,N_24650);
nor U25314 (N_25314,N_24540,N_24693);
xor U25315 (N_25315,N_24621,N_24546);
or U25316 (N_25316,N_24777,N_24549);
xor U25317 (N_25317,N_24897,N_24652);
nand U25318 (N_25318,N_24973,N_24675);
and U25319 (N_25319,N_24592,N_24755);
nor U25320 (N_25320,N_24650,N_24818);
nor U25321 (N_25321,N_24972,N_24987);
nand U25322 (N_25322,N_24840,N_24856);
nand U25323 (N_25323,N_24603,N_24988);
nor U25324 (N_25324,N_24719,N_24513);
nor U25325 (N_25325,N_24758,N_24767);
or U25326 (N_25326,N_24994,N_24959);
nand U25327 (N_25327,N_24954,N_24925);
and U25328 (N_25328,N_24840,N_24594);
nand U25329 (N_25329,N_24673,N_24762);
and U25330 (N_25330,N_24777,N_24892);
or U25331 (N_25331,N_24876,N_24718);
xor U25332 (N_25332,N_24681,N_24973);
nor U25333 (N_25333,N_24837,N_24756);
and U25334 (N_25334,N_24513,N_24551);
or U25335 (N_25335,N_24947,N_24594);
nor U25336 (N_25336,N_24562,N_24605);
or U25337 (N_25337,N_24927,N_24714);
or U25338 (N_25338,N_24654,N_24687);
nor U25339 (N_25339,N_24649,N_24944);
or U25340 (N_25340,N_24543,N_24756);
nand U25341 (N_25341,N_24503,N_24554);
nor U25342 (N_25342,N_24841,N_24985);
or U25343 (N_25343,N_24945,N_24662);
and U25344 (N_25344,N_24656,N_24615);
and U25345 (N_25345,N_24755,N_24623);
nor U25346 (N_25346,N_24792,N_24815);
nor U25347 (N_25347,N_24972,N_24512);
and U25348 (N_25348,N_24938,N_24699);
and U25349 (N_25349,N_24611,N_24843);
xor U25350 (N_25350,N_24622,N_24812);
and U25351 (N_25351,N_24671,N_24602);
nor U25352 (N_25352,N_24846,N_24807);
nor U25353 (N_25353,N_24645,N_24571);
or U25354 (N_25354,N_24554,N_24884);
and U25355 (N_25355,N_24845,N_24982);
nor U25356 (N_25356,N_24888,N_24720);
or U25357 (N_25357,N_24761,N_24607);
nand U25358 (N_25358,N_24943,N_24660);
nand U25359 (N_25359,N_24602,N_24565);
nor U25360 (N_25360,N_24835,N_24946);
nor U25361 (N_25361,N_24755,N_24659);
and U25362 (N_25362,N_24644,N_24802);
or U25363 (N_25363,N_24889,N_24711);
or U25364 (N_25364,N_24711,N_24583);
nor U25365 (N_25365,N_24677,N_24652);
xnor U25366 (N_25366,N_24738,N_24825);
nor U25367 (N_25367,N_24965,N_24665);
or U25368 (N_25368,N_24878,N_24547);
xnor U25369 (N_25369,N_24899,N_24890);
xor U25370 (N_25370,N_24562,N_24903);
nor U25371 (N_25371,N_24626,N_24596);
nor U25372 (N_25372,N_24660,N_24559);
xnor U25373 (N_25373,N_24595,N_24534);
nand U25374 (N_25374,N_24536,N_24834);
and U25375 (N_25375,N_24629,N_24763);
and U25376 (N_25376,N_24565,N_24551);
or U25377 (N_25377,N_24619,N_24546);
nand U25378 (N_25378,N_24880,N_24780);
xnor U25379 (N_25379,N_24611,N_24673);
nor U25380 (N_25380,N_24503,N_24768);
or U25381 (N_25381,N_24781,N_24900);
xor U25382 (N_25382,N_24587,N_24777);
xor U25383 (N_25383,N_24967,N_24699);
nor U25384 (N_25384,N_24674,N_24543);
nor U25385 (N_25385,N_24894,N_24781);
or U25386 (N_25386,N_24615,N_24945);
nor U25387 (N_25387,N_24983,N_24781);
and U25388 (N_25388,N_24518,N_24758);
or U25389 (N_25389,N_24672,N_24737);
xor U25390 (N_25390,N_24874,N_24984);
nand U25391 (N_25391,N_24822,N_24847);
xnor U25392 (N_25392,N_24650,N_24736);
or U25393 (N_25393,N_24696,N_24914);
and U25394 (N_25394,N_24896,N_24946);
and U25395 (N_25395,N_24804,N_24599);
nand U25396 (N_25396,N_24671,N_24642);
nor U25397 (N_25397,N_24534,N_24746);
nand U25398 (N_25398,N_24935,N_24671);
and U25399 (N_25399,N_24689,N_24651);
and U25400 (N_25400,N_24967,N_24867);
nor U25401 (N_25401,N_24800,N_24594);
nor U25402 (N_25402,N_24779,N_24731);
nor U25403 (N_25403,N_24780,N_24727);
or U25404 (N_25404,N_24672,N_24947);
and U25405 (N_25405,N_24845,N_24914);
and U25406 (N_25406,N_24654,N_24698);
nand U25407 (N_25407,N_24856,N_24977);
nand U25408 (N_25408,N_24717,N_24722);
xnor U25409 (N_25409,N_24690,N_24785);
xor U25410 (N_25410,N_24583,N_24899);
nand U25411 (N_25411,N_24860,N_24522);
and U25412 (N_25412,N_24522,N_24576);
and U25413 (N_25413,N_24766,N_24966);
or U25414 (N_25414,N_24558,N_24913);
and U25415 (N_25415,N_24758,N_24813);
or U25416 (N_25416,N_24913,N_24896);
xnor U25417 (N_25417,N_24826,N_24929);
and U25418 (N_25418,N_24899,N_24931);
and U25419 (N_25419,N_24904,N_24686);
nor U25420 (N_25420,N_24721,N_24942);
and U25421 (N_25421,N_24638,N_24605);
or U25422 (N_25422,N_24857,N_24848);
nor U25423 (N_25423,N_24525,N_24744);
nand U25424 (N_25424,N_24814,N_24743);
and U25425 (N_25425,N_24559,N_24856);
or U25426 (N_25426,N_24835,N_24979);
nor U25427 (N_25427,N_24988,N_24974);
or U25428 (N_25428,N_24811,N_24972);
nor U25429 (N_25429,N_24916,N_24680);
nor U25430 (N_25430,N_24515,N_24527);
nor U25431 (N_25431,N_24883,N_24724);
nand U25432 (N_25432,N_24734,N_24661);
or U25433 (N_25433,N_24613,N_24563);
or U25434 (N_25434,N_24927,N_24629);
and U25435 (N_25435,N_24730,N_24889);
xor U25436 (N_25436,N_24519,N_24899);
nand U25437 (N_25437,N_24517,N_24659);
or U25438 (N_25438,N_24983,N_24795);
and U25439 (N_25439,N_24584,N_24672);
or U25440 (N_25440,N_24739,N_24672);
or U25441 (N_25441,N_24882,N_24831);
nand U25442 (N_25442,N_24728,N_24670);
nand U25443 (N_25443,N_24542,N_24721);
xnor U25444 (N_25444,N_24998,N_24960);
and U25445 (N_25445,N_24833,N_24979);
nand U25446 (N_25446,N_24906,N_24553);
nor U25447 (N_25447,N_24601,N_24834);
nand U25448 (N_25448,N_24818,N_24923);
nor U25449 (N_25449,N_24914,N_24910);
nor U25450 (N_25450,N_24563,N_24555);
xor U25451 (N_25451,N_24652,N_24710);
nor U25452 (N_25452,N_24743,N_24501);
and U25453 (N_25453,N_24855,N_24982);
and U25454 (N_25454,N_24568,N_24684);
nor U25455 (N_25455,N_24763,N_24994);
xnor U25456 (N_25456,N_24698,N_24894);
or U25457 (N_25457,N_24617,N_24780);
and U25458 (N_25458,N_24858,N_24765);
and U25459 (N_25459,N_24925,N_24846);
or U25460 (N_25460,N_24944,N_24784);
and U25461 (N_25461,N_24835,N_24632);
xor U25462 (N_25462,N_24954,N_24790);
nor U25463 (N_25463,N_24628,N_24545);
or U25464 (N_25464,N_24803,N_24658);
or U25465 (N_25465,N_24549,N_24555);
or U25466 (N_25466,N_24944,N_24995);
xnor U25467 (N_25467,N_24985,N_24528);
nor U25468 (N_25468,N_24791,N_24853);
xnor U25469 (N_25469,N_24911,N_24517);
nand U25470 (N_25470,N_24949,N_24965);
xnor U25471 (N_25471,N_24523,N_24568);
xnor U25472 (N_25472,N_24956,N_24999);
and U25473 (N_25473,N_24831,N_24644);
and U25474 (N_25474,N_24614,N_24568);
nor U25475 (N_25475,N_24517,N_24800);
xnor U25476 (N_25476,N_24950,N_24672);
nand U25477 (N_25477,N_24555,N_24558);
nand U25478 (N_25478,N_24827,N_24984);
and U25479 (N_25479,N_24934,N_24512);
xor U25480 (N_25480,N_24570,N_24774);
or U25481 (N_25481,N_24974,N_24975);
xor U25482 (N_25482,N_24966,N_24627);
xor U25483 (N_25483,N_24697,N_24727);
and U25484 (N_25484,N_24549,N_24973);
xnor U25485 (N_25485,N_24896,N_24897);
and U25486 (N_25486,N_24867,N_24729);
or U25487 (N_25487,N_24927,N_24690);
xor U25488 (N_25488,N_24934,N_24510);
or U25489 (N_25489,N_24653,N_24626);
xor U25490 (N_25490,N_24661,N_24768);
and U25491 (N_25491,N_24667,N_24973);
xor U25492 (N_25492,N_24766,N_24820);
nor U25493 (N_25493,N_24701,N_24971);
and U25494 (N_25494,N_24945,N_24913);
or U25495 (N_25495,N_24566,N_24848);
and U25496 (N_25496,N_24809,N_24822);
and U25497 (N_25497,N_24829,N_24628);
xnor U25498 (N_25498,N_24718,N_24715);
xnor U25499 (N_25499,N_24768,N_24771);
nor U25500 (N_25500,N_25275,N_25149);
nor U25501 (N_25501,N_25232,N_25058);
nand U25502 (N_25502,N_25363,N_25224);
or U25503 (N_25503,N_25338,N_25208);
or U25504 (N_25504,N_25432,N_25098);
and U25505 (N_25505,N_25274,N_25253);
and U25506 (N_25506,N_25166,N_25152);
nand U25507 (N_25507,N_25291,N_25334);
xor U25508 (N_25508,N_25294,N_25069);
nor U25509 (N_25509,N_25021,N_25056);
nor U25510 (N_25510,N_25127,N_25182);
xor U25511 (N_25511,N_25250,N_25313);
xnor U25512 (N_25512,N_25409,N_25336);
xnor U25513 (N_25513,N_25014,N_25266);
xor U25514 (N_25514,N_25062,N_25343);
or U25515 (N_25515,N_25327,N_25176);
nand U25516 (N_25516,N_25428,N_25395);
nor U25517 (N_25517,N_25196,N_25320);
nand U25518 (N_25518,N_25372,N_25205);
or U25519 (N_25519,N_25457,N_25197);
or U25520 (N_25520,N_25413,N_25431);
or U25521 (N_25521,N_25268,N_25163);
and U25522 (N_25522,N_25033,N_25333);
xor U25523 (N_25523,N_25020,N_25027);
nor U25524 (N_25524,N_25383,N_25341);
xor U25525 (N_25525,N_25499,N_25397);
and U25526 (N_25526,N_25416,N_25439);
nor U25527 (N_25527,N_25311,N_25482);
xnor U25528 (N_25528,N_25084,N_25335);
or U25529 (N_25529,N_25438,N_25353);
and U25530 (N_25530,N_25278,N_25337);
xnor U25531 (N_25531,N_25120,N_25324);
xor U25532 (N_25532,N_25272,N_25219);
and U25533 (N_25533,N_25296,N_25104);
and U25534 (N_25534,N_25032,N_25301);
xnor U25535 (N_25535,N_25436,N_25308);
or U25536 (N_25536,N_25287,N_25461);
and U25537 (N_25537,N_25466,N_25302);
nand U25538 (N_25538,N_25446,N_25183);
and U25539 (N_25539,N_25478,N_25361);
and U25540 (N_25540,N_25359,N_25379);
xor U25541 (N_25541,N_25158,N_25435);
nor U25542 (N_25542,N_25321,N_25083);
or U25543 (N_25543,N_25121,N_25244);
or U25544 (N_25544,N_25420,N_25112);
nand U25545 (N_25545,N_25329,N_25215);
xor U25546 (N_25546,N_25231,N_25087);
xor U25547 (N_25547,N_25270,N_25181);
xor U25548 (N_25548,N_25351,N_25011);
and U25549 (N_25549,N_25368,N_25095);
nor U25550 (N_25550,N_25229,N_25012);
and U25551 (N_25551,N_25496,N_25013);
nand U25552 (N_25552,N_25297,N_25404);
and U25553 (N_25553,N_25285,N_25491);
and U25554 (N_25554,N_25099,N_25042);
nor U25555 (N_25555,N_25249,N_25088);
nor U25556 (N_25556,N_25358,N_25079);
or U25557 (N_25557,N_25106,N_25396);
and U25558 (N_25558,N_25001,N_25154);
nor U25559 (N_25559,N_25109,N_25203);
and U25560 (N_25560,N_25248,N_25188);
nor U25561 (N_25561,N_25452,N_25177);
nor U25562 (N_25562,N_25004,N_25157);
nor U25563 (N_25563,N_25017,N_25172);
and U25564 (N_25564,N_25490,N_25091);
xor U25565 (N_25565,N_25290,N_25492);
nor U25566 (N_25566,N_25068,N_25373);
nand U25567 (N_25567,N_25450,N_25271);
or U25568 (N_25568,N_25073,N_25350);
xor U25569 (N_25569,N_25476,N_25443);
xor U25570 (N_25570,N_25155,N_25118);
xnor U25571 (N_25571,N_25414,N_25047);
and U25572 (N_25572,N_25059,N_25295);
nor U25573 (N_25573,N_25025,N_25424);
xor U25574 (N_25574,N_25200,N_25258);
and U25575 (N_25575,N_25259,N_25326);
or U25576 (N_25576,N_25293,N_25245);
or U25577 (N_25577,N_25470,N_25035);
nand U25578 (N_25578,N_25077,N_25340);
nand U25579 (N_25579,N_25356,N_25233);
nor U25580 (N_25580,N_25008,N_25473);
or U25581 (N_25581,N_25179,N_25137);
nor U25582 (N_25582,N_25255,N_25115);
xor U25583 (N_25583,N_25384,N_25110);
xnor U25584 (N_25584,N_25352,N_25078);
and U25585 (N_25585,N_25211,N_25016);
xor U25586 (N_25586,N_25434,N_25387);
nor U25587 (N_25587,N_25388,N_25116);
xor U25588 (N_25588,N_25031,N_25300);
and U25589 (N_25589,N_25497,N_25082);
and U25590 (N_25590,N_25355,N_25415);
xor U25591 (N_25591,N_25111,N_25080);
nor U25592 (N_25592,N_25280,N_25081);
xnor U25593 (N_25593,N_25173,N_25269);
nand U25594 (N_25594,N_25237,N_25003);
nand U25595 (N_25595,N_25403,N_25367);
xor U25596 (N_25596,N_25010,N_25184);
xor U25597 (N_25597,N_25440,N_25019);
nor U25598 (N_25598,N_25349,N_25228);
or U25599 (N_25599,N_25144,N_25417);
nand U25600 (N_25600,N_25150,N_25028);
xor U25601 (N_25601,N_25227,N_25433);
xnor U25602 (N_25602,N_25444,N_25314);
nor U25603 (N_25603,N_25456,N_25360);
xor U25604 (N_25604,N_25201,N_25463);
nor U25605 (N_25605,N_25283,N_25085);
and U25606 (N_25606,N_25277,N_25276);
nor U25607 (N_25607,N_25328,N_25138);
nor U25608 (N_25608,N_25427,N_25392);
xor U25609 (N_25609,N_25122,N_25286);
nor U25610 (N_25610,N_25223,N_25402);
nor U25611 (N_25611,N_25406,N_25041);
nor U25612 (N_25612,N_25312,N_25487);
nor U25613 (N_25613,N_25412,N_25169);
and U25614 (N_25614,N_25459,N_25040);
or U25615 (N_25615,N_25376,N_25257);
or U25616 (N_25616,N_25374,N_25391);
and U25617 (N_25617,N_25141,N_25394);
xor U25618 (N_25618,N_25030,N_25235);
and U25619 (N_25619,N_25213,N_25485);
nor U25620 (N_25620,N_25174,N_25053);
or U25621 (N_25621,N_25130,N_25316);
xnor U25622 (N_25622,N_25029,N_25217);
xnor U25623 (N_25623,N_25043,N_25400);
nor U25624 (N_25624,N_25153,N_25072);
or U25625 (N_25625,N_25486,N_25411);
xor U25626 (N_25626,N_25075,N_25451);
nand U25627 (N_25627,N_25124,N_25289);
nor U25628 (N_25628,N_25342,N_25045);
or U25629 (N_25629,N_25191,N_25419);
nor U25630 (N_25630,N_25362,N_25151);
nor U25631 (N_25631,N_25318,N_25454);
or U25632 (N_25632,N_25281,N_25306);
xor U25633 (N_25633,N_25418,N_25046);
or U25634 (N_25634,N_25061,N_25117);
nor U25635 (N_25635,N_25195,N_25023);
and U25636 (N_25636,N_25489,N_25168);
nor U25637 (N_25637,N_25243,N_25114);
and U25638 (N_25638,N_25242,N_25399);
xnor U25639 (N_25639,N_25364,N_25134);
and U25640 (N_25640,N_25322,N_25064);
or U25641 (N_25641,N_25299,N_25469);
nand U25642 (N_25642,N_25175,N_25164);
nor U25643 (N_25643,N_25209,N_25140);
nand U25644 (N_25644,N_25128,N_25048);
nor U25645 (N_25645,N_25238,N_25425);
nand U25646 (N_25646,N_25234,N_25484);
or U25647 (N_25647,N_25193,N_25323);
nand U25648 (N_25648,N_25194,N_25057);
or U25649 (N_25649,N_25465,N_25494);
xnor U25650 (N_25650,N_25246,N_25449);
xor U25651 (N_25651,N_25319,N_25462);
or U25652 (N_25652,N_25216,N_25074);
nor U25653 (N_25653,N_25273,N_25345);
or U25654 (N_25654,N_25307,N_25471);
xor U25655 (N_25655,N_25493,N_25050);
and U25656 (N_25656,N_25429,N_25292);
and U25657 (N_25657,N_25220,N_25024);
nor U25658 (N_25658,N_25288,N_25070);
or U25659 (N_25659,N_25148,N_25267);
xor U25660 (N_25660,N_25136,N_25309);
nand U25661 (N_25661,N_25051,N_25063);
and U25662 (N_25662,N_25198,N_25305);
nand U25663 (N_25663,N_25097,N_25065);
nor U25664 (N_25664,N_25093,N_25015);
or U25665 (N_25665,N_25284,N_25398);
xor U25666 (N_25666,N_25421,N_25026);
and U25667 (N_25667,N_25410,N_25139);
nand U25668 (N_25668,N_25039,N_25256);
xnor U25669 (N_25669,N_25365,N_25251);
xnor U25670 (N_25670,N_25007,N_25131);
nand U25671 (N_25671,N_25170,N_25441);
or U25672 (N_25672,N_25218,N_25192);
and U25673 (N_25673,N_25147,N_25422);
and U25674 (N_25674,N_25204,N_25430);
nor U25675 (N_25675,N_25472,N_25142);
or U25676 (N_25676,N_25480,N_25221);
or U25677 (N_25677,N_25185,N_25390);
nor U25678 (N_25678,N_25437,N_25036);
or U25679 (N_25679,N_25060,N_25371);
nor U25680 (N_25680,N_25145,N_25264);
nand U25681 (N_25681,N_25261,N_25006);
xnor U25682 (N_25682,N_25066,N_25389);
nand U25683 (N_25683,N_25222,N_25135);
or U25684 (N_25684,N_25018,N_25186);
or U25685 (N_25685,N_25347,N_25119);
xnor U25686 (N_25686,N_25442,N_25401);
or U25687 (N_25687,N_25005,N_25187);
or U25688 (N_25688,N_25094,N_25468);
nor U25689 (N_25689,N_25393,N_25160);
xnor U25690 (N_25690,N_25178,N_25100);
and U25691 (N_25691,N_25241,N_25202);
nand U25692 (N_25692,N_25113,N_25165);
nor U25693 (N_25693,N_25054,N_25348);
and U25694 (N_25694,N_25086,N_25126);
nor U25695 (N_25695,N_25447,N_25034);
nand U25696 (N_25696,N_25375,N_25146);
nand U25697 (N_25697,N_25252,N_25038);
or U25698 (N_25698,N_25156,N_25262);
or U25699 (N_25699,N_25380,N_25488);
or U25700 (N_25700,N_25423,N_25089);
xnor U25701 (N_25701,N_25239,N_25044);
xnor U25702 (N_25702,N_25049,N_25230);
and U25703 (N_25703,N_25199,N_25369);
xor U25704 (N_25704,N_25214,N_25386);
nand U25705 (N_25705,N_25055,N_25247);
and U25706 (N_25706,N_25096,N_25037);
and U25707 (N_25707,N_25180,N_25107);
or U25708 (N_25708,N_25167,N_25354);
or U25709 (N_25709,N_25240,N_25370);
xor U25710 (N_25710,N_25212,N_25236);
nor U25711 (N_25711,N_25458,N_25317);
and U25712 (N_25712,N_25002,N_25108);
and U25713 (N_25713,N_25298,N_25162);
xor U25714 (N_25714,N_25000,N_25448);
nand U25715 (N_25715,N_25445,N_25331);
xor U25716 (N_25716,N_25226,N_25263);
xor U25717 (N_25717,N_25310,N_25022);
nand U25718 (N_25718,N_25315,N_25123);
nor U25719 (N_25719,N_25426,N_25206);
xor U25720 (N_25720,N_25464,N_25133);
nor U25721 (N_25721,N_25132,N_25210);
nor U25722 (N_25722,N_25143,N_25159);
nor U25723 (N_25723,N_25125,N_25344);
nor U25724 (N_25724,N_25474,N_25103);
or U25725 (N_25725,N_25453,N_25357);
nand U25726 (N_25726,N_25381,N_25102);
or U25727 (N_25727,N_25455,N_25498);
xnor U25728 (N_25728,N_25304,N_25330);
and U25729 (N_25729,N_25408,N_25477);
xor U25730 (N_25730,N_25207,N_25101);
xnor U25731 (N_25731,N_25076,N_25339);
xor U25732 (N_25732,N_25325,N_25303);
or U25733 (N_25733,N_25366,N_25105);
xnor U25734 (N_25734,N_25377,N_25385);
nand U25735 (N_25735,N_25495,N_25279);
xor U25736 (N_25736,N_25479,N_25378);
or U25737 (N_25737,N_25483,N_25052);
or U25738 (N_25738,N_25171,N_25092);
or U25739 (N_25739,N_25332,N_25225);
and U25740 (N_25740,N_25254,N_25481);
and U25741 (N_25741,N_25265,N_25190);
xnor U25742 (N_25742,N_25071,N_25382);
nor U25743 (N_25743,N_25009,N_25189);
and U25744 (N_25744,N_25067,N_25460);
nand U25745 (N_25745,N_25090,N_25467);
xor U25746 (N_25746,N_25346,N_25407);
nor U25747 (N_25747,N_25405,N_25475);
nand U25748 (N_25748,N_25129,N_25282);
nor U25749 (N_25749,N_25260,N_25161);
nand U25750 (N_25750,N_25276,N_25239);
xnor U25751 (N_25751,N_25402,N_25423);
nand U25752 (N_25752,N_25013,N_25061);
nor U25753 (N_25753,N_25151,N_25293);
and U25754 (N_25754,N_25355,N_25169);
nand U25755 (N_25755,N_25198,N_25293);
nor U25756 (N_25756,N_25074,N_25200);
nor U25757 (N_25757,N_25339,N_25395);
and U25758 (N_25758,N_25173,N_25120);
xnor U25759 (N_25759,N_25151,N_25491);
xor U25760 (N_25760,N_25021,N_25302);
nand U25761 (N_25761,N_25218,N_25353);
nand U25762 (N_25762,N_25008,N_25069);
xnor U25763 (N_25763,N_25008,N_25351);
xnor U25764 (N_25764,N_25244,N_25407);
xor U25765 (N_25765,N_25275,N_25036);
or U25766 (N_25766,N_25047,N_25310);
nor U25767 (N_25767,N_25471,N_25198);
nand U25768 (N_25768,N_25258,N_25443);
or U25769 (N_25769,N_25185,N_25045);
nor U25770 (N_25770,N_25323,N_25085);
and U25771 (N_25771,N_25183,N_25447);
or U25772 (N_25772,N_25014,N_25295);
or U25773 (N_25773,N_25165,N_25027);
nor U25774 (N_25774,N_25003,N_25476);
or U25775 (N_25775,N_25389,N_25424);
or U25776 (N_25776,N_25244,N_25260);
xor U25777 (N_25777,N_25059,N_25200);
xnor U25778 (N_25778,N_25227,N_25317);
xnor U25779 (N_25779,N_25036,N_25074);
nor U25780 (N_25780,N_25186,N_25301);
and U25781 (N_25781,N_25459,N_25348);
nand U25782 (N_25782,N_25303,N_25474);
or U25783 (N_25783,N_25042,N_25310);
nand U25784 (N_25784,N_25109,N_25142);
nor U25785 (N_25785,N_25054,N_25200);
nand U25786 (N_25786,N_25365,N_25097);
or U25787 (N_25787,N_25392,N_25013);
nand U25788 (N_25788,N_25046,N_25008);
xnor U25789 (N_25789,N_25159,N_25146);
and U25790 (N_25790,N_25025,N_25169);
nand U25791 (N_25791,N_25479,N_25225);
nand U25792 (N_25792,N_25040,N_25038);
nor U25793 (N_25793,N_25441,N_25366);
and U25794 (N_25794,N_25322,N_25154);
nor U25795 (N_25795,N_25494,N_25400);
xor U25796 (N_25796,N_25267,N_25209);
nor U25797 (N_25797,N_25273,N_25371);
xnor U25798 (N_25798,N_25496,N_25040);
or U25799 (N_25799,N_25125,N_25416);
nor U25800 (N_25800,N_25229,N_25225);
nor U25801 (N_25801,N_25093,N_25404);
xnor U25802 (N_25802,N_25297,N_25491);
or U25803 (N_25803,N_25434,N_25222);
and U25804 (N_25804,N_25280,N_25367);
xor U25805 (N_25805,N_25402,N_25248);
or U25806 (N_25806,N_25083,N_25209);
nor U25807 (N_25807,N_25232,N_25403);
nor U25808 (N_25808,N_25044,N_25215);
or U25809 (N_25809,N_25028,N_25476);
xnor U25810 (N_25810,N_25174,N_25221);
xor U25811 (N_25811,N_25311,N_25361);
xnor U25812 (N_25812,N_25240,N_25252);
and U25813 (N_25813,N_25294,N_25257);
nand U25814 (N_25814,N_25475,N_25165);
xor U25815 (N_25815,N_25088,N_25311);
xor U25816 (N_25816,N_25198,N_25394);
nand U25817 (N_25817,N_25361,N_25417);
xor U25818 (N_25818,N_25251,N_25151);
or U25819 (N_25819,N_25442,N_25062);
xnor U25820 (N_25820,N_25056,N_25004);
nand U25821 (N_25821,N_25460,N_25321);
and U25822 (N_25822,N_25451,N_25400);
nand U25823 (N_25823,N_25008,N_25299);
nand U25824 (N_25824,N_25338,N_25323);
xor U25825 (N_25825,N_25266,N_25137);
nand U25826 (N_25826,N_25462,N_25316);
xor U25827 (N_25827,N_25222,N_25471);
nand U25828 (N_25828,N_25276,N_25063);
and U25829 (N_25829,N_25206,N_25367);
and U25830 (N_25830,N_25226,N_25293);
xnor U25831 (N_25831,N_25470,N_25392);
and U25832 (N_25832,N_25291,N_25498);
and U25833 (N_25833,N_25149,N_25249);
nor U25834 (N_25834,N_25386,N_25449);
or U25835 (N_25835,N_25193,N_25181);
nor U25836 (N_25836,N_25287,N_25104);
xnor U25837 (N_25837,N_25017,N_25336);
xnor U25838 (N_25838,N_25374,N_25191);
xnor U25839 (N_25839,N_25038,N_25407);
nor U25840 (N_25840,N_25410,N_25079);
nor U25841 (N_25841,N_25107,N_25485);
nor U25842 (N_25842,N_25180,N_25114);
nor U25843 (N_25843,N_25414,N_25231);
or U25844 (N_25844,N_25091,N_25075);
and U25845 (N_25845,N_25056,N_25081);
nor U25846 (N_25846,N_25467,N_25426);
xor U25847 (N_25847,N_25372,N_25333);
nand U25848 (N_25848,N_25171,N_25404);
xnor U25849 (N_25849,N_25128,N_25094);
nand U25850 (N_25850,N_25014,N_25325);
and U25851 (N_25851,N_25406,N_25286);
xnor U25852 (N_25852,N_25296,N_25183);
or U25853 (N_25853,N_25457,N_25191);
nor U25854 (N_25854,N_25046,N_25341);
nand U25855 (N_25855,N_25178,N_25446);
xor U25856 (N_25856,N_25198,N_25224);
and U25857 (N_25857,N_25201,N_25380);
nor U25858 (N_25858,N_25044,N_25312);
nor U25859 (N_25859,N_25112,N_25409);
xor U25860 (N_25860,N_25499,N_25330);
and U25861 (N_25861,N_25378,N_25028);
nand U25862 (N_25862,N_25159,N_25141);
xnor U25863 (N_25863,N_25141,N_25163);
xnor U25864 (N_25864,N_25027,N_25329);
xor U25865 (N_25865,N_25392,N_25094);
or U25866 (N_25866,N_25488,N_25308);
and U25867 (N_25867,N_25279,N_25292);
xnor U25868 (N_25868,N_25229,N_25196);
nor U25869 (N_25869,N_25118,N_25427);
or U25870 (N_25870,N_25319,N_25428);
nand U25871 (N_25871,N_25377,N_25093);
and U25872 (N_25872,N_25451,N_25263);
nand U25873 (N_25873,N_25041,N_25254);
nor U25874 (N_25874,N_25296,N_25011);
xor U25875 (N_25875,N_25237,N_25396);
nand U25876 (N_25876,N_25081,N_25368);
xnor U25877 (N_25877,N_25146,N_25294);
nand U25878 (N_25878,N_25083,N_25312);
nand U25879 (N_25879,N_25059,N_25397);
and U25880 (N_25880,N_25057,N_25261);
or U25881 (N_25881,N_25246,N_25430);
nand U25882 (N_25882,N_25094,N_25140);
nor U25883 (N_25883,N_25317,N_25258);
nor U25884 (N_25884,N_25016,N_25394);
or U25885 (N_25885,N_25493,N_25280);
nand U25886 (N_25886,N_25196,N_25016);
nor U25887 (N_25887,N_25060,N_25182);
or U25888 (N_25888,N_25301,N_25467);
xor U25889 (N_25889,N_25437,N_25329);
xor U25890 (N_25890,N_25066,N_25299);
nand U25891 (N_25891,N_25292,N_25164);
and U25892 (N_25892,N_25467,N_25049);
nor U25893 (N_25893,N_25399,N_25425);
and U25894 (N_25894,N_25001,N_25077);
nand U25895 (N_25895,N_25497,N_25313);
or U25896 (N_25896,N_25178,N_25474);
xor U25897 (N_25897,N_25327,N_25305);
or U25898 (N_25898,N_25103,N_25212);
nand U25899 (N_25899,N_25123,N_25324);
xor U25900 (N_25900,N_25395,N_25044);
nor U25901 (N_25901,N_25057,N_25426);
xnor U25902 (N_25902,N_25428,N_25077);
nand U25903 (N_25903,N_25078,N_25150);
nand U25904 (N_25904,N_25413,N_25425);
and U25905 (N_25905,N_25031,N_25009);
nor U25906 (N_25906,N_25413,N_25004);
xor U25907 (N_25907,N_25082,N_25345);
nor U25908 (N_25908,N_25471,N_25337);
xnor U25909 (N_25909,N_25101,N_25067);
or U25910 (N_25910,N_25218,N_25159);
nand U25911 (N_25911,N_25483,N_25034);
nand U25912 (N_25912,N_25391,N_25448);
or U25913 (N_25913,N_25299,N_25330);
nor U25914 (N_25914,N_25166,N_25083);
xor U25915 (N_25915,N_25277,N_25257);
xnor U25916 (N_25916,N_25205,N_25191);
nor U25917 (N_25917,N_25146,N_25075);
or U25918 (N_25918,N_25279,N_25111);
nor U25919 (N_25919,N_25015,N_25188);
nor U25920 (N_25920,N_25150,N_25221);
or U25921 (N_25921,N_25464,N_25331);
or U25922 (N_25922,N_25167,N_25172);
or U25923 (N_25923,N_25318,N_25336);
xnor U25924 (N_25924,N_25084,N_25067);
and U25925 (N_25925,N_25169,N_25138);
nand U25926 (N_25926,N_25163,N_25327);
nand U25927 (N_25927,N_25286,N_25444);
nor U25928 (N_25928,N_25099,N_25238);
xor U25929 (N_25929,N_25301,N_25323);
nor U25930 (N_25930,N_25474,N_25280);
nor U25931 (N_25931,N_25321,N_25489);
or U25932 (N_25932,N_25074,N_25102);
nand U25933 (N_25933,N_25323,N_25147);
and U25934 (N_25934,N_25171,N_25448);
nand U25935 (N_25935,N_25493,N_25266);
and U25936 (N_25936,N_25428,N_25479);
and U25937 (N_25937,N_25110,N_25117);
nand U25938 (N_25938,N_25000,N_25417);
xor U25939 (N_25939,N_25190,N_25141);
and U25940 (N_25940,N_25126,N_25375);
and U25941 (N_25941,N_25386,N_25064);
or U25942 (N_25942,N_25313,N_25477);
nor U25943 (N_25943,N_25062,N_25042);
xnor U25944 (N_25944,N_25407,N_25087);
or U25945 (N_25945,N_25445,N_25442);
and U25946 (N_25946,N_25148,N_25278);
and U25947 (N_25947,N_25306,N_25019);
and U25948 (N_25948,N_25338,N_25090);
xnor U25949 (N_25949,N_25242,N_25102);
or U25950 (N_25950,N_25409,N_25331);
xnor U25951 (N_25951,N_25353,N_25217);
nor U25952 (N_25952,N_25159,N_25069);
or U25953 (N_25953,N_25040,N_25177);
nor U25954 (N_25954,N_25346,N_25352);
or U25955 (N_25955,N_25137,N_25118);
xor U25956 (N_25956,N_25172,N_25297);
nand U25957 (N_25957,N_25430,N_25028);
and U25958 (N_25958,N_25204,N_25223);
nor U25959 (N_25959,N_25314,N_25244);
nor U25960 (N_25960,N_25013,N_25292);
and U25961 (N_25961,N_25390,N_25478);
and U25962 (N_25962,N_25284,N_25259);
or U25963 (N_25963,N_25258,N_25153);
xnor U25964 (N_25964,N_25179,N_25302);
and U25965 (N_25965,N_25429,N_25161);
nor U25966 (N_25966,N_25239,N_25455);
xor U25967 (N_25967,N_25235,N_25159);
xnor U25968 (N_25968,N_25064,N_25447);
and U25969 (N_25969,N_25320,N_25180);
and U25970 (N_25970,N_25399,N_25190);
nand U25971 (N_25971,N_25324,N_25140);
nor U25972 (N_25972,N_25413,N_25187);
or U25973 (N_25973,N_25021,N_25238);
and U25974 (N_25974,N_25029,N_25304);
nor U25975 (N_25975,N_25304,N_25065);
nor U25976 (N_25976,N_25032,N_25157);
nor U25977 (N_25977,N_25053,N_25055);
nor U25978 (N_25978,N_25439,N_25154);
xor U25979 (N_25979,N_25150,N_25098);
nor U25980 (N_25980,N_25424,N_25437);
or U25981 (N_25981,N_25418,N_25324);
nor U25982 (N_25982,N_25273,N_25012);
and U25983 (N_25983,N_25002,N_25070);
and U25984 (N_25984,N_25187,N_25225);
xnor U25985 (N_25985,N_25139,N_25053);
or U25986 (N_25986,N_25393,N_25267);
or U25987 (N_25987,N_25206,N_25352);
or U25988 (N_25988,N_25038,N_25479);
or U25989 (N_25989,N_25305,N_25087);
xnor U25990 (N_25990,N_25231,N_25353);
nand U25991 (N_25991,N_25275,N_25463);
and U25992 (N_25992,N_25492,N_25319);
or U25993 (N_25993,N_25419,N_25154);
and U25994 (N_25994,N_25437,N_25184);
and U25995 (N_25995,N_25359,N_25170);
nand U25996 (N_25996,N_25317,N_25342);
and U25997 (N_25997,N_25072,N_25122);
or U25998 (N_25998,N_25214,N_25437);
xor U25999 (N_25999,N_25281,N_25340);
and U26000 (N_26000,N_25948,N_25952);
and U26001 (N_26001,N_25938,N_25912);
nand U26002 (N_26002,N_25537,N_25949);
and U26003 (N_26003,N_25785,N_25675);
nor U26004 (N_26004,N_25554,N_25534);
xnor U26005 (N_26005,N_25842,N_25862);
or U26006 (N_26006,N_25997,N_25833);
and U26007 (N_26007,N_25893,N_25805);
xor U26008 (N_26008,N_25743,N_25991);
nor U26009 (N_26009,N_25593,N_25959);
xnor U26010 (N_26010,N_25695,N_25773);
nor U26011 (N_26011,N_25998,N_25643);
and U26012 (N_26012,N_25844,N_25741);
xnor U26013 (N_26013,N_25750,N_25798);
and U26014 (N_26014,N_25955,N_25781);
nand U26015 (N_26015,N_25792,N_25674);
and U26016 (N_26016,N_25899,N_25919);
and U26017 (N_26017,N_25562,N_25599);
or U26018 (N_26018,N_25777,N_25865);
xor U26019 (N_26019,N_25589,N_25552);
nor U26020 (N_26020,N_25506,N_25969);
and U26021 (N_26021,N_25718,N_25881);
nand U26022 (N_26022,N_25985,N_25983);
nand U26023 (N_26023,N_25924,N_25531);
nand U26024 (N_26024,N_25713,N_25760);
nand U26025 (N_26025,N_25986,N_25791);
nand U26026 (N_26026,N_25699,N_25730);
nor U26027 (N_26027,N_25512,N_25870);
nand U26028 (N_26028,N_25576,N_25793);
nand U26029 (N_26029,N_25610,N_25858);
nand U26030 (N_26030,N_25748,N_25503);
or U26031 (N_26031,N_25536,N_25529);
xnor U26032 (N_26032,N_25655,N_25634);
or U26033 (N_26033,N_25584,N_25764);
and U26034 (N_26034,N_25664,N_25992);
nor U26035 (N_26035,N_25692,N_25891);
or U26036 (N_26036,N_25690,N_25837);
nand U26037 (N_26037,N_25878,N_25974);
or U26038 (N_26038,N_25619,N_25659);
and U26039 (N_26039,N_25596,N_25590);
xor U26040 (N_26040,N_25587,N_25516);
or U26041 (N_26041,N_25775,N_25539);
nand U26042 (N_26042,N_25910,N_25981);
xnor U26043 (N_26043,N_25823,N_25830);
nand U26044 (N_26044,N_25687,N_25846);
nor U26045 (N_26045,N_25660,N_25567);
nor U26046 (N_26046,N_25714,N_25621);
nor U26047 (N_26047,N_25940,N_25917);
nand U26048 (N_26048,N_25519,N_25950);
xnor U26049 (N_26049,N_25918,N_25591);
nor U26050 (N_26050,N_25926,N_25831);
nand U26051 (N_26051,N_25538,N_25666);
nor U26052 (N_26052,N_25898,N_25696);
nor U26053 (N_26053,N_25670,N_25686);
nor U26054 (N_26054,N_25600,N_25657);
or U26055 (N_26055,N_25649,N_25560);
and U26056 (N_26056,N_25641,N_25611);
or U26057 (N_26057,N_25588,N_25819);
and U26058 (N_26058,N_25580,N_25638);
nand U26059 (N_26059,N_25731,N_25987);
nor U26060 (N_26060,N_25501,N_25715);
nand U26061 (N_26061,N_25541,N_25654);
nand U26062 (N_26062,N_25977,N_25559);
xor U26063 (N_26063,N_25960,N_25635);
or U26064 (N_26064,N_25756,N_25929);
xnor U26065 (N_26065,N_25671,N_25693);
or U26066 (N_26066,N_25704,N_25931);
xnor U26067 (N_26067,N_25609,N_25733);
nand U26068 (N_26068,N_25807,N_25863);
or U26069 (N_26069,N_25749,N_25639);
nand U26070 (N_26070,N_25520,N_25553);
xnor U26071 (N_26071,N_25789,N_25640);
nand U26072 (N_26072,N_25947,N_25669);
nor U26073 (N_26073,N_25927,N_25967);
nand U26074 (N_26074,N_25616,N_25770);
nor U26075 (N_26075,N_25943,N_25677);
or U26076 (N_26076,N_25975,N_25953);
and U26077 (N_26077,N_25883,N_25968);
nand U26078 (N_26078,N_25996,N_25629);
or U26079 (N_26079,N_25982,N_25822);
nand U26080 (N_26080,N_25941,N_25672);
nand U26081 (N_26081,N_25776,N_25916);
or U26082 (N_26082,N_25742,N_25701);
or U26083 (N_26083,N_25608,N_25993);
nand U26084 (N_26084,N_25800,N_25694);
nand U26085 (N_26085,N_25766,N_25772);
nand U26086 (N_26086,N_25737,N_25691);
nand U26087 (N_26087,N_25648,N_25874);
and U26088 (N_26088,N_25747,N_25835);
or U26089 (N_26089,N_25855,N_25966);
nand U26090 (N_26090,N_25888,N_25505);
and U26091 (N_26091,N_25542,N_25845);
and U26092 (N_26092,N_25627,N_25812);
nor U26093 (N_26093,N_25558,N_25951);
nor U26094 (N_26094,N_25540,N_25579);
or U26095 (N_26095,N_25905,N_25592);
nor U26096 (N_26096,N_25502,N_25736);
xnor U26097 (N_26097,N_25607,N_25852);
nand U26098 (N_26098,N_25757,N_25568);
or U26099 (N_26099,N_25957,N_25942);
or U26100 (N_26100,N_25828,N_25826);
nand U26101 (N_26101,N_25525,N_25707);
nand U26102 (N_26102,N_25684,N_25887);
nand U26103 (N_26103,N_25530,N_25988);
or U26104 (N_26104,N_25904,N_25962);
and U26105 (N_26105,N_25509,N_25720);
nand U26106 (N_26106,N_25682,N_25644);
and U26107 (N_26107,N_25866,N_25513);
nand U26108 (N_26108,N_25970,N_25615);
and U26109 (N_26109,N_25788,N_25504);
nand U26110 (N_26110,N_25827,N_25565);
nand U26111 (N_26111,N_25818,N_25532);
and U26112 (N_26112,N_25663,N_25645);
nand U26113 (N_26113,N_25685,N_25595);
nand U26114 (N_26114,N_25528,N_25774);
nor U26115 (N_26115,N_25892,N_25994);
or U26116 (N_26116,N_25586,N_25551);
or U26117 (N_26117,N_25566,N_25976);
and U26118 (N_26118,N_25581,N_25722);
and U26119 (N_26119,N_25879,N_25680);
xor U26120 (N_26120,N_25860,N_25763);
xor U26121 (N_26121,N_25518,N_25739);
xnor U26122 (N_26122,N_25799,N_25729);
nor U26123 (N_26123,N_25758,N_25932);
xnor U26124 (N_26124,N_25900,N_25508);
and U26125 (N_26125,N_25814,N_25698);
xnor U26126 (N_26126,N_25847,N_25582);
nor U26127 (N_26127,N_25618,N_25533);
nand U26128 (N_26128,N_25721,N_25761);
nand U26129 (N_26129,N_25626,N_25738);
xor U26130 (N_26130,N_25875,N_25903);
nor U26131 (N_26131,N_25880,N_25861);
xor U26132 (N_26132,N_25787,N_25995);
or U26133 (N_26133,N_25838,N_25703);
and U26134 (N_26134,N_25744,N_25771);
and U26135 (N_26135,N_25768,N_25765);
nor U26136 (N_26136,N_25697,N_25514);
xor U26137 (N_26137,N_25884,N_25662);
xor U26138 (N_26138,N_25575,N_25825);
and U26139 (N_26139,N_25856,N_25914);
nand U26140 (N_26140,N_25907,N_25719);
xor U26141 (N_26141,N_25762,N_25945);
nand U26142 (N_26142,N_25806,N_25623);
nor U26143 (N_26143,N_25734,N_25613);
nor U26144 (N_26144,N_25958,N_25755);
nand U26145 (N_26145,N_25939,N_25851);
xnor U26146 (N_26146,N_25859,N_25779);
xor U26147 (N_26147,N_25561,N_25889);
xor U26148 (N_26148,N_25711,N_25710);
or U26149 (N_26149,N_25809,N_25658);
nand U26150 (N_26150,N_25795,N_25622);
or U26151 (N_26151,N_25909,N_25667);
nand U26152 (N_26152,N_25548,N_25550);
or U26153 (N_26153,N_25676,N_25632);
xnor U26154 (N_26154,N_25740,N_25563);
nor U26155 (N_26155,N_25601,N_25767);
or U26156 (N_26156,N_25557,N_25937);
nor U26157 (N_26157,N_25813,N_25834);
or U26158 (N_26158,N_25523,N_25935);
or U26159 (N_26159,N_25746,N_25549);
nor U26160 (N_26160,N_25735,N_25517);
xnor U26161 (N_26161,N_25544,N_25728);
or U26162 (N_26162,N_25526,N_25522);
nand U26163 (N_26163,N_25804,N_25602);
nand U26164 (N_26164,N_25606,N_25630);
or U26165 (N_26165,N_25555,N_25612);
nand U26166 (N_26166,N_25751,N_25794);
xnor U26167 (N_26167,N_25702,N_25786);
or U26168 (N_26168,N_25527,N_25843);
nor U26169 (N_26169,N_25688,N_25979);
nor U26170 (N_26170,N_25896,N_25752);
nor U26171 (N_26171,N_25872,N_25535);
nand U26172 (N_26172,N_25871,N_25802);
and U26173 (N_26173,N_25727,N_25857);
nor U26174 (N_26174,N_25853,N_25936);
and U26175 (N_26175,N_25901,N_25642);
nor U26176 (N_26176,N_25574,N_25816);
and U26177 (N_26177,N_25628,N_25652);
or U26178 (N_26178,N_25647,N_25850);
nor U26179 (N_26179,N_25965,N_25913);
or U26180 (N_26180,N_25547,N_25753);
or U26181 (N_26181,N_25933,N_25679);
or U26182 (N_26182,N_25920,N_25716);
nand U26183 (N_26183,N_25815,N_25790);
nand U26184 (N_26184,N_25651,N_25821);
or U26185 (N_26185,N_25709,N_25820);
xnor U26186 (N_26186,N_25603,N_25832);
nor U26187 (N_26187,N_25546,N_25624);
or U26188 (N_26188,N_25572,N_25824);
nand U26189 (N_26189,N_25683,N_25614);
xor U26190 (N_26190,N_25759,N_25700);
or U26191 (N_26191,N_25836,N_25841);
xor U26192 (N_26192,N_25569,N_25978);
nor U26193 (N_26193,N_25573,N_25808);
nand U26194 (N_26194,N_25868,N_25922);
xor U26195 (N_26195,N_25543,N_25902);
or U26196 (N_26196,N_25817,N_25732);
nor U26197 (N_26197,N_25869,N_25625);
nor U26198 (N_26198,N_25811,N_25964);
nor U26199 (N_26199,N_25784,N_25726);
xnor U26200 (N_26200,N_25944,N_25915);
nor U26201 (N_26201,N_25882,N_25597);
nor U26202 (N_26202,N_25585,N_25778);
and U26203 (N_26203,N_25571,N_25673);
and U26204 (N_26204,N_25797,N_25877);
and U26205 (N_26205,N_25849,N_25810);
and U26206 (N_26206,N_25656,N_25653);
nor U26207 (N_26207,N_25973,N_25801);
and U26208 (N_26208,N_25908,N_25854);
nand U26209 (N_26209,N_25598,N_25921);
nand U26210 (N_26210,N_25930,N_25956);
nand U26211 (N_26211,N_25745,N_25990);
nand U26212 (N_26212,N_25620,N_25705);
or U26213 (N_26213,N_25999,N_25681);
or U26214 (N_26214,N_25928,N_25646);
nand U26215 (N_26215,N_25594,N_25724);
xor U26216 (N_26216,N_25840,N_25500);
or U26217 (N_26217,N_25507,N_25617);
and U26218 (N_26218,N_25524,N_25564);
or U26219 (N_26219,N_25848,N_25971);
nand U26220 (N_26220,N_25954,N_25712);
and U26221 (N_26221,N_25665,N_25890);
or U26222 (N_26222,N_25980,N_25637);
nor U26223 (N_26223,N_25708,N_25583);
nand U26224 (N_26224,N_25578,N_25897);
nor U26225 (N_26225,N_25864,N_25961);
nor U26226 (N_26226,N_25782,N_25911);
nand U26227 (N_26227,N_25989,N_25556);
or U26228 (N_26228,N_25650,N_25631);
nand U26229 (N_26229,N_25570,N_25605);
nor U26230 (N_26230,N_25604,N_25725);
and U26231 (N_26231,N_25689,N_25633);
and U26232 (N_26232,N_25515,N_25963);
nand U26233 (N_26233,N_25876,N_25867);
nor U26234 (N_26234,N_25661,N_25803);
nand U26235 (N_26235,N_25668,N_25636);
xor U26236 (N_26236,N_25906,N_25895);
and U26237 (N_26237,N_25946,N_25885);
or U26238 (N_26238,N_25545,N_25706);
nor U26239 (N_26239,N_25717,N_25886);
xnor U26240 (N_26240,N_25769,N_25796);
nor U26241 (N_26241,N_25510,N_25723);
and U26242 (N_26242,N_25925,N_25984);
xnor U26243 (N_26243,N_25678,N_25829);
nand U26244 (N_26244,N_25923,N_25577);
and U26245 (N_26245,N_25511,N_25934);
xnor U26246 (N_26246,N_25754,N_25780);
or U26247 (N_26247,N_25972,N_25873);
and U26248 (N_26248,N_25839,N_25894);
and U26249 (N_26249,N_25521,N_25783);
and U26250 (N_26250,N_25918,N_25609);
or U26251 (N_26251,N_25699,N_25683);
xor U26252 (N_26252,N_25645,N_25561);
and U26253 (N_26253,N_25629,N_25736);
nor U26254 (N_26254,N_25963,N_25716);
xor U26255 (N_26255,N_25866,N_25511);
or U26256 (N_26256,N_25928,N_25992);
nor U26257 (N_26257,N_25962,N_25759);
nand U26258 (N_26258,N_25723,N_25555);
or U26259 (N_26259,N_25548,N_25751);
and U26260 (N_26260,N_25688,N_25984);
nor U26261 (N_26261,N_25625,N_25663);
nor U26262 (N_26262,N_25994,N_25700);
nand U26263 (N_26263,N_25975,N_25826);
or U26264 (N_26264,N_25922,N_25979);
and U26265 (N_26265,N_25507,N_25565);
nand U26266 (N_26266,N_25897,N_25562);
xnor U26267 (N_26267,N_25613,N_25516);
and U26268 (N_26268,N_25707,N_25548);
nor U26269 (N_26269,N_25613,N_25779);
and U26270 (N_26270,N_25557,N_25757);
nor U26271 (N_26271,N_25772,N_25508);
xnor U26272 (N_26272,N_25882,N_25592);
and U26273 (N_26273,N_25849,N_25758);
and U26274 (N_26274,N_25913,N_25904);
or U26275 (N_26275,N_25764,N_25674);
xnor U26276 (N_26276,N_25833,N_25615);
nand U26277 (N_26277,N_25555,N_25725);
or U26278 (N_26278,N_25629,N_25583);
and U26279 (N_26279,N_25825,N_25596);
or U26280 (N_26280,N_25969,N_25670);
or U26281 (N_26281,N_25546,N_25784);
nor U26282 (N_26282,N_25562,N_25641);
or U26283 (N_26283,N_25863,N_25959);
nor U26284 (N_26284,N_25725,N_25818);
nor U26285 (N_26285,N_25791,N_25571);
xnor U26286 (N_26286,N_25575,N_25817);
or U26287 (N_26287,N_25529,N_25828);
or U26288 (N_26288,N_25734,N_25580);
or U26289 (N_26289,N_25858,N_25806);
and U26290 (N_26290,N_25804,N_25998);
and U26291 (N_26291,N_25671,N_25933);
xor U26292 (N_26292,N_25621,N_25701);
or U26293 (N_26293,N_25967,N_25768);
xnor U26294 (N_26294,N_25642,N_25947);
xor U26295 (N_26295,N_25920,N_25646);
and U26296 (N_26296,N_25531,N_25662);
or U26297 (N_26297,N_25814,N_25707);
nand U26298 (N_26298,N_25699,N_25907);
nand U26299 (N_26299,N_25558,N_25542);
and U26300 (N_26300,N_25786,N_25648);
and U26301 (N_26301,N_25710,N_25503);
and U26302 (N_26302,N_25636,N_25865);
or U26303 (N_26303,N_25686,N_25904);
nand U26304 (N_26304,N_25943,N_25740);
nand U26305 (N_26305,N_25580,N_25823);
xnor U26306 (N_26306,N_25946,N_25861);
nor U26307 (N_26307,N_25625,N_25987);
xor U26308 (N_26308,N_25747,N_25766);
nor U26309 (N_26309,N_25971,N_25749);
or U26310 (N_26310,N_25849,N_25771);
and U26311 (N_26311,N_25995,N_25838);
and U26312 (N_26312,N_25890,N_25895);
nand U26313 (N_26313,N_25967,N_25668);
or U26314 (N_26314,N_25600,N_25824);
and U26315 (N_26315,N_25749,N_25836);
or U26316 (N_26316,N_25526,N_25713);
xnor U26317 (N_26317,N_25789,N_25544);
nor U26318 (N_26318,N_25839,N_25609);
nor U26319 (N_26319,N_25514,N_25528);
or U26320 (N_26320,N_25821,N_25696);
or U26321 (N_26321,N_25678,N_25666);
and U26322 (N_26322,N_25805,N_25500);
or U26323 (N_26323,N_25677,N_25820);
nor U26324 (N_26324,N_25731,N_25760);
or U26325 (N_26325,N_25809,N_25912);
or U26326 (N_26326,N_25643,N_25544);
nand U26327 (N_26327,N_25965,N_25505);
nor U26328 (N_26328,N_25644,N_25620);
or U26329 (N_26329,N_25865,N_25736);
nor U26330 (N_26330,N_25877,N_25749);
and U26331 (N_26331,N_25949,N_25963);
nor U26332 (N_26332,N_25585,N_25527);
or U26333 (N_26333,N_25899,N_25868);
nand U26334 (N_26334,N_25777,N_25711);
or U26335 (N_26335,N_25566,N_25991);
or U26336 (N_26336,N_25880,N_25728);
and U26337 (N_26337,N_25562,N_25684);
and U26338 (N_26338,N_25680,N_25671);
nand U26339 (N_26339,N_25914,N_25753);
nand U26340 (N_26340,N_25639,N_25908);
and U26341 (N_26341,N_25947,N_25935);
and U26342 (N_26342,N_25536,N_25698);
xnor U26343 (N_26343,N_25502,N_25551);
and U26344 (N_26344,N_25544,N_25890);
and U26345 (N_26345,N_25788,N_25779);
or U26346 (N_26346,N_25601,N_25965);
or U26347 (N_26347,N_25801,N_25717);
or U26348 (N_26348,N_25970,N_25755);
nand U26349 (N_26349,N_25720,N_25999);
nor U26350 (N_26350,N_25614,N_25823);
or U26351 (N_26351,N_25698,N_25662);
nand U26352 (N_26352,N_25966,N_25935);
nor U26353 (N_26353,N_25841,N_25587);
nor U26354 (N_26354,N_25897,N_25661);
or U26355 (N_26355,N_25684,N_25899);
or U26356 (N_26356,N_25684,N_25694);
and U26357 (N_26357,N_25532,N_25839);
nor U26358 (N_26358,N_25580,N_25627);
and U26359 (N_26359,N_25585,N_25895);
and U26360 (N_26360,N_25697,N_25929);
or U26361 (N_26361,N_25883,N_25850);
nor U26362 (N_26362,N_25555,N_25643);
nor U26363 (N_26363,N_25514,N_25548);
or U26364 (N_26364,N_25579,N_25827);
and U26365 (N_26365,N_25731,N_25732);
nor U26366 (N_26366,N_25751,N_25666);
xor U26367 (N_26367,N_25606,N_25880);
xor U26368 (N_26368,N_25792,N_25775);
or U26369 (N_26369,N_25816,N_25639);
nand U26370 (N_26370,N_25605,N_25516);
or U26371 (N_26371,N_25953,N_25664);
nand U26372 (N_26372,N_25543,N_25771);
nor U26373 (N_26373,N_25513,N_25505);
nor U26374 (N_26374,N_25963,N_25674);
nor U26375 (N_26375,N_25866,N_25936);
or U26376 (N_26376,N_25701,N_25881);
xor U26377 (N_26377,N_25978,N_25689);
nand U26378 (N_26378,N_25934,N_25533);
and U26379 (N_26379,N_25803,N_25754);
nand U26380 (N_26380,N_25747,N_25561);
xnor U26381 (N_26381,N_25766,N_25545);
or U26382 (N_26382,N_25593,N_25767);
nand U26383 (N_26383,N_25536,N_25981);
nand U26384 (N_26384,N_25855,N_25989);
nor U26385 (N_26385,N_25930,N_25684);
or U26386 (N_26386,N_25537,N_25715);
and U26387 (N_26387,N_25960,N_25584);
nor U26388 (N_26388,N_25587,N_25802);
and U26389 (N_26389,N_25603,N_25543);
or U26390 (N_26390,N_25563,N_25897);
and U26391 (N_26391,N_25823,N_25592);
nor U26392 (N_26392,N_25707,N_25901);
and U26393 (N_26393,N_25963,N_25927);
and U26394 (N_26394,N_25666,N_25599);
and U26395 (N_26395,N_25634,N_25625);
xnor U26396 (N_26396,N_25644,N_25870);
nand U26397 (N_26397,N_25559,N_25951);
nand U26398 (N_26398,N_25830,N_25638);
and U26399 (N_26399,N_25947,N_25581);
nor U26400 (N_26400,N_25877,N_25520);
nand U26401 (N_26401,N_25839,N_25746);
nor U26402 (N_26402,N_25797,N_25573);
nand U26403 (N_26403,N_25771,N_25911);
nor U26404 (N_26404,N_25512,N_25609);
nand U26405 (N_26405,N_25624,N_25741);
xnor U26406 (N_26406,N_25525,N_25522);
nand U26407 (N_26407,N_25851,N_25572);
xnor U26408 (N_26408,N_25984,N_25625);
or U26409 (N_26409,N_25735,N_25522);
or U26410 (N_26410,N_25608,N_25714);
nor U26411 (N_26411,N_25551,N_25689);
and U26412 (N_26412,N_25828,N_25701);
or U26413 (N_26413,N_25653,N_25736);
xor U26414 (N_26414,N_25569,N_25737);
nand U26415 (N_26415,N_25928,N_25521);
nor U26416 (N_26416,N_25683,N_25936);
nor U26417 (N_26417,N_25670,N_25906);
nor U26418 (N_26418,N_25722,N_25656);
nand U26419 (N_26419,N_25528,N_25867);
nand U26420 (N_26420,N_25765,N_25537);
xor U26421 (N_26421,N_25905,N_25675);
or U26422 (N_26422,N_25863,N_25528);
nor U26423 (N_26423,N_25714,N_25541);
and U26424 (N_26424,N_25936,N_25727);
and U26425 (N_26425,N_25515,N_25748);
or U26426 (N_26426,N_25829,N_25584);
nand U26427 (N_26427,N_25560,N_25675);
nor U26428 (N_26428,N_25992,N_25891);
nand U26429 (N_26429,N_25560,N_25693);
xor U26430 (N_26430,N_25778,N_25640);
nand U26431 (N_26431,N_25841,N_25768);
nand U26432 (N_26432,N_25996,N_25690);
xor U26433 (N_26433,N_25792,N_25598);
and U26434 (N_26434,N_25920,N_25806);
or U26435 (N_26435,N_25808,N_25903);
or U26436 (N_26436,N_25925,N_25789);
nand U26437 (N_26437,N_25687,N_25566);
nand U26438 (N_26438,N_25608,N_25542);
nor U26439 (N_26439,N_25628,N_25830);
nor U26440 (N_26440,N_25527,N_25591);
nor U26441 (N_26441,N_25799,N_25903);
nand U26442 (N_26442,N_25652,N_25526);
and U26443 (N_26443,N_25525,N_25620);
nor U26444 (N_26444,N_25832,N_25675);
or U26445 (N_26445,N_25851,N_25666);
or U26446 (N_26446,N_25949,N_25894);
xnor U26447 (N_26447,N_25659,N_25934);
or U26448 (N_26448,N_25883,N_25568);
xnor U26449 (N_26449,N_25726,N_25754);
and U26450 (N_26450,N_25694,N_25626);
nand U26451 (N_26451,N_25744,N_25999);
nand U26452 (N_26452,N_25595,N_25713);
nand U26453 (N_26453,N_25920,N_25647);
nand U26454 (N_26454,N_25942,N_25823);
xnor U26455 (N_26455,N_25559,N_25772);
nand U26456 (N_26456,N_25560,N_25860);
nand U26457 (N_26457,N_25843,N_25531);
xnor U26458 (N_26458,N_25919,N_25680);
xnor U26459 (N_26459,N_25650,N_25717);
or U26460 (N_26460,N_25795,N_25732);
or U26461 (N_26461,N_25682,N_25788);
xnor U26462 (N_26462,N_25652,N_25551);
and U26463 (N_26463,N_25858,N_25795);
or U26464 (N_26464,N_25567,N_25988);
nor U26465 (N_26465,N_25976,N_25951);
and U26466 (N_26466,N_25731,N_25868);
xnor U26467 (N_26467,N_25840,N_25780);
and U26468 (N_26468,N_25719,N_25944);
or U26469 (N_26469,N_25599,N_25991);
xnor U26470 (N_26470,N_25504,N_25774);
nand U26471 (N_26471,N_25545,N_25986);
or U26472 (N_26472,N_25819,N_25897);
nor U26473 (N_26473,N_25697,N_25843);
nor U26474 (N_26474,N_25582,N_25923);
nand U26475 (N_26475,N_25606,N_25919);
xnor U26476 (N_26476,N_25781,N_25573);
nand U26477 (N_26477,N_25622,N_25767);
nor U26478 (N_26478,N_25661,N_25619);
and U26479 (N_26479,N_25833,N_25622);
and U26480 (N_26480,N_25911,N_25899);
nor U26481 (N_26481,N_25923,N_25912);
xor U26482 (N_26482,N_25986,N_25719);
xnor U26483 (N_26483,N_25986,N_25525);
nand U26484 (N_26484,N_25688,N_25637);
xor U26485 (N_26485,N_25817,N_25506);
nand U26486 (N_26486,N_25984,N_25963);
nand U26487 (N_26487,N_25635,N_25985);
nor U26488 (N_26488,N_25501,N_25921);
xor U26489 (N_26489,N_25843,N_25659);
or U26490 (N_26490,N_25521,N_25920);
nand U26491 (N_26491,N_25968,N_25554);
xor U26492 (N_26492,N_25626,N_25955);
xnor U26493 (N_26493,N_25933,N_25718);
nand U26494 (N_26494,N_25767,N_25910);
or U26495 (N_26495,N_25932,N_25811);
and U26496 (N_26496,N_25767,N_25674);
nor U26497 (N_26497,N_25923,N_25706);
nand U26498 (N_26498,N_25583,N_25632);
nor U26499 (N_26499,N_25949,N_25778);
nand U26500 (N_26500,N_26227,N_26474);
or U26501 (N_26501,N_26267,N_26386);
nand U26502 (N_26502,N_26122,N_26337);
and U26503 (N_26503,N_26248,N_26446);
nor U26504 (N_26504,N_26418,N_26426);
and U26505 (N_26505,N_26177,N_26154);
xnor U26506 (N_26506,N_26074,N_26489);
nor U26507 (N_26507,N_26187,N_26445);
and U26508 (N_26508,N_26200,N_26109);
or U26509 (N_26509,N_26053,N_26308);
or U26510 (N_26510,N_26498,N_26012);
xnor U26511 (N_26511,N_26338,N_26303);
nor U26512 (N_26512,N_26018,N_26421);
or U26513 (N_26513,N_26372,N_26313);
nor U26514 (N_26514,N_26243,N_26234);
and U26515 (N_26515,N_26136,N_26052);
nand U26516 (N_26516,N_26441,N_26230);
xor U26517 (N_26517,N_26417,N_26468);
nor U26518 (N_26518,N_26183,N_26249);
or U26519 (N_26519,N_26013,N_26022);
xnor U26520 (N_26520,N_26209,N_26063);
and U26521 (N_26521,N_26170,N_26166);
or U26522 (N_26522,N_26329,N_26112);
and U26523 (N_26523,N_26028,N_26151);
xor U26524 (N_26524,N_26195,N_26036);
nand U26525 (N_26525,N_26153,N_26162);
nor U26526 (N_26526,N_26127,N_26078);
xnor U26527 (N_26527,N_26402,N_26497);
xnor U26528 (N_26528,N_26116,N_26269);
or U26529 (N_26529,N_26044,N_26469);
and U26530 (N_26530,N_26293,N_26020);
xor U26531 (N_26531,N_26440,N_26281);
nand U26532 (N_26532,N_26451,N_26081);
nor U26533 (N_26533,N_26365,N_26431);
nand U26534 (N_26534,N_26133,N_26339);
or U26535 (N_26535,N_26367,N_26168);
and U26536 (N_26536,N_26141,N_26150);
nand U26537 (N_26537,N_26377,N_26235);
or U26538 (N_26538,N_26327,N_26427);
xnor U26539 (N_26539,N_26488,N_26123);
xnor U26540 (N_26540,N_26246,N_26399);
xnor U26541 (N_26541,N_26194,N_26450);
nor U26542 (N_26542,N_26341,N_26438);
and U26543 (N_26543,N_26185,N_26199);
xnor U26544 (N_26544,N_26499,N_26077);
nand U26545 (N_26545,N_26137,N_26031);
nand U26546 (N_26546,N_26307,N_26138);
and U26547 (N_26547,N_26203,N_26458);
nor U26548 (N_26548,N_26090,N_26467);
nor U26549 (N_26549,N_26059,N_26221);
or U26550 (N_26550,N_26041,N_26094);
nand U26551 (N_26551,N_26494,N_26482);
xnor U26552 (N_26552,N_26272,N_26120);
nor U26553 (N_26553,N_26315,N_26364);
or U26554 (N_26554,N_26486,N_26299);
nor U26555 (N_26555,N_26210,N_26321);
xnor U26556 (N_26556,N_26245,N_26001);
xor U26557 (N_26557,N_26155,N_26111);
xnor U26558 (N_26558,N_26023,N_26092);
or U26559 (N_26559,N_26217,N_26057);
and U26560 (N_26560,N_26147,N_26007);
and U26561 (N_26561,N_26232,N_26447);
and U26562 (N_26562,N_26056,N_26065);
and U26563 (N_26563,N_26256,N_26385);
or U26564 (N_26564,N_26320,N_26045);
nand U26565 (N_26565,N_26176,N_26242);
or U26566 (N_26566,N_26197,N_26084);
or U26567 (N_26567,N_26139,N_26182);
nor U26568 (N_26568,N_26424,N_26351);
nor U26569 (N_26569,N_26282,N_26072);
xnor U26570 (N_26570,N_26250,N_26205);
or U26571 (N_26571,N_26449,N_26161);
nor U26572 (N_26572,N_26129,N_26042);
or U26573 (N_26573,N_26263,N_26134);
or U26574 (N_26574,N_26037,N_26485);
and U26575 (N_26575,N_26244,N_26291);
nand U26576 (N_26576,N_26214,N_26058);
or U26577 (N_26577,N_26083,N_26419);
or U26578 (N_26578,N_26333,N_26328);
nand U26579 (N_26579,N_26389,N_26379);
or U26580 (N_26580,N_26460,N_26107);
nand U26581 (N_26581,N_26215,N_26343);
and U26582 (N_26582,N_26146,N_26103);
xnor U26583 (N_26583,N_26238,N_26340);
and U26584 (N_26584,N_26411,N_26240);
or U26585 (N_26585,N_26317,N_26278);
or U26586 (N_26586,N_26096,N_26026);
or U26587 (N_26587,N_26178,N_26079);
xor U26588 (N_26588,N_26357,N_26247);
nand U26589 (N_26589,N_26376,N_26188);
or U26590 (N_26590,N_26491,N_26294);
or U26591 (N_26591,N_26190,N_26346);
nor U26592 (N_26592,N_26066,N_26252);
or U26593 (N_26593,N_26395,N_26382);
or U26594 (N_26594,N_26019,N_26212);
and U26595 (N_26595,N_26164,N_26229);
and U26596 (N_26596,N_26470,N_26452);
nand U26597 (N_26597,N_26492,N_26284);
xnor U26598 (N_26598,N_26462,N_26405);
nor U26599 (N_26599,N_26276,N_26118);
xor U26600 (N_26600,N_26442,N_26220);
nand U26601 (N_26601,N_26265,N_26101);
nand U26602 (N_26602,N_26306,N_26174);
nand U26603 (N_26603,N_26145,N_26415);
nand U26604 (N_26604,N_26152,N_26061);
or U26605 (N_26605,N_26075,N_26222);
nand U26606 (N_26606,N_26040,N_26132);
xnor U26607 (N_26607,N_26160,N_26029);
nor U26608 (N_26608,N_26261,N_26448);
xor U26609 (N_26609,N_26373,N_26172);
nor U26610 (N_26610,N_26398,N_26125);
and U26611 (N_26611,N_26097,N_26300);
and U26612 (N_26612,N_26196,N_26356);
xor U26613 (N_26613,N_26404,N_26480);
and U26614 (N_26614,N_26297,N_26102);
nand U26615 (N_26615,N_26105,N_26224);
and U26616 (N_26616,N_26021,N_26016);
and U26617 (N_26617,N_26010,N_26384);
nand U26618 (N_26618,N_26331,N_26143);
nor U26619 (N_26619,N_26428,N_26050);
and U26620 (N_26620,N_26406,N_26085);
or U26621 (N_26621,N_26330,N_26298);
nand U26622 (N_26622,N_26192,N_26181);
and U26623 (N_26623,N_26032,N_26180);
nor U26624 (N_26624,N_26124,N_26251);
nand U26625 (N_26625,N_26173,N_26275);
and U26626 (N_26626,N_26347,N_26439);
and U26627 (N_26627,N_26381,N_26457);
nor U26628 (N_26628,N_26011,N_26416);
and U26629 (N_26629,N_26008,N_26412);
nand U26630 (N_26630,N_26309,N_26495);
nor U26631 (N_26631,N_26403,N_26374);
xnor U26632 (N_26632,N_26466,N_26473);
xnor U26633 (N_26633,N_26068,N_26004);
or U26634 (N_26634,N_26332,N_26336);
and U26635 (N_26635,N_26271,N_26355);
or U26636 (N_26636,N_26034,N_26342);
and U26637 (N_26637,N_26167,N_26024);
xor U26638 (N_26638,N_26359,N_26100);
xor U26639 (N_26639,N_26131,N_26312);
and U26640 (N_26640,N_26006,N_26208);
nand U26641 (N_26641,N_26481,N_26454);
nor U26642 (N_26642,N_26163,N_26483);
or U26643 (N_26643,N_26099,N_26310);
or U26644 (N_26644,N_26360,N_26391);
xor U26645 (N_26645,N_26237,N_26390);
and U26646 (N_26646,N_26005,N_26064);
nor U26647 (N_26647,N_26002,N_26430);
and U26648 (N_26648,N_26423,N_26225);
and U26649 (N_26649,N_26350,N_26219);
and U26650 (N_26650,N_26463,N_26130);
or U26651 (N_26651,N_26396,N_26361);
and U26652 (N_26652,N_26236,N_26478);
and U26653 (N_26653,N_26165,N_26128);
nor U26654 (N_26654,N_26477,N_26273);
xnor U26655 (N_26655,N_26104,N_26098);
nand U26656 (N_26656,N_26397,N_26257);
or U26657 (N_26657,N_26475,N_26290);
nor U26658 (N_26658,N_26093,N_26302);
and U26659 (N_26659,N_26318,N_26211);
nor U26660 (N_26660,N_26201,N_26060);
nand U26661 (N_26661,N_26326,N_26432);
nor U26662 (N_26662,N_26392,N_26435);
and U26663 (N_26663,N_26323,N_26345);
nand U26664 (N_26664,N_26285,N_26433);
or U26665 (N_26665,N_26465,N_26144);
and U26666 (N_26666,N_26216,N_26493);
xnor U26667 (N_26667,N_26264,N_26091);
xor U26668 (N_26668,N_26363,N_26035);
and U26669 (N_26669,N_26292,N_26086);
or U26670 (N_26670,N_26443,N_26179);
xnor U26671 (N_26671,N_26259,N_26378);
xnor U26672 (N_26672,N_26082,N_26262);
and U26673 (N_26673,N_26456,N_26400);
and U26674 (N_26674,N_26157,N_26113);
xor U26675 (N_26675,N_26121,N_26429);
or U26676 (N_26676,N_26142,N_26258);
xnor U26677 (N_26677,N_26095,N_26241);
xnor U26678 (N_26678,N_26476,N_26087);
and U26679 (N_26679,N_26191,N_26062);
and U26680 (N_26680,N_26254,N_26039);
nor U26681 (N_26681,N_26268,N_26410);
xnor U26682 (N_26682,N_26015,N_26231);
and U26683 (N_26683,N_26159,N_26049);
or U26684 (N_26684,N_26393,N_26335);
xnor U26685 (N_26685,N_26289,N_26228);
nand U26686 (N_26686,N_26316,N_26204);
xnor U26687 (N_26687,N_26067,N_26171);
xnor U26688 (N_26688,N_26288,N_26461);
or U26689 (N_26689,N_26000,N_26175);
and U26690 (N_26690,N_26088,N_26149);
nor U26691 (N_26691,N_26354,N_26114);
xnor U26692 (N_26692,N_26353,N_26156);
xnor U26693 (N_26693,N_26301,N_26407);
or U26694 (N_26694,N_26496,N_26383);
and U26695 (N_26695,N_26453,N_26223);
nand U26696 (N_26696,N_26071,N_26368);
xor U26697 (N_26697,N_26305,N_26186);
nor U26698 (N_26698,N_26375,N_26296);
xnor U26699 (N_26699,N_26148,N_26047);
and U26700 (N_26700,N_26193,N_26444);
xnor U26701 (N_26701,N_26348,N_26218);
xnor U26702 (N_26702,N_26295,N_26089);
nor U26703 (N_26703,N_26117,N_26324);
and U26704 (N_26704,N_26408,N_26352);
xnor U26705 (N_26705,N_26110,N_26255);
and U26706 (N_26706,N_26030,N_26051);
nand U26707 (N_26707,N_26119,N_26233);
and U26708 (N_26708,N_26270,N_26490);
or U26709 (N_26709,N_26076,N_26358);
nand U26710 (N_26710,N_26226,N_26207);
or U26711 (N_26711,N_26014,N_26070);
and U26712 (N_26712,N_26319,N_26413);
xor U26713 (N_26713,N_26279,N_26069);
or U26714 (N_26714,N_26033,N_26366);
nand U26715 (N_26715,N_26055,N_26108);
or U26716 (N_26716,N_26038,N_26401);
or U26717 (N_26717,N_26420,N_26169);
or U26718 (N_26718,N_26274,N_26334);
nor U26719 (N_26719,N_26362,N_26371);
xor U26720 (N_26720,N_26283,N_26487);
nand U26721 (N_26721,N_26311,N_26158);
nand U26722 (N_26722,N_26126,N_26414);
and U26723 (N_26723,N_26073,N_26213);
xor U26724 (N_26724,N_26484,N_26206);
nor U26725 (N_26725,N_26314,N_26280);
and U26726 (N_26726,N_26054,N_26239);
xor U26727 (N_26727,N_26344,N_26425);
nor U26728 (N_26728,N_26422,N_26434);
or U26729 (N_26729,N_26017,N_26437);
and U26730 (N_26730,N_26003,N_26080);
nor U26731 (N_26731,N_26369,N_26459);
xor U26732 (N_26732,N_26479,N_26046);
xor U26733 (N_26733,N_26048,N_26106);
and U26734 (N_26734,N_26304,N_26471);
nor U26735 (N_26735,N_26140,N_26009);
and U26736 (N_26736,N_26370,N_26409);
or U26737 (N_26737,N_26325,N_26266);
and U26738 (N_26738,N_26287,N_26388);
nor U26739 (N_26739,N_26025,N_26189);
and U26740 (N_26740,N_26198,N_26286);
nor U26741 (N_26741,N_26277,N_26184);
nor U26742 (N_26742,N_26260,N_26464);
nand U26743 (N_26743,N_26380,N_26436);
nand U26744 (N_26744,N_26322,N_26349);
nor U26745 (N_26745,N_26394,N_26115);
or U26746 (N_26746,N_26472,N_26455);
nand U26747 (N_26747,N_26135,N_26253);
nor U26748 (N_26748,N_26027,N_26043);
nor U26749 (N_26749,N_26202,N_26387);
or U26750 (N_26750,N_26017,N_26413);
nor U26751 (N_26751,N_26013,N_26335);
nand U26752 (N_26752,N_26104,N_26389);
xor U26753 (N_26753,N_26203,N_26118);
xnor U26754 (N_26754,N_26387,N_26048);
or U26755 (N_26755,N_26102,N_26017);
nor U26756 (N_26756,N_26175,N_26045);
nor U26757 (N_26757,N_26332,N_26067);
or U26758 (N_26758,N_26252,N_26389);
nor U26759 (N_26759,N_26416,N_26264);
or U26760 (N_26760,N_26417,N_26231);
and U26761 (N_26761,N_26161,N_26115);
and U26762 (N_26762,N_26208,N_26132);
nand U26763 (N_26763,N_26333,N_26069);
nor U26764 (N_26764,N_26407,N_26251);
xor U26765 (N_26765,N_26378,N_26410);
and U26766 (N_26766,N_26419,N_26198);
and U26767 (N_26767,N_26258,N_26038);
xnor U26768 (N_26768,N_26339,N_26108);
and U26769 (N_26769,N_26470,N_26196);
xnor U26770 (N_26770,N_26323,N_26157);
or U26771 (N_26771,N_26346,N_26221);
or U26772 (N_26772,N_26214,N_26379);
xor U26773 (N_26773,N_26090,N_26434);
nand U26774 (N_26774,N_26118,N_26175);
xor U26775 (N_26775,N_26221,N_26313);
nor U26776 (N_26776,N_26115,N_26072);
nor U26777 (N_26777,N_26365,N_26278);
nor U26778 (N_26778,N_26487,N_26173);
nand U26779 (N_26779,N_26455,N_26467);
xnor U26780 (N_26780,N_26333,N_26045);
or U26781 (N_26781,N_26497,N_26300);
or U26782 (N_26782,N_26454,N_26178);
xor U26783 (N_26783,N_26477,N_26205);
nor U26784 (N_26784,N_26071,N_26430);
and U26785 (N_26785,N_26043,N_26085);
or U26786 (N_26786,N_26355,N_26166);
and U26787 (N_26787,N_26281,N_26404);
and U26788 (N_26788,N_26497,N_26316);
or U26789 (N_26789,N_26384,N_26143);
nand U26790 (N_26790,N_26184,N_26377);
xnor U26791 (N_26791,N_26359,N_26475);
nor U26792 (N_26792,N_26006,N_26468);
nor U26793 (N_26793,N_26374,N_26242);
and U26794 (N_26794,N_26390,N_26184);
and U26795 (N_26795,N_26484,N_26214);
nand U26796 (N_26796,N_26322,N_26491);
and U26797 (N_26797,N_26177,N_26267);
nand U26798 (N_26798,N_26167,N_26075);
or U26799 (N_26799,N_26227,N_26301);
nand U26800 (N_26800,N_26211,N_26140);
nor U26801 (N_26801,N_26000,N_26103);
or U26802 (N_26802,N_26083,N_26381);
and U26803 (N_26803,N_26355,N_26128);
nand U26804 (N_26804,N_26008,N_26166);
and U26805 (N_26805,N_26156,N_26306);
nand U26806 (N_26806,N_26252,N_26499);
nand U26807 (N_26807,N_26324,N_26171);
nand U26808 (N_26808,N_26318,N_26108);
and U26809 (N_26809,N_26348,N_26109);
xnor U26810 (N_26810,N_26423,N_26279);
nand U26811 (N_26811,N_26162,N_26149);
or U26812 (N_26812,N_26472,N_26137);
or U26813 (N_26813,N_26379,N_26254);
and U26814 (N_26814,N_26375,N_26080);
nand U26815 (N_26815,N_26485,N_26350);
or U26816 (N_26816,N_26486,N_26108);
or U26817 (N_26817,N_26174,N_26250);
or U26818 (N_26818,N_26044,N_26482);
nor U26819 (N_26819,N_26403,N_26455);
nand U26820 (N_26820,N_26424,N_26027);
or U26821 (N_26821,N_26471,N_26081);
nor U26822 (N_26822,N_26346,N_26111);
and U26823 (N_26823,N_26351,N_26427);
and U26824 (N_26824,N_26214,N_26351);
nor U26825 (N_26825,N_26456,N_26323);
and U26826 (N_26826,N_26413,N_26227);
xnor U26827 (N_26827,N_26043,N_26345);
and U26828 (N_26828,N_26067,N_26094);
nand U26829 (N_26829,N_26433,N_26200);
and U26830 (N_26830,N_26342,N_26193);
or U26831 (N_26831,N_26163,N_26041);
or U26832 (N_26832,N_26189,N_26065);
xnor U26833 (N_26833,N_26196,N_26039);
xnor U26834 (N_26834,N_26296,N_26367);
and U26835 (N_26835,N_26137,N_26369);
xnor U26836 (N_26836,N_26235,N_26138);
and U26837 (N_26837,N_26244,N_26273);
nand U26838 (N_26838,N_26261,N_26224);
nand U26839 (N_26839,N_26219,N_26084);
nand U26840 (N_26840,N_26434,N_26043);
or U26841 (N_26841,N_26471,N_26489);
nor U26842 (N_26842,N_26379,N_26117);
xnor U26843 (N_26843,N_26218,N_26003);
and U26844 (N_26844,N_26182,N_26196);
nor U26845 (N_26845,N_26443,N_26042);
and U26846 (N_26846,N_26487,N_26350);
or U26847 (N_26847,N_26402,N_26370);
and U26848 (N_26848,N_26361,N_26399);
or U26849 (N_26849,N_26019,N_26061);
xor U26850 (N_26850,N_26187,N_26015);
xor U26851 (N_26851,N_26202,N_26196);
xnor U26852 (N_26852,N_26385,N_26249);
nor U26853 (N_26853,N_26095,N_26298);
xnor U26854 (N_26854,N_26419,N_26120);
nor U26855 (N_26855,N_26493,N_26380);
xnor U26856 (N_26856,N_26441,N_26188);
nor U26857 (N_26857,N_26343,N_26321);
nand U26858 (N_26858,N_26367,N_26304);
nor U26859 (N_26859,N_26051,N_26385);
nor U26860 (N_26860,N_26288,N_26435);
nor U26861 (N_26861,N_26012,N_26135);
or U26862 (N_26862,N_26265,N_26099);
xor U26863 (N_26863,N_26407,N_26278);
or U26864 (N_26864,N_26449,N_26325);
xnor U26865 (N_26865,N_26449,N_26301);
nor U26866 (N_26866,N_26304,N_26233);
nor U26867 (N_26867,N_26158,N_26230);
nor U26868 (N_26868,N_26273,N_26332);
and U26869 (N_26869,N_26452,N_26080);
and U26870 (N_26870,N_26240,N_26053);
nand U26871 (N_26871,N_26206,N_26379);
and U26872 (N_26872,N_26087,N_26024);
nor U26873 (N_26873,N_26427,N_26120);
nand U26874 (N_26874,N_26317,N_26235);
xor U26875 (N_26875,N_26257,N_26490);
and U26876 (N_26876,N_26475,N_26408);
xnor U26877 (N_26877,N_26138,N_26195);
or U26878 (N_26878,N_26124,N_26062);
xor U26879 (N_26879,N_26113,N_26361);
nand U26880 (N_26880,N_26178,N_26253);
nand U26881 (N_26881,N_26313,N_26138);
nand U26882 (N_26882,N_26137,N_26220);
or U26883 (N_26883,N_26137,N_26460);
nor U26884 (N_26884,N_26339,N_26062);
nor U26885 (N_26885,N_26329,N_26102);
nor U26886 (N_26886,N_26013,N_26377);
xor U26887 (N_26887,N_26310,N_26075);
xnor U26888 (N_26888,N_26365,N_26214);
nand U26889 (N_26889,N_26440,N_26014);
nor U26890 (N_26890,N_26300,N_26188);
nand U26891 (N_26891,N_26397,N_26220);
or U26892 (N_26892,N_26265,N_26299);
xnor U26893 (N_26893,N_26374,N_26347);
nand U26894 (N_26894,N_26092,N_26192);
or U26895 (N_26895,N_26022,N_26057);
and U26896 (N_26896,N_26046,N_26190);
xor U26897 (N_26897,N_26308,N_26158);
and U26898 (N_26898,N_26128,N_26085);
or U26899 (N_26899,N_26345,N_26236);
nand U26900 (N_26900,N_26346,N_26198);
xor U26901 (N_26901,N_26495,N_26229);
nor U26902 (N_26902,N_26307,N_26057);
nand U26903 (N_26903,N_26429,N_26309);
or U26904 (N_26904,N_26355,N_26432);
or U26905 (N_26905,N_26390,N_26174);
nand U26906 (N_26906,N_26189,N_26037);
nand U26907 (N_26907,N_26306,N_26038);
and U26908 (N_26908,N_26143,N_26257);
and U26909 (N_26909,N_26022,N_26256);
nor U26910 (N_26910,N_26216,N_26133);
xnor U26911 (N_26911,N_26176,N_26217);
nand U26912 (N_26912,N_26385,N_26222);
or U26913 (N_26913,N_26188,N_26225);
xor U26914 (N_26914,N_26395,N_26349);
and U26915 (N_26915,N_26344,N_26090);
xnor U26916 (N_26916,N_26410,N_26286);
nor U26917 (N_26917,N_26454,N_26190);
and U26918 (N_26918,N_26235,N_26006);
nor U26919 (N_26919,N_26098,N_26365);
nor U26920 (N_26920,N_26389,N_26134);
xor U26921 (N_26921,N_26398,N_26098);
or U26922 (N_26922,N_26044,N_26189);
and U26923 (N_26923,N_26486,N_26392);
and U26924 (N_26924,N_26022,N_26251);
nor U26925 (N_26925,N_26091,N_26165);
or U26926 (N_26926,N_26080,N_26164);
xor U26927 (N_26927,N_26140,N_26317);
nor U26928 (N_26928,N_26050,N_26092);
and U26929 (N_26929,N_26412,N_26026);
or U26930 (N_26930,N_26448,N_26010);
nor U26931 (N_26931,N_26094,N_26199);
nor U26932 (N_26932,N_26267,N_26237);
and U26933 (N_26933,N_26179,N_26324);
xnor U26934 (N_26934,N_26439,N_26385);
xnor U26935 (N_26935,N_26309,N_26230);
or U26936 (N_26936,N_26235,N_26070);
xor U26937 (N_26937,N_26171,N_26019);
and U26938 (N_26938,N_26225,N_26478);
or U26939 (N_26939,N_26390,N_26335);
or U26940 (N_26940,N_26020,N_26466);
nor U26941 (N_26941,N_26434,N_26287);
or U26942 (N_26942,N_26418,N_26083);
and U26943 (N_26943,N_26240,N_26350);
and U26944 (N_26944,N_26311,N_26027);
nor U26945 (N_26945,N_26159,N_26471);
and U26946 (N_26946,N_26005,N_26077);
nand U26947 (N_26947,N_26387,N_26247);
or U26948 (N_26948,N_26209,N_26140);
nand U26949 (N_26949,N_26276,N_26103);
or U26950 (N_26950,N_26204,N_26010);
nor U26951 (N_26951,N_26156,N_26366);
nor U26952 (N_26952,N_26029,N_26265);
nor U26953 (N_26953,N_26100,N_26083);
xor U26954 (N_26954,N_26372,N_26362);
xor U26955 (N_26955,N_26204,N_26048);
and U26956 (N_26956,N_26075,N_26169);
xnor U26957 (N_26957,N_26116,N_26497);
nand U26958 (N_26958,N_26150,N_26174);
nand U26959 (N_26959,N_26291,N_26209);
nand U26960 (N_26960,N_26256,N_26169);
xor U26961 (N_26961,N_26068,N_26496);
xor U26962 (N_26962,N_26360,N_26417);
and U26963 (N_26963,N_26121,N_26489);
nand U26964 (N_26964,N_26088,N_26157);
nand U26965 (N_26965,N_26496,N_26401);
and U26966 (N_26966,N_26104,N_26183);
and U26967 (N_26967,N_26248,N_26239);
nand U26968 (N_26968,N_26435,N_26370);
nand U26969 (N_26969,N_26367,N_26235);
or U26970 (N_26970,N_26387,N_26070);
xor U26971 (N_26971,N_26306,N_26194);
xnor U26972 (N_26972,N_26170,N_26382);
nor U26973 (N_26973,N_26141,N_26332);
nor U26974 (N_26974,N_26206,N_26421);
and U26975 (N_26975,N_26170,N_26173);
nor U26976 (N_26976,N_26076,N_26112);
xor U26977 (N_26977,N_26197,N_26365);
or U26978 (N_26978,N_26058,N_26247);
or U26979 (N_26979,N_26129,N_26226);
and U26980 (N_26980,N_26459,N_26082);
nor U26981 (N_26981,N_26311,N_26110);
nand U26982 (N_26982,N_26328,N_26085);
nand U26983 (N_26983,N_26394,N_26017);
xnor U26984 (N_26984,N_26220,N_26121);
or U26985 (N_26985,N_26477,N_26348);
xnor U26986 (N_26986,N_26174,N_26102);
nand U26987 (N_26987,N_26309,N_26077);
nor U26988 (N_26988,N_26232,N_26165);
or U26989 (N_26989,N_26336,N_26046);
or U26990 (N_26990,N_26039,N_26166);
or U26991 (N_26991,N_26293,N_26009);
and U26992 (N_26992,N_26219,N_26345);
xor U26993 (N_26993,N_26381,N_26179);
xor U26994 (N_26994,N_26335,N_26386);
nand U26995 (N_26995,N_26216,N_26401);
xor U26996 (N_26996,N_26328,N_26277);
or U26997 (N_26997,N_26018,N_26436);
or U26998 (N_26998,N_26406,N_26026);
xor U26999 (N_26999,N_26474,N_26125);
or U27000 (N_27000,N_26512,N_26565);
and U27001 (N_27001,N_26961,N_26771);
nand U27002 (N_27002,N_26605,N_26845);
and U27003 (N_27003,N_26974,N_26611);
or U27004 (N_27004,N_26878,N_26937);
or U27005 (N_27005,N_26622,N_26618);
and U27006 (N_27006,N_26951,N_26986);
xnor U27007 (N_27007,N_26897,N_26922);
nor U27008 (N_27008,N_26969,N_26928);
nor U27009 (N_27009,N_26983,N_26893);
and U27010 (N_27010,N_26890,N_26631);
or U27011 (N_27011,N_26535,N_26901);
and U27012 (N_27012,N_26596,N_26874);
nor U27013 (N_27013,N_26954,N_26613);
nand U27014 (N_27014,N_26573,N_26697);
and U27015 (N_27015,N_26877,N_26673);
nor U27016 (N_27016,N_26526,N_26707);
and U27017 (N_27017,N_26676,N_26637);
xnor U27018 (N_27018,N_26552,N_26876);
or U27019 (N_27019,N_26790,N_26982);
or U27020 (N_27020,N_26515,N_26525);
nand U27021 (N_27021,N_26885,N_26973);
xor U27022 (N_27022,N_26532,N_26595);
and U27023 (N_27023,N_26602,N_26583);
and U27024 (N_27024,N_26628,N_26587);
nor U27025 (N_27025,N_26689,N_26988);
or U27026 (N_27026,N_26608,N_26940);
xnor U27027 (N_27027,N_26540,N_26541);
nand U27028 (N_27028,N_26942,N_26685);
and U27029 (N_27029,N_26609,N_26630);
and U27030 (N_27030,N_26971,N_26764);
nand U27031 (N_27031,N_26506,N_26946);
nor U27032 (N_27032,N_26518,N_26904);
nor U27033 (N_27033,N_26843,N_26776);
and U27034 (N_27034,N_26972,N_26849);
nand U27035 (N_27035,N_26619,N_26690);
nand U27036 (N_27036,N_26510,N_26726);
and U27037 (N_27037,N_26513,N_26669);
nand U27038 (N_27038,N_26538,N_26604);
xnor U27039 (N_27039,N_26746,N_26957);
nand U27040 (N_27040,N_26744,N_26811);
and U27041 (N_27041,N_26570,N_26956);
nand U27042 (N_27042,N_26812,N_26652);
nand U27043 (N_27043,N_26947,N_26994);
and U27044 (N_27044,N_26921,N_26606);
xor U27045 (N_27045,N_26949,N_26634);
or U27046 (N_27046,N_26614,N_26759);
xor U27047 (N_27047,N_26654,N_26722);
nor U27048 (N_27048,N_26700,N_26629);
nand U27049 (N_27049,N_26875,N_26842);
and U27050 (N_27050,N_26585,N_26865);
and U27051 (N_27051,N_26739,N_26985);
xor U27052 (N_27052,N_26660,N_26708);
nor U27053 (N_27053,N_26548,N_26643);
xnor U27054 (N_27054,N_26834,N_26559);
or U27055 (N_27055,N_26657,N_26958);
xnor U27056 (N_27056,N_26650,N_26980);
and U27057 (N_27057,N_26635,N_26888);
or U27058 (N_27058,N_26671,N_26755);
nand U27059 (N_27059,N_26576,N_26826);
or U27060 (N_27060,N_26800,N_26852);
and U27061 (N_27061,N_26765,N_26720);
nor U27062 (N_27062,N_26543,N_26896);
nand U27063 (N_27063,N_26627,N_26717);
xor U27064 (N_27064,N_26616,N_26793);
xnor U27065 (N_27065,N_26775,N_26560);
nor U27066 (N_27066,N_26781,N_26768);
and U27067 (N_27067,N_26655,N_26701);
and U27068 (N_27068,N_26955,N_26796);
nor U27069 (N_27069,N_26822,N_26688);
nand U27070 (N_27070,N_26561,N_26528);
nor U27071 (N_27071,N_26505,N_26626);
xor U27072 (N_27072,N_26913,N_26923);
xnor U27073 (N_27073,N_26572,N_26694);
xnor U27074 (N_27074,N_26967,N_26533);
nor U27075 (N_27075,N_26727,N_26792);
or U27076 (N_27076,N_26715,N_26617);
and U27077 (N_27077,N_26692,N_26522);
nand U27078 (N_27078,N_26906,N_26592);
and U27079 (N_27079,N_26879,N_26911);
and U27080 (N_27080,N_26733,N_26786);
nor U27081 (N_27081,N_26898,N_26502);
nand U27082 (N_27082,N_26615,N_26989);
or U27083 (N_27083,N_26553,N_26732);
nor U27084 (N_27084,N_26659,N_26646);
nand U27085 (N_27085,N_26927,N_26873);
or U27086 (N_27086,N_26806,N_26952);
and U27087 (N_27087,N_26883,N_26704);
nand U27088 (N_27088,N_26943,N_26527);
or U27089 (N_27089,N_26702,N_26953);
nor U27090 (N_27090,N_26820,N_26758);
or U27091 (N_27091,N_26607,N_26871);
or U27092 (N_27092,N_26864,N_26696);
xnor U27093 (N_27093,N_26664,N_26882);
nand U27094 (N_27094,N_26670,N_26537);
and U27095 (N_27095,N_26674,N_26723);
xnor U27096 (N_27096,N_26797,N_26799);
and U27097 (N_27097,N_26810,N_26677);
nand U27098 (N_27098,N_26580,N_26945);
or U27099 (N_27099,N_26567,N_26557);
and U27100 (N_27100,N_26519,N_26935);
nand U27101 (N_27101,N_26760,N_26716);
xnor U27102 (N_27102,N_26860,N_26509);
nand U27103 (N_27103,N_26909,N_26891);
and U27104 (N_27104,N_26839,N_26691);
or U27105 (N_27105,N_26672,N_26915);
xnor U27106 (N_27106,N_26939,N_26962);
nor U27107 (N_27107,N_26802,N_26621);
nor U27108 (N_27108,N_26681,N_26544);
nor U27109 (N_27109,N_26684,N_26597);
and U27110 (N_27110,N_26730,N_26818);
xnor U27111 (N_27111,N_26661,N_26959);
xnor U27112 (N_27112,N_26866,N_26836);
xor U27113 (N_27113,N_26908,N_26718);
or U27114 (N_27114,N_26872,N_26832);
nand U27115 (N_27115,N_26610,N_26554);
and U27116 (N_27116,N_26997,N_26881);
and U27117 (N_27117,N_26821,N_26714);
xor U27118 (N_27118,N_26964,N_26577);
and U27119 (N_27119,N_26749,N_26678);
or U27120 (N_27120,N_26662,N_26644);
xor U27121 (N_27121,N_26777,N_26639);
xnor U27122 (N_27122,N_26601,N_26992);
xor U27123 (N_27123,N_26785,N_26600);
nor U27124 (N_27124,N_26563,N_26903);
nor U27125 (N_27125,N_26582,N_26854);
xnor U27126 (N_27126,N_26679,N_26710);
nor U27127 (N_27127,N_26699,N_26511);
xor U27128 (N_27128,N_26593,N_26977);
and U27129 (N_27129,N_26816,N_26695);
nand U27130 (N_27130,N_26656,N_26584);
and U27131 (N_27131,N_26556,N_26753);
and U27132 (N_27132,N_26675,N_26536);
nor U27133 (N_27133,N_26795,N_26867);
nand U27134 (N_27134,N_26779,N_26682);
or U27135 (N_27135,N_26817,N_26990);
nor U27136 (N_27136,N_26791,N_26902);
nand U27137 (N_27137,N_26514,N_26920);
nand U27138 (N_27138,N_26649,N_26504);
nand U27139 (N_27139,N_26858,N_26719);
and U27140 (N_27140,N_26594,N_26801);
or U27141 (N_27141,N_26666,N_26963);
and U27142 (N_27142,N_26529,N_26516);
nor U27143 (N_27143,N_26778,N_26665);
nand U27144 (N_27144,N_26905,N_26725);
nor U27145 (N_27145,N_26996,N_26924);
or U27146 (N_27146,N_26814,N_26767);
or U27147 (N_27147,N_26706,N_26783);
nor U27148 (N_27148,N_26916,N_26965);
nor U27149 (N_27149,N_26772,N_26633);
nand U27150 (N_27150,N_26741,N_26803);
nand U27151 (N_27151,N_26523,N_26555);
nor U27152 (N_27152,N_26647,N_26500);
or U27153 (N_27153,N_26894,N_26620);
nand U27154 (N_27154,N_26861,N_26762);
nand U27155 (N_27155,N_26931,N_26970);
or U27156 (N_27156,N_26569,N_26912);
xor U27157 (N_27157,N_26848,N_26598);
xnor U27158 (N_27158,N_26827,N_26944);
xor U27159 (N_27159,N_26590,N_26625);
and U27160 (N_27160,N_26987,N_26815);
or U27161 (N_27161,N_26859,N_26805);
or U27162 (N_27162,N_26546,N_26917);
or U27163 (N_27163,N_26507,N_26651);
or U27164 (N_27164,N_26841,N_26641);
nand U27165 (N_27165,N_26591,N_26686);
nand U27166 (N_27166,N_26889,N_26807);
nor U27167 (N_27167,N_26603,N_26551);
xnor U27168 (N_27168,N_26711,N_26794);
and U27169 (N_27169,N_26887,N_26520);
nand U27170 (N_27170,N_26948,N_26539);
xor U27171 (N_27171,N_26774,N_26789);
nor U27172 (N_27172,N_26819,N_26769);
nand U27173 (N_27173,N_26763,N_26929);
or U27174 (N_27174,N_26787,N_26838);
or U27175 (N_27175,N_26825,N_26735);
nor U27176 (N_27176,N_26941,N_26586);
nor U27177 (N_27177,N_26693,N_26574);
nor U27178 (N_27178,N_26534,N_26632);
nor U27179 (N_27179,N_26648,N_26703);
xor U27180 (N_27180,N_26857,N_26738);
nand U27181 (N_27181,N_26809,N_26517);
and U27182 (N_27182,N_26668,N_26578);
nand U27183 (N_27183,N_26895,N_26930);
and U27184 (N_27184,N_26721,N_26743);
and U27185 (N_27185,N_26728,N_26978);
nor U27186 (N_27186,N_26566,N_26784);
xnor U27187 (N_27187,N_26729,N_26521);
and U27188 (N_27188,N_26724,N_26846);
nor U27189 (N_27189,N_26850,N_26575);
nand U27190 (N_27190,N_26562,N_26640);
or U27191 (N_27191,N_26737,N_26868);
or U27192 (N_27192,N_26558,N_26993);
or U27193 (N_27193,N_26835,N_26745);
or U27194 (N_27194,N_26705,N_26663);
xnor U27195 (N_27195,N_26828,N_26804);
xor U27196 (N_27196,N_26831,N_26918);
nor U27197 (N_27197,N_26933,N_26995);
and U27198 (N_27198,N_26748,N_26658);
nor U27199 (N_27199,N_26934,N_26823);
xnor U27200 (N_27200,N_26869,N_26757);
nand U27201 (N_27201,N_26837,N_26742);
nand U27202 (N_27202,N_26736,N_26975);
xnor U27203 (N_27203,N_26564,N_26900);
and U27204 (N_27204,N_26851,N_26960);
or U27205 (N_27205,N_26568,N_26863);
or U27206 (N_27206,N_26549,N_26687);
nor U27207 (N_27207,N_26680,N_26683);
or U27208 (N_27208,N_26919,N_26524);
nand U27209 (N_27209,N_26981,N_26756);
xor U27210 (N_27210,N_26501,N_26645);
nor U27211 (N_27211,N_26926,N_26813);
xor U27212 (N_27212,N_26833,N_26589);
nand U27213 (N_27213,N_26713,N_26581);
nand U27214 (N_27214,N_26766,N_26798);
or U27215 (N_27215,N_26824,N_26880);
xnor U27216 (N_27216,N_26653,N_26886);
xnor U27217 (N_27217,N_26747,N_26508);
nor U27218 (N_27218,N_26579,N_26550);
xor U27219 (N_27219,N_26862,N_26636);
nand U27220 (N_27220,N_26698,N_26731);
xor U27221 (N_27221,N_26936,N_26624);
and U27222 (N_27222,N_26808,N_26853);
nand U27223 (N_27223,N_26991,N_26870);
and U27224 (N_27224,N_26734,N_26892);
xnor U27225 (N_27225,N_26754,N_26938);
xor U27226 (N_27226,N_26782,N_26503);
and U27227 (N_27227,N_26547,N_26840);
nor U27228 (N_27228,N_26999,N_26998);
or U27229 (N_27229,N_26740,N_26984);
xor U27230 (N_27230,N_26530,N_26770);
or U27231 (N_27231,N_26910,N_26979);
nor U27232 (N_27232,N_26642,N_26709);
nor U27233 (N_27233,N_26976,N_26925);
nand U27234 (N_27234,N_26638,N_26542);
xnor U27235 (N_27235,N_26752,N_26968);
or U27236 (N_27236,N_26571,N_26788);
or U27237 (N_27237,N_26830,N_26899);
nand U27238 (N_27238,N_26599,N_26932);
or U27239 (N_27239,N_26750,N_26847);
xnor U27240 (N_27240,N_26623,N_26667);
and U27241 (N_27241,N_26612,N_26844);
and U27242 (N_27242,N_26966,N_26829);
nand U27243 (N_27243,N_26914,N_26588);
xor U27244 (N_27244,N_26751,N_26855);
and U27245 (N_27245,N_26950,N_26907);
nor U27246 (N_27246,N_26531,N_26761);
or U27247 (N_27247,N_26884,N_26773);
nor U27248 (N_27248,N_26780,N_26712);
and U27249 (N_27249,N_26545,N_26856);
nand U27250 (N_27250,N_26953,N_26501);
and U27251 (N_27251,N_26936,N_26616);
and U27252 (N_27252,N_26711,N_26667);
nor U27253 (N_27253,N_26849,N_26860);
nor U27254 (N_27254,N_26531,N_26751);
or U27255 (N_27255,N_26684,N_26905);
or U27256 (N_27256,N_26507,N_26591);
nand U27257 (N_27257,N_26769,N_26888);
xnor U27258 (N_27258,N_26771,N_26988);
nand U27259 (N_27259,N_26879,N_26525);
xnor U27260 (N_27260,N_26509,N_26955);
and U27261 (N_27261,N_26747,N_26694);
and U27262 (N_27262,N_26579,N_26733);
or U27263 (N_27263,N_26826,N_26606);
nor U27264 (N_27264,N_26850,N_26975);
nor U27265 (N_27265,N_26710,N_26623);
xor U27266 (N_27266,N_26770,N_26565);
nand U27267 (N_27267,N_26872,N_26581);
and U27268 (N_27268,N_26542,N_26864);
and U27269 (N_27269,N_26746,N_26653);
nor U27270 (N_27270,N_26778,N_26639);
xnor U27271 (N_27271,N_26792,N_26901);
or U27272 (N_27272,N_26626,N_26646);
xor U27273 (N_27273,N_26926,N_26974);
or U27274 (N_27274,N_26696,N_26993);
and U27275 (N_27275,N_26818,N_26738);
and U27276 (N_27276,N_26800,N_26929);
nor U27277 (N_27277,N_26534,N_26825);
and U27278 (N_27278,N_26763,N_26919);
and U27279 (N_27279,N_26671,N_26525);
or U27280 (N_27280,N_26931,N_26773);
nand U27281 (N_27281,N_26638,N_26775);
nor U27282 (N_27282,N_26626,N_26915);
or U27283 (N_27283,N_26619,N_26961);
nor U27284 (N_27284,N_26826,N_26745);
or U27285 (N_27285,N_26651,N_26950);
nor U27286 (N_27286,N_26775,N_26861);
xor U27287 (N_27287,N_26576,N_26507);
or U27288 (N_27288,N_26854,N_26808);
xor U27289 (N_27289,N_26593,N_26639);
xor U27290 (N_27290,N_26708,N_26817);
xor U27291 (N_27291,N_26767,N_26823);
and U27292 (N_27292,N_26684,N_26965);
or U27293 (N_27293,N_26913,N_26611);
or U27294 (N_27294,N_26920,N_26749);
nand U27295 (N_27295,N_26580,N_26577);
nand U27296 (N_27296,N_26661,N_26951);
or U27297 (N_27297,N_26932,N_26506);
nor U27298 (N_27298,N_26759,N_26991);
and U27299 (N_27299,N_26755,N_26773);
nand U27300 (N_27300,N_26606,N_26952);
and U27301 (N_27301,N_26711,N_26887);
and U27302 (N_27302,N_26791,N_26665);
nor U27303 (N_27303,N_26581,N_26638);
and U27304 (N_27304,N_26792,N_26663);
and U27305 (N_27305,N_26644,N_26564);
xor U27306 (N_27306,N_26882,N_26649);
nor U27307 (N_27307,N_26514,N_26856);
or U27308 (N_27308,N_26778,N_26544);
nor U27309 (N_27309,N_26869,N_26921);
or U27310 (N_27310,N_26895,N_26560);
xnor U27311 (N_27311,N_26874,N_26605);
nand U27312 (N_27312,N_26644,N_26655);
nand U27313 (N_27313,N_26580,N_26899);
nand U27314 (N_27314,N_26615,N_26968);
nor U27315 (N_27315,N_26916,N_26828);
nand U27316 (N_27316,N_26822,N_26513);
nor U27317 (N_27317,N_26698,N_26536);
xnor U27318 (N_27318,N_26891,N_26560);
nand U27319 (N_27319,N_26881,N_26882);
xor U27320 (N_27320,N_26640,N_26909);
nor U27321 (N_27321,N_26531,N_26650);
nand U27322 (N_27322,N_26853,N_26999);
nand U27323 (N_27323,N_26612,N_26520);
xnor U27324 (N_27324,N_26677,N_26821);
or U27325 (N_27325,N_26558,N_26663);
nand U27326 (N_27326,N_26540,N_26549);
and U27327 (N_27327,N_26825,N_26606);
nor U27328 (N_27328,N_26857,N_26995);
nor U27329 (N_27329,N_26956,N_26583);
xnor U27330 (N_27330,N_26547,N_26568);
and U27331 (N_27331,N_26564,N_26543);
or U27332 (N_27332,N_26544,N_26533);
or U27333 (N_27333,N_26696,N_26614);
nor U27334 (N_27334,N_26533,N_26940);
xor U27335 (N_27335,N_26560,N_26712);
xor U27336 (N_27336,N_26694,N_26954);
or U27337 (N_27337,N_26536,N_26808);
or U27338 (N_27338,N_26745,N_26823);
and U27339 (N_27339,N_26573,N_26535);
xnor U27340 (N_27340,N_26808,N_26982);
xor U27341 (N_27341,N_26591,N_26944);
xnor U27342 (N_27342,N_26977,N_26650);
xor U27343 (N_27343,N_26872,N_26805);
nor U27344 (N_27344,N_26546,N_26777);
nand U27345 (N_27345,N_26674,N_26889);
nand U27346 (N_27346,N_26632,N_26559);
nor U27347 (N_27347,N_26882,N_26516);
xnor U27348 (N_27348,N_26925,N_26608);
or U27349 (N_27349,N_26869,N_26858);
nor U27350 (N_27350,N_26906,N_26801);
nand U27351 (N_27351,N_26710,N_26675);
xnor U27352 (N_27352,N_26513,N_26889);
nand U27353 (N_27353,N_26920,N_26530);
nand U27354 (N_27354,N_26822,N_26776);
and U27355 (N_27355,N_26780,N_26946);
nor U27356 (N_27356,N_26801,N_26913);
and U27357 (N_27357,N_26791,N_26746);
nand U27358 (N_27358,N_26901,N_26915);
nand U27359 (N_27359,N_26891,N_26911);
xor U27360 (N_27360,N_26521,N_26782);
xor U27361 (N_27361,N_26974,N_26846);
or U27362 (N_27362,N_26659,N_26673);
and U27363 (N_27363,N_26934,N_26960);
nand U27364 (N_27364,N_26867,N_26687);
nand U27365 (N_27365,N_26842,N_26874);
nor U27366 (N_27366,N_26586,N_26592);
xor U27367 (N_27367,N_26666,N_26829);
or U27368 (N_27368,N_26656,N_26557);
nor U27369 (N_27369,N_26796,N_26925);
nand U27370 (N_27370,N_26567,N_26517);
nor U27371 (N_27371,N_26775,N_26681);
or U27372 (N_27372,N_26813,N_26701);
nor U27373 (N_27373,N_26633,N_26794);
nand U27374 (N_27374,N_26626,N_26963);
xnor U27375 (N_27375,N_26643,N_26737);
xnor U27376 (N_27376,N_26714,N_26943);
xor U27377 (N_27377,N_26835,N_26974);
nor U27378 (N_27378,N_26834,N_26853);
and U27379 (N_27379,N_26531,N_26768);
xor U27380 (N_27380,N_26530,N_26512);
nor U27381 (N_27381,N_26652,N_26847);
and U27382 (N_27382,N_26959,N_26808);
xor U27383 (N_27383,N_26623,N_26727);
nand U27384 (N_27384,N_26707,N_26758);
nor U27385 (N_27385,N_26813,N_26801);
and U27386 (N_27386,N_26649,N_26898);
nor U27387 (N_27387,N_26509,N_26541);
and U27388 (N_27388,N_26772,N_26821);
nand U27389 (N_27389,N_26794,N_26927);
and U27390 (N_27390,N_26945,N_26667);
nand U27391 (N_27391,N_26807,N_26672);
nand U27392 (N_27392,N_26696,N_26656);
nor U27393 (N_27393,N_26693,N_26613);
and U27394 (N_27394,N_26598,N_26974);
and U27395 (N_27395,N_26866,N_26849);
nand U27396 (N_27396,N_26791,N_26624);
nand U27397 (N_27397,N_26575,N_26624);
nor U27398 (N_27398,N_26972,N_26975);
xor U27399 (N_27399,N_26847,N_26619);
nor U27400 (N_27400,N_26830,N_26888);
or U27401 (N_27401,N_26828,N_26922);
and U27402 (N_27402,N_26649,N_26732);
nand U27403 (N_27403,N_26880,N_26536);
or U27404 (N_27404,N_26806,N_26609);
nor U27405 (N_27405,N_26702,N_26666);
nor U27406 (N_27406,N_26994,N_26548);
nand U27407 (N_27407,N_26968,N_26922);
xnor U27408 (N_27408,N_26807,N_26757);
or U27409 (N_27409,N_26808,N_26996);
or U27410 (N_27410,N_26772,N_26659);
and U27411 (N_27411,N_26693,N_26583);
and U27412 (N_27412,N_26859,N_26738);
and U27413 (N_27413,N_26525,N_26647);
nor U27414 (N_27414,N_26935,N_26724);
and U27415 (N_27415,N_26507,N_26804);
nand U27416 (N_27416,N_26613,N_26606);
or U27417 (N_27417,N_26929,N_26646);
nand U27418 (N_27418,N_26560,N_26646);
nor U27419 (N_27419,N_26735,N_26836);
and U27420 (N_27420,N_26518,N_26840);
or U27421 (N_27421,N_26679,N_26529);
or U27422 (N_27422,N_26535,N_26811);
xor U27423 (N_27423,N_26625,N_26822);
and U27424 (N_27424,N_26514,N_26916);
or U27425 (N_27425,N_26697,N_26515);
nand U27426 (N_27426,N_26814,N_26842);
xor U27427 (N_27427,N_26548,N_26505);
nand U27428 (N_27428,N_26997,N_26886);
and U27429 (N_27429,N_26842,N_26701);
or U27430 (N_27430,N_26834,N_26927);
xnor U27431 (N_27431,N_26691,N_26609);
and U27432 (N_27432,N_26577,N_26545);
or U27433 (N_27433,N_26563,N_26589);
nor U27434 (N_27434,N_26716,N_26920);
or U27435 (N_27435,N_26839,N_26582);
xnor U27436 (N_27436,N_26744,N_26545);
nand U27437 (N_27437,N_26612,N_26618);
or U27438 (N_27438,N_26850,N_26644);
and U27439 (N_27439,N_26889,N_26661);
nor U27440 (N_27440,N_26991,N_26595);
xor U27441 (N_27441,N_26767,N_26871);
or U27442 (N_27442,N_26563,N_26580);
or U27443 (N_27443,N_26644,N_26994);
xnor U27444 (N_27444,N_26896,N_26705);
nor U27445 (N_27445,N_26788,N_26910);
and U27446 (N_27446,N_26651,N_26531);
nand U27447 (N_27447,N_26922,N_26752);
and U27448 (N_27448,N_26565,N_26525);
xor U27449 (N_27449,N_26532,N_26748);
nand U27450 (N_27450,N_26563,N_26676);
and U27451 (N_27451,N_26890,N_26591);
and U27452 (N_27452,N_26925,N_26728);
xor U27453 (N_27453,N_26607,N_26818);
xor U27454 (N_27454,N_26748,N_26903);
nor U27455 (N_27455,N_26514,N_26889);
nor U27456 (N_27456,N_26754,N_26597);
nor U27457 (N_27457,N_26648,N_26525);
xnor U27458 (N_27458,N_26743,N_26975);
or U27459 (N_27459,N_26994,N_26741);
nor U27460 (N_27460,N_26832,N_26896);
or U27461 (N_27461,N_26869,N_26642);
or U27462 (N_27462,N_26584,N_26567);
xnor U27463 (N_27463,N_26666,N_26947);
nand U27464 (N_27464,N_26917,N_26924);
nand U27465 (N_27465,N_26900,N_26985);
nor U27466 (N_27466,N_26582,N_26928);
or U27467 (N_27467,N_26745,N_26585);
xor U27468 (N_27468,N_26747,N_26801);
nor U27469 (N_27469,N_26804,N_26599);
nor U27470 (N_27470,N_26503,N_26752);
xor U27471 (N_27471,N_26967,N_26744);
xnor U27472 (N_27472,N_26994,N_26760);
xnor U27473 (N_27473,N_26764,N_26880);
or U27474 (N_27474,N_26890,N_26547);
xor U27475 (N_27475,N_26556,N_26681);
nand U27476 (N_27476,N_26788,N_26609);
nand U27477 (N_27477,N_26545,N_26761);
nor U27478 (N_27478,N_26556,N_26679);
nor U27479 (N_27479,N_26602,N_26885);
nor U27480 (N_27480,N_26781,N_26502);
nand U27481 (N_27481,N_26898,N_26961);
or U27482 (N_27482,N_26794,N_26830);
nor U27483 (N_27483,N_26634,N_26704);
nor U27484 (N_27484,N_26895,N_26834);
or U27485 (N_27485,N_26554,N_26622);
xnor U27486 (N_27486,N_26906,N_26980);
nor U27487 (N_27487,N_26782,N_26815);
nand U27488 (N_27488,N_26992,N_26938);
nand U27489 (N_27489,N_26714,N_26892);
xor U27490 (N_27490,N_26862,N_26925);
xor U27491 (N_27491,N_26586,N_26631);
nor U27492 (N_27492,N_26921,N_26544);
nor U27493 (N_27493,N_26894,N_26769);
nor U27494 (N_27494,N_26979,N_26500);
xor U27495 (N_27495,N_26673,N_26926);
xor U27496 (N_27496,N_26987,N_26902);
nand U27497 (N_27497,N_26736,N_26544);
nor U27498 (N_27498,N_26933,N_26586);
nand U27499 (N_27499,N_26600,N_26643);
nor U27500 (N_27500,N_27270,N_27139);
nor U27501 (N_27501,N_27282,N_27369);
nor U27502 (N_27502,N_27482,N_27303);
nand U27503 (N_27503,N_27127,N_27304);
or U27504 (N_27504,N_27019,N_27310);
nor U27505 (N_27505,N_27147,N_27494);
nand U27506 (N_27506,N_27215,N_27368);
nor U27507 (N_27507,N_27097,N_27119);
and U27508 (N_27508,N_27418,N_27030);
and U27509 (N_27509,N_27212,N_27202);
xnor U27510 (N_27510,N_27098,N_27436);
or U27511 (N_27511,N_27296,N_27474);
xor U27512 (N_27512,N_27092,N_27354);
or U27513 (N_27513,N_27117,N_27286);
nand U27514 (N_27514,N_27166,N_27031);
xor U27515 (N_27515,N_27041,N_27116);
xnor U27516 (N_27516,N_27024,N_27475);
or U27517 (N_27517,N_27471,N_27032);
and U27518 (N_27518,N_27184,N_27143);
xor U27519 (N_27519,N_27292,N_27002);
nor U27520 (N_27520,N_27083,N_27462);
xnor U27521 (N_27521,N_27306,N_27382);
nand U27522 (N_27522,N_27331,N_27342);
or U27523 (N_27523,N_27073,N_27407);
xor U27524 (N_27524,N_27105,N_27273);
nor U27525 (N_27525,N_27063,N_27112);
and U27526 (N_27526,N_27335,N_27185);
and U27527 (N_27527,N_27449,N_27090);
nand U27528 (N_27528,N_27221,N_27069);
or U27529 (N_27529,N_27084,N_27042);
or U27530 (N_27530,N_27037,N_27093);
and U27531 (N_27531,N_27326,N_27114);
and U27532 (N_27532,N_27159,N_27240);
or U27533 (N_27533,N_27197,N_27461);
nand U27534 (N_27534,N_27198,N_27076);
nor U27535 (N_27535,N_27179,N_27386);
and U27536 (N_27536,N_27062,N_27344);
or U27537 (N_27537,N_27200,N_27433);
nor U27538 (N_27538,N_27214,N_27497);
xnor U27539 (N_27539,N_27301,N_27103);
xnor U27540 (N_27540,N_27205,N_27177);
xor U27541 (N_27541,N_27495,N_27350);
and U27542 (N_27542,N_27249,N_27079);
nor U27543 (N_27543,N_27460,N_27291);
or U27544 (N_27544,N_27314,N_27065);
nor U27545 (N_27545,N_27034,N_27142);
nand U27546 (N_27546,N_27104,N_27489);
xor U27547 (N_27547,N_27137,N_27328);
nor U27548 (N_27548,N_27153,N_27053);
and U27549 (N_27549,N_27188,N_27287);
or U27550 (N_27550,N_27237,N_27408);
and U27551 (N_27551,N_27399,N_27472);
and U27552 (N_27552,N_27318,N_27278);
xnor U27553 (N_27553,N_27338,N_27048);
or U27554 (N_27554,N_27036,N_27089);
nor U27555 (N_27555,N_27364,N_27219);
nor U27556 (N_27556,N_27323,N_27280);
nor U27557 (N_27557,N_27252,N_27124);
and U27558 (N_27558,N_27224,N_27411);
or U27559 (N_27559,N_27173,N_27001);
or U27560 (N_27560,N_27220,N_27193);
xnor U27561 (N_27561,N_27014,N_27072);
or U27562 (N_27562,N_27261,N_27426);
nand U27563 (N_27563,N_27035,N_27351);
xor U27564 (N_27564,N_27107,N_27021);
nor U27565 (N_27565,N_27122,N_27458);
nor U27566 (N_27566,N_27447,N_27023);
nor U27567 (N_27567,N_27401,N_27316);
or U27568 (N_27568,N_27181,N_27487);
nand U27569 (N_27569,N_27134,N_27130);
nand U27570 (N_27570,N_27272,N_27123);
or U27571 (N_27571,N_27064,N_27044);
nand U27572 (N_27572,N_27476,N_27319);
or U27573 (N_27573,N_27377,N_27047);
nor U27574 (N_27574,N_27420,N_27321);
and U27575 (N_27575,N_27275,N_27209);
xnor U27576 (N_27576,N_27308,N_27346);
nor U27577 (N_27577,N_27359,N_27235);
or U27578 (N_27578,N_27492,N_27125);
nand U27579 (N_27579,N_27040,N_27102);
nor U27580 (N_27580,N_27467,N_27315);
and U27581 (N_27581,N_27225,N_27080);
nor U27582 (N_27582,N_27329,N_27337);
xor U27583 (N_27583,N_27448,N_27266);
nor U27584 (N_27584,N_27239,N_27496);
nor U27585 (N_27585,N_27330,N_27324);
nand U27586 (N_27586,N_27227,N_27176);
or U27587 (N_27587,N_27478,N_27243);
xor U27588 (N_27588,N_27245,N_27250);
nor U27589 (N_27589,N_27419,N_27012);
or U27590 (N_27590,N_27208,N_27455);
and U27591 (N_27591,N_27480,N_27333);
nand U27592 (N_27592,N_27340,N_27247);
and U27593 (N_27593,N_27135,N_27357);
or U27594 (N_27594,N_27388,N_27484);
or U27595 (N_27595,N_27009,N_27477);
or U27596 (N_27596,N_27425,N_27450);
nand U27597 (N_27597,N_27189,N_27438);
nand U27598 (N_27598,N_27432,N_27441);
and U27599 (N_27599,N_27059,N_27263);
nor U27600 (N_27600,N_27045,N_27375);
or U27601 (N_27601,N_27233,N_27332);
and U27602 (N_27602,N_27336,N_27068);
xnor U27603 (N_27603,N_27171,N_27317);
nor U27604 (N_27604,N_27160,N_27038);
and U27605 (N_27605,N_27196,N_27162);
nor U27606 (N_27606,N_27121,N_27155);
nor U27607 (N_27607,N_27394,N_27352);
or U27608 (N_27608,N_27311,N_27417);
or U27609 (N_27609,N_27051,N_27192);
nand U27610 (N_27610,N_27229,N_27349);
and U27611 (N_27611,N_27404,N_27442);
nor U27612 (N_27612,N_27269,N_27082);
nand U27613 (N_27613,N_27011,N_27046);
and U27614 (N_27614,N_27365,N_27213);
and U27615 (N_27615,N_27183,N_27360);
or U27616 (N_27616,N_27094,N_27446);
nor U27617 (N_27617,N_27279,N_27078);
xnor U27618 (N_27618,N_27416,N_27422);
or U27619 (N_27619,N_27466,N_27099);
nand U27620 (N_27620,N_27115,N_27373);
xnor U27621 (N_27621,N_27445,N_27334);
nor U27622 (N_27622,N_27187,N_27056);
and U27623 (N_27623,N_27085,N_27473);
and U27624 (N_27624,N_27216,N_27148);
xor U27625 (N_27625,N_27295,N_27300);
xor U27626 (N_27626,N_27409,N_27381);
nand U27627 (N_27627,N_27136,N_27271);
nor U27628 (N_27628,N_27405,N_27486);
xnor U27629 (N_27629,N_27383,N_27033);
xnor U27630 (N_27630,N_27015,N_27157);
xor U27631 (N_27631,N_27008,N_27169);
nor U27632 (N_27632,N_27236,N_27452);
nand U27633 (N_27633,N_27234,N_27387);
and U27634 (N_27634,N_27231,N_27353);
xor U27635 (N_27635,N_27457,N_27067);
and U27636 (N_27636,N_27100,N_27361);
nand U27637 (N_27637,N_27043,N_27443);
nand U27638 (N_27638,N_27312,N_27463);
and U27639 (N_27639,N_27451,N_27256);
and U27640 (N_27640,N_27077,N_27400);
or U27641 (N_27641,N_27479,N_27454);
and U27642 (N_27642,N_27459,N_27307);
xnor U27643 (N_27643,N_27228,N_27367);
nand U27644 (N_27644,N_27174,N_27398);
xnor U27645 (N_27645,N_27430,N_27374);
or U27646 (N_27646,N_27022,N_27428);
and U27647 (N_27647,N_27091,N_27293);
or U27648 (N_27648,N_27248,N_27242);
and U27649 (N_27649,N_27003,N_27488);
or U27650 (N_27650,N_27110,N_27362);
or U27651 (N_27651,N_27020,N_27309);
and U27652 (N_27652,N_27406,N_27071);
xor U27653 (N_27653,N_27039,N_27376);
xnor U27654 (N_27654,N_27049,N_27194);
nor U27655 (N_27655,N_27088,N_27289);
nor U27656 (N_27656,N_27027,N_27244);
or U27657 (N_27657,N_27016,N_27253);
nand U27658 (N_27658,N_27058,N_27464);
nor U27659 (N_27659,N_27120,N_27281);
nor U27660 (N_27660,N_27490,N_27060);
nor U27661 (N_27661,N_27028,N_27133);
nor U27662 (N_27662,N_27222,N_27010);
xnor U27663 (N_27663,N_27274,N_27440);
or U27664 (N_27664,N_27156,N_27264);
and U27665 (N_27665,N_27435,N_27207);
or U27666 (N_27666,N_27358,N_27498);
or U27667 (N_27667,N_27203,N_27163);
or U27668 (N_27668,N_27149,N_27017);
and U27669 (N_27669,N_27186,N_27366);
nor U27670 (N_27670,N_27178,N_27070);
and U27671 (N_27671,N_27029,N_27087);
xor U27672 (N_27672,N_27429,N_27283);
and U27673 (N_27673,N_27146,N_27370);
xnor U27674 (N_27674,N_27054,N_27276);
or U27675 (N_27675,N_27439,N_27111);
nand U27676 (N_27676,N_27481,N_27106);
nor U27677 (N_27677,N_27206,N_27493);
and U27678 (N_27678,N_27371,N_27355);
and U27679 (N_27679,N_27129,N_27403);
xor U27680 (N_27680,N_27223,N_27140);
and U27681 (N_27681,N_27285,N_27018);
xor U27682 (N_27682,N_27257,N_27218);
nor U27683 (N_27683,N_27341,N_27182);
xnor U27684 (N_27684,N_27013,N_27158);
or U27685 (N_27685,N_27195,N_27066);
and U27686 (N_27686,N_27232,N_27199);
nand U27687 (N_27687,N_27431,N_27074);
nand U27688 (N_27688,N_27165,N_27101);
nand U27689 (N_27689,N_27005,N_27325);
nand U27690 (N_27690,N_27141,N_27345);
and U27691 (N_27691,N_27412,N_27327);
nor U27692 (N_27692,N_27423,N_27347);
nor U27693 (N_27693,N_27499,N_27131);
nand U27694 (N_27694,N_27230,N_27305);
nor U27695 (N_27695,N_27000,N_27437);
nor U27696 (N_27696,N_27402,N_27161);
nor U27697 (N_27697,N_27421,N_27172);
nor U27698 (N_27698,N_27251,N_27343);
nor U27699 (N_27699,N_27190,N_27095);
and U27700 (N_27700,N_27145,N_27491);
xnor U27701 (N_27701,N_27026,N_27313);
or U27702 (N_27702,N_27210,N_27393);
nand U27703 (N_27703,N_27246,N_27109);
nand U27704 (N_27704,N_27268,N_27086);
nor U27705 (N_27705,N_27175,N_27465);
and U27706 (N_27706,N_27262,N_27372);
nor U27707 (N_27707,N_27164,N_27055);
nor U27708 (N_27708,N_27004,N_27180);
xnor U27709 (N_27709,N_27126,N_27151);
or U27710 (N_27710,N_27456,N_27414);
xor U27711 (N_27711,N_27138,N_27132);
nor U27712 (N_27712,N_27294,N_27469);
or U27713 (N_27713,N_27167,N_27061);
nor U27714 (N_27714,N_27288,N_27396);
or U27715 (N_27715,N_27434,N_27150);
nand U27716 (N_27716,N_27259,N_27241);
xor U27717 (N_27717,N_27384,N_27427);
and U27718 (N_27718,N_27277,N_27297);
xnor U27719 (N_27719,N_27363,N_27152);
or U27720 (N_27720,N_27444,N_27260);
and U27721 (N_27721,N_27392,N_27050);
nor U27722 (N_27722,N_27238,N_27006);
nor U27723 (N_27723,N_27470,N_27254);
xnor U27724 (N_27724,N_27284,N_27385);
and U27725 (N_27725,N_27204,N_27290);
nand U27726 (N_27726,N_27217,N_27211);
xor U27727 (N_27727,N_27397,N_27299);
and U27728 (N_27728,N_27395,N_27302);
nand U27729 (N_27729,N_27007,N_27390);
and U27730 (N_27730,N_27265,N_27424);
nor U27731 (N_27731,N_27154,N_27379);
and U27732 (N_27732,N_27320,N_27380);
nand U27733 (N_27733,N_27453,N_27201);
xor U27734 (N_27734,N_27191,N_27483);
nor U27735 (N_27735,N_27258,N_27144);
or U27736 (N_27736,N_27413,N_27322);
xnor U27737 (N_27737,N_27485,N_27113);
and U27738 (N_27738,N_27128,N_27339);
and U27739 (N_27739,N_27255,N_27025);
and U27740 (N_27740,N_27468,N_27348);
or U27741 (N_27741,N_27391,N_27267);
nor U27742 (N_27742,N_27108,N_27389);
or U27743 (N_27743,N_27378,N_27052);
xnor U27744 (N_27744,N_27075,N_27226);
nor U27745 (N_27745,N_27118,N_27298);
nor U27746 (N_27746,N_27410,N_27081);
nand U27747 (N_27747,N_27170,N_27057);
nand U27748 (N_27748,N_27096,N_27356);
nand U27749 (N_27749,N_27415,N_27168);
and U27750 (N_27750,N_27052,N_27292);
nand U27751 (N_27751,N_27138,N_27394);
or U27752 (N_27752,N_27461,N_27140);
and U27753 (N_27753,N_27053,N_27077);
nand U27754 (N_27754,N_27414,N_27106);
nor U27755 (N_27755,N_27197,N_27482);
xor U27756 (N_27756,N_27321,N_27241);
xor U27757 (N_27757,N_27436,N_27331);
nor U27758 (N_27758,N_27327,N_27012);
or U27759 (N_27759,N_27388,N_27435);
and U27760 (N_27760,N_27478,N_27329);
and U27761 (N_27761,N_27428,N_27019);
and U27762 (N_27762,N_27154,N_27174);
and U27763 (N_27763,N_27197,N_27374);
and U27764 (N_27764,N_27205,N_27333);
and U27765 (N_27765,N_27071,N_27195);
nand U27766 (N_27766,N_27002,N_27165);
and U27767 (N_27767,N_27313,N_27162);
nor U27768 (N_27768,N_27207,N_27083);
nor U27769 (N_27769,N_27105,N_27418);
xnor U27770 (N_27770,N_27015,N_27321);
xor U27771 (N_27771,N_27292,N_27368);
xor U27772 (N_27772,N_27420,N_27083);
nor U27773 (N_27773,N_27002,N_27490);
xor U27774 (N_27774,N_27216,N_27357);
nand U27775 (N_27775,N_27294,N_27228);
nand U27776 (N_27776,N_27184,N_27013);
nand U27777 (N_27777,N_27431,N_27304);
nor U27778 (N_27778,N_27290,N_27242);
xor U27779 (N_27779,N_27110,N_27318);
xor U27780 (N_27780,N_27417,N_27385);
nand U27781 (N_27781,N_27429,N_27340);
xor U27782 (N_27782,N_27132,N_27114);
or U27783 (N_27783,N_27201,N_27231);
nand U27784 (N_27784,N_27469,N_27069);
or U27785 (N_27785,N_27454,N_27084);
nand U27786 (N_27786,N_27461,N_27298);
xor U27787 (N_27787,N_27268,N_27172);
or U27788 (N_27788,N_27205,N_27474);
xnor U27789 (N_27789,N_27462,N_27053);
and U27790 (N_27790,N_27007,N_27055);
or U27791 (N_27791,N_27206,N_27016);
and U27792 (N_27792,N_27443,N_27299);
and U27793 (N_27793,N_27240,N_27099);
nor U27794 (N_27794,N_27337,N_27002);
xor U27795 (N_27795,N_27493,N_27174);
or U27796 (N_27796,N_27224,N_27283);
and U27797 (N_27797,N_27225,N_27102);
and U27798 (N_27798,N_27091,N_27162);
and U27799 (N_27799,N_27382,N_27064);
and U27800 (N_27800,N_27110,N_27255);
or U27801 (N_27801,N_27034,N_27006);
or U27802 (N_27802,N_27040,N_27031);
nor U27803 (N_27803,N_27464,N_27323);
nand U27804 (N_27804,N_27084,N_27372);
xnor U27805 (N_27805,N_27222,N_27012);
xor U27806 (N_27806,N_27347,N_27495);
xnor U27807 (N_27807,N_27363,N_27365);
xor U27808 (N_27808,N_27333,N_27473);
or U27809 (N_27809,N_27081,N_27131);
and U27810 (N_27810,N_27058,N_27072);
nand U27811 (N_27811,N_27043,N_27199);
nand U27812 (N_27812,N_27236,N_27455);
nand U27813 (N_27813,N_27283,N_27124);
xor U27814 (N_27814,N_27442,N_27304);
or U27815 (N_27815,N_27084,N_27450);
and U27816 (N_27816,N_27280,N_27483);
nor U27817 (N_27817,N_27003,N_27332);
nor U27818 (N_27818,N_27457,N_27049);
xnor U27819 (N_27819,N_27383,N_27207);
and U27820 (N_27820,N_27008,N_27182);
and U27821 (N_27821,N_27494,N_27050);
xnor U27822 (N_27822,N_27491,N_27135);
and U27823 (N_27823,N_27493,N_27189);
and U27824 (N_27824,N_27460,N_27267);
and U27825 (N_27825,N_27337,N_27168);
and U27826 (N_27826,N_27310,N_27149);
xor U27827 (N_27827,N_27047,N_27072);
nor U27828 (N_27828,N_27242,N_27144);
and U27829 (N_27829,N_27329,N_27492);
nand U27830 (N_27830,N_27049,N_27103);
xor U27831 (N_27831,N_27017,N_27167);
and U27832 (N_27832,N_27276,N_27450);
xnor U27833 (N_27833,N_27210,N_27335);
nand U27834 (N_27834,N_27403,N_27092);
or U27835 (N_27835,N_27105,N_27189);
nand U27836 (N_27836,N_27466,N_27130);
xor U27837 (N_27837,N_27120,N_27277);
xnor U27838 (N_27838,N_27001,N_27081);
or U27839 (N_27839,N_27463,N_27097);
nand U27840 (N_27840,N_27464,N_27008);
or U27841 (N_27841,N_27443,N_27480);
and U27842 (N_27842,N_27404,N_27348);
nand U27843 (N_27843,N_27135,N_27258);
xnor U27844 (N_27844,N_27185,N_27284);
nor U27845 (N_27845,N_27388,N_27421);
xnor U27846 (N_27846,N_27368,N_27375);
nor U27847 (N_27847,N_27274,N_27194);
or U27848 (N_27848,N_27158,N_27472);
and U27849 (N_27849,N_27217,N_27332);
nor U27850 (N_27850,N_27001,N_27403);
nand U27851 (N_27851,N_27319,N_27295);
and U27852 (N_27852,N_27305,N_27445);
nor U27853 (N_27853,N_27034,N_27235);
or U27854 (N_27854,N_27278,N_27034);
nand U27855 (N_27855,N_27376,N_27195);
nor U27856 (N_27856,N_27341,N_27409);
nor U27857 (N_27857,N_27096,N_27082);
xnor U27858 (N_27858,N_27019,N_27376);
or U27859 (N_27859,N_27177,N_27016);
and U27860 (N_27860,N_27064,N_27484);
nor U27861 (N_27861,N_27181,N_27315);
and U27862 (N_27862,N_27372,N_27102);
and U27863 (N_27863,N_27492,N_27259);
and U27864 (N_27864,N_27420,N_27095);
nor U27865 (N_27865,N_27365,N_27254);
nor U27866 (N_27866,N_27452,N_27313);
or U27867 (N_27867,N_27293,N_27262);
or U27868 (N_27868,N_27435,N_27145);
and U27869 (N_27869,N_27398,N_27362);
nor U27870 (N_27870,N_27072,N_27119);
xnor U27871 (N_27871,N_27458,N_27438);
xor U27872 (N_27872,N_27451,N_27021);
nand U27873 (N_27873,N_27462,N_27337);
and U27874 (N_27874,N_27028,N_27265);
nor U27875 (N_27875,N_27186,N_27157);
or U27876 (N_27876,N_27099,N_27370);
or U27877 (N_27877,N_27095,N_27256);
nor U27878 (N_27878,N_27332,N_27021);
and U27879 (N_27879,N_27470,N_27061);
nand U27880 (N_27880,N_27026,N_27236);
nor U27881 (N_27881,N_27256,N_27316);
nand U27882 (N_27882,N_27095,N_27288);
nor U27883 (N_27883,N_27251,N_27040);
nand U27884 (N_27884,N_27294,N_27286);
nor U27885 (N_27885,N_27163,N_27090);
nand U27886 (N_27886,N_27074,N_27028);
xor U27887 (N_27887,N_27058,N_27469);
nand U27888 (N_27888,N_27121,N_27339);
and U27889 (N_27889,N_27478,N_27207);
nand U27890 (N_27890,N_27196,N_27223);
xnor U27891 (N_27891,N_27472,N_27401);
nor U27892 (N_27892,N_27177,N_27189);
or U27893 (N_27893,N_27046,N_27322);
and U27894 (N_27894,N_27454,N_27048);
nor U27895 (N_27895,N_27371,N_27391);
nand U27896 (N_27896,N_27120,N_27065);
nor U27897 (N_27897,N_27103,N_27419);
or U27898 (N_27898,N_27324,N_27245);
nand U27899 (N_27899,N_27100,N_27366);
or U27900 (N_27900,N_27143,N_27149);
or U27901 (N_27901,N_27381,N_27269);
or U27902 (N_27902,N_27077,N_27184);
nor U27903 (N_27903,N_27143,N_27274);
nand U27904 (N_27904,N_27028,N_27022);
and U27905 (N_27905,N_27422,N_27097);
nor U27906 (N_27906,N_27425,N_27456);
nand U27907 (N_27907,N_27257,N_27163);
nand U27908 (N_27908,N_27319,N_27321);
xor U27909 (N_27909,N_27475,N_27106);
xnor U27910 (N_27910,N_27419,N_27032);
xor U27911 (N_27911,N_27236,N_27281);
nand U27912 (N_27912,N_27203,N_27369);
or U27913 (N_27913,N_27011,N_27112);
xnor U27914 (N_27914,N_27219,N_27235);
nand U27915 (N_27915,N_27032,N_27361);
or U27916 (N_27916,N_27306,N_27119);
nor U27917 (N_27917,N_27287,N_27158);
xor U27918 (N_27918,N_27198,N_27256);
or U27919 (N_27919,N_27403,N_27201);
or U27920 (N_27920,N_27190,N_27284);
xnor U27921 (N_27921,N_27078,N_27145);
nor U27922 (N_27922,N_27433,N_27430);
xnor U27923 (N_27923,N_27413,N_27082);
nor U27924 (N_27924,N_27404,N_27363);
nor U27925 (N_27925,N_27295,N_27293);
or U27926 (N_27926,N_27024,N_27493);
or U27927 (N_27927,N_27252,N_27430);
xor U27928 (N_27928,N_27239,N_27319);
or U27929 (N_27929,N_27370,N_27125);
and U27930 (N_27930,N_27004,N_27401);
and U27931 (N_27931,N_27264,N_27128);
xor U27932 (N_27932,N_27292,N_27134);
nand U27933 (N_27933,N_27028,N_27347);
nand U27934 (N_27934,N_27471,N_27301);
xor U27935 (N_27935,N_27329,N_27403);
nand U27936 (N_27936,N_27157,N_27206);
xor U27937 (N_27937,N_27181,N_27428);
or U27938 (N_27938,N_27071,N_27125);
nor U27939 (N_27939,N_27134,N_27356);
xor U27940 (N_27940,N_27162,N_27066);
or U27941 (N_27941,N_27425,N_27020);
and U27942 (N_27942,N_27107,N_27052);
or U27943 (N_27943,N_27338,N_27453);
xnor U27944 (N_27944,N_27134,N_27412);
and U27945 (N_27945,N_27082,N_27299);
xnor U27946 (N_27946,N_27279,N_27093);
nor U27947 (N_27947,N_27344,N_27329);
and U27948 (N_27948,N_27013,N_27066);
or U27949 (N_27949,N_27306,N_27464);
nand U27950 (N_27950,N_27393,N_27312);
nor U27951 (N_27951,N_27398,N_27479);
nand U27952 (N_27952,N_27198,N_27287);
xnor U27953 (N_27953,N_27442,N_27086);
xnor U27954 (N_27954,N_27346,N_27036);
nand U27955 (N_27955,N_27259,N_27135);
or U27956 (N_27956,N_27325,N_27024);
nor U27957 (N_27957,N_27443,N_27294);
and U27958 (N_27958,N_27352,N_27082);
xor U27959 (N_27959,N_27491,N_27000);
and U27960 (N_27960,N_27351,N_27007);
or U27961 (N_27961,N_27245,N_27054);
or U27962 (N_27962,N_27299,N_27426);
or U27963 (N_27963,N_27186,N_27477);
or U27964 (N_27964,N_27474,N_27209);
nand U27965 (N_27965,N_27295,N_27132);
nor U27966 (N_27966,N_27354,N_27256);
and U27967 (N_27967,N_27166,N_27026);
nand U27968 (N_27968,N_27276,N_27233);
nor U27969 (N_27969,N_27016,N_27461);
and U27970 (N_27970,N_27367,N_27172);
nand U27971 (N_27971,N_27241,N_27288);
and U27972 (N_27972,N_27452,N_27201);
and U27973 (N_27973,N_27150,N_27329);
nand U27974 (N_27974,N_27374,N_27042);
and U27975 (N_27975,N_27156,N_27300);
nor U27976 (N_27976,N_27390,N_27086);
xor U27977 (N_27977,N_27482,N_27149);
nand U27978 (N_27978,N_27210,N_27470);
xor U27979 (N_27979,N_27069,N_27239);
xor U27980 (N_27980,N_27138,N_27182);
nor U27981 (N_27981,N_27145,N_27382);
nand U27982 (N_27982,N_27389,N_27232);
and U27983 (N_27983,N_27409,N_27352);
or U27984 (N_27984,N_27019,N_27358);
and U27985 (N_27985,N_27485,N_27073);
xnor U27986 (N_27986,N_27402,N_27188);
xnor U27987 (N_27987,N_27350,N_27214);
nor U27988 (N_27988,N_27012,N_27382);
and U27989 (N_27989,N_27285,N_27225);
or U27990 (N_27990,N_27106,N_27290);
xnor U27991 (N_27991,N_27380,N_27310);
xnor U27992 (N_27992,N_27229,N_27409);
xor U27993 (N_27993,N_27383,N_27166);
nor U27994 (N_27994,N_27083,N_27342);
nand U27995 (N_27995,N_27226,N_27100);
or U27996 (N_27996,N_27280,N_27166);
or U27997 (N_27997,N_27204,N_27305);
and U27998 (N_27998,N_27016,N_27397);
nand U27999 (N_27999,N_27173,N_27436);
and U28000 (N_28000,N_27525,N_27775);
nor U28001 (N_28001,N_27666,N_27996);
xor U28002 (N_28002,N_27661,N_27536);
or U28003 (N_28003,N_27688,N_27760);
xor U28004 (N_28004,N_27513,N_27514);
and U28005 (N_28005,N_27889,N_27989);
nand U28006 (N_28006,N_27755,N_27560);
nand U28007 (N_28007,N_27736,N_27552);
nand U28008 (N_28008,N_27898,N_27680);
nor U28009 (N_28009,N_27501,N_27977);
xor U28010 (N_28010,N_27551,N_27527);
and U28011 (N_28011,N_27569,N_27772);
nand U28012 (N_28012,N_27553,N_27657);
nor U28013 (N_28013,N_27921,N_27679);
nor U28014 (N_28014,N_27998,N_27927);
and U28015 (N_28015,N_27646,N_27872);
nor U28016 (N_28016,N_27803,N_27531);
nor U28017 (N_28017,N_27521,N_27817);
and U28018 (N_28018,N_27913,N_27693);
nand U28019 (N_28019,N_27503,N_27726);
nand U28020 (N_28020,N_27783,N_27587);
nor U28021 (N_28021,N_27918,N_27846);
nor U28022 (N_28022,N_27548,N_27582);
xor U28023 (N_28023,N_27554,N_27778);
nand U28024 (N_28024,N_27863,N_27792);
and U28025 (N_28025,N_27696,N_27765);
xnor U28026 (N_28026,N_27598,N_27820);
xor U28027 (N_28027,N_27987,N_27647);
nor U28028 (N_28028,N_27723,N_27887);
and U28029 (N_28029,N_27814,N_27859);
or U28030 (N_28030,N_27526,N_27586);
nand U28031 (N_28031,N_27782,N_27896);
or U28032 (N_28032,N_27754,N_27728);
nor U28033 (N_28033,N_27773,N_27707);
xnor U28034 (N_28034,N_27625,N_27881);
xnor U28035 (N_28035,N_27629,N_27664);
and U28036 (N_28036,N_27681,N_27890);
or U28037 (N_28037,N_27861,N_27502);
xor U28038 (N_28038,N_27711,N_27549);
and U28039 (N_28039,N_27836,N_27979);
nor U28040 (N_28040,N_27825,N_27850);
or U28041 (N_28041,N_27784,N_27591);
xor U28042 (N_28042,N_27867,N_27540);
and U28043 (N_28043,N_27518,N_27718);
xnor U28044 (N_28044,N_27749,N_27700);
and U28045 (N_28045,N_27592,N_27758);
xor U28046 (N_28046,N_27577,N_27806);
nor U28047 (N_28047,N_27544,N_27605);
or U28048 (N_28048,N_27877,N_27830);
nand U28049 (N_28049,N_27562,N_27878);
xor U28050 (N_28050,N_27507,N_27858);
nand U28051 (N_28051,N_27505,N_27829);
nor U28052 (N_28052,N_27671,N_27692);
nor U28053 (N_28053,N_27997,N_27737);
nand U28054 (N_28054,N_27766,N_27904);
nor U28055 (N_28055,N_27885,N_27663);
nor U28056 (N_28056,N_27510,N_27866);
nor U28057 (N_28057,N_27988,N_27851);
and U28058 (N_28058,N_27824,N_27500);
nor U28059 (N_28059,N_27807,N_27715);
xnor U28060 (N_28060,N_27788,N_27689);
xor U28061 (N_28061,N_27662,N_27945);
and U28062 (N_28062,N_27897,N_27812);
or U28063 (N_28063,N_27912,N_27798);
or U28064 (N_28064,N_27504,N_27815);
xor U28065 (N_28065,N_27837,N_27741);
and U28066 (N_28066,N_27732,N_27687);
nor U28067 (N_28067,N_27570,N_27771);
nand U28068 (N_28068,N_27805,N_27839);
nor U28069 (N_28069,N_27917,N_27739);
and U28070 (N_28070,N_27966,N_27848);
nor U28071 (N_28071,N_27962,N_27862);
or U28072 (N_28072,N_27516,N_27808);
xor U28073 (N_28073,N_27932,N_27543);
nand U28074 (N_28074,N_27600,N_27992);
nand U28075 (N_28075,N_27734,N_27705);
nor U28076 (N_28076,N_27604,N_27940);
xor U28077 (N_28077,N_27995,N_27937);
nor U28078 (N_28078,N_27642,N_27686);
nand U28079 (N_28079,N_27575,N_27573);
and U28080 (N_28080,N_27909,N_27954);
nand U28081 (N_28081,N_27626,N_27901);
nand U28082 (N_28082,N_27789,N_27742);
and U28083 (N_28083,N_27821,N_27865);
xor U28084 (N_28084,N_27698,N_27910);
or U28085 (N_28085,N_27948,N_27994);
and U28086 (N_28086,N_27709,N_27660);
and U28087 (N_28087,N_27751,N_27975);
nor U28088 (N_28088,N_27740,N_27935);
nand U28089 (N_28089,N_27621,N_27701);
xor U28090 (N_28090,N_27982,N_27614);
or U28091 (N_28091,N_27632,N_27844);
nor U28092 (N_28092,N_27767,N_27941);
or U28093 (N_28093,N_27610,N_27597);
nand U28094 (N_28094,N_27747,N_27984);
and U28095 (N_28095,N_27968,N_27845);
and U28096 (N_28096,N_27923,N_27834);
and U28097 (N_28097,N_27753,N_27716);
nor U28098 (N_28098,N_27894,N_27672);
nand U28099 (N_28099,N_27744,N_27973);
xor U28100 (N_28100,N_27888,N_27731);
xnor U28101 (N_28101,N_27702,N_27602);
and U28102 (N_28102,N_27965,N_27779);
and U28103 (N_28103,N_27777,N_27978);
nor U28104 (N_28104,N_27833,N_27920);
nand U28105 (N_28105,N_27934,N_27883);
nand U28106 (N_28106,N_27704,N_27892);
or U28107 (N_28107,N_27972,N_27931);
xnor U28108 (N_28108,N_27690,N_27761);
nand U28109 (N_28109,N_27607,N_27727);
xor U28110 (N_28110,N_27508,N_27590);
xnor U28111 (N_28111,N_27776,N_27710);
and U28112 (N_28112,N_27627,N_27541);
nor U28113 (N_28113,N_27608,N_27619);
or U28114 (N_28114,N_27944,N_27969);
xor U28115 (N_28115,N_27819,N_27585);
and U28116 (N_28116,N_27787,N_27802);
nand U28117 (N_28117,N_27653,N_27871);
nor U28118 (N_28118,N_27769,N_27724);
and U28119 (N_28119,N_27738,N_27964);
and U28120 (N_28120,N_27799,N_27974);
nor U28121 (N_28121,N_27857,N_27532);
xor U28122 (N_28122,N_27922,N_27869);
nor U28123 (N_28123,N_27643,N_27870);
or U28124 (N_28124,N_27649,N_27603);
nor U28125 (N_28125,N_27622,N_27512);
nand U28126 (N_28126,N_27841,N_27990);
nand U28127 (N_28127,N_27509,N_27804);
xnor U28128 (N_28128,N_27929,N_27623);
or U28129 (N_28129,N_27615,N_27983);
nor U28130 (N_28130,N_27578,N_27659);
xnor U28131 (N_28131,N_27667,N_27564);
nor U28132 (N_28132,N_27524,N_27713);
and U28133 (N_28133,N_27958,N_27900);
nand U28134 (N_28134,N_27847,N_27993);
nand U28135 (N_28135,N_27919,N_27682);
nand U28136 (N_28136,N_27854,N_27949);
nand U28137 (N_28137,N_27832,N_27556);
xnor U28138 (N_28138,N_27624,N_27568);
or U28139 (N_28139,N_27594,N_27907);
or U28140 (N_28140,N_27743,N_27719);
or U28141 (N_28141,N_27547,N_27546);
and U28142 (N_28142,N_27674,N_27899);
nor U28143 (N_28143,N_27538,N_27580);
nand U28144 (N_28144,N_27533,N_27926);
xor U28145 (N_28145,N_27645,N_27786);
and U28146 (N_28146,N_27976,N_27811);
or U28147 (N_28147,N_27635,N_27906);
nor U28148 (N_28148,N_27519,N_27971);
xor U28149 (N_28149,N_27528,N_27567);
nand U28150 (N_28150,N_27764,N_27571);
nand U28151 (N_28151,N_27785,N_27763);
or U28152 (N_28152,N_27565,N_27658);
xor U28153 (N_28153,N_27694,N_27951);
and U28154 (N_28154,N_27612,N_27759);
nand U28155 (N_28155,N_27952,N_27515);
nand U28156 (N_28156,N_27638,N_27818);
nand U28157 (N_28157,N_27566,N_27875);
nand U28158 (N_28158,N_27831,N_27903);
and U28159 (N_28159,N_27796,N_27695);
nand U28160 (N_28160,N_27522,N_27916);
nand U28161 (N_28161,N_27557,N_27529);
nand U28162 (N_28162,N_27616,N_27684);
nor U28163 (N_28163,N_27670,N_27725);
xor U28164 (N_28164,N_27601,N_27746);
xor U28165 (N_28165,N_27947,N_27676);
nor U28166 (N_28166,N_27656,N_27613);
or U28167 (N_28167,N_27697,N_27599);
and U28168 (N_28168,N_27843,N_27930);
nor U28169 (N_28169,N_27581,N_27618);
xnor U28170 (N_28170,N_27595,N_27790);
xor U28171 (N_28171,N_27868,N_27559);
nor U28172 (N_28172,N_27840,N_27712);
nor U28173 (N_28173,N_27644,N_27555);
nor U28174 (N_28174,N_27955,N_27584);
nand U28175 (N_28175,N_27641,N_27908);
nand U28176 (N_28176,N_27780,N_27838);
nor U28177 (N_28177,N_27880,N_27950);
or U28178 (N_28178,N_27856,N_27855);
nor U28179 (N_28179,N_27634,N_27874);
nand U28180 (N_28180,N_27620,N_27762);
and U28181 (N_28181,N_27946,N_27511);
nand U28182 (N_28182,N_27905,N_27828);
xor U28183 (N_28183,N_27722,N_27537);
or U28184 (N_28184,N_27886,N_27640);
nand U28185 (N_28185,N_27520,N_27733);
or U28186 (N_28186,N_27714,N_27823);
nand U28187 (N_28187,N_27650,N_27933);
nor U28188 (N_28188,N_27506,N_27669);
or U28189 (N_28189,N_27652,N_27774);
nand U28190 (N_28190,N_27530,N_27654);
or U28191 (N_28191,N_27579,N_27911);
and U28192 (N_28192,N_27961,N_27963);
nor U28193 (N_28193,N_27835,N_27826);
nand U28194 (N_28194,N_27956,N_27720);
or U28195 (N_28195,N_27985,N_27800);
nor U28196 (N_28196,N_27517,N_27611);
xnor U28197 (N_28197,N_27860,N_27745);
xnor U28198 (N_28198,N_27882,N_27980);
or U28199 (N_28199,N_27879,N_27558);
nor U28200 (N_28200,N_27864,N_27668);
nand U28201 (N_28201,N_27708,N_27574);
xnor U28202 (N_28202,N_27636,N_27563);
and U28203 (N_28203,N_27721,N_27809);
xor U28204 (N_28204,N_27683,N_27545);
nand U28205 (N_28205,N_27730,N_27925);
and U28206 (N_28206,N_27675,N_27827);
or U28207 (N_28207,N_27801,N_27539);
and U28208 (N_28208,N_27967,N_27735);
nor U28209 (N_28209,N_27852,N_27606);
or U28210 (N_28210,N_27842,N_27703);
nand U28211 (N_28211,N_27991,N_27797);
nand U28212 (N_28212,N_27628,N_27884);
nand U28213 (N_28213,N_27588,N_27748);
or U28214 (N_28214,N_27924,N_27609);
and U28215 (N_28215,N_27893,N_27576);
and U28216 (N_28216,N_27943,N_27813);
nand U28217 (N_28217,N_27942,N_27757);
xor U28218 (N_28218,N_27691,N_27928);
nand U28219 (N_28219,N_27593,N_27699);
or U28220 (N_28220,N_27849,N_27639);
and U28221 (N_28221,N_27756,N_27793);
xnor U28222 (N_28222,N_27936,N_27822);
or U28223 (N_28223,N_27902,N_27673);
nand U28224 (N_28224,N_27938,N_27589);
or U28225 (N_28225,N_27953,N_27750);
nor U28226 (N_28226,N_27550,N_27665);
and U28227 (N_28227,N_27523,N_27939);
xnor U28228 (N_28228,N_27542,N_27752);
and U28229 (N_28229,N_27816,N_27637);
nand U28230 (N_28230,N_27791,N_27596);
xnor U28231 (N_28231,N_27915,N_27853);
or U28232 (N_28232,N_27895,N_27631);
or U28233 (N_28233,N_27981,N_27583);
xnor U28234 (N_28234,N_27633,N_27957);
nand U28235 (N_28235,N_27561,N_27678);
nor U28236 (N_28236,N_27534,N_27876);
xnor U28237 (N_28237,N_27648,N_27795);
xor U28238 (N_28238,N_27781,N_27677);
nor U28239 (N_28239,N_27572,N_27794);
xnor U28240 (N_28240,N_27706,N_27810);
nand U28241 (N_28241,N_27655,N_27914);
or U28242 (N_28242,N_27729,N_27959);
nand U28243 (N_28243,N_27685,N_27617);
and U28244 (N_28244,N_27535,N_27891);
nand U28245 (N_28245,N_27768,N_27999);
or U28246 (N_28246,N_27651,N_27873);
xor U28247 (N_28247,N_27630,N_27770);
nand U28248 (N_28248,N_27970,N_27717);
and U28249 (N_28249,N_27986,N_27960);
nor U28250 (N_28250,N_27829,N_27969);
nor U28251 (N_28251,N_27816,N_27789);
xor U28252 (N_28252,N_27504,N_27960);
or U28253 (N_28253,N_27571,N_27956);
or U28254 (N_28254,N_27823,N_27708);
xnor U28255 (N_28255,N_27620,N_27659);
nor U28256 (N_28256,N_27921,N_27657);
nor U28257 (N_28257,N_27893,N_27777);
and U28258 (N_28258,N_27954,N_27675);
and U28259 (N_28259,N_27974,N_27679);
xnor U28260 (N_28260,N_27964,N_27812);
xor U28261 (N_28261,N_27934,N_27686);
or U28262 (N_28262,N_27993,N_27883);
or U28263 (N_28263,N_27841,N_27699);
xor U28264 (N_28264,N_27502,N_27755);
xor U28265 (N_28265,N_27910,N_27762);
or U28266 (N_28266,N_27821,N_27625);
and U28267 (N_28267,N_27534,N_27907);
nor U28268 (N_28268,N_27508,N_27644);
and U28269 (N_28269,N_27904,N_27605);
or U28270 (N_28270,N_27684,N_27593);
nor U28271 (N_28271,N_27718,N_27593);
xnor U28272 (N_28272,N_27821,N_27965);
and U28273 (N_28273,N_27732,N_27946);
and U28274 (N_28274,N_27790,N_27705);
nand U28275 (N_28275,N_27807,N_27953);
nor U28276 (N_28276,N_27995,N_27757);
nand U28277 (N_28277,N_27804,N_27892);
or U28278 (N_28278,N_27506,N_27847);
or U28279 (N_28279,N_27779,N_27801);
or U28280 (N_28280,N_27919,N_27933);
nand U28281 (N_28281,N_27878,N_27898);
nand U28282 (N_28282,N_27739,N_27775);
xor U28283 (N_28283,N_27950,N_27824);
nand U28284 (N_28284,N_27841,N_27607);
nand U28285 (N_28285,N_27700,N_27975);
or U28286 (N_28286,N_27899,N_27610);
nand U28287 (N_28287,N_27680,N_27872);
nand U28288 (N_28288,N_27617,N_27955);
or U28289 (N_28289,N_27625,N_27949);
xor U28290 (N_28290,N_27931,N_27625);
nor U28291 (N_28291,N_27577,N_27870);
or U28292 (N_28292,N_27714,N_27660);
nor U28293 (N_28293,N_27769,N_27511);
or U28294 (N_28294,N_27940,N_27540);
or U28295 (N_28295,N_27707,N_27908);
nand U28296 (N_28296,N_27525,N_27959);
and U28297 (N_28297,N_27662,N_27904);
xor U28298 (N_28298,N_27812,N_27558);
nor U28299 (N_28299,N_27827,N_27930);
xnor U28300 (N_28300,N_27501,N_27832);
nand U28301 (N_28301,N_27722,N_27975);
and U28302 (N_28302,N_27665,N_27924);
or U28303 (N_28303,N_27622,N_27713);
nand U28304 (N_28304,N_27542,N_27652);
xor U28305 (N_28305,N_27658,N_27582);
nor U28306 (N_28306,N_27932,N_27695);
nor U28307 (N_28307,N_27770,N_27587);
nor U28308 (N_28308,N_27598,N_27552);
and U28309 (N_28309,N_27517,N_27948);
or U28310 (N_28310,N_27631,N_27839);
nand U28311 (N_28311,N_27877,N_27977);
xnor U28312 (N_28312,N_27921,N_27604);
nor U28313 (N_28313,N_27989,N_27780);
and U28314 (N_28314,N_27971,N_27894);
and U28315 (N_28315,N_27955,N_27984);
xor U28316 (N_28316,N_27773,N_27901);
xor U28317 (N_28317,N_27759,N_27568);
nand U28318 (N_28318,N_27983,N_27876);
xor U28319 (N_28319,N_27933,N_27541);
xor U28320 (N_28320,N_27956,N_27644);
nand U28321 (N_28321,N_27918,N_27656);
nor U28322 (N_28322,N_27677,N_27824);
nor U28323 (N_28323,N_27505,N_27593);
and U28324 (N_28324,N_27641,N_27706);
or U28325 (N_28325,N_27806,N_27516);
or U28326 (N_28326,N_27849,N_27776);
nor U28327 (N_28327,N_27862,N_27773);
or U28328 (N_28328,N_27504,N_27769);
and U28329 (N_28329,N_27868,N_27717);
xnor U28330 (N_28330,N_27681,N_27746);
nor U28331 (N_28331,N_27889,N_27536);
nand U28332 (N_28332,N_27766,N_27982);
and U28333 (N_28333,N_27521,N_27550);
and U28334 (N_28334,N_27923,N_27815);
nor U28335 (N_28335,N_27926,N_27671);
and U28336 (N_28336,N_27676,N_27599);
or U28337 (N_28337,N_27849,N_27514);
xor U28338 (N_28338,N_27609,N_27960);
and U28339 (N_28339,N_27659,N_27592);
nor U28340 (N_28340,N_27972,N_27965);
xnor U28341 (N_28341,N_27849,N_27932);
nor U28342 (N_28342,N_27680,N_27829);
nor U28343 (N_28343,N_27630,N_27800);
or U28344 (N_28344,N_27560,N_27600);
nor U28345 (N_28345,N_27970,N_27895);
nand U28346 (N_28346,N_27846,N_27851);
nor U28347 (N_28347,N_27927,N_27672);
or U28348 (N_28348,N_27864,N_27628);
nor U28349 (N_28349,N_27704,N_27765);
nor U28350 (N_28350,N_27954,N_27705);
xnor U28351 (N_28351,N_27973,N_27603);
and U28352 (N_28352,N_27972,N_27943);
nor U28353 (N_28353,N_27902,N_27789);
xnor U28354 (N_28354,N_27761,N_27535);
xor U28355 (N_28355,N_27680,N_27540);
xnor U28356 (N_28356,N_27665,N_27976);
or U28357 (N_28357,N_27689,N_27792);
nand U28358 (N_28358,N_27793,N_27961);
xor U28359 (N_28359,N_27534,N_27812);
and U28360 (N_28360,N_27949,N_27991);
and U28361 (N_28361,N_27808,N_27882);
or U28362 (N_28362,N_27858,N_27752);
or U28363 (N_28363,N_27634,N_27796);
or U28364 (N_28364,N_27816,N_27511);
nor U28365 (N_28365,N_27967,N_27520);
nor U28366 (N_28366,N_27629,N_27657);
nor U28367 (N_28367,N_27577,N_27816);
or U28368 (N_28368,N_27550,N_27597);
nor U28369 (N_28369,N_27765,N_27638);
and U28370 (N_28370,N_27667,N_27596);
nor U28371 (N_28371,N_27746,N_27535);
nand U28372 (N_28372,N_27863,N_27656);
nand U28373 (N_28373,N_27751,N_27658);
xor U28374 (N_28374,N_27579,N_27664);
nand U28375 (N_28375,N_27891,N_27962);
nor U28376 (N_28376,N_27678,N_27783);
and U28377 (N_28377,N_27838,N_27667);
nor U28378 (N_28378,N_27752,N_27620);
xor U28379 (N_28379,N_27672,N_27523);
nor U28380 (N_28380,N_27613,N_27612);
nand U28381 (N_28381,N_27925,N_27689);
nor U28382 (N_28382,N_27765,N_27981);
nand U28383 (N_28383,N_27899,N_27679);
and U28384 (N_28384,N_27537,N_27560);
xnor U28385 (N_28385,N_27524,N_27629);
and U28386 (N_28386,N_27669,N_27730);
nor U28387 (N_28387,N_27667,N_27800);
xor U28388 (N_28388,N_27986,N_27859);
nand U28389 (N_28389,N_27737,N_27814);
nor U28390 (N_28390,N_27544,N_27815);
and U28391 (N_28391,N_27575,N_27714);
or U28392 (N_28392,N_27815,N_27814);
or U28393 (N_28393,N_27638,N_27624);
and U28394 (N_28394,N_27795,N_27947);
or U28395 (N_28395,N_27624,N_27577);
and U28396 (N_28396,N_27869,N_27978);
nand U28397 (N_28397,N_27701,N_27967);
xnor U28398 (N_28398,N_27864,N_27538);
and U28399 (N_28399,N_27655,N_27514);
and U28400 (N_28400,N_27923,N_27865);
or U28401 (N_28401,N_27762,N_27867);
and U28402 (N_28402,N_27654,N_27818);
and U28403 (N_28403,N_27928,N_27894);
nand U28404 (N_28404,N_27545,N_27954);
xor U28405 (N_28405,N_27582,N_27968);
nor U28406 (N_28406,N_27721,N_27857);
xnor U28407 (N_28407,N_27542,N_27514);
or U28408 (N_28408,N_27509,N_27779);
nand U28409 (N_28409,N_27766,N_27950);
nor U28410 (N_28410,N_27512,N_27551);
nor U28411 (N_28411,N_27879,N_27874);
nor U28412 (N_28412,N_27900,N_27862);
or U28413 (N_28413,N_27502,N_27532);
or U28414 (N_28414,N_27667,N_27770);
nand U28415 (N_28415,N_27954,N_27829);
or U28416 (N_28416,N_27835,N_27943);
nor U28417 (N_28417,N_27774,N_27576);
or U28418 (N_28418,N_27557,N_27565);
and U28419 (N_28419,N_27856,N_27816);
and U28420 (N_28420,N_27630,N_27511);
xor U28421 (N_28421,N_27953,N_27846);
nor U28422 (N_28422,N_27942,N_27878);
and U28423 (N_28423,N_27676,N_27731);
nand U28424 (N_28424,N_27769,N_27702);
nand U28425 (N_28425,N_27620,N_27950);
nand U28426 (N_28426,N_27616,N_27685);
nand U28427 (N_28427,N_27992,N_27781);
nor U28428 (N_28428,N_27632,N_27794);
nor U28429 (N_28429,N_27764,N_27843);
nor U28430 (N_28430,N_27878,N_27870);
nand U28431 (N_28431,N_27576,N_27882);
or U28432 (N_28432,N_27695,N_27865);
and U28433 (N_28433,N_27729,N_27785);
xnor U28434 (N_28434,N_27927,N_27537);
or U28435 (N_28435,N_27537,N_27652);
and U28436 (N_28436,N_27510,N_27587);
xnor U28437 (N_28437,N_27945,N_27582);
and U28438 (N_28438,N_27582,N_27728);
nand U28439 (N_28439,N_27827,N_27690);
nand U28440 (N_28440,N_27573,N_27975);
and U28441 (N_28441,N_27725,N_27719);
nor U28442 (N_28442,N_27893,N_27788);
and U28443 (N_28443,N_27555,N_27930);
or U28444 (N_28444,N_27645,N_27860);
nand U28445 (N_28445,N_27752,N_27836);
xnor U28446 (N_28446,N_27902,N_27833);
xnor U28447 (N_28447,N_27880,N_27732);
nor U28448 (N_28448,N_27664,N_27517);
nor U28449 (N_28449,N_27518,N_27610);
xor U28450 (N_28450,N_27998,N_27629);
and U28451 (N_28451,N_27501,N_27897);
or U28452 (N_28452,N_27801,N_27838);
or U28453 (N_28453,N_27636,N_27583);
nand U28454 (N_28454,N_27683,N_27816);
nor U28455 (N_28455,N_27904,N_27559);
nand U28456 (N_28456,N_27518,N_27599);
nor U28457 (N_28457,N_27534,N_27898);
or U28458 (N_28458,N_27751,N_27770);
xnor U28459 (N_28459,N_27683,N_27741);
and U28460 (N_28460,N_27509,N_27628);
and U28461 (N_28461,N_27614,N_27905);
nor U28462 (N_28462,N_27806,N_27612);
nor U28463 (N_28463,N_27554,N_27784);
or U28464 (N_28464,N_27659,N_27676);
or U28465 (N_28465,N_27613,N_27942);
nand U28466 (N_28466,N_27858,N_27640);
or U28467 (N_28467,N_27932,N_27991);
xor U28468 (N_28468,N_27586,N_27541);
and U28469 (N_28469,N_27839,N_27574);
and U28470 (N_28470,N_27873,N_27646);
and U28471 (N_28471,N_27817,N_27994);
or U28472 (N_28472,N_27820,N_27897);
nor U28473 (N_28473,N_27795,N_27802);
and U28474 (N_28474,N_27643,N_27746);
nand U28475 (N_28475,N_27823,N_27781);
or U28476 (N_28476,N_27746,N_27562);
and U28477 (N_28477,N_27673,N_27939);
nand U28478 (N_28478,N_27666,N_27612);
xnor U28479 (N_28479,N_27854,N_27682);
nand U28480 (N_28480,N_27946,N_27925);
nor U28481 (N_28481,N_27855,N_27511);
or U28482 (N_28482,N_27598,N_27739);
or U28483 (N_28483,N_27681,N_27775);
and U28484 (N_28484,N_27620,N_27932);
and U28485 (N_28485,N_27735,N_27990);
or U28486 (N_28486,N_27721,N_27505);
xor U28487 (N_28487,N_27513,N_27567);
nor U28488 (N_28488,N_27549,N_27894);
xor U28489 (N_28489,N_27887,N_27614);
nand U28490 (N_28490,N_27725,N_27990);
and U28491 (N_28491,N_27713,N_27754);
xor U28492 (N_28492,N_27878,N_27698);
or U28493 (N_28493,N_27617,N_27593);
nand U28494 (N_28494,N_27702,N_27546);
and U28495 (N_28495,N_27606,N_27773);
xor U28496 (N_28496,N_27772,N_27750);
xor U28497 (N_28497,N_27802,N_27979);
and U28498 (N_28498,N_27991,N_27579);
or U28499 (N_28499,N_27925,N_27644);
or U28500 (N_28500,N_28389,N_28229);
and U28501 (N_28501,N_28423,N_28155);
and U28502 (N_28502,N_28123,N_28365);
nor U28503 (N_28503,N_28476,N_28428);
xor U28504 (N_28504,N_28493,N_28339);
xor U28505 (N_28505,N_28475,N_28099);
nand U28506 (N_28506,N_28296,N_28289);
or U28507 (N_28507,N_28374,N_28252);
and U28508 (N_28508,N_28120,N_28113);
and U28509 (N_28509,N_28197,N_28304);
or U28510 (N_28510,N_28222,N_28178);
and U28511 (N_28511,N_28175,N_28161);
nand U28512 (N_28512,N_28375,N_28379);
nor U28513 (N_28513,N_28395,N_28025);
or U28514 (N_28514,N_28164,N_28263);
or U28515 (N_28515,N_28497,N_28062);
xnor U28516 (N_28516,N_28118,N_28251);
nor U28517 (N_28517,N_28300,N_28483);
and U28518 (N_28518,N_28442,N_28245);
or U28519 (N_28519,N_28079,N_28176);
and U28520 (N_28520,N_28265,N_28319);
and U28521 (N_28521,N_28171,N_28482);
or U28522 (N_28522,N_28328,N_28186);
xor U28523 (N_28523,N_28202,N_28487);
or U28524 (N_28524,N_28080,N_28443);
nand U28525 (N_28525,N_28354,N_28306);
nand U28526 (N_28526,N_28127,N_28036);
and U28527 (N_28527,N_28139,N_28383);
or U28528 (N_28528,N_28371,N_28077);
and U28529 (N_28529,N_28403,N_28478);
nand U28530 (N_28530,N_28350,N_28149);
and U28531 (N_28531,N_28466,N_28221);
or U28532 (N_28532,N_28064,N_28295);
and U28533 (N_28533,N_28154,N_28089);
nor U28534 (N_28534,N_28187,N_28315);
nand U28535 (N_28535,N_28004,N_28196);
or U28536 (N_28536,N_28013,N_28098);
xnor U28537 (N_28537,N_28220,N_28226);
nor U28538 (N_28538,N_28367,N_28150);
xnor U28539 (N_28539,N_28214,N_28384);
nand U28540 (N_28540,N_28006,N_28405);
or U28541 (N_28541,N_28309,N_28049);
nor U28542 (N_28542,N_28185,N_28358);
nand U28543 (N_28543,N_28461,N_28345);
xor U28544 (N_28544,N_28071,N_28417);
xor U28545 (N_28545,N_28302,N_28067);
nand U28546 (N_28546,N_28000,N_28206);
xnor U28547 (N_28547,N_28451,N_28340);
and U28548 (N_28548,N_28117,N_28361);
and U28549 (N_28549,N_28490,N_28174);
xnor U28550 (N_28550,N_28090,N_28468);
and U28551 (N_28551,N_28420,N_28264);
and U28552 (N_28552,N_28135,N_28136);
nand U28553 (N_28553,N_28437,N_28394);
xor U28554 (N_28554,N_28116,N_28481);
xnor U28555 (N_28555,N_28463,N_28054);
xnor U28556 (N_28556,N_28046,N_28391);
nor U28557 (N_28557,N_28179,N_28285);
nand U28558 (N_28558,N_28128,N_28008);
nand U28559 (N_28559,N_28033,N_28291);
and U28560 (N_28560,N_28147,N_28193);
and U28561 (N_28561,N_28381,N_28242);
nand U28562 (N_28562,N_28275,N_28137);
xnor U28563 (N_28563,N_28070,N_28477);
and U28564 (N_28564,N_28225,N_28172);
nor U28565 (N_28565,N_28249,N_28398);
xor U28566 (N_28566,N_28177,N_28074);
nor U28567 (N_28567,N_28409,N_28396);
nor U28568 (N_28568,N_28218,N_28100);
or U28569 (N_28569,N_28151,N_28452);
or U28570 (N_28570,N_28205,N_28407);
and U28571 (N_28571,N_28125,N_28076);
nor U28572 (N_28572,N_28294,N_28274);
xor U28573 (N_28573,N_28037,N_28278);
and U28574 (N_28574,N_28165,N_28181);
or U28575 (N_28575,N_28105,N_28470);
nand U28576 (N_28576,N_28189,N_28082);
xnor U28577 (N_28577,N_28130,N_28232);
or U28578 (N_28578,N_28126,N_28465);
nor U28579 (N_28579,N_28009,N_28303);
and U28580 (N_28580,N_28329,N_28124);
or U28581 (N_28581,N_28106,N_28019);
xnor U28582 (N_28582,N_28364,N_28342);
and U28583 (N_28583,N_28145,N_28148);
and U28584 (N_28584,N_28208,N_28330);
or U28585 (N_28585,N_28388,N_28455);
xor U28586 (N_28586,N_28489,N_28129);
xnor U28587 (N_28587,N_28401,N_28447);
xor U28588 (N_28588,N_28431,N_28277);
nand U28589 (N_28589,N_28404,N_28439);
nand U28590 (N_28590,N_28132,N_28141);
and U28591 (N_28591,N_28473,N_28093);
and U28592 (N_28592,N_28198,N_28188);
nor U28593 (N_28593,N_28212,N_28380);
nor U28594 (N_28594,N_28469,N_28158);
or U28595 (N_28595,N_28255,N_28491);
xor U28596 (N_28596,N_28430,N_28320);
and U28597 (N_28597,N_28238,N_28485);
xnor U28598 (N_28598,N_28055,N_28387);
xor U28599 (N_28599,N_28030,N_28474);
xor U28600 (N_28600,N_28397,N_28060);
nand U28601 (N_28601,N_28167,N_28183);
nor U28602 (N_28602,N_28168,N_28305);
nor U28603 (N_28603,N_28109,N_28085);
xor U28604 (N_28604,N_28243,N_28163);
and U28605 (N_28605,N_28349,N_28402);
and U28606 (N_28606,N_28337,N_28496);
or U28607 (N_28607,N_28072,N_28194);
or U28608 (N_28608,N_28370,N_28223);
or U28609 (N_28609,N_28338,N_28102);
xnor U28610 (N_28610,N_28026,N_28010);
nand U28611 (N_28611,N_28038,N_28312);
nand U28612 (N_28612,N_28453,N_28484);
nand U28613 (N_28613,N_28399,N_28433);
and U28614 (N_28614,N_28081,N_28107);
nor U28615 (N_28615,N_28419,N_28378);
and U28616 (N_28616,N_28045,N_28007);
nor U28617 (N_28617,N_28173,N_28421);
and U28618 (N_28618,N_28052,N_28084);
nor U28619 (N_28619,N_28040,N_28413);
nand U28620 (N_28620,N_28011,N_28133);
xnor U28621 (N_28621,N_28014,N_28231);
nor U28622 (N_28622,N_28385,N_28230);
nand U28623 (N_28623,N_28311,N_28156);
nor U28624 (N_28624,N_28016,N_28024);
nand U28625 (N_28625,N_28333,N_28299);
or U28626 (N_28626,N_28042,N_28191);
nand U28627 (N_28627,N_28012,N_28101);
nor U28628 (N_28628,N_28348,N_28204);
nand U28629 (N_28629,N_28435,N_28332);
and U28630 (N_28630,N_28362,N_28003);
nand U28631 (N_28631,N_28325,N_28103);
and U28632 (N_28632,N_28495,N_28219);
nand U28633 (N_28633,N_28298,N_28432);
or U28634 (N_28634,N_28351,N_28002);
xnor U28635 (N_28635,N_28180,N_28335);
or U28636 (N_28636,N_28479,N_28170);
and U28637 (N_28637,N_28209,N_28440);
nand U28638 (N_28638,N_28237,N_28044);
nand U28639 (N_28639,N_28261,N_28464);
and U28640 (N_28640,N_28092,N_28005);
nand U28641 (N_28641,N_28454,N_28488);
nor U28642 (N_28642,N_28368,N_28160);
nand U28643 (N_28643,N_28213,N_28039);
and U28644 (N_28644,N_28029,N_28192);
xnor U28645 (N_28645,N_28015,N_28057);
nand U28646 (N_28646,N_28043,N_28363);
or U28647 (N_28647,N_28063,N_28115);
xor U28648 (N_28648,N_28224,N_28075);
and U28649 (N_28649,N_28369,N_28091);
and U28650 (N_28650,N_28246,N_28256);
and U28651 (N_28651,N_28492,N_28022);
and U28652 (N_28652,N_28324,N_28462);
nand U28653 (N_28653,N_28244,N_28269);
nand U28654 (N_28654,N_28459,N_28310);
or U28655 (N_28655,N_28271,N_28408);
or U28656 (N_28656,N_28414,N_28283);
nand U28657 (N_28657,N_28078,N_28112);
or U28658 (N_28658,N_28086,N_28235);
xnor U28659 (N_28659,N_28058,N_28066);
nand U28660 (N_28660,N_28153,N_28096);
and U28661 (N_28661,N_28216,N_28434);
xnor U28662 (N_28662,N_28211,N_28203);
and U28663 (N_28663,N_28281,N_28157);
nor U28664 (N_28664,N_28422,N_28268);
xnor U28665 (N_28665,N_28288,N_28047);
nand U28666 (N_28666,N_28190,N_28450);
or U28667 (N_28667,N_28053,N_28201);
or U28668 (N_28668,N_28210,N_28142);
nand U28669 (N_28669,N_28448,N_28144);
nor U28670 (N_28670,N_28444,N_28331);
or U28671 (N_28671,N_28486,N_28138);
nand U28672 (N_28672,N_28095,N_28429);
or U28673 (N_28673,N_28457,N_28286);
nor U28674 (N_28674,N_28412,N_28334);
nand U28675 (N_28675,N_28111,N_28146);
nand U28676 (N_28676,N_28114,N_28480);
nand U28677 (N_28677,N_28366,N_28284);
nand U28678 (N_28678,N_28023,N_28356);
nor U28679 (N_28679,N_28438,N_28327);
and U28680 (N_28680,N_28313,N_28292);
nor U28681 (N_28681,N_28262,N_28272);
nor U28682 (N_28682,N_28372,N_28377);
and U28683 (N_28683,N_28217,N_28241);
nor U28684 (N_28684,N_28359,N_28276);
xor U28685 (N_28685,N_28050,N_28360);
nand U28686 (N_28686,N_28131,N_28068);
xor U28687 (N_28687,N_28498,N_28104);
nand U28688 (N_28688,N_28207,N_28234);
xor U28689 (N_28689,N_28456,N_28308);
xnor U28690 (N_28690,N_28343,N_28254);
and U28691 (N_28691,N_28460,N_28441);
and U28692 (N_28692,N_28357,N_28406);
or U28693 (N_28693,N_28088,N_28400);
nor U28694 (N_28694,N_28065,N_28425);
xnor U28695 (N_28695,N_28059,N_28471);
nand U28696 (N_28696,N_28228,N_28236);
nand U28697 (N_28697,N_28083,N_28307);
nor U28698 (N_28698,N_28373,N_28073);
nand U28699 (N_28699,N_28032,N_28346);
or U28700 (N_28700,N_28411,N_28184);
and U28701 (N_28701,N_28250,N_28143);
and U28702 (N_28702,N_28031,N_28240);
xnor U28703 (N_28703,N_28341,N_28494);
nand U28704 (N_28704,N_28445,N_28293);
or U28705 (N_28705,N_28110,N_28258);
nand U28706 (N_28706,N_28270,N_28227);
nand U28707 (N_28707,N_28027,N_28467);
or U28708 (N_28708,N_28041,N_28061);
nand U28709 (N_28709,N_28169,N_28318);
nand U28710 (N_28710,N_28035,N_28248);
xnor U28711 (N_28711,N_28094,N_28200);
or U28712 (N_28712,N_28314,N_28215);
and U28713 (N_28713,N_28162,N_28279);
nand U28714 (N_28714,N_28233,N_28287);
nor U28715 (N_28715,N_28069,N_28087);
and U28716 (N_28716,N_28273,N_28376);
nand U28717 (N_28717,N_28048,N_28166);
nand U28718 (N_28718,N_28119,N_28056);
xor U28719 (N_28719,N_28321,N_28028);
and U28720 (N_28720,N_28247,N_28436);
xnor U28721 (N_28721,N_28257,N_28122);
nor U28722 (N_28722,N_28317,N_28382);
and U28723 (N_28723,N_28446,N_28410);
nor U28724 (N_28724,N_28297,N_28018);
and U28725 (N_28725,N_28472,N_28449);
nor U28726 (N_28726,N_28239,N_28393);
nor U28727 (N_28727,N_28282,N_28280);
xnor U28728 (N_28728,N_28108,N_28424);
nand U28729 (N_28729,N_28458,N_28353);
nor U28730 (N_28730,N_28195,N_28097);
xor U28731 (N_28731,N_28426,N_28355);
and U28732 (N_28732,N_28352,N_28416);
nor U28733 (N_28733,N_28322,N_28499);
or U28734 (N_28734,N_28347,N_28017);
or U28735 (N_28735,N_28415,N_28386);
or U28736 (N_28736,N_28323,N_28134);
and U28737 (N_28737,N_28140,N_28427);
or U28738 (N_28738,N_28267,N_28253);
and U28739 (N_28739,N_28034,N_28121);
or U28740 (N_28740,N_28051,N_28316);
xnor U28741 (N_28741,N_28021,N_28392);
nand U28742 (N_28742,N_28418,N_28344);
or U28743 (N_28743,N_28290,N_28259);
or U28744 (N_28744,N_28159,N_28152);
and U28745 (N_28745,N_28390,N_28260);
xnor U28746 (N_28746,N_28199,N_28001);
or U28747 (N_28747,N_28266,N_28336);
and U28748 (N_28748,N_28301,N_28020);
or U28749 (N_28749,N_28326,N_28182);
or U28750 (N_28750,N_28475,N_28153);
and U28751 (N_28751,N_28321,N_28113);
and U28752 (N_28752,N_28202,N_28408);
and U28753 (N_28753,N_28363,N_28068);
and U28754 (N_28754,N_28082,N_28335);
nand U28755 (N_28755,N_28032,N_28195);
or U28756 (N_28756,N_28286,N_28111);
xor U28757 (N_28757,N_28047,N_28390);
and U28758 (N_28758,N_28004,N_28014);
or U28759 (N_28759,N_28425,N_28145);
nand U28760 (N_28760,N_28449,N_28193);
xnor U28761 (N_28761,N_28478,N_28017);
nor U28762 (N_28762,N_28462,N_28192);
and U28763 (N_28763,N_28490,N_28477);
nand U28764 (N_28764,N_28135,N_28433);
nand U28765 (N_28765,N_28273,N_28133);
and U28766 (N_28766,N_28474,N_28072);
or U28767 (N_28767,N_28330,N_28425);
xor U28768 (N_28768,N_28093,N_28261);
xnor U28769 (N_28769,N_28414,N_28194);
and U28770 (N_28770,N_28146,N_28268);
xor U28771 (N_28771,N_28068,N_28013);
and U28772 (N_28772,N_28242,N_28180);
and U28773 (N_28773,N_28489,N_28230);
nor U28774 (N_28774,N_28234,N_28324);
and U28775 (N_28775,N_28000,N_28374);
nand U28776 (N_28776,N_28428,N_28103);
xnor U28777 (N_28777,N_28159,N_28093);
nor U28778 (N_28778,N_28461,N_28036);
or U28779 (N_28779,N_28303,N_28324);
and U28780 (N_28780,N_28412,N_28290);
nor U28781 (N_28781,N_28096,N_28137);
xnor U28782 (N_28782,N_28349,N_28203);
or U28783 (N_28783,N_28455,N_28252);
and U28784 (N_28784,N_28149,N_28398);
and U28785 (N_28785,N_28071,N_28234);
nand U28786 (N_28786,N_28005,N_28187);
xnor U28787 (N_28787,N_28038,N_28107);
or U28788 (N_28788,N_28384,N_28281);
nand U28789 (N_28789,N_28344,N_28369);
nand U28790 (N_28790,N_28129,N_28325);
nor U28791 (N_28791,N_28046,N_28435);
xnor U28792 (N_28792,N_28397,N_28200);
or U28793 (N_28793,N_28495,N_28313);
and U28794 (N_28794,N_28371,N_28189);
xnor U28795 (N_28795,N_28101,N_28158);
nor U28796 (N_28796,N_28026,N_28294);
nand U28797 (N_28797,N_28082,N_28331);
nor U28798 (N_28798,N_28309,N_28313);
xor U28799 (N_28799,N_28101,N_28496);
xor U28800 (N_28800,N_28429,N_28006);
nor U28801 (N_28801,N_28307,N_28292);
xnor U28802 (N_28802,N_28008,N_28195);
or U28803 (N_28803,N_28132,N_28337);
and U28804 (N_28804,N_28299,N_28195);
and U28805 (N_28805,N_28436,N_28392);
nor U28806 (N_28806,N_28293,N_28335);
xor U28807 (N_28807,N_28252,N_28326);
and U28808 (N_28808,N_28051,N_28081);
and U28809 (N_28809,N_28412,N_28402);
nor U28810 (N_28810,N_28160,N_28404);
and U28811 (N_28811,N_28072,N_28425);
nand U28812 (N_28812,N_28129,N_28341);
xor U28813 (N_28813,N_28268,N_28092);
or U28814 (N_28814,N_28077,N_28091);
nor U28815 (N_28815,N_28092,N_28458);
nor U28816 (N_28816,N_28332,N_28066);
xor U28817 (N_28817,N_28110,N_28045);
and U28818 (N_28818,N_28039,N_28146);
or U28819 (N_28819,N_28271,N_28494);
or U28820 (N_28820,N_28484,N_28078);
or U28821 (N_28821,N_28351,N_28181);
nand U28822 (N_28822,N_28406,N_28193);
nor U28823 (N_28823,N_28134,N_28023);
xnor U28824 (N_28824,N_28160,N_28039);
or U28825 (N_28825,N_28237,N_28092);
and U28826 (N_28826,N_28369,N_28028);
xor U28827 (N_28827,N_28382,N_28402);
nor U28828 (N_28828,N_28189,N_28304);
xor U28829 (N_28829,N_28321,N_28453);
or U28830 (N_28830,N_28135,N_28037);
or U28831 (N_28831,N_28311,N_28009);
xor U28832 (N_28832,N_28354,N_28099);
and U28833 (N_28833,N_28022,N_28456);
or U28834 (N_28834,N_28342,N_28325);
xor U28835 (N_28835,N_28082,N_28030);
or U28836 (N_28836,N_28389,N_28364);
nor U28837 (N_28837,N_28484,N_28065);
or U28838 (N_28838,N_28088,N_28385);
nor U28839 (N_28839,N_28303,N_28449);
nand U28840 (N_28840,N_28400,N_28050);
nand U28841 (N_28841,N_28036,N_28465);
and U28842 (N_28842,N_28213,N_28248);
xnor U28843 (N_28843,N_28394,N_28315);
and U28844 (N_28844,N_28027,N_28389);
nand U28845 (N_28845,N_28173,N_28003);
xor U28846 (N_28846,N_28466,N_28254);
nand U28847 (N_28847,N_28009,N_28146);
xnor U28848 (N_28848,N_28381,N_28478);
nor U28849 (N_28849,N_28456,N_28228);
xor U28850 (N_28850,N_28090,N_28009);
xnor U28851 (N_28851,N_28483,N_28399);
and U28852 (N_28852,N_28018,N_28471);
xor U28853 (N_28853,N_28458,N_28234);
or U28854 (N_28854,N_28344,N_28333);
nand U28855 (N_28855,N_28042,N_28159);
nand U28856 (N_28856,N_28377,N_28031);
and U28857 (N_28857,N_28042,N_28351);
and U28858 (N_28858,N_28431,N_28424);
nor U28859 (N_28859,N_28101,N_28069);
nor U28860 (N_28860,N_28496,N_28222);
or U28861 (N_28861,N_28313,N_28421);
nor U28862 (N_28862,N_28159,N_28395);
or U28863 (N_28863,N_28020,N_28259);
xor U28864 (N_28864,N_28338,N_28043);
and U28865 (N_28865,N_28427,N_28337);
and U28866 (N_28866,N_28052,N_28158);
and U28867 (N_28867,N_28259,N_28191);
and U28868 (N_28868,N_28142,N_28059);
xnor U28869 (N_28869,N_28405,N_28027);
xor U28870 (N_28870,N_28257,N_28020);
nand U28871 (N_28871,N_28058,N_28345);
nor U28872 (N_28872,N_28181,N_28226);
nand U28873 (N_28873,N_28004,N_28430);
xor U28874 (N_28874,N_28117,N_28456);
nor U28875 (N_28875,N_28105,N_28295);
xnor U28876 (N_28876,N_28237,N_28283);
xor U28877 (N_28877,N_28272,N_28486);
nand U28878 (N_28878,N_28126,N_28430);
and U28879 (N_28879,N_28258,N_28208);
xor U28880 (N_28880,N_28488,N_28222);
xor U28881 (N_28881,N_28052,N_28431);
nor U28882 (N_28882,N_28394,N_28368);
xnor U28883 (N_28883,N_28451,N_28337);
or U28884 (N_28884,N_28474,N_28286);
or U28885 (N_28885,N_28013,N_28080);
nor U28886 (N_28886,N_28495,N_28442);
or U28887 (N_28887,N_28247,N_28468);
or U28888 (N_28888,N_28424,N_28420);
and U28889 (N_28889,N_28489,N_28261);
xor U28890 (N_28890,N_28060,N_28076);
or U28891 (N_28891,N_28317,N_28183);
nand U28892 (N_28892,N_28427,N_28280);
nand U28893 (N_28893,N_28283,N_28304);
or U28894 (N_28894,N_28288,N_28380);
and U28895 (N_28895,N_28485,N_28023);
or U28896 (N_28896,N_28406,N_28142);
or U28897 (N_28897,N_28387,N_28316);
and U28898 (N_28898,N_28259,N_28294);
nand U28899 (N_28899,N_28241,N_28055);
xor U28900 (N_28900,N_28471,N_28429);
nor U28901 (N_28901,N_28095,N_28056);
nand U28902 (N_28902,N_28140,N_28370);
nand U28903 (N_28903,N_28253,N_28234);
or U28904 (N_28904,N_28482,N_28011);
and U28905 (N_28905,N_28299,N_28144);
and U28906 (N_28906,N_28448,N_28238);
and U28907 (N_28907,N_28009,N_28111);
nand U28908 (N_28908,N_28114,N_28204);
and U28909 (N_28909,N_28239,N_28222);
nor U28910 (N_28910,N_28342,N_28447);
and U28911 (N_28911,N_28141,N_28073);
xor U28912 (N_28912,N_28117,N_28400);
or U28913 (N_28913,N_28465,N_28345);
nand U28914 (N_28914,N_28097,N_28011);
xor U28915 (N_28915,N_28285,N_28472);
nor U28916 (N_28916,N_28346,N_28285);
or U28917 (N_28917,N_28274,N_28096);
xor U28918 (N_28918,N_28300,N_28422);
xnor U28919 (N_28919,N_28309,N_28134);
nand U28920 (N_28920,N_28245,N_28286);
and U28921 (N_28921,N_28401,N_28263);
nand U28922 (N_28922,N_28287,N_28359);
nand U28923 (N_28923,N_28475,N_28143);
and U28924 (N_28924,N_28457,N_28493);
or U28925 (N_28925,N_28095,N_28491);
nand U28926 (N_28926,N_28022,N_28309);
and U28927 (N_28927,N_28498,N_28268);
nand U28928 (N_28928,N_28137,N_28054);
xnor U28929 (N_28929,N_28087,N_28013);
and U28930 (N_28930,N_28142,N_28420);
xor U28931 (N_28931,N_28318,N_28218);
nor U28932 (N_28932,N_28236,N_28168);
xor U28933 (N_28933,N_28486,N_28251);
nand U28934 (N_28934,N_28266,N_28355);
and U28935 (N_28935,N_28297,N_28004);
nand U28936 (N_28936,N_28345,N_28294);
nand U28937 (N_28937,N_28122,N_28386);
and U28938 (N_28938,N_28330,N_28072);
nand U28939 (N_28939,N_28459,N_28335);
nor U28940 (N_28940,N_28293,N_28298);
or U28941 (N_28941,N_28494,N_28380);
and U28942 (N_28942,N_28299,N_28445);
nand U28943 (N_28943,N_28007,N_28419);
or U28944 (N_28944,N_28433,N_28218);
and U28945 (N_28945,N_28492,N_28379);
and U28946 (N_28946,N_28145,N_28063);
and U28947 (N_28947,N_28281,N_28117);
and U28948 (N_28948,N_28367,N_28328);
nor U28949 (N_28949,N_28464,N_28458);
and U28950 (N_28950,N_28446,N_28467);
nor U28951 (N_28951,N_28069,N_28466);
nand U28952 (N_28952,N_28165,N_28029);
or U28953 (N_28953,N_28132,N_28490);
or U28954 (N_28954,N_28196,N_28012);
nor U28955 (N_28955,N_28080,N_28120);
nand U28956 (N_28956,N_28074,N_28358);
or U28957 (N_28957,N_28322,N_28013);
and U28958 (N_28958,N_28405,N_28018);
or U28959 (N_28959,N_28047,N_28377);
nand U28960 (N_28960,N_28304,N_28047);
or U28961 (N_28961,N_28231,N_28140);
xor U28962 (N_28962,N_28200,N_28315);
and U28963 (N_28963,N_28024,N_28296);
nor U28964 (N_28964,N_28165,N_28477);
or U28965 (N_28965,N_28301,N_28348);
nor U28966 (N_28966,N_28225,N_28265);
xor U28967 (N_28967,N_28298,N_28103);
xnor U28968 (N_28968,N_28128,N_28235);
or U28969 (N_28969,N_28448,N_28478);
nand U28970 (N_28970,N_28052,N_28388);
xor U28971 (N_28971,N_28421,N_28384);
nand U28972 (N_28972,N_28330,N_28477);
xnor U28973 (N_28973,N_28094,N_28240);
nand U28974 (N_28974,N_28064,N_28169);
nand U28975 (N_28975,N_28104,N_28112);
nand U28976 (N_28976,N_28396,N_28203);
or U28977 (N_28977,N_28388,N_28192);
xnor U28978 (N_28978,N_28092,N_28011);
xnor U28979 (N_28979,N_28326,N_28186);
and U28980 (N_28980,N_28247,N_28365);
nand U28981 (N_28981,N_28472,N_28138);
and U28982 (N_28982,N_28165,N_28360);
xnor U28983 (N_28983,N_28039,N_28448);
or U28984 (N_28984,N_28334,N_28000);
nor U28985 (N_28985,N_28380,N_28255);
and U28986 (N_28986,N_28231,N_28253);
nor U28987 (N_28987,N_28000,N_28104);
or U28988 (N_28988,N_28298,N_28056);
nor U28989 (N_28989,N_28306,N_28466);
or U28990 (N_28990,N_28015,N_28229);
nand U28991 (N_28991,N_28062,N_28498);
nor U28992 (N_28992,N_28483,N_28144);
nor U28993 (N_28993,N_28039,N_28144);
xnor U28994 (N_28994,N_28153,N_28355);
nor U28995 (N_28995,N_28474,N_28400);
xor U28996 (N_28996,N_28245,N_28347);
and U28997 (N_28997,N_28363,N_28489);
nor U28998 (N_28998,N_28057,N_28187);
nand U28999 (N_28999,N_28344,N_28297);
nand U29000 (N_29000,N_28861,N_28934);
nand U29001 (N_29001,N_28613,N_28672);
or U29002 (N_29002,N_28572,N_28587);
xor U29003 (N_29003,N_28599,N_28836);
nand U29004 (N_29004,N_28778,N_28524);
and U29005 (N_29005,N_28787,N_28841);
nand U29006 (N_29006,N_28842,N_28800);
or U29007 (N_29007,N_28973,N_28707);
nand U29008 (N_29008,N_28550,N_28630);
or U29009 (N_29009,N_28935,N_28968);
and U29010 (N_29010,N_28768,N_28575);
or U29011 (N_29011,N_28795,N_28728);
nor U29012 (N_29012,N_28737,N_28964);
or U29013 (N_29013,N_28516,N_28771);
and U29014 (N_29014,N_28643,N_28555);
nand U29015 (N_29015,N_28634,N_28849);
or U29016 (N_29016,N_28767,N_28826);
and U29017 (N_29017,N_28945,N_28981);
nand U29018 (N_29018,N_28631,N_28902);
or U29019 (N_29019,N_28678,N_28822);
nand U29020 (N_29020,N_28788,N_28511);
nand U29021 (N_29021,N_28546,N_28824);
nand U29022 (N_29022,N_28651,N_28814);
and U29023 (N_29023,N_28662,N_28556);
nand U29024 (N_29024,N_28884,N_28959);
nor U29025 (N_29025,N_28649,N_28586);
xnor U29026 (N_29026,N_28920,N_28505);
or U29027 (N_29027,N_28834,N_28817);
and U29028 (N_29028,N_28855,N_28900);
or U29029 (N_29029,N_28607,N_28986);
nor U29030 (N_29030,N_28705,N_28847);
or U29031 (N_29031,N_28955,N_28763);
xnor U29032 (N_29032,N_28840,N_28574);
and U29033 (N_29033,N_28815,N_28681);
nand U29034 (N_29034,N_28548,N_28999);
nor U29035 (N_29035,N_28682,N_28960);
or U29036 (N_29036,N_28906,N_28914);
and U29037 (N_29037,N_28510,N_28989);
or U29038 (N_29038,N_28828,N_28932);
and U29039 (N_29039,N_28810,N_28615);
nand U29040 (N_29040,N_28988,N_28928);
nor U29041 (N_29041,N_28532,N_28783);
or U29042 (N_29042,N_28896,N_28868);
nand U29043 (N_29043,N_28564,N_28991);
xnor U29044 (N_29044,N_28673,N_28745);
and U29045 (N_29045,N_28936,N_28612);
nor U29046 (N_29046,N_28957,N_28799);
nor U29047 (N_29047,N_28692,N_28791);
xnor U29048 (N_29048,N_28753,N_28854);
nor U29049 (N_29049,N_28725,N_28541);
xnor U29050 (N_29050,N_28679,N_28579);
or U29051 (N_29051,N_28827,N_28605);
or U29052 (N_29052,N_28898,N_28711);
and U29053 (N_29053,N_28503,N_28669);
xnor U29054 (N_29054,N_28978,N_28773);
or U29055 (N_29055,N_28919,N_28632);
or U29056 (N_29056,N_28829,N_28922);
or U29057 (N_29057,N_28859,N_28891);
xor U29058 (N_29058,N_28723,N_28789);
xnor U29059 (N_29059,N_28812,N_28543);
nand U29060 (N_29060,N_28941,N_28816);
and U29061 (N_29061,N_28576,N_28756);
nor U29062 (N_29062,N_28916,N_28562);
nor U29063 (N_29063,N_28622,N_28736);
nand U29064 (N_29064,N_28966,N_28792);
and U29065 (N_29065,N_28538,N_28862);
and U29066 (N_29066,N_28933,N_28685);
nor U29067 (N_29067,N_28923,N_28545);
xor U29068 (N_29068,N_28596,N_28666);
or U29069 (N_29069,N_28608,N_28754);
xnor U29070 (N_29070,N_28734,N_28990);
and U29071 (N_29071,N_28652,N_28888);
and U29072 (N_29072,N_28851,N_28775);
or U29073 (N_29073,N_28832,N_28878);
and U29074 (N_29074,N_28951,N_28602);
nand U29075 (N_29075,N_28716,N_28501);
nand U29076 (N_29076,N_28794,N_28589);
and U29077 (N_29077,N_28948,N_28915);
and U29078 (N_29078,N_28944,N_28709);
or U29079 (N_29079,N_28907,N_28661);
and U29080 (N_29080,N_28701,N_28595);
xor U29081 (N_29081,N_28869,N_28557);
nand U29082 (N_29082,N_28648,N_28542);
or U29083 (N_29083,N_28731,N_28887);
and U29084 (N_29084,N_28639,N_28680);
xor U29085 (N_29085,N_28890,N_28979);
nor U29086 (N_29086,N_28885,N_28997);
nor U29087 (N_29087,N_28982,N_28593);
or U29088 (N_29088,N_28892,N_28558);
xor U29089 (N_29089,N_28894,N_28950);
xnor U29090 (N_29090,N_28813,N_28582);
or U29091 (N_29091,N_28811,N_28526);
nand U29092 (N_29092,N_28808,N_28947);
or U29093 (N_29093,N_28688,N_28764);
nor U29094 (N_29094,N_28702,N_28925);
nor U29095 (N_29095,N_28867,N_28893);
and U29096 (N_29096,N_28797,N_28715);
nor U29097 (N_29097,N_28949,N_28776);
or U29098 (N_29098,N_28659,N_28926);
and U29099 (N_29099,N_28992,N_28706);
nor U29100 (N_29100,N_28909,N_28831);
xor U29101 (N_29101,N_28600,N_28694);
nand U29102 (N_29102,N_28803,N_28606);
nor U29103 (N_29103,N_28905,N_28638);
nand U29104 (N_29104,N_28735,N_28512);
xor U29105 (N_29105,N_28712,N_28645);
or U29106 (N_29106,N_28500,N_28640);
nand U29107 (N_29107,N_28618,N_28874);
or U29108 (N_29108,N_28835,N_28713);
or U29109 (N_29109,N_28647,N_28858);
nor U29110 (N_29110,N_28762,N_28969);
nand U29111 (N_29111,N_28733,N_28523);
nand U29112 (N_29112,N_28721,N_28561);
nor U29113 (N_29113,N_28780,N_28646);
nor U29114 (N_29114,N_28747,N_28995);
xnor U29115 (N_29115,N_28876,N_28588);
nand U29116 (N_29116,N_28838,N_28863);
nand U29117 (N_29117,N_28961,N_28577);
xor U29118 (N_29118,N_28509,N_28720);
xor U29119 (N_29119,N_28683,N_28703);
xor U29120 (N_29120,N_28807,N_28921);
nand U29121 (N_29121,N_28774,N_28937);
nor U29122 (N_29122,N_28751,N_28998);
xor U29123 (N_29123,N_28617,N_28690);
nand U29124 (N_29124,N_28585,N_28625);
and U29125 (N_29125,N_28598,N_28530);
xor U29126 (N_29126,N_28603,N_28879);
nand U29127 (N_29127,N_28660,N_28857);
nor U29128 (N_29128,N_28856,N_28699);
nand U29129 (N_29129,N_28686,N_28633);
or U29130 (N_29130,N_28676,N_28804);
or U29131 (N_29131,N_28663,N_28977);
and U29132 (N_29132,N_28980,N_28805);
or U29133 (N_29133,N_28758,N_28962);
nor U29134 (N_29134,N_28818,N_28552);
nor U29135 (N_29135,N_28954,N_28529);
and U29136 (N_29136,N_28965,N_28899);
or U29137 (N_29137,N_28744,N_28740);
nand U29138 (N_29138,N_28996,N_28580);
nor U29139 (N_29139,N_28677,N_28761);
nor U29140 (N_29140,N_28729,N_28940);
nand U29141 (N_29141,N_28911,N_28809);
nor U29142 (N_29142,N_28924,N_28504);
and U29143 (N_29143,N_28777,N_28877);
xnor U29144 (N_29144,N_28732,N_28850);
or U29145 (N_29145,N_28637,N_28704);
nor U29146 (N_29146,N_28687,N_28974);
and U29147 (N_29147,N_28913,N_28938);
nor U29148 (N_29148,N_28628,N_28522);
xor U29149 (N_29149,N_28819,N_28908);
or U29150 (N_29150,N_28570,N_28722);
nor U29151 (N_29151,N_28514,N_28782);
nor U29152 (N_29152,N_28616,N_28527);
xnor U29153 (N_29153,N_28971,N_28610);
and U29154 (N_29154,N_28802,N_28569);
xnor U29155 (N_29155,N_28536,N_28627);
xnor U29156 (N_29156,N_28943,N_28671);
nor U29157 (N_29157,N_28693,N_28845);
and U29158 (N_29158,N_28881,N_28895);
xnor U29159 (N_29159,N_28567,N_28931);
nor U29160 (N_29160,N_28853,N_28559);
nand U29161 (N_29161,N_28691,N_28953);
nor U29162 (N_29162,N_28549,N_28785);
and U29163 (N_29163,N_28872,N_28551);
nor U29164 (N_29164,N_28903,N_28970);
nor U29165 (N_29165,N_28942,N_28609);
xor U29166 (N_29166,N_28604,N_28621);
nand U29167 (N_29167,N_28654,N_28619);
nor U29168 (N_29168,N_28535,N_28518);
xor U29169 (N_29169,N_28839,N_28972);
xor U29170 (N_29170,N_28502,N_28848);
xor U29171 (N_29171,N_28963,N_28865);
nand U29172 (N_29172,N_28650,N_28620);
xor U29173 (N_29173,N_28823,N_28852);
nand U29174 (N_29174,N_28870,N_28521);
nor U29175 (N_29175,N_28750,N_28743);
xnor U29176 (N_29176,N_28539,N_28506);
xnor U29177 (N_29177,N_28533,N_28741);
nand U29178 (N_29178,N_28667,N_28581);
xor U29179 (N_29179,N_28519,N_28565);
or U29180 (N_29180,N_28821,N_28748);
and U29181 (N_29181,N_28534,N_28846);
or U29182 (N_29182,N_28752,N_28742);
and U29183 (N_29183,N_28718,N_28994);
xor U29184 (N_29184,N_28584,N_28985);
or U29185 (N_29185,N_28636,N_28784);
xnor U29186 (N_29186,N_28563,N_28657);
nand U29187 (N_29187,N_28554,N_28537);
nand U29188 (N_29188,N_28871,N_28730);
xor U29189 (N_29189,N_28675,N_28515);
nor U29190 (N_29190,N_28528,N_28553);
nor U29191 (N_29191,N_28765,N_28635);
nand U29192 (N_29192,N_28525,N_28844);
nor U29193 (N_29193,N_28904,N_28983);
xnor U29194 (N_29194,N_28611,N_28755);
or U29195 (N_29195,N_28873,N_28719);
xor U29196 (N_29196,N_28798,N_28759);
nand U29197 (N_29197,N_28739,N_28967);
or U29198 (N_29198,N_28674,N_28830);
and U29199 (N_29199,N_28594,N_28837);
and U29200 (N_29200,N_28927,N_28781);
and U29201 (N_29201,N_28513,N_28626);
xor U29202 (N_29202,N_28749,N_28930);
and U29203 (N_29203,N_28708,N_28727);
xnor U29204 (N_29204,N_28843,N_28786);
nand U29205 (N_29205,N_28958,N_28629);
xor U29206 (N_29206,N_28623,N_28658);
nor U29207 (N_29207,N_28770,N_28917);
nand U29208 (N_29208,N_28897,N_28641);
and U29209 (N_29209,N_28939,N_28796);
or U29210 (N_29210,N_28772,N_28790);
xor U29211 (N_29211,N_28698,N_28726);
or U29212 (N_29212,N_28724,N_28757);
and U29213 (N_29213,N_28882,N_28987);
nor U29214 (N_29214,N_28624,N_28910);
and U29215 (N_29215,N_28929,N_28520);
or U29216 (N_29216,N_28668,N_28825);
or U29217 (N_29217,N_28540,N_28653);
nor U29218 (N_29218,N_28566,N_28591);
nand U29219 (N_29219,N_28597,N_28665);
xnor U29220 (N_29220,N_28889,N_28573);
xor U29221 (N_29221,N_28614,N_28695);
or U29222 (N_29222,N_28993,N_28544);
xnor U29223 (N_29223,N_28766,N_28578);
xnor U29224 (N_29224,N_28601,N_28912);
nand U29225 (N_29225,N_28684,N_28866);
or U29226 (N_29226,N_28714,N_28689);
nor U29227 (N_29227,N_28901,N_28655);
nand U29228 (N_29228,N_28801,N_28590);
and U29229 (N_29229,N_28976,N_28571);
nor U29230 (N_29230,N_28508,N_28746);
xnor U29231 (N_29231,N_28779,N_28517);
nor U29232 (N_29232,N_28880,N_28717);
xor U29233 (N_29233,N_28697,N_28700);
and U29234 (N_29234,N_28860,N_28760);
nand U29235 (N_29235,N_28531,N_28656);
xnor U29236 (N_29236,N_28583,N_28875);
and U29237 (N_29237,N_28886,N_28664);
nor U29238 (N_29238,N_28952,N_28644);
nor U29239 (N_29239,N_28738,N_28806);
xnor U29240 (N_29240,N_28975,N_28864);
nor U29241 (N_29241,N_28820,N_28883);
and U29242 (N_29242,N_28769,N_28547);
nand U29243 (N_29243,N_28833,N_28946);
nand U29244 (N_29244,N_28710,N_28670);
nor U29245 (N_29245,N_28984,N_28918);
and U29246 (N_29246,N_28696,N_28568);
nand U29247 (N_29247,N_28507,N_28560);
or U29248 (N_29248,N_28592,N_28642);
nand U29249 (N_29249,N_28956,N_28793);
nand U29250 (N_29250,N_28545,N_28577);
or U29251 (N_29251,N_28672,N_28886);
xor U29252 (N_29252,N_28521,N_28654);
and U29253 (N_29253,N_28554,N_28747);
or U29254 (N_29254,N_28891,N_28763);
or U29255 (N_29255,N_28718,N_28991);
or U29256 (N_29256,N_28809,N_28650);
nor U29257 (N_29257,N_28900,N_28670);
nor U29258 (N_29258,N_28636,N_28890);
or U29259 (N_29259,N_28628,N_28826);
xor U29260 (N_29260,N_28533,N_28838);
nand U29261 (N_29261,N_28508,N_28694);
and U29262 (N_29262,N_28597,N_28810);
and U29263 (N_29263,N_28710,N_28599);
or U29264 (N_29264,N_28819,N_28729);
xnor U29265 (N_29265,N_28804,N_28520);
nor U29266 (N_29266,N_28762,N_28866);
xor U29267 (N_29267,N_28807,N_28992);
nor U29268 (N_29268,N_28805,N_28920);
nor U29269 (N_29269,N_28509,N_28569);
and U29270 (N_29270,N_28928,N_28649);
and U29271 (N_29271,N_28829,N_28670);
or U29272 (N_29272,N_28572,N_28641);
nor U29273 (N_29273,N_28728,N_28763);
and U29274 (N_29274,N_28592,N_28509);
nand U29275 (N_29275,N_28761,N_28826);
nand U29276 (N_29276,N_28633,N_28688);
or U29277 (N_29277,N_28603,N_28634);
nand U29278 (N_29278,N_28720,N_28760);
and U29279 (N_29279,N_28753,N_28926);
or U29280 (N_29280,N_28863,N_28538);
and U29281 (N_29281,N_28653,N_28982);
nor U29282 (N_29282,N_28658,N_28818);
and U29283 (N_29283,N_28730,N_28985);
nand U29284 (N_29284,N_28886,N_28520);
nand U29285 (N_29285,N_28651,N_28801);
and U29286 (N_29286,N_28642,N_28846);
nand U29287 (N_29287,N_28745,N_28621);
and U29288 (N_29288,N_28907,N_28762);
xor U29289 (N_29289,N_28666,N_28521);
nor U29290 (N_29290,N_28598,N_28827);
and U29291 (N_29291,N_28709,N_28553);
nand U29292 (N_29292,N_28677,N_28989);
nand U29293 (N_29293,N_28595,N_28918);
nor U29294 (N_29294,N_28943,N_28867);
and U29295 (N_29295,N_28621,N_28832);
nor U29296 (N_29296,N_28734,N_28660);
nand U29297 (N_29297,N_28527,N_28757);
or U29298 (N_29298,N_28793,N_28991);
nand U29299 (N_29299,N_28687,N_28813);
nand U29300 (N_29300,N_28672,N_28955);
xor U29301 (N_29301,N_28518,N_28612);
or U29302 (N_29302,N_28914,N_28872);
nor U29303 (N_29303,N_28835,N_28766);
or U29304 (N_29304,N_28954,N_28595);
xnor U29305 (N_29305,N_28925,N_28893);
and U29306 (N_29306,N_28700,N_28888);
or U29307 (N_29307,N_28889,N_28941);
nor U29308 (N_29308,N_28609,N_28973);
or U29309 (N_29309,N_28767,N_28910);
and U29310 (N_29310,N_28826,N_28969);
nand U29311 (N_29311,N_28826,N_28697);
nand U29312 (N_29312,N_28883,N_28894);
xor U29313 (N_29313,N_28775,N_28761);
and U29314 (N_29314,N_28695,N_28938);
xor U29315 (N_29315,N_28893,N_28990);
nand U29316 (N_29316,N_28793,N_28518);
nor U29317 (N_29317,N_28546,N_28613);
nand U29318 (N_29318,N_28913,N_28663);
or U29319 (N_29319,N_28656,N_28714);
and U29320 (N_29320,N_28868,N_28899);
nand U29321 (N_29321,N_28807,N_28869);
xor U29322 (N_29322,N_28620,N_28804);
nor U29323 (N_29323,N_28548,N_28748);
and U29324 (N_29324,N_28884,N_28908);
or U29325 (N_29325,N_28976,N_28540);
or U29326 (N_29326,N_28674,N_28533);
nor U29327 (N_29327,N_28524,N_28689);
or U29328 (N_29328,N_28535,N_28531);
and U29329 (N_29329,N_28767,N_28523);
nand U29330 (N_29330,N_28504,N_28925);
nor U29331 (N_29331,N_28693,N_28799);
or U29332 (N_29332,N_28641,N_28611);
nand U29333 (N_29333,N_28893,N_28550);
or U29334 (N_29334,N_28806,N_28883);
xnor U29335 (N_29335,N_28740,N_28629);
nor U29336 (N_29336,N_28737,N_28910);
nand U29337 (N_29337,N_28728,N_28945);
xnor U29338 (N_29338,N_28966,N_28741);
nand U29339 (N_29339,N_28522,N_28895);
nand U29340 (N_29340,N_28701,N_28803);
or U29341 (N_29341,N_28697,N_28809);
nor U29342 (N_29342,N_28913,N_28834);
or U29343 (N_29343,N_28681,N_28606);
and U29344 (N_29344,N_28815,N_28546);
and U29345 (N_29345,N_28726,N_28920);
and U29346 (N_29346,N_28664,N_28715);
nor U29347 (N_29347,N_28957,N_28801);
xnor U29348 (N_29348,N_28986,N_28868);
xor U29349 (N_29349,N_28573,N_28596);
nand U29350 (N_29350,N_28526,N_28723);
nand U29351 (N_29351,N_28656,N_28553);
nor U29352 (N_29352,N_28785,N_28690);
nand U29353 (N_29353,N_28675,N_28818);
and U29354 (N_29354,N_28913,N_28916);
nor U29355 (N_29355,N_28875,N_28584);
nor U29356 (N_29356,N_28658,N_28866);
or U29357 (N_29357,N_28797,N_28822);
nand U29358 (N_29358,N_28937,N_28948);
xnor U29359 (N_29359,N_28721,N_28855);
xnor U29360 (N_29360,N_28733,N_28659);
nor U29361 (N_29361,N_28783,N_28651);
and U29362 (N_29362,N_28785,N_28966);
xor U29363 (N_29363,N_28828,N_28985);
nand U29364 (N_29364,N_28868,N_28788);
or U29365 (N_29365,N_28592,N_28682);
or U29366 (N_29366,N_28712,N_28594);
xnor U29367 (N_29367,N_28905,N_28790);
xnor U29368 (N_29368,N_28769,N_28914);
or U29369 (N_29369,N_28567,N_28705);
or U29370 (N_29370,N_28909,N_28733);
nor U29371 (N_29371,N_28582,N_28616);
or U29372 (N_29372,N_28810,N_28517);
and U29373 (N_29373,N_28703,N_28857);
nor U29374 (N_29374,N_28520,N_28618);
nand U29375 (N_29375,N_28682,N_28737);
nand U29376 (N_29376,N_28683,N_28995);
and U29377 (N_29377,N_28834,N_28662);
nand U29378 (N_29378,N_28774,N_28884);
nand U29379 (N_29379,N_28619,N_28894);
xnor U29380 (N_29380,N_28904,N_28578);
xor U29381 (N_29381,N_28951,N_28639);
xnor U29382 (N_29382,N_28671,N_28745);
xor U29383 (N_29383,N_28851,N_28511);
or U29384 (N_29384,N_28837,N_28781);
nand U29385 (N_29385,N_28927,N_28690);
nor U29386 (N_29386,N_28918,N_28563);
or U29387 (N_29387,N_28573,N_28708);
nor U29388 (N_29388,N_28550,N_28877);
nand U29389 (N_29389,N_28741,N_28959);
nor U29390 (N_29390,N_28921,N_28941);
nor U29391 (N_29391,N_28720,N_28869);
nor U29392 (N_29392,N_28509,N_28972);
nor U29393 (N_29393,N_28550,N_28616);
xnor U29394 (N_29394,N_28911,N_28549);
or U29395 (N_29395,N_28857,N_28802);
xor U29396 (N_29396,N_28899,N_28881);
nor U29397 (N_29397,N_28751,N_28863);
and U29398 (N_29398,N_28983,N_28923);
nand U29399 (N_29399,N_28788,N_28639);
and U29400 (N_29400,N_28811,N_28708);
and U29401 (N_29401,N_28767,N_28556);
xor U29402 (N_29402,N_28617,N_28526);
nand U29403 (N_29403,N_28673,N_28835);
or U29404 (N_29404,N_28753,N_28552);
xnor U29405 (N_29405,N_28525,N_28690);
or U29406 (N_29406,N_28596,N_28932);
xnor U29407 (N_29407,N_28659,N_28763);
xor U29408 (N_29408,N_28994,N_28509);
and U29409 (N_29409,N_28700,N_28918);
nor U29410 (N_29410,N_28810,N_28939);
xnor U29411 (N_29411,N_28570,N_28767);
nand U29412 (N_29412,N_28547,N_28736);
or U29413 (N_29413,N_28932,N_28963);
and U29414 (N_29414,N_28501,N_28554);
nand U29415 (N_29415,N_28850,N_28522);
and U29416 (N_29416,N_28989,N_28700);
nor U29417 (N_29417,N_28758,N_28756);
nor U29418 (N_29418,N_28723,N_28629);
and U29419 (N_29419,N_28953,N_28512);
or U29420 (N_29420,N_28650,N_28895);
or U29421 (N_29421,N_28859,N_28986);
or U29422 (N_29422,N_28537,N_28538);
nor U29423 (N_29423,N_28504,N_28824);
xor U29424 (N_29424,N_28882,N_28532);
nand U29425 (N_29425,N_28530,N_28862);
nor U29426 (N_29426,N_28511,N_28845);
nand U29427 (N_29427,N_28609,N_28635);
or U29428 (N_29428,N_28962,N_28694);
or U29429 (N_29429,N_28682,N_28841);
nor U29430 (N_29430,N_28686,N_28550);
nor U29431 (N_29431,N_28829,N_28628);
or U29432 (N_29432,N_28592,N_28523);
or U29433 (N_29433,N_28695,N_28992);
nor U29434 (N_29434,N_28787,N_28537);
nor U29435 (N_29435,N_28680,N_28600);
or U29436 (N_29436,N_28941,N_28609);
and U29437 (N_29437,N_28938,N_28787);
and U29438 (N_29438,N_28887,N_28701);
nor U29439 (N_29439,N_28784,N_28731);
nor U29440 (N_29440,N_28731,N_28879);
nor U29441 (N_29441,N_28893,N_28747);
nand U29442 (N_29442,N_28604,N_28626);
nand U29443 (N_29443,N_28796,N_28797);
xor U29444 (N_29444,N_28868,N_28595);
or U29445 (N_29445,N_28505,N_28594);
or U29446 (N_29446,N_28836,N_28714);
nand U29447 (N_29447,N_28627,N_28966);
nand U29448 (N_29448,N_28845,N_28834);
nor U29449 (N_29449,N_28818,N_28567);
nor U29450 (N_29450,N_28932,N_28957);
nor U29451 (N_29451,N_28509,N_28908);
and U29452 (N_29452,N_28562,N_28682);
nand U29453 (N_29453,N_28563,N_28868);
or U29454 (N_29454,N_28919,N_28521);
nor U29455 (N_29455,N_28537,N_28950);
or U29456 (N_29456,N_28765,N_28991);
xnor U29457 (N_29457,N_28698,N_28896);
nor U29458 (N_29458,N_28760,N_28706);
or U29459 (N_29459,N_28879,N_28940);
nor U29460 (N_29460,N_28956,N_28507);
nor U29461 (N_29461,N_28912,N_28812);
nand U29462 (N_29462,N_28540,N_28924);
and U29463 (N_29463,N_28895,N_28621);
or U29464 (N_29464,N_28699,N_28634);
or U29465 (N_29465,N_28761,N_28977);
or U29466 (N_29466,N_28922,N_28620);
nor U29467 (N_29467,N_28953,N_28618);
and U29468 (N_29468,N_28608,N_28707);
nor U29469 (N_29469,N_28745,N_28949);
xor U29470 (N_29470,N_28901,N_28919);
and U29471 (N_29471,N_28901,N_28588);
or U29472 (N_29472,N_28877,N_28914);
or U29473 (N_29473,N_28948,N_28804);
or U29474 (N_29474,N_28826,N_28754);
xnor U29475 (N_29475,N_28503,N_28886);
nor U29476 (N_29476,N_28848,N_28945);
and U29477 (N_29477,N_28520,N_28733);
nand U29478 (N_29478,N_28579,N_28732);
nor U29479 (N_29479,N_28672,N_28892);
and U29480 (N_29480,N_28613,N_28620);
nand U29481 (N_29481,N_28646,N_28602);
nor U29482 (N_29482,N_28821,N_28576);
xor U29483 (N_29483,N_28649,N_28795);
nand U29484 (N_29484,N_28943,N_28862);
and U29485 (N_29485,N_28736,N_28730);
and U29486 (N_29486,N_28907,N_28960);
nand U29487 (N_29487,N_28521,N_28798);
xnor U29488 (N_29488,N_28738,N_28941);
and U29489 (N_29489,N_28763,N_28966);
nand U29490 (N_29490,N_28879,N_28772);
xor U29491 (N_29491,N_28855,N_28851);
and U29492 (N_29492,N_28993,N_28527);
nor U29493 (N_29493,N_28532,N_28924);
nor U29494 (N_29494,N_28822,N_28801);
nor U29495 (N_29495,N_28917,N_28756);
nand U29496 (N_29496,N_28957,N_28638);
nor U29497 (N_29497,N_28590,N_28786);
xor U29498 (N_29498,N_28926,N_28999);
nor U29499 (N_29499,N_28984,N_28938);
and U29500 (N_29500,N_29285,N_29437);
xnor U29501 (N_29501,N_29434,N_29164);
or U29502 (N_29502,N_29299,N_29483);
nor U29503 (N_29503,N_29482,N_29209);
nand U29504 (N_29504,N_29108,N_29348);
nand U29505 (N_29505,N_29467,N_29356);
nand U29506 (N_29506,N_29246,N_29460);
nand U29507 (N_29507,N_29363,N_29110);
or U29508 (N_29508,N_29111,N_29327);
or U29509 (N_29509,N_29249,N_29449);
nor U29510 (N_29510,N_29125,N_29134);
or U29511 (N_29511,N_29095,N_29331);
nor U29512 (N_29512,N_29390,N_29173);
xnor U29513 (N_29513,N_29073,N_29179);
nor U29514 (N_29514,N_29219,N_29212);
nor U29515 (N_29515,N_29038,N_29378);
and U29516 (N_29516,N_29060,N_29191);
and U29517 (N_29517,N_29431,N_29440);
and U29518 (N_29518,N_29372,N_29160);
xnor U29519 (N_29519,N_29308,N_29394);
nand U29520 (N_29520,N_29397,N_29387);
and U29521 (N_29521,N_29093,N_29468);
nand U29522 (N_29522,N_29368,N_29415);
nor U29523 (N_29523,N_29033,N_29315);
nor U29524 (N_29524,N_29251,N_29369);
nand U29525 (N_29525,N_29053,N_29425);
or U29526 (N_29526,N_29446,N_29254);
and U29527 (N_29527,N_29341,N_29463);
or U29528 (N_29528,N_29492,N_29304);
and U29529 (N_29529,N_29079,N_29210);
nand U29530 (N_29530,N_29207,N_29407);
or U29531 (N_29531,N_29114,N_29020);
nand U29532 (N_29532,N_29245,N_29223);
xor U29533 (N_29533,N_29412,N_29213);
and U29534 (N_29534,N_29069,N_29347);
and U29535 (N_29535,N_29025,N_29255);
or U29536 (N_29536,N_29035,N_29433);
nor U29537 (N_29537,N_29211,N_29100);
and U29538 (N_29538,N_29208,N_29154);
and U29539 (N_29539,N_29455,N_29193);
nand U29540 (N_29540,N_29320,N_29247);
nor U29541 (N_29541,N_29082,N_29395);
and U29542 (N_29542,N_29274,N_29126);
nor U29543 (N_29543,N_29480,N_29295);
nor U29544 (N_29544,N_29058,N_29105);
and U29545 (N_29545,N_29004,N_29464);
nor U29546 (N_29546,N_29155,N_29161);
nand U29547 (N_29547,N_29279,N_29199);
xor U29548 (N_29548,N_29250,N_29107);
and U29549 (N_29549,N_29350,N_29151);
and U29550 (N_29550,N_29358,N_29271);
and U29551 (N_29551,N_29143,N_29156);
or U29552 (N_29552,N_29317,N_29198);
nor U29553 (N_29553,N_29090,N_29413);
xor U29554 (N_29554,N_29019,N_29451);
nand U29555 (N_29555,N_29404,N_29051);
nand U29556 (N_29556,N_29041,N_29136);
or U29557 (N_29557,N_29384,N_29221);
and U29558 (N_29558,N_29248,N_29220);
or U29559 (N_29559,N_29287,N_29186);
and U29560 (N_29560,N_29233,N_29008);
xnor U29561 (N_29561,N_29044,N_29086);
and U29562 (N_29562,N_29491,N_29293);
nand U29563 (N_29563,N_29228,N_29040);
nor U29564 (N_29564,N_29229,N_29049);
nand U29565 (N_29565,N_29286,N_29266);
xor U29566 (N_29566,N_29153,N_29351);
and U29567 (N_29567,N_29343,N_29493);
nand U29568 (N_29568,N_29487,N_29311);
nor U29569 (N_29569,N_29381,N_29336);
xnor U29570 (N_29570,N_29195,N_29243);
nand U29571 (N_29571,N_29074,N_29417);
nor U29572 (N_29572,N_29264,N_29022);
or U29573 (N_29573,N_29138,N_29026);
nand U29574 (N_29574,N_29353,N_29080);
xor U29575 (N_29575,N_29300,N_29280);
nor U29576 (N_29576,N_29194,N_29103);
nand U29577 (N_29577,N_29340,N_29326);
nand U29578 (N_29578,N_29135,N_29236);
nor U29579 (N_29579,N_29273,N_29158);
xor U29580 (N_29580,N_29365,N_29032);
xor U29581 (N_29581,N_29106,N_29147);
nor U29582 (N_29582,N_29361,N_29094);
or U29583 (N_29583,N_29054,N_29102);
nor U29584 (N_29584,N_29190,N_29376);
and U29585 (N_29585,N_29104,N_29183);
or U29586 (N_29586,N_29063,N_29206);
and U29587 (N_29587,N_29003,N_29486);
or U29588 (N_29588,N_29024,N_29441);
nand U29589 (N_29589,N_29214,N_29152);
nor U29590 (N_29590,N_29314,N_29442);
xor U29591 (N_29591,N_29338,N_29310);
nor U29592 (N_29592,N_29202,N_29131);
or U29593 (N_29593,N_29130,N_29218);
nand U29594 (N_29594,N_29101,N_29128);
xor U29595 (N_29595,N_29410,N_29276);
and U29596 (N_29596,N_29148,N_29419);
or U29597 (N_29597,N_29252,N_29355);
xor U29598 (N_29598,N_29087,N_29309);
nand U29599 (N_29599,N_29428,N_29169);
xor U29600 (N_29600,N_29119,N_29474);
xor U29601 (N_29601,N_29352,N_29313);
nor U29602 (N_29602,N_29461,N_29129);
and U29603 (N_29603,N_29029,N_29362);
or U29604 (N_29604,N_29132,N_29002);
xnor U29605 (N_29605,N_29364,N_29489);
and U29606 (N_29606,N_29445,N_29027);
nor U29607 (N_29607,N_29188,N_29334);
xnor U29608 (N_29608,N_29477,N_29142);
nand U29609 (N_29609,N_29481,N_29242);
nor U29610 (N_29610,N_29204,N_29373);
and U29611 (N_29611,N_29203,N_29399);
and U29612 (N_29612,N_29490,N_29485);
xor U29613 (N_29613,N_29081,N_29170);
nand U29614 (N_29614,N_29123,N_29330);
and U29615 (N_29615,N_29046,N_29416);
nor U29616 (N_29616,N_29017,N_29388);
and U29617 (N_29617,N_29345,N_29168);
xor U29618 (N_29618,N_29196,N_29393);
nor U29619 (N_29619,N_29201,N_29175);
xnor U29620 (N_29620,N_29016,N_29357);
xnor U29621 (N_29621,N_29262,N_29056);
nand U29622 (N_29622,N_29466,N_29307);
nand U29623 (N_29623,N_29405,N_29075);
and U29624 (N_29624,N_29122,N_29406);
xnor U29625 (N_29625,N_29297,N_29303);
or U29626 (N_29626,N_29064,N_29031);
nand U29627 (N_29627,N_29462,N_29222);
or U29628 (N_29628,N_29414,N_29332);
nor U29629 (N_29629,N_29085,N_29318);
xnor U29630 (N_29630,N_29112,N_29084);
xnor U29631 (N_29631,N_29366,N_29237);
nor U29632 (N_29632,N_29429,N_29167);
and U29633 (N_29633,N_29015,N_29217);
or U29634 (N_29634,N_29234,N_29007);
or U29635 (N_29635,N_29302,N_29200);
and U29636 (N_29636,N_29411,N_29312);
and U29637 (N_29637,N_29178,N_29408);
nand U29638 (N_29638,N_29231,N_29478);
and U29639 (N_29639,N_29071,N_29121);
xor U29640 (N_29640,N_29324,N_29224);
xnor U29641 (N_29641,N_29197,N_29244);
and U29642 (N_29642,N_29037,N_29127);
and U29643 (N_29643,N_29227,N_29113);
or U29644 (N_29644,N_29000,N_29342);
or U29645 (N_29645,N_29281,N_29470);
and U29646 (N_29646,N_29042,N_29070);
nor U29647 (N_29647,N_29141,N_29494);
or U29648 (N_29648,N_29099,N_29055);
or U29649 (N_29649,N_29269,N_29185);
and U29650 (N_29650,N_29339,N_29239);
xor U29651 (N_29651,N_29323,N_29174);
or U29652 (N_29652,N_29473,N_29162);
xnor U29653 (N_29653,N_29306,N_29382);
nor U29654 (N_29654,N_29235,N_29475);
xor U29655 (N_29655,N_29159,N_29459);
nand U29656 (N_29656,N_29010,N_29270);
or U29657 (N_29657,N_29023,N_29497);
nand U29658 (N_29658,N_29157,N_29139);
and U29659 (N_29659,N_29498,N_29275);
xnor U29660 (N_29660,N_29346,N_29439);
nor U29661 (N_29661,N_29253,N_29050);
nand U29662 (N_29662,N_29379,N_29328);
xnor U29663 (N_29663,N_29012,N_29321);
or U29664 (N_29664,N_29165,N_29453);
xnor U29665 (N_29665,N_29215,N_29034);
and U29666 (N_29666,N_29078,N_29265);
nor U29667 (N_29667,N_29177,N_29385);
or U29668 (N_29668,N_29232,N_29120);
and U29669 (N_29669,N_29189,N_29496);
and U29670 (N_29670,N_29182,N_29499);
nor U29671 (N_29671,N_29447,N_29258);
or U29672 (N_29672,N_29421,N_29359);
or U29673 (N_29673,N_29116,N_29171);
nor U29674 (N_29674,N_29396,N_29418);
xnor U29675 (N_29675,N_29284,N_29205);
nand U29676 (N_29676,N_29009,N_29192);
or U29677 (N_29677,N_29146,N_29316);
nor U29678 (N_29678,N_29374,N_29344);
xnor U29679 (N_29679,N_29001,N_29370);
nor U29680 (N_29680,N_29030,N_29013);
and U29681 (N_29681,N_29149,N_29277);
and U29682 (N_29682,N_29319,N_29184);
xor U29683 (N_29683,N_29427,N_29067);
and U29684 (N_29684,N_29292,N_29140);
xor U29685 (N_29685,N_29268,N_29263);
and U29686 (N_29686,N_29450,N_29089);
nand U29687 (N_29687,N_29456,N_29432);
nor U29688 (N_29688,N_29403,N_29371);
nand U29689 (N_29689,N_29062,N_29039);
xor U29690 (N_29690,N_29296,N_29290);
and U29691 (N_29691,N_29057,N_29052);
xor U29692 (N_29692,N_29426,N_29172);
nand U29693 (N_29693,N_29181,N_29045);
xnor U29694 (N_29694,N_29230,N_29150);
and U29695 (N_29695,N_29005,N_29438);
nor U29696 (N_29696,N_29484,N_29325);
xnor U29697 (N_29697,N_29018,N_29435);
nand U29698 (N_29698,N_29430,N_29377);
xnor U29699 (N_29699,N_29322,N_29457);
or U29700 (N_29700,N_29329,N_29241);
or U29701 (N_29701,N_29144,N_29118);
and U29702 (N_29702,N_29226,N_29444);
nor U29703 (N_29703,N_29176,N_29420);
nand U29704 (N_29704,N_29238,N_29036);
xnor U29705 (N_29705,N_29092,N_29028);
and U29706 (N_29706,N_29422,N_29448);
nor U29707 (N_29707,N_29476,N_29360);
nand U29708 (N_29708,N_29458,N_29137);
nand U29709 (N_29709,N_29068,N_29391);
and U29710 (N_29710,N_29257,N_29267);
nor U29711 (N_29711,N_29261,N_29088);
and U29712 (N_29712,N_29349,N_29278);
xor U29713 (N_29713,N_29333,N_29240);
xor U29714 (N_29714,N_29454,N_29452);
nor U29715 (N_29715,N_29259,N_29021);
and U29716 (N_29716,N_29091,N_29187);
xnor U29717 (N_29717,N_29256,N_29166);
nor U29718 (N_29718,N_29260,N_29043);
or U29719 (N_29719,N_29096,N_29282);
or U29720 (N_29720,N_29283,N_29375);
and U29721 (N_29721,N_29098,N_29443);
and U29722 (N_29722,N_29145,N_29180);
nand U29723 (N_29723,N_29048,N_29294);
and U29724 (N_29724,N_29392,N_29124);
nor U29725 (N_29725,N_29401,N_29479);
or U29726 (N_29726,N_29465,N_29409);
nor U29727 (N_29727,N_29301,N_29109);
nand U29728 (N_29728,N_29495,N_29383);
and U29729 (N_29729,N_29469,N_29288);
nand U29730 (N_29730,N_29006,N_29337);
and U29731 (N_29731,N_29077,N_29066);
and U29732 (N_29732,N_29076,N_29059);
xnor U29733 (N_29733,N_29097,N_29163);
and U29734 (N_29734,N_29389,N_29225);
or U29735 (N_29735,N_29065,N_29272);
or U29736 (N_29736,N_29488,N_29289);
and U29737 (N_29737,N_29471,N_29115);
and U29738 (N_29738,N_29291,N_29335);
or U29739 (N_29739,N_29061,N_29400);
or U29740 (N_29740,N_29424,N_29423);
nor U29741 (N_29741,N_29216,N_29047);
nand U29742 (N_29742,N_29386,N_29011);
and U29743 (N_29743,N_29083,N_29398);
nand U29744 (N_29744,N_29380,N_29354);
and U29745 (N_29745,N_29436,N_29298);
nand U29746 (N_29746,N_29133,N_29014);
nand U29747 (N_29747,N_29072,N_29367);
xor U29748 (N_29748,N_29402,N_29305);
or U29749 (N_29749,N_29472,N_29117);
nor U29750 (N_29750,N_29087,N_29033);
or U29751 (N_29751,N_29072,N_29052);
xnor U29752 (N_29752,N_29384,N_29370);
nor U29753 (N_29753,N_29316,N_29180);
nor U29754 (N_29754,N_29048,N_29101);
nor U29755 (N_29755,N_29378,N_29147);
nor U29756 (N_29756,N_29203,N_29009);
or U29757 (N_29757,N_29287,N_29444);
and U29758 (N_29758,N_29280,N_29198);
nor U29759 (N_29759,N_29019,N_29349);
and U29760 (N_29760,N_29309,N_29261);
nor U29761 (N_29761,N_29197,N_29192);
or U29762 (N_29762,N_29360,N_29415);
nand U29763 (N_29763,N_29270,N_29370);
or U29764 (N_29764,N_29228,N_29215);
and U29765 (N_29765,N_29192,N_29279);
and U29766 (N_29766,N_29396,N_29242);
xor U29767 (N_29767,N_29431,N_29057);
and U29768 (N_29768,N_29241,N_29279);
nor U29769 (N_29769,N_29477,N_29011);
and U29770 (N_29770,N_29339,N_29135);
and U29771 (N_29771,N_29289,N_29049);
and U29772 (N_29772,N_29248,N_29409);
nand U29773 (N_29773,N_29263,N_29242);
or U29774 (N_29774,N_29485,N_29190);
nor U29775 (N_29775,N_29189,N_29161);
xor U29776 (N_29776,N_29276,N_29192);
nor U29777 (N_29777,N_29198,N_29158);
nor U29778 (N_29778,N_29313,N_29391);
nor U29779 (N_29779,N_29073,N_29332);
nor U29780 (N_29780,N_29042,N_29324);
nand U29781 (N_29781,N_29208,N_29221);
or U29782 (N_29782,N_29118,N_29274);
or U29783 (N_29783,N_29341,N_29201);
nand U29784 (N_29784,N_29440,N_29155);
or U29785 (N_29785,N_29007,N_29291);
nor U29786 (N_29786,N_29263,N_29001);
nand U29787 (N_29787,N_29041,N_29371);
nand U29788 (N_29788,N_29338,N_29015);
or U29789 (N_29789,N_29129,N_29184);
and U29790 (N_29790,N_29115,N_29252);
nor U29791 (N_29791,N_29241,N_29085);
nand U29792 (N_29792,N_29083,N_29471);
nor U29793 (N_29793,N_29139,N_29467);
xor U29794 (N_29794,N_29186,N_29083);
nand U29795 (N_29795,N_29089,N_29138);
nand U29796 (N_29796,N_29214,N_29158);
and U29797 (N_29797,N_29499,N_29366);
nor U29798 (N_29798,N_29010,N_29370);
or U29799 (N_29799,N_29229,N_29213);
and U29800 (N_29800,N_29344,N_29159);
or U29801 (N_29801,N_29189,N_29219);
and U29802 (N_29802,N_29218,N_29069);
and U29803 (N_29803,N_29004,N_29008);
and U29804 (N_29804,N_29054,N_29316);
nand U29805 (N_29805,N_29160,N_29108);
nor U29806 (N_29806,N_29312,N_29218);
and U29807 (N_29807,N_29448,N_29176);
nor U29808 (N_29808,N_29087,N_29248);
nor U29809 (N_29809,N_29366,N_29421);
and U29810 (N_29810,N_29137,N_29340);
xnor U29811 (N_29811,N_29276,N_29316);
nor U29812 (N_29812,N_29279,N_29293);
nand U29813 (N_29813,N_29139,N_29227);
and U29814 (N_29814,N_29084,N_29086);
xor U29815 (N_29815,N_29181,N_29258);
xnor U29816 (N_29816,N_29303,N_29183);
nand U29817 (N_29817,N_29063,N_29305);
nand U29818 (N_29818,N_29276,N_29262);
and U29819 (N_29819,N_29384,N_29063);
and U29820 (N_29820,N_29213,N_29163);
xor U29821 (N_29821,N_29454,N_29295);
and U29822 (N_29822,N_29161,N_29332);
xor U29823 (N_29823,N_29325,N_29427);
nor U29824 (N_29824,N_29224,N_29185);
xor U29825 (N_29825,N_29215,N_29013);
or U29826 (N_29826,N_29143,N_29138);
and U29827 (N_29827,N_29008,N_29475);
and U29828 (N_29828,N_29132,N_29325);
xnor U29829 (N_29829,N_29232,N_29437);
and U29830 (N_29830,N_29092,N_29160);
or U29831 (N_29831,N_29205,N_29256);
nor U29832 (N_29832,N_29050,N_29110);
xor U29833 (N_29833,N_29134,N_29059);
and U29834 (N_29834,N_29399,N_29117);
and U29835 (N_29835,N_29364,N_29385);
or U29836 (N_29836,N_29293,N_29174);
nor U29837 (N_29837,N_29091,N_29066);
xnor U29838 (N_29838,N_29062,N_29167);
nor U29839 (N_29839,N_29334,N_29082);
nor U29840 (N_29840,N_29482,N_29284);
and U29841 (N_29841,N_29429,N_29369);
nand U29842 (N_29842,N_29170,N_29105);
nor U29843 (N_29843,N_29200,N_29371);
xor U29844 (N_29844,N_29062,N_29281);
and U29845 (N_29845,N_29128,N_29361);
or U29846 (N_29846,N_29209,N_29178);
or U29847 (N_29847,N_29371,N_29114);
or U29848 (N_29848,N_29045,N_29378);
nor U29849 (N_29849,N_29494,N_29326);
nor U29850 (N_29850,N_29233,N_29393);
xor U29851 (N_29851,N_29398,N_29116);
and U29852 (N_29852,N_29093,N_29241);
nor U29853 (N_29853,N_29287,N_29389);
nor U29854 (N_29854,N_29230,N_29182);
xor U29855 (N_29855,N_29199,N_29100);
and U29856 (N_29856,N_29366,N_29063);
xor U29857 (N_29857,N_29475,N_29242);
nand U29858 (N_29858,N_29329,N_29025);
nor U29859 (N_29859,N_29303,N_29328);
nor U29860 (N_29860,N_29420,N_29296);
nand U29861 (N_29861,N_29251,N_29183);
nand U29862 (N_29862,N_29385,N_29192);
nor U29863 (N_29863,N_29403,N_29078);
and U29864 (N_29864,N_29153,N_29268);
xnor U29865 (N_29865,N_29316,N_29476);
nor U29866 (N_29866,N_29251,N_29163);
or U29867 (N_29867,N_29202,N_29438);
xor U29868 (N_29868,N_29002,N_29160);
and U29869 (N_29869,N_29139,N_29347);
nand U29870 (N_29870,N_29100,N_29158);
or U29871 (N_29871,N_29116,N_29388);
xnor U29872 (N_29872,N_29435,N_29150);
xor U29873 (N_29873,N_29246,N_29243);
nand U29874 (N_29874,N_29243,N_29134);
xnor U29875 (N_29875,N_29175,N_29390);
nand U29876 (N_29876,N_29498,N_29005);
nand U29877 (N_29877,N_29063,N_29155);
nand U29878 (N_29878,N_29149,N_29046);
or U29879 (N_29879,N_29133,N_29057);
nand U29880 (N_29880,N_29126,N_29124);
xor U29881 (N_29881,N_29469,N_29480);
or U29882 (N_29882,N_29274,N_29025);
xnor U29883 (N_29883,N_29333,N_29361);
xor U29884 (N_29884,N_29032,N_29111);
and U29885 (N_29885,N_29158,N_29043);
and U29886 (N_29886,N_29215,N_29077);
xnor U29887 (N_29887,N_29422,N_29192);
nor U29888 (N_29888,N_29273,N_29348);
or U29889 (N_29889,N_29481,N_29471);
nor U29890 (N_29890,N_29304,N_29210);
xor U29891 (N_29891,N_29130,N_29056);
xnor U29892 (N_29892,N_29272,N_29383);
or U29893 (N_29893,N_29241,N_29325);
nand U29894 (N_29894,N_29270,N_29063);
nand U29895 (N_29895,N_29023,N_29099);
and U29896 (N_29896,N_29249,N_29014);
xor U29897 (N_29897,N_29127,N_29491);
xor U29898 (N_29898,N_29351,N_29430);
nor U29899 (N_29899,N_29045,N_29211);
and U29900 (N_29900,N_29352,N_29453);
nand U29901 (N_29901,N_29416,N_29326);
and U29902 (N_29902,N_29258,N_29013);
xnor U29903 (N_29903,N_29373,N_29127);
nand U29904 (N_29904,N_29138,N_29084);
or U29905 (N_29905,N_29112,N_29401);
or U29906 (N_29906,N_29004,N_29123);
nand U29907 (N_29907,N_29461,N_29031);
nor U29908 (N_29908,N_29390,N_29230);
nor U29909 (N_29909,N_29321,N_29326);
nand U29910 (N_29910,N_29346,N_29272);
or U29911 (N_29911,N_29432,N_29101);
or U29912 (N_29912,N_29322,N_29139);
xor U29913 (N_29913,N_29331,N_29456);
nand U29914 (N_29914,N_29352,N_29153);
xnor U29915 (N_29915,N_29291,N_29071);
or U29916 (N_29916,N_29255,N_29432);
nand U29917 (N_29917,N_29301,N_29151);
xnor U29918 (N_29918,N_29385,N_29481);
xnor U29919 (N_29919,N_29264,N_29387);
nand U29920 (N_29920,N_29070,N_29150);
or U29921 (N_29921,N_29467,N_29050);
nor U29922 (N_29922,N_29018,N_29413);
and U29923 (N_29923,N_29009,N_29161);
nand U29924 (N_29924,N_29326,N_29368);
and U29925 (N_29925,N_29272,N_29030);
or U29926 (N_29926,N_29470,N_29405);
and U29927 (N_29927,N_29107,N_29281);
nor U29928 (N_29928,N_29365,N_29433);
nand U29929 (N_29929,N_29128,N_29182);
nand U29930 (N_29930,N_29080,N_29049);
and U29931 (N_29931,N_29429,N_29005);
xor U29932 (N_29932,N_29251,N_29080);
nor U29933 (N_29933,N_29490,N_29065);
nand U29934 (N_29934,N_29065,N_29276);
xnor U29935 (N_29935,N_29072,N_29364);
or U29936 (N_29936,N_29001,N_29193);
nor U29937 (N_29937,N_29324,N_29283);
nand U29938 (N_29938,N_29022,N_29184);
nand U29939 (N_29939,N_29174,N_29328);
nor U29940 (N_29940,N_29311,N_29324);
nand U29941 (N_29941,N_29057,N_29264);
nand U29942 (N_29942,N_29080,N_29174);
nor U29943 (N_29943,N_29090,N_29015);
or U29944 (N_29944,N_29426,N_29490);
and U29945 (N_29945,N_29438,N_29073);
nand U29946 (N_29946,N_29203,N_29474);
xnor U29947 (N_29947,N_29265,N_29083);
nor U29948 (N_29948,N_29164,N_29309);
or U29949 (N_29949,N_29175,N_29461);
and U29950 (N_29950,N_29296,N_29114);
nor U29951 (N_29951,N_29226,N_29082);
nor U29952 (N_29952,N_29006,N_29041);
or U29953 (N_29953,N_29200,N_29297);
nor U29954 (N_29954,N_29288,N_29127);
nor U29955 (N_29955,N_29352,N_29320);
nor U29956 (N_29956,N_29302,N_29045);
and U29957 (N_29957,N_29005,N_29033);
nor U29958 (N_29958,N_29335,N_29282);
and U29959 (N_29959,N_29456,N_29299);
nor U29960 (N_29960,N_29276,N_29407);
nand U29961 (N_29961,N_29146,N_29286);
and U29962 (N_29962,N_29253,N_29096);
or U29963 (N_29963,N_29117,N_29180);
xnor U29964 (N_29964,N_29053,N_29048);
xnor U29965 (N_29965,N_29113,N_29241);
xnor U29966 (N_29966,N_29326,N_29017);
nor U29967 (N_29967,N_29310,N_29366);
xnor U29968 (N_29968,N_29206,N_29229);
or U29969 (N_29969,N_29414,N_29145);
or U29970 (N_29970,N_29056,N_29319);
nor U29971 (N_29971,N_29267,N_29101);
and U29972 (N_29972,N_29122,N_29209);
nand U29973 (N_29973,N_29133,N_29367);
and U29974 (N_29974,N_29246,N_29125);
nor U29975 (N_29975,N_29175,N_29071);
or U29976 (N_29976,N_29080,N_29374);
xnor U29977 (N_29977,N_29337,N_29165);
nor U29978 (N_29978,N_29413,N_29300);
and U29979 (N_29979,N_29215,N_29084);
nand U29980 (N_29980,N_29081,N_29381);
xnor U29981 (N_29981,N_29381,N_29020);
nand U29982 (N_29982,N_29025,N_29276);
and U29983 (N_29983,N_29164,N_29067);
or U29984 (N_29984,N_29390,N_29459);
nor U29985 (N_29985,N_29152,N_29169);
nand U29986 (N_29986,N_29472,N_29177);
nor U29987 (N_29987,N_29191,N_29139);
or U29988 (N_29988,N_29366,N_29409);
nor U29989 (N_29989,N_29228,N_29324);
xor U29990 (N_29990,N_29164,N_29374);
nand U29991 (N_29991,N_29481,N_29114);
or U29992 (N_29992,N_29032,N_29014);
nand U29993 (N_29993,N_29431,N_29203);
or U29994 (N_29994,N_29125,N_29462);
nand U29995 (N_29995,N_29225,N_29477);
or U29996 (N_29996,N_29005,N_29395);
nor U29997 (N_29997,N_29266,N_29261);
and U29998 (N_29998,N_29333,N_29401);
nor U29999 (N_29999,N_29095,N_29301);
or UO_0 (O_0,N_29979,N_29944);
nand UO_1 (O_1,N_29671,N_29683);
and UO_2 (O_2,N_29687,N_29584);
or UO_3 (O_3,N_29543,N_29812);
xor UO_4 (O_4,N_29920,N_29679);
xor UO_5 (O_5,N_29990,N_29555);
nor UO_6 (O_6,N_29975,N_29957);
nor UO_7 (O_7,N_29550,N_29757);
xnor UO_8 (O_8,N_29966,N_29904);
xor UO_9 (O_9,N_29621,N_29839);
nor UO_10 (O_10,N_29770,N_29760);
nand UO_11 (O_11,N_29885,N_29766);
nand UO_12 (O_12,N_29559,N_29850);
nor UO_13 (O_13,N_29716,N_29572);
nand UO_14 (O_14,N_29865,N_29593);
xor UO_15 (O_15,N_29703,N_29985);
xnor UO_16 (O_16,N_29519,N_29803);
and UO_17 (O_17,N_29870,N_29750);
nor UO_18 (O_18,N_29704,N_29747);
and UO_19 (O_19,N_29776,N_29767);
nand UO_20 (O_20,N_29748,N_29590);
nor UO_21 (O_21,N_29657,N_29783);
nand UO_22 (O_22,N_29548,N_29591);
xnor UO_23 (O_23,N_29745,N_29749);
and UO_24 (O_24,N_29722,N_29892);
nor UO_25 (O_25,N_29836,N_29582);
xor UO_26 (O_26,N_29815,N_29529);
and UO_27 (O_27,N_29987,N_29670);
nor UO_28 (O_28,N_29717,N_29609);
xnor UO_29 (O_29,N_29965,N_29570);
nor UO_30 (O_30,N_29580,N_29890);
nor UO_31 (O_31,N_29638,N_29739);
nor UO_32 (O_32,N_29505,N_29759);
or UO_33 (O_33,N_29897,N_29787);
nor UO_34 (O_34,N_29614,N_29594);
xor UO_35 (O_35,N_29651,N_29962);
nor UO_36 (O_36,N_29773,N_29964);
xnor UO_37 (O_37,N_29829,N_29700);
nand UO_38 (O_38,N_29845,N_29680);
xor UO_39 (O_39,N_29894,N_29589);
or UO_40 (O_40,N_29627,N_29863);
nand UO_41 (O_41,N_29996,N_29765);
nor UO_42 (O_42,N_29831,N_29856);
nor UO_43 (O_43,N_29713,N_29502);
xor UO_44 (O_44,N_29632,N_29793);
nor UO_45 (O_45,N_29763,N_29697);
nand UO_46 (O_46,N_29661,N_29938);
nand UO_47 (O_47,N_29706,N_29501);
and UO_48 (O_48,N_29654,N_29669);
and UO_49 (O_49,N_29673,N_29796);
and UO_50 (O_50,N_29681,N_29525);
xnor UO_51 (O_51,N_29729,N_29521);
nand UO_52 (O_52,N_29734,N_29574);
or UO_53 (O_53,N_29715,N_29668);
and UO_54 (O_54,N_29616,N_29597);
nor UO_55 (O_55,N_29939,N_29712);
or UO_56 (O_56,N_29823,N_29950);
nor UO_57 (O_57,N_29520,N_29980);
and UO_58 (O_58,N_29694,N_29533);
or UO_59 (O_59,N_29513,N_29549);
and UO_60 (O_60,N_29906,N_29932);
nand UO_61 (O_61,N_29873,N_29608);
xnor UO_62 (O_62,N_29988,N_29725);
nand UO_63 (O_63,N_29804,N_29833);
and UO_64 (O_64,N_29790,N_29561);
or UO_65 (O_65,N_29603,N_29604);
nand UO_66 (O_66,N_29972,N_29951);
nor UO_67 (O_67,N_29620,N_29907);
and UO_68 (O_68,N_29605,N_29779);
or UO_69 (O_69,N_29691,N_29901);
or UO_70 (O_70,N_29995,N_29982);
and UO_71 (O_71,N_29840,N_29948);
xnor UO_72 (O_72,N_29641,N_29688);
nor UO_73 (O_73,N_29586,N_29900);
nand UO_74 (O_74,N_29772,N_29899);
xor UO_75 (O_75,N_29816,N_29913);
and UO_76 (O_76,N_29719,N_29986);
nand UO_77 (O_77,N_29714,N_29931);
and UO_78 (O_78,N_29649,N_29999);
nor UO_79 (O_79,N_29647,N_29784);
or UO_80 (O_80,N_29595,N_29838);
nor UO_81 (O_81,N_29884,N_29699);
nand UO_82 (O_82,N_29507,N_29983);
nor UO_83 (O_83,N_29653,N_29792);
or UO_84 (O_84,N_29510,N_29933);
or UO_85 (O_85,N_29740,N_29943);
nand UO_86 (O_86,N_29882,N_29583);
xnor UO_87 (O_87,N_29678,N_29958);
or UO_88 (O_88,N_29567,N_29924);
xor UO_89 (O_89,N_29600,N_29636);
and UO_90 (O_90,N_29825,N_29676);
or UO_91 (O_91,N_29822,N_29895);
nand UO_92 (O_92,N_29702,N_29728);
nor UO_93 (O_93,N_29707,N_29755);
nor UO_94 (O_94,N_29585,N_29830);
nor UO_95 (O_95,N_29896,N_29746);
nor UO_96 (O_96,N_29841,N_29953);
nand UO_97 (O_97,N_29547,N_29587);
or UO_98 (O_98,N_29859,N_29518);
nand UO_99 (O_99,N_29788,N_29629);
nand UO_100 (O_100,N_29974,N_29733);
xnor UO_101 (O_101,N_29880,N_29743);
and UO_102 (O_102,N_29805,N_29877);
nor UO_103 (O_103,N_29517,N_29886);
xor UO_104 (O_104,N_29613,N_29752);
nand UO_105 (O_105,N_29540,N_29512);
or UO_106 (O_106,N_29709,N_29817);
xor UO_107 (O_107,N_29780,N_29868);
or UO_108 (O_108,N_29558,N_29541);
xnor UO_109 (O_109,N_29837,N_29891);
xnor UO_110 (O_110,N_29564,N_29835);
and UO_111 (O_111,N_29786,N_29644);
and UO_112 (O_112,N_29573,N_29522);
and UO_113 (O_113,N_29961,N_29775);
nand UO_114 (O_114,N_29738,N_29528);
and UO_115 (O_115,N_29970,N_29848);
or UO_116 (O_116,N_29633,N_29861);
nor UO_117 (O_117,N_29727,N_29710);
and UO_118 (O_118,N_29946,N_29610);
nor UO_119 (O_119,N_29864,N_29937);
nor UO_120 (O_120,N_29860,N_29854);
or UO_121 (O_121,N_29640,N_29674);
nand UO_122 (O_122,N_29696,N_29834);
nor UO_123 (O_123,N_29634,N_29802);
xor UO_124 (O_124,N_29735,N_29925);
nor UO_125 (O_125,N_29565,N_29566);
and UO_126 (O_126,N_29628,N_29506);
xor UO_127 (O_127,N_29509,N_29853);
or UO_128 (O_128,N_29508,N_29945);
and UO_129 (O_129,N_29821,N_29797);
nand UO_130 (O_130,N_29579,N_29682);
xor UO_131 (O_131,N_29592,N_29794);
nand UO_132 (O_132,N_29617,N_29826);
nor UO_133 (O_133,N_29523,N_29978);
nand UO_134 (O_134,N_29997,N_29635);
and UO_135 (O_135,N_29720,N_29844);
nor UO_136 (O_136,N_29599,N_29503);
nor UO_137 (O_137,N_29998,N_29562);
or UO_138 (O_138,N_29730,N_29893);
or UO_139 (O_139,N_29539,N_29601);
nor UO_140 (O_140,N_29809,N_29947);
nand UO_141 (O_141,N_29846,N_29832);
and UO_142 (O_142,N_29785,N_29909);
and UO_143 (O_143,N_29511,N_29551);
nor UO_144 (O_144,N_29887,N_29708);
nor UO_145 (O_145,N_29941,N_29981);
or UO_146 (O_146,N_29940,N_29534);
nand UO_147 (O_147,N_29929,N_29935);
or UO_148 (O_148,N_29615,N_29989);
nand UO_149 (O_149,N_29560,N_29910);
nor UO_150 (O_150,N_29955,N_29949);
nand UO_151 (O_151,N_29842,N_29535);
and UO_152 (O_152,N_29642,N_29606);
nor UO_153 (O_153,N_29984,N_29923);
nor UO_154 (O_154,N_29774,N_29820);
or UO_155 (O_155,N_29530,N_29875);
nand UO_156 (O_156,N_29643,N_29928);
or UO_157 (O_157,N_29611,N_29798);
and UO_158 (O_158,N_29905,N_29578);
or UO_159 (O_159,N_29690,N_29898);
nand UO_160 (O_160,N_29667,N_29847);
and UO_161 (O_161,N_29960,N_29568);
nand UO_162 (O_162,N_29542,N_29625);
xnor UO_163 (O_163,N_29992,N_29942);
and UO_164 (O_164,N_29754,N_29652);
nor UO_165 (O_165,N_29655,N_29554);
nor UO_166 (O_166,N_29753,N_29973);
xnor UO_167 (O_167,N_29867,N_29685);
nor UO_168 (O_168,N_29612,N_29824);
nand UO_169 (O_169,N_29806,N_29857);
and UO_170 (O_170,N_29665,N_29721);
xnor UO_171 (O_171,N_29645,N_29675);
and UO_172 (O_172,N_29736,N_29677);
or UO_173 (O_173,N_29919,N_29624);
and UO_174 (O_174,N_29531,N_29827);
or UO_175 (O_175,N_29741,N_29516);
and UO_176 (O_176,N_29618,N_29936);
nand UO_177 (O_177,N_29789,N_29811);
and UO_178 (O_178,N_29956,N_29952);
nor UO_179 (O_179,N_29902,N_29637);
xor UO_180 (O_180,N_29819,N_29814);
and UO_181 (O_181,N_29963,N_29874);
nor UO_182 (O_182,N_29758,N_29810);
nor UO_183 (O_183,N_29571,N_29828);
and UO_184 (O_184,N_29818,N_29879);
or UO_185 (O_185,N_29575,N_29648);
xor UO_186 (O_186,N_29576,N_29777);
or UO_187 (O_187,N_29544,N_29976);
nand UO_188 (O_188,N_29917,N_29791);
xor UO_189 (O_189,N_29514,N_29577);
and UO_190 (O_190,N_29959,N_29663);
nand UO_191 (O_191,N_29532,N_29921);
and UO_192 (O_192,N_29662,N_29598);
nor UO_193 (O_193,N_29813,N_29764);
nand UO_194 (O_194,N_29672,N_29626);
xnor UO_195 (O_195,N_29954,N_29756);
or UO_196 (O_196,N_29927,N_29914);
nor UO_197 (O_197,N_29916,N_29732);
or UO_198 (O_198,N_29744,N_29801);
xor UO_199 (O_199,N_29858,N_29724);
or UO_200 (O_200,N_29903,N_29843);
or UO_201 (O_201,N_29701,N_29698);
xor UO_202 (O_202,N_29500,N_29705);
nand UO_203 (O_203,N_29731,N_29659);
or UO_204 (O_204,N_29751,N_29768);
xor UO_205 (O_205,N_29646,N_29852);
or UO_206 (O_206,N_29851,N_29537);
nand UO_207 (O_207,N_29658,N_29623);
nand UO_208 (O_208,N_29569,N_29855);
nor UO_209 (O_209,N_29869,N_29967);
nor UO_210 (O_210,N_29808,N_29799);
and UO_211 (O_211,N_29588,N_29969);
or UO_212 (O_212,N_29684,N_29556);
or UO_213 (O_213,N_29994,N_29934);
nand UO_214 (O_214,N_29888,N_29631);
and UO_215 (O_215,N_29807,N_29908);
or UO_216 (O_216,N_29602,N_29866);
xnor UO_217 (O_217,N_29883,N_29977);
nor UO_218 (O_218,N_29800,N_29718);
nor UO_219 (O_219,N_29926,N_29607);
or UO_220 (O_220,N_29660,N_29862);
xnor UO_221 (O_221,N_29693,N_29656);
nand UO_222 (O_222,N_29871,N_29689);
xnor UO_223 (O_223,N_29666,N_29918);
and UO_224 (O_224,N_29876,N_29781);
or UO_225 (O_225,N_29915,N_29782);
and UO_226 (O_226,N_29968,N_29664);
xnor UO_227 (O_227,N_29563,N_29504);
nand UO_228 (O_228,N_29849,N_29557);
nand UO_229 (O_229,N_29546,N_29881);
or UO_230 (O_230,N_29545,N_29695);
xnor UO_231 (O_231,N_29930,N_29912);
nand UO_232 (O_232,N_29889,N_29778);
or UO_233 (O_233,N_29872,N_29737);
nand UO_234 (O_234,N_29650,N_29769);
and UO_235 (O_235,N_29991,N_29515);
nand UO_236 (O_236,N_29878,N_29761);
and UO_237 (O_237,N_29742,N_29711);
nor UO_238 (O_238,N_29993,N_29538);
and UO_239 (O_239,N_29524,N_29619);
nand UO_240 (O_240,N_29771,N_29622);
nor UO_241 (O_241,N_29971,N_29596);
and UO_242 (O_242,N_29762,N_29527);
nor UO_243 (O_243,N_29723,N_29581);
and UO_244 (O_244,N_29686,N_29692);
or UO_245 (O_245,N_29536,N_29553);
or UO_246 (O_246,N_29922,N_29911);
and UO_247 (O_247,N_29795,N_29552);
or UO_248 (O_248,N_29630,N_29526);
nor UO_249 (O_249,N_29639,N_29726);
and UO_250 (O_250,N_29859,N_29684);
nand UO_251 (O_251,N_29777,N_29951);
nor UO_252 (O_252,N_29773,N_29889);
nand UO_253 (O_253,N_29958,N_29608);
xnor UO_254 (O_254,N_29684,N_29526);
and UO_255 (O_255,N_29565,N_29923);
nor UO_256 (O_256,N_29627,N_29511);
xnor UO_257 (O_257,N_29752,N_29523);
nand UO_258 (O_258,N_29956,N_29609);
nand UO_259 (O_259,N_29996,N_29680);
nor UO_260 (O_260,N_29620,N_29705);
and UO_261 (O_261,N_29868,N_29977);
xor UO_262 (O_262,N_29775,N_29965);
or UO_263 (O_263,N_29707,N_29509);
nor UO_264 (O_264,N_29776,N_29930);
and UO_265 (O_265,N_29621,N_29737);
xor UO_266 (O_266,N_29986,N_29667);
or UO_267 (O_267,N_29788,N_29970);
nand UO_268 (O_268,N_29866,N_29531);
nor UO_269 (O_269,N_29897,N_29548);
and UO_270 (O_270,N_29790,N_29612);
nor UO_271 (O_271,N_29906,N_29910);
xor UO_272 (O_272,N_29704,N_29577);
xor UO_273 (O_273,N_29849,N_29749);
nor UO_274 (O_274,N_29895,N_29833);
xor UO_275 (O_275,N_29667,N_29815);
nor UO_276 (O_276,N_29680,N_29523);
xor UO_277 (O_277,N_29589,N_29760);
or UO_278 (O_278,N_29797,N_29923);
xnor UO_279 (O_279,N_29923,N_29890);
xor UO_280 (O_280,N_29638,N_29671);
nand UO_281 (O_281,N_29506,N_29585);
and UO_282 (O_282,N_29801,N_29520);
or UO_283 (O_283,N_29697,N_29761);
xnor UO_284 (O_284,N_29763,N_29634);
and UO_285 (O_285,N_29772,N_29877);
and UO_286 (O_286,N_29514,N_29694);
xor UO_287 (O_287,N_29734,N_29798);
nand UO_288 (O_288,N_29736,N_29878);
and UO_289 (O_289,N_29563,N_29929);
nor UO_290 (O_290,N_29647,N_29888);
nand UO_291 (O_291,N_29814,N_29859);
or UO_292 (O_292,N_29731,N_29766);
xor UO_293 (O_293,N_29549,N_29862);
and UO_294 (O_294,N_29630,N_29860);
nor UO_295 (O_295,N_29687,N_29940);
nand UO_296 (O_296,N_29550,N_29669);
xnor UO_297 (O_297,N_29502,N_29686);
xnor UO_298 (O_298,N_29882,N_29635);
nand UO_299 (O_299,N_29788,N_29632);
xnor UO_300 (O_300,N_29800,N_29917);
xor UO_301 (O_301,N_29631,N_29882);
and UO_302 (O_302,N_29578,N_29846);
xnor UO_303 (O_303,N_29960,N_29777);
and UO_304 (O_304,N_29893,N_29636);
xor UO_305 (O_305,N_29838,N_29572);
and UO_306 (O_306,N_29924,N_29970);
nor UO_307 (O_307,N_29996,N_29857);
xor UO_308 (O_308,N_29823,N_29854);
nand UO_309 (O_309,N_29948,N_29660);
nand UO_310 (O_310,N_29594,N_29693);
xnor UO_311 (O_311,N_29582,N_29737);
or UO_312 (O_312,N_29697,N_29796);
and UO_313 (O_313,N_29513,N_29506);
nand UO_314 (O_314,N_29536,N_29671);
and UO_315 (O_315,N_29663,N_29755);
and UO_316 (O_316,N_29611,N_29641);
nor UO_317 (O_317,N_29728,N_29520);
and UO_318 (O_318,N_29576,N_29811);
nand UO_319 (O_319,N_29624,N_29726);
nand UO_320 (O_320,N_29960,N_29781);
or UO_321 (O_321,N_29717,N_29680);
nor UO_322 (O_322,N_29630,N_29941);
nand UO_323 (O_323,N_29821,N_29623);
and UO_324 (O_324,N_29953,N_29529);
nand UO_325 (O_325,N_29853,N_29658);
xnor UO_326 (O_326,N_29644,N_29793);
and UO_327 (O_327,N_29686,N_29885);
nand UO_328 (O_328,N_29923,N_29678);
or UO_329 (O_329,N_29630,N_29676);
or UO_330 (O_330,N_29982,N_29611);
or UO_331 (O_331,N_29725,N_29794);
or UO_332 (O_332,N_29826,N_29756);
or UO_333 (O_333,N_29526,N_29974);
nor UO_334 (O_334,N_29785,N_29827);
nor UO_335 (O_335,N_29826,N_29558);
xor UO_336 (O_336,N_29653,N_29954);
or UO_337 (O_337,N_29855,N_29938);
nand UO_338 (O_338,N_29951,N_29922);
xor UO_339 (O_339,N_29790,N_29528);
or UO_340 (O_340,N_29881,N_29528);
nor UO_341 (O_341,N_29543,N_29710);
xnor UO_342 (O_342,N_29808,N_29956);
and UO_343 (O_343,N_29920,N_29588);
or UO_344 (O_344,N_29688,N_29645);
nor UO_345 (O_345,N_29535,N_29556);
and UO_346 (O_346,N_29957,N_29870);
and UO_347 (O_347,N_29648,N_29526);
xor UO_348 (O_348,N_29645,N_29618);
or UO_349 (O_349,N_29770,N_29618);
xnor UO_350 (O_350,N_29692,N_29516);
or UO_351 (O_351,N_29503,N_29518);
nor UO_352 (O_352,N_29713,N_29904);
and UO_353 (O_353,N_29800,N_29558);
nand UO_354 (O_354,N_29725,N_29811);
and UO_355 (O_355,N_29894,N_29847);
nor UO_356 (O_356,N_29781,N_29520);
and UO_357 (O_357,N_29738,N_29926);
or UO_358 (O_358,N_29695,N_29677);
xor UO_359 (O_359,N_29731,N_29707);
and UO_360 (O_360,N_29845,N_29839);
and UO_361 (O_361,N_29702,N_29968);
and UO_362 (O_362,N_29579,N_29944);
xnor UO_363 (O_363,N_29510,N_29981);
nand UO_364 (O_364,N_29717,N_29743);
or UO_365 (O_365,N_29736,N_29629);
nor UO_366 (O_366,N_29704,N_29661);
nand UO_367 (O_367,N_29657,N_29884);
nor UO_368 (O_368,N_29564,N_29845);
nor UO_369 (O_369,N_29932,N_29993);
and UO_370 (O_370,N_29890,N_29952);
nand UO_371 (O_371,N_29797,N_29697);
or UO_372 (O_372,N_29777,N_29964);
xor UO_373 (O_373,N_29850,N_29685);
nand UO_374 (O_374,N_29614,N_29639);
and UO_375 (O_375,N_29764,N_29891);
xnor UO_376 (O_376,N_29534,N_29883);
nor UO_377 (O_377,N_29506,N_29893);
or UO_378 (O_378,N_29598,N_29757);
or UO_379 (O_379,N_29562,N_29695);
and UO_380 (O_380,N_29838,N_29530);
or UO_381 (O_381,N_29997,N_29993);
or UO_382 (O_382,N_29757,N_29535);
xnor UO_383 (O_383,N_29600,N_29715);
xnor UO_384 (O_384,N_29534,N_29901);
and UO_385 (O_385,N_29563,N_29652);
nor UO_386 (O_386,N_29830,N_29756);
or UO_387 (O_387,N_29635,N_29935);
xor UO_388 (O_388,N_29785,N_29547);
xor UO_389 (O_389,N_29628,N_29877);
and UO_390 (O_390,N_29575,N_29614);
nand UO_391 (O_391,N_29540,N_29687);
or UO_392 (O_392,N_29948,N_29522);
nand UO_393 (O_393,N_29599,N_29701);
nand UO_394 (O_394,N_29827,N_29840);
and UO_395 (O_395,N_29536,N_29787);
nand UO_396 (O_396,N_29834,N_29718);
xor UO_397 (O_397,N_29779,N_29982);
nor UO_398 (O_398,N_29969,N_29931);
and UO_399 (O_399,N_29768,N_29501);
and UO_400 (O_400,N_29517,N_29615);
or UO_401 (O_401,N_29715,N_29958);
or UO_402 (O_402,N_29890,N_29745);
and UO_403 (O_403,N_29828,N_29529);
or UO_404 (O_404,N_29633,N_29528);
nor UO_405 (O_405,N_29904,N_29621);
and UO_406 (O_406,N_29561,N_29967);
or UO_407 (O_407,N_29721,N_29893);
or UO_408 (O_408,N_29631,N_29822);
or UO_409 (O_409,N_29688,N_29596);
xnor UO_410 (O_410,N_29956,N_29901);
nand UO_411 (O_411,N_29849,N_29703);
nor UO_412 (O_412,N_29529,N_29768);
and UO_413 (O_413,N_29909,N_29772);
xor UO_414 (O_414,N_29828,N_29701);
xor UO_415 (O_415,N_29931,N_29627);
nor UO_416 (O_416,N_29711,N_29908);
nand UO_417 (O_417,N_29565,N_29530);
xor UO_418 (O_418,N_29792,N_29875);
xor UO_419 (O_419,N_29639,N_29787);
or UO_420 (O_420,N_29560,N_29915);
xor UO_421 (O_421,N_29571,N_29786);
nor UO_422 (O_422,N_29991,N_29730);
xor UO_423 (O_423,N_29902,N_29512);
xnor UO_424 (O_424,N_29523,N_29747);
and UO_425 (O_425,N_29928,N_29509);
or UO_426 (O_426,N_29565,N_29598);
or UO_427 (O_427,N_29642,N_29607);
and UO_428 (O_428,N_29691,N_29982);
and UO_429 (O_429,N_29770,N_29775);
nand UO_430 (O_430,N_29956,N_29843);
and UO_431 (O_431,N_29773,N_29703);
nand UO_432 (O_432,N_29846,N_29607);
or UO_433 (O_433,N_29546,N_29658);
and UO_434 (O_434,N_29610,N_29771);
nor UO_435 (O_435,N_29672,N_29889);
nand UO_436 (O_436,N_29680,N_29583);
or UO_437 (O_437,N_29708,N_29721);
or UO_438 (O_438,N_29961,N_29659);
or UO_439 (O_439,N_29697,N_29965);
nor UO_440 (O_440,N_29989,N_29921);
and UO_441 (O_441,N_29808,N_29928);
nand UO_442 (O_442,N_29951,N_29816);
xor UO_443 (O_443,N_29575,N_29720);
or UO_444 (O_444,N_29547,N_29557);
xor UO_445 (O_445,N_29722,N_29891);
nor UO_446 (O_446,N_29988,N_29977);
or UO_447 (O_447,N_29984,N_29775);
or UO_448 (O_448,N_29896,N_29978);
and UO_449 (O_449,N_29899,N_29889);
and UO_450 (O_450,N_29533,N_29985);
or UO_451 (O_451,N_29551,N_29894);
and UO_452 (O_452,N_29823,N_29765);
nor UO_453 (O_453,N_29802,N_29757);
nand UO_454 (O_454,N_29539,N_29823);
or UO_455 (O_455,N_29963,N_29717);
and UO_456 (O_456,N_29871,N_29775);
or UO_457 (O_457,N_29765,N_29852);
xnor UO_458 (O_458,N_29960,N_29790);
xor UO_459 (O_459,N_29654,N_29665);
or UO_460 (O_460,N_29590,N_29880);
and UO_461 (O_461,N_29825,N_29829);
nor UO_462 (O_462,N_29954,N_29551);
xor UO_463 (O_463,N_29734,N_29781);
xnor UO_464 (O_464,N_29797,N_29576);
nand UO_465 (O_465,N_29937,N_29500);
and UO_466 (O_466,N_29639,N_29840);
nor UO_467 (O_467,N_29595,N_29638);
nor UO_468 (O_468,N_29843,N_29566);
or UO_469 (O_469,N_29991,N_29680);
nor UO_470 (O_470,N_29602,N_29639);
or UO_471 (O_471,N_29714,N_29589);
xnor UO_472 (O_472,N_29517,N_29916);
xor UO_473 (O_473,N_29929,N_29943);
or UO_474 (O_474,N_29767,N_29613);
and UO_475 (O_475,N_29730,N_29808);
or UO_476 (O_476,N_29912,N_29545);
xor UO_477 (O_477,N_29684,N_29760);
nand UO_478 (O_478,N_29702,N_29943);
xor UO_479 (O_479,N_29564,N_29599);
xor UO_480 (O_480,N_29939,N_29910);
nor UO_481 (O_481,N_29644,N_29953);
or UO_482 (O_482,N_29698,N_29683);
nand UO_483 (O_483,N_29562,N_29812);
or UO_484 (O_484,N_29887,N_29866);
nand UO_485 (O_485,N_29669,N_29590);
nand UO_486 (O_486,N_29723,N_29782);
nand UO_487 (O_487,N_29609,N_29721);
and UO_488 (O_488,N_29962,N_29576);
or UO_489 (O_489,N_29956,N_29748);
nand UO_490 (O_490,N_29891,N_29924);
nor UO_491 (O_491,N_29917,N_29874);
or UO_492 (O_492,N_29900,N_29731);
nand UO_493 (O_493,N_29861,N_29500);
or UO_494 (O_494,N_29860,N_29522);
and UO_495 (O_495,N_29972,N_29581);
nor UO_496 (O_496,N_29667,N_29993);
or UO_497 (O_497,N_29664,N_29555);
nand UO_498 (O_498,N_29882,N_29715);
nor UO_499 (O_499,N_29657,N_29619);
nand UO_500 (O_500,N_29889,N_29929);
xnor UO_501 (O_501,N_29633,N_29512);
and UO_502 (O_502,N_29985,N_29939);
nand UO_503 (O_503,N_29957,N_29530);
nand UO_504 (O_504,N_29617,N_29858);
or UO_505 (O_505,N_29945,N_29979);
and UO_506 (O_506,N_29677,N_29574);
xor UO_507 (O_507,N_29712,N_29957);
xnor UO_508 (O_508,N_29691,N_29559);
or UO_509 (O_509,N_29545,N_29904);
or UO_510 (O_510,N_29873,N_29673);
nand UO_511 (O_511,N_29829,N_29967);
or UO_512 (O_512,N_29736,N_29954);
or UO_513 (O_513,N_29859,N_29666);
or UO_514 (O_514,N_29501,N_29979);
or UO_515 (O_515,N_29817,N_29952);
and UO_516 (O_516,N_29975,N_29801);
and UO_517 (O_517,N_29557,N_29753);
and UO_518 (O_518,N_29768,N_29535);
xnor UO_519 (O_519,N_29683,N_29756);
xnor UO_520 (O_520,N_29783,N_29629);
nor UO_521 (O_521,N_29746,N_29667);
or UO_522 (O_522,N_29849,N_29652);
nor UO_523 (O_523,N_29524,N_29626);
and UO_524 (O_524,N_29661,N_29804);
and UO_525 (O_525,N_29923,N_29768);
nor UO_526 (O_526,N_29505,N_29674);
or UO_527 (O_527,N_29505,N_29663);
and UO_528 (O_528,N_29702,N_29769);
xor UO_529 (O_529,N_29894,N_29731);
nand UO_530 (O_530,N_29832,N_29640);
and UO_531 (O_531,N_29957,N_29756);
xnor UO_532 (O_532,N_29920,N_29506);
xor UO_533 (O_533,N_29675,N_29682);
nor UO_534 (O_534,N_29833,N_29826);
xor UO_535 (O_535,N_29589,N_29873);
nand UO_536 (O_536,N_29521,N_29939);
or UO_537 (O_537,N_29974,N_29874);
nand UO_538 (O_538,N_29636,N_29965);
or UO_539 (O_539,N_29784,N_29606);
nand UO_540 (O_540,N_29609,N_29962);
or UO_541 (O_541,N_29999,N_29865);
nor UO_542 (O_542,N_29592,N_29859);
xnor UO_543 (O_543,N_29621,N_29592);
and UO_544 (O_544,N_29539,N_29724);
xnor UO_545 (O_545,N_29544,N_29765);
and UO_546 (O_546,N_29571,N_29657);
or UO_547 (O_547,N_29765,N_29682);
nor UO_548 (O_548,N_29522,N_29942);
and UO_549 (O_549,N_29641,N_29531);
and UO_550 (O_550,N_29999,N_29974);
xor UO_551 (O_551,N_29720,N_29868);
or UO_552 (O_552,N_29823,N_29625);
and UO_553 (O_553,N_29659,N_29667);
nor UO_554 (O_554,N_29984,N_29840);
or UO_555 (O_555,N_29648,N_29604);
xor UO_556 (O_556,N_29747,N_29616);
and UO_557 (O_557,N_29918,N_29931);
or UO_558 (O_558,N_29820,N_29852);
xnor UO_559 (O_559,N_29689,N_29744);
nor UO_560 (O_560,N_29663,N_29874);
xnor UO_561 (O_561,N_29855,N_29884);
nor UO_562 (O_562,N_29522,N_29989);
and UO_563 (O_563,N_29722,N_29557);
nand UO_564 (O_564,N_29715,N_29708);
and UO_565 (O_565,N_29821,N_29613);
nor UO_566 (O_566,N_29936,N_29801);
nor UO_567 (O_567,N_29808,N_29990);
or UO_568 (O_568,N_29595,N_29850);
xnor UO_569 (O_569,N_29542,N_29981);
nor UO_570 (O_570,N_29867,N_29880);
or UO_571 (O_571,N_29961,N_29869);
xnor UO_572 (O_572,N_29956,N_29669);
nand UO_573 (O_573,N_29628,N_29507);
and UO_574 (O_574,N_29941,N_29806);
nor UO_575 (O_575,N_29752,N_29547);
and UO_576 (O_576,N_29645,N_29870);
xnor UO_577 (O_577,N_29858,N_29609);
nor UO_578 (O_578,N_29917,N_29523);
or UO_579 (O_579,N_29710,N_29960);
nor UO_580 (O_580,N_29519,N_29787);
nand UO_581 (O_581,N_29812,N_29641);
xnor UO_582 (O_582,N_29798,N_29655);
and UO_583 (O_583,N_29501,N_29763);
nor UO_584 (O_584,N_29635,N_29690);
xnor UO_585 (O_585,N_29669,N_29821);
nor UO_586 (O_586,N_29984,N_29740);
and UO_587 (O_587,N_29551,N_29861);
nand UO_588 (O_588,N_29859,N_29527);
or UO_589 (O_589,N_29923,N_29539);
nand UO_590 (O_590,N_29969,N_29674);
nand UO_591 (O_591,N_29697,N_29730);
nor UO_592 (O_592,N_29780,N_29905);
nor UO_593 (O_593,N_29725,N_29585);
or UO_594 (O_594,N_29650,N_29806);
nand UO_595 (O_595,N_29961,N_29899);
and UO_596 (O_596,N_29596,N_29829);
nand UO_597 (O_597,N_29792,N_29860);
xor UO_598 (O_598,N_29762,N_29601);
and UO_599 (O_599,N_29509,N_29954);
nor UO_600 (O_600,N_29636,N_29951);
nor UO_601 (O_601,N_29778,N_29825);
nor UO_602 (O_602,N_29865,N_29877);
nor UO_603 (O_603,N_29983,N_29604);
nor UO_604 (O_604,N_29923,N_29937);
nor UO_605 (O_605,N_29750,N_29589);
or UO_606 (O_606,N_29751,N_29959);
or UO_607 (O_607,N_29812,N_29847);
nand UO_608 (O_608,N_29698,N_29930);
and UO_609 (O_609,N_29856,N_29544);
and UO_610 (O_610,N_29721,N_29734);
or UO_611 (O_611,N_29544,N_29673);
or UO_612 (O_612,N_29849,N_29585);
nor UO_613 (O_613,N_29603,N_29930);
or UO_614 (O_614,N_29666,N_29682);
xor UO_615 (O_615,N_29561,N_29988);
and UO_616 (O_616,N_29654,N_29723);
nand UO_617 (O_617,N_29634,N_29672);
or UO_618 (O_618,N_29881,N_29710);
nor UO_619 (O_619,N_29611,N_29985);
xor UO_620 (O_620,N_29926,N_29625);
nor UO_621 (O_621,N_29938,N_29781);
xnor UO_622 (O_622,N_29589,N_29834);
and UO_623 (O_623,N_29544,N_29524);
nand UO_624 (O_624,N_29593,N_29687);
and UO_625 (O_625,N_29855,N_29750);
xnor UO_626 (O_626,N_29682,N_29789);
xnor UO_627 (O_627,N_29567,N_29889);
nor UO_628 (O_628,N_29866,N_29629);
nor UO_629 (O_629,N_29700,N_29585);
nor UO_630 (O_630,N_29529,N_29955);
nor UO_631 (O_631,N_29540,N_29896);
nand UO_632 (O_632,N_29501,N_29573);
nor UO_633 (O_633,N_29652,N_29957);
nand UO_634 (O_634,N_29506,N_29932);
or UO_635 (O_635,N_29706,N_29639);
xor UO_636 (O_636,N_29914,N_29909);
or UO_637 (O_637,N_29502,N_29977);
xor UO_638 (O_638,N_29869,N_29515);
nand UO_639 (O_639,N_29937,N_29839);
and UO_640 (O_640,N_29629,N_29745);
nor UO_641 (O_641,N_29810,N_29919);
or UO_642 (O_642,N_29543,N_29842);
and UO_643 (O_643,N_29590,N_29851);
xnor UO_644 (O_644,N_29899,N_29816);
nand UO_645 (O_645,N_29954,N_29506);
xnor UO_646 (O_646,N_29717,N_29905);
nand UO_647 (O_647,N_29689,N_29659);
nor UO_648 (O_648,N_29669,N_29711);
or UO_649 (O_649,N_29897,N_29968);
nor UO_650 (O_650,N_29517,N_29733);
and UO_651 (O_651,N_29600,N_29886);
xor UO_652 (O_652,N_29559,N_29943);
and UO_653 (O_653,N_29982,N_29938);
nand UO_654 (O_654,N_29784,N_29826);
and UO_655 (O_655,N_29844,N_29620);
and UO_656 (O_656,N_29823,N_29827);
nor UO_657 (O_657,N_29972,N_29850);
nand UO_658 (O_658,N_29922,N_29736);
nor UO_659 (O_659,N_29886,N_29919);
and UO_660 (O_660,N_29507,N_29696);
and UO_661 (O_661,N_29776,N_29644);
or UO_662 (O_662,N_29941,N_29932);
nand UO_663 (O_663,N_29893,N_29892);
nor UO_664 (O_664,N_29906,N_29638);
nor UO_665 (O_665,N_29651,N_29753);
or UO_666 (O_666,N_29845,N_29977);
xor UO_667 (O_667,N_29836,N_29620);
and UO_668 (O_668,N_29656,N_29507);
or UO_669 (O_669,N_29592,N_29736);
or UO_670 (O_670,N_29901,N_29648);
and UO_671 (O_671,N_29737,N_29919);
or UO_672 (O_672,N_29573,N_29648);
xor UO_673 (O_673,N_29873,N_29963);
or UO_674 (O_674,N_29705,N_29793);
nor UO_675 (O_675,N_29546,N_29794);
or UO_676 (O_676,N_29985,N_29814);
nor UO_677 (O_677,N_29984,N_29905);
xor UO_678 (O_678,N_29599,N_29981);
nand UO_679 (O_679,N_29746,N_29584);
and UO_680 (O_680,N_29653,N_29778);
nor UO_681 (O_681,N_29900,N_29885);
nand UO_682 (O_682,N_29660,N_29779);
xnor UO_683 (O_683,N_29607,N_29662);
nand UO_684 (O_684,N_29525,N_29748);
or UO_685 (O_685,N_29516,N_29519);
nand UO_686 (O_686,N_29688,N_29704);
or UO_687 (O_687,N_29628,N_29726);
and UO_688 (O_688,N_29516,N_29885);
nor UO_689 (O_689,N_29658,N_29920);
or UO_690 (O_690,N_29926,N_29857);
and UO_691 (O_691,N_29527,N_29639);
xnor UO_692 (O_692,N_29575,N_29825);
nor UO_693 (O_693,N_29991,N_29548);
nor UO_694 (O_694,N_29746,N_29768);
xnor UO_695 (O_695,N_29992,N_29552);
nand UO_696 (O_696,N_29891,N_29965);
and UO_697 (O_697,N_29603,N_29685);
nand UO_698 (O_698,N_29692,N_29697);
xor UO_699 (O_699,N_29984,N_29925);
nor UO_700 (O_700,N_29763,N_29527);
nor UO_701 (O_701,N_29631,N_29968);
nor UO_702 (O_702,N_29594,N_29512);
or UO_703 (O_703,N_29724,N_29512);
nor UO_704 (O_704,N_29595,N_29935);
nor UO_705 (O_705,N_29874,N_29881);
or UO_706 (O_706,N_29890,N_29577);
and UO_707 (O_707,N_29550,N_29512);
xor UO_708 (O_708,N_29772,N_29881);
xor UO_709 (O_709,N_29766,N_29726);
nor UO_710 (O_710,N_29860,N_29973);
and UO_711 (O_711,N_29744,N_29804);
or UO_712 (O_712,N_29732,N_29862);
nand UO_713 (O_713,N_29621,N_29594);
xnor UO_714 (O_714,N_29767,N_29701);
or UO_715 (O_715,N_29641,N_29685);
and UO_716 (O_716,N_29688,N_29816);
and UO_717 (O_717,N_29688,N_29655);
or UO_718 (O_718,N_29947,N_29854);
and UO_719 (O_719,N_29612,N_29574);
xnor UO_720 (O_720,N_29849,N_29634);
and UO_721 (O_721,N_29611,N_29832);
and UO_722 (O_722,N_29544,N_29633);
xor UO_723 (O_723,N_29555,N_29773);
nor UO_724 (O_724,N_29918,N_29750);
or UO_725 (O_725,N_29974,N_29514);
or UO_726 (O_726,N_29592,N_29668);
or UO_727 (O_727,N_29977,N_29633);
nand UO_728 (O_728,N_29833,N_29702);
nand UO_729 (O_729,N_29954,N_29533);
and UO_730 (O_730,N_29761,N_29817);
or UO_731 (O_731,N_29544,N_29979);
xnor UO_732 (O_732,N_29582,N_29636);
nor UO_733 (O_733,N_29775,N_29816);
nor UO_734 (O_734,N_29636,N_29864);
nor UO_735 (O_735,N_29651,N_29853);
or UO_736 (O_736,N_29956,N_29819);
or UO_737 (O_737,N_29947,N_29834);
and UO_738 (O_738,N_29934,N_29787);
nand UO_739 (O_739,N_29566,N_29693);
and UO_740 (O_740,N_29995,N_29819);
xor UO_741 (O_741,N_29768,N_29662);
or UO_742 (O_742,N_29762,N_29864);
and UO_743 (O_743,N_29940,N_29902);
nand UO_744 (O_744,N_29938,N_29608);
nor UO_745 (O_745,N_29642,N_29782);
xnor UO_746 (O_746,N_29578,N_29955);
or UO_747 (O_747,N_29719,N_29684);
or UO_748 (O_748,N_29850,N_29703);
and UO_749 (O_749,N_29517,N_29860);
and UO_750 (O_750,N_29706,N_29760);
nand UO_751 (O_751,N_29873,N_29666);
nand UO_752 (O_752,N_29904,N_29900);
xnor UO_753 (O_753,N_29540,N_29676);
nor UO_754 (O_754,N_29819,N_29644);
xor UO_755 (O_755,N_29668,N_29971);
nand UO_756 (O_756,N_29948,N_29658);
or UO_757 (O_757,N_29830,N_29781);
nor UO_758 (O_758,N_29506,N_29668);
nand UO_759 (O_759,N_29699,N_29582);
and UO_760 (O_760,N_29746,N_29907);
xor UO_761 (O_761,N_29890,N_29965);
nand UO_762 (O_762,N_29640,N_29664);
and UO_763 (O_763,N_29895,N_29737);
nand UO_764 (O_764,N_29884,N_29826);
xnor UO_765 (O_765,N_29674,N_29609);
xnor UO_766 (O_766,N_29672,N_29970);
or UO_767 (O_767,N_29883,N_29662);
and UO_768 (O_768,N_29661,N_29561);
and UO_769 (O_769,N_29595,N_29578);
xor UO_770 (O_770,N_29866,N_29710);
or UO_771 (O_771,N_29615,N_29745);
and UO_772 (O_772,N_29757,N_29914);
nor UO_773 (O_773,N_29653,N_29930);
and UO_774 (O_774,N_29529,N_29982);
xnor UO_775 (O_775,N_29684,N_29505);
nand UO_776 (O_776,N_29505,N_29854);
nor UO_777 (O_777,N_29689,N_29911);
xor UO_778 (O_778,N_29615,N_29981);
nand UO_779 (O_779,N_29722,N_29858);
or UO_780 (O_780,N_29531,N_29955);
or UO_781 (O_781,N_29884,N_29755);
xnor UO_782 (O_782,N_29859,N_29630);
or UO_783 (O_783,N_29703,N_29513);
nor UO_784 (O_784,N_29530,N_29730);
nand UO_785 (O_785,N_29772,N_29791);
or UO_786 (O_786,N_29898,N_29743);
and UO_787 (O_787,N_29893,N_29936);
xnor UO_788 (O_788,N_29821,N_29943);
xor UO_789 (O_789,N_29835,N_29895);
and UO_790 (O_790,N_29887,N_29511);
or UO_791 (O_791,N_29620,N_29526);
xor UO_792 (O_792,N_29606,N_29934);
and UO_793 (O_793,N_29581,N_29550);
nor UO_794 (O_794,N_29646,N_29653);
nand UO_795 (O_795,N_29903,N_29769);
or UO_796 (O_796,N_29680,N_29516);
xnor UO_797 (O_797,N_29945,N_29914);
xor UO_798 (O_798,N_29778,N_29510);
nor UO_799 (O_799,N_29522,N_29689);
nand UO_800 (O_800,N_29543,N_29506);
nand UO_801 (O_801,N_29836,N_29608);
nand UO_802 (O_802,N_29505,N_29783);
nand UO_803 (O_803,N_29645,N_29805);
nor UO_804 (O_804,N_29703,N_29951);
xor UO_805 (O_805,N_29556,N_29560);
and UO_806 (O_806,N_29651,N_29883);
nand UO_807 (O_807,N_29559,N_29605);
nor UO_808 (O_808,N_29636,N_29743);
or UO_809 (O_809,N_29964,N_29612);
xor UO_810 (O_810,N_29648,N_29753);
or UO_811 (O_811,N_29902,N_29621);
nor UO_812 (O_812,N_29876,N_29834);
and UO_813 (O_813,N_29551,N_29700);
xor UO_814 (O_814,N_29538,N_29633);
xnor UO_815 (O_815,N_29642,N_29905);
or UO_816 (O_816,N_29611,N_29737);
nand UO_817 (O_817,N_29869,N_29637);
xor UO_818 (O_818,N_29644,N_29595);
xnor UO_819 (O_819,N_29838,N_29805);
and UO_820 (O_820,N_29962,N_29553);
nand UO_821 (O_821,N_29968,N_29526);
nand UO_822 (O_822,N_29595,N_29549);
nand UO_823 (O_823,N_29970,N_29593);
xnor UO_824 (O_824,N_29527,N_29598);
nand UO_825 (O_825,N_29710,N_29697);
nand UO_826 (O_826,N_29872,N_29614);
nand UO_827 (O_827,N_29976,N_29602);
nor UO_828 (O_828,N_29512,N_29631);
and UO_829 (O_829,N_29789,N_29544);
nand UO_830 (O_830,N_29954,N_29914);
nor UO_831 (O_831,N_29795,N_29631);
nor UO_832 (O_832,N_29885,N_29789);
nor UO_833 (O_833,N_29942,N_29956);
or UO_834 (O_834,N_29577,N_29773);
nand UO_835 (O_835,N_29926,N_29575);
xor UO_836 (O_836,N_29584,N_29965);
xnor UO_837 (O_837,N_29703,N_29950);
xor UO_838 (O_838,N_29864,N_29683);
and UO_839 (O_839,N_29641,N_29900);
or UO_840 (O_840,N_29825,N_29616);
xor UO_841 (O_841,N_29840,N_29738);
xor UO_842 (O_842,N_29879,N_29728);
nand UO_843 (O_843,N_29820,N_29602);
xnor UO_844 (O_844,N_29657,N_29999);
and UO_845 (O_845,N_29660,N_29715);
nor UO_846 (O_846,N_29780,N_29554);
xor UO_847 (O_847,N_29870,N_29928);
and UO_848 (O_848,N_29939,N_29647);
nand UO_849 (O_849,N_29838,N_29676);
nand UO_850 (O_850,N_29702,N_29804);
nand UO_851 (O_851,N_29725,N_29693);
nor UO_852 (O_852,N_29901,N_29792);
and UO_853 (O_853,N_29739,N_29720);
nand UO_854 (O_854,N_29585,N_29872);
or UO_855 (O_855,N_29965,N_29542);
nand UO_856 (O_856,N_29688,N_29666);
and UO_857 (O_857,N_29937,N_29871);
or UO_858 (O_858,N_29989,N_29726);
and UO_859 (O_859,N_29568,N_29954);
nand UO_860 (O_860,N_29701,N_29542);
xor UO_861 (O_861,N_29620,N_29954);
and UO_862 (O_862,N_29909,N_29782);
nor UO_863 (O_863,N_29997,N_29662);
nand UO_864 (O_864,N_29873,N_29903);
xnor UO_865 (O_865,N_29986,N_29582);
nor UO_866 (O_866,N_29591,N_29526);
and UO_867 (O_867,N_29715,N_29959);
xnor UO_868 (O_868,N_29953,N_29527);
xor UO_869 (O_869,N_29501,N_29679);
nor UO_870 (O_870,N_29569,N_29848);
nand UO_871 (O_871,N_29782,N_29777);
xor UO_872 (O_872,N_29635,N_29699);
and UO_873 (O_873,N_29599,N_29730);
nor UO_874 (O_874,N_29867,N_29542);
and UO_875 (O_875,N_29631,N_29641);
xnor UO_876 (O_876,N_29641,N_29724);
xor UO_877 (O_877,N_29944,N_29560);
xnor UO_878 (O_878,N_29668,N_29683);
nor UO_879 (O_879,N_29517,N_29826);
nor UO_880 (O_880,N_29969,N_29960);
or UO_881 (O_881,N_29842,N_29671);
and UO_882 (O_882,N_29857,N_29960);
or UO_883 (O_883,N_29919,N_29569);
or UO_884 (O_884,N_29500,N_29875);
or UO_885 (O_885,N_29625,N_29827);
nor UO_886 (O_886,N_29970,N_29835);
and UO_887 (O_887,N_29528,N_29973);
and UO_888 (O_888,N_29656,N_29539);
xor UO_889 (O_889,N_29676,N_29828);
nor UO_890 (O_890,N_29643,N_29947);
nor UO_891 (O_891,N_29632,N_29655);
xor UO_892 (O_892,N_29569,N_29854);
nor UO_893 (O_893,N_29922,N_29974);
or UO_894 (O_894,N_29532,N_29982);
xnor UO_895 (O_895,N_29783,N_29592);
nand UO_896 (O_896,N_29871,N_29598);
nor UO_897 (O_897,N_29885,N_29698);
xnor UO_898 (O_898,N_29950,N_29973);
nand UO_899 (O_899,N_29874,N_29832);
and UO_900 (O_900,N_29954,N_29503);
xnor UO_901 (O_901,N_29700,N_29932);
and UO_902 (O_902,N_29552,N_29757);
nand UO_903 (O_903,N_29898,N_29542);
and UO_904 (O_904,N_29749,N_29964);
and UO_905 (O_905,N_29617,N_29789);
and UO_906 (O_906,N_29512,N_29943);
or UO_907 (O_907,N_29808,N_29702);
nand UO_908 (O_908,N_29857,N_29652);
nand UO_909 (O_909,N_29647,N_29830);
xnor UO_910 (O_910,N_29935,N_29711);
nor UO_911 (O_911,N_29923,N_29576);
or UO_912 (O_912,N_29835,N_29714);
and UO_913 (O_913,N_29657,N_29803);
nor UO_914 (O_914,N_29711,N_29970);
nand UO_915 (O_915,N_29539,N_29753);
or UO_916 (O_916,N_29524,N_29665);
nand UO_917 (O_917,N_29631,N_29806);
xor UO_918 (O_918,N_29790,N_29869);
or UO_919 (O_919,N_29691,N_29779);
nor UO_920 (O_920,N_29762,N_29885);
nor UO_921 (O_921,N_29586,N_29556);
or UO_922 (O_922,N_29798,N_29602);
nor UO_923 (O_923,N_29502,N_29646);
and UO_924 (O_924,N_29684,N_29941);
and UO_925 (O_925,N_29520,N_29624);
nand UO_926 (O_926,N_29885,N_29718);
and UO_927 (O_927,N_29971,N_29682);
nand UO_928 (O_928,N_29568,N_29577);
xor UO_929 (O_929,N_29890,N_29663);
or UO_930 (O_930,N_29852,N_29562);
or UO_931 (O_931,N_29802,N_29931);
or UO_932 (O_932,N_29888,N_29968);
nor UO_933 (O_933,N_29957,N_29789);
nand UO_934 (O_934,N_29990,N_29874);
xor UO_935 (O_935,N_29612,N_29634);
nor UO_936 (O_936,N_29844,N_29664);
and UO_937 (O_937,N_29706,N_29671);
and UO_938 (O_938,N_29637,N_29771);
nor UO_939 (O_939,N_29742,N_29798);
nor UO_940 (O_940,N_29865,N_29869);
or UO_941 (O_941,N_29542,N_29948);
nand UO_942 (O_942,N_29731,N_29557);
nand UO_943 (O_943,N_29501,N_29855);
nand UO_944 (O_944,N_29756,N_29595);
and UO_945 (O_945,N_29864,N_29916);
nor UO_946 (O_946,N_29541,N_29944);
nand UO_947 (O_947,N_29892,N_29623);
or UO_948 (O_948,N_29775,N_29843);
xor UO_949 (O_949,N_29566,N_29671);
nand UO_950 (O_950,N_29541,N_29709);
and UO_951 (O_951,N_29707,N_29753);
nor UO_952 (O_952,N_29908,N_29882);
xor UO_953 (O_953,N_29907,N_29924);
xnor UO_954 (O_954,N_29940,N_29578);
and UO_955 (O_955,N_29779,N_29636);
xnor UO_956 (O_956,N_29783,N_29915);
and UO_957 (O_957,N_29572,N_29649);
nor UO_958 (O_958,N_29699,N_29502);
and UO_959 (O_959,N_29902,N_29801);
nand UO_960 (O_960,N_29621,N_29719);
nor UO_961 (O_961,N_29635,N_29590);
nand UO_962 (O_962,N_29809,N_29824);
and UO_963 (O_963,N_29862,N_29906);
nand UO_964 (O_964,N_29585,N_29688);
nor UO_965 (O_965,N_29849,N_29982);
or UO_966 (O_966,N_29575,N_29781);
or UO_967 (O_967,N_29966,N_29943);
or UO_968 (O_968,N_29965,N_29561);
or UO_969 (O_969,N_29846,N_29898);
nor UO_970 (O_970,N_29946,N_29573);
nor UO_971 (O_971,N_29527,N_29808);
and UO_972 (O_972,N_29870,N_29756);
and UO_973 (O_973,N_29735,N_29622);
and UO_974 (O_974,N_29676,N_29750);
or UO_975 (O_975,N_29613,N_29589);
nor UO_976 (O_976,N_29901,N_29724);
nor UO_977 (O_977,N_29554,N_29973);
nand UO_978 (O_978,N_29703,N_29843);
or UO_979 (O_979,N_29643,N_29966);
and UO_980 (O_980,N_29533,N_29784);
and UO_981 (O_981,N_29889,N_29861);
or UO_982 (O_982,N_29614,N_29593);
xnor UO_983 (O_983,N_29794,N_29909);
nor UO_984 (O_984,N_29506,N_29656);
or UO_985 (O_985,N_29916,N_29737);
xnor UO_986 (O_986,N_29588,N_29636);
or UO_987 (O_987,N_29974,N_29908);
and UO_988 (O_988,N_29961,N_29661);
nand UO_989 (O_989,N_29755,N_29907);
nand UO_990 (O_990,N_29631,N_29679);
and UO_991 (O_991,N_29629,N_29833);
nor UO_992 (O_992,N_29746,N_29751);
and UO_993 (O_993,N_29674,N_29858);
nor UO_994 (O_994,N_29500,N_29578);
and UO_995 (O_995,N_29970,N_29849);
xnor UO_996 (O_996,N_29961,N_29598);
nand UO_997 (O_997,N_29944,N_29994);
or UO_998 (O_998,N_29964,N_29869);
nand UO_999 (O_999,N_29886,N_29525);
nor UO_1000 (O_1000,N_29591,N_29881);
nand UO_1001 (O_1001,N_29807,N_29739);
nand UO_1002 (O_1002,N_29829,N_29811);
or UO_1003 (O_1003,N_29507,N_29780);
or UO_1004 (O_1004,N_29882,N_29563);
xnor UO_1005 (O_1005,N_29828,N_29621);
nor UO_1006 (O_1006,N_29715,N_29996);
or UO_1007 (O_1007,N_29768,N_29683);
or UO_1008 (O_1008,N_29875,N_29888);
and UO_1009 (O_1009,N_29988,N_29594);
xor UO_1010 (O_1010,N_29666,N_29691);
nor UO_1011 (O_1011,N_29513,N_29882);
nand UO_1012 (O_1012,N_29835,N_29681);
xnor UO_1013 (O_1013,N_29824,N_29710);
and UO_1014 (O_1014,N_29862,N_29836);
and UO_1015 (O_1015,N_29824,N_29896);
nand UO_1016 (O_1016,N_29856,N_29725);
nor UO_1017 (O_1017,N_29974,N_29724);
nand UO_1018 (O_1018,N_29626,N_29938);
nand UO_1019 (O_1019,N_29887,N_29599);
nor UO_1020 (O_1020,N_29860,N_29735);
and UO_1021 (O_1021,N_29972,N_29823);
xor UO_1022 (O_1022,N_29822,N_29956);
nand UO_1023 (O_1023,N_29710,N_29859);
nand UO_1024 (O_1024,N_29860,N_29869);
or UO_1025 (O_1025,N_29953,N_29923);
nand UO_1026 (O_1026,N_29518,N_29777);
nand UO_1027 (O_1027,N_29822,N_29873);
and UO_1028 (O_1028,N_29766,N_29757);
and UO_1029 (O_1029,N_29792,N_29797);
or UO_1030 (O_1030,N_29533,N_29780);
or UO_1031 (O_1031,N_29931,N_29944);
or UO_1032 (O_1032,N_29904,N_29843);
nand UO_1033 (O_1033,N_29928,N_29820);
xnor UO_1034 (O_1034,N_29618,N_29740);
xnor UO_1035 (O_1035,N_29613,N_29988);
nor UO_1036 (O_1036,N_29550,N_29825);
nand UO_1037 (O_1037,N_29818,N_29975);
xor UO_1038 (O_1038,N_29595,N_29537);
and UO_1039 (O_1039,N_29845,N_29975);
xor UO_1040 (O_1040,N_29880,N_29512);
and UO_1041 (O_1041,N_29557,N_29628);
xor UO_1042 (O_1042,N_29534,N_29827);
xnor UO_1043 (O_1043,N_29799,N_29796);
and UO_1044 (O_1044,N_29994,N_29523);
nand UO_1045 (O_1045,N_29700,N_29759);
nand UO_1046 (O_1046,N_29975,N_29715);
and UO_1047 (O_1047,N_29838,N_29915);
nor UO_1048 (O_1048,N_29724,N_29669);
and UO_1049 (O_1049,N_29518,N_29986);
and UO_1050 (O_1050,N_29920,N_29928);
nand UO_1051 (O_1051,N_29796,N_29875);
and UO_1052 (O_1052,N_29666,N_29966);
and UO_1053 (O_1053,N_29587,N_29608);
nand UO_1054 (O_1054,N_29948,N_29644);
xor UO_1055 (O_1055,N_29873,N_29574);
and UO_1056 (O_1056,N_29555,N_29684);
nand UO_1057 (O_1057,N_29735,N_29743);
and UO_1058 (O_1058,N_29518,N_29864);
nor UO_1059 (O_1059,N_29835,N_29906);
and UO_1060 (O_1060,N_29898,N_29847);
or UO_1061 (O_1061,N_29930,N_29816);
nand UO_1062 (O_1062,N_29793,N_29809);
and UO_1063 (O_1063,N_29869,N_29831);
nor UO_1064 (O_1064,N_29996,N_29834);
or UO_1065 (O_1065,N_29516,N_29947);
nor UO_1066 (O_1066,N_29722,N_29762);
and UO_1067 (O_1067,N_29724,N_29790);
and UO_1068 (O_1068,N_29712,N_29660);
or UO_1069 (O_1069,N_29926,N_29886);
nor UO_1070 (O_1070,N_29964,N_29602);
xor UO_1071 (O_1071,N_29674,N_29967);
nor UO_1072 (O_1072,N_29560,N_29528);
or UO_1073 (O_1073,N_29972,N_29763);
and UO_1074 (O_1074,N_29966,N_29601);
xor UO_1075 (O_1075,N_29615,N_29942);
and UO_1076 (O_1076,N_29634,N_29520);
and UO_1077 (O_1077,N_29976,N_29958);
and UO_1078 (O_1078,N_29561,N_29654);
and UO_1079 (O_1079,N_29766,N_29793);
nor UO_1080 (O_1080,N_29644,N_29610);
nor UO_1081 (O_1081,N_29930,N_29951);
or UO_1082 (O_1082,N_29594,N_29967);
or UO_1083 (O_1083,N_29894,N_29514);
and UO_1084 (O_1084,N_29764,N_29628);
xnor UO_1085 (O_1085,N_29845,N_29543);
nand UO_1086 (O_1086,N_29978,N_29674);
nor UO_1087 (O_1087,N_29562,N_29731);
nor UO_1088 (O_1088,N_29692,N_29747);
or UO_1089 (O_1089,N_29761,N_29795);
xnor UO_1090 (O_1090,N_29768,N_29668);
nand UO_1091 (O_1091,N_29516,N_29772);
xnor UO_1092 (O_1092,N_29702,N_29835);
nor UO_1093 (O_1093,N_29868,N_29617);
and UO_1094 (O_1094,N_29721,N_29682);
nor UO_1095 (O_1095,N_29694,N_29669);
or UO_1096 (O_1096,N_29783,N_29622);
and UO_1097 (O_1097,N_29871,N_29902);
nor UO_1098 (O_1098,N_29704,N_29675);
nand UO_1099 (O_1099,N_29696,N_29939);
nand UO_1100 (O_1100,N_29807,N_29854);
nand UO_1101 (O_1101,N_29542,N_29731);
xnor UO_1102 (O_1102,N_29885,N_29586);
xnor UO_1103 (O_1103,N_29918,N_29546);
and UO_1104 (O_1104,N_29689,N_29738);
nand UO_1105 (O_1105,N_29896,N_29935);
xnor UO_1106 (O_1106,N_29990,N_29948);
nand UO_1107 (O_1107,N_29796,N_29791);
nand UO_1108 (O_1108,N_29959,N_29683);
nand UO_1109 (O_1109,N_29602,N_29938);
xnor UO_1110 (O_1110,N_29652,N_29771);
and UO_1111 (O_1111,N_29621,N_29711);
xor UO_1112 (O_1112,N_29597,N_29550);
xnor UO_1113 (O_1113,N_29514,N_29844);
nor UO_1114 (O_1114,N_29553,N_29788);
or UO_1115 (O_1115,N_29529,N_29682);
xnor UO_1116 (O_1116,N_29761,N_29513);
and UO_1117 (O_1117,N_29996,N_29811);
or UO_1118 (O_1118,N_29692,N_29566);
xor UO_1119 (O_1119,N_29544,N_29722);
nor UO_1120 (O_1120,N_29596,N_29782);
nor UO_1121 (O_1121,N_29510,N_29625);
and UO_1122 (O_1122,N_29924,N_29798);
nor UO_1123 (O_1123,N_29975,N_29860);
or UO_1124 (O_1124,N_29778,N_29500);
and UO_1125 (O_1125,N_29589,N_29938);
xor UO_1126 (O_1126,N_29692,N_29951);
or UO_1127 (O_1127,N_29537,N_29616);
nand UO_1128 (O_1128,N_29751,N_29996);
or UO_1129 (O_1129,N_29859,N_29891);
or UO_1130 (O_1130,N_29792,N_29921);
nor UO_1131 (O_1131,N_29720,N_29689);
xor UO_1132 (O_1132,N_29732,N_29701);
nor UO_1133 (O_1133,N_29811,N_29730);
or UO_1134 (O_1134,N_29554,N_29523);
nor UO_1135 (O_1135,N_29990,N_29736);
and UO_1136 (O_1136,N_29574,N_29502);
nor UO_1137 (O_1137,N_29553,N_29605);
xnor UO_1138 (O_1138,N_29808,N_29838);
xor UO_1139 (O_1139,N_29594,N_29569);
or UO_1140 (O_1140,N_29880,N_29924);
nand UO_1141 (O_1141,N_29751,N_29806);
and UO_1142 (O_1142,N_29848,N_29839);
nor UO_1143 (O_1143,N_29853,N_29612);
and UO_1144 (O_1144,N_29542,N_29839);
and UO_1145 (O_1145,N_29780,N_29930);
nor UO_1146 (O_1146,N_29689,N_29796);
and UO_1147 (O_1147,N_29919,N_29666);
xnor UO_1148 (O_1148,N_29548,N_29864);
xnor UO_1149 (O_1149,N_29550,N_29572);
xnor UO_1150 (O_1150,N_29642,N_29519);
and UO_1151 (O_1151,N_29888,N_29692);
nor UO_1152 (O_1152,N_29773,N_29520);
and UO_1153 (O_1153,N_29626,N_29899);
and UO_1154 (O_1154,N_29897,N_29668);
and UO_1155 (O_1155,N_29504,N_29683);
xor UO_1156 (O_1156,N_29560,N_29742);
or UO_1157 (O_1157,N_29630,N_29506);
xnor UO_1158 (O_1158,N_29778,N_29900);
nor UO_1159 (O_1159,N_29535,N_29893);
and UO_1160 (O_1160,N_29906,N_29719);
nor UO_1161 (O_1161,N_29943,N_29638);
nor UO_1162 (O_1162,N_29807,N_29516);
and UO_1163 (O_1163,N_29576,N_29506);
and UO_1164 (O_1164,N_29716,N_29839);
xnor UO_1165 (O_1165,N_29997,N_29684);
xor UO_1166 (O_1166,N_29986,N_29757);
or UO_1167 (O_1167,N_29692,N_29626);
xnor UO_1168 (O_1168,N_29600,N_29972);
or UO_1169 (O_1169,N_29971,N_29959);
nand UO_1170 (O_1170,N_29898,N_29795);
xnor UO_1171 (O_1171,N_29511,N_29827);
xor UO_1172 (O_1172,N_29861,N_29906);
xor UO_1173 (O_1173,N_29796,N_29712);
and UO_1174 (O_1174,N_29577,N_29586);
xor UO_1175 (O_1175,N_29912,N_29866);
nand UO_1176 (O_1176,N_29799,N_29933);
or UO_1177 (O_1177,N_29955,N_29945);
or UO_1178 (O_1178,N_29547,N_29888);
nor UO_1179 (O_1179,N_29893,N_29637);
xnor UO_1180 (O_1180,N_29690,N_29623);
nor UO_1181 (O_1181,N_29850,N_29782);
xor UO_1182 (O_1182,N_29924,N_29707);
and UO_1183 (O_1183,N_29910,N_29893);
and UO_1184 (O_1184,N_29614,N_29898);
nand UO_1185 (O_1185,N_29833,N_29791);
xor UO_1186 (O_1186,N_29629,N_29728);
or UO_1187 (O_1187,N_29833,N_29733);
xor UO_1188 (O_1188,N_29583,N_29526);
nand UO_1189 (O_1189,N_29549,N_29733);
nor UO_1190 (O_1190,N_29579,N_29732);
and UO_1191 (O_1191,N_29781,N_29564);
xnor UO_1192 (O_1192,N_29787,N_29876);
or UO_1193 (O_1193,N_29967,N_29832);
xor UO_1194 (O_1194,N_29949,N_29717);
nand UO_1195 (O_1195,N_29521,N_29537);
and UO_1196 (O_1196,N_29546,N_29688);
nand UO_1197 (O_1197,N_29533,N_29965);
nor UO_1198 (O_1198,N_29988,N_29823);
or UO_1199 (O_1199,N_29723,N_29587);
nor UO_1200 (O_1200,N_29951,N_29632);
xor UO_1201 (O_1201,N_29517,N_29750);
or UO_1202 (O_1202,N_29770,N_29829);
and UO_1203 (O_1203,N_29949,N_29522);
xnor UO_1204 (O_1204,N_29584,N_29909);
xnor UO_1205 (O_1205,N_29857,N_29693);
xnor UO_1206 (O_1206,N_29687,N_29917);
or UO_1207 (O_1207,N_29914,N_29653);
nand UO_1208 (O_1208,N_29929,N_29939);
or UO_1209 (O_1209,N_29597,N_29939);
nand UO_1210 (O_1210,N_29696,N_29982);
or UO_1211 (O_1211,N_29671,N_29539);
and UO_1212 (O_1212,N_29787,N_29515);
and UO_1213 (O_1213,N_29901,N_29965);
nor UO_1214 (O_1214,N_29676,N_29595);
nor UO_1215 (O_1215,N_29961,N_29914);
nor UO_1216 (O_1216,N_29954,N_29922);
nand UO_1217 (O_1217,N_29853,N_29794);
and UO_1218 (O_1218,N_29611,N_29515);
and UO_1219 (O_1219,N_29630,N_29823);
nor UO_1220 (O_1220,N_29725,N_29620);
and UO_1221 (O_1221,N_29865,N_29890);
or UO_1222 (O_1222,N_29737,N_29644);
xnor UO_1223 (O_1223,N_29594,N_29562);
xor UO_1224 (O_1224,N_29960,N_29622);
xnor UO_1225 (O_1225,N_29986,N_29893);
or UO_1226 (O_1226,N_29524,N_29937);
or UO_1227 (O_1227,N_29901,N_29846);
xnor UO_1228 (O_1228,N_29642,N_29812);
nand UO_1229 (O_1229,N_29531,N_29943);
or UO_1230 (O_1230,N_29755,N_29744);
nand UO_1231 (O_1231,N_29870,N_29524);
nor UO_1232 (O_1232,N_29523,N_29867);
xnor UO_1233 (O_1233,N_29724,N_29552);
or UO_1234 (O_1234,N_29569,N_29874);
or UO_1235 (O_1235,N_29585,N_29577);
and UO_1236 (O_1236,N_29882,N_29789);
xnor UO_1237 (O_1237,N_29696,N_29581);
nor UO_1238 (O_1238,N_29789,N_29513);
nor UO_1239 (O_1239,N_29873,N_29564);
nand UO_1240 (O_1240,N_29728,N_29876);
xor UO_1241 (O_1241,N_29880,N_29991);
xnor UO_1242 (O_1242,N_29556,N_29537);
or UO_1243 (O_1243,N_29719,N_29724);
xor UO_1244 (O_1244,N_29573,N_29971);
and UO_1245 (O_1245,N_29544,N_29964);
or UO_1246 (O_1246,N_29687,N_29781);
and UO_1247 (O_1247,N_29784,N_29925);
and UO_1248 (O_1248,N_29707,N_29806);
xnor UO_1249 (O_1249,N_29971,N_29690);
and UO_1250 (O_1250,N_29967,N_29940);
or UO_1251 (O_1251,N_29979,N_29973);
xnor UO_1252 (O_1252,N_29798,N_29669);
xnor UO_1253 (O_1253,N_29609,N_29704);
and UO_1254 (O_1254,N_29570,N_29815);
nor UO_1255 (O_1255,N_29980,N_29949);
xor UO_1256 (O_1256,N_29897,N_29951);
nor UO_1257 (O_1257,N_29955,N_29898);
xor UO_1258 (O_1258,N_29670,N_29597);
nand UO_1259 (O_1259,N_29875,N_29723);
xnor UO_1260 (O_1260,N_29712,N_29849);
and UO_1261 (O_1261,N_29766,N_29573);
or UO_1262 (O_1262,N_29620,N_29991);
nor UO_1263 (O_1263,N_29523,N_29778);
xor UO_1264 (O_1264,N_29712,N_29702);
and UO_1265 (O_1265,N_29980,N_29642);
nand UO_1266 (O_1266,N_29614,N_29772);
or UO_1267 (O_1267,N_29743,N_29904);
nor UO_1268 (O_1268,N_29516,N_29918);
or UO_1269 (O_1269,N_29916,N_29882);
nand UO_1270 (O_1270,N_29983,N_29867);
nand UO_1271 (O_1271,N_29843,N_29556);
or UO_1272 (O_1272,N_29501,N_29948);
xor UO_1273 (O_1273,N_29904,N_29615);
and UO_1274 (O_1274,N_29748,N_29762);
nor UO_1275 (O_1275,N_29561,N_29617);
nand UO_1276 (O_1276,N_29864,N_29556);
or UO_1277 (O_1277,N_29815,N_29709);
nand UO_1278 (O_1278,N_29692,N_29945);
xnor UO_1279 (O_1279,N_29601,N_29846);
or UO_1280 (O_1280,N_29590,N_29695);
xor UO_1281 (O_1281,N_29942,N_29714);
nor UO_1282 (O_1282,N_29660,N_29961);
xnor UO_1283 (O_1283,N_29659,N_29859);
and UO_1284 (O_1284,N_29918,N_29775);
or UO_1285 (O_1285,N_29896,N_29617);
nor UO_1286 (O_1286,N_29744,N_29571);
nor UO_1287 (O_1287,N_29962,N_29760);
nor UO_1288 (O_1288,N_29524,N_29815);
and UO_1289 (O_1289,N_29903,N_29942);
and UO_1290 (O_1290,N_29999,N_29734);
or UO_1291 (O_1291,N_29924,N_29836);
or UO_1292 (O_1292,N_29696,N_29952);
nor UO_1293 (O_1293,N_29704,N_29848);
or UO_1294 (O_1294,N_29666,N_29756);
nor UO_1295 (O_1295,N_29910,N_29811);
nand UO_1296 (O_1296,N_29502,N_29664);
nand UO_1297 (O_1297,N_29563,N_29857);
nor UO_1298 (O_1298,N_29567,N_29788);
xnor UO_1299 (O_1299,N_29850,N_29508);
or UO_1300 (O_1300,N_29806,N_29608);
or UO_1301 (O_1301,N_29694,N_29987);
or UO_1302 (O_1302,N_29667,N_29643);
nor UO_1303 (O_1303,N_29925,N_29616);
nor UO_1304 (O_1304,N_29966,N_29903);
xor UO_1305 (O_1305,N_29604,N_29784);
nor UO_1306 (O_1306,N_29714,N_29628);
nor UO_1307 (O_1307,N_29505,N_29514);
nor UO_1308 (O_1308,N_29749,N_29826);
nand UO_1309 (O_1309,N_29737,N_29965);
and UO_1310 (O_1310,N_29724,N_29702);
nand UO_1311 (O_1311,N_29996,N_29966);
or UO_1312 (O_1312,N_29754,N_29930);
xor UO_1313 (O_1313,N_29762,N_29661);
nor UO_1314 (O_1314,N_29816,N_29883);
or UO_1315 (O_1315,N_29567,N_29961);
nand UO_1316 (O_1316,N_29889,N_29656);
nand UO_1317 (O_1317,N_29703,N_29781);
nor UO_1318 (O_1318,N_29968,N_29614);
nor UO_1319 (O_1319,N_29679,N_29721);
nor UO_1320 (O_1320,N_29550,N_29595);
and UO_1321 (O_1321,N_29836,N_29510);
or UO_1322 (O_1322,N_29642,N_29752);
or UO_1323 (O_1323,N_29572,N_29892);
nand UO_1324 (O_1324,N_29952,N_29994);
xnor UO_1325 (O_1325,N_29947,N_29995);
xnor UO_1326 (O_1326,N_29942,N_29729);
nand UO_1327 (O_1327,N_29515,N_29769);
nand UO_1328 (O_1328,N_29959,N_29808);
xnor UO_1329 (O_1329,N_29721,N_29871);
xor UO_1330 (O_1330,N_29575,N_29786);
or UO_1331 (O_1331,N_29845,N_29769);
nor UO_1332 (O_1332,N_29657,N_29889);
or UO_1333 (O_1333,N_29819,N_29509);
and UO_1334 (O_1334,N_29677,N_29983);
xor UO_1335 (O_1335,N_29775,N_29742);
nor UO_1336 (O_1336,N_29911,N_29691);
xor UO_1337 (O_1337,N_29540,N_29824);
and UO_1338 (O_1338,N_29816,N_29734);
or UO_1339 (O_1339,N_29654,N_29861);
xnor UO_1340 (O_1340,N_29931,N_29852);
nand UO_1341 (O_1341,N_29982,N_29646);
and UO_1342 (O_1342,N_29576,N_29732);
xor UO_1343 (O_1343,N_29704,N_29756);
xor UO_1344 (O_1344,N_29707,N_29501);
or UO_1345 (O_1345,N_29647,N_29598);
and UO_1346 (O_1346,N_29970,N_29828);
or UO_1347 (O_1347,N_29850,N_29510);
nand UO_1348 (O_1348,N_29939,N_29758);
nand UO_1349 (O_1349,N_29671,N_29909);
or UO_1350 (O_1350,N_29702,N_29895);
and UO_1351 (O_1351,N_29918,N_29762);
nand UO_1352 (O_1352,N_29788,N_29535);
xnor UO_1353 (O_1353,N_29545,N_29634);
or UO_1354 (O_1354,N_29844,N_29867);
xor UO_1355 (O_1355,N_29866,N_29933);
xor UO_1356 (O_1356,N_29572,N_29756);
or UO_1357 (O_1357,N_29551,N_29616);
and UO_1358 (O_1358,N_29811,N_29632);
or UO_1359 (O_1359,N_29539,N_29622);
nor UO_1360 (O_1360,N_29804,N_29905);
nand UO_1361 (O_1361,N_29522,N_29751);
xor UO_1362 (O_1362,N_29904,N_29988);
and UO_1363 (O_1363,N_29685,N_29505);
xor UO_1364 (O_1364,N_29729,N_29508);
and UO_1365 (O_1365,N_29572,N_29843);
xor UO_1366 (O_1366,N_29624,N_29641);
nor UO_1367 (O_1367,N_29504,N_29567);
xnor UO_1368 (O_1368,N_29981,N_29909);
xnor UO_1369 (O_1369,N_29973,N_29551);
and UO_1370 (O_1370,N_29588,N_29892);
nor UO_1371 (O_1371,N_29906,N_29664);
nor UO_1372 (O_1372,N_29600,N_29657);
nor UO_1373 (O_1373,N_29599,N_29689);
xnor UO_1374 (O_1374,N_29697,N_29899);
and UO_1375 (O_1375,N_29834,N_29759);
or UO_1376 (O_1376,N_29995,N_29595);
nor UO_1377 (O_1377,N_29538,N_29827);
xor UO_1378 (O_1378,N_29934,N_29863);
nand UO_1379 (O_1379,N_29970,N_29773);
nor UO_1380 (O_1380,N_29831,N_29979);
nand UO_1381 (O_1381,N_29544,N_29641);
nor UO_1382 (O_1382,N_29625,N_29862);
and UO_1383 (O_1383,N_29676,N_29974);
and UO_1384 (O_1384,N_29504,N_29957);
nand UO_1385 (O_1385,N_29820,N_29751);
or UO_1386 (O_1386,N_29509,N_29573);
xnor UO_1387 (O_1387,N_29686,N_29511);
or UO_1388 (O_1388,N_29642,N_29845);
nand UO_1389 (O_1389,N_29955,N_29525);
or UO_1390 (O_1390,N_29789,N_29584);
or UO_1391 (O_1391,N_29983,N_29672);
xnor UO_1392 (O_1392,N_29533,N_29653);
and UO_1393 (O_1393,N_29521,N_29774);
nand UO_1394 (O_1394,N_29906,N_29525);
nor UO_1395 (O_1395,N_29601,N_29653);
nand UO_1396 (O_1396,N_29635,N_29996);
nand UO_1397 (O_1397,N_29891,N_29938);
and UO_1398 (O_1398,N_29511,N_29825);
nand UO_1399 (O_1399,N_29570,N_29507);
and UO_1400 (O_1400,N_29628,N_29585);
xnor UO_1401 (O_1401,N_29930,N_29635);
or UO_1402 (O_1402,N_29804,N_29977);
xnor UO_1403 (O_1403,N_29542,N_29746);
nand UO_1404 (O_1404,N_29602,N_29744);
nor UO_1405 (O_1405,N_29957,N_29839);
and UO_1406 (O_1406,N_29788,N_29806);
xnor UO_1407 (O_1407,N_29564,N_29888);
or UO_1408 (O_1408,N_29862,N_29798);
and UO_1409 (O_1409,N_29661,N_29626);
xor UO_1410 (O_1410,N_29532,N_29910);
and UO_1411 (O_1411,N_29830,N_29965);
xor UO_1412 (O_1412,N_29940,N_29843);
xnor UO_1413 (O_1413,N_29886,N_29605);
or UO_1414 (O_1414,N_29953,N_29603);
nor UO_1415 (O_1415,N_29883,N_29943);
or UO_1416 (O_1416,N_29946,N_29535);
and UO_1417 (O_1417,N_29579,N_29856);
or UO_1418 (O_1418,N_29906,N_29909);
and UO_1419 (O_1419,N_29890,N_29964);
and UO_1420 (O_1420,N_29737,N_29923);
or UO_1421 (O_1421,N_29534,N_29696);
and UO_1422 (O_1422,N_29752,N_29710);
xnor UO_1423 (O_1423,N_29947,N_29938);
xnor UO_1424 (O_1424,N_29555,N_29970);
xnor UO_1425 (O_1425,N_29934,N_29614);
xor UO_1426 (O_1426,N_29589,N_29572);
xnor UO_1427 (O_1427,N_29510,N_29573);
nor UO_1428 (O_1428,N_29946,N_29717);
nand UO_1429 (O_1429,N_29742,N_29644);
nor UO_1430 (O_1430,N_29815,N_29592);
and UO_1431 (O_1431,N_29771,N_29888);
nand UO_1432 (O_1432,N_29502,N_29735);
and UO_1433 (O_1433,N_29722,N_29732);
or UO_1434 (O_1434,N_29717,N_29959);
nand UO_1435 (O_1435,N_29835,N_29575);
nand UO_1436 (O_1436,N_29569,N_29560);
or UO_1437 (O_1437,N_29694,N_29633);
nand UO_1438 (O_1438,N_29930,N_29547);
and UO_1439 (O_1439,N_29952,N_29626);
or UO_1440 (O_1440,N_29760,N_29752);
and UO_1441 (O_1441,N_29668,N_29725);
nand UO_1442 (O_1442,N_29945,N_29660);
and UO_1443 (O_1443,N_29620,N_29893);
nor UO_1444 (O_1444,N_29551,N_29825);
xnor UO_1445 (O_1445,N_29974,N_29714);
nor UO_1446 (O_1446,N_29837,N_29678);
and UO_1447 (O_1447,N_29566,N_29520);
and UO_1448 (O_1448,N_29901,N_29949);
xor UO_1449 (O_1449,N_29798,N_29615);
xor UO_1450 (O_1450,N_29623,N_29739);
nor UO_1451 (O_1451,N_29617,N_29872);
nand UO_1452 (O_1452,N_29620,N_29866);
xnor UO_1453 (O_1453,N_29964,N_29637);
nand UO_1454 (O_1454,N_29887,N_29964);
xor UO_1455 (O_1455,N_29813,N_29991);
nand UO_1456 (O_1456,N_29899,N_29522);
and UO_1457 (O_1457,N_29557,N_29621);
nor UO_1458 (O_1458,N_29665,N_29880);
nor UO_1459 (O_1459,N_29696,N_29728);
xor UO_1460 (O_1460,N_29614,N_29954);
nand UO_1461 (O_1461,N_29656,N_29505);
xor UO_1462 (O_1462,N_29700,N_29989);
nand UO_1463 (O_1463,N_29731,N_29521);
xnor UO_1464 (O_1464,N_29782,N_29970);
and UO_1465 (O_1465,N_29542,N_29559);
nand UO_1466 (O_1466,N_29997,N_29596);
nor UO_1467 (O_1467,N_29928,N_29858);
and UO_1468 (O_1468,N_29946,N_29773);
xnor UO_1469 (O_1469,N_29859,N_29680);
nor UO_1470 (O_1470,N_29724,N_29937);
nor UO_1471 (O_1471,N_29535,N_29875);
and UO_1472 (O_1472,N_29719,N_29739);
xor UO_1473 (O_1473,N_29954,N_29982);
nor UO_1474 (O_1474,N_29513,N_29994);
and UO_1475 (O_1475,N_29537,N_29795);
and UO_1476 (O_1476,N_29882,N_29848);
and UO_1477 (O_1477,N_29704,N_29686);
nand UO_1478 (O_1478,N_29713,N_29572);
xnor UO_1479 (O_1479,N_29993,N_29643);
and UO_1480 (O_1480,N_29908,N_29517);
xor UO_1481 (O_1481,N_29529,N_29632);
and UO_1482 (O_1482,N_29856,N_29985);
xnor UO_1483 (O_1483,N_29634,N_29942);
xor UO_1484 (O_1484,N_29774,N_29952);
nand UO_1485 (O_1485,N_29960,N_29529);
and UO_1486 (O_1486,N_29681,N_29574);
nor UO_1487 (O_1487,N_29679,N_29610);
or UO_1488 (O_1488,N_29876,N_29843);
and UO_1489 (O_1489,N_29784,N_29515);
or UO_1490 (O_1490,N_29546,N_29796);
and UO_1491 (O_1491,N_29626,N_29933);
or UO_1492 (O_1492,N_29903,N_29518);
and UO_1493 (O_1493,N_29594,N_29642);
and UO_1494 (O_1494,N_29505,N_29753);
and UO_1495 (O_1495,N_29867,N_29967);
nand UO_1496 (O_1496,N_29930,N_29538);
xnor UO_1497 (O_1497,N_29702,N_29723);
nand UO_1498 (O_1498,N_29773,N_29629);
and UO_1499 (O_1499,N_29656,N_29720);
and UO_1500 (O_1500,N_29724,N_29986);
and UO_1501 (O_1501,N_29830,N_29853);
nor UO_1502 (O_1502,N_29734,N_29685);
and UO_1503 (O_1503,N_29891,N_29721);
nor UO_1504 (O_1504,N_29948,N_29799);
nand UO_1505 (O_1505,N_29526,N_29868);
or UO_1506 (O_1506,N_29559,N_29612);
xor UO_1507 (O_1507,N_29535,N_29814);
or UO_1508 (O_1508,N_29578,N_29572);
xnor UO_1509 (O_1509,N_29620,N_29737);
and UO_1510 (O_1510,N_29782,N_29506);
or UO_1511 (O_1511,N_29734,N_29660);
nor UO_1512 (O_1512,N_29848,N_29812);
and UO_1513 (O_1513,N_29904,N_29835);
and UO_1514 (O_1514,N_29700,N_29929);
or UO_1515 (O_1515,N_29767,N_29739);
nand UO_1516 (O_1516,N_29850,N_29982);
or UO_1517 (O_1517,N_29685,N_29503);
nand UO_1518 (O_1518,N_29705,N_29590);
and UO_1519 (O_1519,N_29977,N_29671);
nand UO_1520 (O_1520,N_29607,N_29530);
or UO_1521 (O_1521,N_29714,N_29808);
nor UO_1522 (O_1522,N_29512,N_29946);
or UO_1523 (O_1523,N_29927,N_29667);
and UO_1524 (O_1524,N_29728,N_29817);
nand UO_1525 (O_1525,N_29645,N_29960);
and UO_1526 (O_1526,N_29598,N_29908);
and UO_1527 (O_1527,N_29577,N_29603);
or UO_1528 (O_1528,N_29580,N_29542);
xor UO_1529 (O_1529,N_29662,N_29725);
nor UO_1530 (O_1530,N_29703,N_29958);
and UO_1531 (O_1531,N_29584,N_29961);
or UO_1532 (O_1532,N_29593,N_29539);
or UO_1533 (O_1533,N_29858,N_29777);
xnor UO_1534 (O_1534,N_29581,N_29930);
or UO_1535 (O_1535,N_29521,N_29582);
xnor UO_1536 (O_1536,N_29570,N_29744);
xor UO_1537 (O_1537,N_29558,N_29593);
nand UO_1538 (O_1538,N_29513,N_29588);
and UO_1539 (O_1539,N_29573,N_29704);
nor UO_1540 (O_1540,N_29792,N_29954);
nor UO_1541 (O_1541,N_29852,N_29892);
xnor UO_1542 (O_1542,N_29708,N_29904);
nand UO_1543 (O_1543,N_29593,N_29952);
xnor UO_1544 (O_1544,N_29598,N_29703);
xor UO_1545 (O_1545,N_29729,N_29664);
nand UO_1546 (O_1546,N_29515,N_29520);
nand UO_1547 (O_1547,N_29517,N_29700);
nand UO_1548 (O_1548,N_29507,N_29902);
nand UO_1549 (O_1549,N_29516,N_29546);
or UO_1550 (O_1550,N_29793,N_29916);
nand UO_1551 (O_1551,N_29846,N_29944);
nand UO_1552 (O_1552,N_29982,N_29711);
nand UO_1553 (O_1553,N_29825,N_29956);
and UO_1554 (O_1554,N_29613,N_29645);
xor UO_1555 (O_1555,N_29678,N_29557);
nor UO_1556 (O_1556,N_29516,N_29941);
nor UO_1557 (O_1557,N_29751,N_29659);
xnor UO_1558 (O_1558,N_29932,N_29577);
or UO_1559 (O_1559,N_29917,N_29817);
xor UO_1560 (O_1560,N_29915,N_29788);
nor UO_1561 (O_1561,N_29663,N_29743);
nand UO_1562 (O_1562,N_29777,N_29846);
nor UO_1563 (O_1563,N_29573,N_29508);
or UO_1564 (O_1564,N_29733,N_29814);
or UO_1565 (O_1565,N_29951,N_29745);
or UO_1566 (O_1566,N_29907,N_29733);
or UO_1567 (O_1567,N_29952,N_29633);
or UO_1568 (O_1568,N_29549,N_29973);
xor UO_1569 (O_1569,N_29702,N_29989);
xor UO_1570 (O_1570,N_29861,N_29844);
nor UO_1571 (O_1571,N_29513,N_29734);
and UO_1572 (O_1572,N_29875,N_29506);
xnor UO_1573 (O_1573,N_29517,N_29952);
or UO_1574 (O_1574,N_29817,N_29522);
nor UO_1575 (O_1575,N_29903,N_29947);
xor UO_1576 (O_1576,N_29950,N_29855);
or UO_1577 (O_1577,N_29983,N_29684);
xnor UO_1578 (O_1578,N_29551,N_29982);
nor UO_1579 (O_1579,N_29726,N_29556);
nand UO_1580 (O_1580,N_29553,N_29527);
xnor UO_1581 (O_1581,N_29977,N_29822);
xor UO_1582 (O_1582,N_29825,N_29916);
xor UO_1583 (O_1583,N_29933,N_29817);
nand UO_1584 (O_1584,N_29939,N_29560);
and UO_1585 (O_1585,N_29788,N_29909);
and UO_1586 (O_1586,N_29721,N_29707);
or UO_1587 (O_1587,N_29718,N_29704);
or UO_1588 (O_1588,N_29721,N_29688);
xor UO_1589 (O_1589,N_29841,N_29732);
xnor UO_1590 (O_1590,N_29936,N_29979);
nor UO_1591 (O_1591,N_29709,N_29623);
nor UO_1592 (O_1592,N_29543,N_29984);
nor UO_1593 (O_1593,N_29919,N_29848);
nand UO_1594 (O_1594,N_29871,N_29991);
or UO_1595 (O_1595,N_29601,N_29566);
xor UO_1596 (O_1596,N_29940,N_29744);
xnor UO_1597 (O_1597,N_29948,N_29822);
nand UO_1598 (O_1598,N_29674,N_29977);
or UO_1599 (O_1599,N_29678,N_29733);
or UO_1600 (O_1600,N_29824,N_29905);
or UO_1601 (O_1601,N_29588,N_29550);
xor UO_1602 (O_1602,N_29867,N_29600);
or UO_1603 (O_1603,N_29527,N_29773);
xnor UO_1604 (O_1604,N_29679,N_29656);
or UO_1605 (O_1605,N_29914,N_29659);
or UO_1606 (O_1606,N_29695,N_29857);
or UO_1607 (O_1607,N_29665,N_29991);
nand UO_1608 (O_1608,N_29680,N_29975);
or UO_1609 (O_1609,N_29851,N_29829);
or UO_1610 (O_1610,N_29885,N_29751);
nand UO_1611 (O_1611,N_29867,N_29768);
or UO_1612 (O_1612,N_29836,N_29880);
nand UO_1613 (O_1613,N_29800,N_29761);
nor UO_1614 (O_1614,N_29680,N_29617);
nand UO_1615 (O_1615,N_29590,N_29657);
xor UO_1616 (O_1616,N_29959,N_29697);
or UO_1617 (O_1617,N_29768,N_29915);
nor UO_1618 (O_1618,N_29510,N_29849);
xnor UO_1619 (O_1619,N_29969,N_29624);
nand UO_1620 (O_1620,N_29572,N_29996);
and UO_1621 (O_1621,N_29816,N_29766);
nand UO_1622 (O_1622,N_29849,N_29691);
or UO_1623 (O_1623,N_29727,N_29763);
and UO_1624 (O_1624,N_29760,N_29779);
nand UO_1625 (O_1625,N_29832,N_29559);
xnor UO_1626 (O_1626,N_29846,N_29590);
nand UO_1627 (O_1627,N_29787,N_29837);
nor UO_1628 (O_1628,N_29958,N_29821);
nand UO_1629 (O_1629,N_29937,N_29942);
xnor UO_1630 (O_1630,N_29801,N_29595);
xor UO_1631 (O_1631,N_29542,N_29734);
and UO_1632 (O_1632,N_29838,N_29959);
nor UO_1633 (O_1633,N_29980,N_29679);
and UO_1634 (O_1634,N_29762,N_29666);
nor UO_1635 (O_1635,N_29973,N_29768);
xnor UO_1636 (O_1636,N_29637,N_29537);
or UO_1637 (O_1637,N_29690,N_29658);
or UO_1638 (O_1638,N_29852,N_29676);
and UO_1639 (O_1639,N_29912,N_29580);
or UO_1640 (O_1640,N_29570,N_29860);
or UO_1641 (O_1641,N_29597,N_29645);
nor UO_1642 (O_1642,N_29966,N_29699);
nand UO_1643 (O_1643,N_29784,N_29634);
nand UO_1644 (O_1644,N_29701,N_29580);
nor UO_1645 (O_1645,N_29586,N_29728);
nor UO_1646 (O_1646,N_29578,N_29716);
nand UO_1647 (O_1647,N_29518,N_29587);
nor UO_1648 (O_1648,N_29675,N_29711);
or UO_1649 (O_1649,N_29920,N_29549);
and UO_1650 (O_1650,N_29782,N_29815);
xor UO_1651 (O_1651,N_29532,N_29843);
nor UO_1652 (O_1652,N_29673,N_29599);
nor UO_1653 (O_1653,N_29927,N_29951);
or UO_1654 (O_1654,N_29903,N_29614);
nor UO_1655 (O_1655,N_29742,N_29549);
nand UO_1656 (O_1656,N_29939,N_29909);
and UO_1657 (O_1657,N_29560,N_29862);
and UO_1658 (O_1658,N_29740,N_29780);
and UO_1659 (O_1659,N_29883,N_29749);
nand UO_1660 (O_1660,N_29943,N_29572);
or UO_1661 (O_1661,N_29835,N_29783);
or UO_1662 (O_1662,N_29879,N_29575);
nand UO_1663 (O_1663,N_29986,N_29674);
nand UO_1664 (O_1664,N_29766,N_29719);
nand UO_1665 (O_1665,N_29932,N_29689);
or UO_1666 (O_1666,N_29586,N_29962);
or UO_1667 (O_1667,N_29706,N_29954);
and UO_1668 (O_1668,N_29719,N_29567);
or UO_1669 (O_1669,N_29534,N_29766);
and UO_1670 (O_1670,N_29937,N_29722);
nand UO_1671 (O_1671,N_29630,N_29595);
and UO_1672 (O_1672,N_29880,N_29658);
nand UO_1673 (O_1673,N_29977,N_29610);
xnor UO_1674 (O_1674,N_29800,N_29719);
and UO_1675 (O_1675,N_29904,N_29571);
and UO_1676 (O_1676,N_29881,N_29505);
xnor UO_1677 (O_1677,N_29556,N_29632);
xnor UO_1678 (O_1678,N_29899,N_29556);
and UO_1679 (O_1679,N_29829,N_29943);
and UO_1680 (O_1680,N_29871,N_29771);
or UO_1681 (O_1681,N_29578,N_29725);
nand UO_1682 (O_1682,N_29656,N_29798);
xnor UO_1683 (O_1683,N_29902,N_29558);
and UO_1684 (O_1684,N_29562,N_29973);
and UO_1685 (O_1685,N_29968,N_29791);
and UO_1686 (O_1686,N_29547,N_29939);
nor UO_1687 (O_1687,N_29664,N_29936);
nand UO_1688 (O_1688,N_29624,N_29536);
or UO_1689 (O_1689,N_29817,N_29747);
xor UO_1690 (O_1690,N_29954,N_29726);
and UO_1691 (O_1691,N_29593,N_29574);
xor UO_1692 (O_1692,N_29588,N_29539);
nand UO_1693 (O_1693,N_29825,N_29659);
or UO_1694 (O_1694,N_29802,N_29883);
nand UO_1695 (O_1695,N_29722,N_29516);
or UO_1696 (O_1696,N_29648,N_29911);
and UO_1697 (O_1697,N_29910,N_29935);
or UO_1698 (O_1698,N_29590,N_29813);
nor UO_1699 (O_1699,N_29926,N_29885);
nand UO_1700 (O_1700,N_29519,N_29763);
xnor UO_1701 (O_1701,N_29593,N_29588);
nor UO_1702 (O_1702,N_29796,N_29895);
nand UO_1703 (O_1703,N_29522,N_29872);
nand UO_1704 (O_1704,N_29959,N_29905);
or UO_1705 (O_1705,N_29825,N_29750);
or UO_1706 (O_1706,N_29792,N_29633);
nor UO_1707 (O_1707,N_29719,N_29536);
or UO_1708 (O_1708,N_29637,N_29738);
nand UO_1709 (O_1709,N_29850,N_29724);
and UO_1710 (O_1710,N_29736,N_29521);
nand UO_1711 (O_1711,N_29797,N_29990);
or UO_1712 (O_1712,N_29644,N_29829);
or UO_1713 (O_1713,N_29748,N_29528);
and UO_1714 (O_1714,N_29925,N_29697);
and UO_1715 (O_1715,N_29749,N_29559);
or UO_1716 (O_1716,N_29846,N_29633);
and UO_1717 (O_1717,N_29896,N_29580);
or UO_1718 (O_1718,N_29828,N_29940);
and UO_1719 (O_1719,N_29981,N_29811);
xnor UO_1720 (O_1720,N_29954,N_29688);
xnor UO_1721 (O_1721,N_29536,N_29523);
nand UO_1722 (O_1722,N_29735,N_29603);
xor UO_1723 (O_1723,N_29690,N_29594);
nor UO_1724 (O_1724,N_29822,N_29758);
xor UO_1725 (O_1725,N_29692,N_29734);
xnor UO_1726 (O_1726,N_29704,N_29822);
nor UO_1727 (O_1727,N_29968,N_29804);
nor UO_1728 (O_1728,N_29624,N_29668);
and UO_1729 (O_1729,N_29733,N_29547);
and UO_1730 (O_1730,N_29917,N_29557);
or UO_1731 (O_1731,N_29691,N_29889);
nand UO_1732 (O_1732,N_29741,N_29923);
nor UO_1733 (O_1733,N_29772,N_29841);
or UO_1734 (O_1734,N_29874,N_29907);
and UO_1735 (O_1735,N_29661,N_29859);
nand UO_1736 (O_1736,N_29755,N_29930);
nand UO_1737 (O_1737,N_29761,N_29959);
or UO_1738 (O_1738,N_29913,N_29609);
and UO_1739 (O_1739,N_29976,N_29917);
xnor UO_1740 (O_1740,N_29548,N_29578);
or UO_1741 (O_1741,N_29860,N_29556);
xnor UO_1742 (O_1742,N_29929,N_29608);
and UO_1743 (O_1743,N_29754,N_29598);
nand UO_1744 (O_1744,N_29828,N_29722);
and UO_1745 (O_1745,N_29605,N_29738);
xnor UO_1746 (O_1746,N_29773,N_29986);
nand UO_1747 (O_1747,N_29871,N_29680);
xor UO_1748 (O_1748,N_29653,N_29897);
xor UO_1749 (O_1749,N_29569,N_29512);
nand UO_1750 (O_1750,N_29845,N_29798);
nor UO_1751 (O_1751,N_29941,N_29714);
and UO_1752 (O_1752,N_29816,N_29828);
nand UO_1753 (O_1753,N_29816,N_29936);
nor UO_1754 (O_1754,N_29949,N_29579);
or UO_1755 (O_1755,N_29691,N_29995);
nor UO_1756 (O_1756,N_29584,N_29819);
or UO_1757 (O_1757,N_29894,N_29571);
and UO_1758 (O_1758,N_29998,N_29838);
nor UO_1759 (O_1759,N_29909,N_29827);
nor UO_1760 (O_1760,N_29550,N_29976);
and UO_1761 (O_1761,N_29968,N_29673);
or UO_1762 (O_1762,N_29688,N_29878);
nand UO_1763 (O_1763,N_29793,N_29590);
or UO_1764 (O_1764,N_29845,N_29662);
nor UO_1765 (O_1765,N_29771,N_29543);
and UO_1766 (O_1766,N_29992,N_29640);
and UO_1767 (O_1767,N_29898,N_29521);
xor UO_1768 (O_1768,N_29572,N_29696);
xor UO_1769 (O_1769,N_29930,N_29818);
xnor UO_1770 (O_1770,N_29998,N_29688);
nor UO_1771 (O_1771,N_29766,N_29822);
nor UO_1772 (O_1772,N_29626,N_29683);
xor UO_1773 (O_1773,N_29917,N_29689);
and UO_1774 (O_1774,N_29808,N_29918);
nand UO_1775 (O_1775,N_29656,N_29764);
or UO_1776 (O_1776,N_29765,N_29720);
and UO_1777 (O_1777,N_29962,N_29995);
nand UO_1778 (O_1778,N_29750,N_29615);
xor UO_1779 (O_1779,N_29697,N_29524);
xor UO_1780 (O_1780,N_29651,N_29819);
xnor UO_1781 (O_1781,N_29560,N_29678);
or UO_1782 (O_1782,N_29788,N_29812);
xor UO_1783 (O_1783,N_29518,N_29742);
xor UO_1784 (O_1784,N_29733,N_29538);
or UO_1785 (O_1785,N_29664,N_29921);
nor UO_1786 (O_1786,N_29631,N_29700);
xnor UO_1787 (O_1787,N_29907,N_29651);
and UO_1788 (O_1788,N_29534,N_29762);
nand UO_1789 (O_1789,N_29622,N_29935);
nand UO_1790 (O_1790,N_29818,N_29911);
and UO_1791 (O_1791,N_29885,N_29955);
nand UO_1792 (O_1792,N_29640,N_29644);
nor UO_1793 (O_1793,N_29801,N_29750);
xor UO_1794 (O_1794,N_29808,N_29769);
and UO_1795 (O_1795,N_29844,N_29790);
and UO_1796 (O_1796,N_29603,N_29945);
or UO_1797 (O_1797,N_29850,N_29908);
xnor UO_1798 (O_1798,N_29541,N_29824);
or UO_1799 (O_1799,N_29774,N_29544);
or UO_1800 (O_1800,N_29693,N_29521);
and UO_1801 (O_1801,N_29631,N_29587);
xnor UO_1802 (O_1802,N_29747,N_29873);
xor UO_1803 (O_1803,N_29592,N_29653);
nor UO_1804 (O_1804,N_29545,N_29618);
nand UO_1805 (O_1805,N_29894,N_29632);
xnor UO_1806 (O_1806,N_29625,N_29830);
nor UO_1807 (O_1807,N_29516,N_29837);
nand UO_1808 (O_1808,N_29888,N_29520);
xor UO_1809 (O_1809,N_29610,N_29886);
nor UO_1810 (O_1810,N_29781,N_29975);
xor UO_1811 (O_1811,N_29571,N_29577);
xor UO_1812 (O_1812,N_29763,N_29793);
xnor UO_1813 (O_1813,N_29796,N_29906);
or UO_1814 (O_1814,N_29751,N_29835);
nor UO_1815 (O_1815,N_29592,N_29851);
or UO_1816 (O_1816,N_29631,N_29670);
xor UO_1817 (O_1817,N_29792,N_29800);
nor UO_1818 (O_1818,N_29828,N_29916);
and UO_1819 (O_1819,N_29646,N_29957);
or UO_1820 (O_1820,N_29812,N_29557);
xor UO_1821 (O_1821,N_29731,N_29676);
nor UO_1822 (O_1822,N_29846,N_29629);
or UO_1823 (O_1823,N_29664,N_29825);
or UO_1824 (O_1824,N_29536,N_29637);
or UO_1825 (O_1825,N_29862,N_29863);
xor UO_1826 (O_1826,N_29611,N_29719);
nor UO_1827 (O_1827,N_29717,N_29884);
and UO_1828 (O_1828,N_29788,N_29960);
xor UO_1829 (O_1829,N_29560,N_29924);
nand UO_1830 (O_1830,N_29682,N_29739);
or UO_1831 (O_1831,N_29610,N_29718);
nor UO_1832 (O_1832,N_29999,N_29803);
nand UO_1833 (O_1833,N_29689,N_29834);
nand UO_1834 (O_1834,N_29834,N_29994);
nor UO_1835 (O_1835,N_29985,N_29822);
or UO_1836 (O_1836,N_29825,N_29939);
nand UO_1837 (O_1837,N_29568,N_29755);
nor UO_1838 (O_1838,N_29633,N_29779);
or UO_1839 (O_1839,N_29755,N_29920);
nor UO_1840 (O_1840,N_29849,N_29565);
and UO_1841 (O_1841,N_29517,N_29682);
nor UO_1842 (O_1842,N_29814,N_29656);
nor UO_1843 (O_1843,N_29984,N_29507);
and UO_1844 (O_1844,N_29980,N_29932);
and UO_1845 (O_1845,N_29761,N_29702);
xor UO_1846 (O_1846,N_29773,N_29940);
and UO_1847 (O_1847,N_29810,N_29872);
xor UO_1848 (O_1848,N_29631,N_29778);
xor UO_1849 (O_1849,N_29544,N_29826);
nand UO_1850 (O_1850,N_29757,N_29665);
nand UO_1851 (O_1851,N_29952,N_29885);
or UO_1852 (O_1852,N_29606,N_29544);
nor UO_1853 (O_1853,N_29627,N_29809);
nand UO_1854 (O_1854,N_29767,N_29885);
xnor UO_1855 (O_1855,N_29934,N_29947);
and UO_1856 (O_1856,N_29750,N_29755);
nor UO_1857 (O_1857,N_29744,N_29616);
or UO_1858 (O_1858,N_29563,N_29953);
xnor UO_1859 (O_1859,N_29838,N_29758);
or UO_1860 (O_1860,N_29530,N_29983);
nor UO_1861 (O_1861,N_29665,N_29556);
and UO_1862 (O_1862,N_29911,N_29801);
or UO_1863 (O_1863,N_29925,N_29945);
nor UO_1864 (O_1864,N_29769,N_29671);
or UO_1865 (O_1865,N_29830,N_29856);
xnor UO_1866 (O_1866,N_29707,N_29929);
nor UO_1867 (O_1867,N_29991,N_29937);
xor UO_1868 (O_1868,N_29991,N_29770);
nor UO_1869 (O_1869,N_29980,N_29619);
nor UO_1870 (O_1870,N_29698,N_29622);
and UO_1871 (O_1871,N_29578,N_29619);
or UO_1872 (O_1872,N_29679,N_29876);
xnor UO_1873 (O_1873,N_29939,N_29515);
nand UO_1874 (O_1874,N_29544,N_29881);
xnor UO_1875 (O_1875,N_29742,N_29962);
nor UO_1876 (O_1876,N_29576,N_29660);
or UO_1877 (O_1877,N_29798,N_29961);
xor UO_1878 (O_1878,N_29522,N_29537);
nand UO_1879 (O_1879,N_29741,N_29652);
and UO_1880 (O_1880,N_29563,N_29813);
xor UO_1881 (O_1881,N_29908,N_29758);
and UO_1882 (O_1882,N_29828,N_29572);
xnor UO_1883 (O_1883,N_29867,N_29524);
nor UO_1884 (O_1884,N_29662,N_29620);
nand UO_1885 (O_1885,N_29500,N_29674);
and UO_1886 (O_1886,N_29595,N_29691);
nor UO_1887 (O_1887,N_29998,N_29829);
xnor UO_1888 (O_1888,N_29783,N_29790);
or UO_1889 (O_1889,N_29829,N_29726);
nor UO_1890 (O_1890,N_29719,N_29873);
nand UO_1891 (O_1891,N_29669,N_29610);
or UO_1892 (O_1892,N_29633,N_29689);
xor UO_1893 (O_1893,N_29824,N_29618);
and UO_1894 (O_1894,N_29617,N_29739);
and UO_1895 (O_1895,N_29767,N_29680);
nand UO_1896 (O_1896,N_29917,N_29923);
xor UO_1897 (O_1897,N_29911,N_29637);
nor UO_1898 (O_1898,N_29555,N_29625);
and UO_1899 (O_1899,N_29744,N_29844);
and UO_1900 (O_1900,N_29915,N_29907);
nor UO_1901 (O_1901,N_29674,N_29823);
or UO_1902 (O_1902,N_29663,N_29939);
and UO_1903 (O_1903,N_29983,N_29916);
nor UO_1904 (O_1904,N_29818,N_29996);
nor UO_1905 (O_1905,N_29596,N_29699);
and UO_1906 (O_1906,N_29616,N_29905);
nor UO_1907 (O_1907,N_29918,N_29922);
and UO_1908 (O_1908,N_29773,N_29537);
or UO_1909 (O_1909,N_29986,N_29764);
or UO_1910 (O_1910,N_29542,N_29665);
and UO_1911 (O_1911,N_29692,N_29565);
nand UO_1912 (O_1912,N_29638,N_29804);
nor UO_1913 (O_1913,N_29818,N_29927);
or UO_1914 (O_1914,N_29957,N_29577);
nor UO_1915 (O_1915,N_29938,N_29555);
or UO_1916 (O_1916,N_29572,N_29782);
xor UO_1917 (O_1917,N_29811,N_29843);
nor UO_1918 (O_1918,N_29815,N_29774);
or UO_1919 (O_1919,N_29768,N_29605);
or UO_1920 (O_1920,N_29977,N_29931);
nor UO_1921 (O_1921,N_29989,N_29622);
nand UO_1922 (O_1922,N_29637,N_29570);
or UO_1923 (O_1923,N_29577,N_29566);
nor UO_1924 (O_1924,N_29785,N_29928);
nor UO_1925 (O_1925,N_29752,N_29707);
nand UO_1926 (O_1926,N_29640,N_29872);
nor UO_1927 (O_1927,N_29605,N_29835);
xnor UO_1928 (O_1928,N_29569,N_29952);
or UO_1929 (O_1929,N_29993,N_29989);
xor UO_1930 (O_1930,N_29968,N_29949);
and UO_1931 (O_1931,N_29936,N_29907);
and UO_1932 (O_1932,N_29682,N_29581);
nor UO_1933 (O_1933,N_29587,N_29726);
and UO_1934 (O_1934,N_29602,N_29664);
or UO_1935 (O_1935,N_29781,N_29957);
nor UO_1936 (O_1936,N_29564,N_29706);
nor UO_1937 (O_1937,N_29824,N_29973);
or UO_1938 (O_1938,N_29772,N_29684);
or UO_1939 (O_1939,N_29755,N_29722);
xor UO_1940 (O_1940,N_29594,N_29610);
xnor UO_1941 (O_1941,N_29945,N_29708);
nor UO_1942 (O_1942,N_29959,N_29878);
and UO_1943 (O_1943,N_29609,N_29702);
xnor UO_1944 (O_1944,N_29850,N_29898);
nand UO_1945 (O_1945,N_29794,N_29743);
nand UO_1946 (O_1946,N_29551,N_29915);
nand UO_1947 (O_1947,N_29574,N_29687);
nor UO_1948 (O_1948,N_29905,N_29876);
nand UO_1949 (O_1949,N_29889,N_29877);
nand UO_1950 (O_1950,N_29754,N_29942);
nand UO_1951 (O_1951,N_29999,N_29696);
nor UO_1952 (O_1952,N_29836,N_29540);
nand UO_1953 (O_1953,N_29506,N_29654);
xor UO_1954 (O_1954,N_29992,N_29780);
nand UO_1955 (O_1955,N_29952,N_29766);
xnor UO_1956 (O_1956,N_29536,N_29694);
nor UO_1957 (O_1957,N_29848,N_29830);
nand UO_1958 (O_1958,N_29787,N_29920);
xnor UO_1959 (O_1959,N_29856,N_29966);
or UO_1960 (O_1960,N_29748,N_29867);
and UO_1961 (O_1961,N_29506,N_29787);
nand UO_1962 (O_1962,N_29745,N_29667);
xnor UO_1963 (O_1963,N_29579,N_29615);
or UO_1964 (O_1964,N_29814,N_29545);
or UO_1965 (O_1965,N_29541,N_29578);
nand UO_1966 (O_1966,N_29601,N_29591);
nand UO_1967 (O_1967,N_29581,N_29519);
nand UO_1968 (O_1968,N_29781,N_29649);
xor UO_1969 (O_1969,N_29865,N_29878);
nand UO_1970 (O_1970,N_29754,N_29984);
nor UO_1971 (O_1971,N_29842,N_29759);
and UO_1972 (O_1972,N_29788,N_29827);
nand UO_1973 (O_1973,N_29995,N_29970);
or UO_1974 (O_1974,N_29984,N_29585);
nand UO_1975 (O_1975,N_29540,N_29784);
or UO_1976 (O_1976,N_29673,N_29790);
and UO_1977 (O_1977,N_29995,N_29830);
and UO_1978 (O_1978,N_29707,N_29993);
and UO_1979 (O_1979,N_29551,N_29751);
xnor UO_1980 (O_1980,N_29754,N_29715);
nand UO_1981 (O_1981,N_29957,N_29963);
and UO_1982 (O_1982,N_29745,N_29860);
xnor UO_1983 (O_1983,N_29859,N_29972);
and UO_1984 (O_1984,N_29744,N_29762);
nor UO_1985 (O_1985,N_29727,N_29625);
and UO_1986 (O_1986,N_29806,N_29565);
and UO_1987 (O_1987,N_29915,N_29728);
nand UO_1988 (O_1988,N_29516,N_29520);
nor UO_1989 (O_1989,N_29638,N_29741);
xor UO_1990 (O_1990,N_29588,N_29626);
or UO_1991 (O_1991,N_29588,N_29679);
xnor UO_1992 (O_1992,N_29646,N_29554);
nor UO_1993 (O_1993,N_29634,N_29795);
nand UO_1994 (O_1994,N_29762,N_29565);
nand UO_1995 (O_1995,N_29689,N_29985);
xor UO_1996 (O_1996,N_29696,N_29825);
and UO_1997 (O_1997,N_29987,N_29579);
and UO_1998 (O_1998,N_29600,N_29991);
or UO_1999 (O_1999,N_29770,N_29565);
nand UO_2000 (O_2000,N_29969,N_29513);
nor UO_2001 (O_2001,N_29862,N_29808);
nand UO_2002 (O_2002,N_29804,N_29986);
and UO_2003 (O_2003,N_29962,N_29735);
xor UO_2004 (O_2004,N_29534,N_29567);
xor UO_2005 (O_2005,N_29880,N_29840);
or UO_2006 (O_2006,N_29776,N_29822);
and UO_2007 (O_2007,N_29929,N_29512);
nand UO_2008 (O_2008,N_29671,N_29538);
and UO_2009 (O_2009,N_29663,N_29872);
nand UO_2010 (O_2010,N_29786,N_29914);
or UO_2011 (O_2011,N_29699,N_29676);
nand UO_2012 (O_2012,N_29731,N_29599);
nand UO_2013 (O_2013,N_29890,N_29768);
or UO_2014 (O_2014,N_29975,N_29568);
and UO_2015 (O_2015,N_29761,N_29597);
xor UO_2016 (O_2016,N_29788,N_29527);
nor UO_2017 (O_2017,N_29565,N_29515);
and UO_2018 (O_2018,N_29750,N_29884);
xnor UO_2019 (O_2019,N_29949,N_29622);
or UO_2020 (O_2020,N_29618,N_29777);
or UO_2021 (O_2021,N_29936,N_29958);
nand UO_2022 (O_2022,N_29715,N_29995);
and UO_2023 (O_2023,N_29578,N_29967);
xnor UO_2024 (O_2024,N_29599,N_29587);
nor UO_2025 (O_2025,N_29599,N_29714);
or UO_2026 (O_2026,N_29971,N_29532);
and UO_2027 (O_2027,N_29837,N_29641);
and UO_2028 (O_2028,N_29987,N_29604);
nor UO_2029 (O_2029,N_29791,N_29573);
nand UO_2030 (O_2030,N_29863,N_29825);
xor UO_2031 (O_2031,N_29871,N_29596);
or UO_2032 (O_2032,N_29786,N_29699);
xnor UO_2033 (O_2033,N_29507,N_29807);
nand UO_2034 (O_2034,N_29627,N_29700);
nor UO_2035 (O_2035,N_29598,N_29561);
and UO_2036 (O_2036,N_29755,N_29976);
nand UO_2037 (O_2037,N_29571,N_29537);
and UO_2038 (O_2038,N_29867,N_29516);
nor UO_2039 (O_2039,N_29608,N_29928);
nor UO_2040 (O_2040,N_29848,N_29659);
nor UO_2041 (O_2041,N_29932,N_29988);
nand UO_2042 (O_2042,N_29537,N_29665);
xor UO_2043 (O_2043,N_29507,N_29756);
xor UO_2044 (O_2044,N_29980,N_29582);
nand UO_2045 (O_2045,N_29930,N_29706);
nand UO_2046 (O_2046,N_29802,N_29645);
nor UO_2047 (O_2047,N_29596,N_29625);
xor UO_2048 (O_2048,N_29616,N_29841);
nor UO_2049 (O_2049,N_29799,N_29501);
and UO_2050 (O_2050,N_29777,N_29564);
or UO_2051 (O_2051,N_29723,N_29745);
or UO_2052 (O_2052,N_29836,N_29597);
nand UO_2053 (O_2053,N_29569,N_29784);
nor UO_2054 (O_2054,N_29650,N_29672);
nor UO_2055 (O_2055,N_29891,N_29643);
or UO_2056 (O_2056,N_29783,N_29676);
xor UO_2057 (O_2057,N_29924,N_29794);
or UO_2058 (O_2058,N_29549,N_29543);
xor UO_2059 (O_2059,N_29743,N_29563);
nand UO_2060 (O_2060,N_29834,N_29924);
nand UO_2061 (O_2061,N_29875,N_29610);
and UO_2062 (O_2062,N_29876,N_29936);
nor UO_2063 (O_2063,N_29690,N_29917);
xor UO_2064 (O_2064,N_29645,N_29874);
and UO_2065 (O_2065,N_29546,N_29627);
and UO_2066 (O_2066,N_29830,N_29665);
nor UO_2067 (O_2067,N_29990,N_29594);
or UO_2068 (O_2068,N_29512,N_29752);
or UO_2069 (O_2069,N_29765,N_29861);
nand UO_2070 (O_2070,N_29543,N_29838);
nor UO_2071 (O_2071,N_29837,N_29603);
xor UO_2072 (O_2072,N_29806,N_29906);
xnor UO_2073 (O_2073,N_29766,N_29999);
or UO_2074 (O_2074,N_29509,N_29998);
and UO_2075 (O_2075,N_29557,N_29874);
or UO_2076 (O_2076,N_29805,N_29738);
nand UO_2077 (O_2077,N_29638,N_29705);
nand UO_2078 (O_2078,N_29678,N_29823);
xnor UO_2079 (O_2079,N_29927,N_29849);
xnor UO_2080 (O_2080,N_29838,N_29644);
or UO_2081 (O_2081,N_29957,N_29541);
and UO_2082 (O_2082,N_29906,N_29863);
and UO_2083 (O_2083,N_29717,N_29753);
xor UO_2084 (O_2084,N_29708,N_29946);
or UO_2085 (O_2085,N_29651,N_29686);
xor UO_2086 (O_2086,N_29650,N_29610);
or UO_2087 (O_2087,N_29617,N_29976);
and UO_2088 (O_2088,N_29696,N_29654);
and UO_2089 (O_2089,N_29900,N_29959);
or UO_2090 (O_2090,N_29542,N_29852);
and UO_2091 (O_2091,N_29518,N_29756);
or UO_2092 (O_2092,N_29519,N_29731);
or UO_2093 (O_2093,N_29724,N_29658);
or UO_2094 (O_2094,N_29765,N_29707);
nand UO_2095 (O_2095,N_29852,N_29950);
nand UO_2096 (O_2096,N_29832,N_29724);
nand UO_2097 (O_2097,N_29978,N_29601);
or UO_2098 (O_2098,N_29716,N_29642);
nand UO_2099 (O_2099,N_29742,N_29624);
nand UO_2100 (O_2100,N_29639,N_29585);
nand UO_2101 (O_2101,N_29656,N_29689);
and UO_2102 (O_2102,N_29885,N_29528);
nand UO_2103 (O_2103,N_29905,N_29919);
nor UO_2104 (O_2104,N_29891,N_29920);
nor UO_2105 (O_2105,N_29582,N_29574);
nand UO_2106 (O_2106,N_29949,N_29747);
xor UO_2107 (O_2107,N_29510,N_29820);
nand UO_2108 (O_2108,N_29689,N_29814);
nand UO_2109 (O_2109,N_29872,N_29722);
xnor UO_2110 (O_2110,N_29922,N_29960);
and UO_2111 (O_2111,N_29990,N_29778);
and UO_2112 (O_2112,N_29698,N_29933);
and UO_2113 (O_2113,N_29570,N_29643);
nand UO_2114 (O_2114,N_29560,N_29802);
nand UO_2115 (O_2115,N_29942,N_29687);
xor UO_2116 (O_2116,N_29826,N_29602);
nor UO_2117 (O_2117,N_29975,N_29995);
or UO_2118 (O_2118,N_29789,N_29606);
nor UO_2119 (O_2119,N_29742,N_29833);
and UO_2120 (O_2120,N_29786,N_29835);
nand UO_2121 (O_2121,N_29976,N_29764);
nor UO_2122 (O_2122,N_29621,N_29517);
and UO_2123 (O_2123,N_29565,N_29603);
and UO_2124 (O_2124,N_29938,N_29963);
or UO_2125 (O_2125,N_29808,N_29965);
nand UO_2126 (O_2126,N_29581,N_29500);
and UO_2127 (O_2127,N_29887,N_29673);
nand UO_2128 (O_2128,N_29732,N_29866);
nor UO_2129 (O_2129,N_29593,N_29524);
nand UO_2130 (O_2130,N_29736,N_29752);
xor UO_2131 (O_2131,N_29910,N_29597);
or UO_2132 (O_2132,N_29605,N_29941);
or UO_2133 (O_2133,N_29780,N_29610);
xnor UO_2134 (O_2134,N_29795,N_29559);
nand UO_2135 (O_2135,N_29668,N_29719);
nor UO_2136 (O_2136,N_29755,N_29712);
and UO_2137 (O_2137,N_29628,N_29627);
and UO_2138 (O_2138,N_29610,N_29619);
nand UO_2139 (O_2139,N_29566,N_29611);
nor UO_2140 (O_2140,N_29985,N_29502);
nand UO_2141 (O_2141,N_29575,N_29640);
and UO_2142 (O_2142,N_29693,N_29529);
nor UO_2143 (O_2143,N_29883,N_29552);
or UO_2144 (O_2144,N_29813,N_29887);
nand UO_2145 (O_2145,N_29573,N_29820);
nor UO_2146 (O_2146,N_29673,N_29719);
or UO_2147 (O_2147,N_29676,N_29664);
nor UO_2148 (O_2148,N_29602,N_29912);
or UO_2149 (O_2149,N_29784,N_29579);
nor UO_2150 (O_2150,N_29887,N_29540);
xor UO_2151 (O_2151,N_29558,N_29516);
or UO_2152 (O_2152,N_29801,N_29632);
nor UO_2153 (O_2153,N_29797,N_29627);
xor UO_2154 (O_2154,N_29526,N_29635);
and UO_2155 (O_2155,N_29569,N_29998);
and UO_2156 (O_2156,N_29653,N_29840);
nor UO_2157 (O_2157,N_29750,N_29661);
xnor UO_2158 (O_2158,N_29534,N_29973);
nand UO_2159 (O_2159,N_29557,N_29676);
xnor UO_2160 (O_2160,N_29761,N_29914);
and UO_2161 (O_2161,N_29572,N_29591);
nand UO_2162 (O_2162,N_29580,N_29676);
nor UO_2163 (O_2163,N_29526,N_29626);
nand UO_2164 (O_2164,N_29631,N_29907);
or UO_2165 (O_2165,N_29565,N_29917);
and UO_2166 (O_2166,N_29850,N_29895);
nor UO_2167 (O_2167,N_29577,N_29706);
nand UO_2168 (O_2168,N_29962,N_29819);
xnor UO_2169 (O_2169,N_29518,N_29768);
nor UO_2170 (O_2170,N_29924,N_29597);
and UO_2171 (O_2171,N_29685,N_29744);
and UO_2172 (O_2172,N_29974,N_29513);
and UO_2173 (O_2173,N_29724,N_29779);
nor UO_2174 (O_2174,N_29772,N_29801);
nand UO_2175 (O_2175,N_29977,N_29687);
and UO_2176 (O_2176,N_29550,N_29511);
nor UO_2177 (O_2177,N_29536,N_29803);
or UO_2178 (O_2178,N_29860,N_29786);
xor UO_2179 (O_2179,N_29713,N_29831);
or UO_2180 (O_2180,N_29622,N_29933);
xor UO_2181 (O_2181,N_29747,N_29604);
nor UO_2182 (O_2182,N_29745,N_29595);
and UO_2183 (O_2183,N_29664,N_29970);
xnor UO_2184 (O_2184,N_29804,N_29562);
or UO_2185 (O_2185,N_29796,N_29995);
nor UO_2186 (O_2186,N_29552,N_29554);
and UO_2187 (O_2187,N_29544,N_29702);
and UO_2188 (O_2188,N_29884,N_29873);
or UO_2189 (O_2189,N_29520,N_29975);
xor UO_2190 (O_2190,N_29764,N_29866);
nor UO_2191 (O_2191,N_29888,N_29827);
or UO_2192 (O_2192,N_29603,N_29720);
nor UO_2193 (O_2193,N_29740,N_29772);
xor UO_2194 (O_2194,N_29622,N_29534);
and UO_2195 (O_2195,N_29631,N_29814);
nand UO_2196 (O_2196,N_29663,N_29576);
or UO_2197 (O_2197,N_29583,N_29969);
and UO_2198 (O_2198,N_29818,N_29540);
and UO_2199 (O_2199,N_29878,N_29646);
and UO_2200 (O_2200,N_29922,N_29505);
xor UO_2201 (O_2201,N_29692,N_29674);
nor UO_2202 (O_2202,N_29822,N_29910);
nand UO_2203 (O_2203,N_29779,N_29863);
or UO_2204 (O_2204,N_29501,N_29966);
nor UO_2205 (O_2205,N_29815,N_29779);
nor UO_2206 (O_2206,N_29519,N_29573);
or UO_2207 (O_2207,N_29707,N_29657);
xor UO_2208 (O_2208,N_29766,N_29916);
and UO_2209 (O_2209,N_29521,N_29821);
nand UO_2210 (O_2210,N_29617,N_29800);
or UO_2211 (O_2211,N_29544,N_29725);
or UO_2212 (O_2212,N_29813,N_29694);
or UO_2213 (O_2213,N_29955,N_29869);
nand UO_2214 (O_2214,N_29622,N_29588);
or UO_2215 (O_2215,N_29756,N_29546);
xnor UO_2216 (O_2216,N_29900,N_29986);
nor UO_2217 (O_2217,N_29513,N_29628);
nor UO_2218 (O_2218,N_29891,N_29712);
and UO_2219 (O_2219,N_29544,N_29971);
nand UO_2220 (O_2220,N_29944,N_29797);
xor UO_2221 (O_2221,N_29831,N_29635);
nand UO_2222 (O_2222,N_29767,N_29802);
xnor UO_2223 (O_2223,N_29811,N_29588);
or UO_2224 (O_2224,N_29648,N_29932);
xnor UO_2225 (O_2225,N_29986,N_29746);
nor UO_2226 (O_2226,N_29769,N_29886);
or UO_2227 (O_2227,N_29956,N_29732);
and UO_2228 (O_2228,N_29899,N_29547);
nor UO_2229 (O_2229,N_29777,N_29606);
nand UO_2230 (O_2230,N_29794,N_29611);
and UO_2231 (O_2231,N_29814,N_29711);
nor UO_2232 (O_2232,N_29517,N_29848);
nor UO_2233 (O_2233,N_29876,N_29802);
and UO_2234 (O_2234,N_29985,N_29958);
nand UO_2235 (O_2235,N_29650,N_29645);
and UO_2236 (O_2236,N_29911,N_29842);
xor UO_2237 (O_2237,N_29691,N_29925);
and UO_2238 (O_2238,N_29853,N_29769);
xor UO_2239 (O_2239,N_29852,N_29746);
or UO_2240 (O_2240,N_29976,N_29537);
nor UO_2241 (O_2241,N_29510,N_29724);
and UO_2242 (O_2242,N_29661,N_29918);
nand UO_2243 (O_2243,N_29618,N_29854);
nor UO_2244 (O_2244,N_29721,N_29598);
xnor UO_2245 (O_2245,N_29586,N_29923);
or UO_2246 (O_2246,N_29936,N_29530);
and UO_2247 (O_2247,N_29518,N_29773);
xor UO_2248 (O_2248,N_29887,N_29921);
xor UO_2249 (O_2249,N_29580,N_29501);
nor UO_2250 (O_2250,N_29846,N_29886);
nor UO_2251 (O_2251,N_29575,N_29667);
nor UO_2252 (O_2252,N_29653,N_29724);
and UO_2253 (O_2253,N_29772,N_29829);
or UO_2254 (O_2254,N_29783,N_29671);
nand UO_2255 (O_2255,N_29791,N_29963);
xnor UO_2256 (O_2256,N_29634,N_29753);
nand UO_2257 (O_2257,N_29562,N_29717);
or UO_2258 (O_2258,N_29675,N_29906);
nand UO_2259 (O_2259,N_29790,N_29682);
or UO_2260 (O_2260,N_29797,N_29805);
xor UO_2261 (O_2261,N_29523,N_29673);
nand UO_2262 (O_2262,N_29886,N_29655);
or UO_2263 (O_2263,N_29893,N_29988);
and UO_2264 (O_2264,N_29958,N_29779);
or UO_2265 (O_2265,N_29928,N_29914);
nor UO_2266 (O_2266,N_29707,N_29548);
nor UO_2267 (O_2267,N_29871,N_29743);
nor UO_2268 (O_2268,N_29555,N_29754);
and UO_2269 (O_2269,N_29873,N_29685);
nand UO_2270 (O_2270,N_29510,N_29894);
xnor UO_2271 (O_2271,N_29657,N_29702);
xnor UO_2272 (O_2272,N_29556,N_29918);
xnor UO_2273 (O_2273,N_29962,N_29558);
xor UO_2274 (O_2274,N_29636,N_29715);
xor UO_2275 (O_2275,N_29699,N_29910);
and UO_2276 (O_2276,N_29544,N_29569);
nand UO_2277 (O_2277,N_29853,N_29764);
xnor UO_2278 (O_2278,N_29712,N_29549);
nor UO_2279 (O_2279,N_29948,N_29787);
nor UO_2280 (O_2280,N_29846,N_29587);
xnor UO_2281 (O_2281,N_29655,N_29583);
and UO_2282 (O_2282,N_29779,N_29585);
or UO_2283 (O_2283,N_29625,N_29658);
nand UO_2284 (O_2284,N_29947,N_29822);
xnor UO_2285 (O_2285,N_29575,N_29669);
xnor UO_2286 (O_2286,N_29671,N_29504);
and UO_2287 (O_2287,N_29710,N_29741);
or UO_2288 (O_2288,N_29600,N_29610);
xnor UO_2289 (O_2289,N_29617,N_29865);
or UO_2290 (O_2290,N_29635,N_29685);
nand UO_2291 (O_2291,N_29876,N_29734);
nor UO_2292 (O_2292,N_29613,N_29803);
and UO_2293 (O_2293,N_29626,N_29925);
and UO_2294 (O_2294,N_29606,N_29646);
xor UO_2295 (O_2295,N_29610,N_29915);
xor UO_2296 (O_2296,N_29590,N_29966);
nor UO_2297 (O_2297,N_29546,N_29748);
or UO_2298 (O_2298,N_29825,N_29699);
and UO_2299 (O_2299,N_29556,N_29511);
xor UO_2300 (O_2300,N_29907,N_29914);
or UO_2301 (O_2301,N_29508,N_29826);
or UO_2302 (O_2302,N_29808,N_29904);
or UO_2303 (O_2303,N_29802,N_29974);
nor UO_2304 (O_2304,N_29771,N_29911);
or UO_2305 (O_2305,N_29998,N_29544);
nor UO_2306 (O_2306,N_29754,N_29668);
and UO_2307 (O_2307,N_29585,N_29647);
nand UO_2308 (O_2308,N_29888,N_29606);
nor UO_2309 (O_2309,N_29739,N_29877);
nor UO_2310 (O_2310,N_29692,N_29680);
nand UO_2311 (O_2311,N_29910,N_29647);
xnor UO_2312 (O_2312,N_29938,N_29769);
or UO_2313 (O_2313,N_29659,N_29924);
xor UO_2314 (O_2314,N_29631,N_29767);
and UO_2315 (O_2315,N_29744,N_29638);
nor UO_2316 (O_2316,N_29583,N_29756);
xor UO_2317 (O_2317,N_29546,N_29977);
nand UO_2318 (O_2318,N_29931,N_29901);
or UO_2319 (O_2319,N_29680,N_29534);
and UO_2320 (O_2320,N_29696,N_29502);
or UO_2321 (O_2321,N_29979,N_29975);
and UO_2322 (O_2322,N_29602,N_29768);
and UO_2323 (O_2323,N_29642,N_29751);
and UO_2324 (O_2324,N_29964,N_29621);
and UO_2325 (O_2325,N_29894,N_29682);
nor UO_2326 (O_2326,N_29772,N_29803);
nand UO_2327 (O_2327,N_29606,N_29717);
and UO_2328 (O_2328,N_29857,N_29947);
or UO_2329 (O_2329,N_29862,N_29664);
xor UO_2330 (O_2330,N_29571,N_29708);
xnor UO_2331 (O_2331,N_29664,N_29960);
xnor UO_2332 (O_2332,N_29670,N_29558);
nor UO_2333 (O_2333,N_29625,N_29824);
nand UO_2334 (O_2334,N_29747,N_29532);
and UO_2335 (O_2335,N_29937,N_29560);
nand UO_2336 (O_2336,N_29755,N_29611);
or UO_2337 (O_2337,N_29776,N_29829);
nor UO_2338 (O_2338,N_29702,N_29668);
nor UO_2339 (O_2339,N_29913,N_29668);
nor UO_2340 (O_2340,N_29834,N_29621);
xnor UO_2341 (O_2341,N_29848,N_29836);
or UO_2342 (O_2342,N_29680,N_29832);
or UO_2343 (O_2343,N_29769,N_29827);
xnor UO_2344 (O_2344,N_29682,N_29699);
xnor UO_2345 (O_2345,N_29770,N_29587);
nand UO_2346 (O_2346,N_29713,N_29984);
or UO_2347 (O_2347,N_29811,N_29962);
xor UO_2348 (O_2348,N_29607,N_29900);
or UO_2349 (O_2349,N_29760,N_29786);
and UO_2350 (O_2350,N_29716,N_29825);
xnor UO_2351 (O_2351,N_29715,N_29529);
or UO_2352 (O_2352,N_29930,N_29952);
and UO_2353 (O_2353,N_29637,N_29944);
xnor UO_2354 (O_2354,N_29566,N_29846);
or UO_2355 (O_2355,N_29758,N_29864);
xor UO_2356 (O_2356,N_29537,N_29966);
or UO_2357 (O_2357,N_29643,N_29877);
nand UO_2358 (O_2358,N_29574,N_29664);
nor UO_2359 (O_2359,N_29617,N_29573);
nand UO_2360 (O_2360,N_29785,N_29943);
nand UO_2361 (O_2361,N_29550,N_29908);
nand UO_2362 (O_2362,N_29656,N_29855);
and UO_2363 (O_2363,N_29511,N_29803);
or UO_2364 (O_2364,N_29965,N_29945);
xor UO_2365 (O_2365,N_29940,N_29536);
nand UO_2366 (O_2366,N_29699,N_29788);
nor UO_2367 (O_2367,N_29722,N_29601);
nor UO_2368 (O_2368,N_29662,N_29766);
xnor UO_2369 (O_2369,N_29867,N_29829);
nand UO_2370 (O_2370,N_29605,N_29533);
and UO_2371 (O_2371,N_29883,N_29831);
nor UO_2372 (O_2372,N_29749,N_29803);
and UO_2373 (O_2373,N_29763,N_29526);
and UO_2374 (O_2374,N_29527,N_29851);
and UO_2375 (O_2375,N_29655,N_29773);
xnor UO_2376 (O_2376,N_29776,N_29523);
xor UO_2377 (O_2377,N_29862,N_29905);
xor UO_2378 (O_2378,N_29867,N_29613);
nand UO_2379 (O_2379,N_29870,N_29563);
xor UO_2380 (O_2380,N_29596,N_29859);
nand UO_2381 (O_2381,N_29687,N_29625);
xor UO_2382 (O_2382,N_29739,N_29503);
xor UO_2383 (O_2383,N_29685,N_29713);
or UO_2384 (O_2384,N_29666,N_29530);
and UO_2385 (O_2385,N_29726,N_29554);
xnor UO_2386 (O_2386,N_29516,N_29905);
and UO_2387 (O_2387,N_29523,N_29790);
nand UO_2388 (O_2388,N_29979,N_29965);
and UO_2389 (O_2389,N_29810,N_29911);
nor UO_2390 (O_2390,N_29720,N_29702);
nor UO_2391 (O_2391,N_29620,N_29873);
xor UO_2392 (O_2392,N_29679,N_29782);
xnor UO_2393 (O_2393,N_29697,N_29926);
and UO_2394 (O_2394,N_29547,N_29814);
or UO_2395 (O_2395,N_29827,N_29509);
and UO_2396 (O_2396,N_29761,N_29789);
and UO_2397 (O_2397,N_29593,N_29823);
nand UO_2398 (O_2398,N_29528,N_29810);
or UO_2399 (O_2399,N_29985,N_29845);
nor UO_2400 (O_2400,N_29873,N_29958);
nand UO_2401 (O_2401,N_29914,N_29503);
and UO_2402 (O_2402,N_29906,N_29980);
nor UO_2403 (O_2403,N_29508,N_29886);
xor UO_2404 (O_2404,N_29677,N_29816);
or UO_2405 (O_2405,N_29551,N_29683);
nor UO_2406 (O_2406,N_29500,N_29646);
xnor UO_2407 (O_2407,N_29520,N_29596);
or UO_2408 (O_2408,N_29723,N_29814);
xor UO_2409 (O_2409,N_29595,N_29503);
or UO_2410 (O_2410,N_29774,N_29978);
nand UO_2411 (O_2411,N_29640,N_29899);
and UO_2412 (O_2412,N_29570,N_29788);
and UO_2413 (O_2413,N_29847,N_29651);
and UO_2414 (O_2414,N_29559,N_29961);
and UO_2415 (O_2415,N_29906,N_29780);
nand UO_2416 (O_2416,N_29723,N_29588);
xnor UO_2417 (O_2417,N_29957,N_29952);
nand UO_2418 (O_2418,N_29753,N_29621);
xor UO_2419 (O_2419,N_29825,N_29700);
nor UO_2420 (O_2420,N_29779,N_29864);
or UO_2421 (O_2421,N_29504,N_29882);
or UO_2422 (O_2422,N_29696,N_29828);
nand UO_2423 (O_2423,N_29934,N_29686);
and UO_2424 (O_2424,N_29802,N_29928);
or UO_2425 (O_2425,N_29556,N_29777);
xor UO_2426 (O_2426,N_29795,N_29975);
or UO_2427 (O_2427,N_29872,N_29599);
and UO_2428 (O_2428,N_29584,N_29817);
nor UO_2429 (O_2429,N_29822,N_29921);
nand UO_2430 (O_2430,N_29794,N_29837);
nand UO_2431 (O_2431,N_29605,N_29907);
xor UO_2432 (O_2432,N_29706,N_29910);
or UO_2433 (O_2433,N_29963,N_29863);
nor UO_2434 (O_2434,N_29558,N_29972);
or UO_2435 (O_2435,N_29857,N_29931);
or UO_2436 (O_2436,N_29548,N_29580);
or UO_2437 (O_2437,N_29707,N_29870);
and UO_2438 (O_2438,N_29518,N_29830);
xnor UO_2439 (O_2439,N_29932,N_29575);
nand UO_2440 (O_2440,N_29542,N_29985);
and UO_2441 (O_2441,N_29756,N_29932);
and UO_2442 (O_2442,N_29576,N_29760);
nor UO_2443 (O_2443,N_29788,N_29865);
nor UO_2444 (O_2444,N_29702,N_29709);
or UO_2445 (O_2445,N_29784,N_29730);
xnor UO_2446 (O_2446,N_29704,N_29860);
or UO_2447 (O_2447,N_29523,N_29671);
xor UO_2448 (O_2448,N_29592,N_29661);
xnor UO_2449 (O_2449,N_29739,N_29569);
xnor UO_2450 (O_2450,N_29617,N_29795);
and UO_2451 (O_2451,N_29799,N_29895);
or UO_2452 (O_2452,N_29578,N_29937);
nand UO_2453 (O_2453,N_29719,N_29624);
nand UO_2454 (O_2454,N_29696,N_29708);
and UO_2455 (O_2455,N_29690,N_29955);
and UO_2456 (O_2456,N_29741,N_29594);
xnor UO_2457 (O_2457,N_29735,N_29731);
or UO_2458 (O_2458,N_29524,N_29611);
nand UO_2459 (O_2459,N_29769,N_29733);
xor UO_2460 (O_2460,N_29789,N_29540);
or UO_2461 (O_2461,N_29578,N_29868);
xor UO_2462 (O_2462,N_29930,N_29904);
and UO_2463 (O_2463,N_29570,N_29599);
or UO_2464 (O_2464,N_29769,N_29726);
xnor UO_2465 (O_2465,N_29927,N_29896);
and UO_2466 (O_2466,N_29943,N_29946);
nor UO_2467 (O_2467,N_29665,N_29652);
and UO_2468 (O_2468,N_29916,N_29980);
nor UO_2469 (O_2469,N_29694,N_29657);
nor UO_2470 (O_2470,N_29833,N_29621);
nor UO_2471 (O_2471,N_29915,N_29795);
nor UO_2472 (O_2472,N_29787,N_29676);
xor UO_2473 (O_2473,N_29753,N_29616);
and UO_2474 (O_2474,N_29806,N_29890);
and UO_2475 (O_2475,N_29996,N_29645);
nand UO_2476 (O_2476,N_29868,N_29836);
nor UO_2477 (O_2477,N_29754,N_29802);
xor UO_2478 (O_2478,N_29768,N_29627);
and UO_2479 (O_2479,N_29654,N_29599);
and UO_2480 (O_2480,N_29754,N_29821);
and UO_2481 (O_2481,N_29808,N_29500);
and UO_2482 (O_2482,N_29805,N_29864);
xnor UO_2483 (O_2483,N_29995,N_29990);
nand UO_2484 (O_2484,N_29879,N_29612);
xor UO_2485 (O_2485,N_29783,N_29735);
or UO_2486 (O_2486,N_29768,N_29967);
nand UO_2487 (O_2487,N_29994,N_29848);
and UO_2488 (O_2488,N_29535,N_29598);
or UO_2489 (O_2489,N_29880,N_29915);
or UO_2490 (O_2490,N_29779,N_29632);
or UO_2491 (O_2491,N_29618,N_29911);
xnor UO_2492 (O_2492,N_29786,N_29721);
xor UO_2493 (O_2493,N_29920,N_29804);
xor UO_2494 (O_2494,N_29803,N_29965);
and UO_2495 (O_2495,N_29764,N_29706);
or UO_2496 (O_2496,N_29786,N_29580);
nor UO_2497 (O_2497,N_29695,N_29884);
nand UO_2498 (O_2498,N_29564,N_29733);
or UO_2499 (O_2499,N_29982,N_29996);
and UO_2500 (O_2500,N_29512,N_29908);
nor UO_2501 (O_2501,N_29838,N_29980);
or UO_2502 (O_2502,N_29530,N_29820);
nand UO_2503 (O_2503,N_29659,N_29543);
and UO_2504 (O_2504,N_29687,N_29968);
xnor UO_2505 (O_2505,N_29569,N_29573);
nor UO_2506 (O_2506,N_29765,N_29877);
xnor UO_2507 (O_2507,N_29939,N_29726);
and UO_2508 (O_2508,N_29811,N_29583);
nand UO_2509 (O_2509,N_29839,N_29907);
or UO_2510 (O_2510,N_29693,N_29701);
and UO_2511 (O_2511,N_29800,N_29515);
xnor UO_2512 (O_2512,N_29966,N_29593);
nand UO_2513 (O_2513,N_29969,N_29786);
or UO_2514 (O_2514,N_29761,N_29561);
xor UO_2515 (O_2515,N_29758,N_29558);
nand UO_2516 (O_2516,N_29744,N_29946);
or UO_2517 (O_2517,N_29539,N_29615);
xnor UO_2518 (O_2518,N_29819,N_29621);
xor UO_2519 (O_2519,N_29787,N_29663);
nor UO_2520 (O_2520,N_29763,N_29554);
xnor UO_2521 (O_2521,N_29581,N_29928);
or UO_2522 (O_2522,N_29674,N_29620);
and UO_2523 (O_2523,N_29811,N_29676);
and UO_2524 (O_2524,N_29594,N_29997);
and UO_2525 (O_2525,N_29511,N_29653);
xor UO_2526 (O_2526,N_29740,N_29985);
nand UO_2527 (O_2527,N_29990,N_29586);
and UO_2528 (O_2528,N_29834,N_29744);
nand UO_2529 (O_2529,N_29588,N_29712);
or UO_2530 (O_2530,N_29756,N_29873);
nand UO_2531 (O_2531,N_29721,N_29620);
and UO_2532 (O_2532,N_29582,N_29687);
nor UO_2533 (O_2533,N_29577,N_29942);
nand UO_2534 (O_2534,N_29548,N_29529);
nand UO_2535 (O_2535,N_29859,N_29763);
nand UO_2536 (O_2536,N_29796,N_29904);
and UO_2537 (O_2537,N_29961,N_29862);
nand UO_2538 (O_2538,N_29736,N_29876);
or UO_2539 (O_2539,N_29522,N_29562);
and UO_2540 (O_2540,N_29577,N_29664);
and UO_2541 (O_2541,N_29652,N_29847);
nand UO_2542 (O_2542,N_29904,N_29752);
and UO_2543 (O_2543,N_29521,N_29975);
nand UO_2544 (O_2544,N_29935,N_29932);
nor UO_2545 (O_2545,N_29525,N_29974);
nand UO_2546 (O_2546,N_29902,N_29820);
or UO_2547 (O_2547,N_29696,N_29992);
or UO_2548 (O_2548,N_29852,N_29505);
nand UO_2549 (O_2549,N_29706,N_29607);
and UO_2550 (O_2550,N_29805,N_29791);
or UO_2551 (O_2551,N_29527,N_29537);
and UO_2552 (O_2552,N_29540,N_29956);
and UO_2553 (O_2553,N_29892,N_29922);
and UO_2554 (O_2554,N_29826,N_29982);
xnor UO_2555 (O_2555,N_29913,N_29528);
xor UO_2556 (O_2556,N_29763,N_29638);
nor UO_2557 (O_2557,N_29524,N_29762);
nor UO_2558 (O_2558,N_29634,N_29669);
nand UO_2559 (O_2559,N_29600,N_29889);
nor UO_2560 (O_2560,N_29615,N_29639);
nor UO_2561 (O_2561,N_29863,N_29933);
xor UO_2562 (O_2562,N_29709,N_29746);
xor UO_2563 (O_2563,N_29513,N_29698);
xor UO_2564 (O_2564,N_29635,N_29502);
nor UO_2565 (O_2565,N_29595,N_29898);
nor UO_2566 (O_2566,N_29738,N_29791);
nand UO_2567 (O_2567,N_29676,N_29836);
or UO_2568 (O_2568,N_29928,N_29589);
nand UO_2569 (O_2569,N_29949,N_29892);
and UO_2570 (O_2570,N_29736,N_29535);
and UO_2571 (O_2571,N_29757,N_29508);
or UO_2572 (O_2572,N_29889,N_29606);
nor UO_2573 (O_2573,N_29938,N_29874);
or UO_2574 (O_2574,N_29628,N_29742);
xor UO_2575 (O_2575,N_29793,N_29786);
xor UO_2576 (O_2576,N_29805,N_29532);
or UO_2577 (O_2577,N_29661,N_29902);
xnor UO_2578 (O_2578,N_29656,N_29610);
or UO_2579 (O_2579,N_29618,N_29907);
and UO_2580 (O_2580,N_29669,N_29623);
xor UO_2581 (O_2581,N_29761,N_29673);
xnor UO_2582 (O_2582,N_29908,N_29884);
xor UO_2583 (O_2583,N_29598,N_29502);
nor UO_2584 (O_2584,N_29884,N_29643);
xor UO_2585 (O_2585,N_29964,N_29688);
and UO_2586 (O_2586,N_29768,N_29820);
nor UO_2587 (O_2587,N_29557,N_29940);
and UO_2588 (O_2588,N_29778,N_29924);
nand UO_2589 (O_2589,N_29657,N_29604);
xor UO_2590 (O_2590,N_29566,N_29841);
nor UO_2591 (O_2591,N_29735,N_29919);
nor UO_2592 (O_2592,N_29562,N_29854);
nand UO_2593 (O_2593,N_29527,N_29842);
or UO_2594 (O_2594,N_29534,N_29942);
or UO_2595 (O_2595,N_29844,N_29939);
and UO_2596 (O_2596,N_29770,N_29527);
xor UO_2597 (O_2597,N_29858,N_29561);
nand UO_2598 (O_2598,N_29900,N_29939);
nand UO_2599 (O_2599,N_29630,N_29817);
nor UO_2600 (O_2600,N_29961,N_29992);
and UO_2601 (O_2601,N_29580,N_29826);
and UO_2602 (O_2602,N_29613,N_29859);
nor UO_2603 (O_2603,N_29699,N_29539);
nand UO_2604 (O_2604,N_29781,N_29979);
nor UO_2605 (O_2605,N_29884,N_29794);
nand UO_2606 (O_2606,N_29683,N_29519);
nand UO_2607 (O_2607,N_29802,N_29701);
nor UO_2608 (O_2608,N_29590,N_29619);
and UO_2609 (O_2609,N_29903,N_29653);
nor UO_2610 (O_2610,N_29932,N_29680);
or UO_2611 (O_2611,N_29643,N_29726);
or UO_2612 (O_2612,N_29690,N_29779);
nand UO_2613 (O_2613,N_29985,N_29545);
or UO_2614 (O_2614,N_29771,N_29934);
xor UO_2615 (O_2615,N_29534,N_29659);
and UO_2616 (O_2616,N_29578,N_29658);
or UO_2617 (O_2617,N_29587,N_29515);
nand UO_2618 (O_2618,N_29882,N_29662);
and UO_2619 (O_2619,N_29573,N_29582);
and UO_2620 (O_2620,N_29749,N_29779);
or UO_2621 (O_2621,N_29838,N_29745);
and UO_2622 (O_2622,N_29509,N_29689);
nand UO_2623 (O_2623,N_29928,N_29827);
nand UO_2624 (O_2624,N_29703,N_29663);
and UO_2625 (O_2625,N_29724,N_29582);
xor UO_2626 (O_2626,N_29684,N_29746);
or UO_2627 (O_2627,N_29534,N_29624);
or UO_2628 (O_2628,N_29704,N_29691);
and UO_2629 (O_2629,N_29888,N_29681);
or UO_2630 (O_2630,N_29646,N_29744);
nand UO_2631 (O_2631,N_29686,N_29942);
nor UO_2632 (O_2632,N_29598,N_29947);
xnor UO_2633 (O_2633,N_29980,N_29890);
and UO_2634 (O_2634,N_29948,N_29905);
or UO_2635 (O_2635,N_29546,N_29903);
or UO_2636 (O_2636,N_29902,N_29655);
or UO_2637 (O_2637,N_29713,N_29866);
and UO_2638 (O_2638,N_29794,N_29547);
nor UO_2639 (O_2639,N_29583,N_29913);
nand UO_2640 (O_2640,N_29942,N_29793);
nand UO_2641 (O_2641,N_29559,N_29878);
or UO_2642 (O_2642,N_29504,N_29783);
or UO_2643 (O_2643,N_29599,N_29868);
and UO_2644 (O_2644,N_29938,N_29880);
xor UO_2645 (O_2645,N_29824,N_29828);
xnor UO_2646 (O_2646,N_29951,N_29762);
and UO_2647 (O_2647,N_29696,N_29970);
or UO_2648 (O_2648,N_29718,N_29882);
xor UO_2649 (O_2649,N_29992,N_29512);
nand UO_2650 (O_2650,N_29510,N_29689);
nand UO_2651 (O_2651,N_29718,N_29542);
xor UO_2652 (O_2652,N_29683,N_29904);
nor UO_2653 (O_2653,N_29670,N_29678);
nand UO_2654 (O_2654,N_29676,N_29840);
or UO_2655 (O_2655,N_29726,N_29666);
nor UO_2656 (O_2656,N_29635,N_29978);
nand UO_2657 (O_2657,N_29672,N_29862);
nor UO_2658 (O_2658,N_29742,N_29525);
and UO_2659 (O_2659,N_29970,N_29712);
and UO_2660 (O_2660,N_29697,N_29973);
nor UO_2661 (O_2661,N_29798,N_29691);
nand UO_2662 (O_2662,N_29548,N_29929);
and UO_2663 (O_2663,N_29594,N_29917);
xnor UO_2664 (O_2664,N_29816,N_29691);
xor UO_2665 (O_2665,N_29880,N_29502);
nand UO_2666 (O_2666,N_29759,N_29905);
nor UO_2667 (O_2667,N_29630,N_29960);
xor UO_2668 (O_2668,N_29929,N_29850);
or UO_2669 (O_2669,N_29919,N_29732);
nor UO_2670 (O_2670,N_29620,N_29611);
nand UO_2671 (O_2671,N_29649,N_29900);
nor UO_2672 (O_2672,N_29849,N_29558);
nand UO_2673 (O_2673,N_29740,N_29581);
nand UO_2674 (O_2674,N_29824,N_29860);
and UO_2675 (O_2675,N_29792,N_29945);
nor UO_2676 (O_2676,N_29768,N_29970);
nand UO_2677 (O_2677,N_29710,N_29673);
and UO_2678 (O_2678,N_29536,N_29635);
nor UO_2679 (O_2679,N_29791,N_29564);
xnor UO_2680 (O_2680,N_29690,N_29693);
xor UO_2681 (O_2681,N_29679,N_29670);
nor UO_2682 (O_2682,N_29895,N_29629);
or UO_2683 (O_2683,N_29885,N_29534);
nand UO_2684 (O_2684,N_29644,N_29851);
or UO_2685 (O_2685,N_29882,N_29831);
and UO_2686 (O_2686,N_29678,N_29939);
nor UO_2687 (O_2687,N_29999,N_29590);
or UO_2688 (O_2688,N_29868,N_29746);
xnor UO_2689 (O_2689,N_29586,N_29607);
xor UO_2690 (O_2690,N_29945,N_29989);
xnor UO_2691 (O_2691,N_29674,N_29673);
or UO_2692 (O_2692,N_29842,N_29533);
and UO_2693 (O_2693,N_29586,N_29860);
xor UO_2694 (O_2694,N_29965,N_29843);
xnor UO_2695 (O_2695,N_29762,N_29516);
nor UO_2696 (O_2696,N_29566,N_29728);
nor UO_2697 (O_2697,N_29742,N_29793);
and UO_2698 (O_2698,N_29896,N_29800);
xor UO_2699 (O_2699,N_29670,N_29948);
xnor UO_2700 (O_2700,N_29745,N_29752);
nand UO_2701 (O_2701,N_29507,N_29658);
or UO_2702 (O_2702,N_29766,N_29669);
or UO_2703 (O_2703,N_29560,N_29535);
nor UO_2704 (O_2704,N_29667,N_29751);
or UO_2705 (O_2705,N_29850,N_29503);
xnor UO_2706 (O_2706,N_29550,N_29696);
and UO_2707 (O_2707,N_29983,N_29873);
and UO_2708 (O_2708,N_29661,N_29564);
nand UO_2709 (O_2709,N_29720,N_29723);
nor UO_2710 (O_2710,N_29994,N_29600);
xor UO_2711 (O_2711,N_29640,N_29802);
nand UO_2712 (O_2712,N_29811,N_29528);
nor UO_2713 (O_2713,N_29878,N_29933);
or UO_2714 (O_2714,N_29732,N_29680);
nand UO_2715 (O_2715,N_29640,N_29552);
or UO_2716 (O_2716,N_29820,N_29512);
nor UO_2717 (O_2717,N_29636,N_29687);
and UO_2718 (O_2718,N_29696,N_29890);
nor UO_2719 (O_2719,N_29738,N_29866);
nand UO_2720 (O_2720,N_29702,N_29905);
xnor UO_2721 (O_2721,N_29702,N_29917);
or UO_2722 (O_2722,N_29888,N_29872);
nor UO_2723 (O_2723,N_29627,N_29804);
xor UO_2724 (O_2724,N_29736,N_29910);
nand UO_2725 (O_2725,N_29893,N_29642);
nand UO_2726 (O_2726,N_29762,N_29859);
or UO_2727 (O_2727,N_29662,N_29968);
xnor UO_2728 (O_2728,N_29970,N_29575);
nand UO_2729 (O_2729,N_29969,N_29575);
nor UO_2730 (O_2730,N_29743,N_29553);
or UO_2731 (O_2731,N_29838,N_29855);
xnor UO_2732 (O_2732,N_29572,N_29820);
or UO_2733 (O_2733,N_29892,N_29606);
xor UO_2734 (O_2734,N_29548,N_29520);
nand UO_2735 (O_2735,N_29699,N_29911);
xor UO_2736 (O_2736,N_29844,N_29722);
or UO_2737 (O_2737,N_29978,N_29857);
and UO_2738 (O_2738,N_29773,N_29925);
nor UO_2739 (O_2739,N_29720,N_29641);
or UO_2740 (O_2740,N_29711,N_29747);
xnor UO_2741 (O_2741,N_29828,N_29800);
nor UO_2742 (O_2742,N_29607,N_29852);
nor UO_2743 (O_2743,N_29710,N_29503);
and UO_2744 (O_2744,N_29872,N_29946);
xor UO_2745 (O_2745,N_29526,N_29831);
or UO_2746 (O_2746,N_29828,N_29837);
or UO_2747 (O_2747,N_29713,N_29525);
or UO_2748 (O_2748,N_29899,N_29819);
xnor UO_2749 (O_2749,N_29775,N_29633);
nor UO_2750 (O_2750,N_29812,N_29745);
and UO_2751 (O_2751,N_29938,N_29654);
xor UO_2752 (O_2752,N_29861,N_29912);
nor UO_2753 (O_2753,N_29982,N_29749);
or UO_2754 (O_2754,N_29745,N_29500);
nand UO_2755 (O_2755,N_29982,N_29705);
nand UO_2756 (O_2756,N_29765,N_29791);
or UO_2757 (O_2757,N_29926,N_29600);
nor UO_2758 (O_2758,N_29789,N_29826);
nor UO_2759 (O_2759,N_29706,N_29692);
nor UO_2760 (O_2760,N_29775,N_29957);
nor UO_2761 (O_2761,N_29572,N_29568);
and UO_2762 (O_2762,N_29795,N_29745);
xnor UO_2763 (O_2763,N_29961,N_29912);
nor UO_2764 (O_2764,N_29963,N_29850);
nor UO_2765 (O_2765,N_29803,N_29541);
or UO_2766 (O_2766,N_29666,N_29997);
xor UO_2767 (O_2767,N_29504,N_29570);
xor UO_2768 (O_2768,N_29948,N_29516);
and UO_2769 (O_2769,N_29919,N_29669);
nor UO_2770 (O_2770,N_29654,N_29535);
or UO_2771 (O_2771,N_29838,N_29600);
or UO_2772 (O_2772,N_29612,N_29763);
nand UO_2773 (O_2773,N_29557,N_29766);
xor UO_2774 (O_2774,N_29796,N_29879);
and UO_2775 (O_2775,N_29586,N_29624);
xnor UO_2776 (O_2776,N_29512,N_29525);
or UO_2777 (O_2777,N_29614,N_29635);
and UO_2778 (O_2778,N_29732,N_29708);
nor UO_2779 (O_2779,N_29582,N_29846);
nand UO_2780 (O_2780,N_29747,N_29712);
nor UO_2781 (O_2781,N_29882,N_29819);
xor UO_2782 (O_2782,N_29886,N_29847);
xnor UO_2783 (O_2783,N_29509,N_29584);
or UO_2784 (O_2784,N_29951,N_29637);
xor UO_2785 (O_2785,N_29604,N_29739);
xnor UO_2786 (O_2786,N_29951,N_29943);
and UO_2787 (O_2787,N_29871,N_29569);
nand UO_2788 (O_2788,N_29531,N_29636);
xnor UO_2789 (O_2789,N_29951,N_29940);
xor UO_2790 (O_2790,N_29702,N_29865);
nand UO_2791 (O_2791,N_29952,N_29584);
nand UO_2792 (O_2792,N_29836,N_29689);
nand UO_2793 (O_2793,N_29718,N_29714);
and UO_2794 (O_2794,N_29751,N_29762);
and UO_2795 (O_2795,N_29544,N_29799);
and UO_2796 (O_2796,N_29806,N_29520);
and UO_2797 (O_2797,N_29522,N_29953);
nand UO_2798 (O_2798,N_29651,N_29501);
xnor UO_2799 (O_2799,N_29515,N_29695);
nand UO_2800 (O_2800,N_29525,N_29892);
xor UO_2801 (O_2801,N_29708,N_29521);
or UO_2802 (O_2802,N_29618,N_29707);
xor UO_2803 (O_2803,N_29674,N_29944);
or UO_2804 (O_2804,N_29616,N_29681);
nor UO_2805 (O_2805,N_29841,N_29645);
xor UO_2806 (O_2806,N_29546,N_29789);
nor UO_2807 (O_2807,N_29996,N_29954);
nor UO_2808 (O_2808,N_29775,N_29550);
or UO_2809 (O_2809,N_29593,N_29923);
and UO_2810 (O_2810,N_29911,N_29575);
nor UO_2811 (O_2811,N_29539,N_29937);
nor UO_2812 (O_2812,N_29694,N_29552);
and UO_2813 (O_2813,N_29925,N_29672);
and UO_2814 (O_2814,N_29563,N_29728);
nand UO_2815 (O_2815,N_29712,N_29874);
nor UO_2816 (O_2816,N_29942,N_29532);
nor UO_2817 (O_2817,N_29523,N_29771);
nor UO_2818 (O_2818,N_29789,N_29852);
nand UO_2819 (O_2819,N_29588,N_29973);
or UO_2820 (O_2820,N_29880,N_29820);
nand UO_2821 (O_2821,N_29957,N_29525);
xor UO_2822 (O_2822,N_29634,N_29598);
nand UO_2823 (O_2823,N_29630,N_29996);
and UO_2824 (O_2824,N_29530,N_29616);
and UO_2825 (O_2825,N_29527,N_29907);
nor UO_2826 (O_2826,N_29773,N_29603);
or UO_2827 (O_2827,N_29639,N_29686);
xor UO_2828 (O_2828,N_29519,N_29866);
xor UO_2829 (O_2829,N_29701,N_29859);
and UO_2830 (O_2830,N_29841,N_29737);
xnor UO_2831 (O_2831,N_29508,N_29776);
xnor UO_2832 (O_2832,N_29702,N_29911);
or UO_2833 (O_2833,N_29851,N_29849);
nand UO_2834 (O_2834,N_29861,N_29585);
nand UO_2835 (O_2835,N_29737,N_29994);
nand UO_2836 (O_2836,N_29598,N_29648);
or UO_2837 (O_2837,N_29760,N_29893);
or UO_2838 (O_2838,N_29613,N_29550);
and UO_2839 (O_2839,N_29944,N_29695);
xnor UO_2840 (O_2840,N_29925,N_29931);
or UO_2841 (O_2841,N_29813,N_29613);
xnor UO_2842 (O_2842,N_29726,N_29709);
nand UO_2843 (O_2843,N_29815,N_29770);
nor UO_2844 (O_2844,N_29837,N_29820);
nor UO_2845 (O_2845,N_29930,N_29856);
or UO_2846 (O_2846,N_29992,N_29815);
nor UO_2847 (O_2847,N_29764,N_29527);
and UO_2848 (O_2848,N_29940,N_29554);
nand UO_2849 (O_2849,N_29661,N_29692);
and UO_2850 (O_2850,N_29903,N_29526);
nand UO_2851 (O_2851,N_29758,N_29979);
nor UO_2852 (O_2852,N_29823,N_29771);
nor UO_2853 (O_2853,N_29905,N_29735);
xnor UO_2854 (O_2854,N_29884,N_29600);
and UO_2855 (O_2855,N_29751,N_29823);
or UO_2856 (O_2856,N_29544,N_29604);
or UO_2857 (O_2857,N_29981,N_29596);
nand UO_2858 (O_2858,N_29578,N_29779);
nand UO_2859 (O_2859,N_29519,N_29725);
nor UO_2860 (O_2860,N_29526,N_29866);
or UO_2861 (O_2861,N_29581,N_29763);
or UO_2862 (O_2862,N_29870,N_29649);
nor UO_2863 (O_2863,N_29545,N_29849);
nand UO_2864 (O_2864,N_29501,N_29848);
nor UO_2865 (O_2865,N_29758,N_29923);
xor UO_2866 (O_2866,N_29602,N_29915);
nor UO_2867 (O_2867,N_29803,N_29866);
nor UO_2868 (O_2868,N_29553,N_29730);
and UO_2869 (O_2869,N_29990,N_29641);
and UO_2870 (O_2870,N_29825,N_29846);
and UO_2871 (O_2871,N_29675,N_29794);
and UO_2872 (O_2872,N_29981,N_29561);
xnor UO_2873 (O_2873,N_29726,N_29513);
nor UO_2874 (O_2874,N_29911,N_29698);
and UO_2875 (O_2875,N_29755,N_29889);
nor UO_2876 (O_2876,N_29960,N_29984);
xor UO_2877 (O_2877,N_29827,N_29681);
nor UO_2878 (O_2878,N_29513,N_29824);
xor UO_2879 (O_2879,N_29562,N_29911);
or UO_2880 (O_2880,N_29691,N_29705);
xnor UO_2881 (O_2881,N_29556,N_29600);
nor UO_2882 (O_2882,N_29891,N_29958);
nand UO_2883 (O_2883,N_29718,N_29764);
nand UO_2884 (O_2884,N_29564,N_29885);
and UO_2885 (O_2885,N_29631,N_29575);
xnor UO_2886 (O_2886,N_29950,N_29559);
and UO_2887 (O_2887,N_29895,N_29517);
xnor UO_2888 (O_2888,N_29862,N_29918);
and UO_2889 (O_2889,N_29703,N_29649);
xnor UO_2890 (O_2890,N_29874,N_29574);
xnor UO_2891 (O_2891,N_29904,N_29909);
or UO_2892 (O_2892,N_29814,N_29554);
xor UO_2893 (O_2893,N_29941,N_29934);
xor UO_2894 (O_2894,N_29692,N_29671);
nor UO_2895 (O_2895,N_29571,N_29901);
nor UO_2896 (O_2896,N_29622,N_29659);
nand UO_2897 (O_2897,N_29513,N_29690);
and UO_2898 (O_2898,N_29791,N_29544);
nand UO_2899 (O_2899,N_29877,N_29603);
and UO_2900 (O_2900,N_29911,N_29916);
nand UO_2901 (O_2901,N_29895,N_29816);
nor UO_2902 (O_2902,N_29682,N_29592);
xnor UO_2903 (O_2903,N_29699,N_29647);
nand UO_2904 (O_2904,N_29700,N_29954);
and UO_2905 (O_2905,N_29588,N_29509);
nand UO_2906 (O_2906,N_29805,N_29618);
xnor UO_2907 (O_2907,N_29790,N_29555);
and UO_2908 (O_2908,N_29732,N_29656);
or UO_2909 (O_2909,N_29563,N_29618);
or UO_2910 (O_2910,N_29823,N_29702);
xor UO_2911 (O_2911,N_29747,N_29746);
or UO_2912 (O_2912,N_29702,N_29935);
or UO_2913 (O_2913,N_29969,N_29776);
and UO_2914 (O_2914,N_29952,N_29848);
nor UO_2915 (O_2915,N_29683,N_29979);
and UO_2916 (O_2916,N_29899,N_29732);
nand UO_2917 (O_2917,N_29590,N_29515);
and UO_2918 (O_2918,N_29573,N_29615);
nand UO_2919 (O_2919,N_29548,N_29738);
and UO_2920 (O_2920,N_29948,N_29618);
or UO_2921 (O_2921,N_29938,N_29518);
or UO_2922 (O_2922,N_29882,N_29841);
xor UO_2923 (O_2923,N_29851,N_29625);
nand UO_2924 (O_2924,N_29879,N_29563);
xor UO_2925 (O_2925,N_29906,N_29504);
nand UO_2926 (O_2926,N_29703,N_29805);
nand UO_2927 (O_2927,N_29865,N_29971);
nand UO_2928 (O_2928,N_29539,N_29556);
xnor UO_2929 (O_2929,N_29992,N_29790);
and UO_2930 (O_2930,N_29942,N_29624);
nor UO_2931 (O_2931,N_29990,N_29899);
nor UO_2932 (O_2932,N_29632,N_29972);
or UO_2933 (O_2933,N_29567,N_29546);
xnor UO_2934 (O_2934,N_29754,N_29661);
xnor UO_2935 (O_2935,N_29901,N_29863);
xnor UO_2936 (O_2936,N_29952,N_29976);
nor UO_2937 (O_2937,N_29624,N_29808);
and UO_2938 (O_2938,N_29773,N_29805);
nor UO_2939 (O_2939,N_29927,N_29953);
or UO_2940 (O_2940,N_29823,N_29687);
and UO_2941 (O_2941,N_29720,N_29614);
xor UO_2942 (O_2942,N_29666,N_29657);
nand UO_2943 (O_2943,N_29769,N_29865);
or UO_2944 (O_2944,N_29542,N_29591);
nor UO_2945 (O_2945,N_29692,N_29665);
or UO_2946 (O_2946,N_29645,N_29824);
or UO_2947 (O_2947,N_29755,N_29814);
and UO_2948 (O_2948,N_29844,N_29626);
and UO_2949 (O_2949,N_29817,N_29632);
nor UO_2950 (O_2950,N_29512,N_29875);
nor UO_2951 (O_2951,N_29779,N_29919);
nand UO_2952 (O_2952,N_29809,N_29582);
and UO_2953 (O_2953,N_29690,N_29880);
nor UO_2954 (O_2954,N_29817,N_29785);
nand UO_2955 (O_2955,N_29796,N_29854);
nand UO_2956 (O_2956,N_29599,N_29752);
or UO_2957 (O_2957,N_29785,N_29550);
nand UO_2958 (O_2958,N_29972,N_29604);
nor UO_2959 (O_2959,N_29798,N_29577);
nand UO_2960 (O_2960,N_29773,N_29640);
nand UO_2961 (O_2961,N_29713,N_29794);
nand UO_2962 (O_2962,N_29931,N_29945);
xnor UO_2963 (O_2963,N_29931,N_29814);
or UO_2964 (O_2964,N_29748,N_29679);
nor UO_2965 (O_2965,N_29712,N_29972);
and UO_2966 (O_2966,N_29702,N_29811);
xor UO_2967 (O_2967,N_29727,N_29600);
xnor UO_2968 (O_2968,N_29837,N_29574);
and UO_2969 (O_2969,N_29862,N_29784);
nor UO_2970 (O_2970,N_29950,N_29958);
xnor UO_2971 (O_2971,N_29534,N_29952);
and UO_2972 (O_2972,N_29748,N_29594);
or UO_2973 (O_2973,N_29602,N_29687);
nor UO_2974 (O_2974,N_29561,N_29500);
nand UO_2975 (O_2975,N_29932,N_29524);
nand UO_2976 (O_2976,N_29650,N_29564);
xor UO_2977 (O_2977,N_29576,N_29776);
nor UO_2978 (O_2978,N_29837,N_29958);
and UO_2979 (O_2979,N_29858,N_29711);
xor UO_2980 (O_2980,N_29628,N_29601);
or UO_2981 (O_2981,N_29931,N_29773);
and UO_2982 (O_2982,N_29517,N_29947);
or UO_2983 (O_2983,N_29677,N_29830);
nor UO_2984 (O_2984,N_29927,N_29628);
nand UO_2985 (O_2985,N_29773,N_29772);
nand UO_2986 (O_2986,N_29910,N_29974);
or UO_2987 (O_2987,N_29824,N_29802);
xor UO_2988 (O_2988,N_29523,N_29873);
xnor UO_2989 (O_2989,N_29863,N_29813);
nand UO_2990 (O_2990,N_29948,N_29733);
nor UO_2991 (O_2991,N_29773,N_29721);
and UO_2992 (O_2992,N_29788,N_29877);
or UO_2993 (O_2993,N_29780,N_29938);
or UO_2994 (O_2994,N_29581,N_29730);
and UO_2995 (O_2995,N_29652,N_29778);
or UO_2996 (O_2996,N_29958,N_29552);
and UO_2997 (O_2997,N_29737,N_29777);
nor UO_2998 (O_2998,N_29626,N_29579);
or UO_2999 (O_2999,N_29975,N_29572);
and UO_3000 (O_3000,N_29951,N_29712);
nor UO_3001 (O_3001,N_29758,N_29613);
xor UO_3002 (O_3002,N_29901,N_29926);
nor UO_3003 (O_3003,N_29543,N_29507);
xnor UO_3004 (O_3004,N_29574,N_29693);
nand UO_3005 (O_3005,N_29996,N_29900);
and UO_3006 (O_3006,N_29930,N_29522);
or UO_3007 (O_3007,N_29630,N_29551);
nand UO_3008 (O_3008,N_29995,N_29833);
or UO_3009 (O_3009,N_29982,N_29785);
xnor UO_3010 (O_3010,N_29516,N_29552);
xnor UO_3011 (O_3011,N_29999,N_29536);
and UO_3012 (O_3012,N_29582,N_29758);
xor UO_3013 (O_3013,N_29840,N_29555);
nand UO_3014 (O_3014,N_29706,N_29536);
nand UO_3015 (O_3015,N_29946,N_29689);
nand UO_3016 (O_3016,N_29551,N_29552);
and UO_3017 (O_3017,N_29890,N_29961);
and UO_3018 (O_3018,N_29518,N_29616);
xor UO_3019 (O_3019,N_29636,N_29545);
nand UO_3020 (O_3020,N_29633,N_29559);
or UO_3021 (O_3021,N_29878,N_29587);
nand UO_3022 (O_3022,N_29714,N_29672);
nor UO_3023 (O_3023,N_29731,N_29514);
xnor UO_3024 (O_3024,N_29765,N_29760);
xnor UO_3025 (O_3025,N_29571,N_29500);
nand UO_3026 (O_3026,N_29711,N_29877);
xor UO_3027 (O_3027,N_29680,N_29580);
nor UO_3028 (O_3028,N_29623,N_29506);
or UO_3029 (O_3029,N_29702,N_29735);
or UO_3030 (O_3030,N_29712,N_29766);
and UO_3031 (O_3031,N_29542,N_29924);
nor UO_3032 (O_3032,N_29844,N_29764);
nand UO_3033 (O_3033,N_29842,N_29703);
nor UO_3034 (O_3034,N_29557,N_29715);
xor UO_3035 (O_3035,N_29740,N_29955);
nand UO_3036 (O_3036,N_29900,N_29859);
xor UO_3037 (O_3037,N_29703,N_29684);
xor UO_3038 (O_3038,N_29730,N_29938);
and UO_3039 (O_3039,N_29659,N_29958);
xor UO_3040 (O_3040,N_29742,N_29576);
nor UO_3041 (O_3041,N_29531,N_29567);
or UO_3042 (O_3042,N_29880,N_29604);
nand UO_3043 (O_3043,N_29933,N_29987);
nor UO_3044 (O_3044,N_29527,N_29510);
and UO_3045 (O_3045,N_29710,N_29599);
xor UO_3046 (O_3046,N_29519,N_29592);
and UO_3047 (O_3047,N_29966,N_29662);
or UO_3048 (O_3048,N_29763,N_29986);
nand UO_3049 (O_3049,N_29635,N_29680);
nor UO_3050 (O_3050,N_29652,N_29746);
nor UO_3051 (O_3051,N_29776,N_29845);
nor UO_3052 (O_3052,N_29994,N_29929);
nor UO_3053 (O_3053,N_29774,N_29545);
and UO_3054 (O_3054,N_29524,N_29872);
nand UO_3055 (O_3055,N_29621,N_29638);
and UO_3056 (O_3056,N_29877,N_29890);
nor UO_3057 (O_3057,N_29564,N_29949);
nor UO_3058 (O_3058,N_29528,N_29803);
nand UO_3059 (O_3059,N_29864,N_29843);
xnor UO_3060 (O_3060,N_29920,N_29964);
and UO_3061 (O_3061,N_29746,N_29641);
xor UO_3062 (O_3062,N_29581,N_29948);
or UO_3063 (O_3063,N_29701,N_29841);
and UO_3064 (O_3064,N_29616,N_29980);
nand UO_3065 (O_3065,N_29583,N_29578);
xnor UO_3066 (O_3066,N_29610,N_29602);
xor UO_3067 (O_3067,N_29543,N_29579);
and UO_3068 (O_3068,N_29541,N_29584);
xnor UO_3069 (O_3069,N_29796,N_29615);
nor UO_3070 (O_3070,N_29761,N_29636);
nand UO_3071 (O_3071,N_29519,N_29979);
nand UO_3072 (O_3072,N_29864,N_29641);
xnor UO_3073 (O_3073,N_29839,N_29589);
nor UO_3074 (O_3074,N_29774,N_29658);
nand UO_3075 (O_3075,N_29799,N_29938);
xor UO_3076 (O_3076,N_29716,N_29691);
nand UO_3077 (O_3077,N_29890,N_29878);
xnor UO_3078 (O_3078,N_29601,N_29554);
and UO_3079 (O_3079,N_29650,N_29759);
nand UO_3080 (O_3080,N_29565,N_29601);
xnor UO_3081 (O_3081,N_29514,N_29763);
nand UO_3082 (O_3082,N_29868,N_29979);
nand UO_3083 (O_3083,N_29732,N_29672);
or UO_3084 (O_3084,N_29627,N_29595);
nand UO_3085 (O_3085,N_29978,N_29947);
or UO_3086 (O_3086,N_29561,N_29770);
nor UO_3087 (O_3087,N_29711,N_29619);
xnor UO_3088 (O_3088,N_29670,N_29686);
nor UO_3089 (O_3089,N_29563,N_29532);
or UO_3090 (O_3090,N_29526,N_29844);
and UO_3091 (O_3091,N_29611,N_29910);
or UO_3092 (O_3092,N_29851,N_29904);
nand UO_3093 (O_3093,N_29800,N_29784);
or UO_3094 (O_3094,N_29604,N_29771);
nand UO_3095 (O_3095,N_29524,N_29534);
and UO_3096 (O_3096,N_29885,N_29841);
nor UO_3097 (O_3097,N_29543,N_29952);
nand UO_3098 (O_3098,N_29606,N_29707);
and UO_3099 (O_3099,N_29919,N_29550);
or UO_3100 (O_3100,N_29951,N_29769);
xor UO_3101 (O_3101,N_29728,N_29510);
nand UO_3102 (O_3102,N_29710,N_29601);
nand UO_3103 (O_3103,N_29959,N_29610);
and UO_3104 (O_3104,N_29982,N_29859);
nand UO_3105 (O_3105,N_29754,N_29537);
xor UO_3106 (O_3106,N_29667,N_29721);
xor UO_3107 (O_3107,N_29607,N_29921);
nor UO_3108 (O_3108,N_29800,N_29553);
xor UO_3109 (O_3109,N_29997,N_29947);
nand UO_3110 (O_3110,N_29785,N_29938);
nor UO_3111 (O_3111,N_29632,N_29735);
nand UO_3112 (O_3112,N_29910,N_29805);
nor UO_3113 (O_3113,N_29691,N_29796);
nand UO_3114 (O_3114,N_29767,N_29710);
and UO_3115 (O_3115,N_29750,N_29675);
and UO_3116 (O_3116,N_29936,N_29582);
xnor UO_3117 (O_3117,N_29748,N_29785);
xnor UO_3118 (O_3118,N_29594,N_29641);
nand UO_3119 (O_3119,N_29892,N_29651);
and UO_3120 (O_3120,N_29960,N_29708);
or UO_3121 (O_3121,N_29598,N_29544);
and UO_3122 (O_3122,N_29531,N_29852);
xor UO_3123 (O_3123,N_29894,N_29854);
and UO_3124 (O_3124,N_29824,N_29851);
nand UO_3125 (O_3125,N_29614,N_29721);
nand UO_3126 (O_3126,N_29568,N_29717);
and UO_3127 (O_3127,N_29638,N_29885);
nor UO_3128 (O_3128,N_29891,N_29615);
and UO_3129 (O_3129,N_29734,N_29724);
nand UO_3130 (O_3130,N_29863,N_29607);
nor UO_3131 (O_3131,N_29536,N_29981);
or UO_3132 (O_3132,N_29880,N_29931);
xnor UO_3133 (O_3133,N_29691,N_29728);
xnor UO_3134 (O_3134,N_29936,N_29943);
or UO_3135 (O_3135,N_29832,N_29968);
xor UO_3136 (O_3136,N_29675,N_29888);
and UO_3137 (O_3137,N_29823,N_29564);
nand UO_3138 (O_3138,N_29948,N_29935);
and UO_3139 (O_3139,N_29722,N_29684);
nor UO_3140 (O_3140,N_29678,N_29760);
xnor UO_3141 (O_3141,N_29967,N_29682);
nand UO_3142 (O_3142,N_29942,N_29575);
and UO_3143 (O_3143,N_29716,N_29924);
or UO_3144 (O_3144,N_29519,N_29783);
or UO_3145 (O_3145,N_29567,N_29707);
or UO_3146 (O_3146,N_29711,N_29602);
nor UO_3147 (O_3147,N_29585,N_29524);
nor UO_3148 (O_3148,N_29999,N_29902);
nand UO_3149 (O_3149,N_29808,N_29539);
or UO_3150 (O_3150,N_29801,N_29674);
and UO_3151 (O_3151,N_29502,N_29931);
or UO_3152 (O_3152,N_29743,N_29769);
or UO_3153 (O_3153,N_29551,N_29590);
nor UO_3154 (O_3154,N_29680,N_29570);
or UO_3155 (O_3155,N_29665,N_29718);
nand UO_3156 (O_3156,N_29694,N_29819);
nand UO_3157 (O_3157,N_29833,N_29780);
and UO_3158 (O_3158,N_29936,N_29799);
nor UO_3159 (O_3159,N_29902,N_29887);
xnor UO_3160 (O_3160,N_29795,N_29866);
nand UO_3161 (O_3161,N_29540,N_29742);
nor UO_3162 (O_3162,N_29620,N_29747);
xnor UO_3163 (O_3163,N_29851,N_29981);
nor UO_3164 (O_3164,N_29911,N_29679);
and UO_3165 (O_3165,N_29579,N_29980);
or UO_3166 (O_3166,N_29653,N_29712);
and UO_3167 (O_3167,N_29839,N_29799);
nor UO_3168 (O_3168,N_29876,N_29955);
and UO_3169 (O_3169,N_29782,N_29795);
and UO_3170 (O_3170,N_29679,N_29829);
xnor UO_3171 (O_3171,N_29515,N_29950);
nor UO_3172 (O_3172,N_29941,N_29649);
nand UO_3173 (O_3173,N_29765,N_29605);
nand UO_3174 (O_3174,N_29577,N_29587);
nor UO_3175 (O_3175,N_29566,N_29593);
or UO_3176 (O_3176,N_29587,N_29657);
xnor UO_3177 (O_3177,N_29984,N_29880);
or UO_3178 (O_3178,N_29784,N_29562);
nor UO_3179 (O_3179,N_29865,N_29777);
nor UO_3180 (O_3180,N_29670,N_29855);
and UO_3181 (O_3181,N_29525,N_29869);
nor UO_3182 (O_3182,N_29828,N_29753);
nor UO_3183 (O_3183,N_29996,N_29734);
nand UO_3184 (O_3184,N_29867,N_29528);
xor UO_3185 (O_3185,N_29964,N_29882);
xnor UO_3186 (O_3186,N_29506,N_29800);
xor UO_3187 (O_3187,N_29868,N_29989);
and UO_3188 (O_3188,N_29922,N_29544);
and UO_3189 (O_3189,N_29845,N_29906);
nand UO_3190 (O_3190,N_29534,N_29704);
or UO_3191 (O_3191,N_29637,N_29582);
nand UO_3192 (O_3192,N_29594,N_29504);
or UO_3193 (O_3193,N_29801,N_29707);
xnor UO_3194 (O_3194,N_29562,N_29885);
or UO_3195 (O_3195,N_29959,N_29509);
nor UO_3196 (O_3196,N_29609,N_29924);
and UO_3197 (O_3197,N_29804,N_29598);
xnor UO_3198 (O_3198,N_29772,N_29657);
nand UO_3199 (O_3199,N_29770,N_29641);
and UO_3200 (O_3200,N_29950,N_29981);
xor UO_3201 (O_3201,N_29694,N_29985);
xnor UO_3202 (O_3202,N_29509,N_29765);
xor UO_3203 (O_3203,N_29858,N_29760);
nand UO_3204 (O_3204,N_29805,N_29529);
xor UO_3205 (O_3205,N_29659,N_29655);
xor UO_3206 (O_3206,N_29677,N_29903);
or UO_3207 (O_3207,N_29811,N_29733);
nor UO_3208 (O_3208,N_29773,N_29875);
nand UO_3209 (O_3209,N_29805,N_29803);
nor UO_3210 (O_3210,N_29525,N_29700);
xnor UO_3211 (O_3211,N_29546,N_29813);
or UO_3212 (O_3212,N_29956,N_29631);
xor UO_3213 (O_3213,N_29740,N_29624);
nand UO_3214 (O_3214,N_29623,N_29644);
nand UO_3215 (O_3215,N_29860,N_29743);
and UO_3216 (O_3216,N_29504,N_29868);
and UO_3217 (O_3217,N_29981,N_29943);
nand UO_3218 (O_3218,N_29580,N_29613);
nand UO_3219 (O_3219,N_29787,N_29817);
nor UO_3220 (O_3220,N_29749,N_29685);
nand UO_3221 (O_3221,N_29751,N_29513);
nand UO_3222 (O_3222,N_29584,N_29942);
xor UO_3223 (O_3223,N_29924,N_29621);
nand UO_3224 (O_3224,N_29629,N_29930);
xor UO_3225 (O_3225,N_29951,N_29883);
nand UO_3226 (O_3226,N_29740,N_29714);
nor UO_3227 (O_3227,N_29675,N_29663);
or UO_3228 (O_3228,N_29691,N_29996);
nand UO_3229 (O_3229,N_29910,N_29793);
nand UO_3230 (O_3230,N_29574,N_29635);
nor UO_3231 (O_3231,N_29677,N_29837);
nand UO_3232 (O_3232,N_29825,N_29501);
nor UO_3233 (O_3233,N_29704,N_29532);
or UO_3234 (O_3234,N_29881,N_29899);
nand UO_3235 (O_3235,N_29787,N_29588);
nor UO_3236 (O_3236,N_29771,N_29684);
or UO_3237 (O_3237,N_29987,N_29596);
and UO_3238 (O_3238,N_29594,N_29604);
nand UO_3239 (O_3239,N_29935,N_29589);
or UO_3240 (O_3240,N_29689,N_29735);
and UO_3241 (O_3241,N_29548,N_29850);
nor UO_3242 (O_3242,N_29744,N_29899);
nand UO_3243 (O_3243,N_29559,N_29730);
and UO_3244 (O_3244,N_29839,N_29855);
and UO_3245 (O_3245,N_29921,N_29839);
xnor UO_3246 (O_3246,N_29923,N_29668);
xnor UO_3247 (O_3247,N_29595,N_29569);
nor UO_3248 (O_3248,N_29577,N_29801);
xnor UO_3249 (O_3249,N_29935,N_29758);
xnor UO_3250 (O_3250,N_29873,N_29970);
nor UO_3251 (O_3251,N_29811,N_29706);
and UO_3252 (O_3252,N_29502,N_29872);
and UO_3253 (O_3253,N_29529,N_29630);
nand UO_3254 (O_3254,N_29590,N_29642);
nand UO_3255 (O_3255,N_29879,N_29955);
or UO_3256 (O_3256,N_29678,N_29570);
nand UO_3257 (O_3257,N_29871,N_29523);
nand UO_3258 (O_3258,N_29586,N_29972);
nand UO_3259 (O_3259,N_29839,N_29919);
and UO_3260 (O_3260,N_29930,N_29747);
nor UO_3261 (O_3261,N_29522,N_29613);
and UO_3262 (O_3262,N_29580,N_29842);
nand UO_3263 (O_3263,N_29708,N_29506);
nor UO_3264 (O_3264,N_29915,N_29555);
or UO_3265 (O_3265,N_29796,N_29908);
xor UO_3266 (O_3266,N_29635,N_29938);
or UO_3267 (O_3267,N_29964,N_29511);
xor UO_3268 (O_3268,N_29825,N_29588);
and UO_3269 (O_3269,N_29837,N_29955);
or UO_3270 (O_3270,N_29979,N_29631);
nor UO_3271 (O_3271,N_29564,N_29771);
nand UO_3272 (O_3272,N_29523,N_29549);
nand UO_3273 (O_3273,N_29821,N_29561);
and UO_3274 (O_3274,N_29840,N_29759);
and UO_3275 (O_3275,N_29990,N_29863);
and UO_3276 (O_3276,N_29898,N_29891);
or UO_3277 (O_3277,N_29573,N_29807);
and UO_3278 (O_3278,N_29788,N_29997);
or UO_3279 (O_3279,N_29960,N_29719);
nor UO_3280 (O_3280,N_29919,N_29597);
xnor UO_3281 (O_3281,N_29678,N_29534);
or UO_3282 (O_3282,N_29965,N_29926);
nand UO_3283 (O_3283,N_29899,N_29827);
nand UO_3284 (O_3284,N_29624,N_29749);
xnor UO_3285 (O_3285,N_29979,N_29609);
xor UO_3286 (O_3286,N_29819,N_29623);
xor UO_3287 (O_3287,N_29636,N_29725);
xor UO_3288 (O_3288,N_29953,N_29577);
and UO_3289 (O_3289,N_29981,N_29530);
xor UO_3290 (O_3290,N_29531,N_29820);
nor UO_3291 (O_3291,N_29596,N_29917);
and UO_3292 (O_3292,N_29721,N_29908);
or UO_3293 (O_3293,N_29517,N_29536);
xnor UO_3294 (O_3294,N_29505,N_29887);
xor UO_3295 (O_3295,N_29698,N_29969);
xnor UO_3296 (O_3296,N_29559,N_29589);
or UO_3297 (O_3297,N_29972,N_29881);
xor UO_3298 (O_3298,N_29826,N_29871);
or UO_3299 (O_3299,N_29504,N_29996);
nor UO_3300 (O_3300,N_29663,N_29646);
nor UO_3301 (O_3301,N_29680,N_29922);
and UO_3302 (O_3302,N_29976,N_29505);
nor UO_3303 (O_3303,N_29733,N_29513);
or UO_3304 (O_3304,N_29945,N_29987);
nor UO_3305 (O_3305,N_29652,N_29543);
and UO_3306 (O_3306,N_29870,N_29834);
nor UO_3307 (O_3307,N_29875,N_29695);
nor UO_3308 (O_3308,N_29724,N_29924);
xor UO_3309 (O_3309,N_29686,N_29619);
nand UO_3310 (O_3310,N_29677,N_29704);
xnor UO_3311 (O_3311,N_29947,N_29552);
and UO_3312 (O_3312,N_29732,N_29943);
nand UO_3313 (O_3313,N_29755,N_29638);
or UO_3314 (O_3314,N_29503,N_29508);
or UO_3315 (O_3315,N_29592,N_29940);
xnor UO_3316 (O_3316,N_29885,N_29886);
xor UO_3317 (O_3317,N_29834,N_29806);
or UO_3318 (O_3318,N_29569,N_29910);
nor UO_3319 (O_3319,N_29816,N_29902);
and UO_3320 (O_3320,N_29826,N_29653);
and UO_3321 (O_3321,N_29511,N_29859);
nand UO_3322 (O_3322,N_29975,N_29820);
and UO_3323 (O_3323,N_29957,N_29539);
xnor UO_3324 (O_3324,N_29797,N_29704);
xnor UO_3325 (O_3325,N_29678,N_29971);
nor UO_3326 (O_3326,N_29584,N_29769);
nor UO_3327 (O_3327,N_29986,N_29880);
xor UO_3328 (O_3328,N_29789,N_29609);
nand UO_3329 (O_3329,N_29546,N_29985);
xnor UO_3330 (O_3330,N_29762,N_29721);
nand UO_3331 (O_3331,N_29935,N_29727);
and UO_3332 (O_3332,N_29894,N_29948);
and UO_3333 (O_3333,N_29734,N_29764);
xnor UO_3334 (O_3334,N_29741,N_29938);
nand UO_3335 (O_3335,N_29696,N_29810);
nand UO_3336 (O_3336,N_29639,N_29954);
or UO_3337 (O_3337,N_29858,N_29659);
nand UO_3338 (O_3338,N_29701,N_29944);
xnor UO_3339 (O_3339,N_29770,N_29795);
or UO_3340 (O_3340,N_29564,N_29749);
nand UO_3341 (O_3341,N_29644,N_29695);
or UO_3342 (O_3342,N_29751,N_29884);
or UO_3343 (O_3343,N_29791,N_29681);
xor UO_3344 (O_3344,N_29814,N_29974);
or UO_3345 (O_3345,N_29627,N_29531);
nor UO_3346 (O_3346,N_29992,N_29855);
or UO_3347 (O_3347,N_29904,N_29608);
xnor UO_3348 (O_3348,N_29801,N_29721);
nand UO_3349 (O_3349,N_29975,N_29659);
and UO_3350 (O_3350,N_29748,N_29704);
or UO_3351 (O_3351,N_29877,N_29863);
nor UO_3352 (O_3352,N_29667,N_29534);
nor UO_3353 (O_3353,N_29832,N_29698);
nand UO_3354 (O_3354,N_29785,N_29562);
nand UO_3355 (O_3355,N_29746,N_29719);
nor UO_3356 (O_3356,N_29988,N_29729);
nor UO_3357 (O_3357,N_29842,N_29877);
nor UO_3358 (O_3358,N_29655,N_29894);
nor UO_3359 (O_3359,N_29563,N_29884);
and UO_3360 (O_3360,N_29620,N_29764);
nand UO_3361 (O_3361,N_29567,N_29691);
or UO_3362 (O_3362,N_29744,N_29855);
xnor UO_3363 (O_3363,N_29658,N_29544);
nor UO_3364 (O_3364,N_29694,N_29592);
and UO_3365 (O_3365,N_29999,N_29566);
and UO_3366 (O_3366,N_29645,N_29550);
or UO_3367 (O_3367,N_29546,N_29524);
xnor UO_3368 (O_3368,N_29810,N_29510);
nor UO_3369 (O_3369,N_29942,N_29503);
nand UO_3370 (O_3370,N_29576,N_29659);
nand UO_3371 (O_3371,N_29653,N_29915);
or UO_3372 (O_3372,N_29824,N_29720);
or UO_3373 (O_3373,N_29797,N_29603);
xnor UO_3374 (O_3374,N_29525,N_29522);
xnor UO_3375 (O_3375,N_29522,N_29741);
or UO_3376 (O_3376,N_29591,N_29589);
nand UO_3377 (O_3377,N_29706,N_29713);
and UO_3378 (O_3378,N_29789,N_29867);
xnor UO_3379 (O_3379,N_29812,N_29882);
xor UO_3380 (O_3380,N_29671,N_29923);
xor UO_3381 (O_3381,N_29887,N_29533);
xnor UO_3382 (O_3382,N_29978,N_29650);
nor UO_3383 (O_3383,N_29671,N_29915);
or UO_3384 (O_3384,N_29965,N_29958);
or UO_3385 (O_3385,N_29865,N_29899);
xor UO_3386 (O_3386,N_29961,N_29514);
nand UO_3387 (O_3387,N_29656,N_29806);
nor UO_3388 (O_3388,N_29803,N_29846);
xor UO_3389 (O_3389,N_29690,N_29652);
nor UO_3390 (O_3390,N_29674,N_29872);
and UO_3391 (O_3391,N_29715,N_29726);
and UO_3392 (O_3392,N_29811,N_29506);
nand UO_3393 (O_3393,N_29664,N_29897);
nand UO_3394 (O_3394,N_29766,N_29815);
and UO_3395 (O_3395,N_29626,N_29774);
or UO_3396 (O_3396,N_29861,N_29674);
nor UO_3397 (O_3397,N_29589,N_29552);
and UO_3398 (O_3398,N_29915,N_29929);
xnor UO_3399 (O_3399,N_29733,N_29601);
or UO_3400 (O_3400,N_29857,N_29585);
and UO_3401 (O_3401,N_29902,N_29826);
or UO_3402 (O_3402,N_29791,N_29946);
nor UO_3403 (O_3403,N_29558,N_29715);
xor UO_3404 (O_3404,N_29848,N_29979);
or UO_3405 (O_3405,N_29592,N_29650);
and UO_3406 (O_3406,N_29567,N_29982);
and UO_3407 (O_3407,N_29978,N_29605);
xor UO_3408 (O_3408,N_29556,N_29968);
or UO_3409 (O_3409,N_29689,N_29691);
nand UO_3410 (O_3410,N_29568,N_29505);
nand UO_3411 (O_3411,N_29703,N_29726);
or UO_3412 (O_3412,N_29842,N_29676);
nand UO_3413 (O_3413,N_29583,N_29768);
or UO_3414 (O_3414,N_29949,N_29856);
nand UO_3415 (O_3415,N_29564,N_29863);
or UO_3416 (O_3416,N_29801,N_29770);
nor UO_3417 (O_3417,N_29779,N_29914);
nor UO_3418 (O_3418,N_29502,N_29715);
or UO_3419 (O_3419,N_29552,N_29959);
nand UO_3420 (O_3420,N_29746,N_29581);
nand UO_3421 (O_3421,N_29607,N_29744);
nor UO_3422 (O_3422,N_29926,N_29764);
and UO_3423 (O_3423,N_29609,N_29708);
nor UO_3424 (O_3424,N_29859,N_29868);
xor UO_3425 (O_3425,N_29743,N_29872);
or UO_3426 (O_3426,N_29647,N_29755);
nand UO_3427 (O_3427,N_29959,N_29730);
nand UO_3428 (O_3428,N_29762,N_29632);
nand UO_3429 (O_3429,N_29806,N_29894);
or UO_3430 (O_3430,N_29622,N_29635);
and UO_3431 (O_3431,N_29867,N_29757);
xnor UO_3432 (O_3432,N_29619,N_29831);
or UO_3433 (O_3433,N_29668,N_29943);
nand UO_3434 (O_3434,N_29640,N_29887);
nand UO_3435 (O_3435,N_29798,N_29595);
and UO_3436 (O_3436,N_29915,N_29682);
nor UO_3437 (O_3437,N_29904,N_29795);
or UO_3438 (O_3438,N_29555,N_29987);
nand UO_3439 (O_3439,N_29791,N_29516);
nand UO_3440 (O_3440,N_29913,N_29514);
xnor UO_3441 (O_3441,N_29530,N_29858);
nor UO_3442 (O_3442,N_29677,N_29542);
or UO_3443 (O_3443,N_29956,N_29715);
and UO_3444 (O_3444,N_29801,N_29875);
or UO_3445 (O_3445,N_29561,N_29697);
nand UO_3446 (O_3446,N_29759,N_29685);
xnor UO_3447 (O_3447,N_29624,N_29913);
nand UO_3448 (O_3448,N_29690,N_29906);
nand UO_3449 (O_3449,N_29955,N_29819);
nor UO_3450 (O_3450,N_29768,N_29878);
and UO_3451 (O_3451,N_29624,N_29774);
or UO_3452 (O_3452,N_29643,N_29963);
or UO_3453 (O_3453,N_29770,N_29769);
xnor UO_3454 (O_3454,N_29902,N_29894);
or UO_3455 (O_3455,N_29598,N_29809);
nand UO_3456 (O_3456,N_29621,N_29926);
or UO_3457 (O_3457,N_29839,N_29867);
and UO_3458 (O_3458,N_29583,N_29643);
nand UO_3459 (O_3459,N_29948,N_29891);
xor UO_3460 (O_3460,N_29805,N_29918);
nand UO_3461 (O_3461,N_29691,N_29791);
or UO_3462 (O_3462,N_29938,N_29757);
nor UO_3463 (O_3463,N_29636,N_29997);
or UO_3464 (O_3464,N_29749,N_29529);
xnor UO_3465 (O_3465,N_29928,N_29726);
xnor UO_3466 (O_3466,N_29757,N_29699);
or UO_3467 (O_3467,N_29739,N_29647);
nor UO_3468 (O_3468,N_29629,N_29905);
and UO_3469 (O_3469,N_29647,N_29771);
xor UO_3470 (O_3470,N_29552,N_29787);
nand UO_3471 (O_3471,N_29561,N_29548);
nand UO_3472 (O_3472,N_29946,N_29881);
nor UO_3473 (O_3473,N_29632,N_29757);
and UO_3474 (O_3474,N_29867,N_29737);
and UO_3475 (O_3475,N_29813,N_29578);
nand UO_3476 (O_3476,N_29707,N_29782);
and UO_3477 (O_3477,N_29735,N_29744);
xor UO_3478 (O_3478,N_29571,N_29933);
xnor UO_3479 (O_3479,N_29639,N_29649);
nor UO_3480 (O_3480,N_29595,N_29923);
nor UO_3481 (O_3481,N_29609,N_29936);
or UO_3482 (O_3482,N_29581,N_29970);
nor UO_3483 (O_3483,N_29844,N_29624);
or UO_3484 (O_3484,N_29771,N_29584);
and UO_3485 (O_3485,N_29652,N_29989);
nor UO_3486 (O_3486,N_29993,N_29510);
xor UO_3487 (O_3487,N_29779,N_29629);
xnor UO_3488 (O_3488,N_29834,N_29812);
and UO_3489 (O_3489,N_29805,N_29507);
nand UO_3490 (O_3490,N_29870,N_29536);
nor UO_3491 (O_3491,N_29885,N_29649);
xor UO_3492 (O_3492,N_29615,N_29769);
and UO_3493 (O_3493,N_29704,N_29870);
nand UO_3494 (O_3494,N_29576,N_29708);
xnor UO_3495 (O_3495,N_29560,N_29932);
and UO_3496 (O_3496,N_29932,N_29536);
and UO_3497 (O_3497,N_29681,N_29820);
nand UO_3498 (O_3498,N_29742,N_29938);
nor UO_3499 (O_3499,N_29746,N_29722);
endmodule