module basic_5000_50000_5000_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_4495,In_3831);
and U1 (N_1,In_3625,In_2004);
nand U2 (N_2,In_2428,In_3656);
and U3 (N_3,In_2397,In_2163);
nand U4 (N_4,In_362,In_2944);
and U5 (N_5,In_2520,In_252);
nor U6 (N_6,In_4414,In_3007);
xor U7 (N_7,In_601,In_3537);
nor U8 (N_8,In_4057,In_2607);
nand U9 (N_9,In_1393,In_4360);
nand U10 (N_10,In_3265,In_1022);
xor U11 (N_11,In_1792,In_4422);
nor U12 (N_12,In_496,In_3660);
nor U13 (N_13,In_2227,In_1424);
nor U14 (N_14,In_2918,In_505);
and U15 (N_15,In_4949,In_4410);
xor U16 (N_16,In_3358,In_4905);
and U17 (N_17,In_4875,In_373);
and U18 (N_18,In_1985,In_3426);
nor U19 (N_19,In_1690,In_2613);
xnor U20 (N_20,In_3251,In_2655);
or U21 (N_21,In_2186,In_2233);
nor U22 (N_22,In_3858,In_3521);
nand U23 (N_23,In_3614,In_2260);
and U24 (N_24,In_1794,In_2787);
and U25 (N_25,In_3244,In_804);
xor U26 (N_26,In_3290,In_1636);
or U27 (N_27,In_4567,In_265);
or U28 (N_28,In_4860,In_1405);
xor U29 (N_29,In_2809,In_3117);
nand U30 (N_30,In_855,In_3338);
and U31 (N_31,In_4008,In_153);
nand U32 (N_32,In_3112,In_3003);
and U33 (N_33,In_1228,In_60);
nand U34 (N_34,In_3565,In_4144);
nor U35 (N_35,In_2189,In_995);
or U36 (N_36,In_4430,In_4336);
nor U37 (N_37,In_2768,In_2465);
and U38 (N_38,In_3506,In_4505);
xnor U39 (N_39,In_4465,In_1944);
xor U40 (N_40,In_2627,In_2468);
nand U41 (N_41,In_2568,In_2120);
or U42 (N_42,In_1302,In_1459);
or U43 (N_43,In_4326,In_114);
nor U44 (N_44,In_4089,In_4285);
and U45 (N_45,In_2179,In_3045);
nand U46 (N_46,In_165,In_3733);
and U47 (N_47,In_664,In_3842);
nor U48 (N_48,In_2467,In_3115);
nor U49 (N_49,In_1036,In_1037);
nor U50 (N_50,In_885,In_4373);
and U51 (N_51,In_4867,In_2068);
nor U52 (N_52,In_1583,In_1127);
and U53 (N_53,In_4247,In_1322);
nand U54 (N_54,In_4684,In_1177);
and U55 (N_55,In_2563,In_1525);
or U56 (N_56,In_143,In_2008);
xor U57 (N_57,In_3905,In_1708);
or U58 (N_58,In_2891,In_3104);
nand U59 (N_59,In_4502,In_4947);
nor U60 (N_60,In_4726,In_3659);
and U61 (N_61,In_1339,In_4850);
xor U62 (N_62,In_923,In_1672);
xor U63 (N_63,In_1745,In_2528);
nand U64 (N_64,In_4718,In_3632);
nor U65 (N_65,In_3712,In_4621);
xnor U66 (N_66,In_2991,In_4912);
nor U67 (N_67,In_3095,In_4538);
nor U68 (N_68,In_4170,In_3339);
and U69 (N_69,In_1810,In_3086);
and U70 (N_70,In_4943,In_964);
nor U71 (N_71,In_4193,In_1232);
or U72 (N_72,In_1924,In_746);
nand U73 (N_73,In_3217,In_1585);
and U74 (N_74,In_2533,In_1046);
nand U75 (N_75,In_3892,In_2405);
and U76 (N_76,In_2660,In_2806);
nor U77 (N_77,In_949,In_2093);
nor U78 (N_78,In_4711,In_3859);
or U79 (N_79,In_1989,In_3765);
and U80 (N_80,In_2170,In_2460);
xnor U81 (N_81,In_172,In_4512);
xor U82 (N_82,In_517,In_2353);
nor U83 (N_83,In_669,In_1088);
nand U84 (N_84,In_3331,In_4289);
nand U85 (N_85,In_3710,In_2683);
xor U86 (N_86,In_1002,In_3300);
and U87 (N_87,In_879,In_3414);
nor U88 (N_88,In_1194,In_4937);
or U89 (N_89,In_2536,In_3566);
nor U90 (N_90,In_4664,In_3243);
nand U91 (N_91,In_3544,In_1237);
nor U92 (N_92,In_2814,In_4794);
nand U93 (N_93,In_139,In_1562);
and U94 (N_94,In_3763,In_1410);
and U95 (N_95,In_1430,In_4442);
xor U96 (N_96,In_1229,In_1192);
nor U97 (N_97,In_203,In_3547);
and U98 (N_98,In_1130,In_1533);
nand U99 (N_99,In_2220,In_4079);
or U100 (N_100,In_385,In_4559);
or U101 (N_101,In_1695,In_1378);
nor U102 (N_102,In_4676,In_3820);
or U103 (N_103,In_3114,In_957);
nor U104 (N_104,In_589,In_3098);
xor U105 (N_105,In_2724,In_3420);
nor U106 (N_106,In_3155,In_4120);
xnor U107 (N_107,In_1581,In_4223);
nand U108 (N_108,In_1815,In_2401);
nand U109 (N_109,In_2129,In_1738);
nand U110 (N_110,In_3536,In_377);
nor U111 (N_111,In_4695,In_3948);
nor U112 (N_112,In_2291,In_1233);
or U113 (N_113,In_2156,In_4760);
nand U114 (N_114,In_1154,In_599);
nor U115 (N_115,In_3514,In_3289);
nand U116 (N_116,In_2750,In_1556);
nand U117 (N_117,In_809,In_616);
nand U118 (N_118,In_2522,In_7);
xor U119 (N_119,In_3951,In_2992);
or U120 (N_120,In_4790,In_711);
or U121 (N_121,In_1915,In_2584);
nor U122 (N_122,In_4513,In_1824);
or U123 (N_123,In_4169,In_3978);
nand U124 (N_124,In_2032,In_2288);
nand U125 (N_125,In_2897,In_2331);
or U126 (N_126,In_3938,In_4549);
nor U127 (N_127,In_886,In_1913);
and U128 (N_128,In_1171,In_1883);
xor U129 (N_129,In_3224,In_77);
nor U130 (N_130,In_4669,In_3286);
and U131 (N_131,In_1015,In_4424);
xnor U132 (N_132,In_1683,In_2682);
xor U133 (N_133,In_3987,In_2577);
nand U134 (N_134,In_3406,In_1251);
nor U135 (N_135,In_4811,In_3277);
nand U136 (N_136,In_877,In_1529);
and U137 (N_137,In_4374,In_2681);
and U138 (N_138,In_872,In_4342);
xor U139 (N_139,In_3337,In_240);
nor U140 (N_140,In_4920,In_4459);
nor U141 (N_141,In_2208,In_1890);
and U142 (N_142,In_1504,In_85);
or U143 (N_143,In_2734,In_4400);
nand U144 (N_144,In_2524,In_4659);
and U145 (N_145,In_132,In_1160);
and U146 (N_146,In_3890,In_445);
nor U147 (N_147,In_1183,In_1618);
nor U148 (N_148,In_4652,In_2035);
nor U149 (N_149,In_3022,In_4443);
nor U150 (N_150,In_1869,In_2138);
xnor U151 (N_151,In_520,In_3245);
nor U152 (N_152,In_2708,In_1575);
and U153 (N_153,In_54,In_1699);
xor U154 (N_154,In_3485,In_4340);
and U155 (N_155,In_3767,In_3852);
or U156 (N_156,In_2791,In_233);
nor U157 (N_157,In_2307,In_1327);
nor U158 (N_158,In_4849,In_777);
nor U159 (N_159,In_2235,In_981);
nand U160 (N_160,In_111,In_3599);
xor U161 (N_161,In_1217,In_334);
nand U162 (N_162,In_3190,In_1244);
nand U163 (N_163,In_2075,In_2966);
nand U164 (N_164,In_3351,In_941);
and U165 (N_165,In_2843,In_3979);
and U166 (N_166,In_83,In_3053);
and U167 (N_167,In_400,In_237);
xor U168 (N_168,In_2476,In_2558);
xnor U169 (N_169,In_2670,In_4011);
nand U170 (N_170,In_2811,In_454);
or U171 (N_171,In_3076,In_4174);
nor U172 (N_172,In_3356,In_34);
nor U173 (N_173,In_2478,In_4069);
nand U174 (N_174,In_4447,In_4451);
nor U175 (N_175,In_3228,In_1920);
nand U176 (N_176,In_1990,In_2596);
nand U177 (N_177,In_51,In_3094);
and U178 (N_178,In_3968,In_486);
nor U179 (N_179,In_3511,In_1628);
and U180 (N_180,In_4387,In_4488);
or U181 (N_181,In_1835,In_906);
nor U182 (N_182,In_4545,In_4017);
and U183 (N_183,In_849,In_3538);
or U184 (N_184,In_4412,In_4118);
or U185 (N_185,In_943,In_4454);
nand U186 (N_186,In_2790,In_3330);
nor U187 (N_187,In_4204,In_3382);
nand U188 (N_188,In_822,In_480);
nand U189 (N_189,In_1467,In_2690);
or U190 (N_190,In_4657,In_3834);
nand U191 (N_191,In_4561,In_3397);
and U192 (N_192,In_1381,In_1145);
xor U193 (N_193,In_2269,In_3383);
xor U194 (N_194,In_2025,In_3605);
and U195 (N_195,In_2244,In_3340);
nor U196 (N_196,In_1742,In_2513);
xnor U197 (N_197,In_1105,In_4093);
or U198 (N_198,In_4745,In_1993);
or U199 (N_199,In_1552,In_1879);
nor U200 (N_200,In_2447,In_3100);
nand U201 (N_201,In_652,In_495);
or U202 (N_202,In_4681,In_3567);
or U203 (N_203,In_3070,In_4101);
or U204 (N_204,In_1468,In_3980);
nand U205 (N_205,In_2411,In_3922);
nor U206 (N_206,In_840,In_810);
or U207 (N_207,In_2862,In_549);
and U208 (N_208,In_1173,In_4496);
xnor U209 (N_209,In_2117,In_870);
xor U210 (N_210,In_4540,In_4484);
and U211 (N_211,In_3046,In_4604);
xnor U212 (N_212,In_627,In_2634);
nor U213 (N_213,In_3012,In_540);
xor U214 (N_214,In_2543,In_1266);
nor U215 (N_215,In_2802,In_1404);
nor U216 (N_216,In_4789,In_1859);
or U217 (N_217,In_498,In_2252);
and U218 (N_218,In_3726,In_2737);
nand U219 (N_219,In_3147,In_2565);
nand U220 (N_220,In_2317,In_1739);
or U221 (N_221,In_3008,In_531);
nor U222 (N_222,In_3924,In_3263);
and U223 (N_223,In_3116,In_4934);
nor U224 (N_224,In_533,In_2329);
nand U225 (N_225,In_1080,In_437);
and U226 (N_226,In_1392,In_2327);
and U227 (N_227,In_3309,In_4721);
xnor U228 (N_228,In_4137,In_3459);
xnor U229 (N_229,In_3199,In_3783);
nand U230 (N_230,In_306,In_1373);
and U231 (N_231,In_1517,In_4059);
nor U232 (N_232,In_2605,In_4861);
or U233 (N_233,In_1945,In_2169);
or U234 (N_234,In_4012,In_2695);
and U235 (N_235,In_898,In_2069);
nand U236 (N_236,In_897,In_3039);
nand U237 (N_237,In_2600,In_3075);
nor U238 (N_238,In_2000,In_4638);
or U239 (N_239,In_157,In_2201);
nor U240 (N_240,In_1694,In_1501);
nor U241 (N_241,In_4113,In_2424);
and U242 (N_242,In_1590,In_1478);
xnor U243 (N_243,In_966,In_3391);
nand U244 (N_244,In_2132,In_2663);
xnor U245 (N_245,In_2335,In_3666);
xnor U246 (N_246,In_4409,In_2902);
nor U247 (N_247,In_996,In_696);
nor U248 (N_248,In_3912,In_2194);
and U249 (N_249,In_4218,In_729);
nor U250 (N_250,In_2475,In_751);
or U251 (N_251,In_2382,In_3713);
and U252 (N_252,In_3664,In_3758);
nor U253 (N_253,In_3734,In_3097);
and U254 (N_254,In_4556,In_2980);
and U255 (N_255,In_1143,In_1819);
or U256 (N_256,In_4839,In_1526);
or U257 (N_257,In_3571,In_3403);
nand U258 (N_258,In_2845,In_4650);
nand U259 (N_259,In_2228,In_2312);
and U260 (N_260,In_395,In_3197);
xnor U261 (N_261,In_4345,In_4837);
nor U262 (N_262,In_2455,In_1941);
or U263 (N_263,In_397,In_3294);
and U264 (N_264,In_3832,In_931);
nor U265 (N_265,In_2204,In_2815);
and U266 (N_266,In_3601,In_2051);
and U267 (N_267,In_1589,In_4994);
nand U268 (N_268,In_390,In_1414);
nand U269 (N_269,In_612,In_4396);
and U270 (N_270,In_3947,In_2904);
xor U271 (N_271,In_4384,In_3207);
nor U272 (N_272,In_1748,In_4797);
nor U273 (N_273,In_3122,In_4622);
or U274 (N_274,In_3668,In_65);
nand U275 (N_275,In_881,In_1316);
nand U276 (N_276,In_3216,In_1781);
xnor U277 (N_277,In_2135,In_633);
xor U278 (N_278,In_972,In_1388);
nor U279 (N_279,In_4583,In_2941);
and U280 (N_280,In_4703,In_1156);
nand U281 (N_281,In_1152,In_4455);
nor U282 (N_282,In_702,In_2757);
nor U283 (N_283,In_4974,In_1721);
xor U284 (N_284,In_3984,In_952);
xnor U285 (N_285,In_1079,In_4748);
or U286 (N_286,In_1651,In_4222);
and U287 (N_287,In_1223,In_3747);
or U288 (N_288,In_3322,In_2693);
xor U289 (N_289,In_2264,In_94);
xor U290 (N_290,In_3646,In_3023);
or U291 (N_291,In_156,In_4448);
nand U292 (N_292,In_3982,In_3066);
nor U293 (N_293,In_4973,In_819);
nor U294 (N_294,In_3755,In_319);
or U295 (N_295,In_3883,In_457);
nand U296 (N_296,In_3901,In_2031);
nor U297 (N_297,In_3176,In_4348);
and U298 (N_298,In_2554,In_1068);
or U299 (N_299,In_2393,In_2174);
xor U300 (N_300,In_4689,In_4720);
nand U301 (N_301,In_4037,In_710);
nand U302 (N_302,In_1007,In_211);
or U303 (N_303,In_3740,In_1818);
or U304 (N_304,In_2951,In_3743);
nand U305 (N_305,In_2416,In_1640);
or U306 (N_306,In_1637,In_554);
or U307 (N_307,In_1216,In_4678);
nand U308 (N_308,In_641,In_1039);
nand U309 (N_309,In_2241,In_1249);
and U310 (N_310,In_1736,In_4584);
and U311 (N_311,In_970,In_2570);
nand U312 (N_312,In_1283,In_3663);
and U313 (N_313,In_1598,In_254);
or U314 (N_314,In_225,In_3840);
nor U315 (N_315,In_4596,In_3665);
nand U316 (N_316,In_1755,In_409);
and U317 (N_317,In_474,In_1831);
or U318 (N_318,In_272,In_4889);
nor U319 (N_319,In_4353,In_2267);
xnor U320 (N_320,In_4461,In_2648);
or U321 (N_321,In_834,In_3815);
nor U322 (N_322,In_246,In_185);
nand U323 (N_323,In_3316,In_2481);
and U324 (N_324,In_1451,In_1867);
nor U325 (N_325,In_3146,In_2721);
nand U326 (N_326,In_4133,In_2136);
or U327 (N_327,In_3453,In_1557);
nand U328 (N_328,In_1433,In_213);
nor U329 (N_329,In_3491,In_2280);
and U330 (N_330,In_3850,In_2567);
or U331 (N_331,In_2827,In_1632);
or U332 (N_332,In_1038,In_4762);
and U333 (N_333,In_663,In_4235);
xor U334 (N_334,In_4368,In_828);
and U335 (N_335,In_3818,In_1827);
or U336 (N_336,In_3962,In_289);
xnor U337 (N_337,In_4243,In_1398);
nand U338 (N_338,In_4315,In_817);
or U339 (N_339,In_2831,In_3841);
nor U340 (N_340,In_170,In_914);
and U341 (N_341,In_4582,In_1826);
nand U342 (N_342,In_1026,In_3024);
or U343 (N_343,In_1276,In_2630);
or U344 (N_344,In_3318,In_988);
and U345 (N_345,In_3510,In_2701);
nand U346 (N_346,In_1485,In_1486);
or U347 (N_347,In_308,In_3178);
or U348 (N_348,In_212,In_1413);
nand U349 (N_349,In_1706,In_3863);
xor U350 (N_350,In_89,In_19);
nor U351 (N_351,In_1545,In_1617);
nand U352 (N_352,In_173,In_451);
or U353 (N_353,In_1462,In_3218);
nand U354 (N_354,In_2836,In_1298);
xor U355 (N_355,In_3560,In_787);
and U356 (N_356,In_4034,In_587);
nor U357 (N_357,In_3191,In_327);
and U358 (N_358,In_2388,In_1278);
nand U359 (N_359,In_2283,In_1855);
nand U360 (N_360,In_4646,In_341);
nand U361 (N_361,In_3684,In_3654);
and U362 (N_362,In_4238,In_1943);
nor U363 (N_363,In_3152,In_2710);
nand U364 (N_364,In_1208,In_896);
nand U365 (N_365,In_2661,In_1875);
xor U366 (N_366,In_2788,In_323);
and U367 (N_367,In_2549,In_1286);
nor U368 (N_368,In_1348,In_3082);
and U369 (N_369,In_4444,In_3241);
nor U370 (N_370,In_39,In_1005);
nand U371 (N_371,In_542,In_2900);
and U372 (N_372,In_2656,In_1889);
or U373 (N_373,In_1375,In_4358);
nor U374 (N_374,In_3535,In_1937);
nor U375 (N_375,In_2527,In_260);
and U376 (N_376,In_4203,In_648);
and U377 (N_377,In_2574,In_2358);
nor U378 (N_378,In_1444,In_2994);
nand U379 (N_379,In_35,In_4744);
nand U380 (N_380,In_785,In_1473);
or U381 (N_381,In_2880,In_3160);
and U382 (N_382,In_1307,In_2311);
and U383 (N_383,In_112,In_1207);
nor U384 (N_384,In_2176,In_1652);
nand U385 (N_385,In_2676,In_2363);
nor U386 (N_386,In_577,In_4385);
nand U387 (N_387,In_2506,In_4408);
or U388 (N_388,In_1484,In_1385);
xor U389 (N_389,In_2961,In_3488);
nor U390 (N_390,In_1508,In_4100);
or U391 (N_391,In_3745,In_1476);
and U392 (N_392,In_1422,In_2866);
nand U393 (N_393,In_4266,In_2453);
xor U394 (N_394,In_1034,In_3764);
nor U395 (N_395,In_1423,In_3078);
xnor U396 (N_396,In_1577,In_3073);
nor U397 (N_397,In_1582,In_3133);
nand U398 (N_398,In_2551,In_3929);
xor U399 (N_399,In_2458,In_1643);
xor U400 (N_400,In_3868,In_3839);
nor U401 (N_401,In_1733,In_497);
xnor U402 (N_402,In_2181,In_1318);
nor U403 (N_403,In_2532,In_4743);
xnor U404 (N_404,In_2833,In_2723);
and U405 (N_405,In_989,In_471);
nand U406 (N_406,In_175,In_4232);
or U407 (N_407,In_3307,In_2081);
nor U408 (N_408,In_4591,In_4195);
and U409 (N_409,In_3748,In_1287);
nor U410 (N_410,In_1456,In_3940);
xnor U411 (N_411,In_2218,In_4719);
or U412 (N_412,In_3205,In_1655);
nand U413 (N_413,In_1479,In_3157);
xnor U414 (N_414,In_1805,In_448);
nor U415 (N_415,In_3349,In_2501);
xor U416 (N_416,In_4571,In_4182);
and U417 (N_417,In_2503,In_1624);
or U418 (N_418,In_3589,In_1193);
and U419 (N_419,In_4736,In_447);
nand U420 (N_420,In_3972,In_684);
nor U421 (N_421,In_1515,In_4548);
xnor U422 (N_422,In_2525,In_3930);
nor U423 (N_423,In_2921,In_571);
xnor U424 (N_424,In_1842,In_2700);
and U425 (N_425,In_2437,In_723);
or U426 (N_426,In_4286,In_4914);
xor U427 (N_427,In_4658,In_3673);
and U428 (N_428,In_1332,In_1976);
and U429 (N_429,In_776,In_1594);
and U430 (N_430,In_420,In_2300);
nand U431 (N_431,In_2145,In_4771);
nand U432 (N_432,In_1849,In_3188);
nor U433 (N_433,In_1190,In_4826);
or U434 (N_434,In_4654,In_3134);
and U435 (N_435,In_1234,In_1481);
nor U436 (N_436,In_3099,In_1984);
xnor U437 (N_437,In_2923,In_55);
or U438 (N_438,In_1917,In_1903);
nand U439 (N_439,In_4466,In_4766);
nand U440 (N_440,In_3125,In_3136);
nand U441 (N_441,In_721,In_243);
nor U442 (N_442,In_2784,In_567);
nor U443 (N_443,In_1259,In_2680);
nor U444 (N_444,In_3903,In_1722);
and U445 (N_445,In_4880,In_3851);
nor U446 (N_446,In_4311,In_291);
nand U447 (N_447,In_1309,In_4388);
nand U448 (N_448,In_1222,In_4969);
xnor U449 (N_449,In_2578,In_3600);
and U450 (N_450,In_4742,In_4499);
nor U451 (N_451,In_1871,In_2745);
nor U452 (N_452,In_1982,In_2215);
or U453 (N_453,In_830,In_2422);
nor U454 (N_454,In_3132,In_2407);
nand U455 (N_455,In_2150,In_2922);
xnor U456 (N_456,In_3556,In_4874);
nor U457 (N_457,In_1914,In_2861);
nand U458 (N_458,In_1773,In_703);
xnor U459 (N_459,In_3135,In_2334);
nor U460 (N_460,In_779,In_1680);
or U461 (N_461,In_791,In_1200);
nor U462 (N_462,In_204,In_2985);
nor U463 (N_463,In_1681,In_1376);
or U464 (N_464,In_716,In_33);
and U465 (N_465,In_2037,In_3282);
xnor U466 (N_466,In_4044,In_4885);
nand U467 (N_467,In_3150,In_4601);
xor U468 (N_468,In_1608,In_1647);
or U469 (N_469,In_2581,In_1621);
xor U470 (N_470,In_3795,In_910);
nand U471 (N_471,In_2521,In_2679);
nor U472 (N_472,In_604,In_297);
nand U473 (N_473,In_1500,In_3472);
or U474 (N_474,In_359,In_3385);
xor U475 (N_475,In_17,In_2418);
xor U476 (N_476,In_4741,In_506);
nor U477 (N_477,In_4832,In_556);
and U478 (N_478,In_4521,In_1098);
and U479 (N_479,In_1053,In_4132);
xnor U480 (N_480,In_4989,In_455);
nand U481 (N_481,In_230,In_3597);
xor U482 (N_482,In_2874,In_1460);
and U483 (N_483,In_944,In_1185);
and U484 (N_484,In_1499,In_3489);
or U485 (N_485,In_747,In_2911);
or U486 (N_486,In_3029,In_660);
nand U487 (N_487,In_4187,In_2064);
nand U488 (N_488,In_2091,In_2841);
xor U489 (N_489,In_3433,In_3492);
xnor U490 (N_490,In_2259,In_2168);
or U491 (N_491,In_3652,In_4476);
nor U492 (N_492,In_2446,In_4634);
and U493 (N_493,In_1319,In_1534);
nand U494 (N_494,In_2638,In_2017);
xor U495 (N_495,In_1936,In_4715);
xnor U496 (N_496,In_4381,In_2413);
xor U497 (N_497,In_1719,In_2909);
or U498 (N_498,In_610,In_2817);
or U499 (N_499,In_1195,In_1956);
or U500 (N_500,In_975,In_2703);
nor U501 (N_501,In_2310,In_2415);
xnor U502 (N_502,In_4570,In_1784);
nor U503 (N_503,In_4341,In_2706);
nor U504 (N_504,In_4968,In_169);
and U505 (N_505,In_620,In_1772);
nand U506 (N_506,In_3914,In_2497);
nand U507 (N_507,In_2870,In_4810);
xnor U508 (N_508,In_851,In_742);
or U509 (N_509,In_1131,In_1573);
nand U510 (N_510,In_4284,In_3631);
nor U511 (N_511,In_1729,In_4526);
or U512 (N_512,In_4647,In_3381);
nand U513 (N_513,In_1400,In_1654);
or U514 (N_514,In_2166,In_2345);
and U515 (N_515,In_1206,In_4095);
or U516 (N_516,In_786,In_3873);
nand U517 (N_517,In_1220,In_3480);
nand U518 (N_518,In_2561,In_4305);
xor U519 (N_519,In_3774,In_1747);
nand U520 (N_520,In_1100,In_4536);
nand U521 (N_521,In_902,In_1735);
and U522 (N_522,In_871,In_1389);
and U523 (N_523,In_3974,In_3750);
xor U524 (N_524,In_762,In_2743);
and U525 (N_525,In_755,In_1093);
and U526 (N_526,In_2119,In_3816);
or U527 (N_527,In_4316,In_1663);
nor U528 (N_528,In_2480,In_816);
or U529 (N_529,In_1726,In_3490);
nand U530 (N_530,In_4806,In_4847);
and U531 (N_531,In_2083,In_4586);
nand U532 (N_532,In_4419,In_4202);
xnor U533 (N_533,In_2935,In_347);
and U534 (N_534,In_376,In_1058);
and U535 (N_535,In_1255,In_1300);
nor U536 (N_536,In_706,In_1288);
and U537 (N_537,In_1704,In_429);
and U538 (N_538,In_761,In_3336);
xor U539 (N_539,In_2188,In_3421);
nand U540 (N_540,In_369,In_825);
nor U541 (N_541,In_1446,In_4249);
nor U542 (N_542,In_3603,In_1689);
or U543 (N_543,In_1112,In_3723);
nand U544 (N_544,In_3362,In_3757);
or U545 (N_545,In_4605,In_3954);
xnor U546 (N_546,In_678,In_158);
nand U547 (N_547,In_3957,In_1983);
xor U548 (N_548,In_1553,In_3293);
nor U549 (N_549,In_1133,In_789);
nand U550 (N_550,In_2603,In_595);
nor U551 (N_551,In_419,In_3255);
nor U552 (N_552,In_3215,In_4824);
or U553 (N_553,In_1971,In_2629);
nand U554 (N_554,In_2301,In_2485);
nor U555 (N_555,In_2212,In_2697);
or U556 (N_556,In_3956,In_608);
or U557 (N_557,In_3028,In_3301);
nor U558 (N_558,In_4066,In_1595);
nor U559 (N_559,In_752,In_4857);
nor U560 (N_560,In_3773,In_4713);
xnor U561 (N_561,In_1843,In_1852);
and U562 (N_562,In_4105,In_2976);
or U563 (N_563,In_463,In_1587);
xor U564 (N_564,In_3159,In_4517);
xnor U565 (N_565,In_3413,In_4062);
nor U566 (N_566,In_2498,In_302);
and U567 (N_567,In_1212,In_1674);
xnor U568 (N_568,In_3281,In_1380);
or U569 (N_569,In_1554,In_4791);
or U570 (N_570,In_1641,In_4094);
nand U571 (N_571,In_3944,In_1676);
nor U572 (N_572,In_739,In_284);
or U573 (N_573,In_1750,In_2942);
nand U574 (N_574,In_4942,In_3074);
nand U575 (N_575,In_1312,In_1325);
or U576 (N_576,In_2190,In_1353);
xor U577 (N_577,In_1138,In_1087);
and U578 (N_578,In_2184,In_434);
and U579 (N_579,In_3708,In_4441);
or U580 (N_580,In_2859,In_3093);
and U581 (N_581,In_1104,In_3055);
nand U582 (N_582,In_2820,In_673);
xor U583 (N_583,In_1242,In_338);
and U584 (N_584,In_2026,In_708);
xor U585 (N_585,In_1110,In_4423);
and U586 (N_586,In_924,In_1001);
xnor U587 (N_587,In_1196,In_2061);
or U588 (N_588,In_4071,In_2107);
nor U589 (N_589,In_3615,In_1987);
or U590 (N_590,In_4082,In_3657);
nand U591 (N_591,In_80,In_4056);
nor U592 (N_592,In_1448,In_2199);
or U593 (N_593,In_1666,In_4878);
nand U594 (N_594,In_4558,In_176);
or U595 (N_595,In_4267,In_4282);
and U596 (N_596,In_4852,In_2540);
nand U597 (N_597,In_2777,In_1108);
and U598 (N_598,In_4722,In_4020);
nor U599 (N_599,In_1292,In_2482);
and U600 (N_600,In_3813,In_1601);
xnor U601 (N_601,In_1365,In_1256);
nand U602 (N_602,In_4515,In_1857);
and U603 (N_603,In_730,In_3447);
and U604 (N_604,In_2553,In_1802);
nor U605 (N_605,In_4581,In_3401);
nand U606 (N_606,In_720,In_1134);
and U607 (N_607,In_2552,In_1331);
or U608 (N_608,In_3539,In_2034);
or U609 (N_609,In_735,In_3314);
or U610 (N_610,In_2637,In_4633);
nor U611 (N_611,In_4568,In_2617);
nand U612 (N_612,In_135,In_674);
xor U613 (N_613,In_4733,In_1544);
or U614 (N_614,In_2869,In_1291);
and U615 (N_615,In_1497,In_3769);
and U616 (N_616,In_3925,In_4783);
nor U617 (N_617,In_4888,In_4687);
nor U618 (N_618,In_2763,In_4840);
xnor U619 (N_619,In_922,In_2056);
nand U620 (N_620,In_1345,In_4420);
nor U621 (N_621,In_355,In_2960);
xnor U622 (N_622,In_4808,In_553);
nor U623 (N_623,In_4925,In_4322);
and U624 (N_624,In_3735,In_4490);
xnor U625 (N_625,In_3044,In_1329);
nand U626 (N_626,In_888,In_2950);
nor U627 (N_627,In_596,In_3430);
nor U628 (N_628,In_856,In_1743);
nand U629 (N_629,In_3194,In_99);
nor U630 (N_630,In_3627,In_3346);
xnor U631 (N_631,In_4323,In_3467);
and U632 (N_632,In_4519,In_1645);
and U633 (N_633,In_593,In_3257);
nor U634 (N_634,In_4225,In_1020);
xnor U635 (N_635,In_3373,In_478);
nor U636 (N_636,In_4356,In_491);
and U637 (N_637,In_1044,In_4916);
and U638 (N_638,In_316,In_412);
xnor U639 (N_639,In_295,In_1519);
or U640 (N_640,In_2005,In_2893);
or U641 (N_641,In_2940,In_4002);
and U642 (N_642,In_208,In_3874);
and U643 (N_643,In_160,In_3766);
nand U644 (N_644,In_1358,In_4127);
nor U645 (N_645,In_628,In_3425);
xnor U646 (N_646,In_4097,In_2423);
xor U647 (N_647,In_4049,In_479);
xnor U648 (N_648,In_4780,In_1246);
nor U649 (N_649,In_2391,In_1516);
nand U650 (N_650,In_4990,In_3949);
or U651 (N_651,In_150,In_381);
nor U652 (N_652,In_642,In_1445);
and U653 (N_653,In_2126,In_3588);
nor U654 (N_654,In_1191,In_261);
nand U655 (N_655,In_339,In_36);
nor U656 (N_656,In_1565,In_481);
or U657 (N_657,In_3378,In_380);
nand U658 (N_658,In_4923,In_1551);
and U659 (N_659,In_288,In_2782);
and U660 (N_660,In_389,In_808);
or U661 (N_661,In_4188,In_2479);
nor U662 (N_662,In_2813,In_2115);
xor U663 (N_663,In_2427,In_3561);
nand U664 (N_664,In_426,In_3681);
xnor U665 (N_665,In_647,In_1107);
nor U666 (N_666,In_2908,In_3173);
nand U667 (N_667,In_1861,In_4055);
or U668 (N_668,In_1043,In_4480);
nand U669 (N_669,In_3405,In_446);
nand U670 (N_670,In_1631,In_806);
or U671 (N_671,In_651,In_3432);
nor U672 (N_672,In_859,In_726);
nand U673 (N_673,In_1838,In_2767);
xnor U674 (N_674,In_2308,In_2125);
nand U675 (N_675,In_1092,In_590);
xor U676 (N_676,In_2798,In_2205);
or U677 (N_677,In_2038,In_1763);
nor U678 (N_678,In_2948,In_2463);
nand U679 (N_679,In_4179,In_232);
or U680 (N_680,In_2538,In_2863);
nand U681 (N_681,In_1986,In_1744);
and U682 (N_682,In_4668,In_456);
nor U683 (N_683,In_2573,In_1542);
nand U684 (N_684,In_3151,In_9);
nor U685 (N_685,In_987,In_97);
or U686 (N_686,In_360,In_650);
and U687 (N_687,In_2343,In_2938);
and U688 (N_688,In_1041,In_1700);
or U689 (N_689,In_1071,In_3179);
or U690 (N_690,In_3350,In_1785);
and U691 (N_691,In_909,In_3808);
or U692 (N_692,In_1095,In_1741);
nand U693 (N_693,In_4590,In_4924);
nor U694 (N_694,In_20,In_2392);
or U695 (N_695,In_403,In_2794);
nor U696 (N_696,In_4228,In_2588);
nand U697 (N_697,In_1673,In_2672);
nor U698 (N_698,In_3760,In_956);
nor U699 (N_699,In_2725,In_1503);
or U700 (N_700,In_4706,In_4196);
nand U701 (N_701,In_274,In_892);
nor U702 (N_702,In_4010,In_3827);
nand U703 (N_703,In_188,In_1873);
xnor U704 (N_704,In_3619,In_2500);
and U705 (N_705,In_3983,In_3476);
nor U706 (N_706,In_4993,In_1257);
xor U707 (N_707,In_4233,In_3035);
nand U708 (N_708,In_4000,In_714);
nand U709 (N_709,In_4177,In_2696);
nand U710 (N_710,In_4427,In_3308);
or U711 (N_711,In_1429,In_42);
xnor U712 (N_712,In_3801,In_4024);
and U713 (N_713,In_3584,In_3742);
nand U714 (N_714,In_4851,In_1066);
nor U715 (N_715,In_4624,In_3123);
or U716 (N_716,In_2175,In_1140);
nand U717 (N_717,In_1779,In_893);
xnor U718 (N_718,In_672,In_4531);
or U719 (N_719,In_1746,In_3071);
xnor U720 (N_720,In_4777,In_2473);
nand U721 (N_721,In_3198,In_4304);
nor U722 (N_722,In_1417,In_659);
or U723 (N_723,In_2726,In_340);
nor U724 (N_724,In_4675,In_3183);
nor U725 (N_725,In_404,In_1884);
or U726 (N_726,In_712,In_4752);
or U727 (N_727,In_1684,In_1203);
xor U728 (N_728,In_1821,In_813);
or U729 (N_729,In_1713,In_4985);
nor U730 (N_730,In_3809,In_3805);
or U731 (N_731,In_4843,In_2624);
or U732 (N_732,In_526,In_698);
nor U733 (N_733,In_4952,In_3047);
xnor U734 (N_734,In_1567,In_2779);
nor U735 (N_735,In_1769,In_1065);
nand U736 (N_736,In_1254,In_2547);
and U737 (N_737,In_1962,In_1841);
or U738 (N_738,In_4522,In_2395);
nand U739 (N_739,In_1111,In_3254);
and U740 (N_740,In_4165,In_1579);
nand U741 (N_741,In_4520,In_1908);
or U742 (N_742,In_2390,In_130);
nor U743 (N_743,In_1075,In_1031);
and U744 (N_744,In_1931,In_3672);
nor U745 (N_745,In_722,In_3129);
nand U746 (N_746,In_2143,In_4793);
nand U747 (N_747,In_2729,In_4456);
and U748 (N_748,In_1929,In_699);
xnor U749 (N_749,In_2742,In_67);
and U750 (N_750,In_4021,In_95);
and U751 (N_751,In_4183,In_4160);
xor U752 (N_752,In_2635,In_4939);
nand U753 (N_753,In_862,In_1153);
nor U754 (N_754,In_1443,In_217);
or U755 (N_755,In_78,In_3048);
nand U756 (N_756,In_3557,In_3269);
nor U757 (N_757,In_3495,In_1607);
or U758 (N_758,In_4630,In_1707);
or U759 (N_759,In_833,In_697);
nor U760 (N_760,In_1797,In_4869);
nand U761 (N_761,In_3162,In_1290);
nand U762 (N_762,In_3608,In_259);
nor U763 (N_763,In_1630,In_3083);
nand U764 (N_764,In_3352,In_982);
nor U765 (N_765,In_3153,In_4898);
nand U766 (N_766,In_6,In_181);
or U767 (N_767,In_2326,In_3860);
or U768 (N_768,In_1170,In_1176);
xor U769 (N_769,In_1528,In_2339);
and U770 (N_770,In_753,In_4121);
nor U771 (N_771,In_3498,In_343);
or U772 (N_772,In_4716,In_4438);
xnor U773 (N_773,In_3806,In_2214);
nand U774 (N_774,In_2594,In_4162);
nand U775 (N_775,In_344,In_1454);
or U776 (N_776,In_2786,In_1960);
and U777 (N_777,In_4158,In_4655);
nor U778 (N_778,In_3004,In_1656);
nand U779 (N_779,In_1771,In_624);
and U780 (N_780,In_1116,In_3899);
nor U781 (N_781,In_192,In_1866);
and U782 (N_782,In_417,In_1399);
nand U783 (N_783,In_2469,In_4468);
nand U784 (N_784,In_2072,In_4439);
nor U785 (N_785,In_3234,In_72);
nor U786 (N_786,In_3921,In_2454);
nand U787 (N_787,In_387,In_4332);
or U788 (N_788,In_740,In_4317);
nor U789 (N_789,In_2077,In_1959);
nand U790 (N_790,In_788,In_990);
or U791 (N_791,In_422,In_958);
or U792 (N_792,In_1117,In_3388);
nand U793 (N_793,In_4140,In_4610);
nand U794 (N_794,In_2387,In_4126);
or U795 (N_795,In_1421,In_2616);
nor U796 (N_796,In_921,In_1425);
xor U797 (N_797,In_3525,In_4701);
nor U798 (N_798,In_4541,In_1390);
nor U799 (N_799,In_1099,In_4792);
nor U800 (N_800,In_1437,In_1754);
nor U801 (N_801,In_3455,In_2585);
or U802 (N_802,In_4064,In_3507);
xnor U803 (N_803,In_523,In_1245);
and U804 (N_804,In_760,In_873);
xor U805 (N_805,In_563,In_1878);
and U806 (N_806,In_2253,In_2067);
nand U807 (N_807,In_1727,In_290);
nand U808 (N_808,In_4616,In_256);
and U809 (N_809,In_3310,In_504);
or U810 (N_810,In_1097,In_600);
and U811 (N_811,In_4485,In_3274);
or U812 (N_812,In_4296,In_1506);
and U813 (N_813,In_4918,In_4046);
nor U814 (N_814,In_913,In_4672);
xnor U815 (N_815,In_4301,In_3640);
nor U816 (N_816,In_2523,In_96);
nand U817 (N_817,In_2677,In_163);
or U818 (N_818,In_1770,In_320);
and U819 (N_819,In_3598,In_992);
xnor U820 (N_820,In_1252,In_4953);
or U821 (N_821,In_3323,In_4546);
or U822 (N_822,In_3232,In_3283);
nand U823 (N_823,In_4904,In_2250);
nand U824 (N_824,In_3370,In_2198);
nand U825 (N_825,In_2292,In_4735);
xor U826 (N_826,In_732,In_1820);
or U827 (N_827,In_1606,In_3823);
and U828 (N_828,In_3669,In_4504);
xor U829 (N_829,In_3728,In_1402);
xnor U830 (N_830,In_3612,In_1083);
and U831 (N_831,In_4343,In_2946);
nand U832 (N_832,In_1811,In_1535);
nand U833 (N_833,In_4050,In_594);
nor U834 (N_834,In_2318,In_4606);
and U835 (N_835,In_904,In_1301);
and U836 (N_836,In_2973,In_44);
xor U837 (N_837,In_3375,In_52);
nand U838 (N_838,In_3275,In_3862);
nand U839 (N_839,In_2494,In_4730);
xnor U840 (N_840,In_3756,In_3389);
nand U841 (N_841,In_4352,In_2699);
and U842 (N_842,In_4329,In_168);
nand U843 (N_843,In_2257,In_3704);
xor U844 (N_844,In_3596,In_4155);
nand U845 (N_845,In_4859,In_3006);
or U846 (N_846,In_3888,In_2749);
nand U847 (N_847,In_4469,In_4143);
nand U848 (N_848,In_4754,In_2442);
or U849 (N_849,In_138,In_1753);
xnor U850 (N_850,In_4492,In_3102);
xor U851 (N_851,In_4751,In_1991);
or U852 (N_852,In_1715,In_3233);
or U853 (N_853,In_3973,In_3379);
and U854 (N_854,In_3670,In_3021);
nor U855 (N_855,In_4554,In_3092);
nand U856 (N_856,In_2007,In_4333);
nor U857 (N_857,In_4288,In_2373);
nor U858 (N_858,In_1675,In_113);
nor U859 (N_859,In_548,In_4507);
and U860 (N_860,In_3923,In_875);
or U861 (N_861,In_2111,In_1395);
nand U862 (N_862,In_3208,In_1055);
or U863 (N_863,In_4390,In_2071);
and U864 (N_864,In_3541,In_1161);
or U865 (N_865,In_1586,In_4908);
nor U866 (N_866,In_4845,In_1045);
nor U867 (N_867,In_3120,In_3812);
or U868 (N_868,In_3068,In_2242);
xnor U869 (N_869,In_4148,In_3204);
nand U870 (N_870,In_425,In_2736);
nand U871 (N_871,In_573,In_853);
xnor U872 (N_872,In_438,In_3877);
xnor U873 (N_873,In_4131,In_1469);
and U874 (N_874,In_4933,In_3468);
and U875 (N_875,In_3732,In_1299);
xnor U876 (N_876,In_458,In_2968);
or U877 (N_877,In_4769,In_911);
nor U878 (N_878,In_1980,In_2741);
and U879 (N_879,In_950,In_3887);
xor U880 (N_880,In_1150,In_2152);
xor U881 (N_881,In_3849,In_693);
or U882 (N_882,In_1239,In_4803);
xnor U883 (N_883,In_2847,In_3916);
nor U884 (N_884,In_4940,In_4178);
nor U885 (N_885,In_475,In_4481);
xnor U886 (N_886,In_2967,In_1856);
xnor U887 (N_887,In_4136,In_182);
xor U888 (N_888,In_1447,In_3229);
or U889 (N_889,In_4452,In_2740);
xor U890 (N_890,In_4173,In_570);
nor U891 (N_891,In_3287,In_1480);
and U892 (N_892,In_700,In_62);
and U893 (N_893,In_2773,In_2229);
xnor U894 (N_894,In_489,In_4821);
xnor U895 (N_895,In_3449,In_4068);
xor U896 (N_896,In_649,In_948);
xnor U897 (N_897,In_2901,In_4216);
nor U898 (N_898,In_2094,In_1916);
nand U899 (N_899,In_103,In_3342);
and U900 (N_900,In_1243,In_736);
nand U901 (N_901,In_3679,In_741);
or U902 (N_902,In_2796,In_2575);
nor U903 (N_903,In_2457,In_349);
nand U904 (N_904,In_315,In_3678);
nand U905 (N_905,In_3088,In_1870);
nor U906 (N_906,In_3580,In_1279);
xor U907 (N_907,In_4346,In_2088);
and U908 (N_908,In_782,In_3653);
nand U909 (N_909,In_1211,In_4578);
xnor U910 (N_910,In_4280,In_622);
and U911 (N_911,In_365,In_472);
nand U912 (N_912,In_4892,In_3288);
or U913 (N_913,In_4479,In_3211);
nor U914 (N_914,In_3206,In_4367);
and U915 (N_915,In_1450,In_1409);
and U916 (N_916,In_3969,In_2104);
or U917 (N_917,In_724,In_882);
nor U918 (N_918,In_3611,In_3909);
or U919 (N_919,In_2456,In_938);
nor U920 (N_920,In_4128,In_1578);
nor U921 (N_921,In_3651,In_1209);
or U922 (N_922,In_92,In_4260);
nand U923 (N_923,In_1284,In_1004);
xnor U924 (N_924,In_2160,In_4328);
xnor U925 (N_925,In_14,In_655);
and U926 (N_926,In_4897,In_1258);
and U927 (N_927,In_1961,In_4081);
and U928 (N_928,In_3484,In_309);
and U929 (N_929,In_4798,In_2436);
xnor U930 (N_930,In_4391,In_546);
nor U931 (N_931,In_1240,In_268);
and U932 (N_932,In_4524,In_3238);
nand U933 (N_933,In_4248,In_4159);
or U934 (N_934,In_1662,In_4598);
nand U935 (N_935,In_4911,In_3680);
or U936 (N_936,In_1701,In_4324);
or U937 (N_937,In_947,In_4489);
nand U938 (N_938,In_1397,In_214);
and U939 (N_939,In_623,In_1762);
and U940 (N_940,In_2360,In_1619);
nor U941 (N_941,In_631,In_3546);
xor U942 (N_942,In_1714,In_3649);
nand U943 (N_943,In_2516,In_2402);
nand U944 (N_944,In_4413,In_1854);
nor U945 (N_945,In_832,In_4253);
and U946 (N_946,In_1471,In_3910);
nor U947 (N_947,In_2370,In_4516);
nor U948 (N_948,In_2421,In_1812);
and U949 (N_949,In_3416,In_1540);
and U950 (N_950,In_1297,In_609);
or U951 (N_951,In_483,In_1434);
xnor U952 (N_952,In_3941,In_4318);
and U953 (N_953,In_0,In_2643);
or U954 (N_954,In_3276,In_1507);
xor U955 (N_955,In_1988,In_4838);
and U956 (N_956,In_3744,In_2599);
and U957 (N_957,In_3508,In_2556);
and U958 (N_958,In_4255,In_4307);
nand U959 (N_959,In_1386,In_3701);
and U960 (N_960,In_2758,In_1896);
nand U961 (N_961,In_3977,In_4740);
nor U962 (N_962,In_410,In_4096);
and U963 (N_963,In_3717,In_3196);
xor U964 (N_964,In_2274,In_1756);
nand U965 (N_965,In_3542,In_4431);
nor U966 (N_966,In_4417,In_3248);
xor U967 (N_967,In_3699,In_2730);
xnor U968 (N_968,In_863,In_3486);
or U969 (N_969,In_4001,In_1546);
nand U970 (N_970,In_3780,In_2349);
xnor U971 (N_971,In_4572,In_2450);
and U972 (N_972,In_2183,In_1649);
and U973 (N_973,In_1267,In_2571);
xnor U974 (N_974,In_1558,In_4913);
or U975 (N_975,In_2849,In_1218);
nor U976 (N_976,In_928,In_1474);
nor U977 (N_977,In_1648,In_2844);
xnor U978 (N_978,In_1767,In_2419);
or U979 (N_979,In_2112,In_3145);
xor U980 (N_980,In_4903,In_775);
nand U981 (N_981,In_1151,In_2688);
or U982 (N_982,In_1691,In_4835);
xor U983 (N_983,In_3478,In_1804);
nor U984 (N_984,In_2082,In_4960);
nor U985 (N_985,In_267,In_4950);
and U986 (N_986,In_3847,In_2230);
or U987 (N_987,In_1149,In_3235);
and U988 (N_988,In_3797,In_591);
nand U989 (N_989,In_4707,In_1817);
or U990 (N_990,In_2364,In_3437);
or U991 (N_991,In_2073,In_1470);
and U992 (N_992,In_4070,In_4252);
or U993 (N_993,In_2853,In_558);
xnor U994 (N_994,In_4135,In_424);
xnor U995 (N_995,In_101,In_2202);
and U996 (N_996,In_317,In_1947);
nor U997 (N_997,In_4593,In_3616);
nand U998 (N_998,In_2876,In_2712);
nor U999 (N_999,In_3623,In_4380);
or U1000 (N_1000,In_3647,In_1074);
and U1001 (N_1001,N_66,In_1814);
xor U1002 (N_1002,In_3754,In_4970);
and U1003 (N_1003,In_3955,In_4313);
or U1004 (N_1004,In_1604,In_71);
nor U1005 (N_1005,N_141,In_768);
nand U1006 (N_1006,In_1795,In_3996);
xor U1007 (N_1007,In_4779,In_1505);
and U1008 (N_1008,In_234,In_2486);
or U1009 (N_1009,In_3593,N_196);
nand U1010 (N_1010,N_558,In_4979);
or U1011 (N_1011,In_1186,In_3650);
nor U1012 (N_1012,In_469,In_3463);
xnor U1013 (N_1013,In_124,N_618);
nor U1014 (N_1014,N_518,In_557);
xor U1015 (N_1015,N_836,N_56);
and U1016 (N_1016,In_842,In_2338);
and U1017 (N_1017,In_1342,N_864);
xnor U1018 (N_1018,In_3299,In_3749);
xor U1019 (N_1019,In_2792,N_432);
nor U1020 (N_1020,In_4723,In_2261);
or U1021 (N_1021,In_3465,In_1603);
and U1022 (N_1022,N_326,In_4146);
and U1023 (N_1023,In_1184,N_692);
xor U1024 (N_1024,N_611,In_487);
nor U1025 (N_1025,In_1269,N_482);
and U1026 (N_1026,N_505,In_2717);
nor U1027 (N_1027,In_4210,In_1761);
nand U1028 (N_1028,In_4366,In_3648);
and U1029 (N_1029,In_2033,In_1052);
nand U1030 (N_1030,In_4542,In_467);
or U1031 (N_1031,N_148,In_1644);
and U1032 (N_1032,N_718,In_939);
xnor U1033 (N_1033,In_2914,In_1146);
xnor U1034 (N_1034,In_4256,In_3724);
nor U1035 (N_1035,N_435,In_4415);
nand U1036 (N_1036,In_508,In_4161);
nor U1037 (N_1037,In_3474,In_4436);
nor U1038 (N_1038,N_925,In_528);
nand U1039 (N_1039,In_4951,N_295);
nor U1040 (N_1040,In_3419,In_1268);
xnor U1041 (N_1041,In_2101,In_3493);
and U1042 (N_1042,In_2917,N_194);
nor U1043 (N_1043,In_197,In_1786);
xnor U1044 (N_1044,N_761,In_1349);
nor U1045 (N_1045,In_1303,In_2671);
or U1046 (N_1046,N_341,In_304);
nand U1047 (N_1047,N_468,In_2276);
nand U1048 (N_1048,In_3810,In_4931);
nor U1049 (N_1049,N_225,In_757);
xor U1050 (N_1050,In_4123,N_690);
xnor U1051 (N_1051,In_976,In_1096);
nand U1052 (N_1052,In_4312,N_990);
and U1053 (N_1053,In_4917,In_4809);
nor U1054 (N_1054,In_3250,N_300);
or U1055 (N_1055,In_1967,In_4434);
nor U1056 (N_1056,N_856,In_4764);
nand U1057 (N_1057,In_275,In_2888);
nor U1058 (N_1058,N_731,In_3264);
nor U1059 (N_1059,In_231,In_1070);
and U1060 (N_1060,N_830,In_249);
xor U1061 (N_1061,In_1027,In_4245);
or U1062 (N_1062,In_1803,N_70);
xnor U1063 (N_1063,In_2040,N_60);
nand U1064 (N_1064,N_844,In_4755);
nand U1065 (N_1065,N_985,In_492);
or U1066 (N_1066,In_428,In_271);
nor U1067 (N_1067,In_1024,In_1369);
and U1068 (N_1068,In_206,In_3483);
xnor U1069 (N_1069,In_4310,N_269);
and U1070 (N_1070,In_2114,In_820);
or U1071 (N_1071,In_4661,In_2240);
and U1072 (N_1072,N_255,In_4948);
nor U1073 (N_1073,In_1688,In_3261);
nor U1074 (N_1074,In_2496,N_799);
nor U1075 (N_1075,In_2593,N_358);
xor U1076 (N_1076,In_1035,In_2381);
or U1077 (N_1077,In_3575,N_414);
or U1078 (N_1078,In_1121,N_397);
or U1079 (N_1079,In_569,In_405);
or U1080 (N_1080,In_3552,In_1089);
or U1081 (N_1081,In_353,In_2766);
xor U1082 (N_1082,In_4275,In_1106);
and U1083 (N_1083,In_482,In_4747);
or U1084 (N_1084,In_2019,In_929);
xnor U1085 (N_1085,In_3165,In_2582);
nand U1086 (N_1086,N_521,In_4254);
nand U1087 (N_1087,In_476,In_3270);
and U1088 (N_1088,N_510,N_697);
nor U1089 (N_1089,N_699,In_901);
nand U1090 (N_1090,N_224,In_1697);
nor U1091 (N_1091,In_4446,N_152);
or U1092 (N_1092,In_2002,In_2271);
or U1093 (N_1093,In_1782,In_1530);
xor U1094 (N_1094,In_4965,In_846);
and U1095 (N_1095,In_452,In_1572);
nor U1096 (N_1096,In_4125,In_3829);
nand U1097 (N_1097,In_2864,In_4980);
xnor U1098 (N_1098,In_4820,In_1541);
or U1099 (N_1099,In_665,In_2238);
xor U1100 (N_1100,In_3020,In_894);
nor U1101 (N_1101,In_4620,In_3927);
xor U1102 (N_1102,In_979,In_1830);
nand U1103 (N_1103,In_1457,In_2780);
nand U1104 (N_1104,In_4404,In_4961);
xnor U1105 (N_1105,In_224,In_3700);
nor U1106 (N_1106,N_956,In_1682);
or U1107 (N_1107,In_707,In_3671);
xnor U1108 (N_1108,In_1514,In_818);
xor U1109 (N_1109,In_3607,N_606);
and U1110 (N_1110,In_3707,In_4022);
nand U1111 (N_1111,In_1521,In_4429);
nand U1112 (N_1112,In_4116,In_4398);
xnor U1113 (N_1113,In_4209,In_3784);
nand U1114 (N_1114,In_1759,In_1328);
and U1115 (N_1115,In_743,In_615);
nand U1116 (N_1116,In_4362,In_3473);
or U1117 (N_1117,N_166,N_987);
nor U1118 (N_1118,In_3168,In_159);
xor U1119 (N_1119,In_1274,In_3900);
nor U1120 (N_1120,In_2664,N_444);
nor U1121 (N_1121,In_3915,N_461);
or U1122 (N_1122,In_2323,N_979);
and U1123 (N_1123,In_731,In_2386);
or U1124 (N_1124,N_794,N_156);
nor U1125 (N_1125,In_4091,N_639);
or U1126 (N_1126,In_4691,N_913);
and U1127 (N_1127,In_4608,N_620);
and U1128 (N_1128,In_379,In_109);
or U1129 (N_1129,In_4184,In_2622);
nor U1130 (N_1130,N_455,N_945);
xor U1131 (N_1131,In_4812,In_3920);
xor U1132 (N_1132,In_4663,N_471);
and U1133 (N_1133,In_210,In_3986);
or U1134 (N_1134,N_952,In_1549);
or U1135 (N_1135,In_2014,N_737);
nor U1136 (N_1136,In_3487,In_149);
nor U1137 (N_1137,In_2210,In_3807);
nor U1138 (N_1138,In_2225,N_357);
xor U1139 (N_1139,In_2598,In_1665);
nor U1140 (N_1140,N_874,In_2895);
nand U1141 (N_1141,In_3943,In_621);
nand U1142 (N_1142,In_3554,In_263);
xnor U1143 (N_1143,N_745,N_299);
or U1144 (N_1144,In_4440,N_212);
nand U1145 (N_1145,N_450,In_602);
nand U1146 (N_1146,In_4023,In_3002);
xor U1147 (N_1147,In_1895,N_105);
nor U1148 (N_1148,In_484,In_3154);
nand U1149 (N_1149,In_1791,N_429);
and U1150 (N_1150,In_550,In_2816);
xnor U1151 (N_1151,In_3770,N_719);
or U1152 (N_1152,In_3803,In_4180);
nor U1153 (N_1153,In_2192,In_4045);
and U1154 (N_1154,In_1354,In_3242);
nand U1155 (N_1155,In_2842,In_592);
xnor U1156 (N_1156,N_851,In_4959);
and U1157 (N_1157,In_3942,In_280);
or U1158 (N_1158,In_3693,In_2080);
nand U1159 (N_1159,In_998,N_792);
or U1160 (N_1160,In_1686,In_2065);
or U1161 (N_1161,In_1368,In_2167);
xor U1162 (N_1162,In_4462,In_1650);
nor U1163 (N_1163,In_1627,In_277);
or U1164 (N_1164,N_619,In_4864);
or U1165 (N_1165,In_4108,In_4103);
xnor U1166 (N_1166,In_1366,In_108);
xor U1167 (N_1167,In_574,N_680);
and U1168 (N_1168,In_346,In_1048);
and U1169 (N_1169,In_2507,In_2512);
and U1170 (N_1170,N_971,In_104);
nand U1171 (N_1171,In_3718,In_2828);
xnor U1172 (N_1172,In_4592,In_2927);
xnor U1173 (N_1173,N_251,N_642);
nor U1174 (N_1174,In_1261,In_4152);
nand U1175 (N_1175,In_733,In_543);
nor U1176 (N_1176,In_2526,N_806);
xor U1177 (N_1177,In_658,In_1789);
nor U1178 (N_1178,N_716,In_4297);
or U1179 (N_1179,In_3121,In_3602);
nor U1180 (N_1180,N_183,In_4106);
and U1181 (N_1181,N_169,In_18);
nor U1182 (N_1182,In_4731,In_2193);
xor U1183 (N_1183,In_368,In_3457);
nor U1184 (N_1184,In_1461,In_3470);
nor U1185 (N_1185,In_541,In_4799);
and U1186 (N_1186,In_3551,In_3838);
nor U1187 (N_1187,In_4842,In_3332);
nand U1188 (N_1188,In_4763,In_4694);
or U1189 (N_1189,In_3266,In_255);
or U1190 (N_1190,N_858,N_706);
xnor U1191 (N_1191,In_4533,In_358);
or U1192 (N_1192,In_2604,In_12);
or U1193 (N_1193,In_4576,In_4628);
and U1194 (N_1194,N_782,In_3637);
nand U1195 (N_1195,N_968,N_949);
and U1196 (N_1196,In_3882,In_4163);
nand U1197 (N_1197,N_420,In_3219);
or U1198 (N_1198,In_3558,In_4039);
nand U1199 (N_1199,In_2959,In_2544);
nand U1200 (N_1200,In_3360,In_1776);
nor U1201 (N_1201,In_3775,In_4027);
and U1202 (N_1202,In_2887,In_133);
nand U1203 (N_1203,In_2537,N_556);
nand U1204 (N_1204,In_2925,In_1364);
xor U1205 (N_1205,In_2084,In_1494);
xor U1206 (N_1206,In_796,In_2835);
xnor U1207 (N_1207,N_770,N_648);
nand U1208 (N_1208,N_74,In_2356);
and U1209 (N_1209,In_2499,In_1102);
nor U1210 (N_1210,In_3771,In_2118);
xnor U1211 (N_1211,N_986,In_3469);
xnor U1212 (N_1212,In_2385,In_3072);
xnor U1213 (N_1213,N_17,In_161);
or U1214 (N_1214,In_4725,In_3497);
nand U1215 (N_1215,In_503,N_386);
nor U1216 (N_1216,In_4003,In_3110);
and U1217 (N_1217,In_2711,N_131);
nand U1218 (N_1218,In_3913,In_2678);
and U1219 (N_1219,N_139,N_602);
nand U1220 (N_1220,In_3865,In_1696);
xnor U1221 (N_1221,In_709,In_4299);
xor U1222 (N_1222,In_1888,N_531);
nand U1223 (N_1223,In_1539,In_1934);
and U1224 (N_1224,In_519,In_1592);
nor U1225 (N_1225,N_629,In_3848);
or U1226 (N_1226,In_2649,In_4349);
nor U1227 (N_1227,In_48,In_3200);
nand U1228 (N_1228,In_1213,N_264);
xor U1229 (N_1229,In_3052,N_304);
xnor U1230 (N_1230,In_4501,In_430);
and U1231 (N_1231,In_1845,N_94);
nand U1232 (N_1232,In_3434,In_848);
nor U1233 (N_1233,N_523,N_587);
nand U1234 (N_1234,In_4251,In_4319);
nand U1235 (N_1235,N_434,In_171);
nand U1236 (N_1236,In_614,In_4320);
nor U1237 (N_1237,In_1938,In_310);
nand U1238 (N_1238,In_2995,N_286);
nor U1239 (N_1239,N_490,N_624);
nor U1240 (N_1240,In_4909,In_2012);
xor U1241 (N_1241,In_2131,In_2203);
or U1242 (N_1242,In_3009,In_179);
and U1243 (N_1243,In_64,In_3635);
or U1244 (N_1244,N_484,N_989);
or U1245 (N_1245,In_1009,In_3785);
or U1246 (N_1246,In_4379,N_265);
xor U1247 (N_1247,In_162,In_3448);
nand U1248 (N_1248,In_1907,N_599);
nor U1249 (N_1249,In_4724,In_1882);
and U1250 (N_1250,N_786,In_919);
xor U1251 (N_1251,In_3644,N_721);
nand U1252 (N_1252,N_134,In_3328);
xnor U1253 (N_1253,In_869,N_702);
or U1254 (N_1254,N_634,In_3239);
and U1255 (N_1255,In_2546,In_3423);
and U1256 (N_1256,In_324,In_3751);
nor U1257 (N_1257,In_3213,In_4921);
or U1258 (N_1258,N_100,In_436);
nand U1259 (N_1259,In_2772,In_4683);
xnor U1260 (N_1260,N_753,In_4901);
xnor U1261 (N_1261,N_938,N_104);
or U1262 (N_1262,N_859,In_3582);
and U1263 (N_1263,N_364,In_1315);
nand U1264 (N_1264,In_2224,In_352);
xor U1265 (N_1265,In_2302,In_2462);
xnor U1266 (N_1266,N_193,N_550);
xnor U1267 (N_1267,In_1262,In_2965);
xor U1268 (N_1268,N_992,N_390);
xnor U1269 (N_1269,In_3137,In_2978);
nand U1270 (N_1270,In_2196,N_958);
or U1271 (N_1271,In_2438,In_3458);
or U1272 (N_1272,In_3417,In_4528);
and U1273 (N_1273,N_34,In_4882);
xnor U1274 (N_1274,N_3,In_3396);
and U1275 (N_1275,N_749,In_131);
nor U1276 (N_1276,N_325,N_542);
and U1277 (N_1277,In_226,In_2324);
xor U1278 (N_1278,In_269,In_2896);
nand U1279 (N_1279,In_1377,N_124);
nand U1280 (N_1280,In_1226,In_3844);
and U1281 (N_1281,In_2219,In_3800);
and U1282 (N_1282,In_2760,In_845);
xnor U1283 (N_1283,In_2134,In_2410);
nand U1284 (N_1284,In_2367,N_919);
nor U1285 (N_1285,In_4261,In_3195);
and U1286 (N_1286,In_8,N_372);
nor U1287 (N_1287,In_1886,In_3361);
nor U1288 (N_1288,In_3063,In_3706);
and U1289 (N_1289,In_3524,In_235);
and U1290 (N_1290,In_3908,In_1751);
or U1291 (N_1291,N_494,In_2046);
xor U1292 (N_1292,In_257,In_229);
nand U1293 (N_1293,In_4784,In_1766);
nor U1294 (N_1294,In_223,In_117);
xor U1295 (N_1295,In_2651,In_367);
and U1296 (N_1296,N_184,N_103);
and U1297 (N_1297,In_314,In_584);
nor U1298 (N_1298,In_2795,N_839);
or U1299 (N_1299,In_24,In_3390);
and U1300 (N_1300,In_3410,In_3353);
and U1301 (N_1301,In_1778,In_2720);
or U1302 (N_1302,N_248,In_1136);
xnor U1303 (N_1303,In_605,In_1248);
and U1304 (N_1304,In_1877,N_873);
xnor U1305 (N_1305,In_715,In_991);
nor U1306 (N_1306,In_2409,In_2389);
nand U1307 (N_1307,In_2857,N_669);
nand U1308 (N_1308,N_149,In_1165);
xor U1309 (N_1309,In_2105,In_1357);
nor U1310 (N_1310,In_4403,N_978);
nor U1311 (N_1311,N_532,In_4250);
or U1312 (N_1312,In_691,In_1396);
and U1313 (N_1313,In_1067,In_4124);
nor U1314 (N_1314,In_1296,In_2732);
nand U1315 (N_1315,In_1737,In_415);
or U1316 (N_1316,In_5,N_24);
or U1317 (N_1317,N_768,In_580);
xor U1318 (N_1318,N_203,In_2865);
xnor U1319 (N_1319,In_382,In_965);
nor U1320 (N_1320,In_3259,N_11);
xor U1321 (N_1321,In_4569,In_4998);
and U1322 (N_1322,In_298,In_69);
xor U1323 (N_1323,In_634,In_1906);
or U1324 (N_1324,In_1851,In_858);
nand U1325 (N_1325,N_22,N_840);
nand U1326 (N_1326,N_464,In_4768);
or U1327 (N_1327,In_3504,N_457);
and U1328 (N_1328,In_2510,In_1334);
xnor U1329 (N_1329,N_182,In_1418);
nand U1330 (N_1330,N_381,In_2275);
and U1331 (N_1331,In_3967,N_557);
or U1332 (N_1332,N_337,In_3609);
nor U1333 (N_1333,In_3705,In_2947);
nor U1334 (N_1334,In_671,In_2180);
nor U1335 (N_1335,N_573,In_719);
and U1336 (N_1336,In_183,N_678);
and U1337 (N_1337,In_758,In_2149);
xnor U1338 (N_1338,In_1823,In_2785);
xor U1339 (N_1339,In_3880,In_2414);
xor U1340 (N_1340,N_356,In_2892);
nand U1341 (N_1341,In_1548,In_3989);
nand U1342 (N_1342,In_1502,In_2823);
or U1343 (N_1343,In_4085,In_607);
and U1344 (N_1344,In_2074,In_485);
and U1345 (N_1345,N_637,In_3174);
and U1346 (N_1346,N_942,In_4643);
or U1347 (N_1347,In_2086,N_15);
or U1348 (N_1348,In_1725,N_76);
nor U1349 (N_1349,In_123,N_379);
nand U1350 (N_1350,N_6,In_216);
and U1351 (N_1351,In_466,In_4274);
xor U1352 (N_1352,N_489,N_388);
nand U1353 (N_1353,N_297,In_962);
xor U1354 (N_1354,In_1731,In_3335);
and U1355 (N_1355,In_3087,In_354);
nand U1356 (N_1356,In_3689,N_69);
nand U1357 (N_1357,In_3431,In_3686);
nand U1358 (N_1358,In_357,In_927);
nor U1359 (N_1359,N_0,N_578);
or U1360 (N_1360,N_694,N_90);
nand U1361 (N_1361,In_1010,N_188);
nor U1362 (N_1362,In_1668,N_422);
nor U1363 (N_1363,In_1868,In_4191);
xor U1364 (N_1364,In_1925,In_3527);
nor U1365 (N_1365,N_628,N_899);
or U1366 (N_1366,N_107,In_2931);
xnor U1367 (N_1367,N_190,N_598);
nand U1368 (N_1368,N_758,In_2130);
nor U1369 (N_1369,N_54,In_87);
or U1370 (N_1370,In_953,In_2408);
xnor U1371 (N_1371,In_2542,N_539);
nor U1372 (N_1372,In_1615,N_983);
or U1373 (N_1373,In_1180,In_860);
or U1374 (N_1374,In_2029,In_1482);
xnor U1375 (N_1375,N_347,In_1757);
and U1376 (N_1376,In_4963,In_1709);
and U1377 (N_1377,In_1238,In_4192);
nor U1378 (N_1378,In_3826,In_3440);
or U1379 (N_1379,In_1881,In_2216);
nand U1380 (N_1380,In_1427,In_2620);
xnor U1381 (N_1381,In_4445,In_414);
and U1382 (N_1382,N_130,N_174);
and U1383 (N_1383,In_2559,In_2615);
or U1384 (N_1384,In_1543,In_4753);
nand U1385 (N_1385,In_530,In_4119);
or U1386 (N_1386,N_389,In_1602);
nand U1387 (N_1387,N_809,In_174);
or U1388 (N_1388,In_4927,In_1042);
xnor U1389 (N_1389,N_155,In_955);
nand U1390 (N_1390,In_1963,N_41);
nor U1391 (N_1391,In_3581,In_2383);
or U1392 (N_1392,In_432,N_926);
nor U1393 (N_1393,In_513,In_4166);
nand U1394 (N_1394,In_4717,In_4276);
and U1395 (N_1395,In_3501,In_4936);
or U1396 (N_1396,In_4983,In_4006);
nor U1397 (N_1397,In_75,In_4088);
nor U1398 (N_1398,In_4594,In_1060);
or U1399 (N_1399,N_52,In_2650);
xor U1400 (N_1400,In_765,N_908);
nand U1401 (N_1401,N_538,N_377);
or U1402 (N_1402,In_146,In_1477);
or U1403 (N_1403,In_725,N_446);
nor U1404 (N_1404,In_4051,N_805);
xor U1405 (N_1405,In_127,In_2846);
or U1406 (N_1406,In_1094,N_613);
and U1407 (N_1407,In_1076,In_2090);
and U1408 (N_1408,In_374,In_993);
nand U1409 (N_1409,In_3260,In_98);
and U1410 (N_1410,In_2151,In_3886);
nor U1411 (N_1411,In_4168,N_572);
nand U1412 (N_1412,In_857,In_4139);
and U1413 (N_1413,N_95,N_272);
nor U1414 (N_1414,In_2207,In_3530);
nand U1415 (N_1415,N_730,N_544);
nand U1416 (N_1416,In_2662,In_2346);
and U1417 (N_1417,In_2013,In_1892);
xor U1418 (N_1418,In_3643,In_3441);
nand U1419 (N_1419,In_1387,In_4817);
or U1420 (N_1420,In_2848,In_462);
nor U1421 (N_1421,N_652,N_800);
and U1422 (N_1422,In_1432,In_4355);
nand U1423 (N_1423,In_3721,In_4383);
nor U1424 (N_1424,In_3515,In_2399);
and U1425 (N_1425,In_1320,In_3477);
and U1426 (N_1426,In_2248,In_4997);
xnor U1427 (N_1427,N_853,N_832);
and U1428 (N_1428,In_215,In_2981);
nor U1429 (N_1429,In_2359,In_4629);
or U1430 (N_1430,In_1524,In_4612);
or U1431 (N_1431,In_2009,In_1488);
and U1432 (N_1432,In_771,In_2316);
nor U1433 (N_1433,In_4482,In_3730);
or U1434 (N_1434,N_884,N_458);
xor U1435 (N_1435,In_1351,In_4432);
xor U1436 (N_1436,In_1610,N_273);
nand U1437 (N_1437,In_3144,In_3446);
or U1438 (N_1438,In_2783,In_3482);
nand U1439 (N_1439,N_740,N_252);
nand U1440 (N_1440,In_3630,In_1168);
nand U1441 (N_1441,In_1716,N_362);
nor U1442 (N_1442,In_282,In_3548);
or U1443 (N_1443,In_4231,In_3280);
xnor U1444 (N_1444,In_4984,In_666);
nor U1445 (N_1445,N_877,In_1128);
or U1446 (N_1446,In_748,In_2137);
nor U1447 (N_1447,In_90,In_3533);
nor U1448 (N_1448,In_2350,N_478);
nor U1449 (N_1449,In_4208,In_4645);
nand U1450 (N_1450,N_376,In_2052);
nand U1451 (N_1451,In_1355,N_401);
nand U1452 (N_1452,In_431,In_4181);
or U1453 (N_1453,In_3127,In_2020);
nor U1454 (N_1454,In_3411,In_3881);
or U1455 (N_1455,In_4077,N_951);
xnor U1456 (N_1456,In_3141,In_4651);
and U1457 (N_1457,In_4378,In_2778);
nand U1458 (N_1458,In_2039,In_3348);
nand U1459 (N_1459,N_659,In_1441);
nand U1460 (N_1460,In_4896,N_650);
or U1461 (N_1461,In_1670,N_274);
nand U1462 (N_1462,In_4660,In_4564);
xnor U1463 (N_1463,In_3976,N_453);
nor U1464 (N_1464,In_4015,In_959);
xnor U1465 (N_1465,In_1082,N_807);
nor U1466 (N_1466,In_3369,N_240);
and U1467 (N_1467,In_3570,N_46);
and U1468 (N_1468,N_201,In_3794);
xnor U1469 (N_1469,In_3879,In_3341);
nor U1470 (N_1470,In_3777,In_4428);
nor U1471 (N_1471,In_2342,In_4982);
xor U1472 (N_1472,N_279,In_3563);
nand U1473 (N_1473,In_2139,N_672);
or U1474 (N_1474,In_4457,In_2059);
and U1475 (N_1475,In_836,In_3519);
nor U1476 (N_1476,In_2952,In_1667);
nor U1477 (N_1477,In_632,In_3231);
nand U1478 (N_1478,In_4321,N_865);
nand U1479 (N_1479,In_518,In_2926);
nand U1480 (N_1480,In_521,In_4844);
nand U1481 (N_1481,In_4030,In_3454);
or U1482 (N_1482,N_734,In_3438);
nand U1483 (N_1483,N_173,In_3343);
xor U1484 (N_1484,In_3412,N_448);
or U1485 (N_1485,In_4,In_3658);
or U1486 (N_1486,In_1620,In_2534);
and U1487 (N_1487,In_2444,N_305);
nand U1488 (N_1488,In_4474,In_2658);
or U1489 (N_1489,In_2669,N_684);
nand U1490 (N_1490,In_1115,N_953);
and U1491 (N_1491,N_608,N_666);
or U1492 (N_1492,N_895,In_3392);
nand U1493 (N_1493,In_4632,In_383);
and U1494 (N_1494,In_2015,In_2278);
nor U1495 (N_1495,In_3043,N_436);
xor U1496 (N_1496,N_147,N_423);
or U1497 (N_1497,N_197,In_3456);
xor U1498 (N_1498,N_822,In_3526);
xor U1499 (N_1499,In_1816,In_1172);
nand U1500 (N_1500,In_4074,N_698);
or U1501 (N_1501,In_4788,In_1014);
or U1502 (N_1502,N_691,In_4392);
or U1503 (N_1503,In_2045,In_1305);
xor U1504 (N_1504,In_4607,In_579);
nand U1505 (N_1505,In_3011,N_565);
nand U1506 (N_1506,In_619,In_3090);
xnor U1507 (N_1507,In_3906,In_1862);
nor U1508 (N_1508,In_278,In_3503);
and U1509 (N_1509,In_2255,In_2550);
or U1510 (N_1510,In_1900,N_933);
nor U1511 (N_1511,In_4038,In_1806);
and U1512 (N_1512,In_134,In_1970);
nand U1513 (N_1513,In_1016,In_1148);
nand U1514 (N_1514,N_667,In_2239);
nand U1515 (N_1515,In_4778,In_13);
nor U1516 (N_1516,In_705,N_932);
and U1517 (N_1517,In_4615,In_1911);
or U1518 (N_1518,In_1800,N_586);
nor U1519 (N_1519,N_199,In_1808);
xnor U1520 (N_1520,In_4816,In_2340);
xnor U1521 (N_1521,In_4084,N_247);
nand U1522 (N_1522,In_3036,N_370);
xor U1523 (N_1523,In_2328,N_821);
xor U1524 (N_1524,In_4727,In_2640);
nand U1525 (N_1525,N_45,N_889);
nand U1526 (N_1526,N_36,N_344);
or U1527 (N_1527,N_917,In_977);
nor U1528 (N_1528,N_592,N_496);
nor U1529 (N_1529,In_635,In_3249);
and U1530 (N_1530,In_3661,N_413);
xor U1531 (N_1531,N_393,In_3592);
nor U1532 (N_1532,In_3374,In_4239);
and U1533 (N_1533,In_2306,In_1711);
xnor U1534 (N_1534,In_4025,N_43);
nor U1535 (N_1535,In_1760,In_4956);
or U1536 (N_1536,In_2398,In_3694);
nor U1537 (N_1537,In_2474,N_798);
or U1538 (N_1538,N_528,N_564);
xor U1539 (N_1539,N_729,In_406);
and U1540 (N_1540,N_540,In_4494);
or U1541 (N_1541,In_3702,N_1);
nand U1542 (N_1542,In_3988,In_4369);
nand U1543 (N_1543,In_4009,N_513);
and U1544 (N_1544,N_855,N_767);
nor U1545 (N_1545,In_2070,In_4518);
or U1546 (N_1546,N_186,In_4978);
and U1547 (N_1547,In_294,In_3819);
or U1548 (N_1548,In_4215,N_395);
xor U1549 (N_1549,In_3371,In_2489);
nand U1550 (N_1550,In_3329,In_1141);
nor U1551 (N_1551,N_600,In_4772);
and U1552 (N_1552,In_2636,In_144);
nor U1553 (N_1553,In_4437,In_2804);
and U1554 (N_1554,In_738,In_4574);
nand U1555 (N_1555,In_2110,In_2018);
or U1556 (N_1556,In_2491,In_4372);
xnor U1557 (N_1557,In_1580,N_449);
nor U1558 (N_1558,N_75,In_3321);
nand U1559 (N_1559,In_4421,N_363);
xor U1560 (N_1560,In_2404,In_4527);
nand U1561 (N_1561,In_3937,In_3407);
or U1562 (N_1562,In_4200,In_792);
xnor U1563 (N_1563,In_2265,N_715);
xnor U1564 (N_1564,In_3512,In_4714);
xnor U1565 (N_1565,In_2380,In_568);
nand U1566 (N_1566,In_1142,In_1837);
nor U1567 (N_1567,N_890,N_529);
or U1568 (N_1568,N_220,In_4016);
nand U1569 (N_1569,In_1157,In_4883);
or U1570 (N_1570,In_1050,In_2369);
xnor U1571 (N_1571,In_3409,In_2840);
or U1572 (N_1572,In_2733,N_319);
and U1573 (N_1573,In_1059,In_2006);
xor U1574 (N_1574,N_61,N_21);
and U1575 (N_1575,In_4737,In_895);
or U1576 (N_1576,In_2281,In_2362);
or U1577 (N_1577,In_2989,In_3001);
xnor U1578 (N_1578,In_2759,N_151);
xnor U1579 (N_1579,In_1513,N_7);
nor U1580 (N_1580,In_3518,In_1560);
nand U1581 (N_1581,In_1265,In_3408);
xor U1582 (N_1582,In_201,In_4241);
and U1583 (N_1583,In_366,In_1047);
nand U1584 (N_1584,N_845,In_3845);
nand U1585 (N_1585,In_2826,N_625);
and U1586 (N_1586,In_3297,In_1012);
nand U1587 (N_1587,In_3394,N_115);
nand U1588 (N_1588,In_903,In_1049);
and U1589 (N_1589,N_391,In_3499);
nand U1590 (N_1590,In_2294,N_627);
nand U1591 (N_1591,In_2354,In_2365);
or U1592 (N_1592,In_3445,In_1201);
or U1593 (N_1593,N_13,N_663);
or U1594 (N_1594,N_29,In_4357);
xor U1595 (N_1595,In_2433,In_3303);
xnor U1596 (N_1596,In_920,In_1231);
nand U1597 (N_1597,In_4395,In_2127);
nand U1598 (N_1598,In_4220,In_3246);
xor U1599 (N_1599,In_1496,In_2121);
xor U1600 (N_1600,In_750,N_310);
nor U1601 (N_1601,In_2614,In_4014);
nand U1602 (N_1602,In_4111,In_4467);
or U1603 (N_1603,In_3325,N_421);
and U1604 (N_1604,In_1796,In_4560);
nand U1605 (N_1605,In_4382,In_954);
and U1606 (N_1606,In_3415,In_2564);
nor U1607 (N_1607,In_4677,N_964);
nand U1608 (N_1608,N_918,In_4032);
and U1609 (N_1609,N_128,In_2221);
nand U1610 (N_1610,In_3221,In_2030);
xnor U1611 (N_1611,N_957,In_3825);
or U1612 (N_1612,N_207,N_339);
and U1613 (N_1613,In_694,In_477);
nor U1614 (N_1614,In_3946,In_3496);
and U1615 (N_1615,In_4058,In_198);
nand U1616 (N_1616,N_311,In_926);
xnor U1617 (N_1617,In_3793,In_2085);
or U1618 (N_1618,N_717,In_2144);
or U1619 (N_1619,N_187,In_4371);
and U1620 (N_1620,In_4087,N_208);
nor U1621 (N_1621,In_4151,In_337);
or U1622 (N_1622,In_960,In_1023);
and U1623 (N_1623,In_30,In_119);
nand U1624 (N_1624,In_2735,N_289);
xnor U1625 (N_1625,N_331,In_4264);
or U1626 (N_1626,In_4278,In_3464);
or U1627 (N_1627,In_2576,N_85);
and U1628 (N_1628,N_451,N_560);
or U1629 (N_1629,In_4804,In_1669);
or U1630 (N_1630,In_4227,In_2325);
and U1631 (N_1631,N_132,N_841);
xor U1632 (N_1632,N_507,In_4327);
nor U1633 (N_1633,In_2285,N_427);
and U1634 (N_1634,In_1836,In_4609);
nand U1635 (N_1635,In_247,In_2771);
xor U1636 (N_1636,In_4986,N_293);
and U1637 (N_1637,In_1953,In_737);
nor U1638 (N_1638,In_3027,In_391);
xor U1639 (N_1639,N_862,In_2053);
nand U1640 (N_1640,In_1090,In_3796);
and U1641 (N_1641,In_3202,N_563);
and U1642 (N_1642,In_4107,In_864);
or U1643 (N_1643,In_974,In_221);
nand U1644 (N_1644,In_2305,In_2872);
xor U1645 (N_1645,N_178,In_248);
and U1646 (N_1646,In_1910,N_246);
or U1647 (N_1647,In_2592,In_3345);
xor U1648 (N_1648,In_4164,In_997);
xnor U1649 (N_1649,In_2915,In_790);
xnor U1650 (N_1650,N_688,In_3327);
nand U1651 (N_1651,In_2591,In_3292);
nor U1652 (N_1652,In_2631,N_834);
nand U1653 (N_1653,N_476,In_228);
nor U1654 (N_1654,In_2694,In_2601);
xor U1655 (N_1655,In_4265,In_264);
nor U1656 (N_1656,In_209,N_323);
xor U1657 (N_1657,In_4919,In_837);
and U1658 (N_1658,N_522,In_299);
and U1659 (N_1659,In_3149,In_1436);
nor U1660 (N_1660,N_477,In_3715);
xor U1661 (N_1661,In_1285,In_2076);
and U1662 (N_1662,In_3781,In_3108);
or U1663 (N_1663,In_22,In_407);
nor U1664 (N_1664,N_741,N_771);
nand U1665 (N_1665,In_2412,In_3427);
nand U1666 (N_1666,In_2472,In_1280);
nor U1667 (N_1667,In_1317,In_1705);
and U1668 (N_1668,N_713,N_837);
nor U1669 (N_1669,In_3372,In_3109);
and U1670 (N_1670,In_581,In_345);
xor U1671 (N_1671,N_399,In_1021);
xnor U1672 (N_1672,N_819,In_4026);
nor U1673 (N_1673,In_3494,N_575);
or U1674 (N_1674,N_551,In_1902);
and U1675 (N_1675,N_160,In_4354);
nand U1676 (N_1676,In_166,In_2932);
and U1677 (N_1677,In_4699,In_167);
and U1678 (N_1678,In_3857,In_4995);
xor U1679 (N_1679,In_1382,In_1591);
xor U1680 (N_1680,In_2003,In_1547);
nand U1681 (N_1681,In_1458,N_447);
and U1682 (N_1682,In_1356,In_891);
nand U1683 (N_1683,In_141,N_744);
xnor U1684 (N_1684,In_2211,N_562);
nand U1685 (N_1685,In_918,In_686);
nand U1686 (N_1686,In_3990,In_908);
xor U1687 (N_1687,N_525,In_189);
and U1688 (N_1688,In_3867,N_739);
nor U1689 (N_1689,In_4879,In_3685);
and U1690 (N_1690,In_2907,In_4761);
or U1691 (N_1691,N_256,N_135);
or U1692 (N_1692,In_3203,In_2449);
nand U1693 (N_1693,In_3258,In_3185);
xor U1694 (N_1694,In_2879,In_690);
and U1695 (N_1695,In_2754,N_316);
xnor U1696 (N_1696,N_646,In_780);
nand U1697 (N_1697,In_219,In_4493);
and U1698 (N_1698,In_653,In_4926);
and U1699 (N_1699,In_2586,N_641);
and U1700 (N_1700,N_206,In_3256);
nor U1701 (N_1701,N_725,N_343);
and U1702 (N_1702,N_313,In_1950);
nand U1703 (N_1703,In_28,In_326);
and U1704 (N_1704,N_870,N_519);
nor U1705 (N_1705,In_205,In_2429);
nand U1706 (N_1706,N_732,In_2953);
xnor U1707 (N_1707,N_479,In_4555);
and U1708 (N_1708,In_4098,In_50);
nand U1709 (N_1709,In_1966,In_583);
and U1710 (N_1710,N_910,In_1408);
and U1711 (N_1711,In_1571,In_2824);
nor U1712 (N_1712,In_4295,In_814);
or U1713 (N_1713,N_567,N_676);
nand U1714 (N_1714,In_2886,In_3424);
nor U1715 (N_1715,In_4259,N_733);
nand U1716 (N_1716,N_533,In_120);
nand U1717 (N_1717,In_2470,In_2860);
and U1718 (N_1718,N_585,In_4028);
xnor U1719 (N_1719,N_164,In_2434);
and U1720 (N_1720,In_3436,In_2719);
nand U1721 (N_1721,In_2738,In_866);
xnor U1722 (N_1722,N_354,In_105);
xor U1723 (N_1723,In_946,In_2987);
or U1724 (N_1724,In_4814,In_3606);
nand U1725 (N_1725,N_660,In_4642);
nor U1726 (N_1726,N_928,In_2641);
nor U1727 (N_1727,N_722,N_260);
and U1728 (N_1728,In_281,In_3719);
or U1729 (N_1729,In_3091,In_3067);
nor U1730 (N_1730,In_1162,In_3516);
and U1731 (N_1731,In_270,In_3779);
nand U1732 (N_1732,In_4258,N_221);
and U1733 (N_1733,In_488,In_2752);
nor U1734 (N_1734,In_4471,N_571);
xnor U1735 (N_1735,In_3450,N_89);
nand U1736 (N_1736,N_647,N_108);
or U1737 (N_1737,N_842,In_2054);
xor U1738 (N_1738,In_15,In_2313);
xor U1739 (N_1739,In_2979,N_993);
nor U1740 (N_1740,N_665,In_3999);
and U1741 (N_1741,In_2172,In_4262);
or U1742 (N_1742,In_1979,In_3230);
nand U1743 (N_1743,N_270,In_3950);
nand U1744 (N_1744,In_443,N_893);
and U1745 (N_1745,In_88,In_3931);
and U1746 (N_1746,N_157,N_312);
and U1747 (N_1747,N_765,In_2011);
and U1748 (N_1748,In_450,In_1532);
nor U1749 (N_1749,In_999,In_3313);
and U1750 (N_1750,N_541,In_152);
nor U1751 (N_1751,In_1612,In_2511);
nor U1752 (N_1752,In_3861,In_4603);
xnor U1753 (N_1753,In_4893,In_1343);
or U1754 (N_1754,N_213,In_93);
and U1755 (N_1755,In_2464,In_1030);
nand U1756 (N_1756,In_4887,In_3404);
nor U1757 (N_1757,N_32,In_1614);
and U1758 (N_1758,In_2580,In_1749);
and U1759 (N_1759,In_3124,In_3181);
nand U1760 (N_1760,In_1909,N_875);
and U1761 (N_1761,N_960,N_83);
xnor U1762 (N_1762,N_580,In_3720);
xor U1763 (N_1763,In_1646,N_57);
or U1764 (N_1764,N_39,In_797);
xor U1765 (N_1765,In_4700,In_1310);
and U1766 (N_1766,N_772,In_2337);
and U1767 (N_1767,N_561,In_4435);
and U1768 (N_1768,N_336,In_2505);
nor U1769 (N_1769,In_2270,In_778);
and U1770 (N_1770,In_2273,N_250);
nor U1771 (N_1771,In_3319,N_371);
or U1772 (N_1772,In_2236,In_3610);
nor U1773 (N_1773,N_488,In_2583);
nand U1774 (N_1774,In_3991,In_3667);
nor U1775 (N_1775,N_162,In_1415);
xor U1776 (N_1776,In_2928,In_2268);
xor U1777 (N_1777,In_53,N_700);
nor U1778 (N_1778,In_514,N_176);
nand U1779 (N_1779,In_515,In_1638);
xnor U1780 (N_1780,In_905,N_318);
nand U1781 (N_1781,In_1119,In_2850);
or U1782 (N_1782,In_4866,In_1426);
nor U1783 (N_1783,In_4073,In_2197);
nor U1784 (N_1784,In_2366,In_940);
and U1785 (N_1785,N_995,N_662);
or U1786 (N_1786,N_911,N_584);
or U1787 (N_1787,In_2698,N_902);
xnor U1788 (N_1788,In_4303,In_3355);
xor U1789 (N_1789,In_1372,In_1452);
xor U1790 (N_1790,N_335,In_4836);
nor U1791 (N_1791,In_4153,In_3959);
or U1792 (N_1792,In_2747,In_126);
or U1793 (N_1793,In_4696,In_3268);
or U1794 (N_1794,In_4891,In_46);
nor U1795 (N_1795,In_1596,In_1940);
or U1796 (N_1796,N_415,In_3);
nor U1797 (N_1797,In_4201,N_671);
nand U1798 (N_1798,In_578,In_490);
or U1799 (N_1799,In_3272,In_1787);
or U1800 (N_1800,In_3253,In_4199);
and U1801 (N_1801,In_2562,In_3583);
xor U1802 (N_1802,In_773,In_2142);
or U1803 (N_1803,In_2279,N_499);
nand U1804 (N_1804,In_3252,N_355);
xnor U1805 (N_1805,In_4279,In_867);
nor U1806 (N_1806,In_4450,In_2258);
xnor U1807 (N_1807,In_1181,In_1992);
nor U1808 (N_1808,In_2645,In_4801);
xnor U1809 (N_1809,In_4272,In_2448);
and U1810 (N_1810,In_4287,In_3479);
nor U1811 (N_1811,In_985,In_3013);
or U1812 (N_1812,In_413,N_292);
xor U1813 (N_1813,In_3574,In_2231);
xnor U1814 (N_1814,In_1692,In_1954);
nand U1815 (N_1815,In_3549,In_1981);
xnor U1816 (N_1816,In_4597,N_615);
or U1817 (N_1817,N_287,In_2262);
nand U1818 (N_1818,In_2102,N_632);
xnor U1819 (N_1819,N_789,In_4865);
nand U1820 (N_1820,In_1019,In_2162);
and U1821 (N_1821,In_4563,In_4690);
nor U1822 (N_1822,In_1197,In_3786);
and U1823 (N_1823,In_2560,In_932);
xor U1824 (N_1824,N_110,In_3872);
nand U1825 (N_1825,In_266,N_781);
nand U1826 (N_1826,In_2839,In_4217);
nor U1827 (N_1827,In_4774,In_4631);
xnor U1828 (N_1828,In_4975,In_3119);
or U1829 (N_1829,N_894,In_1679);
xor U1830 (N_1830,In_106,In_2187);
nand U1831 (N_1831,In_1561,In_843);
and U1832 (N_1832,In_4575,N_460);
or U1833 (N_1833,In_1069,In_4290);
nor U1834 (N_1834,In_2982,In_1880);
and U1835 (N_1835,N_872,In_2722);
and U1836 (N_1836,In_4122,In_2016);
or U1837 (N_1837,In_1933,N_44);
nor U1838 (N_1838,In_1798,N_143);
and U1839 (N_1839,N_59,In_2466);
xor U1840 (N_1840,N_400,In_811);
nor U1841 (N_1841,In_3418,In_3107);
xnor U1842 (N_1842,N_746,In_2079);
xor U1843 (N_1843,In_3126,In_2964);
and U1844 (N_1844,N_681,In_4483);
and U1845 (N_1845,N_824,N_614);
nor U1846 (N_1846,In_4004,In_1333);
nand U1847 (N_1847,In_640,In_4134);
nor U1848 (N_1848,In_4767,In_582);
nor U1849 (N_1849,In_4041,In_4829);
nand U1850 (N_1850,In_3854,In_2894);
xnor U1851 (N_1851,In_2103,N_569);
nor U1852 (N_1852,In_2851,In_4205);
or U1853 (N_1853,In_236,In_2877);
nor U1854 (N_1854,N_217,In_1335);
nand U1855 (N_1855,N_535,N_654);
or U1856 (N_1856,In_1235,In_826);
xor U1857 (N_1857,In_4665,In_3828);
nor U1858 (N_1858,In_2822,In_3326);
or U1859 (N_1859,N_950,In_838);
and U1860 (N_1860,N_511,N_467);
nor U1861 (N_1861,N_439,N_80);
nand U1862 (N_1862,N_617,N_545);
and U1863 (N_1863,In_3393,In_2062);
or U1864 (N_1864,In_4475,In_4708);
nand U1865 (N_1865,In_4641,In_321);
and U1866 (N_1866,In_2984,In_1710);
nor U1867 (N_1867,In_242,In_2731);
nor U1868 (N_1868,N_200,In_1122);
xnor U1869 (N_1869,In_4928,In_2021);
or U1870 (N_1870,In_2739,N_596);
nand U1871 (N_1871,In_2375,In_1998);
or U1872 (N_1872,In_3855,N_259);
or U1873 (N_1873,In_1569,In_3790);
xnor U1874 (N_1874,In_4331,In_3961);
nor U1875 (N_1875,In_4298,N_181);
nor U1876 (N_1876,In_4682,In_1442);
or U1877 (N_1877,N_81,In_61);
nor U1878 (N_1878,In_3032,N_321);
nor U1879 (N_1879,In_4618,In_3128);
and U1880 (N_1880,In_560,N_306);
xor U1881 (N_1881,In_3509,In_3148);
and U1882 (N_1882,In_3752,In_4551);
and U1883 (N_1883,In_3084,In_2140);
nor U1884 (N_1884,In_2147,In_3500);
and U1885 (N_1885,In_4351,In_3187);
nor U1886 (N_1886,N_253,In_835);
and U1887 (N_1887,In_468,In_3919);
or U1888 (N_1888,In_3591,In_1227);
nor U1889 (N_1889,N_752,In_178);
xor U1890 (N_1890,N_175,N_644);
and U1891 (N_1891,In_292,In_1498);
xor U1892 (N_1892,In_772,In_1179);
or U1893 (N_1893,In_884,In_2652);
or U1894 (N_1894,In_597,In_3683);
xor U1895 (N_1895,In_1466,In_118);
or U1896 (N_1896,In_2852,In_2234);
xnor U1897 (N_1897,In_3970,In_1304);
nand U1898 (N_1898,In_1006,In_2797);
xnor U1899 (N_1899,In_4529,In_4377);
xnor U1900 (N_1900,In_2182,In_2493);
nor U1901 (N_1901,N_167,In_1899);
nand U1902 (N_1902,In_4781,In_795);
xnor U1903 (N_1903,In_2508,In_880);
or U1904 (N_1904,In_1712,In_3768);
or U1905 (N_1905,In_4712,In_2675);
nand U1906 (N_1906,In_680,In_2762);
nor U1907 (N_1907,In_2217,In_296);
nand U1908 (N_1908,In_2993,N_574);
or U1909 (N_1909,In_3738,In_4043);
and U1910 (N_1910,In_3059,In_1371);
nor U1911 (N_1911,In_1661,In_1927);
and U1912 (N_1912,In_1807,In_2805);
xor U1913 (N_1913,In_942,N_687);
xor U1914 (N_1914,In_4831,In_4363);
xor U1915 (N_1915,In_3014,In_1574);
nor U1916 (N_1916,In_3062,In_2459);
nand U1917 (N_1917,In_3065,In_3305);
nor U1918 (N_1918,In_356,N_944);
nor U1919 (N_1919,N_117,N_904);
nor U1920 (N_1920,N_4,In_4063);
nor U1921 (N_1921,N_920,In_1957);
and U1922 (N_1922,In_4636,In_1401);
nor U1923 (N_1923,In_2133,In_1777);
xnor U1924 (N_1924,In_2642,N_622);
nand U1925 (N_1925,In_844,In_1483);
nand U1926 (N_1926,In_137,In_4562);
nor U1927 (N_1927,N_298,In_2113);
nand U1928 (N_1928,In_4550,In_1033);
and U1929 (N_1929,In_2776,In_2899);
nand U1930 (N_1930,In_1406,In_4728);
xnor U1931 (N_1931,In_470,In_2246);
and U1932 (N_1932,In_2800,In_522);
and U1933 (N_1933,In_994,N_981);
xor U1934 (N_1934,N_686,In_2898);
nor U1935 (N_1935,In_2303,N_163);
nand U1936 (N_1936,In_2639,In_441);
and U1937 (N_1937,In_2509,In_200);
nand U1938 (N_1938,In_4176,In_4666);
and U1939 (N_1939,N_508,N_465);
xor U1940 (N_1940,N_416,In_3753);
xor U1941 (N_1941,N_113,In_2858);
nand U1942 (N_1942,N_288,In_3311);
nand U1943 (N_1943,In_4602,N_275);
xor U1944 (N_1944,N_441,In_1949);
and U1945 (N_1945,N_387,In_1834);
or U1946 (N_1946,In_4614,In_4890);
nor U1947 (N_1947,N_498,In_4477);
and U1948 (N_1948,In_1563,In_802);
nor U1949 (N_1949,In_1166,In_4334);
and U1950 (N_1950,In_3138,In_3891);
xnor U1951 (N_1951,In_2347,In_3080);
and U1952 (N_1952,In_3641,In_1520);
nand U1953 (N_1953,In_4640,N_37);
nor U1954 (N_1954,N_452,N_492);
or U1955 (N_1955,In_1155,In_4910);
nor U1956 (N_1956,In_1559,In_510);
nor U1957 (N_1957,N_237,In_10);
xnor U1958 (N_1958,In_3037,In_3579);
nand U1959 (N_1959,In_4393,N_764);
xor U1960 (N_1960,In_2254,In_3054);
nor U1961 (N_1961,In_4693,In_2569);
nor U1962 (N_1962,In_2602,In_4770);
xor U1963 (N_1963,N_227,In_2319);
or U1964 (N_1964,N_649,In_4895);
nand U1965 (N_1965,N_314,In_1174);
nand U1966 (N_1966,In_4613,In_3788);
and U1967 (N_1967,N_68,N_675);
nand U1968 (N_1968,In_2990,In_3926);
xor U1969 (N_1969,N_977,In_1144);
nand U1970 (N_1970,In_4370,In_3960);
and U1971 (N_1971,In_3843,In_4566);
nor U1972 (N_1972,In_1061,In_4053);
or U1973 (N_1973,In_1338,In_2666);
and U1974 (N_1974,In_1876,N_140);
and U1975 (N_1975,N_914,In_286);
or U1976 (N_1976,N_268,In_1270);
and U1977 (N_1977,N_146,In_4075);
or U1978 (N_1978,In_1639,In_3935);
nand U1979 (N_1979,In_537,N_750);
or U1980 (N_1980,In_3267,N_759);
xor U1981 (N_1981,N_929,In_3621);
nand U1982 (N_1982,N_801,In_3814);
or U1983 (N_1983,N_348,In_575);
nand U1984 (N_1984,N_982,In_3363);
xor U1985 (N_1985,In_2793,In_2881);
xnor U1986 (N_1986,In_336,N_796);
nand U1987 (N_1987,In_983,In_1158);
nor U1988 (N_1988,In_764,In_2519);
and U1989 (N_1989,In_70,In_1626);
or U1990 (N_1990,In_2243,N_338);
or U1991 (N_1991,In_3030,In_388);
or U1992 (N_1992,In_1584,In_917);
and U1993 (N_1993,N_847,In_2997);
and U1994 (N_1994,N_320,In_3746);
or U1995 (N_1995,In_331,In_770);
nor U1996 (N_1996,In_3633,In_2812);
nand U1997 (N_1997,In_1362,In_677);
and U1998 (N_1998,In_1865,In_937);
xor U1999 (N_1999,N_991,In_2704);
and U2000 (N_2000,In_4972,In_2432);
and U2001 (N_2001,N_122,N_233);
or U2002 (N_2002,N_1666,N_1698);
nand U2003 (N_2003,In_279,N_1028);
nor U2004 (N_2004,In_2,N_25);
and U2005 (N_2005,N_946,In_973);
xor U2006 (N_2006,In_3676,N_1262);
nand U2007 (N_2007,In_2919,N_42);
nor U2008 (N_2008,N_1580,In_4242);
nor U2009 (N_2009,In_1032,In_3792);
xnor U2010 (N_2010,N_1999,In_4765);
and U2011 (N_2011,In_4941,N_1812);
xnor U2012 (N_2012,In_831,In_2854);
nor U2013 (N_2013,In_1994,In_1897);
or U2014 (N_2014,In_3359,In_1282);
nor U2015 (N_2015,N_1743,N_1946);
xnor U2016 (N_2016,N_1068,In_1702);
xnor U2017 (N_2017,N_1438,In_4987);
and U2018 (N_2018,N_215,In_2171);
and U2019 (N_2019,In_3169,N_500);
or U2020 (N_2020,N_1491,N_1710);
nand U2021 (N_2021,In_2087,In_984);
nor U2022 (N_2022,N_850,N_1356);
nand U2023 (N_2023,In_1350,N_1344);
xnor U2024 (N_2024,In_102,N_1218);
and U2025 (N_2025,N_345,N_1521);
or U2026 (N_2026,In_473,In_1182);
nand U2027 (N_2027,N_1430,N_1335);
nand U2028 (N_2028,In_3992,N_527);
xor U2029 (N_2029,In_2657,N_1486);
or U2030 (N_2030,N_1602,In_2403);
nand U2031 (N_2031,In_2769,In_2875);
nor U2032 (N_2032,In_626,In_2920);
and U2033 (N_2033,In_3452,In_1163);
nor U2034 (N_2034,In_285,In_3051);
xor U2035 (N_2035,In_2492,N_502);
and U2036 (N_2036,In_1225,In_544);
xnor U2037 (N_2037,N_1185,In_2048);
and U2038 (N_2038,N_1914,In_4460);
and U2039 (N_2039,In_4625,In_3399);
and U2040 (N_2040,In_945,In_4172);
and U2041 (N_2041,N_1865,In_3545);
nor U2042 (N_2042,N_1053,In_1056);
nor U2043 (N_2043,N_661,N_1747);
nor U2044 (N_2044,In_3817,N_97);
or U2045 (N_2045,N_1131,N_1951);
or U2046 (N_2046,In_3884,In_3236);
nand U2047 (N_2047,In_4270,In_4229);
nand U2048 (N_2048,N_209,In_1260);
nand U2049 (N_2049,In_449,N_469);
xor U2050 (N_2050,N_1687,In_3995);
xnor U2051 (N_2051,In_335,N_133);
nor U2052 (N_2052,In_2684,In_3060);
and U2053 (N_2053,N_1682,N_1174);
nand U2054 (N_2054,In_2157,In_3049);
nor U2055 (N_2055,N_442,N_1460);
nand U2056 (N_2056,N_1990,In_3170);
and U2057 (N_2057,N_1154,N_1412);
nand U2058 (N_2058,N_72,N_640);
xnor U2059 (N_2059,In_2999,In_2937);
or U2060 (N_2060,In_1758,N_888);
and U2061 (N_2061,N_549,N_1340);
nor U2062 (N_2062,In_1391,In_2063);
or U2063 (N_2063,N_12,N_1357);
nand U2064 (N_2064,N_14,In_2913);
xnor U2065 (N_2065,In_2610,In_1214);
nor U2066 (N_2066,In_4588,In_4932);
or U2067 (N_2067,N_939,N_1288);
nor U2068 (N_2068,In_1440,In_1809);
nand U2069 (N_2069,In_1271,In_399);
and U2070 (N_2070,N_1187,N_1668);
or U2071 (N_2071,In_4782,In_238);
nand U2072 (N_2072,In_1642,N_1448);
xor U2073 (N_2073,In_1029,In_1275);
and U2074 (N_2074,N_1007,In_1657);
and U2075 (N_2075,In_2986,N_947);
nor U2076 (N_2076,In_2089,N_1182);
and U2077 (N_2077,N_1127,N_1504);
nor U2078 (N_2078,In_2439,In_1717);
nand U2079 (N_2079,N_360,N_1258);
and U2080 (N_2080,N_854,In_2667);
or U2081 (N_2081,In_1537,In_4306);
nor U2082 (N_2082,In_2296,N_1853);
xnor U2083 (N_2083,In_351,N_1327);
nand U2084 (N_2084,N_138,In_2336);
nor U2085 (N_2085,N_626,N_1518);
or U2086 (N_2086,N_1786,In_58);
xor U2087 (N_2087,N_486,N_1027);
xor U2088 (N_2088,In_1040,N_1933);
or U2089 (N_2089,In_2247,N_1114);
and U2090 (N_2090,N_515,In_4129);
nand U2091 (N_2091,In_1923,N_1723);
nand U2092 (N_2092,N_210,N_583);
nor U2093 (N_2093,N_481,N_1221);
xnor U2094 (N_2094,N_534,N_755);
and U2095 (N_2095,N_1211,In_4186);
and U2096 (N_2096,N_1202,N_1032);
nor U2097 (N_2097,N_2,N_1557);
and U2098 (N_2098,In_361,N_30);
and U2099 (N_2099,N_1167,In_3853);
nor U2100 (N_2100,N_1598,In_4807);
nor U2101 (N_2101,N_1330,N_1847);
nor U2102 (N_2102,In_1844,N_843);
or U2103 (N_2103,In_1263,N_512);
and U2104 (N_2104,In_1419,In_1912);
and U2105 (N_2105,N_1308,In_2970);
nand U2106 (N_2106,In_2829,N_1015);
nor U2107 (N_2107,In_3789,In_915);
xor U2108 (N_2108,N_1189,In_511);
nor U2109 (N_2109,In_1084,In_1780);
or U2110 (N_2110,In_2293,N_1453);
or U2111 (N_2111,N_1966,In_3953);
nand U2112 (N_2112,N_1246,N_1214);
and U2113 (N_2113,N_1768,N_1183);
or U2114 (N_2114,In_2718,In_3822);
and U2115 (N_2115,In_4464,In_683);
or U2116 (N_2116,In_4957,N_975);
nor U2117 (N_2117,N_1284,N_1950);
and U2118 (N_2118,In_2541,N_1061);
nand U2119 (N_2119,N_1299,N_1538);
xnor U2120 (N_2120,N_1199,N_1215);
xor U2121 (N_2121,N_1461,N_689);
and U2122 (N_2122,In_1018,N_1592);
nor U2123 (N_2123,In_262,N_1177);
and U2124 (N_2124,In_193,N_595);
nand U2125 (N_2125,N_590,N_1331);
nand U2126 (N_2126,N_1248,N_1004);
nand U2127 (N_2127,In_3703,N_165);
or U2128 (N_2128,N_1393,N_1144);
nor U2129 (N_2129,In_3064,In_3481);
or U2130 (N_2130,In_4671,In_439);
nor U2131 (N_2131,N_1540,In_3222);
xnor U2132 (N_2132,In_4680,In_2010);
xnor U2133 (N_2133,N_1235,N_1827);
and U2134 (N_2134,N_1281,In_3354);
and U2135 (N_2135,In_4906,In_4399);
nand U2136 (N_2136,In_500,In_588);
and U2137 (N_2137,N_1120,N_1336);
nand U2138 (N_2138,In_3038,In_4092);
or U2139 (N_2139,In_4815,N_885);
nor U2140 (N_2140,N_475,N_988);
nand U2141 (N_2141,N_1316,In_2889);
xnor U2142 (N_2142,N_1625,In_2632);
nor U2143 (N_2143,N_1569,N_724);
and U2144 (N_2144,In_440,N_1473);
and U2145 (N_2145,N_1632,In_1969);
and U2146 (N_2146,In_2078,N_1022);
xor U2147 (N_2147,N_1194,N_1509);
nand U2148 (N_2148,N_1887,N_1888);
xnor U2149 (N_2149,N_974,N_238);
or U2150 (N_2150,N_1361,N_257);
and U2151 (N_2151,In_3041,N_1526);
and U2152 (N_2152,In_4234,N_1434);
and U2153 (N_2153,N_695,In_4870);
or U2154 (N_2154,In_1730,N_1241);
and U2155 (N_2155,N_1806,In_2099);
nor U2156 (N_2156,In_3077,In_3576);
nand U2157 (N_2157,N_1721,In_4138);
or U2158 (N_2158,In_3324,In_301);
nor U2159 (N_2159,N_1819,N_1346);
nand U2160 (N_2160,N_1195,In_3475);
and U2161 (N_2161,N_9,N_930);
nor U2162 (N_2162,In_2905,In_43);
and U2163 (N_2163,In_3428,N_1717);
nor U2164 (N_2164,In_4339,In_3634);
xnor U2165 (N_2165,In_31,In_4577);
xor U2166 (N_2166,N_1096,In_643);
xor U2167 (N_2167,N_431,N_1209);
xor U2168 (N_2168,N_1444,N_1441);
nand U2169 (N_2169,In_3291,In_3212);
and U2170 (N_2170,In_2963,In_4040);
or U2171 (N_2171,N_35,N_1103);
and U2172 (N_2172,In_2789,In_82);
nor U2173 (N_2173,N_1776,In_1846);
xor U2174 (N_2174,In_3402,In_1367);
or U2175 (N_2175,In_4876,N_150);
nor U2176 (N_2176,In_1801,In_3164);
nor U2177 (N_2177,In_1118,In_4656);
nand U2178 (N_2178,In_2299,N_616);
and U2179 (N_2179,N_1677,N_1571);
nand U2180 (N_2180,In_378,N_1086);
nor U2181 (N_2181,N_470,N_909);
nor U2182 (N_2182,N_912,In_3636);
nand U2183 (N_2183,In_963,In_4822);
nand U2184 (N_2184,N_1132,In_3451);
or U2185 (N_2185,In_1412,In_3553);
or U2186 (N_2186,In_4060,N_428);
xnor U2187 (N_2187,In_1219,In_4498);
or U2188 (N_2188,In_547,N_954);
nand U2189 (N_2189,In_3285,N_1880);
nand U2190 (N_2190,In_3543,In_3386);
xnor U2191 (N_2191,N_1379,In_4365);
and U2192 (N_2192,In_3885,In_1633);
nor U2193 (N_2193,In_3798,In_3695);
nor U2194 (N_2194,N_555,In_681);
and U2195 (N_2195,In_4855,N_1635);
xnor U2196 (N_2196,N_1146,In_4219);
xor U2197 (N_2197,In_4930,In_4375);
nand U2198 (N_2198,In_3682,In_4411);
or U2199 (N_2199,N_1186,N_262);
nand U2200 (N_2200,N_1525,N_1275);
nand U2201 (N_2201,N_1111,N_934);
and U2202 (N_2202,In_2890,N_1133);
xnor U2203 (N_2203,In_3759,In_1660);
nand U2204 (N_2204,In_4156,N_1590);
and U2205 (N_2205,In_1139,N_504);
nand U2206 (N_2206,N_1934,In_1829);
and U2207 (N_2207,N_1077,N_1549);
or U2208 (N_2208,N_1554,N_1296);
and U2209 (N_2209,In_534,N_1319);
xor U2210 (N_2210,N_1545,In_769);
or U2211 (N_2211,N_1947,N_1309);
or U2212 (N_2212,N_1727,In_2673);
or U2213 (N_2213,In_781,In_4359);
and U2214 (N_2214,N_1232,In_4981);
nor U2215 (N_2215,In_4472,N_1205);
xor U2216 (N_2216,In_2548,In_3247);
nor U2217 (N_2217,N_1979,N_1919);
or U2218 (N_2218,In_4224,N_664);
or U2219 (N_2219,N_923,In_3505);
and U2220 (N_2220,N_1739,In_3837);
or U2221 (N_2221,In_1003,In_245);
nand U2222 (N_2222,N_1909,N_1588);
xor U2223 (N_2223,N_501,N_736);
nand U2224 (N_2224,N_1793,N_1210);
or U2225 (N_2225,In_1685,N_559);
or U2226 (N_2226,In_2933,N_1551);
nor U2227 (N_2227,N_1064,N_1041);
nor U2228 (N_2228,In_2873,N_222);
nand U2229 (N_2229,N_1570,In_4543);
and U2230 (N_2230,N_1409,N_1069);
and U2231 (N_2231,In_4230,N_601);
nor U2232 (N_2232,N_189,In_2287);
and U2233 (N_2233,N_1115,In_2368);
or U2234 (N_2234,In_1858,In_617);
and U2235 (N_2235,N_1302,In_3674);
and U2236 (N_2236,In_4877,N_1906);
nand U2237 (N_2237,N_1529,N_1977);
nand U2238 (N_2238,In_4626,In_2949);
nor U2239 (N_2239,N_1782,N_1586);
and U2240 (N_2240,N_1901,In_2153);
xnor U2241 (N_2241,In_4072,In_4386);
and U2242 (N_2242,N_1458,N_711);
nand U2243 (N_2243,In_4048,In_4637);
or U2244 (N_2244,N_1672,N_1832);
or U2245 (N_2245,In_636,N_1321);
xor U2246 (N_2246,N_1603,N_1980);
nand U2247 (N_2247,N_1324,N_1137);
nor U2248 (N_2248,In_2837,In_4863);
xor U2249 (N_2249,N_1607,N_835);
xnor U2250 (N_2250,In_2058,In_1370);
or U2251 (N_2251,N_714,In_3911);
xor U2252 (N_2252,In_1995,In_312);
and U2253 (N_2253,N_361,N_1043);
and U2254 (N_2254,In_2124,In_4302);
xnor U2255 (N_2255,In_66,In_3945);
nand U2256 (N_2256,In_3180,In_4361);
or U2257 (N_2257,N_1584,In_3727);
xnor U2258 (N_2258,N_180,In_2529);
nand U2259 (N_2259,In_1273,In_1840);
and U2260 (N_2260,In_2495,In_1928);
xnor U2261 (N_2261,N_1534,N_1255);
or U2262 (N_2262,In_3010,N_426);
xnor U2263 (N_2263,N_1003,In_4825);
nor U2264 (N_2264,In_3400,N_1965);
xor U2265 (N_2265,In_4685,N_1799);
and U2266 (N_2266,N_1542,N_1937);
xor U2267 (N_2267,N_1972,N_963);
nand U2268 (N_2268,In_821,N_774);
and U2269 (N_2269,In_3058,N_1879);
xnor U2270 (N_2270,N_1796,N_1969);
nand U2271 (N_2271,In_4894,N_1396);
nand U2272 (N_2272,N_1629,N_1333);
nor U2273 (N_2273,N_1341,N_1599);
nor U2274 (N_2274,In_3907,In_662);
and U2275 (N_2275,In_4486,In_1659);
nor U2276 (N_2276,N_424,In_1324);
and U2277 (N_2277,In_1159,In_692);
xor U2278 (N_2278,In_244,In_4036);
or U2279 (N_2279,N_301,N_1121);
nand U2280 (N_2280,N_408,In_2372);
or U2281 (N_2281,N_1314,In_2298);
and U2282 (N_2282,N_1926,N_1092);
nor U2283 (N_2283,In_2096,N_27);
or U2284 (N_2284,N_1217,In_4854);
xor U2285 (N_2285,In_4698,N_892);
or U2286 (N_2286,In_3573,In_459);
or U2287 (N_2287,In_4147,In_1253);
nor U2288 (N_2288,In_402,N_1463);
or U2289 (N_2289,N_866,In_2924);
nand U2290 (N_2290,In_1693,N_594);
nor U2291 (N_2291,In_3262,In_618);
nor U2292 (N_2292,In_1293,N_332);
nand U2293 (N_2293,In_2996,N_1113);
nor U2294 (N_2294,In_3223,In_1918);
or U2295 (N_2295,N_962,N_924);
nand U2296 (N_2296,In_3875,N_1225);
nand U2297 (N_2297,N_1544,N_1732);
or U2298 (N_2298,N_803,N_1274);
xnor U2299 (N_2299,N_1696,In_1308);
and U2300 (N_2300,N_1454,In_1740);
or U2301 (N_2301,In_805,N_568);
nand U2302 (N_2302,N_1385,In_2263);
and U2303 (N_2303,In_2348,In_1832);
nand U2304 (N_2304,N_1746,In_1438);
xnor U2305 (N_2305,In_2818,In_1930);
nor U2306 (N_2306,In_3688,N_1814);
nand U2307 (N_2307,N_1078,In_1169);
nand U2308 (N_2308,In_3189,N_1135);
nor U2309 (N_2309,N_366,N_1443);
or U2310 (N_2310,In_273,In_978);
nand U2311 (N_2311,N_1013,N_1143);
nand U2312 (N_2312,In_4686,N_1943);
nor U2313 (N_2313,N_1469,In_4552);
xor U2314 (N_2314,N_161,In_4977);
or U2315 (N_2315,In_1522,In_2707);
nor U2316 (N_2316,In_3529,N_1236);
and U2317 (N_2317,In_1374,In_1799);
nand U2318 (N_2318,N_1936,In_4746);
nor U2319 (N_2319,In_3895,In_1775);
or U2320 (N_2320,N_1589,N_876);
nand U2321 (N_2321,In_3620,N_1725);
nand U2322 (N_2322,In_442,N_1522);
or U2323 (N_2323,In_3466,N_1971);
or U2324 (N_2324,In_4491,N_1403);
nand U2325 (N_2325,N_1406,In_2295);
or U2326 (N_2326,In_1946,In_2530);
nand U2327 (N_2327,In_1863,In_824);
or U2328 (N_2328,In_2974,N_1613);
or U2329 (N_2329,N_1708,N_657);
nand U2330 (N_2330,In_2028,In_392);
xnor U2331 (N_2331,In_4902,N_1291);
and U2332 (N_2332,N_1101,N_1911);
xor U2333 (N_2333,In_4157,N_793);
or U2334 (N_2334,N_1636,In_4029);
nand U2335 (N_2335,In_2597,N_218);
nand U2336 (N_2336,In_4796,N_1987);
or U2337 (N_2337,N_1305,N_867);
or U2338 (N_2338,In_4738,In_184);
and U2339 (N_2339,In_3655,N_638);
xor U2340 (N_2340,In_1204,In_4237);
and U2341 (N_2341,In_2595,In_3347);
nand U2342 (N_2342,N_1596,N_1724);
xnor U2343 (N_2343,In_2249,In_2514);
nor U2344 (N_2344,In_1853,N_462);
nor U2345 (N_2345,N_651,In_2400);
or U2346 (N_2346,N_1026,N_1678);
nand U2347 (N_2347,N_1998,In_766);
xor U2348 (N_2348,N_1719,In_1965);
nor U2349 (N_2349,N_198,In_4185);
xnor U2350 (N_2350,N_177,N_1849);
nand U2351 (N_2351,N_1432,In_1147);
and U2352 (N_2352,N_1051,N_84);
xor U2353 (N_2353,N_116,In_26);
nand U2354 (N_2354,N_1134,N_114);
or U2355 (N_2355,N_1565,In_3772);
nand U2356 (N_2356,N_1978,In_2705);
and U2357 (N_2357,N_1052,In_2713);
or U2358 (N_2358,N_91,N_1711);
nor U2359 (N_2359,N_948,N_1238);
xnor U2360 (N_2360,In_3312,N_1764);
or U2361 (N_2361,N_1997,In_516);
nand U2362 (N_2362,N_1834,In_3018);
or U2363 (N_2363,N_1422,N_1754);
nor U2364 (N_2364,N_430,In_1236);
xor U2365 (N_2365,In_538,In_287);
or U2366 (N_2366,N_1560,In_4463);
nor U2367 (N_2367,N_1342,In_1765);
nor U2368 (N_2368,In_1435,In_2557);
nor U2369 (N_2369,In_29,N_1824);
xor U2370 (N_2370,In_767,In_3645);
and U2371 (N_2371,In_3163,N_1332);
nor U2372 (N_2372,N_1644,N_1485);
or U2373 (N_2373,In_164,N_1239);
nand U2374 (N_2374,In_4547,N_1964);
nor U2375 (N_2375,In_3531,In_79);
xnor U2376 (N_2376,In_325,In_3096);
nor U2377 (N_2377,In_2178,In_100);
nor U2378 (N_2378,N_1271,N_1345);
or U2379 (N_2379,N_994,N_1074);
xnor U2380 (N_2380,In_1178,N_760);
xnor U2381 (N_2381,In_3376,In_1813);
or U2382 (N_2382,N_849,N_1651);
nor U2383 (N_2383,N_879,N_473);
xnor U2384 (N_2384,In_3804,In_4802);
xnor U2385 (N_2385,In_4007,In_3778);
nand U2386 (N_2386,N_1117,N_1142);
or U2387 (N_2387,In_2256,In_935);
nor U2388 (N_2388,N_1566,N_1381);
or U2389 (N_2389,N_1456,N_281);
xnor U2390 (N_2390,N_1794,In_3182);
xor U2391 (N_2391,N_5,In_4033);
nor U2392 (N_2392,In_3364,In_220);
and U2393 (N_2393,N_1820,N_1197);
nand U2394 (N_2394,In_207,In_3896);
xnor U2395 (N_2395,N_380,In_1613);
or U2396 (N_2396,N_1270,In_1114);
or U2397 (N_2397,N_144,N_1815);
or U2398 (N_2398,In_2487,In_3000);
nand U2399 (N_2399,In_1123,In_4704);
and U2400 (N_2400,In_4497,In_3439);
nor U2401 (N_2401,N_463,In_603);
or U2402 (N_2402,N_1905,N_823);
nand U2403 (N_2403,N_906,N_1140);
nor U2404 (N_2404,In_1576,In_551);
and U2405 (N_2405,N_1156,In_2049);
and U2406 (N_2406,In_3186,N_1645);
and U2407 (N_2407,N_966,In_2765);
xnor U2408 (N_2408,In_2173,In_2977);
or U2409 (N_2409,In_2929,In_4732);
nand U2410 (N_2410,N_1104,N_1488);
and U2411 (N_2411,N_1956,N_1399);
xor U2412 (N_2412,In_155,N_26);
nand U2413 (N_2413,In_2001,N_417);
nand U2414 (N_2414,N_1541,In_3761);
and U2415 (N_2415,In_1752,N_1600);
or U2416 (N_2416,In_4702,In_4226);
or U2417 (N_2417,N_1714,N_1272);
nor U2418 (N_2418,In_1718,In_1487);
and U2419 (N_2419,N_1301,N_1400);
xor U2420 (N_2420,N_1172,N_1046);
nand U2421 (N_2421,In_799,In_1341);
and U2422 (N_2422,N_228,N_1647);
xor U2423 (N_2423,N_1470,N_1242);
xnor U2424 (N_2424,In_4635,N_1896);
nor U2425 (N_2425,In_2177,N_214);
or U2426 (N_2426,In_525,In_3595);
nor U2427 (N_2427,In_4929,N_757);
nor U2428 (N_2428,In_2930,In_4709);
xor U2429 (N_2429,In_933,N_1577);
or U2430 (N_2430,N_236,In_3105);
nor U2431 (N_2431,N_1213,N_1553);
and U2432 (N_2432,In_2245,In_2753);
and U2433 (N_2433,N_192,N_64);
nor U2434 (N_2434,In_1935,In_566);
xnor U2435 (N_2435,N_1108,N_1907);
xor U2436 (N_2436,N_1037,N_1353);
or U2437 (N_2437,In_3799,N_1160);
nor U2438 (N_2438,In_4899,N_1079);
nor U2439 (N_2439,In_128,In_1512);
xor U2440 (N_2440,In_2799,In_4207);
nor U2441 (N_2441,In_3081,N_239);
xnor U2442 (N_2442,In_1359,In_1850);
xor U2443 (N_2443,N_1377,N_509);
xnor U2444 (N_2444,N_886,In_2756);
and U2445 (N_2445,N_1506,N_1110);
nand U2446 (N_2446,In_3089,In_3460);
or U2447 (N_2447,N_1705,N_1548);
nor U2448 (N_2448,In_2161,In_2517);
or U2449 (N_2449,In_2155,N_1912);
or U2450 (N_2450,N_1829,N_788);
nor U2451 (N_2451,In_2971,N_623);
or U2452 (N_2452,In_3894,In_4881);
or U2453 (N_2453,In_2957,In_1188);
and U2454 (N_2454,N_1428,In_4833);
nor U2455 (N_2455,N_153,In_2023);
and U2456 (N_2456,N_1038,In_883);
and U2457 (N_2457,In_1600,In_1013);
nor U2458 (N_2458,N_333,N_296);
xnor U2459 (N_2459,N_1479,In_2426);
nor U2460 (N_2460,In_639,N_334);
or U2461 (N_2461,In_2109,In_4347);
xor U2462 (N_2462,N_1920,In_2659);
or U2463 (N_2463,In_1384,N_1451);
or U2464 (N_2464,N_1066,In_3638);
or U2465 (N_2465,N_329,In_930);
nand U2466 (N_2466,N_1646,In_3791);
or U2467 (N_2467,In_1593,N_1136);
xnor U2468 (N_2468,N_1848,N_1856);
xnor U2469 (N_2469,In_40,N_1392);
and U2470 (N_2470,In_763,N_965);
and U2471 (N_2471,In_4775,In_4530);
nor U2472 (N_2472,N_1372,N_1750);
nor U2473 (N_2473,N_820,In_850);
xor U2474 (N_2474,N_579,In_3227);
and U2475 (N_2475,N_1253,In_1768);
and U2476 (N_2476,In_1550,N_1628);
nand U2477 (N_2477,N_1830,In_4418);
or U2478 (N_2478,In_2539,In_3171);
nand U2479 (N_2479,N_394,N_735);
xnor U2480 (N_2480,N_1763,In_4344);
and U2481 (N_2481,N_1928,In_1465);
xnor U2482 (N_2482,In_1028,N_547);
nor U2483 (N_2483,N_1884,N_1550);
nand U2484 (N_2484,In_1978,N_1620);
and U2485 (N_2485,In_1955,In_253);
xnor U2486 (N_2486,N_1735,N_658);
nor U2487 (N_2487,N_1945,N_1637);
nor U2488 (N_2488,In_3824,N_878);
or U2489 (N_2489,In_107,In_4858);
nor U2490 (N_2490,In_364,In_564);
or U2491 (N_2491,In_2808,In_1847);
nand U2492 (N_2492,In_4453,N_419);
nand U2493 (N_2493,N_1365,In_4244);
nand U2494 (N_2494,In_1491,N_1123);
nand U2495 (N_2495,N_790,N_1921);
xor U2496 (N_2496,N_303,In_1874);
or U2497 (N_2497,N_1497,In_2685);
nand U2498 (N_2498,N_1967,In_1996);
nor U2499 (N_2499,N_973,N_1514);
or U2500 (N_2500,In_4458,N_1075);
nor U2501 (N_2501,In_1629,In_2654);
xnor U2502 (N_2502,N_1910,N_58);
nand U2503 (N_2503,In_1885,N_101);
or U2504 (N_2504,In_4500,N_1944);
nor U2505 (N_2505,In_2668,In_734);
and U2506 (N_2506,N_922,N_1690);
xnor U2507 (N_2507,N_566,N_815);
nand U2508 (N_2508,N_1975,N_195);
xor U2509 (N_2509,In_1189,In_465);
and U2510 (N_2510,In_865,N_802);
nand U2511 (N_2511,N_1675,N_677);
or U2512 (N_2512,In_4787,In_4589);
nand U2513 (N_2513,N_1080,In_2647);
and U2514 (N_2514,In_2146,N_1761);
xnor U2515 (N_2515,N_1073,In_3344);
nand U2516 (N_2516,N_1020,In_4756);
nor U2517 (N_2517,In_4402,N_1427);
nor U2518 (N_2518,N_1366,N_1036);
nor U2519 (N_2519,N_1055,N_1962);
nor U2520 (N_2520,In_713,In_2098);
or U2521 (N_2521,In_936,In_1199);
and U2522 (N_2522,In_971,In_661);
xor U2523 (N_2523,N_309,N_1658);
xor U2524 (N_2524,N_1181,N_1034);
xnor U2525 (N_2525,In_630,N_999);
or U2526 (N_2526,In_1247,In_803);
nand U2527 (N_2527,In_4149,N_1759);
nor U2528 (N_2528,In_2884,N_709);
and U2529 (N_2529,N_1067,N_1012);
nand U2530 (N_2530,In_4394,In_2321);
nand U2531 (N_2531,In_2686,N_1722);
and U2532 (N_2532,N_1559,In_1164);
xnor U2533 (N_2533,In_4697,N_1462);
nor U2534 (N_2534,In_4325,N_1268);
and U2535 (N_2535,N_1499,In_1428);
and U2536 (N_2536,In_841,N_1476);
and U2537 (N_2537,In_4145,In_3101);
nand U2538 (N_2538,N_1107,N_290);
nor U2539 (N_2539,In_887,N_1401);
xnor U2540 (N_2540,In_350,N_1394);
nand U2541 (N_2541,N_1991,In_3398);
nand U2542 (N_2542,N_1940,In_4416);
xor U2543 (N_2543,N_1556,N_1699);
nand U2544 (N_2544,In_3042,In_56);
nand U2545 (N_2545,N_418,N_612);
nor U2546 (N_2546,N_1371,N_172);
or U2547 (N_2547,In_1536,In_2606);
xnor U2548 (N_2548,In_2226,In_47);
nand U2549 (N_2549,N_1733,In_3271);
xnor U2550 (N_2550,N_1405,In_793);
nand U2551 (N_2551,N_1343,N_1851);
xor U2552 (N_2552,N_980,N_673);
nand U2553 (N_2553,In_3626,In_4846);
or U2554 (N_2554,N_1622,N_961);
or U2555 (N_2555,In_606,N_1091);
xor U2556 (N_2556,In_1379,N_1621);
xor U2557 (N_2557,In_4758,In_1822);
and U2558 (N_2558,In_4397,In_565);
and U2559 (N_2559,N_743,N_1859);
or U2560 (N_2560,N_1895,N_1611);
and U2561 (N_2561,In_1078,In_1306);
nand U2562 (N_2562,N_703,N_191);
nand U2563 (N_2563,N_1164,N_226);
xnor U2564 (N_2564,In_3302,N_1654);
or U2565 (N_2565,N_1623,N_340);
nand U2566 (N_2566,In_4856,In_951);
nor U2567 (N_2567,N_526,In_1972);
or U2568 (N_2568,In_576,N_548);
xor U2569 (N_2569,N_244,In_4221);
or U2570 (N_2570,N_254,In_2653);
nand U2571 (N_2571,N_1230,In_3870);
xor U2572 (N_2572,N_382,In_1057);
and U2573 (N_2573,N_1822,N_1520);
nor U2574 (N_2574,N_1869,N_633);
nand U2575 (N_2575,In_3111,In_1671);
or U2576 (N_2576,In_3833,In_4823);
or U2577 (N_2577,In_4644,N_943);
xnor U2578 (N_2578,In_4786,In_2417);
xnor U2579 (N_2579,In_2518,In_2357);
nor U2580 (N_2580,In_4389,In_1828);
or U2581 (N_2581,N_168,N_996);
xor U2582 (N_2582,N_1630,In_4619);
nor U2583 (N_2583,In_1864,N_1384);
or U2584 (N_2584,N_1701,N_1835);
nand U2585 (N_2585,In_186,N_871);
or U2586 (N_2586,N_307,In_1566);
or U2587 (N_2587,N_1858,N_78);
xor U2588 (N_2588,N_491,In_2770);
and U2589 (N_2589,N_1147,In_4401);
or U2590 (N_2590,In_3898,In_1538);
nand U2591 (N_2591,In_3220,N_1840);
xor U2592 (N_2592,N_88,N_1318);
and U2593 (N_2593,N_1347,N_1983);
nor U2594 (N_2594,N_328,In_2158);
nor U2595 (N_2595,In_527,N_1585);
xnor U2596 (N_2596,N_787,N_1673);
nand U2597 (N_2597,In_552,N_1150);
xnor U2598 (N_2598,In_4213,In_1518);
or U2599 (N_2599,N_1358,N_710);
or U2600 (N_2600,In_1531,In_3687);
or U2601 (N_2601,In_1732,In_868);
nand U2602 (N_2602,N_1706,N_1558);
nor U2603 (N_2603,N_1938,In_3442);
or U2604 (N_2604,In_1383,N_1265);
nor U2605 (N_2605,N_1527,In_2579);
or U2606 (N_2606,N_349,N_826);
xor U2607 (N_2607,N_1665,In_4114);
nand U2608 (N_2608,N_514,N_1811);
nand U2609 (N_2609,N_123,N_445);
or U2610 (N_2610,N_125,N_1583);
or U2611 (N_2611,N_1165,In_2461);
and U2612 (N_2612,In_1230,N_1874);
nand U2613 (N_2613,In_2122,N_1900);
xor U2614 (N_2614,In_925,N_1257);
and U2615 (N_2615,N_1085,In_4102);
or U2616 (N_2616,N_1457,In_2504);
nand U2617 (N_2617,In_140,N_1289);
xnor U2618 (N_2618,In_3864,In_2042);
nand U2619 (N_2619,In_4886,N_1389);
nor U2620 (N_2620,In_1125,In_2625);
nor U2621 (N_2621,In_4749,In_2222);
xnor U2622 (N_2622,N_1065,N_1349);
or U2623 (N_2623,N_1810,N_1813);
and U2624 (N_2624,In_4109,In_1449);
nand U2625 (N_2625,In_561,N_720);
nor U2626 (N_2626,In_3787,N_1414);
and U2627 (N_2627,In_460,In_3691);
nor U2628 (N_2628,N_315,N_136);
nand U2629 (N_2629,In_3033,In_2315);
xor U2630 (N_2630,N_1563,N_1280);
and U2631 (N_2631,N_352,In_2344);
nor U2632 (N_2632,In_1588,In_676);
nand U2633 (N_2633,In_4828,N_243);
nor U2634 (N_2634,N_127,N_1390);
and U2635 (N_2635,N_1249,In_313);
nand U2636 (N_2636,N_1126,N_1790);
or U2637 (N_2637,N_756,N_410);
nor U2638 (N_2638,In_2709,In_4470);
or U2639 (N_2639,In_4872,N_1844);
and U2640 (N_2640,In_4862,N_778);
and U2641 (N_2641,N_1391,N_1843);
and U2642 (N_2642,In_1132,N_1561);
nand U2643 (N_2643,In_1360,N_630);
nor U2644 (N_2644,N_1304,N_294);
nor U2645 (N_2645,In_1337,In_3017);
xnor U2646 (N_2646,In_1344,N_346);
nor U2647 (N_2647,In_1764,N_1395);
nor U2648 (N_2648,N_342,In_3934);
or U2649 (N_2649,N_1420,In_3739);
nand U2650 (N_2650,In_3594,N_1818);
and U2651 (N_2651,N_705,In_657);
nand U2652 (N_2652,In_4283,N_1686);
nand U2653 (N_2653,N_1298,N_285);
or U2654 (N_2654,N_1269,In_4112);
or U2655 (N_2655,In_784,N_1741);
and U2656 (N_2656,N_882,N_1639);
and U2657 (N_2657,N_1208,In_421);
xor U2658 (N_2658,N_1247,N_120);
or U2659 (N_2659,In_4350,In_1000);
xnor U2660 (N_2660,N_483,In_1788);
and U2661 (N_2661,N_51,N_1503);
and U2662 (N_2662,In_3711,N_459);
and U2663 (N_2663,N_1715,N_1035);
nor U2664 (N_2664,In_3279,In_986);
nor U2665 (N_2665,In_2988,In_4154);
and U2666 (N_2666,N_668,In_718);
and U2667 (N_2667,In_4268,In_4585);
nor U2668 (N_2668,In_1463,N_597);
nand U2669 (N_2669,In_4364,N_1720);
or U2670 (N_2670,In_1774,In_148);
nand U2671 (N_2671,In_916,N_576);
or U2672 (N_2672,In_1272,In_3471);
or U2673 (N_2673,In_49,In_3586);
or U2674 (N_2674,N_1376,In_4996);
nor U2675 (N_2675,N_1626,In_2962);
and U2676 (N_2676,In_1568,In_4966);
xnor U2677 (N_2677,N_216,In_1294);
nand U2678 (N_2678,N_1388,In_3578);
or U2679 (N_2679,N_1446,In_2807);
xor U2680 (N_2680,In_682,N_1661);
nor U2681 (N_2681,In_4508,N_402);
nand U2682 (N_2682,N_1130,N_1712);
or U2683 (N_2683,In_23,In_4212);
nor U2684 (N_2684,In_3298,In_3061);
and U2685 (N_2685,In_3975,N_1716);
or U2686 (N_2686,N_1765,N_1286);
and U2687 (N_2687,In_687,In_3731);
xor U2688 (N_2688,In_4757,In_4945);
or U2689 (N_2689,In_2148,N_936);
nor U2690 (N_2690,N_92,In_3997);
nand U2691 (N_2691,In_536,In_1527);
and U2692 (N_2692,In_1509,In_2903);
and U2693 (N_2693,N_1693,N_1816);
nor U2694 (N_2694,In_371,In_2185);
and U2695 (N_2695,In_1495,N_440);
and U2696 (N_2696,N_1994,N_869);
nand U2697 (N_2697,N_1162,N_1198);
nand U2698 (N_2698,N_1726,In_847);
nand U2699 (N_2699,N_1317,N_1295);
or U2700 (N_2700,N_1587,In_4236);
xor U2701 (N_2701,In_1403,In_4473);
or U2702 (N_2702,N_185,N_1109);
and U2703 (N_2703,In_4734,In_276);
nor U2704 (N_2704,N_816,In_2755);
and U2705 (N_2705,In_839,N_1303);
nor U2706 (N_2706,N_1122,In_1295);
nor U2707 (N_2707,N_1823,In_2488);
or U2708 (N_2708,N_55,In_4175);
or U2709 (N_2709,In_250,In_1064);
and U2710 (N_2710,In_4759,In_3273);
and U2711 (N_2711,In_2801,In_1958);
xnor U2712 (N_2712,In_386,N_1846);
and U2713 (N_2713,N_1060,In_2687);
xnor U2714 (N_2714,N_1228,N_1576);
xor U2715 (N_2715,In_4868,In_2100);
nand U2716 (N_2716,In_1475,N_1713);
and U2717 (N_2717,N_670,N_1307);
nor U2718 (N_2718,In_3889,In_4750);
and U2719 (N_2719,In_4338,In_1724);
nand U2720 (N_2720,N_1374,N_40);
or U2721 (N_2721,N_1493,In_435);
and U2722 (N_2722,In_384,In_1921);
and U2723 (N_2723,N_249,N_1993);
and U2724 (N_2724,N_1828,N_1019);
nand U2725 (N_2725,N_777,In_1124);
xor U2726 (N_2726,In_3572,In_2702);
xnor U2727 (N_2727,N_1788,N_1312);
xnor U2728 (N_2728,In_823,In_4579);
nor U2729 (N_2729,In_76,In_3917);
or U2730 (N_2730,In_800,In_3958);
nor U2731 (N_2731,N_1125,N_1736);
or U2732 (N_2732,In_1103,In_3590);
nand U2733 (N_2733,In_876,In_3696);
nor U2734 (N_2734,In_4065,In_2882);
nand U2735 (N_2735,In_4830,In_3981);
nand U2736 (N_2736,N_1157,N_1989);
and U2737 (N_2737,In_1616,N_112);
nand U2738 (N_2738,In_1833,In_1311);
nand U2739 (N_2739,N_530,N_1283);
nand U2740 (N_2740,In_3040,N_605);
or U2741 (N_2741,In_1464,N_517);
and U2742 (N_2742,N_48,N_1694);
xor U2743 (N_2743,In_4308,N_1753);
nand U2744 (N_2744,In_4907,In_2955);
or U2745 (N_2745,N_1568,In_4019);
and U2746 (N_2746,In_3522,N_972);
xnor U2747 (N_2747,N_1158,In_854);
nor U2748 (N_2748,In_3698,N_1883);
nor U2749 (N_2749,N_106,In_1340);
or U2750 (N_2750,In_4954,In_2715);
nand U2751 (N_2751,In_3835,N_1293);
nor U2752 (N_2752,N_935,N_437);
nor U2753 (N_2753,N_1031,In_1455);
nand U2754 (N_2754,N_1942,N_1515);
and U2755 (N_2755,In_2781,N_374);
nand U2756 (N_2756,N_881,N_1697);
or U2757 (N_2757,In_2484,In_45);
or U2758 (N_2758,In_744,In_3613);
nand U2759 (N_2759,In_2320,In_668);
and U2760 (N_2760,In_4211,N_121);
and U2761 (N_2761,N_1128,N_828);
and U2762 (N_2762,In_3897,N_456);
nor U2763 (N_2763,N_1730,N_1633);
or U2764 (N_2764,In_3315,N_905);
xnor U2765 (N_2765,In_2555,N_263);
nand U2766 (N_2766,In_4197,N_582);
or U2767 (N_2767,N_1161,N_1572);
xor U2768 (N_2768,N_1378,In_1241);
nand U2769 (N_2769,N_1649,N_643);
xor U2770 (N_2770,In_2910,In_3902);
nand U2771 (N_2771,In_717,N_1908);
nand U2772 (N_2772,N_589,N_1260);
and U2773 (N_2773,In_2885,N_82);
nand U2774 (N_2774,N_1523,N_655);
nand U2775 (N_2775,In_2232,N_880);
nor U2776 (N_2776,N_696,N_1996);
xor U2777 (N_2777,In_4115,In_3306);
xnor U2778 (N_2778,N_827,N_1924);
xor U2779 (N_2779,In_16,In_899);
nand U2780 (N_2780,In_499,N_1662);
or U2781 (N_2781,In_1135,In_749);
nand U2782 (N_2782,N_159,In_1063);
xnor U2783 (N_2783,In_3019,In_2716);
and U2784 (N_2784,In_2916,N_1294);
nand U2785 (N_2785,N_1676,N_1017);
nor U2786 (N_2786,N_87,In_2810);
nor U2787 (N_2787,In_199,In_2332);
xor U2788 (N_2788,N_1494,N_232);
nor U2789 (N_2789,In_2154,N_385);
nor U2790 (N_2790,In_2855,N_635);
xnor U2791 (N_2791,N_1870,N_1787);
or U2792 (N_2792,In_4967,N_897);
and U2793 (N_2793,N_1973,N_102);
nand U2794 (N_2794,N_1878,In_2746);
or U2795 (N_2795,N_230,In_1926);
nand U2796 (N_2796,N_412,In_759);
nand U2797 (N_2797,In_1081,In_4510);
and U2798 (N_2798,N_1624,N_261);
nand U2799 (N_2799,N_863,N_1216);
nor U2800 (N_2800,N_267,N_1871);
nor U2801 (N_2801,In_3333,N_751);
xor U2802 (N_2802,In_1210,N_1429);
nand U2803 (N_2803,N_1684,In_2803);
or U2804 (N_2804,In_2041,In_967);
and U2805 (N_2805,In_2024,In_4813);
nand U2806 (N_2806,In_3528,N_1373);
or U2807 (N_2807,In_2945,N_1882);
or U2808 (N_2808,N_1709,N_487);
xor U2809 (N_2809,N_1718,N_727);
nor U2810 (N_2810,N_1175,N_1423);
or U2811 (N_2811,N_1837,In_3295);
nor U2812 (N_2812,In_2490,In_3555);
xor U2813 (N_2813,In_1250,N_1839);
nand U2814 (N_2814,In_1891,N_1119);
nor U2815 (N_2815,In_2284,In_2764);
and U2816 (N_2816,In_110,N_1227);
nor U2817 (N_2817,In_4080,N_1155);
and U2818 (N_2818,N_959,In_196);
nand U2819 (N_2819,N_1664,In_2304);
xnor U2820 (N_2820,In_2440,N_1703);
xnor U2821 (N_2821,In_180,In_398);
or U2822 (N_2822,N_546,In_4922);
and U2823 (N_2823,In_1790,N_1968);
nand U2824 (N_2824,N_245,In_4600);
and U2825 (N_2825,N_1263,N_780);
or U2826 (N_2826,In_529,N_997);
nand U2827 (N_2827,N_1141,N_1098);
and U2828 (N_2828,In_348,In_1126);
nor U2829 (N_2829,In_1086,N_1616);
nand U2830 (N_2830,N_808,In_3965);
and U2831 (N_2831,In_4425,In_2431);
nand U2832 (N_2832,In_4557,N_1159);
or U2833 (N_2833,N_1862,N_50);
and U2834 (N_2834,N_280,N_1350);
nor U2835 (N_2835,N_896,N_1760);
nor U2836 (N_2836,N_1354,In_2619);
nor U2837 (N_2837,In_187,In_57);
nor U2838 (N_2838,N_1893,N_126);
xor U2839 (N_2839,N_1203,N_62);
xnor U2840 (N_2840,In_4841,In_4117);
and U2841 (N_2841,N_1014,In_667);
and U2842 (N_2842,In_4739,In_311);
nor U2843 (N_2843,N_282,N_1801);
nor U2844 (N_2844,In_4405,In_227);
or U2845 (N_2845,N_1960,In_4573);
nand U2846 (N_2846,In_3304,In_3963);
nand U2847 (N_2847,N_1452,N_903);
xnor U2848 (N_2848,N_1219,In_3139);
and U2849 (N_2849,In_3520,N_1707);
xor U2850 (N_2850,N_1875,N_1807);
nand U2851 (N_2851,N_1751,N_704);
or U2852 (N_2852,N_1925,N_1511);
xnor U2853 (N_2853,In_1017,N_223);
xor U2854 (N_2854,N_1510,In_2314);
xnor U2855 (N_2855,In_68,In_3069);
nand U2856 (N_2856,In_3015,In_73);
xnor U2857 (N_2857,N_795,In_4271);
xnor U2858 (N_2858,In_625,N_495);
nand U2859 (N_2859,N_581,N_1868);
or U2860 (N_2860,In_4171,In_1321);
and U2861 (N_2861,In_3384,In_507);
xnor U2862 (N_2862,In_4955,N_1054);
nor U2863 (N_2863,N_1437,N_1328);
nor U2864 (N_2864,N_1821,N_1657);
xor U2865 (N_2865,In_3762,N_1490);
and U2866 (N_2866,In_4104,In_1313);
and U2867 (N_2867,N_1088,N_229);
nor U2868 (N_2868,In_4544,N_1169);
or U2869 (N_2869,N_1582,In_689);
and U2870 (N_2870,N_708,N_1421);
xnor U2871 (N_2871,In_1609,In_27);
xor U2872 (N_2872,In_4776,In_586);
or U2873 (N_2873,N_1770,In_145);
nor U2874 (N_2874,In_1611,N_784);
nor U2875 (N_2875,N_1808,In_1658);
nor U2876 (N_2876,In_2047,In_2452);
and U2877 (N_2877,In_2095,N_1757);
and U2878 (N_2878,In_695,In_191);
xor U2879 (N_2879,In_4246,In_258);
xnor U2880 (N_2880,N_1922,In_827);
or U2881 (N_2881,N_1867,N_472);
xnor U2882 (N_2882,In_1664,In_2159);
and U2883 (N_2883,In_4167,N_1891);
xnor U2884 (N_2884,N_1546,N_1408);
and U2885 (N_2885,In_2191,N_852);
or U2886 (N_2886,In_572,In_142);
nand U2887 (N_2887,In_815,In_4150);
and U2888 (N_2888,N_931,In_646);
xor U2889 (N_2889,N_1370,N_1042);
nand U2890 (N_2890,N_883,In_2871);
and U2891 (N_2891,In_968,In_1062);
nor U2892 (N_2892,N_137,In_3585);
nor U2893 (N_2893,In_4679,N_1889);
nand U2894 (N_2894,In_4534,In_330);
and U2895 (N_2895,In_147,In_3387);
nand U2896 (N_2896,In_222,In_1363);
or U2897 (N_2897,In_2483,N_1474);
nor U2898 (N_2898,In_1264,N_384);
or U2899 (N_2899,N_405,N_1171);
or U2900 (N_2900,N_1660,N_967);
and U2901 (N_2901,In_3167,In_3932);
nor U2902 (N_2902,In_32,In_2200);
nand U2903 (N_2903,N_1826,N_1338);
or U2904 (N_2904,N_1190,N_353);
or U2905 (N_2905,N_1817,In_4539);
or U2906 (N_2906,N_1831,N_1986);
nor U2907 (N_2907,In_464,N_1352);
and U2908 (N_2908,N_1948,N_848);
and U2909 (N_2909,In_218,In_1051);
or U2910 (N_2910,N_898,N_728);
or U2911 (N_2911,In_889,N_8);
or U2912 (N_2912,In_4291,N_1659);
or U2913 (N_2913,In_728,N_707);
nand U2914 (N_2914,In_3184,N_1591);
and U2915 (N_2915,N_1595,In_3802);
and U2916 (N_2916,In_1887,N_955);
xor U2917 (N_2917,In_444,In_3985);
xnor U2918 (N_2918,In_4873,In_283);
and U2919 (N_2919,N_1482,N_1226);
xor U2920 (N_2920,N_1173,N_1502);
nor U2921 (N_2921,N_723,N_308);
xor U2922 (N_2922,N_111,N_1581);
or U2923 (N_2923,In_21,N_1415);
and U2924 (N_2924,In_3192,N_86);
and U2925 (N_2925,N_235,N_1082);
xor U2926 (N_2926,N_1471,N_1507);
nor U2927 (N_2927,N_1916,N_49);
and U2928 (N_2928,N_1683,N_1923);
or U2929 (N_2929,N_1774,In_2050);
nor U2930 (N_2930,N_1532,In_1894);
and U2931 (N_2931,In_1492,N_976);
and U2932 (N_2932,N_1913,In_2621);
and U2933 (N_2933,In_3050,In_4335);
xor U2934 (N_2934,In_3918,In_2435);
xor U2935 (N_2935,In_2396,N_1981);
xnor U2936 (N_2936,N_365,In_493);
xnor U2937 (N_2937,In_2609,N_1894);
or U2938 (N_2938,In_3624,N_1508);
xnor U2939 (N_2939,In_4834,In_3532);
or U2940 (N_2940,In_1635,In_3177);
or U2941 (N_2941,In_2535,In_251);
nor U2942 (N_2942,In_59,N_1982);
and U2943 (N_2943,In_2912,In_2943);
nor U2944 (N_2944,N_1855,N_211);
xor U2945 (N_2945,In_670,In_4293);
xor U2946 (N_2946,N_940,N_392);
and U2947 (N_2947,In_411,In_4627);
or U2948 (N_2948,In_1077,In_122);
nor U2949 (N_2949,N_937,In_3869);
and U2950 (N_2950,N_302,N_16);
xnor U2951 (N_2951,N_1477,In_3830);
xnor U2952 (N_2952,N_1857,In_4785);
and U2953 (N_2953,In_1973,In_3540);
nand U2954 (N_2954,In_4673,In_3056);
nor U2955 (N_2955,N_1496,In_3821);
xor U2956 (N_2956,N_1212,N_1297);
xnor U2957 (N_2957,N_1885,N_1652);
and U2958 (N_2958,N_1930,N_1375);
xnor U2959 (N_2959,N_1285,N_1279);
xor U2960 (N_2960,N_28,N_1329);
or U2961 (N_2961,In_1898,N_1555);
nor U2962 (N_2962,N_1917,N_1148);
xor U2963 (N_2963,In_4623,In_3106);
nand U2964 (N_2964,In_3893,In_136);
nor U2965 (N_2965,N_1223,N_1995);
and U2966 (N_2966,In_370,N_170);
or U2967 (N_2967,N_375,In_194);
nand U2968 (N_2968,N_754,N_1483);
and U2969 (N_2969,In_333,N_857);
nor U2970 (N_2970,In_4962,N_1500);
xnor U2971 (N_2971,N_1791,N_1619);
nor U2972 (N_2972,In_2954,N_1145);
nand U2973 (N_2973,N_1355,N_204);
and U2974 (N_2974,N_1685,In_2289);
or U2975 (N_2975,N_1431,In_2744);
xnor U2976 (N_2976,In_3296,In_2384);
and U2977 (N_2977,N_1094,N_1850);
and U2978 (N_2978,N_1610,In_2430);
and U2979 (N_2979,In_1361,N_1902);
xnor U2980 (N_2980,N_359,In_545);
nor U2981 (N_2981,N_1692,In_3103);
and U2982 (N_2982,In_638,N_607);
or U2983 (N_2983,N_291,N_1618);
nor U2984 (N_2984,In_4240,In_2341);
and U2985 (N_2985,N_1364,In_4013);
nor U2986 (N_2986,N_1047,N_1410);
xor U2987 (N_2987,N_887,N_118);
or U2988 (N_2988,N_1233,N_1903);
nand U2989 (N_2989,In_3278,N_1833);
and U2990 (N_2990,In_1120,In_4805);
or U2991 (N_2991,N_1918,In_2477);
or U2992 (N_2992,In_1416,In_2728);
or U2993 (N_2993,N_1193,In_3564);
and U2994 (N_2994,In_4999,In_3998);
or U2995 (N_2995,In_322,N_506);
nand U2996 (N_2996,In_2714,N_1881);
nor U2997 (N_2997,N_1778,In_177);
xnor U2998 (N_2998,In_2727,N_915);
nor U2999 (N_2999,In_1678,In_2589);
xor U3000 (N_3000,In_2587,N_2191);
or U3001 (N_3001,N_2718,N_2187);
nor U3002 (N_3002,N_1594,In_688);
or U3003 (N_3003,N_2937,N_2810);
and U3004 (N_3004,In_4617,N_2279);
or U3005 (N_3005,N_2915,N_1049);
xor U3006 (N_3006,N_2401,In_502);
xnor U3007 (N_3007,N_2498,N_831);
xor U3008 (N_3008,In_4189,N_2665);
or U3009 (N_3009,In_3005,N_2836);
and U3010 (N_3010,N_1535,N_1450);
xnor U3011 (N_3011,N_2411,N_2041);
xor U3012 (N_3012,In_3782,N_1313);
and U3013 (N_3013,In_2983,N_2595);
nand U3014 (N_3014,N_2701,In_3461);
nor U3015 (N_3015,In_3367,N_2061);
and U3016 (N_3016,N_2634,N_2102);
and U3017 (N_3017,N_2643,N_1877);
or U3018 (N_3018,N_2824,In_1215);
or U3019 (N_3019,N_1383,N_2173);
xor U3020 (N_3020,N_1536,N_2576);
xor U3021 (N_3021,N_480,N_1597);
nor U3022 (N_3022,In_4005,N_2787);
xnor U3023 (N_3023,N_2543,N_2329);
nand U3024 (N_3024,N_119,N_2039);
xnor U3025 (N_3025,N_1688,N_2563);
nand U3026 (N_3026,N_2302,N_1039);
and U3027 (N_3027,N_2445,In_637);
nand U3028 (N_3028,N_1044,N_2670);
nor U3029 (N_3029,N_2094,N_2831);
nor U3030 (N_3030,In_241,N_2929);
or U3031 (N_3031,In_2618,N_2327);
nand U3032 (N_3032,N_2381,N_1320);
xor U3033 (N_3033,In_4848,In_4692);
xnor U3034 (N_3034,N_2351,In_1167);
xor U3035 (N_3035,N_2172,N_2713);
or U3036 (N_3036,N_2660,N_1517);
or U3037 (N_3037,In_393,N_2141);
nand U3038 (N_3038,N_2273,N_2434);
nand U3039 (N_3039,N_2516,N_2507);
nor U3040 (N_3040,N_2520,N_1564);
and U3041 (N_3041,N_2237,N_2842);
and U3042 (N_3042,N_2571,In_679);
xnor U3043 (N_3043,N_1480,In_1952);
xor U3044 (N_3044,N_2573,N_2437);
and U3045 (N_3045,N_2878,N_2217);
nor U3046 (N_3046,N_2201,N_2154);
nor U3047 (N_3047,N_1528,N_2422);
nand U3048 (N_3048,In_4061,In_2333);
nor U3049 (N_3049,In_3161,In_4487);
nor U3050 (N_3050,In_512,N_2231);
or U3051 (N_3051,N_2555,N_1640);
nand U3052 (N_3052,In_2106,In_812);
nor U3053 (N_3053,N_2879,N_2916);
nor U3054 (N_3054,N_2817,N_2835);
xnor U3055 (N_3055,N_2129,N_1206);
and U3056 (N_3056,In_3836,N_454);
and U3057 (N_3057,N_2751,N_2234);
or U3058 (N_3058,N_276,N_2250);
nand U3059 (N_3059,N_1369,N_683);
nand U3060 (N_3060,In_2277,N_2823);
or U3061 (N_3061,N_2395,In_115);
or U3062 (N_3062,N_179,N_769);
xnor U3063 (N_3063,N_2865,N_2413);
and U3064 (N_3064,In_2856,In_1728);
nand U3065 (N_3065,N_1653,N_2448);
nand U3066 (N_3066,In_4449,N_1886);
nor U3067 (N_3067,N_2305,In_3642);
and U3068 (N_3068,N_998,N_1207);
nor U3069 (N_3069,N_2248,N_1866);
nor U3070 (N_3070,N_2761,N_520);
nand U3071 (N_3071,N_1398,N_2006);
xor U3072 (N_3072,N_2811,N_2236);
nor U3073 (N_3073,N_2615,N_2648);
xnor U3074 (N_3074,N_2574,N_2725);
xnor U3075 (N_3075,In_3118,N_1439);
nor U3076 (N_3076,In_2644,N_20);
nand U3077 (N_3077,In_1634,N_2075);
and U3078 (N_3078,In_1054,N_2745);
nand U3079 (N_3079,N_2923,N_2085);
and U3080 (N_3080,N_1976,N_2024);
nor U3081 (N_3081,In_3639,N_2209);
nor U3082 (N_3082,In_4611,In_2934);
nand U3083 (N_3083,N_2832,N_2055);
and U3084 (N_3084,N_2051,N_2157);
xor U3085 (N_3085,In_890,In_2394);
nand U3086 (N_3086,In_2936,N_2802);
nand U3087 (N_3087,N_1087,N_2686);
or U3088 (N_3088,N_588,N_2876);
or U3089 (N_3089,N_2944,N_2928);
or U3090 (N_3090,N_2506,N_1970);
xor U3091 (N_3091,N_2920,N_810);
xor U3092 (N_3092,In_2164,N_2440);
nand U3093 (N_3093,N_861,N_553);
nand U3094 (N_3094,N_2753,N_2567);
nand U3095 (N_3095,N_1105,N_1040);
or U3096 (N_3096,N_2330,N_2957);
nand U3097 (N_3097,N_1744,In_3193);
nand U3098 (N_3098,N_1737,N_1435);
and U3099 (N_3099,N_2796,In_1597);
xor U3100 (N_3100,N_1838,N_2511);
nand U3101 (N_3101,N_2277,N_2941);
xnor U3102 (N_3102,N_1845,In_3513);
nor U3103 (N_3103,N_1234,N_2491);
or U3104 (N_3104,N_776,N_2599);
nand U3105 (N_3105,In_4257,N_2866);
xnor U3106 (N_3106,In_1901,N_2949);
nor U3107 (N_3107,N_2793,N_2123);
or U3108 (N_3108,N_2292,In_2206);
xor U3109 (N_3109,N_2240,N_2142);
xnor U3110 (N_3110,N_406,In_3057);
or U3111 (N_3111,N_2453,In_4523);
and U3112 (N_3112,N_2977,N_2334);
and U3113 (N_3113,In_3675,In_3618);
or U3114 (N_3114,In_2044,N_1005);
xor U3115 (N_3115,N_1861,N_2781);
nand U3116 (N_3116,N_2698,N_2723);
nand U3117 (N_3117,N_2553,N_2467);
or U3118 (N_3118,N_2961,N_2077);
nor U3119 (N_3119,In_1073,In_3569);
nand U3120 (N_3120,In_3237,In_539);
nand U3121 (N_3121,N_2103,N_1192);
nor U3122 (N_3122,N_2729,N_2451);
nand U3123 (N_3123,In_4130,N_1949);
xor U3124 (N_3124,N_1670,N_682);
xor U3125 (N_3125,N_2286,N_1612);
and U3126 (N_3126,In_3158,In_4535);
nand U3127 (N_3127,In_783,In_1289);
nand U3128 (N_3128,N_2073,N_1152);
nand U3129 (N_3129,N_1863,N_2748);
xnor U3130 (N_3130,N_2684,N_1057);
xnor U3131 (N_3131,In_2451,In_3629);
xnor U3132 (N_3132,N_2934,N_2825);
nor U3133 (N_3133,N_2689,N_2795);
nand U3134 (N_3134,N_2387,In_3722);
nand U3135 (N_3135,N_2532,N_2518);
nor U3136 (N_3136,In_3716,N_1784);
or U3137 (N_3137,In_1411,N_2079);
and U3138 (N_3138,N_817,In_2969);
xor U3139 (N_3139,N_2220,N_1671);
xor U3140 (N_3140,N_2140,In_2322);
xnor U3141 (N_3141,In_1939,N_1954);
and U3142 (N_3142,N_2295,In_4976);
nor U3143 (N_3143,N_1359,In_4532);
and U3144 (N_3144,N_2497,N_1326);
or U3145 (N_3145,N_1898,N_2486);
nand U3146 (N_3146,N_2890,N_438);
nor U3147 (N_3147,N_2343,In_2692);
nor U3148 (N_3148,N_1100,In_1948);
xor U3149 (N_3149,N_2534,In_2566);
xor U3150 (N_3150,N_330,N_2303);
and U3151 (N_3151,In_3964,N_2042);
nor U3152 (N_3152,N_10,N_2537);
nand U3153 (N_3153,N_1766,N_443);
nand U3154 (N_3154,N_2913,N_2827);
or U3155 (N_3155,N_2533,N_2531);
nor U3156 (N_3156,N_2312,N_2025);
or U3157 (N_3157,N_2695,N_2671);
nand U3158 (N_3158,N_2225,N_2180);
and U3159 (N_3159,N_2444,N_2148);
nor U3160 (N_3160,N_2526,N_2114);
xnor U3161 (N_3161,N_1935,N_2956);
nor U3162 (N_3162,N_2134,N_685);
nand U3163 (N_3163,N_2251,N_2710);
xnor U3164 (N_3164,N_2580,In_2425);
nand U3165 (N_3165,N_1634,N_2262);
nand U3166 (N_3166,N_425,N_2138);
nor U3167 (N_3167,In_154,N_2308);
xnor U3168 (N_3168,N_2649,In_4853);
or U3169 (N_3169,N_2121,N_2124);
nand U3170 (N_3170,N_1609,In_3776);
or U3171 (N_3171,N_2931,N_1201);
nor U3172 (N_3172,N_2959,N_2336);
xnor U3173 (N_3173,N_1939,N_2485);
xor U3174 (N_3174,N_2664,N_2523);
and U3175 (N_3175,N_2493,N_2552);
xor U3176 (N_3176,N_591,N_2669);
nand U3177 (N_3177,N_1311,N_2822);
nor U3178 (N_3178,N_2095,N_2742);
and U3179 (N_3179,N_2906,N_1196);
or U3180 (N_3180,N_2510,N_2622);
nand U3181 (N_3181,N_2979,N_2712);
or U3182 (N_3182,N_2963,N_2460);
nor U3183 (N_3183,N_2791,N_825);
xnor U3184 (N_3184,N_1689,N_38);
xnor U3185 (N_3185,N_536,N_2128);
xnor U3186 (N_3186,N_2219,In_969);
nor U3187 (N_3187,N_1745,N_2113);
nand U3188 (N_3188,N_2015,In_1942);
nor U3189 (N_3189,In_685,In_4263);
or U3190 (N_3190,In_2376,N_2133);
nor U3191 (N_3191,N_79,N_2800);
and U3192 (N_3192,N_1178,N_2386);
nand U3193 (N_3193,N_1240,N_1779);
and U3194 (N_3194,N_2194,N_2776);
nand U3195 (N_3195,N_2631,N_2206);
xnor U3196 (N_3196,N_1229,N_2736);
and U3197 (N_3197,N_2702,N_2354);
and U3198 (N_3198,N_2394,N_2784);
and U3199 (N_3199,N_2424,N_2179);
nor U3200 (N_3200,In_3928,In_4688);
xnor U3201 (N_3201,N_404,N_900);
nand U3202 (N_3202,In_3587,N_2366);
nand U3203 (N_3203,N_2368,N_1738);
xor U3204 (N_3204,N_96,N_109);
or U3205 (N_3205,N_2834,N_2570);
nand U3206 (N_3206,N_2380,In_4674);
or U3207 (N_3207,N_2400,N_969);
xnor U3208 (N_3208,N_2714,N_2975);
xnor U3209 (N_3209,N_1501,N_1095);
and U3210 (N_3210,In_1407,N_2252);
xor U3211 (N_3211,N_2243,N_2969);
nor U3212 (N_3212,N_2650,N_1695);
xnor U3213 (N_3213,In_4506,N_1641);
or U3214 (N_3214,In_2128,N_373);
and U3215 (N_3215,N_2188,N_485);
xor U3216 (N_3216,N_2029,N_2964);
nor U3217 (N_3217,N_1890,In_41);
or U3218 (N_3218,N_1959,N_2358);
or U3219 (N_3219,In_3365,N_2398);
nor U3220 (N_3220,N_2848,N_283);
or U3221 (N_3221,In_4099,In_116);
xor U3222 (N_3222,N_2788,N_2760);
nand U3223 (N_3223,N_2829,N_921);
or U3224 (N_3224,N_2938,N_2363);
nand U3225 (N_3225,N_2849,In_2351);
and U3226 (N_3226,In_3444,N_1440);
nor U3227 (N_3227,N_1578,N_2218);
nor U3228 (N_3228,N_2636,N_2283);
xor U3229 (N_3229,N_2630,N_145);
nor U3230 (N_3230,N_1418,In_372);
or U3231 (N_3231,In_878,In_86);
nor U3232 (N_3232,N_2734,In_4964);
or U3233 (N_3233,N_2266,N_2060);
or U3234 (N_3234,N_2983,In_1472);
and U3235 (N_3235,N_503,N_2036);
nor U3236 (N_3236,N_2259,In_4509);
xnor U3237 (N_3237,N_2372,N_2820);
and U3238 (N_3238,In_2237,In_3443);
xnor U3239 (N_3239,In_4639,N_2645);
xnor U3240 (N_3240,N_1734,N_1322);
xnor U3241 (N_3241,N_2586,N_2681);
and U3242 (N_3242,N_2668,N_2462);
xnor U3243 (N_3243,In_2612,N_2682);
or U3244 (N_3244,In_416,N_2030);
nor U3245 (N_3245,In_2374,In_2251);
xor U3246 (N_3246,N_1200,N_2322);
xor U3247 (N_3247,N_2005,N_1656);
xnor U3248 (N_3248,In_202,N_1310);
nand U3249 (N_3249,In_4648,N_2821);
nand U3250 (N_3250,In_427,N_2228);
nand U3251 (N_3251,In_418,N_2373);
and U3252 (N_3252,In_1109,N_1397);
and U3253 (N_3253,In_3225,N_2458);
nand U3254 (N_3254,In_1326,N_1543);
xor U3255 (N_3255,N_2272,In_3662);
or U3256 (N_3256,In_2378,In_2022);
xor U3257 (N_3257,N_2309,In_3952);
nand U3258 (N_3258,In_2626,N_2126);
nand U3259 (N_3259,N_1363,In_4042);
or U3260 (N_3260,N_2973,N_2799);
xor U3261 (N_3261,In_3534,N_2089);
nor U3262 (N_3262,N_2608,N_1899);
and U3263 (N_3263,N_2321,N_2542);
nor U3264 (N_3264,N_2709,N_2293);
and U3265 (N_3265,N_474,N_2346);
or U3266 (N_3266,N_2442,N_2285);
and U3267 (N_3267,N_2167,N_2757);
and U3268 (N_3268,N_2319,N_398);
or U3269 (N_3269,N_2903,N_2994);
and U3270 (N_3270,N_916,N_2813);
nor U3271 (N_3271,In_4142,N_2098);
and U3272 (N_3272,N_1360,N_891);
or U3273 (N_3273,In_1129,N_2160);
and U3274 (N_3274,In_1085,N_2728);
xnor U3275 (N_3275,N_219,N_2026);
and U3276 (N_3276,In_4662,N_2951);
or U3277 (N_3277,N_2450,N_2290);
xnor U3278 (N_3278,N_2633,In_2055);
nor U3279 (N_3279,In_2819,In_3320);
or U3280 (N_3280,In_1687,N_2299);
nor U3281 (N_3281,N_2474,In_2297);
xor U3282 (N_3282,N_2816,N_2461);
nor U3283 (N_3283,N_970,N_2490);
nand U3284 (N_3284,N_1413,N_2410);
nand U3285 (N_3285,In_2355,N_610);
nor U3286 (N_3286,N_1524,N_2769);
nand U3287 (N_3287,In_4292,N_2530);
or U3288 (N_3288,N_2361,In_807);
xor U3289 (N_3289,In_4376,N_2628);
nand U3290 (N_3290,N_2274,In_4110);
nand U3291 (N_3291,N_1072,In_656);
nand U3292 (N_3292,N_2018,N_2280);
nand U3293 (N_3293,N_846,N_2624);
and U3294 (N_3294,In_3523,N_2384);
or U3295 (N_3295,N_1873,N_2184);
xor U3296 (N_3296,In_3856,N_2893);
and U3297 (N_3297,N_2655,N_2884);
and U3298 (N_3298,N_2502,N_2875);
xnor U3299 (N_3299,N_775,N_2264);
nor U3300 (N_3300,N_1781,N_2014);
xnor U3301 (N_3301,N_2902,N_2642);
and U3302 (N_3302,In_4206,In_4194);
xnor U3303 (N_3303,N_2770,N_2174);
nand U3304 (N_3304,In_4090,N_1112);
or U3305 (N_3305,In_1860,In_2441);
nor U3306 (N_3306,N_2706,N_2877);
xnor U3307 (N_3307,In_4653,N_2189);
nand U3308 (N_3308,N_367,N_552);
xnor U3309 (N_3309,N_2847,In_2066);
nand U3310 (N_3310,N_2207,N_2159);
nor U3311 (N_3311,N_1777,N_2694);
nor U3312 (N_3312,N_1251,N_2318);
nand U3313 (N_3313,N_2221,N_2943);
nor U3314 (N_3314,In_1008,N_1992);
and U3315 (N_3315,N_2888,N_2499);
nand U3316 (N_3316,N_2214,N_2013);
xnor U3317 (N_3317,N_284,N_1492);
nor U3318 (N_3318,In_1330,N_33);
nand U3319 (N_3319,In_4938,N_1011);
xor U3320 (N_3320,In_675,N_2166);
nor U3321 (N_3321,N_2646,In_1346);
nand U3322 (N_3322,N_2635,In_1137);
or U3323 (N_3323,N_2211,N_1277);
nor U3324 (N_3324,N_1244,N_1752);
xor U3325 (N_3325,N_2261,In_74);
and U3326 (N_3326,N_2116,In_2502);
nor U3327 (N_3327,In_2043,In_3377);
or U3328 (N_3328,N_2339,N_2362);
or U3329 (N_3329,N_1700,N_1605);
and U3330 (N_3330,N_1006,N_1854);
nor U3331 (N_3331,N_1138,N_2317);
nand U3332 (N_3332,N_2156,N_2340);
or U3333 (N_3333,N_2487,In_1323);
nand U3334 (N_3334,N_2854,N_2609);
xor U3335 (N_3335,In_2057,N_2350);
nor U3336 (N_3336,In_2998,In_4818);
nor U3337 (N_3337,N_2925,N_2222);
nand U3338 (N_3338,N_2165,N_2953);
or U3339 (N_3339,N_2040,N_2476);
nor U3340 (N_3340,N_2764,N_1118);
and U3341 (N_3341,In_2282,N_2550);
or U3342 (N_3342,N_2226,N_378);
nand U3343 (N_3343,In_1281,N_1567);
nand U3344 (N_3344,N_2454,N_2972);
nor U3345 (N_3345,N_2995,In_2165);
nor U3346 (N_3346,In_4587,N_2417);
or U3347 (N_3347,In_4031,In_2572);
or U3348 (N_3348,N_2700,N_2275);
nand U3349 (N_3349,N_2047,N_2338);
nand U3350 (N_3350,N_2805,In_1091);
and U3351 (N_3351,In_1872,N_1876);
xor U3352 (N_3352,In_3517,In_2027);
or U3353 (N_3353,N_2270,N_1404);
and U3354 (N_3354,N_1380,N_2864);
nand U3355 (N_3355,N_1772,N_2420);
nand U3356 (N_3356,N_2023,N_2775);
nand U3357 (N_3357,N_369,N_1315);
or U3358 (N_3358,N_2672,N_2300);
xnor U3359 (N_3359,N_2464,N_2600);
nor U3360 (N_3360,In_2060,N_2431);
nand U3361 (N_3361,N_2790,N_2780);
nor U3362 (N_3362,N_324,N_2939);
nor U3363 (N_3363,N_1464,N_1099);
and U3364 (N_3364,In_745,N_2948);
xor U3365 (N_3365,In_900,N_2845);
xnor U3366 (N_3366,N_2607,N_2565);
or U3367 (N_3367,N_1655,N_2038);
and U3368 (N_3368,N_2053,N_927);
or U3369 (N_3369,In_2213,N_2731);
or U3370 (N_3370,N_2955,In_3210);
and U3371 (N_3371,N_2383,N_241);
xor U3372 (N_3372,In_4503,In_4309);
or U3373 (N_3373,N_2662,N_1593);
nand U3374 (N_3374,N_2057,N_762);
and U3375 (N_3375,N_2200,N_2626);
nand U3376 (N_3376,N_2679,N_2096);
xor U3377 (N_3377,N_2144,N_2656);
nand U3378 (N_3378,N_791,N_2181);
xor U3379 (N_3379,N_2687,In_3131);
and U3380 (N_3380,N_2078,N_2425);
nor U3381 (N_3381,N_2732,N_322);
nand U3382 (N_3382,N_1417,N_411);
and U3383 (N_3383,N_1484,In_300);
nand U3384 (N_3384,In_2975,N_2120);
nand U3385 (N_3385,N_2724,N_1058);
nor U3386 (N_3386,N_2899,In_1905);
and U3387 (N_3387,N_2750,N_2204);
or U3388 (N_3388,N_2109,N_1539);
nand U3389 (N_3389,N_2898,N_1941);
and U3390 (N_3390,In_2116,N_1614);
and U3391 (N_3391,N_2162,N_53);
nand U3392 (N_3392,N_2999,N_1731);
and U3393 (N_3393,In_2633,N_1904);
nand U3394 (N_3394,N_2716,N_1426);
nand U3395 (N_3395,N_2858,N_2612);
xor U3396 (N_3396,In_1510,N_1465);
nor U3397 (N_3397,N_2560,N_2766);
nor U3398 (N_3398,N_2301,N_1081);
nand U3399 (N_3399,N_2064,N_2564);
nor U3400 (N_3400,N_2756,In_151);
nor U3401 (N_3401,N_2418,N_1780);
and U3402 (N_3402,N_2987,N_2069);
nand U3403 (N_3403,N_2389,N_2406);
nor U3404 (N_3404,N_1059,N_2562);
xor U3405 (N_3405,N_1030,N_1222);
and U3406 (N_3406,N_1323,N_2117);
nor U3407 (N_3407,N_2314,In_1011);
or U3408 (N_3408,N_2508,N_2441);
and U3409 (N_3409,N_2774,N_2494);
or U3410 (N_3410,N_2143,In_4884);
and U3411 (N_3411,In_2223,N_154);
or U3412 (N_3412,In_1202,N_2000);
and U3413 (N_3413,N_2328,N_1455);
nand U3414 (N_3414,In_1431,N_1224);
nand U3415 (N_3415,In_1205,N_2203);
xnor U3416 (N_3416,In_3628,In_3172);
nor U3417 (N_3417,N_2763,In_3936);
and U3418 (N_3418,N_2512,In_494);
or U3419 (N_3419,N_2183,In_453);
nand U3420 (N_3420,In_423,In_2420);
and U3421 (N_3421,In_2036,In_3994);
or U3422 (N_3422,N_2492,N_1674);
and U3423 (N_3423,N_1574,N_2151);
nand U3424 (N_3424,N_403,N_142);
or U3425 (N_3425,N_2349,N_258);
and U3426 (N_3426,N_1023,In_1175);
nand U3427 (N_3427,N_2323,N_2254);
or U3428 (N_3428,N_537,In_4946);
nor U3429 (N_3429,In_3113,In_2371);
and U3430 (N_3430,N_1481,N_1436);
or U3431 (N_3431,In_4971,In_1653);
xnor U3432 (N_3432,In_2443,In_2471);
or U3433 (N_3433,N_2068,N_2632);
nor U3434 (N_3434,N_1742,In_2751);
xor U3435 (N_3435,In_4337,In_4330);
nor U3436 (N_3436,N_129,N_2479);
nor U3437 (N_3437,N_2032,In_3622);
xor U3438 (N_3438,In_84,N_1447);
and U3439 (N_3439,In_3846,N_2347);
or U3440 (N_3440,N_2653,In_3142);
and U3441 (N_3441,N_2489,N_2074);
xnor U3442 (N_3442,N_1016,In_654);
xor U3443 (N_3443,N_1056,N_2045);
and U3444 (N_3444,N_2396,In_3966);
xnor U3445 (N_3445,N_1407,In_318);
and U3446 (N_3446,N_1606,N_2837);
and U3447 (N_3447,N_604,N_2707);
or U3448 (N_3448,N_2112,In_4433);
nor U3449 (N_3449,N_2178,N_2895);
and U3450 (N_3450,N_1767,In_375);
nand U3451 (N_3451,In_239,N_2841);
xnor U3452 (N_3452,N_2990,N_2744);
xnor U3453 (N_3453,N_2894,In_4988);
or U3454 (N_3454,In_934,In_2838);
or U3455 (N_3455,N_2659,N_171);
or U3456 (N_3456,In_2361,N_2629);
and U3457 (N_3457,In_2689,N_2661);
or U3458 (N_3458,N_2310,In_1453);
or U3459 (N_3459,N_2551,In_3993);
nor U3460 (N_3460,N_2145,N_2572);
nor U3461 (N_3461,N_907,N_2455);
nor U3462 (N_3462,In_861,N_2883);
xor U3463 (N_3463,In_1999,N_516);
or U3464 (N_3464,N_2940,N_2465);
and U3465 (N_3465,N_1387,N_2307);
nor U3466 (N_3466,N_2288,N_2620);
xnor U3467 (N_3467,N_2027,In_3714);
nor U3468 (N_3468,N_2088,N_2348);
nand U3469 (N_3469,N_1552,N_2762);
and U3470 (N_3470,N_2536,N_773);
xnor U3471 (N_3471,N_2130,N_2613);
or U3472 (N_3472,N_2860,N_813);
nand U3473 (N_3473,N_804,In_2195);
nand U3474 (N_3474,In_195,N_2247);
nand U3475 (N_3475,N_2598,N_2367);
or U3476 (N_3476,In_509,N_1050);
nand U3477 (N_3477,N_65,N_2426);
nor U3478 (N_3478,N_2127,In_329);
nor U3479 (N_3479,In_2867,N_2245);
xnor U3480 (N_3480,N_2101,N_1419);
or U3481 (N_3481,N_2887,N_1045);
nand U3482 (N_3482,In_125,N_1029);
nor U3483 (N_3483,N_2066,In_1523);
nor U3484 (N_3484,In_3368,N_2678);
or U3485 (N_3485,N_2924,In_2832);
xnor U3486 (N_3486,In_1555,N_653);
nor U3487 (N_3487,In_2590,N_2830);
xnor U3488 (N_3488,N_2765,N_2812);
and U3489 (N_3489,N_2404,N_2927);
xor U3490 (N_3490,N_2720,In_2266);
and U3491 (N_3491,N_2808,N_2087);
nor U3492 (N_3492,N_2423,N_2717);
or U3493 (N_3493,In_3226,N_2647);
nand U3494 (N_3494,In_2531,N_2281);
xor U3495 (N_3495,In_1420,N_2752);
nand U3496 (N_3496,N_1337,N_2984);
nand U3497 (N_3497,N_2554,N_1804);
xnor U3498 (N_3498,N_2447,N_2480);
or U3499 (N_3499,N_2185,N_2054);
nand U3500 (N_3500,N_1797,N_2873);
nor U3501 (N_3501,In_2290,N_2594);
nand U3502 (N_3502,N_1798,N_1008);
and U3503 (N_3503,N_783,N_2390);
and U3504 (N_3504,N_2909,In_1025);
and U3505 (N_3505,In_63,N_1579);
nor U3506 (N_3506,N_2777,N_2149);
or U3507 (N_3507,N_2846,N_1513);
nor U3508 (N_3508,N_1292,In_1904);
nor U3509 (N_3509,N_2577,N_603);
and U3510 (N_3510,N_67,N_2735);
or U3511 (N_3511,N_2388,In_293);
and U3512 (N_3512,N_2779,N_2749);
and U3513 (N_3513,N_748,N_2311);
nor U3514 (N_3514,N_2320,N_2269);
and U3515 (N_3515,N_2409,N_2839);
nand U3516 (N_3516,In_2665,N_554);
or U3517 (N_3517,N_1795,N_1300);
and U3518 (N_3518,N_2164,N_1151);
and U3519 (N_3519,N_2227,In_3725);
or U3520 (N_3520,In_4083,N_2155);
nand U3521 (N_3521,In_3462,In_3214);
and U3522 (N_3522,N_2680,In_11);
xor U3523 (N_3523,N_1601,N_747);
and U3524 (N_3524,In_907,N_317);
or U3525 (N_3525,N_2132,N_2699);
or U3526 (N_3526,N_2058,N_1783);
and U3527 (N_3527,N_2991,N_2676);
nor U3528 (N_3528,N_2965,N_2996);
xor U3529 (N_3529,N_2559,In_704);
nor U3530 (N_3530,N_2119,N_2654);
and U3531 (N_3531,N_941,N_1089);
xor U3532 (N_3532,In_3697,N_2801);
nand U3533 (N_3533,N_2070,N_2538);
or U3534 (N_3534,In_3357,N_2582);
nand U3535 (N_3535,N_2342,In_4800);
nand U3536 (N_3536,In_2445,N_1749);
nand U3537 (N_3537,N_570,In_3876);
nand U3538 (N_3538,N_2168,N_593);
nand U3539 (N_3539,N_2456,N_2606);
xor U3540 (N_3540,In_912,In_1490);
nand U3541 (N_3541,In_461,In_2209);
nor U3542 (N_3542,N_2978,In_4580);
or U3543 (N_3543,N_2782,N_2100);
nor U3544 (N_3544,N_2627,N_2104);
and U3545 (N_3545,N_1021,N_2276);
and U3546 (N_3546,N_2405,N_2067);
xnor U3547 (N_3547,N_1955,In_2515);
xor U3548 (N_3548,N_2584,In_2379);
or U3549 (N_3549,N_524,N_1267);
nand U3550 (N_3550,N_2605,N_2558);
or U3551 (N_3551,N_2541,In_3166);
nor U3552 (N_3552,In_1,N_2110);
xor U3553 (N_3553,In_4277,N_2284);
xor U3554 (N_3554,N_2048,In_1720);
nor U3555 (N_3555,N_2786,N_1627);
xnor U3556 (N_3556,In_4406,N_1180);
xnor U3557 (N_3557,In_2825,In_2939);
or U3558 (N_3558,In_3025,N_1489);
or U3559 (N_3559,In_3284,N_2242);
nor U3560 (N_3560,N_2031,N_1367);
xor U3561 (N_3561,N_2803,N_2549);
and U3562 (N_3562,In_4944,In_3736);
and U3563 (N_3563,In_3380,N_679);
nand U3564 (N_3564,N_2910,N_2806);
and U3565 (N_3565,N_2408,N_2282);
xor U3566 (N_3566,In_1977,N_1259);
nor U3567 (N_3567,N_2807,N_2675);
nand U3568 (N_3568,N_2998,N_1243);
nand U3569 (N_3569,N_2674,N_1728);
nor U3570 (N_3570,In_3971,N_2602);
and U3571 (N_3571,N_2375,N_2954);
xor U3572 (N_3572,N_2980,N_266);
or U3573 (N_3573,In_2092,N_779);
nand U3574 (N_3574,N_2341,N_2976);
and U3575 (N_3575,N_2125,N_2889);
xnor U3576 (N_3576,In_3209,N_2547);
xnor U3577 (N_3577,N_2974,N_1416);
nor U3578 (N_3578,N_2880,N_2759);
xnor U3579 (N_3579,In_3878,N_2020);
and U3580 (N_3580,N_2271,N_2357);
nor U3581 (N_3581,N_2019,N_1220);
xnor U3582 (N_3582,In_2309,N_2746);
or U3583 (N_3583,N_2637,N_1424);
or U3584 (N_3584,N_2484,In_1570);
xnor U3585 (N_3585,N_2593,N_2090);
and U3586 (N_3586,N_1116,N_2215);
nand U3587 (N_3587,In_2330,N_1650);
nand U3588 (N_3588,In_1974,N_2967);
nor U3589 (N_3589,N_1071,N_2016);
or U3590 (N_3590,N_2152,N_2419);
and U3591 (N_3591,N_2131,In_1511);
nand U3592 (N_3592,N_2483,N_2768);
or U3593 (N_3593,N_158,N_2727);
nor U3594 (N_3594,N_984,N_1519);
nand U3595 (N_3595,N_1245,N_71);
xor U3596 (N_3596,N_1149,In_1698);
nor U3597 (N_3597,N_2871,N_2002);
or U3598 (N_3598,In_342,N_2260);
and U3599 (N_3599,N_2028,In_1703);
xor U3600 (N_3600,N_1351,N_2828);
xnor U3601 (N_3601,N_636,N_2108);
nor U3602 (N_3602,N_277,N_1487);
and U3603 (N_3603,N_1748,In_2774);
nand U3604 (N_3604,N_2238,N_2106);
or U3605 (N_3605,N_2666,In_4599);
nand U3606 (N_3606,In_562,In_4273);
nor U3607 (N_3607,In_3677,In_2097);
nor U3608 (N_3608,N_2092,In_3604);
nor U3609 (N_3609,N_1530,N_2912);
nor U3610 (N_3610,In_3502,In_3550);
nand U3611 (N_3611,In_1605,N_2084);
nor U3612 (N_3612,N_2050,N_2402);
nor U3613 (N_3613,N_2958,N_2640);
and U3614 (N_3614,N_1334,N_2107);
nand U3615 (N_3615,In_4992,In_2972);
nand U3616 (N_3616,N_2919,N_2950);
xnor U3617 (N_3617,In_2123,N_2478);
nand U3618 (N_3618,In_4314,In_2406);
nand U3619 (N_3619,N_2591,In_2611);
and U3620 (N_3620,In_4054,N_2470);
or U3621 (N_3621,N_1669,N_2851);
and U3622 (N_3622,N_2176,N_2268);
nor U3623 (N_3623,In_3692,N_2374);
and U3624 (N_3624,N_2004,N_2326);
xnor U3625 (N_3625,N_2677,N_2052);
nor U3626 (N_3626,In_4667,N_1010);
nand U3627 (N_3627,N_2192,N_1617);
nor U3628 (N_3628,In_1489,N_2150);
nand U3629 (N_3629,N_2618,N_2287);
and U3630 (N_3630,In_4076,In_645);
nor U3631 (N_3631,N_2071,N_2738);
nor U3632 (N_3632,In_2834,N_1191);
and U3633 (N_3633,N_1102,N_1002);
and U3634 (N_3634,N_2575,In_3016);
or U3635 (N_3635,N_2115,N_2869);
nor U3636 (N_3636,N_2267,N_2205);
or U3637 (N_3637,N_2517,N_2603);
and U3638 (N_3638,N_2244,N_2697);
and U3639 (N_3639,In_644,N_2667);
or U3640 (N_3640,N_2797,N_1516);
xnor U3641 (N_3641,N_1402,N_1505);
and U3642 (N_3642,N_2414,In_4511);
nor U3643 (N_3643,N_2833,In_4078);
xnor U3644 (N_3644,N_1368,In_3175);
and U3645 (N_3645,N_2239,N_1472);
nand U3646 (N_3646,In_852,N_2583);
nand U3647 (N_3647,N_2773,N_2170);
or U3648 (N_3648,N_2504,N_2838);
nor U3649 (N_3649,N_1974,N_2692);
or U3650 (N_3650,N_2885,In_3435);
and U3651 (N_3651,N_2193,N_1740);
nand U3652 (N_3652,N_2468,In_190);
or U3653 (N_3653,In_4478,N_2278);
or U3654 (N_3654,In_4991,In_3866);
nand U3655 (N_3655,N_1231,In_4190);
xnor U3656 (N_3656,N_1691,In_2748);
nor U3657 (N_3657,In_305,N_2359);
nand U3658 (N_3658,N_838,N_2224);
nor U3659 (N_3659,N_2561,In_1964);
or U3660 (N_3660,N_1445,N_2171);
nor U3661 (N_3661,N_2003,N_2989);
or U3662 (N_3662,N_2435,N_2719);
xor U3663 (N_3663,N_2616,In_303);
xnor U3664 (N_3664,N_1153,N_1250);
nor U3665 (N_3665,In_4595,N_2535);
and U3666 (N_3666,N_1809,N_785);
xor U3667 (N_3667,In_1825,N_2315);
nand U3668 (N_3668,N_2376,N_2072);
nand U3669 (N_3669,N_1755,N_2496);
nand U3670 (N_3670,N_1789,N_2588);
and U3671 (N_3671,N_2993,N_1872);
nor U3672 (N_3672,N_2914,In_754);
and U3673 (N_3673,N_278,N_1927);
nor U3674 (N_3674,In_4407,N_2438);
xor U3675 (N_3675,N_2352,In_2878);
and U3676 (N_3676,In_4705,N_1264);
xnor U3677 (N_3677,N_1792,N_2046);
and U3678 (N_3678,N_1076,N_868);
nand U3679 (N_3679,N_1988,In_2868);
nor U3680 (N_3680,N_2882,N_2495);
nand U3681 (N_3681,N_2708,N_2062);
and U3682 (N_3682,In_3317,N_2579);
xor U3683 (N_3683,N_2639,N_1176);
and U3684 (N_3684,N_2874,N_1531);
xor U3685 (N_3685,N_2625,N_383);
nor U3686 (N_3686,In_3422,N_1276);
nand U3687 (N_3687,N_2545,N_2500);
xnor U3688 (N_3688,In_25,N_63);
nand U3689 (N_3689,N_1915,N_2457);
and U3690 (N_3690,In_363,N_2809);
and U3691 (N_3691,In_332,N_2962);
and U3692 (N_3692,N_2522,In_501);
nand U3693 (N_3693,In_2646,In_1848);
nand U3694 (N_3694,N_2223,N_1681);
xor U3695 (N_3695,N_18,N_2332);
nand U3696 (N_3696,N_2663,N_2982);
and U3697 (N_3697,N_1785,N_2241);
nor U3698 (N_3698,N_2093,N_2146);
nand U3699 (N_3699,N_1773,N_2099);
nand U3700 (N_3700,In_4819,N_1261);
nand U3701 (N_3701,N_2988,N_2852);
and U3702 (N_3702,N_2657,In_4710);
or U3703 (N_3703,In_1734,N_1254);
nor U3704 (N_3704,In_3031,N_231);
nand U3705 (N_3705,In_829,N_2355);
and U3706 (N_3706,N_2514,In_1187);
xnor U3707 (N_3707,N_351,N_2365);
and U3708 (N_3708,N_2548,N_2216);
nand U3709 (N_3709,N_2900,In_1599);
and U3710 (N_3710,N_1188,N_2289);
xnor U3711 (N_3711,In_1932,N_2377);
xnor U3712 (N_3712,In_4649,N_2638);
or U3713 (N_3713,N_2688,N_1468);
nand U3714 (N_3714,In_4052,N_818);
nand U3715 (N_3715,In_3240,In_874);
nand U3716 (N_3716,In_3871,N_2443);
nand U3717 (N_3717,N_2233,N_2743);
nand U3718 (N_3718,N_1000,N_726);
or U3719 (N_3719,N_2397,In_1951);
xnor U3720 (N_3720,N_2917,N_1018);
xor U3721 (N_3721,In_4935,In_3143);
nor U3722 (N_3722,In_1314,N_2399);
nor U3723 (N_3723,N_2379,N_1184);
and U3724 (N_3724,N_2076,N_2169);
xnor U3725 (N_3725,In_3568,N_1615);
nor U3726 (N_3726,N_2519,N_2739);
and U3727 (N_3727,N_1179,N_901);
xor U3728 (N_3728,In_3085,N_2585);
and U3729 (N_3729,N_2952,In_4047);
or U3730 (N_3730,N_2685,N_2304);
and U3731 (N_3731,N_1106,N_2798);
nor U3732 (N_3732,In_559,N_2641);
or U3733 (N_3733,N_2673,In_3026);
nand U3734 (N_3734,N_234,N_2196);
nor U3735 (N_3735,N_2393,N_2696);
or U3736 (N_3736,In_4900,N_2291);
and U3737 (N_3737,N_2540,N_2158);
nand U3738 (N_3738,N_1642,N_2693);
and U3739 (N_3739,N_31,N_2022);
xor U3740 (N_3740,N_2059,N_2111);
or U3741 (N_3741,In_4795,In_4553);
or U3742 (N_3742,N_1325,In_2141);
and U3743 (N_3743,N_433,In_3741);
nand U3744 (N_3744,In_2906,N_2246);
nor U3745 (N_3745,N_2870,N_2981);
nor U3746 (N_3746,N_2546,N_2370);
and U3747 (N_3747,N_2080,N_1282);
or U3748 (N_3748,N_2081,In_3709);
nand U3749 (N_3749,N_693,In_585);
xor U3750 (N_3750,N_2892,N_1048);
xor U3751 (N_3751,N_2255,In_4871);
nand U3752 (N_3752,N_2007,N_2597);
xor U3753 (N_3753,N_2011,N_1663);
nor U3754 (N_3754,In_4294,In_2272);
nand U3755 (N_3755,N_712,N_2012);
and U3756 (N_3756,N_2477,N_2566);
nand U3757 (N_3757,N_1533,N_497);
nor U3758 (N_3758,In_1997,N_860);
or U3759 (N_3759,In_1893,N_2475);
and U3760 (N_3760,N_2446,N_2918);
nor U3761 (N_3761,In_3156,In_433);
xor U3762 (N_3762,N_2415,N_2353);
nor U3763 (N_3763,N_2992,N_2683);
or U3764 (N_3764,N_814,N_2826);
or U3765 (N_3765,N_2872,In_2623);
or U3766 (N_3766,N_1573,In_4773);
nor U3767 (N_3767,N_2230,N_1512);
and U3768 (N_3768,N_2086,N_1864);
nand U3769 (N_3769,N_2056,N_2711);
or U3770 (N_3770,N_1097,In_4281);
or U3771 (N_3771,N_2905,N_2345);
xnor U3772 (N_3772,In_2286,N_2213);
xnor U3773 (N_3773,In_774,N_2921);
nand U3774 (N_3774,N_2590,In_3617);
xnor U3775 (N_3775,N_2235,N_2946);
nand U3776 (N_3776,N_2175,N_543);
and U3777 (N_3777,N_2758,N_2568);
xnor U3778 (N_3778,In_1968,N_1348);
nand U3779 (N_3779,N_1362,N_2190);
xor U3780 (N_3780,N_2298,In_2691);
nand U3781 (N_3781,N_2371,In_801);
and U3782 (N_3782,N_2843,In_611);
nand U3783 (N_3783,N_2741,In_613);
and U3784 (N_3784,In_1622,N_2137);
xnor U3785 (N_3785,N_2364,N_1953);
nand U3786 (N_3786,In_3562,N_2258);
nand U3787 (N_3787,N_1124,N_811);
or U3788 (N_3788,In_1224,N_2378);
or U3789 (N_3789,N_2610,N_2922);
xnor U3790 (N_3790,N_47,N_2896);
and U3791 (N_3791,N_2589,N_2737);
nand U3792 (N_3792,N_1433,In_1564);
nand U3793 (N_3793,In_4915,N_2966);
xnor U3794 (N_3794,In_3939,In_1198);
nand U3795 (N_3795,N_812,N_23);
nand U3796 (N_3796,In_3034,N_2256);
and U3797 (N_3797,N_2935,N_1237);
or U3798 (N_3798,In_129,In_394);
nand U3799 (N_3799,In_598,N_1170);
and U3800 (N_3800,In_794,N_2930);
and U3801 (N_3801,N_2369,N_674);
or U3802 (N_3802,In_4525,In_1625);
and U3803 (N_3803,N_2853,N_2482);
and U3804 (N_3804,N_2932,N_2436);
xnor U3805 (N_3805,N_2970,In_401);
nand U3806 (N_3806,N_2556,N_2897);
or U3807 (N_3807,N_1631,In_121);
xnor U3808 (N_3808,N_1800,N_2771);
nor U3809 (N_3809,N_2986,N_1704);
or U3810 (N_3810,In_1336,N_2430);
nand U3811 (N_3811,N_2407,N_2198);
nor U3812 (N_3812,N_1608,In_1839);
or U3813 (N_3813,N_2163,N_2008);
or U3814 (N_3814,N_2539,N_205);
xor U3815 (N_3815,N_2623,N_1769);
or U3816 (N_3816,In_798,N_2815);
and U3817 (N_3817,N_2867,N_2105);
nand U3818 (N_3818,N_2433,N_2515);
nand U3819 (N_3819,N_98,N_1449);
or U3820 (N_3820,N_2715,In_2377);
or U3821 (N_3821,N_738,N_2153);
nand U3822 (N_3822,N_1478,N_2968);
and U3823 (N_3823,N_1805,N_1961);
and U3824 (N_3824,N_2644,N_2199);
nor U3825 (N_3825,N_2063,N_1897);
xnor U3826 (N_3826,N_2265,N_2428);
and U3827 (N_3827,N_1163,In_3577);
nand U3828 (N_3828,N_701,N_2427);
nor U3829 (N_3829,N_1024,N_2850);
or U3830 (N_3830,In_408,N_1957);
or U3831 (N_3831,In_2761,In_3429);
or U3832 (N_3832,In_2608,N_2416);
or U3833 (N_3833,In_4426,N_631);
nor U3834 (N_3834,N_2356,In_1919);
nor U3835 (N_3835,N_2557,N_2229);
nor U3836 (N_3836,N_2232,N_1952);
and U3837 (N_3837,N_2049,In_2821);
and U3838 (N_3838,N_2703,N_2818);
nand U3839 (N_3839,N_2509,In_3079);
xnor U3840 (N_3840,N_2333,N_2471);
and U3841 (N_3841,In_3201,N_2604);
xor U3842 (N_3842,N_2294,N_2587);
nand U3843 (N_3843,N_2862,N_1756);
nand U3844 (N_3844,In_2883,N_2936);
nor U3845 (N_3845,N_1411,N_1459);
or U3846 (N_3846,In_1347,In_555);
and U3847 (N_3847,N_1842,In_1783);
nand U3848 (N_3848,N_2296,In_727);
nor U3849 (N_3849,N_2439,In_2830);
nand U3850 (N_3850,N_2740,N_2316);
and U3851 (N_3851,N_2501,N_1852);
nor U3852 (N_3852,N_2596,N_2891);
nor U3853 (N_3853,N_2044,N_2592);
and U3854 (N_3854,In_1072,In_4958);
nor U3855 (N_3855,N_2933,N_1266);
or U3856 (N_3856,N_2581,N_2473);
or U3857 (N_3857,In_2352,N_1166);
and U3858 (N_3858,In_961,N_2886);
xor U3859 (N_3859,N_1547,N_1129);
and U3860 (N_3860,N_2721,N_2202);
xor U3861 (N_3861,N_2452,N_2469);
or U3862 (N_3862,N_368,In_3729);
nor U3863 (N_3863,N_2253,N_2360);
xnor U3864 (N_3864,N_2382,N_1083);
and U3865 (N_3865,In_4035,In_1677);
nor U3866 (N_3866,N_2182,In_4141);
or U3867 (N_3867,N_99,N_2208);
or U3868 (N_3868,N_2306,N_2009);
nor U3869 (N_3869,N_2135,N_1929);
and U3870 (N_3870,In_1101,In_4086);
nor U3871 (N_3871,N_1638,N_1963);
xor U3872 (N_3872,N_2652,N_2525);
nand U3873 (N_3873,N_2614,N_2335);
and U3874 (N_3874,N_2945,N_2527);
nor U3875 (N_3875,N_2091,N_2403);
or U3876 (N_3876,N_2263,In_4198);
nor U3877 (N_3877,N_1256,In_2958);
nor U3878 (N_3878,N_1762,N_407);
and U3879 (N_3879,N_2097,N_2449);
and U3880 (N_3880,N_2792,N_1984);
xnor U3881 (N_3881,In_2775,In_1277);
and U3882 (N_3882,N_2840,N_2035);
or U3883 (N_3883,N_1062,N_2249);
nor U3884 (N_3884,N_77,N_1537);
or U3885 (N_3885,In_38,In_1221);
xor U3886 (N_3886,N_1758,N_1841);
or U3887 (N_3887,N_2911,N_2082);
nand U3888 (N_3888,N_2726,N_2857);
and U3889 (N_3889,N_1892,N_1729);
nand U3890 (N_3890,N_2844,N_1475);
xnor U3891 (N_3891,N_1679,N_1425);
and U3892 (N_3892,N_2488,N_327);
nand U3893 (N_3893,N_2619,In_1493);
nand U3894 (N_3894,N_2651,N_1252);
nor U3895 (N_3895,In_3140,In_2545);
and U3896 (N_3896,In_524,N_1643);
and U3897 (N_3897,In_1922,N_1339);
nand U3898 (N_3898,N_1139,N_2544);
xor U3899 (N_3899,In_1975,N_1498);
and U3900 (N_3900,N_1562,N_2017);
nand U3901 (N_3901,N_2459,N_2997);
xor U3902 (N_3902,N_1070,N_2385);
xor U3903 (N_3903,N_609,N_2481);
and U3904 (N_3904,In_532,In_3559);
nand U3905 (N_3905,In_4565,N_2907);
nand U3906 (N_3906,N_2926,N_1467);
and U3907 (N_3907,N_2021,N_2621);
or U3908 (N_3908,N_2617,N_2861);
or U3909 (N_3909,N_1836,N_2043);
nand U3910 (N_3910,N_2794,N_2804);
xor U3911 (N_3911,In_756,In_307);
nand U3912 (N_3912,N_2034,N_2690);
nand U3913 (N_3913,N_2297,N_396);
nand U3914 (N_3914,In_1723,N_2863);
xnor U3915 (N_3915,N_2755,In_3395);
nor U3916 (N_3916,N_2754,N_1771);
nor U3917 (N_3917,N_1604,N_1958);
xnor U3918 (N_3918,N_1860,In_3737);
and U3919 (N_3919,In_91,N_833);
nor U3920 (N_3920,N_766,N_1702);
nand U3921 (N_3921,N_2658,In_328);
and U3922 (N_3922,In_3904,N_2083);
xnor U3923 (N_3923,N_1033,N_2324);
and U3924 (N_3924,In_3130,N_1803);
xnor U3925 (N_3925,N_1442,N_2421);
nand U3926 (N_3926,N_2337,In_3366);
and U3927 (N_3927,N_2722,In_1623);
and U3928 (N_3928,N_2505,N_1273);
and U3929 (N_3929,N_2033,N_2578);
and U3930 (N_3930,In_4827,N_2778);
nor U3931 (N_3931,In_4514,N_1466);
or U3932 (N_3932,N_2186,N_1648);
or U3933 (N_3933,In_1352,N_2212);
nor U3934 (N_3934,In_629,N_2985);
or U3935 (N_3935,N_829,N_2521);
nor U3936 (N_3936,N_742,In_2674);
and U3937 (N_3937,N_2010,N_2611);
xor U3938 (N_3938,N_2814,N_2942);
xnor U3939 (N_3939,N_2529,N_1931);
xnor U3940 (N_3940,N_1025,N_2001);
xor U3941 (N_3941,In_3811,N_242);
nand U3942 (N_3942,N_2210,In_701);
nor U3943 (N_3943,N_1825,N_2313);
nor U3944 (N_3944,N_2947,In_4670);
nor U3945 (N_3945,In_4537,N_1680);
nand U3946 (N_3946,N_2569,N_2513);
and U3947 (N_3947,N_1093,N_2859);
and U3948 (N_3948,N_2856,In_4067);
nand U3949 (N_3949,N_1306,N_93);
or U3950 (N_3950,In_396,In_4729);
nand U3951 (N_3951,N_1290,N_409);
xnor U3952 (N_3952,N_1287,N_1278);
nor U3953 (N_3953,In_3334,N_1495);
nor U3954 (N_3954,N_1802,N_656);
or U3955 (N_3955,N_2412,N_2819);
or U3956 (N_3956,N_2197,N_2855);
xnor U3957 (N_3957,N_2429,In_4269);
nor U3958 (N_3958,N_2971,N_2472);
nand U3959 (N_3959,N_1386,N_493);
or U3960 (N_3960,In_2956,N_2177);
or U3961 (N_3961,N_2705,In_1113);
nand U3962 (N_3962,N_2065,N_2691);
and U3963 (N_3963,N_2767,In_3933);
nand U3964 (N_3964,N_2432,In_4214);
and U3965 (N_3965,In_535,In_1394);
or U3966 (N_3966,N_2139,N_2524);
or U3967 (N_3967,N_73,N_2344);
nor U3968 (N_3968,N_1090,N_2704);
or U3969 (N_3969,N_1204,N_2136);
or U3970 (N_3970,N_2391,N_1985);
nor U3971 (N_3971,N_2901,N_19);
or U3972 (N_3972,In_4018,N_2195);
xnor U3973 (N_3973,N_1667,N_202);
nor U3974 (N_3974,In_81,N_1009);
or U3975 (N_3975,N_2785,N_2960);
xnor U3976 (N_3976,N_2118,N_2747);
nor U3977 (N_3977,N_2733,In_1793);
or U3978 (N_3978,N_2789,N_797);
or U3979 (N_3979,N_1001,N_2730);
nor U3980 (N_3980,N_2161,N_621);
or U3981 (N_3981,N_2463,N_2147);
or U3982 (N_3982,N_1063,N_2908);
nand U3983 (N_3983,N_2325,N_763);
or U3984 (N_3984,N_2881,N_2772);
nor U3985 (N_3985,In_2108,N_466);
and U3986 (N_3986,N_577,N_2122);
nor U3987 (N_3987,In_980,N_1932);
and U3988 (N_3988,N_2037,N_645);
nor U3989 (N_3989,N_2257,N_2331);
nand U3990 (N_3990,N_2601,In_4300);
nor U3991 (N_3991,In_1439,N_350);
or U3992 (N_3992,N_1168,N_2783);
or U3993 (N_3993,In_2628,N_2904);
or U3994 (N_3994,In_3690,N_1575);
and U3995 (N_3995,N_2528,N_2392);
nand U3996 (N_3996,N_2466,N_271);
and U3997 (N_3997,N_2868,N_2503);
nand U3998 (N_3998,N_1382,In_37);
and U3999 (N_3999,N_1084,N_1775);
nand U4000 (N_4000,N_3777,N_3395);
xor U4001 (N_4001,N_3961,N_3585);
nand U4002 (N_4002,N_3093,N_3931);
xor U4003 (N_4003,N_3211,N_3023);
xor U4004 (N_4004,N_3915,N_3392);
nor U4005 (N_4005,N_3889,N_3874);
xor U4006 (N_4006,N_3759,N_3029);
nand U4007 (N_4007,N_3198,N_3255);
xor U4008 (N_4008,N_3057,N_3106);
nand U4009 (N_4009,N_3166,N_3210);
and U4010 (N_4010,N_3489,N_3682);
and U4011 (N_4011,N_3216,N_3923);
xnor U4012 (N_4012,N_3340,N_3007);
and U4013 (N_4013,N_3970,N_3206);
xor U4014 (N_4014,N_3573,N_3997);
or U4015 (N_4015,N_3227,N_3209);
and U4016 (N_4016,N_3688,N_3911);
nand U4017 (N_4017,N_3313,N_3734);
nand U4018 (N_4018,N_3384,N_3017);
nand U4019 (N_4019,N_3813,N_3707);
nor U4020 (N_4020,N_3197,N_3827);
xnor U4021 (N_4021,N_3596,N_3870);
xnor U4022 (N_4022,N_3620,N_3611);
nor U4023 (N_4023,N_3043,N_3304);
xnor U4024 (N_4024,N_3971,N_3276);
xnor U4025 (N_4025,N_3804,N_3951);
nand U4026 (N_4026,N_3268,N_3549);
nor U4027 (N_4027,N_3231,N_3075);
and U4028 (N_4028,N_3912,N_3645);
xor U4029 (N_4029,N_3321,N_3507);
nor U4030 (N_4030,N_3287,N_3969);
nand U4031 (N_4031,N_3862,N_3687);
nor U4032 (N_4032,N_3570,N_3629);
nand U4033 (N_4033,N_3792,N_3134);
nor U4034 (N_4034,N_3218,N_3882);
nor U4035 (N_4035,N_3035,N_3715);
and U4036 (N_4036,N_3562,N_3581);
nand U4037 (N_4037,N_3431,N_3642);
and U4038 (N_4038,N_3014,N_3101);
and U4039 (N_4039,N_3930,N_3040);
nand U4040 (N_4040,N_3621,N_3797);
and U4041 (N_4041,N_3213,N_3836);
and U4042 (N_4042,N_3244,N_3354);
nor U4043 (N_4043,N_3180,N_3714);
xnor U4044 (N_4044,N_3730,N_3439);
or U4045 (N_4045,N_3731,N_3718);
nand U4046 (N_4046,N_3584,N_3194);
xnor U4047 (N_4047,N_3772,N_3551);
xnor U4048 (N_4048,N_3579,N_3236);
or U4049 (N_4049,N_3095,N_3401);
nor U4050 (N_4050,N_3146,N_3670);
nor U4051 (N_4051,N_3619,N_3233);
xor U4052 (N_4052,N_3954,N_3447);
xnor U4053 (N_4053,N_3950,N_3665);
or U4054 (N_4054,N_3494,N_3186);
nor U4055 (N_4055,N_3434,N_3164);
and U4056 (N_4056,N_3791,N_3527);
and U4057 (N_4057,N_3632,N_3280);
nor U4058 (N_4058,N_3099,N_3187);
and U4059 (N_4059,N_3863,N_3992);
or U4060 (N_4060,N_3639,N_3808);
and U4061 (N_4061,N_3638,N_3351);
and U4062 (N_4062,N_3208,N_3427);
or U4063 (N_4063,N_3408,N_3429);
xor U4064 (N_4064,N_3964,N_3633);
or U4065 (N_4065,N_3842,N_3116);
nand U4066 (N_4066,N_3534,N_3524);
nor U4067 (N_4067,N_3936,N_3695);
and U4068 (N_4068,N_3024,N_3848);
nand U4069 (N_4069,N_3540,N_3531);
and U4070 (N_4070,N_3283,N_3366);
and U4071 (N_4071,N_3382,N_3523);
and U4072 (N_4072,N_3428,N_3205);
or U4073 (N_4073,N_3067,N_3819);
or U4074 (N_4074,N_3991,N_3312);
nand U4075 (N_4075,N_3650,N_3722);
or U4076 (N_4076,N_3050,N_3379);
nand U4077 (N_4077,N_3945,N_3663);
and U4078 (N_4078,N_3617,N_3886);
and U4079 (N_4079,N_3595,N_3114);
or U4080 (N_4080,N_3156,N_3577);
xnor U4081 (N_4081,N_3770,N_3193);
xor U4082 (N_4082,N_3583,N_3168);
or U4083 (N_4083,N_3301,N_3248);
nor U4084 (N_4084,N_3451,N_3824);
and U4085 (N_4085,N_3752,N_3421);
nor U4086 (N_4086,N_3165,N_3151);
or U4087 (N_4087,N_3604,N_3601);
nand U4088 (N_4088,N_3440,N_3615);
nor U4089 (N_4089,N_3348,N_3191);
or U4090 (N_4090,N_3190,N_3933);
and U4091 (N_4091,N_3826,N_3341);
nand U4092 (N_4092,N_3884,N_3511);
or U4093 (N_4093,N_3022,N_3793);
xor U4094 (N_4094,N_3393,N_3122);
xnor U4095 (N_4095,N_3185,N_3655);
xnor U4096 (N_4096,N_3012,N_3653);
nand U4097 (N_4097,N_3605,N_3018);
or U4098 (N_4098,N_3569,N_3820);
or U4099 (N_4099,N_3060,N_3973);
nand U4100 (N_4100,N_3952,N_3356);
or U4101 (N_4101,N_3253,N_3436);
nand U4102 (N_4102,N_3654,N_3861);
nor U4103 (N_4103,N_3815,N_3533);
and U4104 (N_4104,N_3674,N_3140);
xor U4105 (N_4105,N_3956,N_3976);
or U4106 (N_4106,N_3322,N_3821);
and U4107 (N_4107,N_3337,N_3291);
xnor U4108 (N_4108,N_3360,N_3631);
or U4109 (N_4109,N_3495,N_3331);
nor U4110 (N_4110,N_3542,N_3152);
xnor U4111 (N_4111,N_3153,N_3525);
nand U4112 (N_4112,N_3479,N_3526);
nor U4113 (N_4113,N_3296,N_3069);
or U4114 (N_4114,N_3309,N_3786);
nor U4115 (N_4115,N_3377,N_3941);
or U4116 (N_4116,N_3618,N_3090);
and U4117 (N_4117,N_3726,N_3626);
nor U4118 (N_4118,N_3809,N_3795);
xor U4119 (N_4119,N_3072,N_3838);
nor U4120 (N_4120,N_3728,N_3405);
xor U4121 (N_4121,N_3025,N_3582);
or U4122 (N_4122,N_3940,N_3052);
and U4123 (N_4123,N_3219,N_3516);
nand U4124 (N_4124,N_3753,N_3671);
or U4125 (N_4125,N_3009,N_3318);
xor U4126 (N_4126,N_3323,N_3594);
nor U4127 (N_4127,N_3675,N_3725);
nand U4128 (N_4128,N_3935,N_3999);
or U4129 (N_4129,N_3471,N_3747);
or U4130 (N_4130,N_3097,N_3710);
or U4131 (N_4131,N_3649,N_3282);
xnor U4132 (N_4132,N_3857,N_3470);
and U4133 (N_4133,N_3108,N_3648);
or U4134 (N_4134,N_3664,N_3727);
xnor U4135 (N_4135,N_3887,N_3363);
and U4136 (N_4136,N_3817,N_3736);
nand U4137 (N_4137,N_3254,N_3472);
nand U4138 (N_4138,N_3738,N_3442);
and U4139 (N_4139,N_3102,N_3659);
and U4140 (N_4140,N_3741,N_3981);
xnor U4141 (N_4141,N_3799,N_3200);
or U4142 (N_4142,N_3705,N_3011);
nor U4143 (N_4143,N_3368,N_3775);
nor U4144 (N_4144,N_3089,N_3499);
nor U4145 (N_4145,N_3580,N_3910);
and U4146 (N_4146,N_3238,N_3880);
xor U4147 (N_4147,N_3466,N_3157);
or U4148 (N_4148,N_3832,N_3702);
and U4149 (N_4149,N_3873,N_3708);
nor U4150 (N_4150,N_3426,N_3774);
and U4151 (N_4151,N_3845,N_3415);
nor U4152 (N_4152,N_3587,N_3693);
and U4153 (N_4153,N_3539,N_3719);
or U4154 (N_4154,N_3563,N_3765);
or U4155 (N_4155,N_3487,N_3481);
nor U4156 (N_4156,N_3703,N_3243);
or U4157 (N_4157,N_3257,N_3504);
or U4158 (N_4158,N_3085,N_3171);
or U4159 (N_4159,N_3637,N_3225);
nand U4160 (N_4160,N_3432,N_3757);
nor U4161 (N_4161,N_3875,N_3537);
nand U4162 (N_4162,N_3541,N_3158);
nor U4163 (N_4163,N_3742,N_3139);
and U4164 (N_4164,N_3297,N_3602);
and U4165 (N_4165,N_3983,N_3364);
and U4166 (N_4166,N_3810,N_3691);
nand U4167 (N_4167,N_3801,N_3914);
xor U4168 (N_4168,N_3790,N_3656);
or U4169 (N_4169,N_3685,N_3482);
xor U4170 (N_4170,N_3262,N_3686);
or U4171 (N_4171,N_3333,N_3054);
and U4172 (N_4172,N_3572,N_3419);
nand U4173 (N_4173,N_3651,N_3555);
or U4174 (N_4174,N_3247,N_3294);
and U4175 (N_4175,N_3070,N_3724);
xnor U4176 (N_4176,N_3975,N_3589);
nand U4177 (N_4177,N_3925,N_3942);
or U4178 (N_4178,N_3369,N_3055);
xor U4179 (N_4179,N_3561,N_3167);
xor U4180 (N_4180,N_3111,N_3982);
nand U4181 (N_4181,N_3899,N_3916);
nand U4182 (N_4182,N_3173,N_3657);
nor U4183 (N_4183,N_3529,N_3400);
and U4184 (N_4184,N_3452,N_3199);
nor U4185 (N_4185,N_3755,N_3266);
xnor U4186 (N_4186,N_3937,N_3444);
nor U4187 (N_4187,N_3240,N_3943);
or U4188 (N_4188,N_3934,N_3127);
xnor U4189 (N_4189,N_3994,N_3635);
or U4190 (N_4190,N_3928,N_3978);
xor U4191 (N_4191,N_3796,N_3966);
nor U4192 (N_4192,N_3739,N_3087);
xnor U4193 (N_4193,N_3386,N_3279);
nand U4194 (N_4194,N_3763,N_3315);
nor U4195 (N_4195,N_3559,N_3132);
nand U4196 (N_4196,N_3397,N_3335);
xor U4197 (N_4197,N_3113,N_3803);
and U4198 (N_4198,N_3455,N_3798);
or U4199 (N_4199,N_3460,N_3996);
or U4200 (N_4200,N_3105,N_3096);
and U4201 (N_4201,N_3032,N_3987);
or U4202 (N_4202,N_3290,N_3141);
nor U4203 (N_4203,N_3438,N_3958);
xor U4204 (N_4204,N_3418,N_3359);
and U4205 (N_4205,N_3372,N_3729);
and U4206 (N_4206,N_3036,N_3258);
or U4207 (N_4207,N_3092,N_3647);
nand U4208 (N_4208,N_3867,N_3713);
xnor U4209 (N_4209,N_3010,N_3574);
and U4210 (N_4210,N_3136,N_3061);
xnor U4211 (N_4211,N_3365,N_3284);
xor U4212 (N_4212,N_3142,N_3027);
nor U4213 (N_4213,N_3998,N_3417);
xor U4214 (N_4214,N_3163,N_3450);
or U4215 (N_4215,N_3130,N_3303);
nor U4216 (N_4216,N_3610,N_3362);
xnor U4217 (N_4217,N_3669,N_3864);
nand U4218 (N_4218,N_3004,N_3678);
and U4219 (N_4219,N_3245,N_3016);
xnor U4220 (N_4220,N_3546,N_3062);
and U4221 (N_4221,N_3381,N_3298);
and U4222 (N_4222,N_3921,N_3552);
xnor U4223 (N_4223,N_3039,N_3850);
nor U4224 (N_4224,N_3847,N_3672);
nand U4225 (N_4225,N_3906,N_3962);
nand U4226 (N_4226,N_3249,N_3586);
xnor U4227 (N_4227,N_3890,N_3338);
or U4228 (N_4228,N_3094,N_3330);
or U4229 (N_4229,N_3776,N_3184);
xor U4230 (N_4230,N_3474,N_3512);
nor U4231 (N_4231,N_3506,N_3128);
xnor U4232 (N_4232,N_3517,N_3215);
or U4233 (N_4233,N_3929,N_3042);
nor U4234 (N_4234,N_3344,N_3353);
and U4235 (N_4235,N_3501,N_3289);
nor U4236 (N_4236,N_3980,N_3046);
nand U4237 (N_4237,N_3679,N_3723);
xnor U4238 (N_4238,N_3411,N_3737);
nor U4239 (N_4239,N_3006,N_3144);
nand U4240 (N_4240,N_3783,N_3545);
nor U4241 (N_4241,N_3558,N_3608);
nand U4242 (N_4242,N_3860,N_3868);
nor U4243 (N_4243,N_3049,N_3876);
and U4244 (N_4244,N_3782,N_3835);
nand U4245 (N_4245,N_3424,N_3456);
and U4246 (N_4246,N_3399,N_3091);
and U4247 (N_4247,N_3410,N_3402);
nand U4248 (N_4248,N_3837,N_3104);
and U4249 (N_4249,N_3878,N_3483);
nand U4250 (N_4250,N_3079,N_3217);
and U4251 (N_4251,N_3480,N_3661);
and U4252 (N_4252,N_3858,N_3473);
or U4253 (N_4253,N_3469,N_3175);
and U4254 (N_4254,N_3636,N_3412);
or U4255 (N_4255,N_3993,N_3073);
and U4256 (N_4256,N_3492,N_3242);
or U4257 (N_4257,N_3885,N_3274);
xnor U4258 (N_4258,N_3320,N_3750);
nor U4259 (N_4259,N_3148,N_3853);
and U4260 (N_4260,N_3192,N_3989);
and U4261 (N_4261,N_3521,N_3021);
nor U4262 (N_4262,N_3735,N_3390);
or U4263 (N_4263,N_3683,N_3214);
nor U4264 (N_4264,N_3267,N_3423);
xor U4265 (N_4265,N_3273,N_3047);
or U4266 (N_4266,N_3646,N_3960);
nand U4267 (N_4267,N_3232,N_3893);
xor U4268 (N_4268,N_3311,N_3121);
or U4269 (N_4269,N_3324,N_3556);
or U4270 (N_4270,N_3712,N_3917);
nand U4271 (N_4271,N_3038,N_3743);
or U4272 (N_4272,N_3454,N_3909);
or U4273 (N_4273,N_3869,N_3900);
nand U4274 (N_4274,N_3627,N_3644);
nor U4275 (N_4275,N_3446,N_3371);
and U4276 (N_4276,N_3566,N_3908);
xor U4277 (N_4277,N_3677,N_3448);
xor U4278 (N_4278,N_3302,N_3462);
nand U4279 (N_4279,N_3008,N_3204);
nand U4280 (N_4280,N_3293,N_3147);
and U4281 (N_4281,N_3547,N_3787);
nor U4282 (N_4282,N_3385,N_3319);
nand U4283 (N_4283,N_3325,N_3203);
xnor U4284 (N_4284,N_3491,N_3905);
and U4285 (N_4285,N_3391,N_3565);
or U4286 (N_4286,N_3828,N_3932);
xor U4287 (N_4287,N_3918,N_3388);
or U4288 (N_4288,N_3031,N_3532);
and U4289 (N_4289,N_3575,N_3334);
nand U4290 (N_4290,N_3907,N_3414);
and U4291 (N_4291,N_3189,N_3475);
or U4292 (N_4292,N_3652,N_3676);
xor U4293 (N_4293,N_3990,N_3550);
nand U4294 (N_4294,N_3126,N_3241);
nand U4295 (N_4295,N_3856,N_3896);
nand U4296 (N_4296,N_3510,N_3985);
or U4297 (N_4297,N_3224,N_3201);
or U4298 (N_4298,N_3272,N_3564);
or U4299 (N_4299,N_3433,N_3490);
xnor U4300 (N_4300,N_3100,N_3894);
nand U4301 (N_4301,N_3308,N_3922);
and U4302 (N_4302,N_3328,N_3083);
nor U4303 (N_4303,N_3784,N_3955);
nand U4304 (N_4304,N_3058,N_3361);
xor U4305 (N_4305,N_3508,N_3785);
nand U4306 (N_4306,N_3305,N_3680);
xor U4307 (N_4307,N_3053,N_3196);
nand U4308 (N_4308,N_3711,N_3409);
and U4309 (N_4309,N_3179,N_3430);
nor U4310 (N_4310,N_3768,N_3716);
nand U4311 (N_4311,N_3051,N_3329);
and U4312 (N_4312,N_3700,N_3746);
nand U4313 (N_4313,N_3265,N_3854);
nor U4314 (N_4314,N_3221,N_3903);
xor U4315 (N_4315,N_3295,N_3063);
nand U4316 (N_4316,N_3749,N_3769);
nor U4317 (N_4317,N_3355,N_3263);
nand U4318 (N_4318,N_3098,N_3269);
xnor U4319 (N_4319,N_3706,N_3172);
xnor U4320 (N_4320,N_3468,N_3948);
or U4321 (N_4321,N_3453,N_3115);
nand U4322 (N_4322,N_3692,N_3476);
nand U4323 (N_4323,N_3464,N_3614);
and U4324 (N_4324,N_3939,N_3522);
nor U4325 (N_4325,N_3045,N_3314);
and U4326 (N_4326,N_3270,N_3543);
xnor U4327 (N_4327,N_3957,N_3839);
or U4328 (N_4328,N_3041,N_3000);
nor U4329 (N_4329,N_3326,N_3946);
xnor U4330 (N_4330,N_3814,N_3502);
nand U4331 (N_4331,N_3252,N_3159);
nor U4332 (N_4332,N_3513,N_3968);
xnor U4333 (N_4333,N_3235,N_3065);
nor U4334 (N_4334,N_3034,N_3953);
nor U4335 (N_4335,N_3124,N_3924);
or U4336 (N_4336,N_3250,N_3779);
or U4337 (N_4337,N_3744,N_3441);
and U4338 (N_4338,N_3223,N_3855);
nand U4339 (N_4339,N_3398,N_3264);
xnor U4340 (N_4340,N_3578,N_3699);
or U4341 (N_4341,N_3299,N_3979);
nor U4342 (N_4342,N_3500,N_3086);
and U4343 (N_4343,N_3904,N_3503);
and U4344 (N_4344,N_3288,N_3458);
nand U4345 (N_4345,N_3913,N_3001);
nor U4346 (N_4346,N_3155,N_3959);
or U4347 (N_4347,N_3222,N_3228);
and U4348 (N_4348,N_3628,N_3133);
xor U4349 (N_4349,N_3285,N_3622);
xor U4350 (N_4350,N_3177,N_3780);
and U4351 (N_4351,N_3135,N_3275);
xnor U4352 (N_4352,N_3033,N_3843);
nand U4353 (N_4353,N_3681,N_3781);
and U4354 (N_4354,N_3689,N_3237);
nor U4355 (N_4355,N_3963,N_3816);
nand U4356 (N_4356,N_3081,N_3745);
or U4357 (N_4357,N_3920,N_3407);
nand U4358 (N_4358,N_3778,N_3349);
nand U4359 (N_4359,N_3493,N_3212);
or U4360 (N_4360,N_3117,N_3339);
and U4361 (N_4361,N_3892,N_3463);
xnor U4362 (N_4362,N_3457,N_3600);
or U4363 (N_4363,N_3343,N_3256);
xor U4364 (N_4364,N_3771,N_3760);
or U4365 (N_4365,N_3641,N_3352);
nand U4366 (N_4366,N_3088,N_3733);
xnor U4367 (N_4367,N_3536,N_3883);
and U4368 (N_4368,N_3327,N_3310);
nand U4369 (N_4369,N_3740,N_3514);
and U4370 (N_4370,N_3478,N_3557);
nand U4371 (N_4371,N_3110,N_3413);
xnor U4372 (N_4372,N_3891,N_3926);
nand U4373 (N_4373,N_3292,N_3422);
xor U4374 (N_4374,N_3420,N_3938);
or U4375 (N_4375,N_3554,N_3183);
nor U4376 (N_4376,N_3066,N_3278);
nand U4377 (N_4377,N_3251,N_3571);
xnor U4378 (N_4378,N_3766,N_3181);
nand U4379 (N_4379,N_3840,N_3825);
xnor U4380 (N_4380,N_3897,N_3013);
nand U4381 (N_4381,N_3612,N_3865);
and U4382 (N_4382,N_3380,N_3317);
nand U4383 (N_4383,N_3174,N_3849);
xor U4384 (N_4384,N_3528,N_3350);
and U4385 (N_4385,N_3149,N_3220);
nor U4386 (N_4386,N_3496,N_3300);
nand U4387 (N_4387,N_3965,N_3986);
or U4388 (N_4388,N_3901,N_3841);
nor U4389 (N_4389,N_3668,N_3028);
or U4390 (N_4390,N_3030,N_3666);
nor U4391 (N_4391,N_3118,N_3445);
nor U4392 (N_4392,N_3509,N_3176);
or U4393 (N_4393,N_3520,N_3103);
nor U4394 (N_4394,N_3375,N_3123);
or U4395 (N_4395,N_3698,N_3623);
and U4396 (N_4396,N_3342,N_3435);
or U4397 (N_4397,N_3597,N_3829);
xor U4398 (N_4398,N_3044,N_3800);
and U4399 (N_4399,N_3129,N_3277);
nor U4400 (N_4400,N_3788,N_3530);
nor U4401 (N_4401,N_3690,N_3673);
and U4402 (N_4402,N_3138,N_3367);
and U4403 (N_4403,N_3701,N_3515);
nor U4404 (N_4404,N_3588,N_3467);
or U4405 (N_4405,N_3347,N_3425);
xor U4406 (N_4406,N_3947,N_3188);
nor U4407 (N_4407,N_3567,N_3376);
nand U4408 (N_4408,N_3229,N_3560);
nand U4409 (N_4409,N_3684,N_3852);
nor U4410 (N_4410,N_3443,N_3059);
and U4411 (N_4411,N_3281,N_3003);
xor U4412 (N_4412,N_3773,N_3406);
or U4413 (N_4413,N_3593,N_3357);
xor U4414 (N_4414,N_3387,N_3161);
or U4415 (N_4415,N_3370,N_3078);
xnor U4416 (N_4416,N_3592,N_3316);
and U4417 (N_4417,N_3071,N_3606);
nor U4418 (N_4418,N_3396,N_3607);
nand U4419 (N_4419,N_3833,N_3169);
xnor U4420 (N_4420,N_3084,N_3806);
or U4421 (N_4421,N_3259,N_3662);
nand U4422 (N_4422,N_3544,N_3389);
nand U4423 (N_4423,N_3919,N_3872);
or U4424 (N_4424,N_3568,N_3972);
nor U4425 (N_4425,N_3548,N_3271);
nand U4426 (N_4426,N_3851,N_3643);
xnor U4427 (N_4427,N_3477,N_3178);
and U4428 (N_4428,N_3346,N_3859);
xor U4429 (N_4429,N_3764,N_3076);
nor U4430 (N_4430,N_3404,N_3634);
nand U4431 (N_4431,N_3498,N_3020);
nand U4432 (N_4432,N_3373,N_3812);
xor U4433 (N_4433,N_3107,N_3871);
nand U4434 (N_4434,N_3505,N_3603);
and U4435 (N_4435,N_3162,N_3286);
nand U4436 (N_4436,N_3082,N_3761);
or U4437 (N_4437,N_3944,N_3137);
and U4438 (N_4438,N_3754,N_3459);
nor U4439 (N_4439,N_3844,N_3239);
or U4440 (N_4440,N_3056,N_3336);
and U4441 (N_4441,N_3794,N_3616);
and U4442 (N_4442,N_3732,N_3120);
or U4443 (N_4443,N_3709,N_3226);
nand U4444 (N_4444,N_3625,N_3658);
nand U4445 (N_4445,N_3202,N_3306);
xor U4446 (N_4446,N_3465,N_3307);
or U4447 (N_4447,N_3704,N_3805);
nand U4448 (N_4448,N_3888,N_3074);
or U4449 (N_4449,N_3519,N_3416);
and U4450 (N_4450,N_3374,N_3758);
nor U4451 (N_4451,N_3260,N_3019);
or U4452 (N_4452,N_3437,N_3037);
xnor U4453 (N_4453,N_3640,N_3895);
xnor U4454 (N_4454,N_3624,N_3576);
or U4455 (N_4455,N_3154,N_3488);
nand U4456 (N_4456,N_3720,N_3898);
nor U4457 (N_4457,N_3112,N_3846);
and U4458 (N_4458,N_3881,N_3160);
or U4459 (N_4459,N_3394,N_3064);
nand U4460 (N_4460,N_3026,N_3802);
xor U4461 (N_4461,N_3598,N_3717);
and U4462 (N_4462,N_3822,N_3080);
and U4463 (N_4463,N_3807,N_3131);
or U4464 (N_4464,N_3345,N_3261);
and U4465 (N_4465,N_3630,N_3984);
or U4466 (N_4466,N_3762,N_3553);
nand U4467 (N_4467,N_3830,N_3077);
and U4468 (N_4468,N_3756,N_3332);
xor U4469 (N_4469,N_3449,N_3484);
xnor U4470 (N_4470,N_3879,N_3048);
xnor U4471 (N_4471,N_3974,N_3246);
and U4472 (N_4472,N_3949,N_3697);
and U4473 (N_4473,N_3789,N_3818);
or U4474 (N_4474,N_3877,N_3015);
nand U4475 (N_4475,N_3748,N_3599);
or U4476 (N_4476,N_3109,N_3497);
and U4477 (N_4477,N_3721,N_3461);
nand U4478 (N_4478,N_3767,N_3613);
nand U4479 (N_4479,N_3195,N_3182);
xor U4480 (N_4480,N_3234,N_3358);
and U4481 (N_4481,N_3518,N_3145);
nand U4482 (N_4482,N_3811,N_3831);
nand U4483 (N_4483,N_3834,N_3143);
xnor U4484 (N_4484,N_3538,N_3486);
and U4485 (N_4485,N_3002,N_3660);
nor U4486 (N_4486,N_3823,N_3125);
nor U4487 (N_4487,N_3383,N_3694);
or U4488 (N_4488,N_3590,N_3378);
nand U4489 (N_4489,N_3230,N_3170);
nand U4490 (N_4490,N_3403,N_3119);
or U4491 (N_4491,N_3207,N_3667);
nand U4492 (N_4492,N_3927,N_3995);
or U4493 (N_4493,N_3988,N_3068);
or U4494 (N_4494,N_3150,N_3751);
or U4495 (N_4495,N_3535,N_3902);
and U4496 (N_4496,N_3005,N_3609);
and U4497 (N_4497,N_3977,N_3485);
nor U4498 (N_4498,N_3866,N_3967);
nand U4499 (N_4499,N_3591,N_3696);
nor U4500 (N_4500,N_3495,N_3646);
nand U4501 (N_4501,N_3403,N_3330);
nor U4502 (N_4502,N_3982,N_3309);
and U4503 (N_4503,N_3404,N_3411);
or U4504 (N_4504,N_3835,N_3962);
and U4505 (N_4505,N_3585,N_3014);
xor U4506 (N_4506,N_3813,N_3415);
xor U4507 (N_4507,N_3493,N_3394);
nor U4508 (N_4508,N_3674,N_3500);
xor U4509 (N_4509,N_3428,N_3710);
nand U4510 (N_4510,N_3921,N_3417);
xor U4511 (N_4511,N_3608,N_3203);
or U4512 (N_4512,N_3245,N_3852);
and U4513 (N_4513,N_3638,N_3116);
nand U4514 (N_4514,N_3622,N_3571);
or U4515 (N_4515,N_3384,N_3085);
or U4516 (N_4516,N_3481,N_3108);
nand U4517 (N_4517,N_3696,N_3950);
xor U4518 (N_4518,N_3764,N_3724);
and U4519 (N_4519,N_3472,N_3966);
xor U4520 (N_4520,N_3419,N_3496);
nand U4521 (N_4521,N_3280,N_3868);
nor U4522 (N_4522,N_3181,N_3115);
xor U4523 (N_4523,N_3525,N_3632);
nand U4524 (N_4524,N_3967,N_3412);
and U4525 (N_4525,N_3973,N_3291);
and U4526 (N_4526,N_3220,N_3592);
or U4527 (N_4527,N_3866,N_3316);
and U4528 (N_4528,N_3938,N_3592);
nor U4529 (N_4529,N_3357,N_3168);
or U4530 (N_4530,N_3450,N_3997);
nor U4531 (N_4531,N_3516,N_3296);
xor U4532 (N_4532,N_3527,N_3992);
and U4533 (N_4533,N_3375,N_3314);
and U4534 (N_4534,N_3481,N_3619);
nand U4535 (N_4535,N_3691,N_3234);
or U4536 (N_4536,N_3182,N_3247);
nor U4537 (N_4537,N_3848,N_3761);
and U4538 (N_4538,N_3797,N_3505);
or U4539 (N_4539,N_3908,N_3857);
or U4540 (N_4540,N_3702,N_3222);
nand U4541 (N_4541,N_3974,N_3255);
or U4542 (N_4542,N_3914,N_3203);
xor U4543 (N_4543,N_3146,N_3296);
nand U4544 (N_4544,N_3410,N_3548);
or U4545 (N_4545,N_3302,N_3258);
and U4546 (N_4546,N_3416,N_3199);
nand U4547 (N_4547,N_3094,N_3815);
and U4548 (N_4548,N_3072,N_3873);
or U4549 (N_4549,N_3286,N_3157);
nor U4550 (N_4550,N_3005,N_3346);
and U4551 (N_4551,N_3178,N_3359);
or U4552 (N_4552,N_3946,N_3078);
or U4553 (N_4553,N_3229,N_3703);
and U4554 (N_4554,N_3524,N_3984);
nor U4555 (N_4555,N_3812,N_3399);
and U4556 (N_4556,N_3768,N_3441);
nor U4557 (N_4557,N_3750,N_3421);
nand U4558 (N_4558,N_3664,N_3402);
and U4559 (N_4559,N_3427,N_3345);
nor U4560 (N_4560,N_3456,N_3411);
nor U4561 (N_4561,N_3024,N_3134);
and U4562 (N_4562,N_3581,N_3809);
nor U4563 (N_4563,N_3977,N_3334);
nor U4564 (N_4564,N_3996,N_3852);
or U4565 (N_4565,N_3112,N_3858);
or U4566 (N_4566,N_3508,N_3618);
and U4567 (N_4567,N_3532,N_3811);
nor U4568 (N_4568,N_3156,N_3152);
xnor U4569 (N_4569,N_3598,N_3205);
nand U4570 (N_4570,N_3496,N_3066);
xor U4571 (N_4571,N_3139,N_3906);
nand U4572 (N_4572,N_3395,N_3653);
nand U4573 (N_4573,N_3714,N_3335);
and U4574 (N_4574,N_3701,N_3275);
nor U4575 (N_4575,N_3543,N_3154);
and U4576 (N_4576,N_3656,N_3965);
and U4577 (N_4577,N_3700,N_3364);
nor U4578 (N_4578,N_3562,N_3236);
nand U4579 (N_4579,N_3503,N_3279);
or U4580 (N_4580,N_3080,N_3598);
nor U4581 (N_4581,N_3586,N_3010);
and U4582 (N_4582,N_3566,N_3871);
nor U4583 (N_4583,N_3957,N_3636);
nand U4584 (N_4584,N_3420,N_3809);
xnor U4585 (N_4585,N_3652,N_3946);
xor U4586 (N_4586,N_3975,N_3149);
nor U4587 (N_4587,N_3343,N_3467);
xor U4588 (N_4588,N_3846,N_3332);
xnor U4589 (N_4589,N_3347,N_3988);
nor U4590 (N_4590,N_3319,N_3483);
and U4591 (N_4591,N_3074,N_3952);
or U4592 (N_4592,N_3369,N_3704);
nor U4593 (N_4593,N_3715,N_3928);
xor U4594 (N_4594,N_3337,N_3471);
nor U4595 (N_4595,N_3258,N_3092);
or U4596 (N_4596,N_3314,N_3744);
nor U4597 (N_4597,N_3537,N_3763);
nand U4598 (N_4598,N_3623,N_3695);
nand U4599 (N_4599,N_3421,N_3070);
or U4600 (N_4600,N_3882,N_3047);
and U4601 (N_4601,N_3473,N_3933);
and U4602 (N_4602,N_3656,N_3483);
xnor U4603 (N_4603,N_3308,N_3752);
nor U4604 (N_4604,N_3963,N_3949);
and U4605 (N_4605,N_3389,N_3003);
nand U4606 (N_4606,N_3986,N_3940);
or U4607 (N_4607,N_3557,N_3566);
xor U4608 (N_4608,N_3589,N_3844);
nand U4609 (N_4609,N_3035,N_3756);
xor U4610 (N_4610,N_3502,N_3158);
xnor U4611 (N_4611,N_3105,N_3820);
nand U4612 (N_4612,N_3990,N_3036);
nor U4613 (N_4613,N_3044,N_3825);
and U4614 (N_4614,N_3845,N_3260);
xnor U4615 (N_4615,N_3454,N_3487);
nand U4616 (N_4616,N_3118,N_3776);
nor U4617 (N_4617,N_3484,N_3644);
and U4618 (N_4618,N_3546,N_3442);
xnor U4619 (N_4619,N_3586,N_3401);
and U4620 (N_4620,N_3653,N_3423);
xnor U4621 (N_4621,N_3012,N_3281);
or U4622 (N_4622,N_3113,N_3065);
nor U4623 (N_4623,N_3425,N_3030);
or U4624 (N_4624,N_3332,N_3892);
xnor U4625 (N_4625,N_3415,N_3293);
nand U4626 (N_4626,N_3014,N_3690);
and U4627 (N_4627,N_3802,N_3282);
xnor U4628 (N_4628,N_3198,N_3894);
and U4629 (N_4629,N_3988,N_3425);
xnor U4630 (N_4630,N_3906,N_3386);
nand U4631 (N_4631,N_3032,N_3209);
or U4632 (N_4632,N_3456,N_3253);
nand U4633 (N_4633,N_3526,N_3646);
xnor U4634 (N_4634,N_3950,N_3475);
xnor U4635 (N_4635,N_3472,N_3484);
nand U4636 (N_4636,N_3696,N_3278);
and U4637 (N_4637,N_3622,N_3143);
xor U4638 (N_4638,N_3589,N_3704);
nand U4639 (N_4639,N_3936,N_3285);
and U4640 (N_4640,N_3980,N_3590);
nand U4641 (N_4641,N_3074,N_3213);
and U4642 (N_4642,N_3659,N_3214);
nand U4643 (N_4643,N_3264,N_3399);
and U4644 (N_4644,N_3055,N_3309);
xor U4645 (N_4645,N_3401,N_3404);
xor U4646 (N_4646,N_3473,N_3792);
nor U4647 (N_4647,N_3219,N_3268);
nand U4648 (N_4648,N_3381,N_3074);
or U4649 (N_4649,N_3959,N_3282);
xnor U4650 (N_4650,N_3853,N_3118);
xnor U4651 (N_4651,N_3614,N_3345);
nor U4652 (N_4652,N_3810,N_3588);
nor U4653 (N_4653,N_3761,N_3223);
and U4654 (N_4654,N_3813,N_3335);
or U4655 (N_4655,N_3218,N_3588);
xor U4656 (N_4656,N_3345,N_3240);
or U4657 (N_4657,N_3977,N_3293);
or U4658 (N_4658,N_3124,N_3941);
nor U4659 (N_4659,N_3344,N_3695);
or U4660 (N_4660,N_3689,N_3430);
and U4661 (N_4661,N_3860,N_3863);
nor U4662 (N_4662,N_3750,N_3558);
xnor U4663 (N_4663,N_3949,N_3277);
nor U4664 (N_4664,N_3046,N_3389);
nand U4665 (N_4665,N_3762,N_3053);
nand U4666 (N_4666,N_3129,N_3118);
or U4667 (N_4667,N_3948,N_3738);
or U4668 (N_4668,N_3709,N_3563);
xor U4669 (N_4669,N_3369,N_3737);
and U4670 (N_4670,N_3997,N_3984);
or U4671 (N_4671,N_3378,N_3910);
nor U4672 (N_4672,N_3578,N_3032);
xnor U4673 (N_4673,N_3187,N_3928);
nand U4674 (N_4674,N_3554,N_3593);
nor U4675 (N_4675,N_3478,N_3816);
or U4676 (N_4676,N_3906,N_3437);
and U4677 (N_4677,N_3616,N_3853);
and U4678 (N_4678,N_3827,N_3628);
xor U4679 (N_4679,N_3939,N_3368);
xnor U4680 (N_4680,N_3942,N_3462);
or U4681 (N_4681,N_3285,N_3327);
or U4682 (N_4682,N_3876,N_3411);
and U4683 (N_4683,N_3182,N_3786);
or U4684 (N_4684,N_3213,N_3091);
or U4685 (N_4685,N_3635,N_3196);
xor U4686 (N_4686,N_3435,N_3592);
or U4687 (N_4687,N_3695,N_3502);
nand U4688 (N_4688,N_3022,N_3014);
or U4689 (N_4689,N_3036,N_3125);
or U4690 (N_4690,N_3429,N_3136);
or U4691 (N_4691,N_3788,N_3806);
nand U4692 (N_4692,N_3741,N_3160);
or U4693 (N_4693,N_3531,N_3411);
or U4694 (N_4694,N_3877,N_3755);
nand U4695 (N_4695,N_3749,N_3629);
and U4696 (N_4696,N_3605,N_3926);
nor U4697 (N_4697,N_3451,N_3595);
nand U4698 (N_4698,N_3975,N_3087);
and U4699 (N_4699,N_3565,N_3052);
or U4700 (N_4700,N_3621,N_3995);
nand U4701 (N_4701,N_3149,N_3145);
nand U4702 (N_4702,N_3794,N_3008);
or U4703 (N_4703,N_3806,N_3254);
or U4704 (N_4704,N_3128,N_3919);
xnor U4705 (N_4705,N_3370,N_3787);
and U4706 (N_4706,N_3252,N_3751);
nor U4707 (N_4707,N_3550,N_3829);
nor U4708 (N_4708,N_3587,N_3867);
xor U4709 (N_4709,N_3352,N_3793);
nand U4710 (N_4710,N_3181,N_3635);
or U4711 (N_4711,N_3736,N_3102);
nand U4712 (N_4712,N_3749,N_3035);
and U4713 (N_4713,N_3626,N_3679);
and U4714 (N_4714,N_3146,N_3846);
nor U4715 (N_4715,N_3855,N_3171);
and U4716 (N_4716,N_3955,N_3554);
or U4717 (N_4717,N_3281,N_3336);
and U4718 (N_4718,N_3995,N_3151);
nor U4719 (N_4719,N_3540,N_3226);
nor U4720 (N_4720,N_3502,N_3135);
nand U4721 (N_4721,N_3447,N_3196);
xnor U4722 (N_4722,N_3684,N_3404);
and U4723 (N_4723,N_3704,N_3689);
and U4724 (N_4724,N_3187,N_3921);
and U4725 (N_4725,N_3853,N_3414);
xnor U4726 (N_4726,N_3637,N_3899);
xnor U4727 (N_4727,N_3339,N_3401);
and U4728 (N_4728,N_3470,N_3458);
nor U4729 (N_4729,N_3598,N_3426);
nand U4730 (N_4730,N_3598,N_3269);
nand U4731 (N_4731,N_3236,N_3827);
or U4732 (N_4732,N_3577,N_3337);
or U4733 (N_4733,N_3027,N_3549);
nor U4734 (N_4734,N_3780,N_3381);
xnor U4735 (N_4735,N_3470,N_3450);
or U4736 (N_4736,N_3569,N_3378);
nand U4737 (N_4737,N_3170,N_3314);
and U4738 (N_4738,N_3372,N_3281);
and U4739 (N_4739,N_3214,N_3918);
xnor U4740 (N_4740,N_3812,N_3277);
nand U4741 (N_4741,N_3271,N_3458);
or U4742 (N_4742,N_3251,N_3782);
and U4743 (N_4743,N_3809,N_3189);
and U4744 (N_4744,N_3061,N_3310);
or U4745 (N_4745,N_3775,N_3099);
or U4746 (N_4746,N_3476,N_3913);
xor U4747 (N_4747,N_3985,N_3341);
xor U4748 (N_4748,N_3962,N_3001);
nor U4749 (N_4749,N_3389,N_3531);
or U4750 (N_4750,N_3202,N_3863);
nor U4751 (N_4751,N_3829,N_3911);
nand U4752 (N_4752,N_3926,N_3228);
xnor U4753 (N_4753,N_3380,N_3517);
nand U4754 (N_4754,N_3890,N_3891);
and U4755 (N_4755,N_3089,N_3684);
and U4756 (N_4756,N_3935,N_3747);
nor U4757 (N_4757,N_3816,N_3614);
nor U4758 (N_4758,N_3538,N_3091);
nand U4759 (N_4759,N_3648,N_3057);
or U4760 (N_4760,N_3383,N_3385);
nor U4761 (N_4761,N_3003,N_3188);
or U4762 (N_4762,N_3970,N_3343);
or U4763 (N_4763,N_3005,N_3891);
nor U4764 (N_4764,N_3386,N_3657);
xor U4765 (N_4765,N_3497,N_3725);
or U4766 (N_4766,N_3643,N_3794);
nand U4767 (N_4767,N_3050,N_3624);
xor U4768 (N_4768,N_3427,N_3093);
nor U4769 (N_4769,N_3259,N_3529);
nand U4770 (N_4770,N_3547,N_3251);
and U4771 (N_4771,N_3498,N_3430);
or U4772 (N_4772,N_3079,N_3067);
nor U4773 (N_4773,N_3455,N_3076);
or U4774 (N_4774,N_3612,N_3583);
xnor U4775 (N_4775,N_3234,N_3904);
xnor U4776 (N_4776,N_3422,N_3813);
xor U4777 (N_4777,N_3122,N_3617);
nor U4778 (N_4778,N_3385,N_3640);
xor U4779 (N_4779,N_3778,N_3769);
or U4780 (N_4780,N_3160,N_3206);
nand U4781 (N_4781,N_3901,N_3203);
xnor U4782 (N_4782,N_3745,N_3797);
nand U4783 (N_4783,N_3544,N_3752);
xnor U4784 (N_4784,N_3110,N_3575);
or U4785 (N_4785,N_3603,N_3769);
nand U4786 (N_4786,N_3300,N_3930);
nor U4787 (N_4787,N_3300,N_3631);
and U4788 (N_4788,N_3116,N_3844);
or U4789 (N_4789,N_3327,N_3323);
xnor U4790 (N_4790,N_3051,N_3441);
xnor U4791 (N_4791,N_3845,N_3944);
nand U4792 (N_4792,N_3288,N_3317);
nand U4793 (N_4793,N_3091,N_3325);
or U4794 (N_4794,N_3535,N_3754);
nand U4795 (N_4795,N_3175,N_3126);
or U4796 (N_4796,N_3174,N_3952);
xnor U4797 (N_4797,N_3688,N_3642);
or U4798 (N_4798,N_3257,N_3387);
and U4799 (N_4799,N_3314,N_3055);
nand U4800 (N_4800,N_3778,N_3565);
nor U4801 (N_4801,N_3149,N_3517);
or U4802 (N_4802,N_3084,N_3079);
and U4803 (N_4803,N_3040,N_3522);
nor U4804 (N_4804,N_3394,N_3141);
nor U4805 (N_4805,N_3363,N_3655);
nor U4806 (N_4806,N_3372,N_3669);
or U4807 (N_4807,N_3096,N_3999);
xor U4808 (N_4808,N_3698,N_3932);
xnor U4809 (N_4809,N_3046,N_3901);
nor U4810 (N_4810,N_3458,N_3144);
xnor U4811 (N_4811,N_3911,N_3946);
and U4812 (N_4812,N_3778,N_3242);
and U4813 (N_4813,N_3928,N_3452);
nor U4814 (N_4814,N_3934,N_3853);
xor U4815 (N_4815,N_3860,N_3208);
and U4816 (N_4816,N_3857,N_3104);
xor U4817 (N_4817,N_3073,N_3316);
nor U4818 (N_4818,N_3769,N_3903);
nor U4819 (N_4819,N_3853,N_3686);
nand U4820 (N_4820,N_3636,N_3048);
nor U4821 (N_4821,N_3538,N_3601);
nand U4822 (N_4822,N_3729,N_3262);
nor U4823 (N_4823,N_3570,N_3461);
and U4824 (N_4824,N_3184,N_3277);
nor U4825 (N_4825,N_3355,N_3504);
nor U4826 (N_4826,N_3660,N_3822);
nand U4827 (N_4827,N_3632,N_3694);
xnor U4828 (N_4828,N_3431,N_3710);
or U4829 (N_4829,N_3501,N_3700);
nand U4830 (N_4830,N_3687,N_3376);
xor U4831 (N_4831,N_3103,N_3427);
nand U4832 (N_4832,N_3333,N_3755);
or U4833 (N_4833,N_3253,N_3363);
and U4834 (N_4834,N_3154,N_3242);
and U4835 (N_4835,N_3757,N_3380);
nand U4836 (N_4836,N_3012,N_3312);
xnor U4837 (N_4837,N_3040,N_3302);
and U4838 (N_4838,N_3739,N_3717);
and U4839 (N_4839,N_3501,N_3849);
and U4840 (N_4840,N_3058,N_3093);
nand U4841 (N_4841,N_3543,N_3366);
or U4842 (N_4842,N_3467,N_3459);
nand U4843 (N_4843,N_3456,N_3218);
xor U4844 (N_4844,N_3596,N_3545);
and U4845 (N_4845,N_3572,N_3137);
nor U4846 (N_4846,N_3758,N_3590);
nor U4847 (N_4847,N_3241,N_3356);
and U4848 (N_4848,N_3859,N_3496);
xnor U4849 (N_4849,N_3742,N_3252);
and U4850 (N_4850,N_3883,N_3283);
or U4851 (N_4851,N_3559,N_3064);
and U4852 (N_4852,N_3243,N_3625);
xor U4853 (N_4853,N_3439,N_3166);
nand U4854 (N_4854,N_3910,N_3205);
xor U4855 (N_4855,N_3663,N_3101);
and U4856 (N_4856,N_3354,N_3276);
nand U4857 (N_4857,N_3164,N_3715);
nand U4858 (N_4858,N_3337,N_3260);
nand U4859 (N_4859,N_3422,N_3731);
nor U4860 (N_4860,N_3575,N_3990);
or U4861 (N_4861,N_3476,N_3721);
or U4862 (N_4862,N_3382,N_3595);
nand U4863 (N_4863,N_3077,N_3073);
or U4864 (N_4864,N_3240,N_3469);
nand U4865 (N_4865,N_3731,N_3255);
nand U4866 (N_4866,N_3831,N_3141);
or U4867 (N_4867,N_3289,N_3693);
xor U4868 (N_4868,N_3674,N_3579);
nand U4869 (N_4869,N_3112,N_3217);
or U4870 (N_4870,N_3037,N_3718);
nand U4871 (N_4871,N_3442,N_3671);
nor U4872 (N_4872,N_3143,N_3589);
nor U4873 (N_4873,N_3354,N_3147);
nor U4874 (N_4874,N_3368,N_3530);
nor U4875 (N_4875,N_3025,N_3808);
xnor U4876 (N_4876,N_3167,N_3925);
nor U4877 (N_4877,N_3822,N_3884);
xnor U4878 (N_4878,N_3054,N_3822);
nor U4879 (N_4879,N_3415,N_3902);
nor U4880 (N_4880,N_3536,N_3382);
xor U4881 (N_4881,N_3470,N_3824);
xnor U4882 (N_4882,N_3508,N_3231);
and U4883 (N_4883,N_3342,N_3792);
nor U4884 (N_4884,N_3870,N_3025);
xnor U4885 (N_4885,N_3162,N_3741);
nand U4886 (N_4886,N_3070,N_3075);
xor U4887 (N_4887,N_3333,N_3652);
nand U4888 (N_4888,N_3037,N_3405);
nor U4889 (N_4889,N_3684,N_3460);
xnor U4890 (N_4890,N_3628,N_3178);
and U4891 (N_4891,N_3959,N_3232);
nand U4892 (N_4892,N_3895,N_3931);
or U4893 (N_4893,N_3536,N_3188);
and U4894 (N_4894,N_3783,N_3284);
or U4895 (N_4895,N_3182,N_3646);
and U4896 (N_4896,N_3181,N_3488);
or U4897 (N_4897,N_3628,N_3015);
nand U4898 (N_4898,N_3219,N_3439);
and U4899 (N_4899,N_3597,N_3718);
nand U4900 (N_4900,N_3428,N_3079);
nand U4901 (N_4901,N_3277,N_3449);
and U4902 (N_4902,N_3611,N_3516);
nor U4903 (N_4903,N_3470,N_3383);
nand U4904 (N_4904,N_3733,N_3189);
and U4905 (N_4905,N_3378,N_3718);
and U4906 (N_4906,N_3929,N_3437);
or U4907 (N_4907,N_3021,N_3834);
nand U4908 (N_4908,N_3563,N_3554);
or U4909 (N_4909,N_3430,N_3747);
xor U4910 (N_4910,N_3640,N_3219);
and U4911 (N_4911,N_3162,N_3501);
and U4912 (N_4912,N_3773,N_3045);
nor U4913 (N_4913,N_3549,N_3858);
nor U4914 (N_4914,N_3778,N_3572);
or U4915 (N_4915,N_3716,N_3994);
nand U4916 (N_4916,N_3821,N_3956);
xnor U4917 (N_4917,N_3953,N_3414);
nand U4918 (N_4918,N_3038,N_3016);
nand U4919 (N_4919,N_3066,N_3418);
and U4920 (N_4920,N_3740,N_3635);
xnor U4921 (N_4921,N_3433,N_3621);
or U4922 (N_4922,N_3842,N_3336);
and U4923 (N_4923,N_3298,N_3499);
nor U4924 (N_4924,N_3843,N_3643);
nor U4925 (N_4925,N_3057,N_3745);
and U4926 (N_4926,N_3771,N_3775);
or U4927 (N_4927,N_3730,N_3231);
nor U4928 (N_4928,N_3902,N_3683);
xor U4929 (N_4929,N_3450,N_3824);
and U4930 (N_4930,N_3834,N_3825);
xnor U4931 (N_4931,N_3020,N_3961);
or U4932 (N_4932,N_3198,N_3161);
nand U4933 (N_4933,N_3503,N_3772);
nand U4934 (N_4934,N_3139,N_3806);
or U4935 (N_4935,N_3133,N_3001);
or U4936 (N_4936,N_3515,N_3920);
xnor U4937 (N_4937,N_3578,N_3775);
nand U4938 (N_4938,N_3202,N_3072);
nand U4939 (N_4939,N_3537,N_3072);
nand U4940 (N_4940,N_3465,N_3658);
nor U4941 (N_4941,N_3324,N_3208);
xor U4942 (N_4942,N_3334,N_3394);
and U4943 (N_4943,N_3526,N_3809);
or U4944 (N_4944,N_3171,N_3017);
or U4945 (N_4945,N_3375,N_3419);
nor U4946 (N_4946,N_3204,N_3821);
or U4947 (N_4947,N_3383,N_3666);
xnor U4948 (N_4948,N_3177,N_3378);
xnor U4949 (N_4949,N_3898,N_3342);
and U4950 (N_4950,N_3806,N_3306);
nand U4951 (N_4951,N_3210,N_3543);
xnor U4952 (N_4952,N_3458,N_3697);
nand U4953 (N_4953,N_3542,N_3297);
xor U4954 (N_4954,N_3919,N_3370);
or U4955 (N_4955,N_3126,N_3377);
nor U4956 (N_4956,N_3382,N_3870);
nand U4957 (N_4957,N_3284,N_3293);
nand U4958 (N_4958,N_3076,N_3797);
and U4959 (N_4959,N_3597,N_3583);
nor U4960 (N_4960,N_3827,N_3004);
nor U4961 (N_4961,N_3303,N_3986);
and U4962 (N_4962,N_3100,N_3218);
xor U4963 (N_4963,N_3909,N_3715);
and U4964 (N_4964,N_3283,N_3269);
nand U4965 (N_4965,N_3072,N_3174);
and U4966 (N_4966,N_3069,N_3432);
nand U4967 (N_4967,N_3167,N_3746);
or U4968 (N_4968,N_3078,N_3775);
and U4969 (N_4969,N_3355,N_3765);
or U4970 (N_4970,N_3046,N_3346);
nand U4971 (N_4971,N_3227,N_3612);
xnor U4972 (N_4972,N_3733,N_3033);
or U4973 (N_4973,N_3862,N_3502);
nor U4974 (N_4974,N_3602,N_3421);
nand U4975 (N_4975,N_3525,N_3947);
nand U4976 (N_4976,N_3726,N_3305);
nor U4977 (N_4977,N_3196,N_3472);
or U4978 (N_4978,N_3098,N_3956);
xor U4979 (N_4979,N_3001,N_3328);
or U4980 (N_4980,N_3703,N_3200);
nand U4981 (N_4981,N_3756,N_3819);
and U4982 (N_4982,N_3171,N_3401);
and U4983 (N_4983,N_3361,N_3151);
and U4984 (N_4984,N_3041,N_3179);
and U4985 (N_4985,N_3322,N_3593);
nand U4986 (N_4986,N_3922,N_3538);
or U4987 (N_4987,N_3065,N_3273);
and U4988 (N_4988,N_3227,N_3206);
nand U4989 (N_4989,N_3886,N_3288);
xnor U4990 (N_4990,N_3710,N_3119);
or U4991 (N_4991,N_3399,N_3894);
nor U4992 (N_4992,N_3396,N_3984);
or U4993 (N_4993,N_3569,N_3459);
nand U4994 (N_4994,N_3515,N_3714);
or U4995 (N_4995,N_3298,N_3214);
nor U4996 (N_4996,N_3161,N_3904);
nand U4997 (N_4997,N_3499,N_3492);
or U4998 (N_4998,N_3743,N_3283);
nand U4999 (N_4999,N_3936,N_3341);
and U5000 (N_5000,N_4807,N_4919);
nand U5001 (N_5001,N_4637,N_4423);
or U5002 (N_5002,N_4710,N_4259);
nor U5003 (N_5003,N_4439,N_4231);
nor U5004 (N_5004,N_4274,N_4188);
nor U5005 (N_5005,N_4918,N_4435);
or U5006 (N_5006,N_4263,N_4327);
or U5007 (N_5007,N_4788,N_4754);
or U5008 (N_5008,N_4258,N_4548);
xnor U5009 (N_5009,N_4238,N_4074);
nor U5010 (N_5010,N_4309,N_4532);
nor U5011 (N_5011,N_4154,N_4666);
xnor U5012 (N_5012,N_4393,N_4332);
and U5013 (N_5013,N_4727,N_4494);
nor U5014 (N_5014,N_4275,N_4511);
xor U5015 (N_5015,N_4976,N_4142);
nor U5016 (N_5016,N_4036,N_4159);
or U5017 (N_5017,N_4396,N_4767);
or U5018 (N_5018,N_4877,N_4001);
nand U5019 (N_5019,N_4051,N_4530);
nor U5020 (N_5020,N_4834,N_4146);
or U5021 (N_5021,N_4787,N_4007);
xor U5022 (N_5022,N_4640,N_4186);
nand U5023 (N_5023,N_4481,N_4264);
or U5024 (N_5024,N_4080,N_4639);
or U5025 (N_5025,N_4443,N_4453);
nand U5026 (N_5026,N_4362,N_4868);
and U5027 (N_5027,N_4971,N_4020);
and U5028 (N_5028,N_4909,N_4880);
and U5029 (N_5029,N_4827,N_4270);
and U5030 (N_5030,N_4706,N_4529);
nor U5031 (N_5031,N_4300,N_4345);
nor U5032 (N_5032,N_4504,N_4391);
or U5033 (N_5033,N_4670,N_4780);
xnor U5034 (N_5034,N_4601,N_4165);
and U5035 (N_5035,N_4024,N_4629);
xnor U5036 (N_5036,N_4568,N_4874);
nor U5037 (N_5037,N_4075,N_4506);
nor U5038 (N_5038,N_4779,N_4851);
xor U5039 (N_5039,N_4731,N_4552);
nor U5040 (N_5040,N_4286,N_4096);
or U5041 (N_5041,N_4943,N_4321);
xor U5042 (N_5042,N_4092,N_4658);
and U5043 (N_5043,N_4931,N_4041);
nor U5044 (N_5044,N_4246,N_4108);
and U5045 (N_5045,N_4642,N_4760);
nor U5046 (N_5046,N_4336,N_4355);
nor U5047 (N_5047,N_4324,N_4547);
nand U5048 (N_5048,N_4945,N_4408);
or U5049 (N_5049,N_4442,N_4955);
and U5050 (N_5050,N_4837,N_4800);
xnor U5051 (N_5051,N_4618,N_4312);
and U5052 (N_5052,N_4737,N_4215);
nor U5053 (N_5053,N_4615,N_4609);
nor U5054 (N_5054,N_4746,N_4383);
and U5055 (N_5055,N_4303,N_4052);
and U5056 (N_5056,N_4673,N_4112);
nand U5057 (N_5057,N_4822,N_4451);
nand U5058 (N_5058,N_4008,N_4645);
nor U5059 (N_5059,N_4330,N_4992);
nor U5060 (N_5060,N_4400,N_4516);
xnor U5061 (N_5061,N_4952,N_4221);
nand U5062 (N_5062,N_4891,N_4354);
or U5063 (N_5063,N_4683,N_4218);
nor U5064 (N_5064,N_4871,N_4241);
nand U5065 (N_5065,N_4331,N_4985);
and U5066 (N_5066,N_4882,N_4253);
and U5067 (N_5067,N_4464,N_4963);
or U5068 (N_5068,N_4729,N_4411);
nand U5069 (N_5069,N_4922,N_4693);
nor U5070 (N_5070,N_4082,N_4187);
nand U5071 (N_5071,N_4974,N_4026);
nor U5072 (N_5072,N_4098,N_4404);
or U5073 (N_5073,N_4541,N_4296);
or U5074 (N_5074,N_4424,N_4513);
nor U5075 (N_5075,N_4222,N_4197);
nand U5076 (N_5076,N_4009,N_4267);
nand U5077 (N_5077,N_4405,N_4755);
nor U5078 (N_5078,N_4695,N_4194);
nor U5079 (N_5079,N_4913,N_4198);
or U5080 (N_5080,N_4519,N_4703);
nor U5081 (N_5081,N_4826,N_4845);
nand U5082 (N_5082,N_4697,N_4564);
nor U5083 (N_5083,N_4229,N_4998);
nor U5084 (N_5084,N_4179,N_4230);
nand U5085 (N_5085,N_4203,N_4164);
nor U5086 (N_5086,N_4531,N_4722);
nand U5087 (N_5087,N_4941,N_4561);
and U5088 (N_5088,N_4557,N_4343);
nor U5089 (N_5089,N_4433,N_4589);
xor U5090 (N_5090,N_4202,N_4853);
or U5091 (N_5091,N_4757,N_4797);
or U5092 (N_5092,N_4820,N_4635);
or U5093 (N_5093,N_4338,N_4269);
nand U5094 (N_5094,N_4887,N_4386);
or U5095 (N_5095,N_4591,N_4223);
nand U5096 (N_5096,N_4518,N_4648);
and U5097 (N_5097,N_4682,N_4255);
or U5098 (N_5098,N_4058,N_4633);
and U5099 (N_5099,N_4091,N_4958);
and U5100 (N_5100,N_4875,N_4921);
xor U5101 (N_5101,N_4679,N_4720);
xor U5102 (N_5102,N_4749,N_4260);
nand U5103 (N_5103,N_4669,N_4342);
and U5104 (N_5104,N_4616,N_4782);
and U5105 (N_5105,N_4284,N_4212);
nand U5106 (N_5106,N_4016,N_4733);
and U5107 (N_5107,N_4103,N_4719);
and U5108 (N_5108,N_4527,N_4128);
and U5109 (N_5109,N_4276,N_4625);
and U5110 (N_5110,N_4297,N_4524);
nor U5111 (N_5111,N_4318,N_4996);
or U5112 (N_5112,N_4674,N_4018);
or U5113 (N_5113,N_4388,N_4378);
xnor U5114 (N_5114,N_4621,N_4774);
xnor U5115 (N_5115,N_4474,N_4569);
nor U5116 (N_5116,N_4975,N_4254);
or U5117 (N_5117,N_4499,N_4002);
xnor U5118 (N_5118,N_4023,N_4847);
or U5119 (N_5119,N_4725,N_4028);
xor U5120 (N_5120,N_4896,N_4636);
and U5121 (N_5121,N_4859,N_4039);
nand U5122 (N_5122,N_4129,N_4624);
and U5123 (N_5123,N_4649,N_4872);
xnor U5124 (N_5124,N_4910,N_4549);
xnor U5125 (N_5125,N_4619,N_4173);
or U5126 (N_5126,N_4661,N_4644);
and U5127 (N_5127,N_4415,N_4858);
xor U5128 (N_5128,N_4436,N_4938);
or U5129 (N_5129,N_4337,N_4614);
xor U5130 (N_5130,N_4145,N_4643);
xor U5131 (N_5131,N_4430,N_4956);
xnor U5132 (N_5132,N_4340,N_4207);
nor U5133 (N_5133,N_4457,N_4768);
nand U5134 (N_5134,N_4756,N_4984);
nand U5135 (N_5135,N_4503,N_4438);
nand U5136 (N_5136,N_4791,N_4929);
nand U5137 (N_5137,N_4521,N_4077);
xnor U5138 (N_5138,N_4397,N_4377);
nor U5139 (N_5139,N_4283,N_4116);
and U5140 (N_5140,N_4199,N_4361);
or U5141 (N_5141,N_4067,N_4470);
nor U5142 (N_5142,N_4533,N_4983);
nand U5143 (N_5143,N_4315,N_4884);
nor U5144 (N_5144,N_4599,N_4932);
nor U5145 (N_5145,N_4817,N_4209);
nor U5146 (N_5146,N_4565,N_4492);
nand U5147 (N_5147,N_4476,N_4402);
xnor U5148 (N_5148,N_4416,N_4831);
nor U5149 (N_5149,N_4803,N_4718);
xnor U5150 (N_5150,N_4449,N_4178);
xnor U5151 (N_5151,N_4429,N_4764);
nor U5152 (N_5152,N_4582,N_4546);
xnor U5153 (N_5153,N_4201,N_4678);
nand U5154 (N_5154,N_4814,N_4211);
or U5155 (N_5155,N_4395,N_4272);
or U5156 (N_5156,N_4551,N_4409);
nor U5157 (N_5157,N_4226,N_4627);
and U5158 (N_5158,N_4224,N_4789);
nand U5159 (N_5159,N_4192,N_4538);
nor U5160 (N_5160,N_4792,N_4843);
nor U5161 (N_5161,N_4256,N_4239);
nor U5162 (N_5162,N_4333,N_4182);
and U5163 (N_5163,N_4157,N_4371);
and U5164 (N_5164,N_4496,N_4497);
and U5165 (N_5165,N_4559,N_4364);
and U5166 (N_5166,N_4341,N_4195);
and U5167 (N_5167,N_4136,N_4988);
and U5168 (N_5168,N_4890,N_4328);
nor U5169 (N_5169,N_4765,N_4054);
or U5170 (N_5170,N_4786,N_4382);
nand U5171 (N_5171,N_4110,N_4581);
nor U5172 (N_5172,N_4857,N_4403);
xnor U5173 (N_5173,N_4596,N_4401);
and U5174 (N_5174,N_4536,N_4427);
or U5175 (N_5175,N_4964,N_4991);
nor U5176 (N_5176,N_4465,N_4268);
nor U5177 (N_5177,N_4721,N_4111);
or U5178 (N_5178,N_4204,N_4356);
nor U5179 (N_5179,N_4161,N_4942);
and U5180 (N_5180,N_4933,N_4227);
xnor U5181 (N_5181,N_4479,N_4773);
and U5182 (N_5182,N_4793,N_4808);
nor U5183 (N_5183,N_4713,N_4795);
nor U5184 (N_5184,N_4273,N_4978);
and U5185 (N_5185,N_4305,N_4667);
and U5186 (N_5186,N_4567,N_4243);
nor U5187 (N_5187,N_4593,N_4155);
or U5188 (N_5188,N_4486,N_4540);
xor U5189 (N_5189,N_4372,N_4171);
or U5190 (N_5190,N_4122,N_4245);
and U5191 (N_5191,N_4537,N_4135);
and U5192 (N_5192,N_4021,N_4612);
nor U5193 (N_5193,N_4707,N_4414);
xor U5194 (N_5194,N_4004,N_4708);
xor U5195 (N_5195,N_4118,N_4047);
nor U5196 (N_5196,N_4132,N_4189);
and U5197 (N_5197,N_4799,N_4630);
xnor U5198 (N_5198,N_4784,N_4698);
xor U5199 (N_5199,N_4883,N_4689);
nor U5200 (N_5200,N_4033,N_4855);
or U5201 (N_5201,N_4715,N_4937);
xor U5202 (N_5202,N_4390,N_4736);
and U5203 (N_5203,N_4291,N_4086);
nand U5204 (N_5204,N_4174,N_4545);
xnor U5205 (N_5205,N_4908,N_4282);
nand U5206 (N_5206,N_4448,N_4166);
nand U5207 (N_5207,N_4526,N_4761);
nand U5208 (N_5208,N_4989,N_4571);
nand U5209 (N_5209,N_4461,N_4995);
or U5210 (N_5210,N_4510,N_4700);
nor U5211 (N_5211,N_4322,N_4613);
nor U5212 (N_5212,N_4688,N_4592);
nor U5213 (N_5213,N_4830,N_4914);
or U5214 (N_5214,N_4158,N_4732);
xnor U5215 (N_5215,N_4452,N_4347);
and U5216 (N_5216,N_4946,N_4864);
nor U5217 (N_5217,N_4081,N_4957);
xor U5218 (N_5218,N_4980,N_4090);
and U5219 (N_5219,N_4894,N_4242);
or U5220 (N_5220,N_4570,N_4912);
xor U5221 (N_5221,N_4939,N_4346);
xnor U5222 (N_5222,N_4251,N_4394);
nand U5223 (N_5223,N_4917,N_4467);
and U5224 (N_5224,N_4063,N_4121);
nor U5225 (N_5225,N_4660,N_4087);
xnor U5226 (N_5226,N_4723,N_4664);
and U5227 (N_5227,N_4934,N_4078);
nor U5228 (N_5228,N_4953,N_4307);
and U5229 (N_5229,N_4901,N_4022);
xor U5230 (N_5230,N_4823,N_4233);
xnor U5231 (N_5231,N_4055,N_4576);
xnor U5232 (N_5232,N_4508,N_4102);
xnor U5233 (N_5233,N_4017,N_4359);
xor U5234 (N_5234,N_4480,N_4498);
or U5235 (N_5235,N_4056,N_4804);
and U5236 (N_5236,N_4954,N_4675);
or U5237 (N_5237,N_4100,N_4292);
nor U5238 (N_5238,N_4869,N_4595);
or U5239 (N_5239,N_4965,N_4131);
or U5240 (N_5240,N_4960,N_4515);
xor U5241 (N_5241,N_4025,N_4907);
xor U5242 (N_5242,N_4622,N_4947);
xor U5243 (N_5243,N_4994,N_4177);
and U5244 (N_5244,N_4728,N_4083);
and U5245 (N_5245,N_4176,N_4517);
xor U5246 (N_5246,N_4191,N_4902);
nor U5247 (N_5247,N_4073,N_4127);
and U5248 (N_5248,N_4387,N_4232);
xnor U5249 (N_5249,N_4316,N_4977);
nand U5250 (N_5250,N_4997,N_4865);
and U5251 (N_5251,N_4590,N_4419);
nor U5252 (N_5252,N_4167,N_4839);
xor U5253 (N_5253,N_4454,N_4878);
or U5254 (N_5254,N_4248,N_4088);
and U5255 (N_5255,N_4488,N_4069);
or U5256 (N_5256,N_4962,N_4811);
or U5257 (N_5257,N_4428,N_4420);
and U5258 (N_5258,N_4152,N_4717);
xnor U5259 (N_5259,N_4656,N_4329);
nor U5260 (N_5260,N_4586,N_4691);
nor U5261 (N_5261,N_4061,N_4425);
nand U5262 (N_5262,N_4062,N_4588);
and U5263 (N_5263,N_4308,N_4970);
and U5264 (N_5264,N_4969,N_4948);
xor U5265 (N_5265,N_4915,N_4860);
xor U5266 (N_5266,N_4287,N_4175);
and U5267 (N_5267,N_4072,N_4003);
nor U5268 (N_5268,N_4751,N_4841);
xnor U5269 (N_5269,N_4099,N_4353);
nand U5270 (N_5270,N_4213,N_4881);
nand U5271 (N_5271,N_4904,N_4348);
nand U5272 (N_5272,N_4846,N_4686);
nand U5273 (N_5273,N_4982,N_4898);
nand U5274 (N_5274,N_4575,N_4936);
and U5275 (N_5275,N_4631,N_4628);
nand U5276 (N_5276,N_4785,N_4577);
xnor U5277 (N_5277,N_4462,N_4863);
and U5278 (N_5278,N_4271,N_4893);
nor U5279 (N_5279,N_4876,N_4059);
or U5280 (N_5280,N_4665,N_4298);
or U5281 (N_5281,N_4641,N_4133);
xnor U5282 (N_5282,N_4279,N_4434);
xor U5283 (N_5283,N_4743,N_4472);
and U5284 (N_5284,N_4815,N_4240);
nor U5285 (N_5285,N_4469,N_4037);
nor U5286 (N_5286,N_4053,N_4999);
or U5287 (N_5287,N_4237,N_4745);
xor U5288 (N_5288,N_4852,N_4701);
nor U5289 (N_5289,N_4543,N_4357);
xor U5290 (N_5290,N_4185,N_4304);
nand U5291 (N_5291,N_4558,N_4873);
nand U5292 (N_5292,N_4770,N_4006);
or U5293 (N_5293,N_4854,N_4553);
and U5294 (N_5294,N_4038,N_4079);
nor U5295 (N_5295,N_4825,N_4200);
or U5296 (N_5296,N_4677,N_4801);
nor U5297 (N_5297,N_4832,N_4778);
or U5298 (N_5298,N_4542,N_4680);
and U5299 (N_5299,N_4013,N_4716);
and U5300 (N_5300,N_4153,N_4280);
xnor U5301 (N_5301,N_4911,N_4849);
nor U5302 (N_5302,N_4149,N_4810);
nor U5303 (N_5303,N_4375,N_4950);
and U5304 (N_5304,N_4306,N_4712);
nor U5305 (N_5305,N_4181,N_4012);
and U5306 (N_5306,N_4769,N_4216);
and U5307 (N_5307,N_4466,N_4651);
nor U5308 (N_5308,N_4489,N_4699);
xnor U5309 (N_5309,N_4335,N_4410);
or U5310 (N_5310,N_4011,N_4456);
or U5311 (N_5311,N_4889,N_4478);
nand U5312 (N_5312,N_4125,N_4587);
nor U5313 (N_5313,N_4668,N_4295);
and U5314 (N_5314,N_4603,N_4611);
nand U5315 (N_5315,N_4605,N_4490);
nand U5316 (N_5316,N_4487,N_4724);
nor U5317 (N_5317,N_4373,N_4030);
or U5318 (N_5318,N_4981,N_4663);
xor U5319 (N_5319,N_4119,N_4068);
nor U5320 (N_5320,N_4168,N_4608);
nor U5321 (N_5321,N_4585,N_4126);
or U5322 (N_5322,N_4406,N_4398);
or U5323 (N_5323,N_4836,N_4250);
and U5324 (N_5324,N_4654,N_4685);
xnor U5325 (N_5325,N_4326,N_4554);
nand U5326 (N_5326,N_4967,N_4535);
and U5327 (N_5327,N_4709,N_4702);
nand U5328 (N_5328,N_4010,N_4389);
nand U5329 (N_5329,N_4925,N_4225);
nand U5330 (N_5330,N_4899,N_4812);
nor U5331 (N_5331,N_4281,N_4838);
nand U5332 (N_5332,N_4109,N_4824);
xor U5333 (N_5333,N_4123,N_4446);
or U5334 (N_5334,N_4892,N_4562);
or U5335 (N_5335,N_4045,N_4106);
and U5336 (N_5336,N_4924,N_4450);
nor U5337 (N_5337,N_4048,N_4726);
nand U5338 (N_5338,N_4762,N_4520);
or U5339 (N_5339,N_4431,N_4502);
nor U5340 (N_5340,N_4818,N_4206);
xnor U5341 (N_5341,N_4060,N_4509);
and U5342 (N_5342,N_4501,N_4169);
nand U5343 (N_5343,N_4781,N_4217);
nand U5344 (N_5344,N_4319,N_4027);
or U5345 (N_5345,N_4042,N_4692);
xnor U5346 (N_5346,N_4150,N_4374);
and U5347 (N_5347,N_4987,N_4819);
and U5348 (N_5348,N_4783,N_4413);
or U5349 (N_5349,N_4927,N_4031);
nand U5350 (N_5350,N_4714,N_4370);
nand U5351 (N_5351,N_4655,N_4244);
or U5352 (N_5352,N_4311,N_4441);
xor U5353 (N_5353,N_4744,N_4813);
or U5354 (N_5354,N_4638,N_4228);
nor U5355 (N_5355,N_4445,N_4986);
nor U5356 (N_5356,N_4475,N_4437);
and U5357 (N_5357,N_4493,N_4935);
nor U5358 (N_5358,N_4285,N_4208);
nor U5359 (N_5359,N_4463,N_4634);
nand U5360 (N_5360,N_4339,N_4694);
nor U5361 (N_5361,N_4385,N_4358);
or U5362 (N_5362,N_4777,N_4951);
xnor U5363 (N_5363,N_4623,N_4742);
or U5364 (N_5364,N_4015,N_4866);
nand U5365 (N_5365,N_4289,N_4447);
and U5366 (N_5366,N_4104,N_4617);
xnor U5367 (N_5367,N_4138,N_4095);
nand U5368 (N_5368,N_4484,N_4426);
and U5369 (N_5369,N_4870,N_4580);
and U5370 (N_5370,N_4829,N_4848);
xor U5371 (N_5371,N_4930,N_4172);
or U5372 (N_5372,N_4966,N_4143);
nor U5373 (N_5373,N_4500,N_4560);
or U5374 (N_5374,N_4730,N_4805);
xor U5375 (N_5375,N_4076,N_4798);
xnor U5376 (N_5376,N_4886,N_4193);
or U5377 (N_5377,N_4990,N_4302);
nor U5378 (N_5378,N_4835,N_4584);
or U5379 (N_5379,N_4879,N_4662);
and U5380 (N_5380,N_4210,N_4763);
nand U5381 (N_5381,N_4771,N_4392);
and U5382 (N_5382,N_4294,N_4979);
or U5383 (N_5383,N_4905,N_4748);
or U5384 (N_5384,N_4170,N_4652);
or U5385 (N_5385,N_4514,N_4366);
nand U5386 (N_5386,N_4759,N_4632);
or U5387 (N_5387,N_4741,N_4850);
nor U5388 (N_5388,N_4190,N_4089);
nand U5389 (N_5389,N_4101,N_4626);
or U5390 (N_5390,N_4897,N_4029);
nand U5391 (N_5391,N_4120,N_4610);
or U5392 (N_5392,N_4035,N_4539);
nand U5393 (N_5393,N_4117,N_4566);
xor U5394 (N_5394,N_4459,N_4350);
or U5395 (N_5395,N_4418,N_4040);
nor U5396 (N_5396,N_4057,N_4512);
nand U5397 (N_5397,N_4816,N_4278);
nand U5398 (N_5398,N_4923,N_4766);
and U5399 (N_5399,N_4162,N_4473);
nand U5400 (N_5400,N_4252,N_4525);
xnor U5401 (N_5401,N_4365,N_4672);
nor U5402 (N_5402,N_4093,N_4050);
nand U5403 (N_5403,N_4114,N_4344);
xor U5404 (N_5404,N_4351,N_4944);
nand U5405 (N_5405,N_4180,N_4972);
or U5406 (N_5406,N_4650,N_4140);
nand U5407 (N_5407,N_4034,N_4758);
xnor U5408 (N_5408,N_4776,N_4468);
nand U5409 (N_5409,N_4184,N_4740);
nand U5410 (N_5410,N_4219,N_4477);
nand U5411 (N_5411,N_4113,N_4973);
and U5412 (N_5412,N_4115,N_4412);
or U5413 (N_5413,N_4070,N_4676);
nor U5414 (N_5414,N_4071,N_4750);
or U5415 (N_5415,N_4085,N_4097);
xnor U5416 (N_5416,N_4407,N_4363);
and U5417 (N_5417,N_4753,N_4043);
nor U5418 (N_5418,N_4705,N_4421);
xor U5419 (N_5419,N_4775,N_4735);
nor U5420 (N_5420,N_4888,N_4885);
nor U5421 (N_5421,N_4739,N_4014);
or U5422 (N_5422,N_4752,N_4861);
nor U5423 (N_5423,N_4594,N_4288);
nor U5424 (N_5424,N_4578,N_4968);
nand U5425 (N_5425,N_4368,N_4379);
nand U5426 (N_5426,N_4455,N_4507);
and U5427 (N_5427,N_4310,N_4606);
or U5428 (N_5428,N_4959,N_4840);
xor U5429 (N_5429,N_4137,N_4671);
xor U5430 (N_5430,N_4598,N_4065);
or U5431 (N_5431,N_4600,N_4380);
nand U5432 (N_5432,N_4044,N_4163);
and U5433 (N_5433,N_4597,N_4144);
or U5434 (N_5434,N_4471,N_4417);
nand U5435 (N_5435,N_4602,N_4659);
nand U5436 (N_5436,N_4794,N_4604);
nand U5437 (N_5437,N_4005,N_4066);
xor U5438 (N_5438,N_4928,N_4690);
or U5439 (N_5439,N_4993,N_4681);
nor U5440 (N_5440,N_4796,N_4105);
or U5441 (N_5441,N_4367,N_4842);
or U5442 (N_5442,N_4124,N_4563);
nand U5443 (N_5443,N_4360,N_4483);
or U5444 (N_5444,N_4139,N_4369);
nor U5445 (N_5445,N_4234,N_4828);
or U5446 (N_5446,N_4376,N_4903);
nand U5447 (N_5447,N_4747,N_4572);
nor U5448 (N_5448,N_4214,N_4019);
nor U5449 (N_5449,N_4647,N_4205);
or U5450 (N_5450,N_4916,N_4196);
and U5451 (N_5451,N_4049,N_4032);
and U5452 (N_5452,N_4352,N_4249);
or U5453 (N_5453,N_4064,N_4148);
and U5454 (N_5454,N_4528,N_4134);
or U5455 (N_5455,N_4574,N_4802);
nor U5456 (N_5456,N_4806,N_4550);
xor U5457 (N_5457,N_4940,N_4491);
or U5458 (N_5458,N_4949,N_4325);
nand U5459 (N_5459,N_4314,N_4607);
nor U5460 (N_5460,N_4301,N_4183);
xor U5461 (N_5461,N_4313,N_4856);
nand U5462 (N_5462,N_4809,N_4653);
xor U5463 (N_5463,N_4084,N_4257);
and U5464 (N_5464,N_4920,N_4147);
nor U5465 (N_5465,N_4220,N_4381);
or U5466 (N_5466,N_4247,N_4460);
and U5467 (N_5467,N_4000,N_4265);
nor U5468 (N_5468,N_4862,N_4151);
xor U5469 (N_5469,N_4687,N_4620);
or U5470 (N_5470,N_4734,N_4573);
and U5471 (N_5471,N_4833,N_4160);
nor U5472 (N_5472,N_4317,N_4556);
nand U5473 (N_5473,N_4349,N_4495);
and U5474 (N_5474,N_4646,N_4299);
nor U5475 (N_5475,N_4821,N_4900);
nand U5476 (N_5476,N_4440,N_4141);
or U5477 (N_5477,N_4867,N_4277);
nor U5478 (N_5478,N_4444,N_4579);
nor U5479 (N_5479,N_4290,N_4458);
nand U5480 (N_5480,N_4293,N_4534);
nand U5481 (N_5481,N_4704,N_4485);
xor U5482 (N_5482,N_4156,N_4384);
xor U5483 (N_5483,N_4926,N_4844);
xnor U5484 (N_5484,N_4235,N_4684);
and U5485 (N_5485,N_4522,N_4505);
and U5486 (N_5486,N_4790,N_4334);
xor U5487 (N_5487,N_4523,N_4772);
nand U5488 (N_5488,N_4657,N_4323);
or U5489 (N_5489,N_4236,N_4696);
xor U5490 (N_5490,N_4320,N_4482);
and U5491 (N_5491,N_4261,N_4094);
and U5492 (N_5492,N_4961,N_4046);
nor U5493 (N_5493,N_4432,N_4422);
xor U5494 (N_5494,N_4711,N_4130);
and U5495 (N_5495,N_4555,N_4262);
or U5496 (N_5496,N_4906,N_4583);
nor U5497 (N_5497,N_4107,N_4895);
and U5498 (N_5498,N_4544,N_4399);
xor U5499 (N_5499,N_4738,N_4266);
xor U5500 (N_5500,N_4728,N_4830);
nor U5501 (N_5501,N_4120,N_4471);
and U5502 (N_5502,N_4923,N_4142);
nor U5503 (N_5503,N_4127,N_4767);
nand U5504 (N_5504,N_4048,N_4691);
and U5505 (N_5505,N_4031,N_4378);
nor U5506 (N_5506,N_4035,N_4012);
or U5507 (N_5507,N_4576,N_4780);
and U5508 (N_5508,N_4126,N_4067);
nand U5509 (N_5509,N_4973,N_4404);
xnor U5510 (N_5510,N_4932,N_4564);
or U5511 (N_5511,N_4659,N_4495);
xor U5512 (N_5512,N_4500,N_4831);
nor U5513 (N_5513,N_4842,N_4518);
xor U5514 (N_5514,N_4609,N_4910);
and U5515 (N_5515,N_4919,N_4753);
and U5516 (N_5516,N_4549,N_4845);
xnor U5517 (N_5517,N_4953,N_4555);
and U5518 (N_5518,N_4051,N_4236);
or U5519 (N_5519,N_4152,N_4871);
and U5520 (N_5520,N_4908,N_4654);
nor U5521 (N_5521,N_4753,N_4678);
nand U5522 (N_5522,N_4617,N_4336);
nor U5523 (N_5523,N_4331,N_4326);
nor U5524 (N_5524,N_4047,N_4914);
nor U5525 (N_5525,N_4629,N_4081);
nor U5526 (N_5526,N_4288,N_4555);
or U5527 (N_5527,N_4202,N_4606);
and U5528 (N_5528,N_4660,N_4656);
xor U5529 (N_5529,N_4165,N_4906);
xnor U5530 (N_5530,N_4581,N_4550);
xnor U5531 (N_5531,N_4263,N_4808);
nor U5532 (N_5532,N_4391,N_4536);
nor U5533 (N_5533,N_4773,N_4170);
and U5534 (N_5534,N_4333,N_4617);
or U5535 (N_5535,N_4682,N_4403);
nor U5536 (N_5536,N_4113,N_4283);
or U5537 (N_5537,N_4864,N_4865);
nand U5538 (N_5538,N_4997,N_4756);
or U5539 (N_5539,N_4207,N_4298);
and U5540 (N_5540,N_4014,N_4276);
xor U5541 (N_5541,N_4654,N_4117);
or U5542 (N_5542,N_4152,N_4574);
and U5543 (N_5543,N_4574,N_4451);
or U5544 (N_5544,N_4217,N_4270);
nor U5545 (N_5545,N_4186,N_4972);
nand U5546 (N_5546,N_4192,N_4367);
and U5547 (N_5547,N_4681,N_4319);
or U5548 (N_5548,N_4076,N_4315);
nor U5549 (N_5549,N_4330,N_4715);
nand U5550 (N_5550,N_4733,N_4655);
or U5551 (N_5551,N_4450,N_4234);
or U5552 (N_5552,N_4066,N_4772);
nand U5553 (N_5553,N_4260,N_4118);
nand U5554 (N_5554,N_4777,N_4564);
nor U5555 (N_5555,N_4286,N_4940);
xnor U5556 (N_5556,N_4751,N_4567);
and U5557 (N_5557,N_4326,N_4577);
or U5558 (N_5558,N_4101,N_4560);
xor U5559 (N_5559,N_4499,N_4870);
nor U5560 (N_5560,N_4700,N_4637);
xor U5561 (N_5561,N_4444,N_4663);
or U5562 (N_5562,N_4738,N_4079);
xnor U5563 (N_5563,N_4201,N_4846);
and U5564 (N_5564,N_4777,N_4722);
nand U5565 (N_5565,N_4207,N_4076);
nor U5566 (N_5566,N_4741,N_4926);
or U5567 (N_5567,N_4512,N_4379);
nand U5568 (N_5568,N_4834,N_4006);
xor U5569 (N_5569,N_4866,N_4855);
nor U5570 (N_5570,N_4399,N_4963);
nand U5571 (N_5571,N_4976,N_4908);
nand U5572 (N_5572,N_4400,N_4869);
and U5573 (N_5573,N_4765,N_4886);
or U5574 (N_5574,N_4202,N_4509);
or U5575 (N_5575,N_4419,N_4629);
nand U5576 (N_5576,N_4623,N_4890);
xor U5577 (N_5577,N_4005,N_4663);
nor U5578 (N_5578,N_4779,N_4283);
xnor U5579 (N_5579,N_4007,N_4353);
and U5580 (N_5580,N_4068,N_4323);
xor U5581 (N_5581,N_4607,N_4977);
or U5582 (N_5582,N_4509,N_4176);
and U5583 (N_5583,N_4838,N_4014);
nor U5584 (N_5584,N_4911,N_4407);
nand U5585 (N_5585,N_4687,N_4268);
nand U5586 (N_5586,N_4777,N_4631);
xor U5587 (N_5587,N_4176,N_4805);
and U5588 (N_5588,N_4272,N_4176);
and U5589 (N_5589,N_4437,N_4927);
nand U5590 (N_5590,N_4163,N_4118);
nor U5591 (N_5591,N_4033,N_4143);
nand U5592 (N_5592,N_4066,N_4715);
or U5593 (N_5593,N_4288,N_4546);
nand U5594 (N_5594,N_4877,N_4104);
or U5595 (N_5595,N_4881,N_4135);
or U5596 (N_5596,N_4830,N_4176);
xnor U5597 (N_5597,N_4898,N_4422);
or U5598 (N_5598,N_4508,N_4684);
or U5599 (N_5599,N_4076,N_4531);
nor U5600 (N_5600,N_4588,N_4071);
and U5601 (N_5601,N_4075,N_4182);
nor U5602 (N_5602,N_4721,N_4962);
nand U5603 (N_5603,N_4548,N_4457);
and U5604 (N_5604,N_4827,N_4392);
nand U5605 (N_5605,N_4993,N_4309);
and U5606 (N_5606,N_4606,N_4704);
nand U5607 (N_5607,N_4925,N_4555);
or U5608 (N_5608,N_4125,N_4392);
and U5609 (N_5609,N_4884,N_4245);
or U5610 (N_5610,N_4688,N_4510);
nand U5611 (N_5611,N_4655,N_4515);
xnor U5612 (N_5612,N_4238,N_4480);
or U5613 (N_5613,N_4045,N_4467);
nor U5614 (N_5614,N_4543,N_4474);
or U5615 (N_5615,N_4063,N_4779);
or U5616 (N_5616,N_4207,N_4219);
nand U5617 (N_5617,N_4690,N_4530);
xor U5618 (N_5618,N_4489,N_4637);
and U5619 (N_5619,N_4444,N_4372);
and U5620 (N_5620,N_4908,N_4538);
nand U5621 (N_5621,N_4561,N_4395);
nand U5622 (N_5622,N_4250,N_4553);
and U5623 (N_5623,N_4318,N_4385);
nand U5624 (N_5624,N_4729,N_4795);
nor U5625 (N_5625,N_4912,N_4803);
nand U5626 (N_5626,N_4073,N_4542);
and U5627 (N_5627,N_4308,N_4602);
xnor U5628 (N_5628,N_4822,N_4853);
and U5629 (N_5629,N_4624,N_4130);
nor U5630 (N_5630,N_4396,N_4049);
or U5631 (N_5631,N_4077,N_4474);
or U5632 (N_5632,N_4112,N_4291);
nand U5633 (N_5633,N_4616,N_4545);
xor U5634 (N_5634,N_4105,N_4992);
xor U5635 (N_5635,N_4720,N_4525);
nand U5636 (N_5636,N_4089,N_4660);
or U5637 (N_5637,N_4884,N_4232);
or U5638 (N_5638,N_4133,N_4310);
xor U5639 (N_5639,N_4089,N_4854);
nor U5640 (N_5640,N_4334,N_4142);
and U5641 (N_5641,N_4585,N_4705);
and U5642 (N_5642,N_4673,N_4131);
xor U5643 (N_5643,N_4169,N_4812);
or U5644 (N_5644,N_4876,N_4367);
nand U5645 (N_5645,N_4313,N_4779);
or U5646 (N_5646,N_4665,N_4813);
or U5647 (N_5647,N_4482,N_4048);
xnor U5648 (N_5648,N_4831,N_4936);
or U5649 (N_5649,N_4678,N_4856);
xnor U5650 (N_5650,N_4962,N_4322);
or U5651 (N_5651,N_4277,N_4963);
nand U5652 (N_5652,N_4780,N_4459);
or U5653 (N_5653,N_4234,N_4985);
xor U5654 (N_5654,N_4163,N_4444);
and U5655 (N_5655,N_4447,N_4239);
and U5656 (N_5656,N_4526,N_4374);
xnor U5657 (N_5657,N_4378,N_4706);
nand U5658 (N_5658,N_4016,N_4936);
or U5659 (N_5659,N_4674,N_4316);
and U5660 (N_5660,N_4355,N_4305);
or U5661 (N_5661,N_4449,N_4988);
xor U5662 (N_5662,N_4614,N_4232);
and U5663 (N_5663,N_4081,N_4182);
or U5664 (N_5664,N_4184,N_4716);
nand U5665 (N_5665,N_4045,N_4068);
nor U5666 (N_5666,N_4783,N_4220);
nor U5667 (N_5667,N_4510,N_4237);
nor U5668 (N_5668,N_4527,N_4444);
nor U5669 (N_5669,N_4519,N_4924);
or U5670 (N_5670,N_4017,N_4867);
xor U5671 (N_5671,N_4953,N_4140);
nand U5672 (N_5672,N_4806,N_4997);
or U5673 (N_5673,N_4437,N_4133);
or U5674 (N_5674,N_4574,N_4504);
and U5675 (N_5675,N_4450,N_4878);
nand U5676 (N_5676,N_4891,N_4665);
and U5677 (N_5677,N_4615,N_4130);
xor U5678 (N_5678,N_4543,N_4337);
and U5679 (N_5679,N_4986,N_4388);
xnor U5680 (N_5680,N_4152,N_4325);
or U5681 (N_5681,N_4215,N_4375);
xnor U5682 (N_5682,N_4823,N_4472);
nor U5683 (N_5683,N_4049,N_4311);
and U5684 (N_5684,N_4395,N_4762);
and U5685 (N_5685,N_4764,N_4273);
or U5686 (N_5686,N_4420,N_4282);
xor U5687 (N_5687,N_4831,N_4289);
nand U5688 (N_5688,N_4349,N_4526);
nor U5689 (N_5689,N_4433,N_4791);
nand U5690 (N_5690,N_4506,N_4300);
xnor U5691 (N_5691,N_4595,N_4276);
and U5692 (N_5692,N_4614,N_4128);
and U5693 (N_5693,N_4823,N_4393);
nand U5694 (N_5694,N_4618,N_4119);
xor U5695 (N_5695,N_4442,N_4609);
or U5696 (N_5696,N_4581,N_4309);
nor U5697 (N_5697,N_4394,N_4023);
nand U5698 (N_5698,N_4218,N_4510);
or U5699 (N_5699,N_4490,N_4409);
nand U5700 (N_5700,N_4877,N_4223);
nand U5701 (N_5701,N_4028,N_4246);
and U5702 (N_5702,N_4160,N_4805);
and U5703 (N_5703,N_4930,N_4229);
nand U5704 (N_5704,N_4805,N_4258);
or U5705 (N_5705,N_4580,N_4791);
and U5706 (N_5706,N_4772,N_4392);
xnor U5707 (N_5707,N_4987,N_4316);
and U5708 (N_5708,N_4210,N_4208);
xor U5709 (N_5709,N_4599,N_4082);
nand U5710 (N_5710,N_4205,N_4890);
and U5711 (N_5711,N_4365,N_4314);
and U5712 (N_5712,N_4746,N_4657);
xnor U5713 (N_5713,N_4437,N_4664);
nand U5714 (N_5714,N_4387,N_4681);
xnor U5715 (N_5715,N_4740,N_4866);
nand U5716 (N_5716,N_4544,N_4517);
nor U5717 (N_5717,N_4372,N_4520);
xor U5718 (N_5718,N_4478,N_4515);
xnor U5719 (N_5719,N_4285,N_4949);
xnor U5720 (N_5720,N_4906,N_4613);
nand U5721 (N_5721,N_4212,N_4085);
and U5722 (N_5722,N_4317,N_4302);
and U5723 (N_5723,N_4570,N_4091);
xnor U5724 (N_5724,N_4583,N_4654);
nand U5725 (N_5725,N_4230,N_4368);
nor U5726 (N_5726,N_4940,N_4951);
or U5727 (N_5727,N_4474,N_4831);
nor U5728 (N_5728,N_4030,N_4556);
nand U5729 (N_5729,N_4014,N_4091);
nand U5730 (N_5730,N_4905,N_4639);
nor U5731 (N_5731,N_4678,N_4881);
nor U5732 (N_5732,N_4510,N_4371);
nor U5733 (N_5733,N_4892,N_4101);
or U5734 (N_5734,N_4125,N_4030);
nand U5735 (N_5735,N_4275,N_4734);
xnor U5736 (N_5736,N_4683,N_4854);
nand U5737 (N_5737,N_4870,N_4455);
and U5738 (N_5738,N_4784,N_4258);
nand U5739 (N_5739,N_4331,N_4413);
nand U5740 (N_5740,N_4790,N_4378);
and U5741 (N_5741,N_4686,N_4663);
xor U5742 (N_5742,N_4542,N_4033);
and U5743 (N_5743,N_4414,N_4737);
xnor U5744 (N_5744,N_4881,N_4046);
and U5745 (N_5745,N_4050,N_4340);
or U5746 (N_5746,N_4890,N_4137);
and U5747 (N_5747,N_4086,N_4407);
and U5748 (N_5748,N_4145,N_4060);
nor U5749 (N_5749,N_4900,N_4780);
nor U5750 (N_5750,N_4021,N_4906);
and U5751 (N_5751,N_4948,N_4424);
or U5752 (N_5752,N_4701,N_4417);
xor U5753 (N_5753,N_4854,N_4004);
nand U5754 (N_5754,N_4289,N_4549);
nand U5755 (N_5755,N_4533,N_4239);
xnor U5756 (N_5756,N_4423,N_4640);
nand U5757 (N_5757,N_4941,N_4918);
nand U5758 (N_5758,N_4294,N_4873);
nand U5759 (N_5759,N_4722,N_4986);
nor U5760 (N_5760,N_4449,N_4730);
nor U5761 (N_5761,N_4988,N_4465);
nor U5762 (N_5762,N_4205,N_4216);
nor U5763 (N_5763,N_4180,N_4808);
and U5764 (N_5764,N_4642,N_4315);
nor U5765 (N_5765,N_4764,N_4874);
and U5766 (N_5766,N_4334,N_4702);
nand U5767 (N_5767,N_4542,N_4277);
or U5768 (N_5768,N_4656,N_4021);
nor U5769 (N_5769,N_4276,N_4545);
nand U5770 (N_5770,N_4099,N_4919);
xor U5771 (N_5771,N_4691,N_4002);
xnor U5772 (N_5772,N_4880,N_4983);
xor U5773 (N_5773,N_4929,N_4843);
xor U5774 (N_5774,N_4044,N_4724);
nand U5775 (N_5775,N_4723,N_4895);
and U5776 (N_5776,N_4023,N_4257);
and U5777 (N_5777,N_4299,N_4682);
nor U5778 (N_5778,N_4977,N_4076);
nor U5779 (N_5779,N_4879,N_4016);
or U5780 (N_5780,N_4283,N_4730);
or U5781 (N_5781,N_4807,N_4401);
nor U5782 (N_5782,N_4929,N_4345);
nand U5783 (N_5783,N_4569,N_4798);
and U5784 (N_5784,N_4904,N_4810);
nor U5785 (N_5785,N_4163,N_4506);
and U5786 (N_5786,N_4388,N_4984);
nor U5787 (N_5787,N_4623,N_4424);
and U5788 (N_5788,N_4069,N_4612);
nand U5789 (N_5789,N_4843,N_4063);
nor U5790 (N_5790,N_4035,N_4407);
and U5791 (N_5791,N_4177,N_4963);
xor U5792 (N_5792,N_4630,N_4407);
xnor U5793 (N_5793,N_4731,N_4595);
xnor U5794 (N_5794,N_4484,N_4368);
and U5795 (N_5795,N_4064,N_4038);
and U5796 (N_5796,N_4770,N_4653);
or U5797 (N_5797,N_4072,N_4430);
and U5798 (N_5798,N_4353,N_4684);
and U5799 (N_5799,N_4773,N_4523);
nand U5800 (N_5800,N_4586,N_4147);
and U5801 (N_5801,N_4301,N_4843);
nand U5802 (N_5802,N_4206,N_4821);
or U5803 (N_5803,N_4991,N_4015);
xnor U5804 (N_5804,N_4761,N_4701);
nor U5805 (N_5805,N_4751,N_4415);
nor U5806 (N_5806,N_4972,N_4127);
and U5807 (N_5807,N_4107,N_4666);
nor U5808 (N_5808,N_4044,N_4191);
nand U5809 (N_5809,N_4113,N_4605);
nor U5810 (N_5810,N_4476,N_4185);
nor U5811 (N_5811,N_4872,N_4401);
nand U5812 (N_5812,N_4495,N_4459);
or U5813 (N_5813,N_4076,N_4547);
and U5814 (N_5814,N_4646,N_4398);
and U5815 (N_5815,N_4393,N_4756);
xnor U5816 (N_5816,N_4831,N_4681);
nand U5817 (N_5817,N_4096,N_4845);
and U5818 (N_5818,N_4010,N_4109);
nor U5819 (N_5819,N_4909,N_4803);
xnor U5820 (N_5820,N_4496,N_4736);
nand U5821 (N_5821,N_4850,N_4717);
nand U5822 (N_5822,N_4707,N_4515);
xnor U5823 (N_5823,N_4241,N_4918);
or U5824 (N_5824,N_4900,N_4665);
nor U5825 (N_5825,N_4006,N_4149);
xnor U5826 (N_5826,N_4209,N_4421);
or U5827 (N_5827,N_4240,N_4622);
xnor U5828 (N_5828,N_4885,N_4878);
xor U5829 (N_5829,N_4384,N_4336);
and U5830 (N_5830,N_4872,N_4416);
or U5831 (N_5831,N_4609,N_4390);
xor U5832 (N_5832,N_4520,N_4074);
and U5833 (N_5833,N_4623,N_4768);
xor U5834 (N_5834,N_4784,N_4318);
xnor U5835 (N_5835,N_4311,N_4144);
nor U5836 (N_5836,N_4384,N_4832);
and U5837 (N_5837,N_4497,N_4246);
or U5838 (N_5838,N_4996,N_4287);
nand U5839 (N_5839,N_4615,N_4119);
nand U5840 (N_5840,N_4423,N_4837);
xnor U5841 (N_5841,N_4650,N_4417);
nand U5842 (N_5842,N_4379,N_4698);
nor U5843 (N_5843,N_4941,N_4198);
xor U5844 (N_5844,N_4969,N_4177);
nor U5845 (N_5845,N_4637,N_4697);
and U5846 (N_5846,N_4899,N_4575);
nand U5847 (N_5847,N_4496,N_4768);
and U5848 (N_5848,N_4630,N_4160);
xnor U5849 (N_5849,N_4812,N_4589);
xnor U5850 (N_5850,N_4154,N_4069);
nor U5851 (N_5851,N_4797,N_4348);
or U5852 (N_5852,N_4480,N_4849);
or U5853 (N_5853,N_4132,N_4199);
nand U5854 (N_5854,N_4088,N_4312);
and U5855 (N_5855,N_4226,N_4277);
xnor U5856 (N_5856,N_4491,N_4265);
nor U5857 (N_5857,N_4889,N_4927);
nand U5858 (N_5858,N_4045,N_4086);
nor U5859 (N_5859,N_4185,N_4075);
nand U5860 (N_5860,N_4181,N_4837);
nand U5861 (N_5861,N_4791,N_4003);
nor U5862 (N_5862,N_4656,N_4045);
or U5863 (N_5863,N_4472,N_4739);
nor U5864 (N_5864,N_4532,N_4412);
or U5865 (N_5865,N_4699,N_4323);
or U5866 (N_5866,N_4278,N_4093);
nand U5867 (N_5867,N_4903,N_4306);
xnor U5868 (N_5868,N_4690,N_4846);
nor U5869 (N_5869,N_4338,N_4782);
nand U5870 (N_5870,N_4813,N_4408);
xor U5871 (N_5871,N_4697,N_4768);
xor U5872 (N_5872,N_4967,N_4136);
nor U5873 (N_5873,N_4027,N_4469);
nor U5874 (N_5874,N_4498,N_4729);
xor U5875 (N_5875,N_4567,N_4305);
or U5876 (N_5876,N_4153,N_4291);
nand U5877 (N_5877,N_4344,N_4624);
or U5878 (N_5878,N_4196,N_4708);
or U5879 (N_5879,N_4641,N_4225);
nor U5880 (N_5880,N_4494,N_4217);
xnor U5881 (N_5881,N_4799,N_4621);
xor U5882 (N_5882,N_4917,N_4598);
and U5883 (N_5883,N_4071,N_4014);
xor U5884 (N_5884,N_4176,N_4152);
and U5885 (N_5885,N_4436,N_4947);
or U5886 (N_5886,N_4450,N_4119);
or U5887 (N_5887,N_4922,N_4343);
xnor U5888 (N_5888,N_4937,N_4640);
and U5889 (N_5889,N_4671,N_4630);
xnor U5890 (N_5890,N_4821,N_4237);
or U5891 (N_5891,N_4465,N_4489);
or U5892 (N_5892,N_4557,N_4511);
and U5893 (N_5893,N_4475,N_4664);
and U5894 (N_5894,N_4222,N_4499);
xnor U5895 (N_5895,N_4886,N_4803);
nand U5896 (N_5896,N_4530,N_4440);
or U5897 (N_5897,N_4267,N_4948);
xnor U5898 (N_5898,N_4120,N_4968);
and U5899 (N_5899,N_4613,N_4583);
or U5900 (N_5900,N_4393,N_4672);
nor U5901 (N_5901,N_4223,N_4636);
nand U5902 (N_5902,N_4030,N_4349);
or U5903 (N_5903,N_4447,N_4445);
and U5904 (N_5904,N_4576,N_4586);
nand U5905 (N_5905,N_4474,N_4221);
nand U5906 (N_5906,N_4866,N_4707);
and U5907 (N_5907,N_4134,N_4822);
nand U5908 (N_5908,N_4638,N_4360);
nor U5909 (N_5909,N_4216,N_4867);
and U5910 (N_5910,N_4880,N_4065);
nor U5911 (N_5911,N_4982,N_4046);
nand U5912 (N_5912,N_4385,N_4742);
nor U5913 (N_5913,N_4136,N_4482);
and U5914 (N_5914,N_4453,N_4034);
and U5915 (N_5915,N_4231,N_4157);
and U5916 (N_5916,N_4642,N_4811);
and U5917 (N_5917,N_4703,N_4805);
nand U5918 (N_5918,N_4336,N_4340);
nand U5919 (N_5919,N_4223,N_4570);
or U5920 (N_5920,N_4937,N_4895);
nor U5921 (N_5921,N_4715,N_4048);
xor U5922 (N_5922,N_4274,N_4606);
or U5923 (N_5923,N_4795,N_4637);
xnor U5924 (N_5924,N_4168,N_4950);
nand U5925 (N_5925,N_4909,N_4683);
and U5926 (N_5926,N_4193,N_4138);
nand U5927 (N_5927,N_4061,N_4053);
xnor U5928 (N_5928,N_4039,N_4185);
or U5929 (N_5929,N_4044,N_4081);
and U5930 (N_5930,N_4860,N_4602);
and U5931 (N_5931,N_4977,N_4635);
and U5932 (N_5932,N_4231,N_4249);
nor U5933 (N_5933,N_4890,N_4577);
and U5934 (N_5934,N_4130,N_4159);
nand U5935 (N_5935,N_4915,N_4869);
and U5936 (N_5936,N_4166,N_4807);
and U5937 (N_5937,N_4219,N_4229);
and U5938 (N_5938,N_4255,N_4952);
and U5939 (N_5939,N_4370,N_4595);
nor U5940 (N_5940,N_4949,N_4954);
xor U5941 (N_5941,N_4683,N_4242);
or U5942 (N_5942,N_4267,N_4313);
and U5943 (N_5943,N_4228,N_4356);
nand U5944 (N_5944,N_4599,N_4128);
nor U5945 (N_5945,N_4344,N_4684);
nand U5946 (N_5946,N_4806,N_4628);
nor U5947 (N_5947,N_4917,N_4988);
nor U5948 (N_5948,N_4916,N_4439);
nor U5949 (N_5949,N_4450,N_4153);
nor U5950 (N_5950,N_4560,N_4910);
nand U5951 (N_5951,N_4613,N_4198);
or U5952 (N_5952,N_4881,N_4784);
nand U5953 (N_5953,N_4771,N_4233);
nand U5954 (N_5954,N_4298,N_4719);
nand U5955 (N_5955,N_4333,N_4829);
or U5956 (N_5956,N_4226,N_4000);
and U5957 (N_5957,N_4699,N_4120);
nand U5958 (N_5958,N_4890,N_4396);
or U5959 (N_5959,N_4478,N_4966);
and U5960 (N_5960,N_4121,N_4782);
xnor U5961 (N_5961,N_4066,N_4838);
nand U5962 (N_5962,N_4773,N_4986);
or U5963 (N_5963,N_4238,N_4126);
nand U5964 (N_5964,N_4939,N_4755);
and U5965 (N_5965,N_4371,N_4263);
or U5966 (N_5966,N_4843,N_4174);
or U5967 (N_5967,N_4087,N_4476);
and U5968 (N_5968,N_4719,N_4401);
or U5969 (N_5969,N_4605,N_4607);
xor U5970 (N_5970,N_4555,N_4263);
nor U5971 (N_5971,N_4808,N_4501);
xnor U5972 (N_5972,N_4191,N_4423);
or U5973 (N_5973,N_4765,N_4741);
nor U5974 (N_5974,N_4974,N_4341);
nor U5975 (N_5975,N_4581,N_4868);
or U5976 (N_5976,N_4961,N_4301);
nand U5977 (N_5977,N_4716,N_4251);
nand U5978 (N_5978,N_4036,N_4430);
or U5979 (N_5979,N_4957,N_4420);
nor U5980 (N_5980,N_4386,N_4192);
or U5981 (N_5981,N_4031,N_4795);
xor U5982 (N_5982,N_4960,N_4526);
nor U5983 (N_5983,N_4864,N_4907);
nand U5984 (N_5984,N_4850,N_4290);
xor U5985 (N_5985,N_4915,N_4293);
xnor U5986 (N_5986,N_4723,N_4629);
and U5987 (N_5987,N_4004,N_4740);
nand U5988 (N_5988,N_4210,N_4937);
nand U5989 (N_5989,N_4915,N_4312);
or U5990 (N_5990,N_4392,N_4179);
nor U5991 (N_5991,N_4685,N_4308);
or U5992 (N_5992,N_4578,N_4854);
and U5993 (N_5993,N_4670,N_4728);
or U5994 (N_5994,N_4481,N_4175);
and U5995 (N_5995,N_4928,N_4421);
nor U5996 (N_5996,N_4495,N_4080);
nor U5997 (N_5997,N_4155,N_4437);
nor U5998 (N_5998,N_4539,N_4812);
nor U5999 (N_5999,N_4799,N_4591);
and U6000 (N_6000,N_5099,N_5747);
and U6001 (N_6001,N_5948,N_5861);
or U6002 (N_6002,N_5674,N_5720);
nand U6003 (N_6003,N_5909,N_5539);
nand U6004 (N_6004,N_5911,N_5477);
xnor U6005 (N_6005,N_5405,N_5855);
nor U6006 (N_6006,N_5061,N_5520);
xor U6007 (N_6007,N_5191,N_5093);
nand U6008 (N_6008,N_5599,N_5961);
xor U6009 (N_6009,N_5046,N_5661);
nand U6010 (N_6010,N_5514,N_5915);
and U6011 (N_6011,N_5100,N_5389);
nand U6012 (N_6012,N_5551,N_5614);
or U6013 (N_6013,N_5459,N_5872);
xnor U6014 (N_6014,N_5194,N_5347);
nand U6015 (N_6015,N_5225,N_5836);
nor U6016 (N_6016,N_5509,N_5688);
or U6017 (N_6017,N_5937,N_5779);
nand U6018 (N_6018,N_5935,N_5698);
nor U6019 (N_6019,N_5247,N_5657);
nor U6020 (N_6020,N_5110,N_5232);
nand U6021 (N_6021,N_5679,N_5017);
and U6022 (N_6022,N_5324,N_5150);
nand U6023 (N_6023,N_5702,N_5335);
xor U6024 (N_6024,N_5580,N_5781);
xor U6025 (N_6025,N_5873,N_5859);
or U6026 (N_6026,N_5486,N_5808);
nand U6027 (N_6027,N_5211,N_5549);
nor U6028 (N_6028,N_5140,N_5226);
or U6029 (N_6029,N_5920,N_5256);
nor U6030 (N_6030,N_5812,N_5913);
xnor U6031 (N_6031,N_5999,N_5399);
nor U6032 (N_6032,N_5758,N_5972);
nor U6033 (N_6033,N_5036,N_5690);
nand U6034 (N_6034,N_5381,N_5723);
and U6035 (N_6035,N_5178,N_5451);
xnor U6036 (N_6036,N_5768,N_5939);
or U6037 (N_6037,N_5914,N_5184);
xnor U6038 (N_6038,N_5671,N_5057);
nor U6039 (N_6039,N_5642,N_5414);
nor U6040 (N_6040,N_5689,N_5553);
nand U6041 (N_6041,N_5111,N_5994);
nor U6042 (N_6042,N_5884,N_5002);
nand U6043 (N_6043,N_5653,N_5052);
and U6044 (N_6044,N_5415,N_5432);
and U6045 (N_6045,N_5359,N_5395);
xnor U6046 (N_6046,N_5265,N_5814);
and U6047 (N_6047,N_5740,N_5803);
or U6048 (N_6048,N_5439,N_5020);
nand U6049 (N_6049,N_5841,N_5524);
or U6050 (N_6050,N_5336,N_5673);
or U6051 (N_6051,N_5217,N_5101);
or U6052 (N_6052,N_5648,N_5953);
and U6053 (N_6053,N_5148,N_5259);
nor U6054 (N_6054,N_5638,N_5132);
and U6055 (N_6055,N_5511,N_5936);
or U6056 (N_6056,N_5607,N_5300);
nor U6057 (N_6057,N_5561,N_5367);
xnor U6058 (N_6058,N_5840,N_5233);
nand U6059 (N_6059,N_5312,N_5971);
and U6060 (N_6060,N_5856,N_5446);
nand U6061 (N_6061,N_5675,N_5450);
nand U6062 (N_6062,N_5786,N_5290);
and U6063 (N_6063,N_5379,N_5942);
nand U6064 (N_6064,N_5402,N_5600);
nor U6065 (N_6065,N_5230,N_5275);
and U6066 (N_6066,N_5572,N_5918);
nor U6067 (N_6067,N_5727,N_5717);
xor U6068 (N_6068,N_5502,N_5202);
and U6069 (N_6069,N_5408,N_5162);
or U6070 (N_6070,N_5000,N_5550);
and U6071 (N_6071,N_5737,N_5476);
nand U6072 (N_6072,N_5512,N_5606);
nand U6073 (N_6073,N_5033,N_5910);
and U6074 (N_6074,N_5388,N_5351);
or U6075 (N_6075,N_5806,N_5927);
xor U6076 (N_6076,N_5505,N_5004);
and U6077 (N_6077,N_5579,N_5445);
and U6078 (N_6078,N_5237,N_5097);
or U6079 (N_6079,N_5266,N_5308);
nor U6080 (N_6080,N_5537,N_5921);
nand U6081 (N_6081,N_5822,N_5789);
xor U6082 (N_6082,N_5147,N_5243);
nor U6083 (N_6083,N_5650,N_5294);
and U6084 (N_6084,N_5656,N_5299);
or U6085 (N_6085,N_5382,N_5339);
and U6086 (N_6086,N_5213,N_5930);
and U6087 (N_6087,N_5397,N_5531);
nand U6088 (N_6088,N_5115,N_5494);
nor U6089 (N_6089,N_5021,N_5493);
or U6090 (N_6090,N_5257,N_5070);
or U6091 (N_6091,N_5757,N_5102);
or U6092 (N_6092,N_5536,N_5680);
or U6093 (N_6093,N_5354,N_5499);
nor U6094 (N_6094,N_5584,N_5318);
or U6095 (N_6095,N_5570,N_5797);
or U6096 (N_6096,N_5203,N_5108);
and U6097 (N_6097,N_5124,N_5876);
nand U6098 (N_6098,N_5443,N_5331);
nand U6099 (N_6099,N_5252,N_5413);
nor U6100 (N_6100,N_5363,N_5007);
nor U6101 (N_6101,N_5933,N_5681);
nor U6102 (N_6102,N_5277,N_5463);
or U6103 (N_6103,N_5907,N_5134);
or U6104 (N_6104,N_5672,N_5605);
nor U6105 (N_6105,N_5869,N_5562);
xnor U6106 (N_6106,N_5498,N_5922);
xor U6107 (N_6107,N_5692,N_5372);
or U6108 (N_6108,N_5555,N_5842);
nor U6109 (N_6109,N_5902,N_5894);
nand U6110 (N_6110,N_5709,N_5712);
nor U6111 (N_6111,N_5079,N_5711);
nor U6112 (N_6112,N_5542,N_5938);
xnor U6113 (N_6113,N_5954,N_5436);
and U6114 (N_6114,N_5546,N_5851);
and U6115 (N_6115,N_5992,N_5391);
nor U6116 (N_6116,N_5510,N_5329);
xor U6117 (N_6117,N_5538,N_5297);
nor U6118 (N_6118,N_5323,N_5192);
and U6119 (N_6119,N_5287,N_5305);
and U6120 (N_6120,N_5077,N_5665);
nand U6121 (N_6121,N_5107,N_5283);
nand U6122 (N_6122,N_5713,N_5645);
or U6123 (N_6123,N_5949,N_5398);
and U6124 (N_6124,N_5258,N_5978);
nand U6125 (N_6125,N_5205,N_5094);
or U6126 (N_6126,N_5288,N_5343);
nand U6127 (N_6127,N_5249,N_5633);
xor U6128 (N_6128,N_5787,N_5635);
nor U6129 (N_6129,N_5261,N_5559);
xor U6130 (N_6130,N_5401,N_5044);
xor U6131 (N_6131,N_5892,N_5652);
xnor U6132 (N_6132,N_5874,N_5532);
nor U6133 (N_6133,N_5478,N_5885);
or U6134 (N_6134,N_5696,N_5990);
nor U6135 (N_6135,N_5955,N_5291);
xor U6136 (N_6136,N_5271,N_5304);
nor U6137 (N_6137,N_5188,N_5278);
nand U6138 (N_6138,N_5228,N_5736);
or U6139 (N_6139,N_5164,N_5734);
or U6140 (N_6140,N_5507,N_5500);
and U6141 (N_6141,N_5015,N_5270);
xor U6142 (N_6142,N_5001,N_5926);
nor U6143 (N_6143,N_5566,N_5867);
xor U6144 (N_6144,N_5752,N_5785);
nor U6145 (N_6145,N_5160,N_5461);
or U6146 (N_6146,N_5651,N_5835);
nand U6147 (N_6147,N_5362,N_5344);
nor U6148 (N_6148,N_5898,N_5545);
nor U6149 (N_6149,N_5594,N_5845);
nor U6150 (N_6150,N_5464,N_5325);
nand U6151 (N_6151,N_5619,N_5573);
or U6152 (N_6152,N_5313,N_5056);
or U6153 (N_6153,N_5706,N_5967);
and U6154 (N_6154,N_5172,N_5274);
nand U6155 (N_6155,N_5438,N_5714);
xnor U6156 (N_6156,N_5603,N_5832);
nand U6157 (N_6157,N_5602,N_5468);
nor U6158 (N_6158,N_5063,N_5941);
nor U6159 (N_6159,N_5014,N_5624);
and U6160 (N_6160,N_5460,N_5701);
nor U6161 (N_6161,N_5114,N_5149);
and U6162 (N_6162,N_5116,N_5010);
xor U6163 (N_6163,N_5593,N_5043);
or U6164 (N_6164,N_5189,N_5098);
and U6165 (N_6165,N_5534,N_5637);
nand U6166 (N_6166,N_5868,N_5142);
or U6167 (N_6167,N_5728,N_5170);
nand U6168 (N_6168,N_5667,N_5658);
or U6169 (N_6169,N_5360,N_5893);
or U6170 (N_6170,N_5073,N_5771);
xor U6171 (N_6171,N_5206,N_5660);
and U6172 (N_6172,N_5678,N_5458);
xor U6173 (N_6173,N_5337,N_5826);
and U6174 (N_6174,N_5361,N_5628);
nand U6175 (N_6175,N_5794,N_5253);
xnor U6176 (N_6176,N_5374,N_5197);
nand U6177 (N_6177,N_5846,N_5899);
xor U6178 (N_6178,N_5547,N_5370);
nor U6179 (N_6179,N_5557,N_5519);
nand U6180 (N_6180,N_5818,N_5407);
nor U6181 (N_6181,N_5770,N_5267);
xnor U6182 (N_6182,N_5783,N_5541);
and U6183 (N_6183,N_5490,N_5364);
nand U6184 (N_6184,N_5754,N_5819);
nor U6185 (N_6185,N_5923,N_5453);
nor U6186 (N_6186,N_5905,N_5138);
and U6187 (N_6187,N_5581,N_5244);
nor U6188 (N_6188,N_5383,N_5090);
xnor U6189 (N_6189,N_5946,N_5141);
and U6190 (N_6190,N_5743,N_5292);
and U6191 (N_6191,N_5222,N_5966);
or U6192 (N_6192,N_5465,N_5621);
nor U6193 (N_6193,N_5179,N_5106);
or U6194 (N_6194,N_5231,N_5066);
or U6195 (N_6195,N_5729,N_5227);
and U6196 (N_6196,N_5055,N_5957);
nand U6197 (N_6197,N_5617,N_5326);
xnor U6198 (N_6198,N_5322,N_5423);
nor U6199 (N_6199,N_5577,N_5289);
or U6200 (N_6200,N_5775,N_5040);
xor U6201 (N_6201,N_5136,N_5609);
or U6202 (N_6202,N_5622,N_5760);
and U6203 (N_6203,N_5129,N_5295);
and U6204 (N_6204,N_5366,N_5377);
xor U6205 (N_6205,N_5151,N_5041);
or U6206 (N_6206,N_5823,N_5442);
nand U6207 (N_6207,N_5240,N_5176);
and U6208 (N_6208,N_5615,N_5422);
and U6209 (N_6209,N_5683,N_5332);
xnor U6210 (N_6210,N_5521,N_5054);
nor U6211 (N_6211,N_5485,N_5597);
and U6212 (N_6212,N_5234,N_5175);
and U6213 (N_6213,N_5641,N_5153);
nand U6214 (N_6214,N_5092,N_5068);
xor U6215 (N_6215,N_5693,N_5083);
and U6216 (N_6216,N_5356,N_5034);
nor U6217 (N_6217,N_5601,N_5810);
or U6218 (N_6218,N_5582,N_5871);
or U6219 (N_6219,N_5437,N_5384);
and U6220 (N_6220,N_5302,N_5748);
or U6221 (N_6221,N_5492,N_5654);
nand U6222 (N_6222,N_5242,N_5908);
and U6223 (N_6223,N_5236,N_5973);
xnor U6224 (N_6224,N_5375,N_5462);
xor U6225 (N_6225,N_5281,N_5625);
nor U6226 (N_6226,N_5944,N_5260);
or U6227 (N_6227,N_5403,N_5865);
xnor U6228 (N_6228,N_5454,N_5119);
and U6229 (N_6229,N_5396,N_5032);
or U6230 (N_6230,N_5181,N_5746);
nor U6231 (N_6231,N_5345,N_5889);
xnor U6232 (N_6232,N_5997,N_5307);
or U6233 (N_6233,N_5982,N_5880);
and U6234 (N_6234,N_5440,N_5739);
xor U6235 (N_6235,N_5655,N_5756);
xor U6236 (N_6236,N_5251,N_5528);
and U6237 (N_6237,N_5365,N_5996);
and U6238 (N_6238,N_5755,N_5863);
or U6239 (N_6239,N_5145,N_5012);
or U6240 (N_6240,N_5103,N_5470);
nor U6241 (N_6241,N_5167,N_5799);
and U6242 (N_6242,N_5790,N_5328);
nand U6243 (N_6243,N_5137,N_5455);
nor U6244 (N_6244,N_5722,N_5029);
or U6245 (N_6245,N_5919,N_5829);
nand U6246 (N_6246,N_5612,N_5346);
nor U6247 (N_6247,N_5724,N_5050);
nand U6248 (N_6248,N_5903,N_5418);
nand U6249 (N_6249,N_5338,N_5086);
or U6250 (N_6250,N_5207,N_5424);
nand U6251 (N_6251,N_5084,N_5730);
nand U6252 (N_6252,N_5540,N_5820);
nor U6253 (N_6253,N_5031,N_5198);
or U6254 (N_6254,N_5262,N_5472);
nand U6255 (N_6255,N_5725,N_5122);
nand U6256 (N_6256,N_5870,N_5830);
or U6257 (N_6257,N_5616,N_5357);
or U6258 (N_6258,N_5471,N_5591);
nor U6259 (N_6259,N_5831,N_5852);
nor U6260 (N_6260,N_5199,N_5105);
nor U6261 (N_6261,N_5595,N_5159);
xnor U6262 (N_6262,N_5604,N_5989);
and U6263 (N_6263,N_5157,N_5699);
nand U6264 (N_6264,N_5135,N_5774);
or U6265 (N_6265,N_5028,N_5934);
nand U6266 (N_6266,N_5828,N_5089);
nor U6267 (N_6267,N_5890,N_5864);
nand U6268 (N_6268,N_5793,N_5535);
nand U6269 (N_6269,N_5548,N_5763);
nor U6270 (N_6270,N_5798,N_5895);
or U6271 (N_6271,N_5080,N_5986);
and U6272 (N_6272,N_5517,N_5805);
xor U6273 (N_6273,N_5759,N_5045);
nor U6274 (N_6274,N_5051,N_5904);
nand U6275 (N_6275,N_5522,N_5221);
or U6276 (N_6276,N_5005,N_5639);
nor U6277 (N_6277,N_5296,N_5879);
nand U6278 (N_6278,N_5587,N_5506);
nand U6279 (N_6279,N_5195,N_5596);
xnor U6280 (N_6280,N_5087,N_5686);
nor U6281 (N_6281,N_5881,N_5480);
nor U6282 (N_6282,N_5069,N_5386);
nand U6283 (N_6283,N_5024,N_5750);
nor U6284 (N_6284,N_5816,N_5428);
or U6285 (N_6285,N_5039,N_5104);
and U6286 (N_6286,N_5065,N_5960);
and U6287 (N_6287,N_5780,N_5109);
xor U6288 (N_6288,N_5769,N_5404);
nand U6289 (N_6289,N_5564,N_5761);
and U6290 (N_6290,N_5254,N_5825);
xor U6291 (N_6291,N_5710,N_5659);
and U6292 (N_6292,N_5647,N_5072);
nor U6293 (N_6293,N_5788,N_5877);
nor U6294 (N_6294,N_5215,N_5394);
and U6295 (N_6295,N_5117,N_5742);
xor U6296 (N_6296,N_5161,N_5618);
and U6297 (N_6297,N_5013,N_5764);
nor U6298 (N_6298,N_5554,N_5139);
or U6299 (N_6299,N_5177,N_5390);
and U6300 (N_6300,N_5127,N_5456);
nor U6301 (N_6301,N_5662,N_5449);
and U6302 (N_6302,N_5526,N_5316);
xnor U6303 (N_6303,N_5062,N_5860);
nor U6304 (N_6304,N_5035,N_5800);
or U6305 (N_6305,N_5269,N_5417);
nand U6306 (N_6306,N_5410,N_5058);
xnor U6307 (N_6307,N_5687,N_5563);
or U6308 (N_6308,N_5556,N_5976);
nor U6309 (N_6309,N_5782,N_5833);
or U6310 (N_6310,N_5518,N_5917);
nand U6311 (N_6311,N_5513,N_5112);
or U6312 (N_6312,N_5796,N_5025);
xnor U6313 (N_6313,N_5060,N_5285);
and U6314 (N_6314,N_5216,N_5427);
xnor U6315 (N_6315,N_5421,N_5441);
and U6316 (N_6316,N_5218,N_5169);
and U6317 (N_6317,N_5610,N_5118);
nand U6318 (N_6318,N_5631,N_5916);
nand U6319 (N_6319,N_5314,N_5590);
nand U6320 (N_6320,N_5821,N_5987);
and U6321 (N_6321,N_5053,N_5575);
nand U6322 (N_6322,N_5406,N_5968);
nand U6323 (N_6323,N_5945,N_5074);
and U6324 (N_6324,N_5355,N_5726);
nor U6325 (N_6325,N_5174,N_5484);
xnor U6326 (N_6326,N_5738,N_5668);
nand U6327 (N_6327,N_5896,N_5802);
nand U6328 (N_6328,N_5317,N_5886);
nand U6329 (N_6329,N_5773,N_5489);
xor U6330 (N_6330,N_5088,N_5574);
and U6331 (N_6331,N_5705,N_5282);
nand U6332 (N_6332,N_5980,N_5447);
nor U6333 (N_6333,N_5011,N_5611);
xor U6334 (N_6334,N_5026,N_5320);
nor U6335 (N_6335,N_5848,N_5984);
or U6336 (N_6336,N_5183,N_5928);
nor U6337 (N_6337,N_5995,N_5731);
or U6338 (N_6338,N_5670,N_5970);
nor U6339 (N_6339,N_5646,N_5223);
nand U6340 (N_6340,N_5200,N_5196);
and U6341 (N_6341,N_5838,N_5327);
nor U6342 (N_6342,N_5762,N_5027);
or U6343 (N_6343,N_5416,N_5208);
nor U6344 (N_6344,N_5804,N_5630);
xnor U6345 (N_6345,N_5636,N_5481);
or U6346 (N_6346,N_5900,N_5071);
nand U6347 (N_6347,N_5733,N_5634);
or U6348 (N_6348,N_5629,N_5981);
or U6349 (N_6349,N_5286,N_5947);
nor U6350 (N_6350,N_5201,N_5568);
xor U6351 (N_6351,N_5473,N_5883);
xor U6352 (N_6352,N_5047,N_5745);
nor U6353 (N_6353,N_5358,N_5588);
or U6354 (N_6354,N_5479,N_5085);
xor U6355 (N_6355,N_5315,N_5235);
xor U6356 (N_6356,N_5452,N_5697);
nor U6357 (N_6357,N_5224,N_5887);
nand U6358 (N_6358,N_5154,N_5158);
xor U6359 (N_6359,N_5279,N_5964);
nor U6360 (N_6360,N_5019,N_5369);
nand U6361 (N_6361,N_5801,N_5246);
nor U6362 (N_6362,N_5817,N_5969);
nor U6363 (N_6363,N_5951,N_5784);
or U6364 (N_6364,N_5932,N_5263);
and U6365 (N_6365,N_5735,N_5430);
nor U6366 (N_6366,N_5393,N_5273);
nand U6367 (N_6367,N_5583,N_5623);
nor U6368 (N_6368,N_5349,N_5700);
and U6369 (N_6369,N_5501,N_5979);
or U6370 (N_6370,N_5018,N_5125);
nor U6371 (N_6371,N_5685,N_5210);
or U6372 (N_6372,N_5993,N_5677);
nor U6373 (N_6373,N_5608,N_5857);
xnor U6374 (N_6374,N_5182,N_5854);
xor U6375 (N_6375,N_5212,N_5844);
nor U6376 (N_6376,N_5766,N_5839);
xnor U6377 (N_6377,N_5578,N_5156);
nor U6378 (N_6378,N_5626,N_5704);
or U6379 (N_6379,N_5525,N_5076);
nand U6380 (N_6380,N_5741,N_5301);
and U6381 (N_6381,N_5190,N_5715);
and U6382 (N_6382,N_5544,N_5988);
or U6383 (N_6383,N_5882,N_5264);
and U6384 (N_6384,N_5813,N_5592);
xnor U6385 (N_6385,N_5952,N_5380);
nor U6386 (N_6386,N_5448,N_5483);
nand U6387 (N_6387,N_5891,N_5250);
nor U6388 (N_6388,N_5425,N_5732);
nand U6389 (N_6389,N_5186,N_5962);
nand U6390 (N_6390,N_5306,N_5400);
nand U6391 (N_6391,N_5632,N_5589);
nor U6392 (N_6392,N_5530,N_5834);
nand U6393 (N_6393,N_5837,N_5508);
and U6394 (N_6394,N_5807,N_5385);
nand U6395 (N_6395,N_5009,N_5875);
xor U6396 (N_6396,N_5878,N_5310);
nor U6397 (N_6397,N_5049,N_5113);
nand U6398 (N_6398,N_5912,N_5411);
nor U6399 (N_6399,N_5245,N_5958);
nor U6400 (N_6400,N_5691,N_5791);
xor U6401 (N_6401,N_5173,N_5703);
and U6402 (N_6402,N_5977,N_5795);
nor U6403 (N_6403,N_5219,N_5241);
xor U6404 (N_6404,N_5168,N_5131);
nand U6405 (N_6405,N_5931,N_5866);
nand U6406 (N_6406,N_5558,N_5862);
nor U6407 (N_6407,N_5180,N_5187);
or U6408 (N_6408,N_5644,N_5482);
and U6409 (N_6409,N_5497,N_5515);
or U6410 (N_6410,N_5853,N_5321);
nand U6411 (N_6411,N_5037,N_5420);
xnor U6412 (N_6412,N_5682,N_5412);
xnor U6413 (N_6413,N_5695,N_5133);
and U6414 (N_6414,N_5123,N_5293);
nand U6415 (N_6415,N_5749,N_5214);
and U6416 (N_6416,N_5006,N_5716);
or U6417 (N_6417,N_5008,N_5815);
or U6418 (N_6418,N_5333,N_5824);
nor U6419 (N_6419,N_5620,N_5444);
nor U6420 (N_6420,N_5664,N_5897);
and U6421 (N_6421,N_5466,N_5409);
nand U6422 (N_6422,N_5434,N_5376);
xnor U6423 (N_6423,N_5827,N_5003);
nor U6424 (N_6424,N_5585,N_5503);
or U6425 (N_6425,N_5811,N_5567);
xor U6426 (N_6426,N_5248,N_5925);
or U6427 (N_6427,N_5901,N_5627);
xor U6428 (N_6428,N_5023,N_5598);
nand U6429 (N_6429,N_5858,N_5469);
nor U6430 (N_6430,N_5030,N_5718);
nor U6431 (N_6431,N_5560,N_5330);
nor U6432 (N_6432,N_5371,N_5983);
nor U6433 (N_6433,N_5956,N_5091);
nor U6434 (N_6434,N_5684,N_5341);
and U6435 (N_6435,N_5940,N_5950);
xor U6436 (N_6436,N_5613,N_5075);
nor U6437 (N_6437,N_5435,N_5719);
and U6438 (N_6438,N_5708,N_5965);
nor U6439 (N_6439,N_5943,N_5998);
and U6440 (N_6440,N_5569,N_5504);
or U6441 (N_6441,N_5533,N_5171);
or U6442 (N_6442,N_5185,N_5694);
xor U6443 (N_6443,N_5272,N_5906);
xor U6444 (N_6444,N_5963,N_5143);
nand U6445 (N_6445,N_5543,N_5527);
xnor U6446 (N_6446,N_5663,N_5204);
or U6447 (N_6447,N_5765,N_5120);
xnor U6448 (N_6448,N_5319,N_5340);
and U6449 (N_6449,N_5744,N_5342);
nand U6450 (N_6450,N_5419,N_5529);
nand U6451 (N_6451,N_5640,N_5268);
and U6452 (N_6452,N_5146,N_5843);
and U6453 (N_6453,N_5433,N_5643);
and U6454 (N_6454,N_5776,N_5166);
or U6455 (N_6455,N_5850,N_5516);
nor U6456 (N_6456,N_5847,N_5487);
or U6457 (N_6457,N_5128,N_5392);
or U6458 (N_6458,N_5474,N_5144);
nor U6459 (N_6459,N_5163,N_5707);
nand U6460 (N_6460,N_5467,N_5239);
or U6461 (N_6461,N_5121,N_5975);
and U6462 (N_6462,N_5586,N_5255);
nor U6463 (N_6463,N_5495,N_5067);
and U6464 (N_6464,N_5751,N_5849);
xnor U6465 (N_6465,N_5929,N_5078);
nand U6466 (N_6466,N_5311,N_5048);
nand U6467 (N_6467,N_5353,N_5016);
and U6468 (N_6468,N_5038,N_5238);
and U6469 (N_6469,N_5152,N_5373);
nand U6470 (N_6470,N_5042,N_5309);
or U6471 (N_6471,N_5491,N_5378);
or U6472 (N_6472,N_5022,N_5523);
nand U6473 (N_6473,N_5303,N_5126);
and U6474 (N_6474,N_5280,N_5334);
and U6475 (N_6475,N_5096,N_5777);
xnor U6476 (N_6476,N_5298,N_5778);
and U6477 (N_6477,N_5350,N_5426);
and U6478 (N_6478,N_5368,N_5387);
and U6479 (N_6479,N_5985,N_5155);
and U6480 (N_6480,N_5888,N_5082);
and U6481 (N_6481,N_5229,N_5721);
nor U6482 (N_6482,N_5475,N_5809);
xnor U6483 (N_6483,N_5095,N_5792);
xor U6484 (N_6484,N_5130,N_5220);
or U6485 (N_6485,N_5676,N_5193);
or U6486 (N_6486,N_5571,N_5496);
or U6487 (N_6487,N_5276,N_5209);
xnor U6488 (N_6488,N_5457,N_5666);
and U6489 (N_6489,N_5552,N_5959);
and U6490 (N_6490,N_5064,N_5767);
xnor U6491 (N_6491,N_5991,N_5565);
and U6492 (N_6492,N_5352,N_5576);
xnor U6493 (N_6493,N_5348,N_5924);
and U6494 (N_6494,N_5081,N_5974);
or U6495 (N_6495,N_5649,N_5488);
nand U6496 (N_6496,N_5669,N_5429);
nor U6497 (N_6497,N_5284,N_5431);
or U6498 (N_6498,N_5059,N_5753);
nor U6499 (N_6499,N_5772,N_5165);
nand U6500 (N_6500,N_5883,N_5716);
or U6501 (N_6501,N_5012,N_5359);
xnor U6502 (N_6502,N_5420,N_5497);
nand U6503 (N_6503,N_5176,N_5490);
xor U6504 (N_6504,N_5374,N_5405);
and U6505 (N_6505,N_5160,N_5308);
nand U6506 (N_6506,N_5367,N_5624);
xor U6507 (N_6507,N_5144,N_5425);
xnor U6508 (N_6508,N_5019,N_5166);
xor U6509 (N_6509,N_5854,N_5630);
nand U6510 (N_6510,N_5209,N_5625);
xor U6511 (N_6511,N_5426,N_5222);
nor U6512 (N_6512,N_5913,N_5233);
and U6513 (N_6513,N_5444,N_5608);
xor U6514 (N_6514,N_5212,N_5281);
nand U6515 (N_6515,N_5974,N_5197);
nor U6516 (N_6516,N_5409,N_5366);
or U6517 (N_6517,N_5818,N_5202);
xnor U6518 (N_6518,N_5541,N_5040);
nor U6519 (N_6519,N_5380,N_5911);
xnor U6520 (N_6520,N_5680,N_5829);
nand U6521 (N_6521,N_5398,N_5163);
nand U6522 (N_6522,N_5506,N_5061);
nand U6523 (N_6523,N_5722,N_5960);
xnor U6524 (N_6524,N_5803,N_5476);
nand U6525 (N_6525,N_5086,N_5870);
nor U6526 (N_6526,N_5310,N_5452);
and U6527 (N_6527,N_5917,N_5413);
and U6528 (N_6528,N_5982,N_5824);
xnor U6529 (N_6529,N_5109,N_5630);
and U6530 (N_6530,N_5064,N_5789);
or U6531 (N_6531,N_5597,N_5653);
and U6532 (N_6532,N_5876,N_5678);
or U6533 (N_6533,N_5778,N_5287);
nor U6534 (N_6534,N_5059,N_5161);
xor U6535 (N_6535,N_5438,N_5968);
xor U6536 (N_6536,N_5326,N_5346);
xor U6537 (N_6537,N_5688,N_5185);
nor U6538 (N_6538,N_5386,N_5299);
or U6539 (N_6539,N_5380,N_5754);
and U6540 (N_6540,N_5022,N_5728);
nand U6541 (N_6541,N_5273,N_5488);
xnor U6542 (N_6542,N_5463,N_5116);
xor U6543 (N_6543,N_5487,N_5491);
nor U6544 (N_6544,N_5386,N_5507);
or U6545 (N_6545,N_5823,N_5562);
and U6546 (N_6546,N_5410,N_5721);
or U6547 (N_6547,N_5358,N_5338);
and U6548 (N_6548,N_5153,N_5797);
and U6549 (N_6549,N_5542,N_5826);
nand U6550 (N_6550,N_5277,N_5477);
nor U6551 (N_6551,N_5819,N_5010);
xnor U6552 (N_6552,N_5518,N_5330);
nand U6553 (N_6553,N_5507,N_5346);
nand U6554 (N_6554,N_5789,N_5250);
or U6555 (N_6555,N_5192,N_5842);
nand U6556 (N_6556,N_5861,N_5405);
nor U6557 (N_6557,N_5161,N_5993);
nand U6558 (N_6558,N_5361,N_5870);
xor U6559 (N_6559,N_5904,N_5934);
xnor U6560 (N_6560,N_5144,N_5332);
nand U6561 (N_6561,N_5224,N_5604);
or U6562 (N_6562,N_5131,N_5065);
and U6563 (N_6563,N_5870,N_5619);
xnor U6564 (N_6564,N_5694,N_5600);
nor U6565 (N_6565,N_5664,N_5115);
or U6566 (N_6566,N_5252,N_5964);
nor U6567 (N_6567,N_5806,N_5549);
nand U6568 (N_6568,N_5451,N_5457);
xor U6569 (N_6569,N_5005,N_5559);
nand U6570 (N_6570,N_5141,N_5441);
and U6571 (N_6571,N_5822,N_5731);
nand U6572 (N_6572,N_5994,N_5404);
xor U6573 (N_6573,N_5123,N_5750);
nand U6574 (N_6574,N_5657,N_5522);
or U6575 (N_6575,N_5204,N_5018);
xor U6576 (N_6576,N_5480,N_5737);
nor U6577 (N_6577,N_5187,N_5511);
or U6578 (N_6578,N_5326,N_5106);
xor U6579 (N_6579,N_5187,N_5936);
and U6580 (N_6580,N_5187,N_5247);
or U6581 (N_6581,N_5467,N_5836);
nor U6582 (N_6582,N_5024,N_5582);
nand U6583 (N_6583,N_5524,N_5999);
or U6584 (N_6584,N_5353,N_5693);
and U6585 (N_6585,N_5378,N_5484);
xnor U6586 (N_6586,N_5474,N_5347);
xnor U6587 (N_6587,N_5553,N_5254);
or U6588 (N_6588,N_5012,N_5854);
nor U6589 (N_6589,N_5405,N_5484);
nor U6590 (N_6590,N_5688,N_5605);
and U6591 (N_6591,N_5667,N_5796);
and U6592 (N_6592,N_5851,N_5070);
and U6593 (N_6593,N_5062,N_5727);
nand U6594 (N_6594,N_5718,N_5886);
xnor U6595 (N_6595,N_5797,N_5541);
nand U6596 (N_6596,N_5239,N_5949);
nor U6597 (N_6597,N_5795,N_5190);
xnor U6598 (N_6598,N_5718,N_5717);
xor U6599 (N_6599,N_5667,N_5590);
and U6600 (N_6600,N_5942,N_5712);
nand U6601 (N_6601,N_5917,N_5530);
or U6602 (N_6602,N_5194,N_5772);
xor U6603 (N_6603,N_5827,N_5886);
nand U6604 (N_6604,N_5728,N_5603);
and U6605 (N_6605,N_5300,N_5157);
nand U6606 (N_6606,N_5843,N_5005);
xor U6607 (N_6607,N_5922,N_5555);
nand U6608 (N_6608,N_5267,N_5650);
or U6609 (N_6609,N_5072,N_5151);
nand U6610 (N_6610,N_5317,N_5209);
and U6611 (N_6611,N_5206,N_5880);
and U6612 (N_6612,N_5832,N_5794);
or U6613 (N_6613,N_5384,N_5260);
xnor U6614 (N_6614,N_5580,N_5376);
nor U6615 (N_6615,N_5533,N_5479);
or U6616 (N_6616,N_5367,N_5469);
and U6617 (N_6617,N_5034,N_5733);
xor U6618 (N_6618,N_5979,N_5880);
xnor U6619 (N_6619,N_5229,N_5946);
or U6620 (N_6620,N_5192,N_5698);
xor U6621 (N_6621,N_5491,N_5757);
or U6622 (N_6622,N_5574,N_5049);
and U6623 (N_6623,N_5226,N_5455);
or U6624 (N_6624,N_5123,N_5095);
and U6625 (N_6625,N_5763,N_5130);
or U6626 (N_6626,N_5486,N_5359);
nor U6627 (N_6627,N_5994,N_5568);
nand U6628 (N_6628,N_5709,N_5338);
or U6629 (N_6629,N_5414,N_5431);
or U6630 (N_6630,N_5833,N_5788);
nor U6631 (N_6631,N_5136,N_5059);
and U6632 (N_6632,N_5032,N_5149);
nand U6633 (N_6633,N_5360,N_5402);
xnor U6634 (N_6634,N_5764,N_5406);
nand U6635 (N_6635,N_5080,N_5566);
nor U6636 (N_6636,N_5434,N_5757);
or U6637 (N_6637,N_5416,N_5481);
xor U6638 (N_6638,N_5834,N_5329);
or U6639 (N_6639,N_5402,N_5950);
or U6640 (N_6640,N_5132,N_5762);
nor U6641 (N_6641,N_5674,N_5276);
and U6642 (N_6642,N_5806,N_5672);
xor U6643 (N_6643,N_5619,N_5252);
and U6644 (N_6644,N_5108,N_5567);
nor U6645 (N_6645,N_5057,N_5792);
nand U6646 (N_6646,N_5693,N_5544);
nand U6647 (N_6647,N_5560,N_5773);
or U6648 (N_6648,N_5371,N_5630);
nand U6649 (N_6649,N_5976,N_5483);
and U6650 (N_6650,N_5008,N_5781);
xor U6651 (N_6651,N_5241,N_5200);
xnor U6652 (N_6652,N_5091,N_5004);
nand U6653 (N_6653,N_5664,N_5241);
and U6654 (N_6654,N_5281,N_5572);
or U6655 (N_6655,N_5993,N_5256);
or U6656 (N_6656,N_5181,N_5774);
nor U6657 (N_6657,N_5220,N_5999);
or U6658 (N_6658,N_5276,N_5905);
xor U6659 (N_6659,N_5663,N_5080);
nand U6660 (N_6660,N_5344,N_5779);
nor U6661 (N_6661,N_5971,N_5704);
xor U6662 (N_6662,N_5552,N_5780);
xor U6663 (N_6663,N_5070,N_5802);
nor U6664 (N_6664,N_5145,N_5520);
nor U6665 (N_6665,N_5981,N_5174);
and U6666 (N_6666,N_5595,N_5139);
or U6667 (N_6667,N_5188,N_5701);
nand U6668 (N_6668,N_5177,N_5887);
nand U6669 (N_6669,N_5725,N_5220);
nor U6670 (N_6670,N_5208,N_5350);
xnor U6671 (N_6671,N_5543,N_5459);
nor U6672 (N_6672,N_5179,N_5877);
nand U6673 (N_6673,N_5199,N_5148);
xor U6674 (N_6674,N_5949,N_5433);
xor U6675 (N_6675,N_5951,N_5738);
or U6676 (N_6676,N_5883,N_5210);
and U6677 (N_6677,N_5569,N_5443);
or U6678 (N_6678,N_5171,N_5062);
or U6679 (N_6679,N_5254,N_5692);
xor U6680 (N_6680,N_5672,N_5664);
xnor U6681 (N_6681,N_5565,N_5913);
nor U6682 (N_6682,N_5898,N_5049);
xor U6683 (N_6683,N_5633,N_5310);
or U6684 (N_6684,N_5486,N_5870);
nor U6685 (N_6685,N_5669,N_5125);
and U6686 (N_6686,N_5591,N_5470);
xnor U6687 (N_6687,N_5763,N_5570);
or U6688 (N_6688,N_5632,N_5601);
or U6689 (N_6689,N_5092,N_5832);
nor U6690 (N_6690,N_5635,N_5064);
nand U6691 (N_6691,N_5102,N_5972);
nor U6692 (N_6692,N_5684,N_5061);
or U6693 (N_6693,N_5414,N_5692);
or U6694 (N_6694,N_5251,N_5732);
or U6695 (N_6695,N_5866,N_5893);
or U6696 (N_6696,N_5393,N_5847);
nand U6697 (N_6697,N_5031,N_5056);
nand U6698 (N_6698,N_5952,N_5425);
and U6699 (N_6699,N_5387,N_5393);
xnor U6700 (N_6700,N_5193,N_5347);
nor U6701 (N_6701,N_5222,N_5534);
and U6702 (N_6702,N_5691,N_5552);
or U6703 (N_6703,N_5169,N_5769);
xnor U6704 (N_6704,N_5167,N_5656);
nand U6705 (N_6705,N_5035,N_5978);
xor U6706 (N_6706,N_5979,N_5874);
xor U6707 (N_6707,N_5185,N_5221);
or U6708 (N_6708,N_5751,N_5819);
nor U6709 (N_6709,N_5433,N_5321);
xor U6710 (N_6710,N_5113,N_5986);
nor U6711 (N_6711,N_5927,N_5374);
or U6712 (N_6712,N_5702,N_5556);
nor U6713 (N_6713,N_5463,N_5902);
nand U6714 (N_6714,N_5282,N_5672);
nand U6715 (N_6715,N_5014,N_5851);
nand U6716 (N_6716,N_5741,N_5454);
nor U6717 (N_6717,N_5971,N_5626);
nor U6718 (N_6718,N_5369,N_5245);
or U6719 (N_6719,N_5857,N_5890);
nor U6720 (N_6720,N_5480,N_5065);
nor U6721 (N_6721,N_5605,N_5390);
xor U6722 (N_6722,N_5237,N_5001);
nor U6723 (N_6723,N_5526,N_5774);
or U6724 (N_6724,N_5193,N_5487);
nand U6725 (N_6725,N_5590,N_5053);
and U6726 (N_6726,N_5158,N_5923);
nand U6727 (N_6727,N_5554,N_5416);
nand U6728 (N_6728,N_5225,N_5073);
and U6729 (N_6729,N_5623,N_5009);
nand U6730 (N_6730,N_5871,N_5760);
nand U6731 (N_6731,N_5456,N_5673);
or U6732 (N_6732,N_5592,N_5644);
or U6733 (N_6733,N_5796,N_5483);
nor U6734 (N_6734,N_5488,N_5431);
and U6735 (N_6735,N_5513,N_5766);
nand U6736 (N_6736,N_5147,N_5212);
and U6737 (N_6737,N_5458,N_5260);
and U6738 (N_6738,N_5050,N_5537);
xor U6739 (N_6739,N_5292,N_5481);
nand U6740 (N_6740,N_5162,N_5125);
or U6741 (N_6741,N_5508,N_5141);
nand U6742 (N_6742,N_5630,N_5168);
nand U6743 (N_6743,N_5004,N_5883);
or U6744 (N_6744,N_5807,N_5372);
nor U6745 (N_6745,N_5360,N_5299);
xor U6746 (N_6746,N_5786,N_5998);
xor U6747 (N_6747,N_5194,N_5912);
nor U6748 (N_6748,N_5781,N_5272);
nand U6749 (N_6749,N_5559,N_5807);
nand U6750 (N_6750,N_5608,N_5698);
xor U6751 (N_6751,N_5880,N_5942);
nor U6752 (N_6752,N_5150,N_5741);
and U6753 (N_6753,N_5771,N_5301);
and U6754 (N_6754,N_5896,N_5389);
or U6755 (N_6755,N_5221,N_5848);
xnor U6756 (N_6756,N_5772,N_5763);
and U6757 (N_6757,N_5170,N_5979);
xor U6758 (N_6758,N_5361,N_5491);
nand U6759 (N_6759,N_5521,N_5490);
nand U6760 (N_6760,N_5905,N_5706);
xor U6761 (N_6761,N_5966,N_5971);
and U6762 (N_6762,N_5645,N_5953);
nand U6763 (N_6763,N_5698,N_5762);
and U6764 (N_6764,N_5729,N_5713);
nor U6765 (N_6765,N_5550,N_5935);
nor U6766 (N_6766,N_5745,N_5905);
or U6767 (N_6767,N_5865,N_5982);
nand U6768 (N_6768,N_5413,N_5650);
nor U6769 (N_6769,N_5436,N_5050);
or U6770 (N_6770,N_5121,N_5081);
nor U6771 (N_6771,N_5942,N_5008);
xnor U6772 (N_6772,N_5057,N_5370);
or U6773 (N_6773,N_5267,N_5477);
nand U6774 (N_6774,N_5107,N_5733);
or U6775 (N_6775,N_5486,N_5007);
and U6776 (N_6776,N_5681,N_5903);
nor U6777 (N_6777,N_5092,N_5216);
nor U6778 (N_6778,N_5672,N_5044);
nand U6779 (N_6779,N_5331,N_5913);
xor U6780 (N_6780,N_5892,N_5124);
and U6781 (N_6781,N_5399,N_5818);
and U6782 (N_6782,N_5186,N_5212);
nor U6783 (N_6783,N_5469,N_5487);
nand U6784 (N_6784,N_5519,N_5479);
nand U6785 (N_6785,N_5385,N_5114);
nand U6786 (N_6786,N_5525,N_5016);
or U6787 (N_6787,N_5187,N_5033);
or U6788 (N_6788,N_5275,N_5376);
xor U6789 (N_6789,N_5774,N_5517);
xnor U6790 (N_6790,N_5685,N_5368);
and U6791 (N_6791,N_5740,N_5490);
xnor U6792 (N_6792,N_5750,N_5654);
or U6793 (N_6793,N_5711,N_5652);
or U6794 (N_6794,N_5977,N_5733);
or U6795 (N_6795,N_5009,N_5162);
nor U6796 (N_6796,N_5380,N_5167);
xnor U6797 (N_6797,N_5461,N_5843);
and U6798 (N_6798,N_5658,N_5801);
and U6799 (N_6799,N_5850,N_5707);
or U6800 (N_6800,N_5969,N_5928);
nor U6801 (N_6801,N_5552,N_5781);
xnor U6802 (N_6802,N_5095,N_5479);
nor U6803 (N_6803,N_5440,N_5334);
nor U6804 (N_6804,N_5582,N_5495);
or U6805 (N_6805,N_5426,N_5370);
xnor U6806 (N_6806,N_5422,N_5659);
and U6807 (N_6807,N_5547,N_5368);
or U6808 (N_6808,N_5919,N_5598);
xnor U6809 (N_6809,N_5078,N_5603);
nor U6810 (N_6810,N_5449,N_5633);
nand U6811 (N_6811,N_5944,N_5953);
and U6812 (N_6812,N_5600,N_5579);
nand U6813 (N_6813,N_5977,N_5394);
or U6814 (N_6814,N_5905,N_5902);
nor U6815 (N_6815,N_5468,N_5699);
or U6816 (N_6816,N_5010,N_5199);
or U6817 (N_6817,N_5602,N_5731);
or U6818 (N_6818,N_5986,N_5475);
nand U6819 (N_6819,N_5807,N_5156);
and U6820 (N_6820,N_5150,N_5696);
xnor U6821 (N_6821,N_5005,N_5863);
nor U6822 (N_6822,N_5798,N_5552);
nor U6823 (N_6823,N_5768,N_5147);
or U6824 (N_6824,N_5584,N_5461);
and U6825 (N_6825,N_5655,N_5895);
nand U6826 (N_6826,N_5601,N_5458);
or U6827 (N_6827,N_5207,N_5485);
nand U6828 (N_6828,N_5749,N_5628);
nand U6829 (N_6829,N_5773,N_5051);
and U6830 (N_6830,N_5472,N_5445);
nand U6831 (N_6831,N_5317,N_5982);
and U6832 (N_6832,N_5667,N_5073);
nand U6833 (N_6833,N_5703,N_5239);
nor U6834 (N_6834,N_5411,N_5102);
nor U6835 (N_6835,N_5889,N_5222);
and U6836 (N_6836,N_5228,N_5254);
nand U6837 (N_6837,N_5218,N_5312);
nor U6838 (N_6838,N_5254,N_5881);
nor U6839 (N_6839,N_5029,N_5217);
and U6840 (N_6840,N_5543,N_5000);
or U6841 (N_6841,N_5169,N_5946);
or U6842 (N_6842,N_5515,N_5852);
and U6843 (N_6843,N_5367,N_5107);
nand U6844 (N_6844,N_5839,N_5589);
xnor U6845 (N_6845,N_5610,N_5916);
and U6846 (N_6846,N_5643,N_5463);
and U6847 (N_6847,N_5373,N_5141);
or U6848 (N_6848,N_5720,N_5560);
nor U6849 (N_6849,N_5743,N_5465);
and U6850 (N_6850,N_5210,N_5920);
nor U6851 (N_6851,N_5968,N_5795);
nor U6852 (N_6852,N_5530,N_5414);
nand U6853 (N_6853,N_5506,N_5807);
or U6854 (N_6854,N_5685,N_5743);
nand U6855 (N_6855,N_5362,N_5697);
and U6856 (N_6856,N_5886,N_5426);
nor U6857 (N_6857,N_5587,N_5480);
or U6858 (N_6858,N_5607,N_5966);
xnor U6859 (N_6859,N_5688,N_5774);
nand U6860 (N_6860,N_5353,N_5600);
and U6861 (N_6861,N_5455,N_5240);
and U6862 (N_6862,N_5416,N_5392);
nand U6863 (N_6863,N_5890,N_5412);
or U6864 (N_6864,N_5251,N_5231);
and U6865 (N_6865,N_5029,N_5688);
xor U6866 (N_6866,N_5074,N_5920);
or U6867 (N_6867,N_5220,N_5427);
nand U6868 (N_6868,N_5101,N_5221);
or U6869 (N_6869,N_5232,N_5280);
or U6870 (N_6870,N_5898,N_5098);
nand U6871 (N_6871,N_5450,N_5987);
nor U6872 (N_6872,N_5019,N_5537);
and U6873 (N_6873,N_5996,N_5841);
and U6874 (N_6874,N_5819,N_5689);
xnor U6875 (N_6875,N_5009,N_5453);
xnor U6876 (N_6876,N_5199,N_5651);
nand U6877 (N_6877,N_5109,N_5374);
and U6878 (N_6878,N_5729,N_5839);
nand U6879 (N_6879,N_5140,N_5464);
or U6880 (N_6880,N_5922,N_5072);
nand U6881 (N_6881,N_5140,N_5485);
and U6882 (N_6882,N_5193,N_5430);
and U6883 (N_6883,N_5953,N_5327);
or U6884 (N_6884,N_5455,N_5747);
nand U6885 (N_6885,N_5491,N_5370);
and U6886 (N_6886,N_5553,N_5778);
or U6887 (N_6887,N_5657,N_5802);
and U6888 (N_6888,N_5468,N_5311);
nand U6889 (N_6889,N_5894,N_5162);
nand U6890 (N_6890,N_5556,N_5107);
xor U6891 (N_6891,N_5249,N_5462);
xor U6892 (N_6892,N_5933,N_5616);
nand U6893 (N_6893,N_5965,N_5819);
and U6894 (N_6894,N_5345,N_5065);
nand U6895 (N_6895,N_5093,N_5755);
nor U6896 (N_6896,N_5705,N_5608);
or U6897 (N_6897,N_5559,N_5995);
nand U6898 (N_6898,N_5646,N_5088);
or U6899 (N_6899,N_5427,N_5726);
xnor U6900 (N_6900,N_5169,N_5003);
and U6901 (N_6901,N_5394,N_5861);
and U6902 (N_6902,N_5865,N_5308);
and U6903 (N_6903,N_5123,N_5714);
nand U6904 (N_6904,N_5540,N_5842);
nor U6905 (N_6905,N_5551,N_5065);
nand U6906 (N_6906,N_5215,N_5284);
or U6907 (N_6907,N_5365,N_5308);
nor U6908 (N_6908,N_5537,N_5025);
nor U6909 (N_6909,N_5930,N_5450);
and U6910 (N_6910,N_5804,N_5088);
nor U6911 (N_6911,N_5627,N_5909);
nand U6912 (N_6912,N_5778,N_5244);
nand U6913 (N_6913,N_5740,N_5360);
xor U6914 (N_6914,N_5995,N_5323);
or U6915 (N_6915,N_5756,N_5905);
nor U6916 (N_6916,N_5589,N_5554);
and U6917 (N_6917,N_5028,N_5544);
or U6918 (N_6918,N_5763,N_5363);
nor U6919 (N_6919,N_5148,N_5078);
xnor U6920 (N_6920,N_5604,N_5736);
xnor U6921 (N_6921,N_5461,N_5497);
xnor U6922 (N_6922,N_5120,N_5695);
and U6923 (N_6923,N_5962,N_5105);
or U6924 (N_6924,N_5846,N_5212);
nand U6925 (N_6925,N_5762,N_5455);
xor U6926 (N_6926,N_5833,N_5736);
or U6927 (N_6927,N_5613,N_5784);
nor U6928 (N_6928,N_5912,N_5904);
xnor U6929 (N_6929,N_5639,N_5741);
and U6930 (N_6930,N_5990,N_5043);
nor U6931 (N_6931,N_5183,N_5110);
xor U6932 (N_6932,N_5823,N_5738);
nor U6933 (N_6933,N_5317,N_5710);
nor U6934 (N_6934,N_5385,N_5051);
and U6935 (N_6935,N_5747,N_5487);
and U6936 (N_6936,N_5872,N_5116);
nor U6937 (N_6937,N_5260,N_5585);
nand U6938 (N_6938,N_5191,N_5673);
or U6939 (N_6939,N_5247,N_5351);
and U6940 (N_6940,N_5782,N_5203);
or U6941 (N_6941,N_5791,N_5899);
or U6942 (N_6942,N_5980,N_5730);
and U6943 (N_6943,N_5050,N_5539);
nor U6944 (N_6944,N_5334,N_5650);
or U6945 (N_6945,N_5379,N_5418);
nor U6946 (N_6946,N_5888,N_5288);
xnor U6947 (N_6947,N_5421,N_5355);
nand U6948 (N_6948,N_5349,N_5049);
or U6949 (N_6949,N_5407,N_5410);
and U6950 (N_6950,N_5446,N_5164);
nand U6951 (N_6951,N_5985,N_5251);
xor U6952 (N_6952,N_5219,N_5611);
nor U6953 (N_6953,N_5567,N_5354);
or U6954 (N_6954,N_5669,N_5747);
or U6955 (N_6955,N_5921,N_5941);
nor U6956 (N_6956,N_5405,N_5698);
nor U6957 (N_6957,N_5753,N_5253);
and U6958 (N_6958,N_5861,N_5373);
nor U6959 (N_6959,N_5989,N_5180);
or U6960 (N_6960,N_5759,N_5329);
or U6961 (N_6961,N_5979,N_5023);
nor U6962 (N_6962,N_5546,N_5084);
nand U6963 (N_6963,N_5075,N_5962);
or U6964 (N_6964,N_5958,N_5079);
xnor U6965 (N_6965,N_5051,N_5403);
nand U6966 (N_6966,N_5916,N_5001);
or U6967 (N_6967,N_5955,N_5109);
xor U6968 (N_6968,N_5474,N_5499);
xnor U6969 (N_6969,N_5989,N_5537);
nand U6970 (N_6970,N_5442,N_5615);
or U6971 (N_6971,N_5594,N_5104);
and U6972 (N_6972,N_5755,N_5099);
xnor U6973 (N_6973,N_5694,N_5276);
and U6974 (N_6974,N_5186,N_5514);
nand U6975 (N_6975,N_5943,N_5655);
nand U6976 (N_6976,N_5436,N_5406);
and U6977 (N_6977,N_5923,N_5525);
and U6978 (N_6978,N_5717,N_5937);
or U6979 (N_6979,N_5605,N_5293);
or U6980 (N_6980,N_5524,N_5180);
xor U6981 (N_6981,N_5908,N_5560);
nor U6982 (N_6982,N_5287,N_5534);
nor U6983 (N_6983,N_5829,N_5817);
nand U6984 (N_6984,N_5726,N_5841);
or U6985 (N_6985,N_5483,N_5744);
nand U6986 (N_6986,N_5924,N_5045);
or U6987 (N_6987,N_5837,N_5996);
nor U6988 (N_6988,N_5244,N_5641);
xor U6989 (N_6989,N_5185,N_5430);
nor U6990 (N_6990,N_5327,N_5574);
nor U6991 (N_6991,N_5336,N_5956);
xnor U6992 (N_6992,N_5561,N_5166);
nor U6993 (N_6993,N_5654,N_5883);
and U6994 (N_6994,N_5169,N_5420);
xnor U6995 (N_6995,N_5559,N_5257);
nor U6996 (N_6996,N_5824,N_5680);
or U6997 (N_6997,N_5915,N_5459);
xor U6998 (N_6998,N_5971,N_5068);
and U6999 (N_6999,N_5407,N_5483);
xnor U7000 (N_7000,N_6261,N_6459);
nand U7001 (N_7001,N_6381,N_6766);
xnor U7002 (N_7002,N_6882,N_6278);
and U7003 (N_7003,N_6761,N_6888);
xor U7004 (N_7004,N_6854,N_6560);
nor U7005 (N_7005,N_6818,N_6338);
xnor U7006 (N_7006,N_6250,N_6443);
nand U7007 (N_7007,N_6603,N_6624);
nor U7008 (N_7008,N_6478,N_6101);
xnor U7009 (N_7009,N_6294,N_6680);
or U7010 (N_7010,N_6308,N_6215);
or U7011 (N_7011,N_6061,N_6553);
nor U7012 (N_7012,N_6040,N_6451);
or U7013 (N_7013,N_6442,N_6685);
and U7014 (N_7014,N_6024,N_6924);
nand U7015 (N_7015,N_6281,N_6028);
nor U7016 (N_7016,N_6765,N_6592);
nor U7017 (N_7017,N_6333,N_6594);
or U7018 (N_7018,N_6244,N_6686);
or U7019 (N_7019,N_6944,N_6626);
and U7020 (N_7020,N_6589,N_6260);
or U7021 (N_7021,N_6007,N_6668);
nor U7022 (N_7022,N_6386,N_6325);
nand U7023 (N_7023,N_6331,N_6519);
and U7024 (N_7024,N_6552,N_6688);
and U7025 (N_7025,N_6005,N_6873);
nand U7026 (N_7026,N_6817,N_6931);
or U7027 (N_7027,N_6890,N_6081);
nor U7028 (N_7028,N_6727,N_6164);
nand U7029 (N_7029,N_6191,N_6088);
nor U7030 (N_7030,N_6228,N_6365);
xor U7031 (N_7031,N_6324,N_6133);
or U7032 (N_7032,N_6900,N_6906);
nand U7033 (N_7033,N_6437,N_6558);
nor U7034 (N_7034,N_6729,N_6086);
or U7035 (N_7035,N_6463,N_6482);
and U7036 (N_7036,N_6207,N_6841);
and U7037 (N_7037,N_6779,N_6090);
xor U7038 (N_7038,N_6557,N_6837);
nand U7039 (N_7039,N_6726,N_6327);
and U7040 (N_7040,N_6960,N_6607);
nand U7041 (N_7041,N_6132,N_6982);
and U7042 (N_7042,N_6067,N_6747);
nor U7043 (N_7043,N_6857,N_6827);
nand U7044 (N_7044,N_6000,N_6606);
or U7045 (N_7045,N_6149,N_6919);
or U7046 (N_7046,N_6600,N_6499);
or U7047 (N_7047,N_6450,N_6613);
or U7048 (N_7048,N_6108,N_6427);
xor U7049 (N_7049,N_6990,N_6929);
and U7050 (N_7050,N_6051,N_6484);
nor U7051 (N_7051,N_6263,N_6513);
or U7052 (N_7052,N_6409,N_6050);
nand U7053 (N_7053,N_6676,N_6908);
xor U7054 (N_7054,N_6605,N_6312);
and U7055 (N_7055,N_6104,N_6710);
and U7056 (N_7056,N_6678,N_6912);
xor U7057 (N_7057,N_6737,N_6847);
xor U7058 (N_7058,N_6255,N_6355);
nor U7059 (N_7059,N_6099,N_6823);
and U7060 (N_7060,N_6885,N_6269);
xor U7061 (N_7061,N_6839,N_6423);
or U7062 (N_7062,N_6042,N_6136);
or U7063 (N_7063,N_6800,N_6881);
and U7064 (N_7064,N_6523,N_6148);
xor U7065 (N_7065,N_6073,N_6614);
or U7066 (N_7066,N_6543,N_6539);
nand U7067 (N_7067,N_6282,N_6198);
or U7068 (N_7068,N_6682,N_6230);
or U7069 (N_7069,N_6638,N_6271);
xor U7070 (N_7070,N_6524,N_6774);
xor U7071 (N_7071,N_6563,N_6011);
xnor U7072 (N_7072,N_6618,N_6397);
xnor U7073 (N_7073,N_6569,N_6803);
or U7074 (N_7074,N_6385,N_6240);
nand U7075 (N_7075,N_6852,N_6712);
nor U7076 (N_7076,N_6374,N_6573);
nand U7077 (N_7077,N_6856,N_6227);
nor U7078 (N_7078,N_6345,N_6498);
or U7079 (N_7079,N_6755,N_6163);
and U7080 (N_7080,N_6771,N_6453);
nor U7081 (N_7081,N_6257,N_6611);
and U7082 (N_7082,N_6320,N_6902);
or U7083 (N_7083,N_6899,N_6997);
and U7084 (N_7084,N_6448,N_6217);
or U7085 (N_7085,N_6256,N_6445);
or U7086 (N_7086,N_6077,N_6936);
xor U7087 (N_7087,N_6702,N_6113);
xor U7088 (N_7088,N_6930,N_6041);
and U7089 (N_7089,N_6705,N_6641);
nor U7090 (N_7090,N_6231,N_6928);
and U7091 (N_7091,N_6279,N_6330);
or U7092 (N_7092,N_6336,N_6435);
nand U7093 (N_7093,N_6440,N_6200);
nor U7094 (N_7094,N_6939,N_6938);
nor U7095 (N_7095,N_6877,N_6143);
and U7096 (N_7096,N_6984,N_6358);
xor U7097 (N_7097,N_6203,N_6674);
xnor U7098 (N_7098,N_6408,N_6768);
and U7099 (N_7099,N_6842,N_6627);
nor U7100 (N_7100,N_6623,N_6103);
xnor U7101 (N_7101,N_6152,N_6883);
xnor U7102 (N_7102,N_6068,N_6597);
xnor U7103 (N_7103,N_6154,N_6910);
or U7104 (N_7104,N_6047,N_6760);
nor U7105 (N_7105,N_6617,N_6106);
xor U7106 (N_7106,N_6695,N_6652);
nand U7107 (N_7107,N_6978,N_6654);
or U7108 (N_7108,N_6959,N_6075);
nand U7109 (N_7109,N_6773,N_6117);
and U7110 (N_7110,N_6575,N_6532);
or U7111 (N_7111,N_6535,N_6080);
or U7112 (N_7112,N_6981,N_6977);
or U7113 (N_7113,N_6403,N_6826);
xnor U7114 (N_7114,N_6446,N_6790);
nand U7115 (N_7115,N_6322,N_6033);
nand U7116 (N_7116,N_6147,N_6848);
or U7117 (N_7117,N_6961,N_6964);
and U7118 (N_7118,N_6340,N_6292);
nand U7119 (N_7119,N_6366,N_6302);
xor U7120 (N_7120,N_6684,N_6130);
nand U7121 (N_7121,N_6965,N_6807);
xor U7122 (N_7122,N_6515,N_6780);
xor U7123 (N_7123,N_6677,N_6027);
or U7124 (N_7124,N_6329,N_6886);
nand U7125 (N_7125,N_6180,N_6493);
xnor U7126 (N_7126,N_6082,N_6031);
nor U7127 (N_7127,N_6315,N_6376);
xor U7128 (N_7128,N_6884,N_6661);
and U7129 (N_7129,N_6742,N_6782);
nand U7130 (N_7130,N_6013,N_6943);
nand U7131 (N_7131,N_6540,N_6879);
xor U7132 (N_7132,N_6212,N_6811);
and U7133 (N_7133,N_6173,N_6290);
nor U7134 (N_7134,N_6194,N_6794);
nor U7135 (N_7135,N_6192,N_6361);
or U7136 (N_7136,N_6660,N_6916);
and U7137 (N_7137,N_6574,N_6467);
xor U7138 (N_7138,N_6470,N_6893);
xnor U7139 (N_7139,N_6021,N_6752);
nand U7140 (N_7140,N_6395,N_6022);
and U7141 (N_7141,N_6145,N_6599);
xnor U7142 (N_7142,N_6183,N_6349);
or U7143 (N_7143,N_6556,N_6764);
and U7144 (N_7144,N_6375,N_6236);
or U7145 (N_7145,N_6647,N_6527);
and U7146 (N_7146,N_6797,N_6009);
nand U7147 (N_7147,N_6283,N_6251);
or U7148 (N_7148,N_6016,N_6551);
nand U7149 (N_7149,N_6485,N_6970);
nor U7150 (N_7150,N_6867,N_6604);
xnor U7151 (N_7151,N_6500,N_6469);
xor U7152 (N_7152,N_6602,N_6105);
xnor U7153 (N_7153,N_6962,N_6023);
and U7154 (N_7154,N_6418,N_6190);
or U7155 (N_7155,N_6872,N_6341);
or U7156 (N_7156,N_6111,N_6400);
nand U7157 (N_7157,N_6026,N_6744);
and U7158 (N_7158,N_6037,N_6460);
nor U7159 (N_7159,N_6541,N_6998);
xnor U7160 (N_7160,N_6206,N_6757);
nand U7161 (N_7161,N_6436,N_6006);
nor U7162 (N_7162,N_6741,N_6896);
or U7163 (N_7163,N_6276,N_6428);
nand U7164 (N_7164,N_6795,N_6734);
and U7165 (N_7165,N_6656,N_6703);
xor U7166 (N_7166,N_6550,N_6792);
and U7167 (N_7167,N_6304,N_6243);
xor U7168 (N_7168,N_6536,N_6490);
nor U7169 (N_7169,N_6268,N_6628);
nand U7170 (N_7170,N_6559,N_6252);
xor U7171 (N_7171,N_6064,N_6922);
nor U7172 (N_7172,N_6706,N_6522);
xor U7173 (N_7173,N_6226,N_6415);
nand U7174 (N_7174,N_6321,N_6286);
and U7175 (N_7175,N_6237,N_6667);
or U7176 (N_7176,N_6275,N_6620);
or U7177 (N_7177,N_6564,N_6732);
or U7178 (N_7178,N_6870,N_6967);
or U7179 (N_7179,N_6004,N_6949);
nand U7180 (N_7180,N_6335,N_6404);
nand U7181 (N_7181,N_6505,N_6363);
xor U7182 (N_7182,N_6351,N_6270);
nand U7183 (N_7183,N_6093,N_6076);
xor U7184 (N_7184,N_6865,N_6581);
nor U7185 (N_7185,N_6071,N_6831);
xnor U7186 (N_7186,N_6772,N_6402);
xnor U7187 (N_7187,N_6239,N_6861);
xor U7188 (N_7188,N_6196,N_6158);
and U7189 (N_7189,N_6339,N_6974);
nand U7190 (N_7190,N_6935,N_6185);
xnor U7191 (N_7191,N_6489,N_6993);
nand U7192 (N_7192,N_6430,N_6254);
nor U7193 (N_7193,N_6208,N_6018);
or U7194 (N_7194,N_6666,N_6631);
and U7195 (N_7195,N_6801,N_6516);
and U7196 (N_7196,N_6472,N_6991);
nor U7197 (N_7197,N_6548,N_6019);
nor U7198 (N_7198,N_6700,N_6462);
and U7199 (N_7199,N_6120,N_6504);
or U7200 (N_7200,N_6380,N_6770);
nand U7201 (N_7201,N_6642,N_6114);
or U7202 (N_7202,N_6025,N_6074);
nand U7203 (N_7203,N_6131,N_6649);
nor U7204 (N_7204,N_6781,N_6512);
nand U7205 (N_7205,N_6287,N_6864);
and U7206 (N_7206,N_6394,N_6029);
and U7207 (N_7207,N_6305,N_6775);
and U7208 (N_7208,N_6123,N_6220);
and U7209 (N_7209,N_6937,N_6921);
and U7210 (N_7210,N_6739,N_6083);
nor U7211 (N_7211,N_6384,N_6788);
nor U7212 (N_7212,N_6014,N_6895);
and U7213 (N_7213,N_6079,N_6116);
and U7214 (N_7214,N_6311,N_6332);
or U7215 (N_7215,N_6644,N_6139);
nand U7216 (N_7216,N_6791,N_6671);
nand U7217 (N_7217,N_6946,N_6502);
and U7218 (N_7218,N_6348,N_6537);
and U7219 (N_7219,N_6566,N_6588);
xor U7220 (N_7220,N_6480,N_6357);
nor U7221 (N_7221,N_6822,N_6291);
nand U7222 (N_7222,N_6650,N_6951);
xnor U7223 (N_7223,N_6314,N_6187);
and U7224 (N_7224,N_6048,N_6653);
nor U7225 (N_7225,N_6479,N_6802);
xor U7226 (N_7226,N_6030,N_6683);
xnor U7227 (N_7227,N_6927,N_6957);
xnor U7228 (N_7228,N_6326,N_6989);
xnor U7229 (N_7229,N_6776,N_6941);
and U7230 (N_7230,N_6115,N_6932);
and U7231 (N_7231,N_6054,N_6232);
xor U7232 (N_7232,N_6669,N_6001);
xnor U7233 (N_7233,N_6576,N_6621);
or U7234 (N_7234,N_6298,N_6369);
nand U7235 (N_7235,N_6643,N_6751);
nand U7236 (N_7236,N_6595,N_6720);
or U7237 (N_7237,N_6417,N_6561);
xor U7238 (N_7238,N_6749,N_6307);
nor U7239 (N_7239,N_6619,N_6722);
or U7240 (N_7240,N_6640,N_6306);
or U7241 (N_7241,N_6663,N_6988);
nor U7242 (N_7242,N_6264,N_6309);
nand U7243 (N_7243,N_6630,N_6942);
xor U7244 (N_7244,N_6044,N_6495);
or U7245 (N_7245,N_6161,N_6034);
or U7246 (N_7246,N_6863,N_6904);
xor U7247 (N_7247,N_6247,N_6983);
xnor U7248 (N_7248,N_6659,N_6828);
xnor U7249 (N_7249,N_6065,N_6151);
or U7250 (N_7250,N_6477,N_6918);
nor U7251 (N_7251,N_6060,N_6850);
nor U7252 (N_7252,N_6214,N_6353);
or U7253 (N_7253,N_6182,N_6238);
or U7254 (N_7254,N_6692,N_6109);
nor U7255 (N_7255,N_6032,N_6150);
xnor U7256 (N_7256,N_6923,N_6137);
or U7257 (N_7257,N_6473,N_6517);
xor U7258 (N_7258,N_6999,N_6963);
or U7259 (N_7259,N_6288,N_6907);
xor U7260 (N_7260,N_6160,N_6610);
nand U7261 (N_7261,N_6429,N_6509);
xnor U7262 (N_7262,N_6945,N_6745);
or U7263 (N_7263,N_6176,N_6531);
nor U7264 (N_7264,N_6723,N_6750);
or U7265 (N_7265,N_6319,N_6112);
xor U7266 (N_7266,N_6748,N_6608);
nand U7267 (N_7267,N_6177,N_6213);
or U7268 (N_7268,N_6897,N_6249);
nor U7269 (N_7269,N_6169,N_6736);
or U7270 (N_7270,N_6815,N_6107);
nand U7271 (N_7271,N_6475,N_6438);
xor U7272 (N_7272,N_6805,N_6334);
and U7273 (N_7273,N_6809,N_6832);
nor U7274 (N_7274,N_6549,N_6052);
nand U7275 (N_7275,N_6796,N_6952);
nand U7276 (N_7276,N_6492,N_6259);
and U7277 (N_7277,N_6586,N_6843);
and U7278 (N_7278,N_6778,N_6078);
xnor U7279 (N_7279,N_6222,N_6426);
nand U7280 (N_7280,N_6799,N_6211);
xor U7281 (N_7281,N_6303,N_6830);
nand U7282 (N_7282,N_6425,N_6759);
or U7283 (N_7283,N_6398,N_6233);
nand U7284 (N_7284,N_6368,N_6789);
xor U7285 (N_7285,N_6582,N_6609);
nand U7286 (N_7286,N_6672,N_6954);
xnor U7287 (N_7287,N_6777,N_6804);
and U7288 (N_7288,N_6393,N_6063);
xnor U7289 (N_7289,N_6934,N_6691);
and U7290 (N_7290,N_6178,N_6645);
nand U7291 (N_7291,N_6346,N_6411);
or U7292 (N_7292,N_6915,N_6844);
nor U7293 (N_7293,N_6209,N_6992);
or U7294 (N_7294,N_6465,N_6849);
xnor U7295 (N_7295,N_6138,N_6171);
or U7296 (N_7296,N_6940,N_6547);
or U7297 (N_7297,N_6468,N_6474);
nand U7298 (N_7298,N_6892,N_6205);
nor U7299 (N_7299,N_6568,N_6825);
nand U7300 (N_7300,N_6784,N_6184);
or U7301 (N_7301,N_6267,N_6210);
and U7302 (N_7302,N_6901,N_6410);
nor U7303 (N_7303,N_6987,N_6891);
xnor U7304 (N_7304,N_6554,N_6874);
and U7305 (N_7305,N_6481,N_6265);
or U7306 (N_7306,N_6914,N_6382);
or U7307 (N_7307,N_6293,N_6199);
nor U7308 (N_7308,N_6506,N_6053);
xnor U7309 (N_7309,N_6420,N_6412);
or U7310 (N_7310,N_6360,N_6534);
nor U7311 (N_7311,N_6616,N_6170);
or U7312 (N_7312,N_6717,N_6679);
and U7313 (N_7313,N_6181,N_6097);
and U7314 (N_7314,N_6058,N_6711);
xor U7315 (N_7315,N_6371,N_6494);
or U7316 (N_7316,N_6740,N_6066);
or U7317 (N_7317,N_6503,N_6003);
or U7318 (N_7318,N_6461,N_6887);
and U7319 (N_7319,N_6359,N_6508);
and U7320 (N_7320,N_6567,N_6488);
nand U7321 (N_7321,N_6414,N_6769);
nand U7322 (N_7322,N_6284,N_6419);
or U7323 (N_7323,N_6625,N_6853);
and U7324 (N_7324,N_6793,N_6144);
nor U7325 (N_7325,N_6172,N_6570);
and U7326 (N_7326,N_6925,N_6675);
and U7327 (N_7327,N_6471,N_6578);
nor U7328 (N_7328,N_6447,N_6693);
nand U7329 (N_7329,N_6980,N_6615);
or U7330 (N_7330,N_6202,N_6094);
nand U7331 (N_7331,N_6846,N_6836);
xnor U7332 (N_7332,N_6175,N_6407);
or U7333 (N_7333,N_6008,N_6622);
nor U7334 (N_7334,N_6153,N_6225);
and U7335 (N_7335,N_6406,N_6687);
nand U7336 (N_7336,N_6898,N_6069);
and U7337 (N_7337,N_6584,N_6728);
nor U7338 (N_7338,N_6089,N_6452);
nand U7339 (N_7339,N_6601,N_6218);
xnor U7340 (N_7340,N_6421,N_6388);
xor U7341 (N_7341,N_6310,N_6708);
or U7342 (N_7342,N_6234,N_6973);
or U7343 (N_7343,N_6317,N_6986);
nor U7344 (N_7344,N_6223,N_6903);
nor U7345 (N_7345,N_6562,N_6819);
or U7346 (N_7346,N_6084,N_6933);
or U7347 (N_7347,N_6721,N_6894);
and U7348 (N_7348,N_6253,N_6070);
xor U7349 (N_7349,N_6313,N_6201);
nand U7350 (N_7350,N_6373,N_6344);
xor U7351 (N_7351,N_6483,N_6441);
xor U7352 (N_7352,N_6783,N_6690);
or U7353 (N_7353,N_6392,N_6119);
nand U7354 (N_7354,N_6612,N_6416);
or U7355 (N_7355,N_6920,N_6354);
or U7356 (N_7356,N_6100,N_6698);
nand U7357 (N_7357,N_6646,N_6162);
nand U7358 (N_7358,N_6141,N_6216);
xnor U7359 (N_7359,N_6718,N_6681);
or U7360 (N_7360,N_6289,N_6431);
and U7361 (N_7361,N_6510,N_6533);
xor U7362 (N_7362,N_6166,N_6458);
and U7363 (N_7363,N_6422,N_6958);
nor U7364 (N_7364,N_6528,N_6829);
or U7365 (N_7365,N_6731,N_6555);
nor U7366 (N_7366,N_6015,N_6753);
nor U7367 (N_7367,N_6456,N_6525);
or U7368 (N_7368,N_6806,N_6996);
nand U7369 (N_7369,N_6714,N_6277);
nand U7370 (N_7370,N_6128,N_6087);
nand U7371 (N_7371,N_6098,N_6219);
nor U7372 (N_7372,N_6636,N_6969);
and U7373 (N_7373,N_6501,N_6689);
xor U7374 (N_7374,N_6585,N_6948);
nand U7375 (N_7375,N_6091,N_6972);
and U7376 (N_7376,N_6529,N_6496);
or U7377 (N_7377,N_6057,N_6020);
and U7378 (N_7378,N_6860,N_6713);
xor U7379 (N_7379,N_6632,N_6658);
xnor U7380 (N_7380,N_6814,N_6035);
or U7381 (N_7381,N_6491,N_6186);
nor U7382 (N_7382,N_6657,N_6059);
or U7383 (N_7383,N_6204,N_6629);
or U7384 (N_7384,N_6486,N_6968);
xor U7385 (N_7385,N_6296,N_6167);
nor U7386 (N_7386,N_6285,N_6518);
or U7387 (N_7387,N_6762,N_6590);
or U7388 (N_7388,N_6125,N_6579);
or U7389 (N_7389,N_6118,N_6580);
nand U7390 (N_7390,N_6174,N_6242);
nand U7391 (N_7391,N_6110,N_6146);
nor U7392 (N_7392,N_6347,N_6538);
xor U7393 (N_7393,N_6372,N_6572);
and U7394 (N_7394,N_6545,N_6730);
xor U7395 (N_7395,N_6159,N_6639);
nand U7396 (N_7396,N_6917,N_6055);
nand U7397 (N_7397,N_6995,N_6966);
nand U7398 (N_7398,N_6295,N_6043);
or U7399 (N_7399,N_6197,N_6245);
nor U7400 (N_7400,N_6858,N_6845);
nor U7401 (N_7401,N_6168,N_6840);
nand U7402 (N_7402,N_6135,N_6155);
nor U7403 (N_7403,N_6913,N_6868);
and U7404 (N_7404,N_6707,N_6648);
and U7405 (N_7405,N_6716,N_6432);
and U7406 (N_7406,N_6140,N_6002);
and U7407 (N_7407,N_6763,N_6454);
nand U7408 (N_7408,N_6122,N_6129);
nand U7409 (N_7409,N_6274,N_6511);
nor U7410 (N_7410,N_6591,N_6039);
and U7411 (N_7411,N_6514,N_6821);
nor U7412 (N_7412,N_6318,N_6379);
and U7413 (N_7413,N_6362,N_6449);
and U7414 (N_7414,N_6655,N_6010);
or U7415 (N_7415,N_6994,N_6405);
and U7416 (N_7416,N_6062,N_6662);
xor U7417 (N_7417,N_6012,N_6634);
and U7418 (N_7418,N_6670,N_6221);
and U7419 (N_7419,N_6880,N_6049);
xor U7420 (N_7420,N_6577,N_6851);
nor U7421 (N_7421,N_6754,N_6719);
nor U7422 (N_7422,N_6387,N_6300);
and U7423 (N_7423,N_6072,N_6424);
nand U7424 (N_7424,N_6188,N_6724);
and U7425 (N_7425,N_6497,N_6808);
xnor U7426 (N_7426,N_6866,N_6950);
and U7427 (N_7427,N_6975,N_6869);
nor U7428 (N_7428,N_6598,N_6299);
nand U7429 (N_7429,N_6466,N_6633);
xnor U7430 (N_7430,N_6258,N_6673);
nand U7431 (N_7431,N_6521,N_6810);
nand U7432 (N_7432,N_6694,N_6127);
xnor U7433 (N_7433,N_6838,N_6095);
nand U7434 (N_7434,N_6979,N_6241);
nor U7435 (N_7435,N_6377,N_6816);
nor U7436 (N_7436,N_6142,N_6767);
nand U7437 (N_7437,N_6735,N_6248);
xnor U7438 (N_7438,N_6664,N_6985);
and U7439 (N_7439,N_6905,N_6725);
and U7440 (N_7440,N_6096,N_6911);
nand U7441 (N_7441,N_6544,N_6056);
nor U7442 (N_7442,N_6526,N_6704);
and U7443 (N_7443,N_6343,N_6571);
or U7444 (N_7444,N_6546,N_6102);
and U7445 (N_7445,N_6738,N_6875);
nand U7446 (N_7446,N_6017,N_6715);
nor U7447 (N_7447,N_6045,N_6947);
and U7448 (N_7448,N_6507,N_6812);
nand U7449 (N_7449,N_6195,N_6593);
nand U7450 (N_7450,N_6396,N_6487);
and U7451 (N_7451,N_6337,N_6476);
or U7452 (N_7452,N_6637,N_6383);
xor U7453 (N_7453,N_6701,N_6157);
nor U7454 (N_7454,N_6189,N_6297);
and U7455 (N_7455,N_6364,N_6651);
and U7456 (N_7456,N_6746,N_6798);
nand U7457 (N_7457,N_6280,N_6824);
nor U7458 (N_7458,N_6820,N_6266);
nand U7459 (N_7459,N_6956,N_6699);
nor U7460 (N_7460,N_6262,N_6587);
nand U7461 (N_7461,N_6124,N_6156);
and U7462 (N_7462,N_6036,N_6328);
nand U7463 (N_7463,N_6342,N_6976);
and U7464 (N_7464,N_6833,N_6378);
or U7465 (N_7465,N_6953,N_6835);
and U7466 (N_7466,N_6390,N_6444);
and U7467 (N_7467,N_6596,N_6758);
xor U7468 (N_7468,N_6389,N_6583);
or U7469 (N_7469,N_6391,N_6696);
xor U7470 (N_7470,N_6876,N_6224);
nand U7471 (N_7471,N_6370,N_6743);
or U7472 (N_7472,N_6179,N_6756);
nor U7473 (N_7473,N_6092,N_6229);
or U7474 (N_7474,N_6530,N_6520);
or U7475 (N_7475,N_6542,N_6786);
nand U7476 (N_7476,N_6457,N_6235);
or U7477 (N_7477,N_6787,N_6165);
xnor U7478 (N_7478,N_6871,N_6665);
or U7479 (N_7479,N_6434,N_6352);
nand U7480 (N_7480,N_6909,N_6926);
and U7481 (N_7481,N_6246,N_6038);
nor U7482 (N_7482,N_6323,N_6433);
nand U7483 (N_7483,N_6134,N_6439);
xnor U7484 (N_7484,N_6367,N_6272);
or U7485 (N_7485,N_6971,N_6878);
or U7486 (N_7486,N_6733,N_6813);
nand U7487 (N_7487,N_6859,N_6955);
and U7488 (N_7488,N_6085,N_6565);
nor U7489 (N_7489,N_6046,N_6785);
and U7490 (N_7490,N_6862,N_6121);
or U7491 (N_7491,N_6709,N_6413);
and U7492 (N_7492,N_6301,N_6316);
nor U7493 (N_7493,N_6273,N_6635);
nand U7494 (N_7494,N_6855,N_6193);
or U7495 (N_7495,N_6697,N_6401);
nand U7496 (N_7496,N_6889,N_6834);
nor U7497 (N_7497,N_6126,N_6356);
nor U7498 (N_7498,N_6350,N_6464);
nor U7499 (N_7499,N_6455,N_6399);
nor U7500 (N_7500,N_6613,N_6997);
and U7501 (N_7501,N_6935,N_6705);
nand U7502 (N_7502,N_6663,N_6939);
and U7503 (N_7503,N_6483,N_6566);
or U7504 (N_7504,N_6643,N_6517);
and U7505 (N_7505,N_6739,N_6172);
xor U7506 (N_7506,N_6168,N_6080);
nand U7507 (N_7507,N_6574,N_6932);
nand U7508 (N_7508,N_6251,N_6778);
and U7509 (N_7509,N_6138,N_6250);
nor U7510 (N_7510,N_6123,N_6293);
or U7511 (N_7511,N_6223,N_6472);
nor U7512 (N_7512,N_6997,N_6366);
nand U7513 (N_7513,N_6007,N_6427);
nand U7514 (N_7514,N_6694,N_6326);
nand U7515 (N_7515,N_6799,N_6950);
or U7516 (N_7516,N_6746,N_6908);
nor U7517 (N_7517,N_6516,N_6606);
xnor U7518 (N_7518,N_6236,N_6847);
nor U7519 (N_7519,N_6677,N_6933);
xor U7520 (N_7520,N_6143,N_6416);
or U7521 (N_7521,N_6293,N_6549);
and U7522 (N_7522,N_6699,N_6409);
xor U7523 (N_7523,N_6486,N_6440);
or U7524 (N_7524,N_6758,N_6396);
nand U7525 (N_7525,N_6713,N_6826);
nor U7526 (N_7526,N_6293,N_6722);
or U7527 (N_7527,N_6046,N_6313);
or U7528 (N_7528,N_6134,N_6536);
xnor U7529 (N_7529,N_6750,N_6053);
or U7530 (N_7530,N_6122,N_6921);
nand U7531 (N_7531,N_6554,N_6795);
and U7532 (N_7532,N_6834,N_6421);
nand U7533 (N_7533,N_6625,N_6903);
xor U7534 (N_7534,N_6255,N_6862);
xnor U7535 (N_7535,N_6064,N_6026);
or U7536 (N_7536,N_6317,N_6638);
nor U7537 (N_7537,N_6394,N_6911);
and U7538 (N_7538,N_6170,N_6012);
or U7539 (N_7539,N_6574,N_6491);
xor U7540 (N_7540,N_6536,N_6042);
or U7541 (N_7541,N_6305,N_6270);
nor U7542 (N_7542,N_6738,N_6029);
xor U7543 (N_7543,N_6118,N_6246);
or U7544 (N_7544,N_6844,N_6913);
xnor U7545 (N_7545,N_6245,N_6584);
and U7546 (N_7546,N_6606,N_6858);
and U7547 (N_7547,N_6299,N_6343);
nor U7548 (N_7548,N_6670,N_6902);
nor U7549 (N_7549,N_6799,N_6149);
nor U7550 (N_7550,N_6689,N_6323);
nor U7551 (N_7551,N_6162,N_6722);
and U7552 (N_7552,N_6774,N_6656);
nand U7553 (N_7553,N_6874,N_6383);
and U7554 (N_7554,N_6695,N_6600);
and U7555 (N_7555,N_6003,N_6581);
and U7556 (N_7556,N_6730,N_6993);
xor U7557 (N_7557,N_6813,N_6462);
or U7558 (N_7558,N_6686,N_6320);
nor U7559 (N_7559,N_6238,N_6901);
nand U7560 (N_7560,N_6735,N_6677);
nor U7561 (N_7561,N_6415,N_6202);
or U7562 (N_7562,N_6197,N_6687);
nand U7563 (N_7563,N_6830,N_6812);
or U7564 (N_7564,N_6344,N_6721);
xnor U7565 (N_7565,N_6118,N_6805);
nand U7566 (N_7566,N_6930,N_6488);
and U7567 (N_7567,N_6657,N_6441);
and U7568 (N_7568,N_6807,N_6505);
and U7569 (N_7569,N_6809,N_6046);
nor U7570 (N_7570,N_6760,N_6074);
nand U7571 (N_7571,N_6315,N_6246);
xor U7572 (N_7572,N_6846,N_6411);
nand U7573 (N_7573,N_6902,N_6199);
or U7574 (N_7574,N_6259,N_6415);
xor U7575 (N_7575,N_6963,N_6191);
and U7576 (N_7576,N_6656,N_6224);
xor U7577 (N_7577,N_6873,N_6558);
or U7578 (N_7578,N_6607,N_6720);
and U7579 (N_7579,N_6045,N_6831);
or U7580 (N_7580,N_6381,N_6609);
or U7581 (N_7581,N_6915,N_6726);
xnor U7582 (N_7582,N_6061,N_6433);
and U7583 (N_7583,N_6252,N_6137);
and U7584 (N_7584,N_6208,N_6232);
and U7585 (N_7585,N_6814,N_6286);
nand U7586 (N_7586,N_6627,N_6861);
nor U7587 (N_7587,N_6170,N_6566);
or U7588 (N_7588,N_6713,N_6805);
xnor U7589 (N_7589,N_6157,N_6782);
nor U7590 (N_7590,N_6394,N_6424);
nor U7591 (N_7591,N_6856,N_6155);
and U7592 (N_7592,N_6059,N_6643);
xnor U7593 (N_7593,N_6289,N_6120);
or U7594 (N_7594,N_6466,N_6182);
nand U7595 (N_7595,N_6586,N_6650);
and U7596 (N_7596,N_6855,N_6089);
xnor U7597 (N_7597,N_6326,N_6250);
or U7598 (N_7598,N_6839,N_6373);
and U7599 (N_7599,N_6796,N_6085);
and U7600 (N_7600,N_6146,N_6015);
or U7601 (N_7601,N_6725,N_6744);
and U7602 (N_7602,N_6145,N_6983);
and U7603 (N_7603,N_6906,N_6640);
or U7604 (N_7604,N_6218,N_6110);
xor U7605 (N_7605,N_6894,N_6945);
and U7606 (N_7606,N_6281,N_6070);
and U7607 (N_7607,N_6772,N_6801);
nand U7608 (N_7608,N_6265,N_6311);
or U7609 (N_7609,N_6013,N_6936);
nor U7610 (N_7610,N_6791,N_6587);
xnor U7611 (N_7611,N_6614,N_6371);
xnor U7612 (N_7612,N_6807,N_6708);
or U7613 (N_7613,N_6135,N_6262);
and U7614 (N_7614,N_6358,N_6273);
or U7615 (N_7615,N_6952,N_6917);
nor U7616 (N_7616,N_6482,N_6443);
and U7617 (N_7617,N_6570,N_6753);
or U7618 (N_7618,N_6411,N_6025);
or U7619 (N_7619,N_6670,N_6787);
xor U7620 (N_7620,N_6989,N_6799);
and U7621 (N_7621,N_6563,N_6762);
xor U7622 (N_7622,N_6981,N_6748);
xor U7623 (N_7623,N_6120,N_6130);
xor U7624 (N_7624,N_6769,N_6105);
and U7625 (N_7625,N_6948,N_6942);
and U7626 (N_7626,N_6489,N_6101);
xor U7627 (N_7627,N_6897,N_6386);
xnor U7628 (N_7628,N_6420,N_6164);
nor U7629 (N_7629,N_6024,N_6443);
nand U7630 (N_7630,N_6346,N_6094);
nand U7631 (N_7631,N_6585,N_6682);
or U7632 (N_7632,N_6760,N_6704);
xnor U7633 (N_7633,N_6074,N_6318);
xnor U7634 (N_7634,N_6894,N_6196);
nor U7635 (N_7635,N_6429,N_6169);
xnor U7636 (N_7636,N_6958,N_6537);
nor U7637 (N_7637,N_6042,N_6982);
nand U7638 (N_7638,N_6068,N_6836);
or U7639 (N_7639,N_6308,N_6266);
xnor U7640 (N_7640,N_6023,N_6828);
or U7641 (N_7641,N_6702,N_6974);
and U7642 (N_7642,N_6753,N_6055);
nor U7643 (N_7643,N_6265,N_6849);
nand U7644 (N_7644,N_6966,N_6016);
xnor U7645 (N_7645,N_6273,N_6718);
nor U7646 (N_7646,N_6834,N_6928);
xor U7647 (N_7647,N_6911,N_6689);
nor U7648 (N_7648,N_6945,N_6129);
or U7649 (N_7649,N_6593,N_6112);
nand U7650 (N_7650,N_6537,N_6647);
or U7651 (N_7651,N_6197,N_6951);
nor U7652 (N_7652,N_6252,N_6555);
nand U7653 (N_7653,N_6148,N_6490);
nor U7654 (N_7654,N_6466,N_6082);
nor U7655 (N_7655,N_6307,N_6054);
nor U7656 (N_7656,N_6702,N_6328);
and U7657 (N_7657,N_6454,N_6996);
and U7658 (N_7658,N_6522,N_6868);
and U7659 (N_7659,N_6738,N_6463);
xnor U7660 (N_7660,N_6553,N_6856);
nor U7661 (N_7661,N_6725,N_6563);
and U7662 (N_7662,N_6515,N_6572);
xnor U7663 (N_7663,N_6167,N_6505);
and U7664 (N_7664,N_6204,N_6155);
and U7665 (N_7665,N_6790,N_6252);
xor U7666 (N_7666,N_6087,N_6299);
or U7667 (N_7667,N_6844,N_6481);
nand U7668 (N_7668,N_6410,N_6116);
or U7669 (N_7669,N_6768,N_6516);
or U7670 (N_7670,N_6653,N_6031);
or U7671 (N_7671,N_6367,N_6118);
or U7672 (N_7672,N_6800,N_6605);
nand U7673 (N_7673,N_6198,N_6457);
and U7674 (N_7674,N_6718,N_6047);
or U7675 (N_7675,N_6035,N_6094);
nand U7676 (N_7676,N_6912,N_6675);
nand U7677 (N_7677,N_6215,N_6380);
nor U7678 (N_7678,N_6206,N_6192);
and U7679 (N_7679,N_6594,N_6936);
and U7680 (N_7680,N_6514,N_6186);
and U7681 (N_7681,N_6563,N_6057);
or U7682 (N_7682,N_6047,N_6107);
xnor U7683 (N_7683,N_6471,N_6504);
nand U7684 (N_7684,N_6992,N_6615);
and U7685 (N_7685,N_6217,N_6666);
nor U7686 (N_7686,N_6697,N_6369);
nand U7687 (N_7687,N_6866,N_6777);
xnor U7688 (N_7688,N_6964,N_6269);
xnor U7689 (N_7689,N_6104,N_6404);
or U7690 (N_7690,N_6100,N_6732);
nand U7691 (N_7691,N_6008,N_6062);
or U7692 (N_7692,N_6038,N_6753);
and U7693 (N_7693,N_6447,N_6465);
nor U7694 (N_7694,N_6503,N_6658);
nand U7695 (N_7695,N_6218,N_6891);
and U7696 (N_7696,N_6468,N_6418);
nor U7697 (N_7697,N_6298,N_6258);
or U7698 (N_7698,N_6022,N_6980);
xor U7699 (N_7699,N_6452,N_6379);
nor U7700 (N_7700,N_6302,N_6867);
xnor U7701 (N_7701,N_6420,N_6185);
nand U7702 (N_7702,N_6662,N_6258);
xnor U7703 (N_7703,N_6597,N_6400);
or U7704 (N_7704,N_6774,N_6344);
nand U7705 (N_7705,N_6035,N_6238);
nand U7706 (N_7706,N_6587,N_6334);
and U7707 (N_7707,N_6392,N_6715);
xnor U7708 (N_7708,N_6005,N_6046);
and U7709 (N_7709,N_6018,N_6038);
nor U7710 (N_7710,N_6531,N_6978);
xnor U7711 (N_7711,N_6476,N_6342);
xor U7712 (N_7712,N_6578,N_6747);
nand U7713 (N_7713,N_6900,N_6984);
nand U7714 (N_7714,N_6073,N_6411);
nor U7715 (N_7715,N_6140,N_6806);
or U7716 (N_7716,N_6987,N_6579);
and U7717 (N_7717,N_6193,N_6152);
nor U7718 (N_7718,N_6125,N_6334);
xor U7719 (N_7719,N_6396,N_6381);
or U7720 (N_7720,N_6554,N_6565);
and U7721 (N_7721,N_6261,N_6078);
or U7722 (N_7722,N_6720,N_6140);
xor U7723 (N_7723,N_6670,N_6236);
xnor U7724 (N_7724,N_6897,N_6065);
and U7725 (N_7725,N_6549,N_6466);
nor U7726 (N_7726,N_6634,N_6623);
and U7727 (N_7727,N_6105,N_6698);
or U7728 (N_7728,N_6846,N_6638);
nor U7729 (N_7729,N_6699,N_6358);
nand U7730 (N_7730,N_6369,N_6642);
nand U7731 (N_7731,N_6394,N_6579);
nand U7732 (N_7732,N_6838,N_6842);
nor U7733 (N_7733,N_6462,N_6374);
nor U7734 (N_7734,N_6674,N_6850);
nor U7735 (N_7735,N_6867,N_6128);
xnor U7736 (N_7736,N_6619,N_6458);
xnor U7737 (N_7737,N_6685,N_6573);
and U7738 (N_7738,N_6251,N_6103);
xor U7739 (N_7739,N_6559,N_6186);
nor U7740 (N_7740,N_6271,N_6260);
and U7741 (N_7741,N_6127,N_6628);
or U7742 (N_7742,N_6361,N_6889);
or U7743 (N_7743,N_6243,N_6141);
or U7744 (N_7744,N_6820,N_6965);
or U7745 (N_7745,N_6973,N_6661);
xor U7746 (N_7746,N_6980,N_6857);
xnor U7747 (N_7747,N_6303,N_6805);
or U7748 (N_7748,N_6226,N_6154);
nand U7749 (N_7749,N_6533,N_6158);
xor U7750 (N_7750,N_6313,N_6019);
nand U7751 (N_7751,N_6648,N_6810);
nor U7752 (N_7752,N_6996,N_6117);
nand U7753 (N_7753,N_6010,N_6865);
or U7754 (N_7754,N_6353,N_6063);
or U7755 (N_7755,N_6757,N_6197);
xnor U7756 (N_7756,N_6743,N_6336);
nor U7757 (N_7757,N_6364,N_6231);
or U7758 (N_7758,N_6298,N_6061);
xnor U7759 (N_7759,N_6338,N_6000);
and U7760 (N_7760,N_6724,N_6168);
nor U7761 (N_7761,N_6246,N_6702);
or U7762 (N_7762,N_6671,N_6940);
xnor U7763 (N_7763,N_6877,N_6278);
xor U7764 (N_7764,N_6117,N_6971);
and U7765 (N_7765,N_6599,N_6114);
and U7766 (N_7766,N_6756,N_6592);
or U7767 (N_7767,N_6862,N_6322);
nand U7768 (N_7768,N_6823,N_6702);
nand U7769 (N_7769,N_6493,N_6414);
xnor U7770 (N_7770,N_6168,N_6923);
nand U7771 (N_7771,N_6591,N_6393);
and U7772 (N_7772,N_6316,N_6433);
nor U7773 (N_7773,N_6028,N_6251);
nor U7774 (N_7774,N_6440,N_6805);
xnor U7775 (N_7775,N_6304,N_6735);
xnor U7776 (N_7776,N_6908,N_6483);
nor U7777 (N_7777,N_6397,N_6670);
and U7778 (N_7778,N_6849,N_6883);
nand U7779 (N_7779,N_6207,N_6256);
nand U7780 (N_7780,N_6702,N_6981);
nand U7781 (N_7781,N_6624,N_6403);
or U7782 (N_7782,N_6720,N_6003);
xnor U7783 (N_7783,N_6078,N_6354);
xnor U7784 (N_7784,N_6934,N_6810);
nand U7785 (N_7785,N_6407,N_6466);
and U7786 (N_7786,N_6675,N_6546);
nor U7787 (N_7787,N_6475,N_6666);
and U7788 (N_7788,N_6886,N_6264);
or U7789 (N_7789,N_6232,N_6216);
or U7790 (N_7790,N_6945,N_6342);
and U7791 (N_7791,N_6039,N_6164);
or U7792 (N_7792,N_6109,N_6925);
or U7793 (N_7793,N_6298,N_6262);
xor U7794 (N_7794,N_6894,N_6729);
nand U7795 (N_7795,N_6573,N_6199);
or U7796 (N_7796,N_6299,N_6206);
nor U7797 (N_7797,N_6307,N_6304);
nor U7798 (N_7798,N_6424,N_6406);
nor U7799 (N_7799,N_6903,N_6614);
nor U7800 (N_7800,N_6024,N_6167);
xor U7801 (N_7801,N_6929,N_6059);
nand U7802 (N_7802,N_6737,N_6751);
nand U7803 (N_7803,N_6033,N_6149);
or U7804 (N_7804,N_6949,N_6263);
xor U7805 (N_7805,N_6144,N_6556);
xnor U7806 (N_7806,N_6746,N_6923);
xnor U7807 (N_7807,N_6515,N_6517);
nand U7808 (N_7808,N_6600,N_6320);
xor U7809 (N_7809,N_6798,N_6954);
nor U7810 (N_7810,N_6956,N_6407);
xor U7811 (N_7811,N_6290,N_6595);
and U7812 (N_7812,N_6782,N_6298);
nor U7813 (N_7813,N_6084,N_6462);
and U7814 (N_7814,N_6734,N_6200);
and U7815 (N_7815,N_6992,N_6083);
nor U7816 (N_7816,N_6209,N_6902);
xnor U7817 (N_7817,N_6027,N_6271);
and U7818 (N_7818,N_6940,N_6794);
and U7819 (N_7819,N_6581,N_6784);
or U7820 (N_7820,N_6640,N_6972);
nor U7821 (N_7821,N_6788,N_6284);
nand U7822 (N_7822,N_6089,N_6615);
and U7823 (N_7823,N_6003,N_6699);
or U7824 (N_7824,N_6514,N_6673);
and U7825 (N_7825,N_6095,N_6064);
nand U7826 (N_7826,N_6504,N_6052);
or U7827 (N_7827,N_6907,N_6544);
and U7828 (N_7828,N_6065,N_6997);
nand U7829 (N_7829,N_6732,N_6802);
nand U7830 (N_7830,N_6718,N_6635);
or U7831 (N_7831,N_6616,N_6953);
or U7832 (N_7832,N_6788,N_6140);
or U7833 (N_7833,N_6153,N_6218);
nor U7834 (N_7834,N_6020,N_6881);
or U7835 (N_7835,N_6047,N_6900);
and U7836 (N_7836,N_6497,N_6042);
xor U7837 (N_7837,N_6743,N_6876);
nor U7838 (N_7838,N_6688,N_6261);
and U7839 (N_7839,N_6181,N_6561);
nor U7840 (N_7840,N_6457,N_6693);
nor U7841 (N_7841,N_6384,N_6174);
nor U7842 (N_7842,N_6182,N_6055);
nor U7843 (N_7843,N_6823,N_6891);
xnor U7844 (N_7844,N_6029,N_6485);
or U7845 (N_7845,N_6440,N_6393);
or U7846 (N_7846,N_6607,N_6285);
or U7847 (N_7847,N_6077,N_6810);
nand U7848 (N_7848,N_6805,N_6999);
nor U7849 (N_7849,N_6034,N_6116);
xor U7850 (N_7850,N_6487,N_6739);
nor U7851 (N_7851,N_6093,N_6184);
nor U7852 (N_7852,N_6274,N_6421);
nand U7853 (N_7853,N_6381,N_6282);
or U7854 (N_7854,N_6754,N_6548);
and U7855 (N_7855,N_6929,N_6343);
or U7856 (N_7856,N_6067,N_6641);
nor U7857 (N_7857,N_6796,N_6382);
xnor U7858 (N_7858,N_6337,N_6970);
or U7859 (N_7859,N_6094,N_6700);
or U7860 (N_7860,N_6839,N_6054);
nor U7861 (N_7861,N_6818,N_6053);
or U7862 (N_7862,N_6041,N_6920);
nand U7863 (N_7863,N_6860,N_6862);
xor U7864 (N_7864,N_6049,N_6384);
nand U7865 (N_7865,N_6817,N_6328);
and U7866 (N_7866,N_6154,N_6095);
nand U7867 (N_7867,N_6186,N_6303);
or U7868 (N_7868,N_6799,N_6905);
and U7869 (N_7869,N_6579,N_6262);
nor U7870 (N_7870,N_6708,N_6255);
nor U7871 (N_7871,N_6342,N_6706);
nor U7872 (N_7872,N_6018,N_6102);
nand U7873 (N_7873,N_6753,N_6676);
nand U7874 (N_7874,N_6761,N_6165);
or U7875 (N_7875,N_6648,N_6040);
nor U7876 (N_7876,N_6360,N_6578);
nand U7877 (N_7877,N_6677,N_6052);
and U7878 (N_7878,N_6573,N_6602);
xor U7879 (N_7879,N_6953,N_6587);
nand U7880 (N_7880,N_6516,N_6688);
and U7881 (N_7881,N_6841,N_6546);
xor U7882 (N_7882,N_6558,N_6858);
xnor U7883 (N_7883,N_6354,N_6627);
xnor U7884 (N_7884,N_6207,N_6213);
or U7885 (N_7885,N_6001,N_6741);
or U7886 (N_7886,N_6921,N_6539);
nor U7887 (N_7887,N_6274,N_6856);
and U7888 (N_7888,N_6751,N_6575);
and U7889 (N_7889,N_6479,N_6616);
nor U7890 (N_7890,N_6484,N_6751);
xor U7891 (N_7891,N_6316,N_6400);
nand U7892 (N_7892,N_6614,N_6958);
nand U7893 (N_7893,N_6143,N_6456);
nor U7894 (N_7894,N_6235,N_6983);
nand U7895 (N_7895,N_6110,N_6078);
and U7896 (N_7896,N_6971,N_6089);
and U7897 (N_7897,N_6496,N_6121);
nor U7898 (N_7898,N_6412,N_6846);
nand U7899 (N_7899,N_6088,N_6060);
nand U7900 (N_7900,N_6344,N_6521);
nand U7901 (N_7901,N_6267,N_6685);
xor U7902 (N_7902,N_6530,N_6909);
xor U7903 (N_7903,N_6219,N_6997);
or U7904 (N_7904,N_6596,N_6083);
xor U7905 (N_7905,N_6458,N_6091);
and U7906 (N_7906,N_6636,N_6033);
nand U7907 (N_7907,N_6408,N_6108);
nor U7908 (N_7908,N_6738,N_6511);
or U7909 (N_7909,N_6950,N_6808);
nand U7910 (N_7910,N_6380,N_6320);
and U7911 (N_7911,N_6494,N_6786);
and U7912 (N_7912,N_6349,N_6485);
nand U7913 (N_7913,N_6020,N_6673);
or U7914 (N_7914,N_6754,N_6214);
nor U7915 (N_7915,N_6584,N_6447);
xnor U7916 (N_7916,N_6698,N_6116);
nand U7917 (N_7917,N_6957,N_6967);
xnor U7918 (N_7918,N_6809,N_6922);
or U7919 (N_7919,N_6381,N_6070);
xor U7920 (N_7920,N_6431,N_6382);
xor U7921 (N_7921,N_6320,N_6068);
xor U7922 (N_7922,N_6294,N_6633);
and U7923 (N_7923,N_6264,N_6937);
or U7924 (N_7924,N_6044,N_6320);
xnor U7925 (N_7925,N_6305,N_6473);
nand U7926 (N_7926,N_6883,N_6953);
xor U7927 (N_7927,N_6783,N_6099);
or U7928 (N_7928,N_6828,N_6992);
nand U7929 (N_7929,N_6760,N_6859);
or U7930 (N_7930,N_6338,N_6628);
and U7931 (N_7931,N_6998,N_6655);
nand U7932 (N_7932,N_6051,N_6264);
and U7933 (N_7933,N_6582,N_6614);
and U7934 (N_7934,N_6610,N_6665);
or U7935 (N_7935,N_6384,N_6531);
and U7936 (N_7936,N_6118,N_6430);
and U7937 (N_7937,N_6789,N_6110);
nand U7938 (N_7938,N_6546,N_6913);
nor U7939 (N_7939,N_6755,N_6584);
nor U7940 (N_7940,N_6360,N_6190);
or U7941 (N_7941,N_6920,N_6256);
nor U7942 (N_7942,N_6872,N_6038);
nor U7943 (N_7943,N_6973,N_6808);
nor U7944 (N_7944,N_6331,N_6939);
or U7945 (N_7945,N_6831,N_6762);
nor U7946 (N_7946,N_6443,N_6891);
nor U7947 (N_7947,N_6829,N_6798);
nor U7948 (N_7948,N_6662,N_6399);
nor U7949 (N_7949,N_6533,N_6897);
nand U7950 (N_7950,N_6946,N_6555);
nand U7951 (N_7951,N_6132,N_6235);
and U7952 (N_7952,N_6136,N_6812);
nand U7953 (N_7953,N_6202,N_6463);
nor U7954 (N_7954,N_6460,N_6776);
nand U7955 (N_7955,N_6604,N_6655);
and U7956 (N_7956,N_6991,N_6834);
and U7957 (N_7957,N_6043,N_6838);
and U7958 (N_7958,N_6436,N_6338);
xor U7959 (N_7959,N_6792,N_6474);
or U7960 (N_7960,N_6524,N_6384);
nand U7961 (N_7961,N_6151,N_6387);
or U7962 (N_7962,N_6397,N_6839);
or U7963 (N_7963,N_6639,N_6442);
xor U7964 (N_7964,N_6624,N_6234);
or U7965 (N_7965,N_6284,N_6198);
and U7966 (N_7966,N_6138,N_6865);
nand U7967 (N_7967,N_6369,N_6601);
or U7968 (N_7968,N_6975,N_6665);
xnor U7969 (N_7969,N_6987,N_6532);
nor U7970 (N_7970,N_6712,N_6152);
and U7971 (N_7971,N_6500,N_6689);
xnor U7972 (N_7972,N_6116,N_6505);
nand U7973 (N_7973,N_6242,N_6233);
nor U7974 (N_7974,N_6131,N_6578);
or U7975 (N_7975,N_6096,N_6661);
and U7976 (N_7976,N_6303,N_6152);
xnor U7977 (N_7977,N_6475,N_6680);
xnor U7978 (N_7978,N_6085,N_6553);
nor U7979 (N_7979,N_6741,N_6473);
nand U7980 (N_7980,N_6876,N_6582);
and U7981 (N_7981,N_6234,N_6238);
or U7982 (N_7982,N_6464,N_6878);
nor U7983 (N_7983,N_6496,N_6823);
and U7984 (N_7984,N_6359,N_6410);
nor U7985 (N_7985,N_6736,N_6035);
nor U7986 (N_7986,N_6138,N_6121);
nor U7987 (N_7987,N_6793,N_6017);
and U7988 (N_7988,N_6914,N_6322);
nor U7989 (N_7989,N_6087,N_6770);
or U7990 (N_7990,N_6940,N_6490);
or U7991 (N_7991,N_6781,N_6988);
nor U7992 (N_7992,N_6119,N_6581);
nand U7993 (N_7993,N_6550,N_6419);
or U7994 (N_7994,N_6524,N_6051);
nor U7995 (N_7995,N_6442,N_6543);
or U7996 (N_7996,N_6777,N_6200);
xnor U7997 (N_7997,N_6949,N_6960);
or U7998 (N_7998,N_6368,N_6120);
or U7999 (N_7999,N_6983,N_6085);
xor U8000 (N_8000,N_7006,N_7882);
nand U8001 (N_8001,N_7237,N_7011);
nor U8002 (N_8002,N_7950,N_7132);
xor U8003 (N_8003,N_7574,N_7088);
or U8004 (N_8004,N_7009,N_7197);
xor U8005 (N_8005,N_7502,N_7525);
xnor U8006 (N_8006,N_7356,N_7640);
xnor U8007 (N_8007,N_7351,N_7572);
nor U8008 (N_8008,N_7083,N_7823);
and U8009 (N_8009,N_7493,N_7171);
nand U8010 (N_8010,N_7863,N_7535);
and U8011 (N_8011,N_7016,N_7759);
or U8012 (N_8012,N_7213,N_7783);
and U8013 (N_8013,N_7624,N_7837);
nor U8014 (N_8014,N_7076,N_7658);
nor U8015 (N_8015,N_7769,N_7753);
nor U8016 (N_8016,N_7177,N_7565);
xor U8017 (N_8017,N_7944,N_7548);
and U8018 (N_8018,N_7465,N_7097);
or U8019 (N_8019,N_7614,N_7650);
or U8020 (N_8020,N_7071,N_7516);
and U8021 (N_8021,N_7741,N_7233);
nor U8022 (N_8022,N_7072,N_7259);
nor U8023 (N_8023,N_7904,N_7090);
xor U8024 (N_8024,N_7252,N_7727);
nand U8025 (N_8025,N_7571,N_7915);
xor U8026 (N_8026,N_7219,N_7334);
or U8027 (N_8027,N_7651,N_7507);
nor U8028 (N_8028,N_7275,N_7964);
xor U8029 (N_8029,N_7587,N_7223);
nor U8030 (N_8030,N_7668,N_7919);
and U8031 (N_8031,N_7362,N_7924);
xor U8032 (N_8032,N_7940,N_7390);
or U8033 (N_8033,N_7411,N_7128);
nor U8034 (N_8034,N_7291,N_7894);
or U8035 (N_8035,N_7646,N_7506);
nand U8036 (N_8036,N_7500,N_7639);
and U8037 (N_8037,N_7157,N_7939);
xnor U8038 (N_8038,N_7768,N_7248);
and U8039 (N_8039,N_7671,N_7274);
xnor U8040 (N_8040,N_7361,N_7193);
nand U8041 (N_8041,N_7024,N_7210);
or U8042 (N_8042,N_7819,N_7613);
nand U8043 (N_8043,N_7874,N_7696);
xor U8044 (N_8044,N_7693,N_7773);
nand U8045 (N_8045,N_7730,N_7562);
nand U8046 (N_8046,N_7568,N_7710);
xnor U8047 (N_8047,N_7486,N_7691);
xnor U8048 (N_8048,N_7342,N_7972);
nand U8049 (N_8049,N_7776,N_7198);
and U8050 (N_8050,N_7902,N_7531);
nand U8051 (N_8051,N_7281,N_7401);
nand U8052 (N_8052,N_7364,N_7181);
and U8053 (N_8053,N_7133,N_7810);
xnor U8054 (N_8054,N_7293,N_7993);
xnor U8055 (N_8055,N_7517,N_7942);
nand U8056 (N_8056,N_7510,N_7109);
xor U8057 (N_8057,N_7876,N_7995);
and U8058 (N_8058,N_7630,N_7604);
nand U8059 (N_8059,N_7108,N_7688);
and U8060 (N_8060,N_7106,N_7699);
xnor U8061 (N_8061,N_7179,N_7384);
and U8062 (N_8062,N_7468,N_7854);
and U8063 (N_8063,N_7170,N_7448);
nor U8064 (N_8064,N_7138,N_7519);
nand U8065 (N_8065,N_7841,N_7946);
and U8066 (N_8066,N_7878,N_7005);
nor U8067 (N_8067,N_7709,N_7609);
nor U8068 (N_8068,N_7185,N_7247);
xor U8069 (N_8069,N_7827,N_7272);
xnor U8070 (N_8070,N_7323,N_7853);
or U8071 (N_8071,N_7402,N_7620);
or U8072 (N_8072,N_7897,N_7503);
nand U8073 (N_8073,N_7811,N_7117);
nand U8074 (N_8074,N_7920,N_7616);
nand U8075 (N_8075,N_7560,N_7752);
xnor U8076 (N_8076,N_7726,N_7798);
nor U8077 (N_8077,N_7637,N_7784);
nor U8078 (N_8078,N_7887,N_7733);
xnor U8079 (N_8079,N_7343,N_7721);
xnor U8080 (N_8080,N_7393,N_7154);
or U8081 (N_8081,N_7771,N_7834);
nand U8082 (N_8082,N_7822,N_7421);
nor U8083 (N_8083,N_7976,N_7400);
nor U8084 (N_8084,N_7675,N_7447);
xnor U8085 (N_8085,N_7102,N_7778);
or U8086 (N_8086,N_7360,N_7672);
nor U8087 (N_8087,N_7595,N_7387);
and U8088 (N_8088,N_7461,N_7349);
xor U8089 (N_8089,N_7842,N_7655);
or U8090 (N_8090,N_7278,N_7427);
or U8091 (N_8091,N_7756,N_7328);
nand U8092 (N_8092,N_7282,N_7222);
and U8093 (N_8093,N_7289,N_7934);
and U8094 (N_8094,N_7182,N_7977);
and U8095 (N_8095,N_7330,N_7473);
nor U8096 (N_8096,N_7445,N_7497);
nand U8097 (N_8097,N_7744,N_7828);
xor U8098 (N_8098,N_7591,N_7000);
and U8099 (N_8099,N_7514,N_7437);
and U8100 (N_8100,N_7286,N_7664);
or U8101 (N_8101,N_7186,N_7829);
nand U8102 (N_8102,N_7321,N_7116);
or U8103 (N_8103,N_7423,N_7340);
nand U8104 (N_8104,N_7312,N_7202);
xnor U8105 (N_8105,N_7736,N_7795);
or U8106 (N_8106,N_7835,N_7295);
nand U8107 (N_8107,N_7431,N_7788);
and U8108 (N_8108,N_7697,N_7978);
or U8109 (N_8109,N_7406,N_7062);
or U8110 (N_8110,N_7412,N_7196);
xnor U8111 (N_8111,N_7002,N_7831);
xor U8112 (N_8112,N_7504,N_7945);
and U8113 (N_8113,N_7618,N_7948);
nand U8114 (N_8114,N_7283,N_7305);
or U8115 (N_8115,N_7512,N_7112);
nand U8116 (N_8116,N_7382,N_7377);
nor U8117 (N_8117,N_7596,N_7253);
or U8118 (N_8118,N_7395,N_7054);
nand U8119 (N_8119,N_7523,N_7466);
nor U8120 (N_8120,N_7801,N_7234);
nor U8121 (N_8121,N_7178,N_7634);
nor U8122 (N_8122,N_7747,N_7107);
xnor U8123 (N_8123,N_7173,N_7714);
xor U8124 (N_8124,N_7856,N_7872);
nand U8125 (N_8125,N_7398,N_7861);
nand U8126 (N_8126,N_7557,N_7513);
or U8127 (N_8127,N_7965,N_7600);
xor U8128 (N_8128,N_7036,N_7492);
xor U8129 (N_8129,N_7996,N_7467);
or U8130 (N_8130,N_7292,N_7212);
xor U8131 (N_8131,N_7937,N_7383);
or U8132 (N_8132,N_7674,N_7552);
nor U8133 (N_8133,N_7297,N_7839);
nand U8134 (N_8134,N_7900,N_7542);
or U8135 (N_8135,N_7702,N_7215);
xor U8136 (N_8136,N_7718,N_7781);
or U8137 (N_8137,N_7392,N_7802);
nor U8138 (N_8138,N_7898,N_7724);
xor U8139 (N_8139,N_7405,N_7124);
xor U8140 (N_8140,N_7589,N_7815);
nand U8141 (N_8141,N_7063,N_7416);
nor U8142 (N_8142,N_7713,N_7374);
nand U8143 (N_8143,N_7187,N_7914);
or U8144 (N_8144,N_7949,N_7916);
xnor U8145 (N_8145,N_7137,N_7419);
nor U8146 (N_8146,N_7532,N_7229);
and U8147 (N_8147,N_7855,N_7449);
xor U8148 (N_8148,N_7812,N_7807);
nand U8149 (N_8149,N_7205,N_7808);
nor U8150 (N_8150,N_7318,N_7287);
nor U8151 (N_8151,N_7873,N_7539);
or U8152 (N_8152,N_7564,N_7300);
nor U8153 (N_8153,N_7796,N_7055);
nand U8154 (N_8154,N_7598,N_7586);
and U8155 (N_8155,N_7344,N_7067);
xnor U8156 (N_8156,N_7594,N_7742);
and U8157 (N_8157,N_7679,N_7734);
and U8158 (N_8158,N_7520,N_7308);
nand U8159 (N_8159,N_7188,N_7424);
nor U8160 (N_8160,N_7845,N_7498);
nor U8161 (N_8161,N_7105,N_7337);
and U8162 (N_8162,N_7022,N_7317);
or U8163 (N_8163,N_7460,N_7869);
nor U8164 (N_8164,N_7652,N_7032);
or U8165 (N_8165,N_7254,N_7908);
or U8166 (N_8166,N_7723,N_7456);
nor U8167 (N_8167,N_7785,N_7943);
and U8168 (N_8168,N_7870,N_7388);
or U8169 (N_8169,N_7010,N_7896);
nor U8170 (N_8170,N_7825,N_7249);
nor U8171 (N_8171,N_7732,N_7541);
nor U8172 (N_8172,N_7754,N_7617);
nand U8173 (N_8173,N_7826,N_7947);
or U8174 (N_8174,N_7214,N_7569);
xor U8175 (N_8175,N_7482,N_7765);
and U8176 (N_8176,N_7566,N_7306);
xor U8177 (N_8177,N_7065,N_7687);
or U8178 (N_8178,N_7255,N_7122);
or U8179 (N_8179,N_7716,N_7103);
and U8180 (N_8180,N_7068,N_7313);
and U8181 (N_8181,N_7030,N_7974);
xnor U8182 (N_8182,N_7073,N_7550);
and U8183 (N_8183,N_7701,N_7459);
nand U8184 (N_8184,N_7151,N_7141);
xor U8185 (N_8185,N_7487,N_7602);
and U8186 (N_8186,N_7803,N_7867);
or U8187 (N_8187,N_7866,N_7140);
xnor U8188 (N_8188,N_7100,N_7200);
nor U8189 (N_8189,N_7139,N_7649);
or U8190 (N_8190,N_7985,N_7003);
nor U8191 (N_8191,N_7986,N_7775);
nor U8192 (N_8192,N_7787,N_7150);
or U8193 (N_8193,N_7891,N_7893);
nand U8194 (N_8194,N_7911,N_7251);
and U8195 (N_8195,N_7066,N_7925);
and U8196 (N_8196,N_7797,N_7537);
and U8197 (N_8197,N_7017,N_7126);
nand U8198 (N_8198,N_7846,N_7739);
or U8199 (N_8199,N_7556,N_7399);
nand U8200 (N_8200,N_7533,N_7260);
xor U8201 (N_8201,N_7115,N_7147);
xor U8202 (N_8202,N_7669,N_7429);
and U8203 (N_8203,N_7485,N_7757);
nand U8204 (N_8204,N_7385,N_7546);
nor U8205 (N_8205,N_7087,N_7654);
and U8206 (N_8206,N_7368,N_7766);
xnor U8207 (N_8207,N_7019,N_7816);
nor U8208 (N_8208,N_7121,N_7064);
and U8209 (N_8209,N_7134,N_7983);
nand U8210 (N_8210,N_7645,N_7501);
nand U8211 (N_8211,N_7026,N_7098);
nand U8212 (N_8212,N_7998,N_7127);
or U8213 (N_8213,N_7425,N_7489);
xor U8214 (N_8214,N_7909,N_7074);
or U8215 (N_8215,N_7712,N_7989);
nor U8216 (N_8216,N_7875,N_7376);
and U8217 (N_8217,N_7369,N_7833);
nor U8218 (N_8218,N_7021,N_7667);
or U8219 (N_8219,N_7167,N_7404);
nor U8220 (N_8220,N_7800,N_7973);
nor U8221 (N_8221,N_7070,N_7892);
or U8222 (N_8222,N_7371,N_7346);
or U8223 (N_8223,N_7216,N_7610);
and U8224 (N_8224,N_7967,N_7131);
nand U8225 (N_8225,N_7307,N_7125);
nor U8226 (N_8226,N_7325,N_7051);
or U8227 (N_8227,N_7761,N_7962);
nand U8228 (N_8228,N_7695,N_7991);
or U8229 (N_8229,N_7298,N_7397);
nor U8230 (N_8230,N_7824,N_7958);
nand U8231 (N_8231,N_7806,N_7320);
nand U8232 (N_8232,N_7414,N_7015);
xnor U8233 (N_8233,N_7242,N_7581);
xnor U8234 (N_8234,N_7077,N_7271);
nand U8235 (N_8235,N_7220,N_7160);
and U8236 (N_8236,N_7358,N_7938);
nand U8237 (N_8237,N_7590,N_7844);
xnor U8238 (N_8238,N_7379,N_7577);
or U8239 (N_8239,N_7430,N_7623);
and U8240 (N_8240,N_7886,N_7391);
and U8241 (N_8241,N_7035,N_7027);
nand U8242 (N_8242,N_7082,N_7339);
nand U8243 (N_8243,N_7481,N_7365);
nor U8244 (N_8244,N_7984,N_7890);
and U8245 (N_8245,N_7615,N_7558);
and U8246 (N_8246,N_7464,N_7114);
nand U8247 (N_8247,N_7540,N_7698);
and U8248 (N_8248,N_7599,N_7740);
nor U8249 (N_8249,N_7849,N_7673);
xnor U8250 (N_8250,N_7791,N_7959);
nand U8251 (N_8251,N_7746,N_7932);
xnor U8252 (N_8252,N_7903,N_7149);
xor U8253 (N_8253,N_7162,N_7415);
nor U8254 (N_8254,N_7034,N_7232);
nor U8255 (N_8255,N_7593,N_7881);
and U8256 (N_8256,N_7013,N_7207);
xnor U8257 (N_8257,N_7536,N_7191);
or U8258 (N_8258,N_7491,N_7299);
nand U8259 (N_8259,N_7889,N_7643);
and U8260 (N_8260,N_7910,N_7858);
or U8261 (N_8261,N_7789,N_7621);
or U8262 (N_8262,N_7471,N_7172);
nand U8263 (N_8263,N_7864,N_7622);
or U8264 (N_8264,N_7917,N_7555);
xor U8265 (N_8265,N_7711,N_7608);
xor U8266 (N_8266,N_7857,N_7585);
nand U8267 (N_8267,N_7031,N_7575);
nor U8268 (N_8268,N_7331,N_7145);
and U8269 (N_8269,N_7053,N_7078);
or U8270 (N_8270,N_7877,N_7373);
xnor U8271 (N_8271,N_7276,N_7790);
xnor U8272 (N_8272,N_7745,N_7014);
nand U8273 (N_8273,N_7583,N_7158);
or U8274 (N_8274,N_7143,N_7079);
nor U8275 (N_8275,N_7280,N_7152);
nand U8276 (N_8276,N_7352,N_7244);
or U8277 (N_8277,N_7472,N_7111);
xor U8278 (N_8278,N_7256,N_7224);
or U8279 (N_8279,N_7963,N_7901);
or U8280 (N_8280,N_7641,N_7928);
or U8281 (N_8281,N_7439,N_7168);
xnor U8282 (N_8282,N_7868,N_7326);
and U8283 (N_8283,N_7047,N_7250);
nor U8284 (N_8284,N_7495,N_7436);
and U8285 (N_8285,N_7852,N_7408);
nor U8286 (N_8286,N_7567,N_7403);
nand U8287 (N_8287,N_7763,N_7023);
nor U8288 (N_8288,N_7341,N_7678);
nand U8289 (N_8289,N_7060,N_7970);
and U8290 (N_8290,N_7029,N_7941);
xnor U8291 (N_8291,N_7476,N_7189);
nor U8292 (N_8292,N_7821,N_7129);
nand U8293 (N_8293,N_7838,N_7239);
xnor U8294 (N_8294,N_7680,N_7549);
nor U8295 (N_8295,N_7478,N_7426);
nand U8296 (N_8296,N_7534,N_7729);
nand U8297 (N_8297,N_7428,N_7619);
nand U8298 (N_8298,N_7386,N_7367);
and U8299 (N_8299,N_7451,N_7530);
nor U8300 (N_8300,N_7725,N_7442);
xnor U8301 (N_8301,N_7153,N_7095);
or U8302 (N_8302,N_7483,N_7770);
nor U8303 (N_8303,N_7545,N_7319);
xor U8304 (N_8304,N_7665,N_7777);
nand U8305 (N_8305,N_7518,N_7443);
and U8306 (N_8306,N_7332,N_7632);
nand U8307 (N_8307,N_7551,N_7288);
nor U8308 (N_8308,N_7039,N_7372);
nor U8309 (N_8309,N_7380,N_7666);
xnor U8310 (N_8310,N_7235,N_7161);
or U8311 (N_8311,N_7311,N_7850);
nand U8312 (N_8312,N_7052,N_7302);
nor U8313 (N_8313,N_7538,N_7041);
and U8314 (N_8314,N_7862,N_7028);
and U8315 (N_8315,N_7146,N_7413);
and U8316 (N_8316,N_7452,N_7042);
nor U8317 (N_8317,N_7056,N_7199);
and U8318 (N_8318,N_7592,N_7262);
or U8319 (N_8319,N_7694,N_7304);
nor U8320 (N_8320,N_7166,N_7720);
or U8321 (N_8321,N_7273,N_7044);
nand U8322 (N_8322,N_7774,N_7059);
nand U8323 (N_8323,N_7159,N_7907);
and U8324 (N_8324,N_7099,N_7851);
nand U8325 (N_8325,N_7814,N_7316);
and U8326 (N_8326,N_7327,N_7926);
xnor U8327 (N_8327,N_7290,N_7496);
or U8328 (N_8328,N_7999,N_7389);
nor U8329 (N_8329,N_7164,N_7279);
nor U8330 (N_8330,N_7156,N_7792);
xnor U8331 (N_8331,N_7463,N_7221);
nor U8332 (N_8332,N_7410,N_7264);
nand U8333 (N_8333,N_7809,N_7971);
nor U8334 (N_8334,N_7012,N_7936);
xor U8335 (N_8335,N_7227,N_7190);
nor U8336 (N_8336,N_7576,N_7681);
xor U8337 (N_8337,N_7582,N_7018);
nor U8338 (N_8338,N_7089,N_7335);
and U8339 (N_8339,N_7847,N_7040);
and U8340 (N_8340,N_7081,N_7350);
or U8341 (N_8341,N_7057,N_7584);
and U8342 (N_8342,N_7285,N_7277);
or U8343 (N_8343,N_7123,N_7750);
or U8344 (N_8344,N_7440,N_7001);
xor U8345 (N_8345,N_7764,N_7644);
or U8346 (N_8346,N_7155,N_7357);
and U8347 (N_8347,N_7930,N_7135);
or U8348 (N_8348,N_7657,N_7267);
nand U8349 (N_8349,N_7755,N_7084);
and U8350 (N_8350,N_7884,N_7960);
and U8351 (N_8351,N_7647,N_7240);
or U8352 (N_8352,N_7455,N_7762);
and U8353 (N_8353,N_7441,N_7458);
nor U8354 (N_8354,N_7597,N_7772);
or U8355 (N_8355,N_7961,N_7469);
or U8356 (N_8356,N_7148,N_7830);
nor U8357 (N_8357,N_7048,N_7580);
and U8358 (N_8358,N_7075,N_7025);
or U8359 (N_8359,N_7923,N_7050);
nand U8360 (N_8360,N_7080,N_7524);
xor U8361 (N_8361,N_7987,N_7348);
nand U8362 (N_8362,N_7782,N_7284);
nor U8363 (N_8363,N_7686,N_7092);
nor U8364 (N_8364,N_7879,N_7366);
or U8365 (N_8365,N_7049,N_7660);
and U8366 (N_8366,N_7638,N_7499);
nand U8367 (N_8367,N_7130,N_7663);
or U8368 (N_8368,N_7354,N_7484);
xnor U8369 (N_8369,N_7194,N_7636);
or U8370 (N_8370,N_7954,N_7743);
or U8371 (N_8371,N_7969,N_7329);
xnor U8372 (N_8372,N_7046,N_7118);
or U8373 (N_8373,N_7929,N_7888);
and U8374 (N_8374,N_7922,N_7848);
nor U8375 (N_8375,N_7832,N_7918);
nand U8376 (N_8376,N_7885,N_7905);
or U8377 (N_8377,N_7715,N_7760);
and U8378 (N_8378,N_7091,N_7038);
nand U8379 (N_8379,N_7611,N_7037);
nand U8380 (N_8380,N_7268,N_7626);
xnor U8381 (N_8381,N_7511,N_7955);
nor U8382 (N_8382,N_7957,N_7509);
xnor U8383 (N_8383,N_7722,N_7605);
xor U8384 (N_8384,N_7805,N_7804);
or U8385 (N_8385,N_7422,N_7642);
nor U8386 (N_8386,N_7980,N_7488);
or U8387 (N_8387,N_7899,N_7336);
nand U8388 (N_8388,N_7997,N_7236);
xor U8389 (N_8389,N_7526,N_7378);
xnor U8390 (N_8390,N_7407,N_7375);
xnor U8391 (N_8391,N_7270,N_7561);
and U8392 (N_8392,N_7738,N_7004);
or U8393 (N_8393,N_7975,N_7692);
or U8394 (N_8394,N_7201,N_7203);
xor U8395 (N_8395,N_7007,N_7749);
or U8396 (N_8396,N_7226,N_7880);
nand U8397 (N_8397,N_7184,N_7935);
nand U8398 (N_8398,N_7629,N_7707);
nor U8399 (N_8399,N_7981,N_7717);
or U8400 (N_8400,N_7607,N_7952);
or U8401 (N_8401,N_7633,N_7438);
or U8402 (N_8402,N_7865,N_7982);
nand U8403 (N_8403,N_7208,N_7093);
nor U8404 (N_8404,N_7677,N_7310);
xnor U8405 (N_8405,N_7435,N_7860);
nand U8406 (N_8406,N_7176,N_7522);
or U8407 (N_8407,N_7450,N_7094);
nor U8408 (N_8408,N_7751,N_7058);
xnor U8409 (N_8409,N_7779,N_7956);
xor U8410 (N_8410,N_7113,N_7813);
nor U8411 (N_8411,N_7477,N_7353);
nand U8412 (N_8412,N_7470,N_7136);
nor U8413 (N_8413,N_7183,N_7676);
xor U8414 (N_8414,N_7246,N_7144);
xor U8415 (N_8415,N_7453,N_7338);
nand U8416 (N_8416,N_7480,N_7301);
and U8417 (N_8417,N_7793,N_7912);
nand U8418 (N_8418,N_7990,N_7931);
nor U8419 (N_8419,N_7968,N_7119);
or U8420 (N_8420,N_7418,N_7043);
nor U8421 (N_8421,N_7799,N_7490);
nand U8422 (N_8422,N_7370,N_7554);
nand U8423 (N_8423,N_7101,N_7840);
or U8424 (N_8424,N_7359,N_7748);
xnor U8425 (N_8425,N_7355,N_7728);
and U8426 (N_8426,N_7085,N_7994);
nand U8427 (N_8427,N_7527,N_7767);
xor U8428 (N_8428,N_7559,N_7110);
nor U8429 (N_8429,N_7653,N_7601);
nor U8430 (N_8430,N_7225,N_7457);
and U8431 (N_8431,N_7434,N_7794);
and U8432 (N_8432,N_7008,N_7818);
nand U8433 (N_8433,N_7737,N_7309);
or U8434 (N_8434,N_7494,N_7913);
and U8435 (N_8435,N_7921,N_7104);
nand U8436 (N_8436,N_7603,N_7261);
nor U8437 (N_8437,N_7979,N_7883);
or U8438 (N_8438,N_7579,N_7069);
or U8439 (N_8439,N_7553,N_7521);
nand U8440 (N_8440,N_7690,N_7175);
nand U8441 (N_8441,N_7238,N_7474);
nor U8442 (N_8442,N_7966,N_7685);
or U8443 (N_8443,N_7927,N_7363);
nand U8444 (N_8444,N_7217,N_7731);
or U8445 (N_8445,N_7479,N_7120);
xnor U8446 (N_8446,N_7394,N_7836);
or U8447 (N_8447,N_7528,N_7263);
nor U8448 (N_8448,N_7780,N_7700);
and U8449 (N_8449,N_7446,N_7169);
or U8450 (N_8450,N_7704,N_7563);
nor U8451 (N_8451,N_7988,N_7241);
xnor U8452 (N_8452,N_7661,N_7662);
and U8453 (N_8453,N_7195,N_7269);
nor U8454 (N_8454,N_7211,N_7515);
xor U8455 (N_8455,N_7871,N_7670);
or U8456 (N_8456,N_7612,N_7296);
and U8457 (N_8457,N_7228,N_7906);
nand U8458 (N_8458,N_7345,N_7020);
and U8459 (N_8459,N_7475,N_7180);
or U8460 (N_8460,N_7543,N_7529);
and U8461 (N_8461,N_7409,N_7547);
xor U8462 (N_8462,N_7735,N_7315);
nand U8463 (N_8463,N_7820,N_7508);
and U8464 (N_8464,N_7933,N_7682);
and U8465 (N_8465,N_7454,N_7659);
or U8466 (N_8466,N_7462,N_7684);
xnor U8467 (N_8467,N_7631,N_7347);
xnor U8468 (N_8468,N_7708,N_7265);
or U8469 (N_8469,N_7817,N_7045);
nand U8470 (N_8470,N_7420,N_7656);
nor U8471 (N_8471,N_7174,N_7895);
or U8472 (N_8472,N_7433,N_7206);
nand U8473 (N_8473,N_7627,N_7231);
nor U8474 (N_8474,N_7544,N_7843);
and U8475 (N_8475,N_7396,N_7322);
or U8476 (N_8476,N_7683,N_7786);
and U8477 (N_8477,N_7625,N_7204);
nand U8478 (N_8478,N_7689,N_7505);
and U8479 (N_8479,N_7417,N_7588);
nand U8480 (N_8480,N_7294,N_7061);
and U8481 (N_8481,N_7706,N_7258);
nand U8482 (N_8482,N_7953,N_7992);
and U8483 (N_8483,N_7705,N_7444);
or U8484 (N_8484,N_7606,N_7230);
and U8485 (N_8485,N_7324,N_7381);
and U8486 (N_8486,N_7163,N_7209);
nand U8487 (N_8487,N_7703,N_7635);
xor U8488 (N_8488,N_7257,N_7570);
or U8489 (N_8489,N_7192,N_7245);
xor U8490 (N_8490,N_7086,N_7303);
xnor U8491 (N_8491,N_7573,N_7951);
nor U8492 (N_8492,N_7096,N_7218);
or U8493 (N_8493,N_7648,N_7758);
or U8494 (N_8494,N_7142,N_7033);
nor U8495 (N_8495,N_7314,N_7266);
xnor U8496 (N_8496,N_7719,N_7859);
and U8497 (N_8497,N_7578,N_7333);
nand U8498 (N_8498,N_7165,N_7243);
or U8499 (N_8499,N_7432,N_7628);
and U8500 (N_8500,N_7077,N_7513);
nand U8501 (N_8501,N_7946,N_7047);
nor U8502 (N_8502,N_7381,N_7516);
and U8503 (N_8503,N_7373,N_7424);
and U8504 (N_8504,N_7763,N_7719);
or U8505 (N_8505,N_7550,N_7160);
and U8506 (N_8506,N_7065,N_7812);
nand U8507 (N_8507,N_7474,N_7333);
nor U8508 (N_8508,N_7490,N_7398);
or U8509 (N_8509,N_7076,N_7861);
or U8510 (N_8510,N_7779,N_7097);
nor U8511 (N_8511,N_7335,N_7270);
or U8512 (N_8512,N_7742,N_7905);
and U8513 (N_8513,N_7822,N_7731);
nand U8514 (N_8514,N_7846,N_7326);
nand U8515 (N_8515,N_7244,N_7812);
or U8516 (N_8516,N_7942,N_7948);
or U8517 (N_8517,N_7876,N_7465);
or U8518 (N_8518,N_7877,N_7972);
nor U8519 (N_8519,N_7356,N_7062);
or U8520 (N_8520,N_7443,N_7246);
or U8521 (N_8521,N_7048,N_7768);
or U8522 (N_8522,N_7098,N_7288);
nor U8523 (N_8523,N_7017,N_7949);
nand U8524 (N_8524,N_7201,N_7579);
nand U8525 (N_8525,N_7459,N_7178);
and U8526 (N_8526,N_7158,N_7010);
xnor U8527 (N_8527,N_7832,N_7381);
nand U8528 (N_8528,N_7176,N_7334);
and U8529 (N_8529,N_7468,N_7422);
and U8530 (N_8530,N_7631,N_7643);
nor U8531 (N_8531,N_7051,N_7524);
nand U8532 (N_8532,N_7471,N_7208);
xnor U8533 (N_8533,N_7818,N_7628);
nand U8534 (N_8534,N_7076,N_7077);
and U8535 (N_8535,N_7714,N_7148);
xor U8536 (N_8536,N_7241,N_7787);
nand U8537 (N_8537,N_7975,N_7570);
xor U8538 (N_8538,N_7761,N_7848);
and U8539 (N_8539,N_7699,N_7271);
xnor U8540 (N_8540,N_7435,N_7548);
or U8541 (N_8541,N_7506,N_7956);
and U8542 (N_8542,N_7160,N_7027);
or U8543 (N_8543,N_7143,N_7961);
nand U8544 (N_8544,N_7143,N_7907);
or U8545 (N_8545,N_7141,N_7227);
nand U8546 (N_8546,N_7608,N_7654);
xnor U8547 (N_8547,N_7489,N_7093);
xor U8548 (N_8548,N_7478,N_7379);
and U8549 (N_8549,N_7734,N_7065);
and U8550 (N_8550,N_7816,N_7002);
or U8551 (N_8551,N_7909,N_7545);
or U8552 (N_8552,N_7901,N_7411);
xor U8553 (N_8553,N_7030,N_7081);
nor U8554 (N_8554,N_7758,N_7732);
xor U8555 (N_8555,N_7607,N_7377);
and U8556 (N_8556,N_7697,N_7441);
nand U8557 (N_8557,N_7617,N_7660);
or U8558 (N_8558,N_7359,N_7683);
xor U8559 (N_8559,N_7060,N_7380);
and U8560 (N_8560,N_7518,N_7841);
or U8561 (N_8561,N_7701,N_7230);
nand U8562 (N_8562,N_7169,N_7797);
and U8563 (N_8563,N_7954,N_7814);
nor U8564 (N_8564,N_7147,N_7400);
or U8565 (N_8565,N_7763,N_7929);
and U8566 (N_8566,N_7725,N_7910);
xnor U8567 (N_8567,N_7745,N_7054);
nor U8568 (N_8568,N_7766,N_7375);
xor U8569 (N_8569,N_7161,N_7356);
or U8570 (N_8570,N_7531,N_7194);
nand U8571 (N_8571,N_7716,N_7290);
or U8572 (N_8572,N_7809,N_7687);
or U8573 (N_8573,N_7472,N_7016);
nand U8574 (N_8574,N_7835,N_7075);
and U8575 (N_8575,N_7223,N_7648);
and U8576 (N_8576,N_7383,N_7322);
xnor U8577 (N_8577,N_7326,N_7368);
and U8578 (N_8578,N_7770,N_7115);
xnor U8579 (N_8579,N_7978,N_7219);
xnor U8580 (N_8580,N_7427,N_7299);
or U8581 (N_8581,N_7230,N_7969);
nand U8582 (N_8582,N_7180,N_7076);
and U8583 (N_8583,N_7155,N_7105);
nor U8584 (N_8584,N_7542,N_7953);
and U8585 (N_8585,N_7800,N_7803);
nand U8586 (N_8586,N_7578,N_7612);
or U8587 (N_8587,N_7376,N_7321);
nor U8588 (N_8588,N_7037,N_7368);
and U8589 (N_8589,N_7801,N_7318);
and U8590 (N_8590,N_7260,N_7149);
or U8591 (N_8591,N_7448,N_7419);
and U8592 (N_8592,N_7954,N_7199);
nand U8593 (N_8593,N_7385,N_7852);
or U8594 (N_8594,N_7428,N_7598);
xor U8595 (N_8595,N_7456,N_7885);
and U8596 (N_8596,N_7743,N_7852);
nand U8597 (N_8597,N_7230,N_7077);
or U8598 (N_8598,N_7506,N_7825);
nand U8599 (N_8599,N_7917,N_7067);
and U8600 (N_8600,N_7061,N_7211);
and U8601 (N_8601,N_7414,N_7569);
or U8602 (N_8602,N_7200,N_7599);
and U8603 (N_8603,N_7636,N_7375);
xor U8604 (N_8604,N_7915,N_7191);
and U8605 (N_8605,N_7341,N_7242);
nand U8606 (N_8606,N_7183,N_7721);
nor U8607 (N_8607,N_7642,N_7046);
and U8608 (N_8608,N_7027,N_7159);
nor U8609 (N_8609,N_7719,N_7421);
xnor U8610 (N_8610,N_7592,N_7096);
xor U8611 (N_8611,N_7100,N_7207);
and U8612 (N_8612,N_7728,N_7265);
xnor U8613 (N_8613,N_7334,N_7163);
and U8614 (N_8614,N_7898,N_7814);
xor U8615 (N_8615,N_7907,N_7455);
and U8616 (N_8616,N_7659,N_7002);
and U8617 (N_8617,N_7283,N_7881);
or U8618 (N_8618,N_7350,N_7627);
or U8619 (N_8619,N_7889,N_7362);
nand U8620 (N_8620,N_7845,N_7974);
xnor U8621 (N_8621,N_7194,N_7450);
and U8622 (N_8622,N_7082,N_7999);
or U8623 (N_8623,N_7797,N_7461);
xnor U8624 (N_8624,N_7785,N_7538);
xor U8625 (N_8625,N_7205,N_7684);
nor U8626 (N_8626,N_7025,N_7027);
nor U8627 (N_8627,N_7463,N_7648);
nor U8628 (N_8628,N_7958,N_7940);
and U8629 (N_8629,N_7163,N_7765);
nor U8630 (N_8630,N_7162,N_7754);
or U8631 (N_8631,N_7733,N_7301);
xor U8632 (N_8632,N_7819,N_7285);
nor U8633 (N_8633,N_7413,N_7964);
xor U8634 (N_8634,N_7650,N_7633);
nor U8635 (N_8635,N_7061,N_7986);
and U8636 (N_8636,N_7058,N_7155);
nand U8637 (N_8637,N_7969,N_7828);
xnor U8638 (N_8638,N_7788,N_7002);
and U8639 (N_8639,N_7382,N_7023);
or U8640 (N_8640,N_7593,N_7282);
and U8641 (N_8641,N_7047,N_7452);
nor U8642 (N_8642,N_7530,N_7363);
xor U8643 (N_8643,N_7803,N_7761);
nor U8644 (N_8644,N_7965,N_7442);
xnor U8645 (N_8645,N_7646,N_7156);
nor U8646 (N_8646,N_7989,N_7343);
and U8647 (N_8647,N_7114,N_7043);
nor U8648 (N_8648,N_7165,N_7446);
xnor U8649 (N_8649,N_7069,N_7443);
xnor U8650 (N_8650,N_7534,N_7270);
and U8651 (N_8651,N_7001,N_7312);
nor U8652 (N_8652,N_7190,N_7013);
xor U8653 (N_8653,N_7001,N_7982);
xnor U8654 (N_8654,N_7260,N_7438);
nor U8655 (N_8655,N_7533,N_7020);
and U8656 (N_8656,N_7677,N_7833);
nand U8657 (N_8657,N_7996,N_7031);
xnor U8658 (N_8658,N_7249,N_7837);
or U8659 (N_8659,N_7400,N_7299);
xor U8660 (N_8660,N_7735,N_7714);
nand U8661 (N_8661,N_7112,N_7049);
nand U8662 (N_8662,N_7695,N_7529);
and U8663 (N_8663,N_7600,N_7043);
nand U8664 (N_8664,N_7764,N_7097);
or U8665 (N_8665,N_7202,N_7059);
nand U8666 (N_8666,N_7142,N_7327);
and U8667 (N_8667,N_7736,N_7796);
nor U8668 (N_8668,N_7851,N_7372);
nor U8669 (N_8669,N_7581,N_7941);
and U8670 (N_8670,N_7960,N_7470);
nand U8671 (N_8671,N_7607,N_7328);
and U8672 (N_8672,N_7352,N_7880);
nor U8673 (N_8673,N_7440,N_7452);
and U8674 (N_8674,N_7621,N_7355);
nand U8675 (N_8675,N_7068,N_7958);
or U8676 (N_8676,N_7820,N_7380);
or U8677 (N_8677,N_7484,N_7575);
xor U8678 (N_8678,N_7043,N_7191);
and U8679 (N_8679,N_7466,N_7240);
or U8680 (N_8680,N_7361,N_7057);
nand U8681 (N_8681,N_7653,N_7640);
nor U8682 (N_8682,N_7672,N_7114);
nand U8683 (N_8683,N_7247,N_7979);
or U8684 (N_8684,N_7544,N_7074);
and U8685 (N_8685,N_7054,N_7719);
and U8686 (N_8686,N_7637,N_7940);
and U8687 (N_8687,N_7341,N_7066);
or U8688 (N_8688,N_7953,N_7420);
xor U8689 (N_8689,N_7524,N_7457);
nor U8690 (N_8690,N_7828,N_7993);
xor U8691 (N_8691,N_7987,N_7775);
nand U8692 (N_8692,N_7285,N_7587);
and U8693 (N_8693,N_7596,N_7681);
nor U8694 (N_8694,N_7759,N_7044);
nand U8695 (N_8695,N_7655,N_7766);
or U8696 (N_8696,N_7054,N_7646);
xnor U8697 (N_8697,N_7077,N_7079);
and U8698 (N_8698,N_7342,N_7056);
nand U8699 (N_8699,N_7877,N_7843);
nand U8700 (N_8700,N_7169,N_7458);
or U8701 (N_8701,N_7926,N_7849);
or U8702 (N_8702,N_7543,N_7434);
nand U8703 (N_8703,N_7889,N_7548);
xnor U8704 (N_8704,N_7524,N_7854);
or U8705 (N_8705,N_7990,N_7496);
xnor U8706 (N_8706,N_7196,N_7978);
nand U8707 (N_8707,N_7491,N_7484);
or U8708 (N_8708,N_7205,N_7698);
nor U8709 (N_8709,N_7421,N_7431);
nor U8710 (N_8710,N_7633,N_7170);
and U8711 (N_8711,N_7345,N_7499);
nand U8712 (N_8712,N_7200,N_7135);
xor U8713 (N_8713,N_7215,N_7451);
and U8714 (N_8714,N_7460,N_7211);
or U8715 (N_8715,N_7063,N_7542);
and U8716 (N_8716,N_7540,N_7996);
and U8717 (N_8717,N_7099,N_7175);
nor U8718 (N_8718,N_7000,N_7562);
and U8719 (N_8719,N_7049,N_7366);
nor U8720 (N_8720,N_7665,N_7283);
nor U8721 (N_8721,N_7160,N_7596);
nand U8722 (N_8722,N_7994,N_7454);
and U8723 (N_8723,N_7418,N_7758);
nand U8724 (N_8724,N_7008,N_7474);
and U8725 (N_8725,N_7607,N_7708);
and U8726 (N_8726,N_7345,N_7615);
nor U8727 (N_8727,N_7048,N_7512);
or U8728 (N_8728,N_7475,N_7925);
or U8729 (N_8729,N_7647,N_7399);
nand U8730 (N_8730,N_7192,N_7546);
nor U8731 (N_8731,N_7954,N_7336);
nor U8732 (N_8732,N_7526,N_7545);
nor U8733 (N_8733,N_7828,N_7234);
nand U8734 (N_8734,N_7994,N_7360);
nand U8735 (N_8735,N_7589,N_7031);
nor U8736 (N_8736,N_7324,N_7325);
xor U8737 (N_8737,N_7231,N_7150);
nand U8738 (N_8738,N_7011,N_7445);
xnor U8739 (N_8739,N_7038,N_7931);
nor U8740 (N_8740,N_7476,N_7042);
or U8741 (N_8741,N_7640,N_7825);
or U8742 (N_8742,N_7789,N_7165);
nand U8743 (N_8743,N_7433,N_7443);
nand U8744 (N_8744,N_7463,N_7510);
or U8745 (N_8745,N_7143,N_7777);
xnor U8746 (N_8746,N_7527,N_7202);
xor U8747 (N_8747,N_7857,N_7596);
nor U8748 (N_8748,N_7208,N_7218);
xnor U8749 (N_8749,N_7925,N_7229);
and U8750 (N_8750,N_7809,N_7581);
or U8751 (N_8751,N_7421,N_7773);
nor U8752 (N_8752,N_7744,N_7297);
and U8753 (N_8753,N_7136,N_7803);
xor U8754 (N_8754,N_7724,N_7115);
nor U8755 (N_8755,N_7336,N_7820);
or U8756 (N_8756,N_7170,N_7715);
nand U8757 (N_8757,N_7908,N_7576);
xnor U8758 (N_8758,N_7888,N_7692);
and U8759 (N_8759,N_7358,N_7512);
nand U8760 (N_8760,N_7127,N_7178);
or U8761 (N_8761,N_7511,N_7153);
xor U8762 (N_8762,N_7071,N_7279);
and U8763 (N_8763,N_7448,N_7239);
xnor U8764 (N_8764,N_7430,N_7233);
and U8765 (N_8765,N_7088,N_7603);
nor U8766 (N_8766,N_7647,N_7699);
and U8767 (N_8767,N_7672,N_7082);
nor U8768 (N_8768,N_7670,N_7798);
and U8769 (N_8769,N_7614,N_7647);
and U8770 (N_8770,N_7693,N_7884);
or U8771 (N_8771,N_7260,N_7616);
or U8772 (N_8772,N_7044,N_7590);
nand U8773 (N_8773,N_7901,N_7566);
or U8774 (N_8774,N_7706,N_7089);
nor U8775 (N_8775,N_7189,N_7653);
and U8776 (N_8776,N_7001,N_7549);
xnor U8777 (N_8777,N_7118,N_7774);
nor U8778 (N_8778,N_7282,N_7967);
xor U8779 (N_8779,N_7586,N_7780);
or U8780 (N_8780,N_7482,N_7139);
xnor U8781 (N_8781,N_7142,N_7716);
or U8782 (N_8782,N_7034,N_7598);
and U8783 (N_8783,N_7546,N_7725);
or U8784 (N_8784,N_7545,N_7298);
nor U8785 (N_8785,N_7356,N_7349);
or U8786 (N_8786,N_7933,N_7275);
nor U8787 (N_8787,N_7599,N_7217);
or U8788 (N_8788,N_7081,N_7228);
and U8789 (N_8789,N_7690,N_7584);
nand U8790 (N_8790,N_7445,N_7168);
or U8791 (N_8791,N_7306,N_7626);
xnor U8792 (N_8792,N_7023,N_7602);
and U8793 (N_8793,N_7487,N_7425);
xor U8794 (N_8794,N_7722,N_7679);
nand U8795 (N_8795,N_7414,N_7107);
and U8796 (N_8796,N_7061,N_7203);
and U8797 (N_8797,N_7487,N_7279);
xor U8798 (N_8798,N_7847,N_7961);
and U8799 (N_8799,N_7558,N_7052);
nor U8800 (N_8800,N_7055,N_7107);
nor U8801 (N_8801,N_7790,N_7640);
or U8802 (N_8802,N_7695,N_7614);
and U8803 (N_8803,N_7003,N_7740);
xor U8804 (N_8804,N_7753,N_7015);
nand U8805 (N_8805,N_7444,N_7795);
and U8806 (N_8806,N_7145,N_7406);
nor U8807 (N_8807,N_7827,N_7754);
xnor U8808 (N_8808,N_7320,N_7424);
and U8809 (N_8809,N_7166,N_7161);
and U8810 (N_8810,N_7998,N_7860);
or U8811 (N_8811,N_7822,N_7967);
nor U8812 (N_8812,N_7500,N_7344);
nand U8813 (N_8813,N_7098,N_7325);
nor U8814 (N_8814,N_7900,N_7396);
xor U8815 (N_8815,N_7835,N_7666);
nor U8816 (N_8816,N_7050,N_7307);
nor U8817 (N_8817,N_7216,N_7691);
nand U8818 (N_8818,N_7955,N_7227);
or U8819 (N_8819,N_7458,N_7983);
nand U8820 (N_8820,N_7626,N_7892);
and U8821 (N_8821,N_7203,N_7718);
and U8822 (N_8822,N_7489,N_7060);
or U8823 (N_8823,N_7290,N_7591);
or U8824 (N_8824,N_7967,N_7806);
nor U8825 (N_8825,N_7721,N_7683);
nor U8826 (N_8826,N_7713,N_7104);
xor U8827 (N_8827,N_7607,N_7654);
or U8828 (N_8828,N_7998,N_7379);
xor U8829 (N_8829,N_7838,N_7455);
and U8830 (N_8830,N_7313,N_7706);
nand U8831 (N_8831,N_7294,N_7269);
or U8832 (N_8832,N_7662,N_7134);
and U8833 (N_8833,N_7814,N_7522);
and U8834 (N_8834,N_7903,N_7691);
nor U8835 (N_8835,N_7742,N_7211);
nor U8836 (N_8836,N_7361,N_7012);
xor U8837 (N_8837,N_7711,N_7620);
and U8838 (N_8838,N_7368,N_7507);
xnor U8839 (N_8839,N_7670,N_7869);
nand U8840 (N_8840,N_7471,N_7549);
or U8841 (N_8841,N_7350,N_7773);
nand U8842 (N_8842,N_7845,N_7783);
or U8843 (N_8843,N_7363,N_7951);
xor U8844 (N_8844,N_7088,N_7797);
nor U8845 (N_8845,N_7171,N_7515);
nand U8846 (N_8846,N_7474,N_7108);
xnor U8847 (N_8847,N_7887,N_7191);
nand U8848 (N_8848,N_7425,N_7145);
and U8849 (N_8849,N_7980,N_7398);
and U8850 (N_8850,N_7331,N_7291);
or U8851 (N_8851,N_7849,N_7546);
or U8852 (N_8852,N_7549,N_7767);
or U8853 (N_8853,N_7315,N_7609);
nand U8854 (N_8854,N_7519,N_7205);
xnor U8855 (N_8855,N_7489,N_7389);
and U8856 (N_8856,N_7897,N_7033);
and U8857 (N_8857,N_7606,N_7559);
xnor U8858 (N_8858,N_7583,N_7596);
xnor U8859 (N_8859,N_7696,N_7737);
or U8860 (N_8860,N_7745,N_7868);
xnor U8861 (N_8861,N_7853,N_7329);
and U8862 (N_8862,N_7693,N_7414);
and U8863 (N_8863,N_7839,N_7254);
xnor U8864 (N_8864,N_7926,N_7435);
nor U8865 (N_8865,N_7183,N_7205);
xnor U8866 (N_8866,N_7781,N_7590);
xnor U8867 (N_8867,N_7290,N_7619);
or U8868 (N_8868,N_7458,N_7409);
nor U8869 (N_8869,N_7404,N_7063);
and U8870 (N_8870,N_7815,N_7003);
nor U8871 (N_8871,N_7294,N_7817);
nor U8872 (N_8872,N_7779,N_7419);
nor U8873 (N_8873,N_7404,N_7505);
or U8874 (N_8874,N_7109,N_7795);
nand U8875 (N_8875,N_7615,N_7535);
and U8876 (N_8876,N_7102,N_7046);
xor U8877 (N_8877,N_7190,N_7780);
nor U8878 (N_8878,N_7081,N_7443);
and U8879 (N_8879,N_7927,N_7530);
nand U8880 (N_8880,N_7817,N_7417);
and U8881 (N_8881,N_7983,N_7481);
nand U8882 (N_8882,N_7284,N_7842);
nand U8883 (N_8883,N_7859,N_7899);
nand U8884 (N_8884,N_7792,N_7464);
xor U8885 (N_8885,N_7908,N_7912);
xor U8886 (N_8886,N_7323,N_7029);
nor U8887 (N_8887,N_7363,N_7511);
and U8888 (N_8888,N_7410,N_7093);
xor U8889 (N_8889,N_7259,N_7017);
or U8890 (N_8890,N_7694,N_7770);
nand U8891 (N_8891,N_7382,N_7101);
and U8892 (N_8892,N_7337,N_7469);
nand U8893 (N_8893,N_7135,N_7099);
xnor U8894 (N_8894,N_7974,N_7486);
nand U8895 (N_8895,N_7629,N_7599);
nand U8896 (N_8896,N_7122,N_7477);
xor U8897 (N_8897,N_7851,N_7836);
and U8898 (N_8898,N_7725,N_7890);
xor U8899 (N_8899,N_7849,N_7447);
xnor U8900 (N_8900,N_7850,N_7009);
nand U8901 (N_8901,N_7449,N_7615);
nand U8902 (N_8902,N_7942,N_7547);
and U8903 (N_8903,N_7190,N_7322);
and U8904 (N_8904,N_7226,N_7715);
nor U8905 (N_8905,N_7664,N_7310);
nor U8906 (N_8906,N_7425,N_7942);
and U8907 (N_8907,N_7452,N_7696);
nor U8908 (N_8908,N_7004,N_7812);
and U8909 (N_8909,N_7813,N_7698);
nor U8910 (N_8910,N_7516,N_7646);
xnor U8911 (N_8911,N_7728,N_7161);
or U8912 (N_8912,N_7555,N_7103);
nand U8913 (N_8913,N_7715,N_7858);
nand U8914 (N_8914,N_7492,N_7509);
nor U8915 (N_8915,N_7497,N_7369);
nand U8916 (N_8916,N_7738,N_7287);
and U8917 (N_8917,N_7422,N_7972);
xor U8918 (N_8918,N_7703,N_7837);
xor U8919 (N_8919,N_7585,N_7881);
or U8920 (N_8920,N_7365,N_7850);
nand U8921 (N_8921,N_7463,N_7849);
nand U8922 (N_8922,N_7650,N_7956);
xnor U8923 (N_8923,N_7162,N_7123);
and U8924 (N_8924,N_7636,N_7347);
and U8925 (N_8925,N_7856,N_7458);
nor U8926 (N_8926,N_7226,N_7118);
xor U8927 (N_8927,N_7362,N_7545);
nor U8928 (N_8928,N_7445,N_7004);
nor U8929 (N_8929,N_7930,N_7424);
and U8930 (N_8930,N_7575,N_7374);
xnor U8931 (N_8931,N_7290,N_7045);
xnor U8932 (N_8932,N_7567,N_7634);
and U8933 (N_8933,N_7219,N_7577);
xor U8934 (N_8934,N_7447,N_7373);
or U8935 (N_8935,N_7923,N_7873);
nor U8936 (N_8936,N_7937,N_7443);
and U8937 (N_8937,N_7186,N_7322);
nor U8938 (N_8938,N_7207,N_7146);
nor U8939 (N_8939,N_7099,N_7934);
xor U8940 (N_8940,N_7501,N_7770);
or U8941 (N_8941,N_7561,N_7763);
nor U8942 (N_8942,N_7602,N_7846);
nor U8943 (N_8943,N_7216,N_7382);
nor U8944 (N_8944,N_7997,N_7307);
nor U8945 (N_8945,N_7965,N_7210);
nor U8946 (N_8946,N_7900,N_7050);
nor U8947 (N_8947,N_7156,N_7244);
or U8948 (N_8948,N_7524,N_7774);
and U8949 (N_8949,N_7288,N_7061);
xnor U8950 (N_8950,N_7044,N_7694);
or U8951 (N_8951,N_7857,N_7305);
xnor U8952 (N_8952,N_7557,N_7261);
and U8953 (N_8953,N_7012,N_7027);
nor U8954 (N_8954,N_7032,N_7064);
or U8955 (N_8955,N_7240,N_7588);
nand U8956 (N_8956,N_7453,N_7587);
nand U8957 (N_8957,N_7844,N_7915);
nand U8958 (N_8958,N_7215,N_7648);
nor U8959 (N_8959,N_7072,N_7800);
xor U8960 (N_8960,N_7857,N_7804);
nor U8961 (N_8961,N_7131,N_7046);
nand U8962 (N_8962,N_7382,N_7322);
nor U8963 (N_8963,N_7717,N_7120);
or U8964 (N_8964,N_7450,N_7087);
nor U8965 (N_8965,N_7409,N_7281);
or U8966 (N_8966,N_7640,N_7377);
nor U8967 (N_8967,N_7939,N_7607);
xor U8968 (N_8968,N_7184,N_7518);
nor U8969 (N_8969,N_7982,N_7108);
nor U8970 (N_8970,N_7910,N_7591);
or U8971 (N_8971,N_7507,N_7553);
xnor U8972 (N_8972,N_7435,N_7871);
nor U8973 (N_8973,N_7078,N_7619);
nand U8974 (N_8974,N_7877,N_7588);
nand U8975 (N_8975,N_7301,N_7333);
nand U8976 (N_8976,N_7722,N_7863);
xor U8977 (N_8977,N_7852,N_7249);
xor U8978 (N_8978,N_7473,N_7695);
nand U8979 (N_8979,N_7905,N_7434);
nor U8980 (N_8980,N_7543,N_7125);
or U8981 (N_8981,N_7896,N_7812);
nand U8982 (N_8982,N_7597,N_7519);
or U8983 (N_8983,N_7870,N_7742);
or U8984 (N_8984,N_7509,N_7663);
xor U8985 (N_8985,N_7852,N_7454);
nor U8986 (N_8986,N_7036,N_7353);
or U8987 (N_8987,N_7306,N_7774);
xor U8988 (N_8988,N_7764,N_7888);
and U8989 (N_8989,N_7634,N_7811);
xor U8990 (N_8990,N_7969,N_7045);
nor U8991 (N_8991,N_7074,N_7278);
xor U8992 (N_8992,N_7800,N_7361);
xnor U8993 (N_8993,N_7172,N_7357);
nand U8994 (N_8994,N_7521,N_7644);
or U8995 (N_8995,N_7302,N_7144);
and U8996 (N_8996,N_7560,N_7931);
and U8997 (N_8997,N_7181,N_7667);
or U8998 (N_8998,N_7596,N_7135);
or U8999 (N_8999,N_7989,N_7675);
or U9000 (N_9000,N_8873,N_8240);
nor U9001 (N_9001,N_8563,N_8609);
nand U9002 (N_9002,N_8279,N_8364);
nand U9003 (N_9003,N_8166,N_8742);
and U9004 (N_9004,N_8352,N_8865);
xnor U9005 (N_9005,N_8646,N_8186);
and U9006 (N_9006,N_8158,N_8581);
nor U9007 (N_9007,N_8263,N_8714);
nor U9008 (N_9008,N_8383,N_8586);
or U9009 (N_9009,N_8784,N_8132);
nand U9010 (N_9010,N_8244,N_8533);
xor U9011 (N_9011,N_8971,N_8256);
and U9012 (N_9012,N_8621,N_8718);
nand U9013 (N_9013,N_8031,N_8973);
and U9014 (N_9014,N_8068,N_8937);
nor U9015 (N_9015,N_8974,N_8192);
and U9016 (N_9016,N_8443,N_8866);
nand U9017 (N_9017,N_8819,N_8765);
or U9018 (N_9018,N_8537,N_8982);
or U9019 (N_9019,N_8618,N_8454);
nand U9020 (N_9020,N_8408,N_8853);
nand U9021 (N_9021,N_8874,N_8938);
and U9022 (N_9022,N_8835,N_8210);
nand U9023 (N_9023,N_8350,N_8074);
nor U9024 (N_9024,N_8117,N_8374);
xor U9025 (N_9025,N_8947,N_8107);
nand U9026 (N_9026,N_8859,N_8562);
or U9027 (N_9027,N_8486,N_8410);
and U9028 (N_9028,N_8401,N_8257);
nand U9029 (N_9029,N_8536,N_8530);
and U9030 (N_9030,N_8936,N_8990);
or U9031 (N_9031,N_8312,N_8195);
nand U9032 (N_9032,N_8558,N_8962);
nand U9033 (N_9033,N_8333,N_8125);
or U9034 (N_9034,N_8073,N_8612);
or U9035 (N_9035,N_8918,N_8392);
xor U9036 (N_9036,N_8991,N_8684);
nor U9037 (N_9037,N_8395,N_8721);
nand U9038 (N_9038,N_8082,N_8453);
xnor U9039 (N_9039,N_8177,N_8541);
and U9040 (N_9040,N_8067,N_8850);
nand U9041 (N_9041,N_8596,N_8422);
xnor U9042 (N_9042,N_8003,N_8292);
or U9043 (N_9043,N_8844,N_8245);
or U9044 (N_9044,N_8092,N_8522);
or U9045 (N_9045,N_8012,N_8322);
nor U9046 (N_9046,N_8431,N_8281);
nand U9047 (N_9047,N_8911,N_8801);
nand U9048 (N_9048,N_8269,N_8775);
nand U9049 (N_9049,N_8923,N_8642);
and U9050 (N_9050,N_8371,N_8075);
nand U9051 (N_9051,N_8808,N_8055);
xor U9052 (N_9052,N_8899,N_8216);
and U9053 (N_9053,N_8314,N_8193);
nand U9054 (N_9054,N_8429,N_8298);
xnor U9055 (N_9055,N_8228,N_8397);
or U9056 (N_9056,N_8128,N_8437);
xnor U9057 (N_9057,N_8731,N_8488);
xnor U9058 (N_9058,N_8348,N_8878);
nand U9059 (N_9059,N_8421,N_8542);
nand U9060 (N_9060,N_8243,N_8782);
nor U9061 (N_9061,N_8223,N_8551);
and U9062 (N_9062,N_8020,N_8707);
or U9063 (N_9063,N_8423,N_8978);
xor U9064 (N_9064,N_8072,N_8110);
nor U9065 (N_9065,N_8643,N_8798);
or U9066 (N_9066,N_8828,N_8597);
nor U9067 (N_9067,N_8008,N_8890);
and U9068 (N_9068,N_8685,N_8458);
or U9069 (N_9069,N_8066,N_8553);
nand U9070 (N_9070,N_8199,N_8550);
xnor U9071 (N_9071,N_8354,N_8334);
and U9072 (N_9072,N_8864,N_8776);
nor U9073 (N_9073,N_8888,N_8797);
or U9074 (N_9074,N_8062,N_8709);
and U9075 (N_9075,N_8140,N_8121);
nor U9076 (N_9076,N_8701,N_8834);
nand U9077 (N_9077,N_8104,N_8206);
xnor U9078 (N_9078,N_8357,N_8813);
or U9079 (N_9079,N_8254,N_8208);
nor U9080 (N_9080,N_8788,N_8069);
nand U9081 (N_9081,N_8001,N_8483);
xor U9082 (N_9082,N_8341,N_8291);
nand U9083 (N_9083,N_8297,N_8559);
and U9084 (N_9084,N_8419,N_8149);
nand U9085 (N_9085,N_8303,N_8496);
nand U9086 (N_9086,N_8146,N_8887);
nor U9087 (N_9087,N_8764,N_8520);
or U9088 (N_9088,N_8921,N_8668);
nand U9089 (N_9089,N_8239,N_8157);
xor U9090 (N_9090,N_8638,N_8954);
and U9091 (N_9091,N_8089,N_8085);
and U9092 (N_9092,N_8424,N_8077);
nor U9093 (N_9093,N_8466,N_8296);
nand U9094 (N_9094,N_8889,N_8736);
nor U9095 (N_9095,N_8109,N_8343);
nand U9096 (N_9096,N_8628,N_8368);
or U9097 (N_9097,N_8960,N_8529);
and U9098 (N_9098,N_8926,N_8826);
xnor U9099 (N_9099,N_8829,N_8599);
xor U9100 (N_9100,N_8572,N_8142);
or U9101 (N_9101,N_8474,N_8703);
and U9102 (N_9102,N_8927,N_8169);
xor U9103 (N_9103,N_8189,N_8699);
or U9104 (N_9104,N_8323,N_8795);
or U9105 (N_9105,N_8601,N_8747);
nand U9106 (N_9106,N_8482,N_8715);
and U9107 (N_9107,N_8970,N_8151);
or U9108 (N_9108,N_8886,N_8574);
and U9109 (N_9109,N_8955,N_8958);
and U9110 (N_9110,N_8002,N_8913);
and U9111 (N_9111,N_8857,N_8118);
or U9112 (N_9112,N_8019,N_8552);
nor U9113 (N_9113,N_8783,N_8630);
nand U9114 (N_9114,N_8076,N_8037);
nor U9115 (N_9115,N_8875,N_8016);
nand U9116 (N_9116,N_8900,N_8847);
xnor U9117 (N_9117,N_8344,N_8375);
and U9118 (N_9118,N_8238,N_8578);
xor U9119 (N_9119,N_8227,N_8675);
xnor U9120 (N_9120,N_8723,N_8674);
nand U9121 (N_9121,N_8162,N_8617);
nand U9122 (N_9122,N_8061,N_8382);
and U9123 (N_9123,N_8017,N_8155);
or U9124 (N_9124,N_8535,N_8274);
xor U9125 (N_9125,N_8464,N_8204);
or U9126 (N_9126,N_8439,N_8745);
xor U9127 (N_9127,N_8141,N_8667);
nor U9128 (N_9128,N_8187,N_8841);
or U9129 (N_9129,N_8613,N_8388);
or U9130 (N_9130,N_8372,N_8655);
or U9131 (N_9131,N_8241,N_8262);
nor U9132 (N_9132,N_8659,N_8778);
xor U9133 (N_9133,N_8676,N_8988);
nand U9134 (N_9134,N_8404,N_8105);
xnor U9135 (N_9135,N_8846,N_8758);
nand U9136 (N_9136,N_8839,N_8734);
or U9137 (N_9137,N_8179,N_8907);
xor U9138 (N_9138,N_8218,N_8205);
or U9139 (N_9139,N_8825,N_8221);
nor U9140 (N_9140,N_8318,N_8898);
and U9141 (N_9141,N_8048,N_8827);
or U9142 (N_9142,N_8370,N_8175);
xnor U9143 (N_9143,N_8702,N_8527);
xor U9144 (N_9144,N_8147,N_8051);
nand U9145 (N_9145,N_8097,N_8081);
or U9146 (N_9146,N_8268,N_8363);
nor U9147 (N_9147,N_8906,N_8603);
xnor U9148 (N_9148,N_8405,N_8891);
xor U9149 (N_9149,N_8038,N_8159);
xnor U9150 (N_9150,N_8126,N_8090);
xor U9151 (N_9151,N_8411,N_8261);
and U9152 (N_9152,N_8315,N_8237);
or U9153 (N_9153,N_8884,N_8079);
xor U9154 (N_9154,N_8696,N_8943);
xor U9155 (N_9155,N_8852,N_8418);
nand U9156 (N_9156,N_8903,N_8133);
xor U9157 (N_9157,N_8649,N_8508);
xor U9158 (N_9158,N_8108,N_8058);
nor U9159 (N_9159,N_8904,N_8285);
nand U9160 (N_9160,N_8420,N_8456);
nand U9161 (N_9161,N_8755,N_8815);
nand U9162 (N_9162,N_8014,N_8230);
nor U9163 (N_9163,N_8650,N_8623);
nor U9164 (N_9164,N_8768,N_8682);
xor U9165 (N_9165,N_8789,N_8346);
or U9166 (N_9166,N_8821,N_8272);
and U9167 (N_9167,N_8180,N_8743);
xnor U9168 (N_9168,N_8120,N_8447);
and U9169 (N_9169,N_8662,N_8403);
xnor U9170 (N_9170,N_8331,N_8358);
xnor U9171 (N_9171,N_8928,N_8722);
xnor U9172 (N_9172,N_8931,N_8573);
and U9173 (N_9173,N_8495,N_8994);
nand U9174 (N_9174,N_8507,N_8693);
nand U9175 (N_9175,N_8521,N_8705);
xnor U9176 (N_9176,N_8996,N_8417);
or U9177 (N_9177,N_8164,N_8381);
xnor U9178 (N_9178,N_8373,N_8610);
nor U9179 (N_9179,N_8746,N_8248);
nand U9180 (N_9180,N_8637,N_8644);
nor U9181 (N_9181,N_8202,N_8930);
nor U9182 (N_9182,N_8983,N_8629);
and U9183 (N_9183,N_8356,N_8391);
nor U9184 (N_9184,N_8332,N_8934);
xor U9185 (N_9185,N_8673,N_8490);
xor U9186 (N_9186,N_8690,N_8964);
xnor U9187 (N_9187,N_8760,N_8099);
xor U9188 (N_9188,N_8152,N_8479);
or U9189 (N_9189,N_8432,N_8213);
or U9190 (N_9190,N_8459,N_8176);
nor U9191 (N_9191,N_8716,N_8987);
or U9192 (N_9192,N_8582,N_8605);
or U9193 (N_9193,N_8489,N_8124);
or U9194 (N_9194,N_8294,N_8992);
nor U9195 (N_9195,N_8013,N_8880);
xor U9196 (N_9196,N_8499,N_8883);
nand U9197 (N_9197,N_8035,N_8531);
xnor U9198 (N_9198,N_8896,N_8113);
xnor U9199 (N_9199,N_8135,N_8103);
nor U9200 (N_9200,N_8895,N_8519);
nand U9201 (N_9201,N_8044,N_8328);
or U9202 (N_9202,N_8807,N_8950);
or U9203 (N_9203,N_8565,N_8953);
or U9204 (N_9204,N_8589,N_8756);
xnor U9205 (N_9205,N_8145,N_8280);
xor U9206 (N_9206,N_8774,N_8339);
nor U9207 (N_9207,N_8590,N_8652);
or U9208 (N_9208,N_8029,N_8452);
and U9209 (N_9209,N_8377,N_8881);
nand U9210 (N_9210,N_8564,N_8338);
or U9211 (N_9211,N_8800,N_8446);
nand U9212 (N_9212,N_8185,N_8567);
or U9213 (N_9213,N_8704,N_8033);
and U9214 (N_9214,N_8049,N_8448);
and U9215 (N_9215,N_8426,N_8050);
nand U9216 (N_9216,N_8376,N_8409);
nor U9217 (N_9217,N_8608,N_8476);
and U9218 (N_9218,N_8487,N_8095);
or U9219 (N_9219,N_8053,N_8413);
xnor U9220 (N_9220,N_8198,N_8604);
xnor U9221 (N_9221,N_8860,N_8047);
and U9222 (N_9222,N_8912,N_8143);
or U9223 (N_9223,N_8647,N_8538);
and U9224 (N_9224,N_8326,N_8752);
nand U9225 (N_9225,N_8870,N_8136);
nor U9226 (N_9226,N_8270,N_8009);
and U9227 (N_9227,N_8390,N_8689);
nand U9228 (N_9228,N_8127,N_8654);
or U9229 (N_9229,N_8727,N_8161);
and U9230 (N_9230,N_8319,N_8299);
nand U9231 (N_9231,N_8024,N_8060);
nor U9232 (N_9232,N_8871,N_8710);
and U9233 (N_9233,N_8036,N_8730);
or U9234 (N_9234,N_8657,N_8342);
or U9235 (N_9235,N_8571,N_8465);
and U9236 (N_9236,N_8570,N_8767);
xnor U9237 (N_9237,N_8949,N_8516);
xnor U9238 (N_9238,N_8335,N_8639);
or U9239 (N_9239,N_8919,N_8796);
nor U9240 (N_9240,N_8394,N_8641);
nor U9241 (N_9241,N_8023,N_8098);
or U9242 (N_9242,N_8168,N_8330);
and U9243 (N_9243,N_8384,N_8816);
nand U9244 (N_9244,N_8719,N_8380);
nand U9245 (N_9245,N_8977,N_8810);
nor U9246 (N_9246,N_8043,N_8428);
and U9247 (N_9247,N_8946,N_8144);
nand U9248 (N_9248,N_8620,N_8026);
nand U9249 (N_9249,N_8004,N_8347);
and U9250 (N_9250,N_8739,N_8733);
and U9251 (N_9251,N_8304,N_8378);
xor U9252 (N_9252,N_8430,N_8300);
or U9253 (N_9253,N_8728,N_8985);
nor U9254 (N_9254,N_8713,N_8324);
and U9255 (N_9255,N_8267,N_8306);
or U9256 (N_9256,N_8400,N_8498);
nor U9257 (N_9257,N_8809,N_8307);
and U9258 (N_9258,N_8259,N_8100);
and U9259 (N_9259,N_8305,N_8515);
and U9260 (N_9260,N_8525,N_8389);
nor U9261 (N_9261,N_8678,N_8735);
nand U9262 (N_9262,N_8595,N_8818);
and U9263 (N_9263,N_8472,N_8271);
and U9264 (N_9264,N_8225,N_8969);
nand U9265 (N_9265,N_8242,N_8648);
nor U9266 (N_9266,N_8741,N_8308);
and U9267 (N_9267,N_8406,N_8577);
or U9268 (N_9268,N_8138,N_8961);
xnor U9269 (N_9269,N_8027,N_8065);
or U9270 (N_9270,N_8700,N_8777);
or U9271 (N_9271,N_8369,N_8264);
and U9272 (N_9272,N_8967,N_8708);
and U9273 (N_9273,N_8956,N_8683);
nand U9274 (N_9274,N_8740,N_8951);
and U9275 (N_9275,N_8467,N_8687);
and U9276 (N_9276,N_8284,N_8633);
and U9277 (N_9277,N_8514,N_8790);
nor U9278 (N_9278,N_8500,N_8131);
nor U9279 (N_9279,N_8313,N_8509);
nor U9280 (N_9280,N_8836,N_8606);
nor U9281 (N_9281,N_8444,N_8814);
and U9282 (N_9282,N_8286,N_8056);
xnor U9283 (N_9283,N_8367,N_8032);
nor U9284 (N_9284,N_8902,N_8779);
nand U9285 (N_9285,N_8653,N_8167);
and U9286 (N_9286,N_8897,N_8576);
or U9287 (N_9287,N_8822,N_8692);
nand U9288 (N_9288,N_8503,N_8207);
nand U9289 (N_9289,N_8671,N_8882);
or U9290 (N_9290,N_8030,N_8805);
xnor U9291 (N_9291,N_8018,N_8183);
and U9292 (N_9292,N_8402,N_8720);
nor U9293 (N_9293,N_8909,N_8753);
and U9294 (N_9294,N_8959,N_8084);
nor U9295 (N_9295,N_8115,N_8288);
xor U9296 (N_9296,N_8477,N_8366);
and U9297 (N_9297,N_8669,N_8282);
and U9298 (N_9298,N_8759,N_8194);
nand U9299 (N_9299,N_8915,N_8794);
nor U9300 (N_9300,N_8566,N_8658);
and U9301 (N_9301,N_8554,N_8114);
or U9302 (N_9302,N_8712,N_8598);
nand U9303 (N_9303,N_8594,N_8484);
xor U9304 (N_9304,N_8433,N_8894);
xnor U9305 (N_9305,N_8359,N_8632);
and U9306 (N_9306,N_8224,N_8000);
or U9307 (N_9307,N_8501,N_8635);
and U9308 (N_9308,N_8436,N_8340);
or U9309 (N_9309,N_8449,N_8737);
xor U9310 (N_9310,N_8711,N_8833);
xnor U9311 (N_9311,N_8532,N_8276);
xor U9312 (N_9312,N_8247,N_8217);
or U9313 (N_9313,N_8924,N_8851);
xor U9314 (N_9314,N_8945,N_8111);
and U9315 (N_9315,N_8320,N_8455);
xor U9316 (N_9316,N_8989,N_8602);
and U9317 (N_9317,N_8670,N_8510);
nand U9318 (N_9318,N_8511,N_8694);
nand U9319 (N_9319,N_8491,N_8627);
nand U9320 (N_9320,N_8150,N_8780);
nand U9321 (N_9321,N_8770,N_8748);
nor U9322 (N_9322,N_8252,N_8492);
and U9323 (N_9323,N_8544,N_8517);
or U9324 (N_9324,N_8824,N_8993);
or U9325 (N_9325,N_8512,N_8998);
nor U9326 (N_9326,N_8942,N_8485);
xor U9327 (N_9327,N_8080,N_8697);
nor U9328 (N_9328,N_8539,N_8568);
nand U9329 (N_9329,N_8309,N_8434);
nand U9330 (N_9330,N_8787,N_8840);
and U9331 (N_9331,N_8278,N_8025);
and U9332 (N_9332,N_8817,N_8679);
xor U9333 (N_9333,N_8385,N_8325);
xnor U9334 (N_9334,N_8616,N_8277);
or U9335 (N_9335,N_8656,N_8792);
xor U9336 (N_9336,N_8624,N_8526);
or U9337 (N_9337,N_8349,N_8995);
and U9338 (N_9338,N_8914,N_8178);
or U9339 (N_9339,N_8929,N_8588);
or U9340 (N_9340,N_8321,N_8414);
nand U9341 (N_9341,N_8773,N_8717);
nor U9342 (N_9342,N_8087,N_8327);
and U9343 (N_9343,N_8130,N_8876);
nand U9344 (N_9344,N_8469,N_8010);
nand U9345 (N_9345,N_8845,N_8457);
nor U9346 (N_9346,N_8663,N_8106);
nor U9347 (N_9347,N_8830,N_8462);
nand U9348 (N_9348,N_8337,N_8122);
nand U9349 (N_9349,N_8052,N_8137);
xor U9350 (N_9350,N_8083,N_8148);
or U9351 (N_9351,N_8078,N_8965);
nor U9352 (N_9352,N_8494,N_8171);
nor U9353 (N_9353,N_8255,N_8732);
nor U9354 (N_9354,N_8011,N_8856);
nand U9355 (N_9355,N_8849,N_8258);
xnor U9356 (N_9356,N_8651,N_8063);
xnor U9357 (N_9357,N_8772,N_8173);
nand U9358 (N_9358,N_8948,N_8398);
nor U9359 (N_9359,N_8972,N_8353);
xor U9360 (N_9360,N_8139,N_8226);
and U9361 (N_9361,N_8569,N_8540);
nor U9362 (N_9362,N_8600,N_8631);
nand U9363 (N_9363,N_8028,N_8831);
xnor U9364 (N_9364,N_8762,N_8253);
and U9365 (N_9365,N_8980,N_8212);
xor U9366 (N_9366,N_8005,N_8265);
nand U9367 (N_9367,N_8698,N_8441);
nor U9368 (N_9368,N_8619,N_8917);
and U9369 (N_9369,N_8435,N_8592);
and U9370 (N_9370,N_8665,N_8231);
xor U9371 (N_9371,N_8399,N_8607);
and U9372 (N_9372,N_8916,N_8680);
nor U9373 (N_9373,N_8811,N_8843);
nand U9374 (N_9374,N_8283,N_8666);
nor U9375 (N_9375,N_8952,N_8611);
nor U9376 (N_9376,N_8505,N_8726);
xnor U9377 (N_9377,N_8094,N_8160);
or U9378 (N_9378,N_8345,N_8473);
or U9379 (N_9379,N_8287,N_8855);
or U9380 (N_9380,N_8200,N_8935);
xor U9381 (N_9381,N_8636,N_8556);
and U9382 (N_9382,N_8064,N_8034);
or U9383 (N_9383,N_8986,N_8260);
xnor U9384 (N_9384,N_8196,N_8555);
or U9385 (N_9385,N_8806,N_8006);
nand U9386 (N_9386,N_8351,N_8761);
xor U9387 (N_9387,N_8233,N_8744);
nor U9388 (N_9388,N_8944,N_8999);
nand U9389 (N_9389,N_8749,N_8686);
and U9390 (N_9390,N_8119,N_8425);
nor U9391 (N_9391,N_8549,N_8548);
or U9392 (N_9392,N_8387,N_8672);
nand U9393 (N_9393,N_8275,N_8738);
nand U9394 (N_9394,N_8664,N_8250);
and U9395 (N_9395,N_8976,N_8892);
xnor U9396 (N_9396,N_8766,N_8725);
xor U9397 (N_9397,N_8963,N_8979);
or U9398 (N_9398,N_8893,N_8393);
nand U9399 (N_9399,N_8751,N_8416);
or U9400 (N_9400,N_8071,N_8862);
xor U9401 (N_9401,N_8781,N_8518);
nand U9402 (N_9402,N_8932,N_8706);
nor U9403 (N_9403,N_8771,N_8156);
or U9404 (N_9404,N_8724,N_8182);
or U9405 (N_9405,N_8645,N_8188);
and U9406 (N_9406,N_8475,N_8869);
xor U9407 (N_9407,N_8868,N_8848);
nor U9408 (N_9408,N_8925,N_8534);
and U9409 (N_9409,N_8203,N_8301);
nand U9410 (N_9410,N_8181,N_8445);
nand U9411 (N_9411,N_8386,N_8547);
and U9412 (N_9412,N_8471,N_8593);
nand U9413 (N_9413,N_8506,N_8634);
nand U9414 (N_9414,N_8799,N_8622);
and U9415 (N_9415,N_8407,N_8640);
or U9416 (N_9416,N_8046,N_8513);
xor U9417 (N_9417,N_8804,N_8625);
xor U9418 (N_9418,N_8172,N_8872);
nand U9419 (N_9419,N_8229,N_8191);
xor U9420 (N_9420,N_8219,N_8863);
nand U9421 (N_9421,N_8316,N_8129);
and U9422 (N_9422,N_8584,N_8901);
and U9423 (N_9423,N_8102,N_8546);
nand U9424 (N_9424,N_8174,N_8587);
nand U9425 (N_9425,N_8396,N_8163);
xor U9426 (N_9426,N_8302,N_8585);
nand U9427 (N_9427,N_8677,N_8750);
nand U9428 (N_9428,N_8802,N_8088);
xnor U9429 (N_9429,N_8523,N_8170);
nand U9430 (N_9430,N_8123,N_8201);
and U9431 (N_9431,N_8543,N_8045);
nor U9432 (N_9432,N_8468,N_8310);
nand U9433 (N_9433,N_8478,N_8463);
xnor U9434 (N_9434,N_8688,N_8729);
nor U9435 (N_9435,N_8661,N_8215);
and U9436 (N_9436,N_8222,N_8355);
nand U9437 (N_9437,N_8560,N_8450);
or U9438 (N_9438,N_8154,N_8093);
nand U9439 (N_9439,N_8438,N_8691);
xnor U9440 (N_9440,N_8480,N_8317);
nand U9441 (N_9441,N_8528,N_8838);
or U9442 (N_9442,N_8412,N_8545);
nor U9443 (N_9443,N_8885,N_8365);
xor U9444 (N_9444,N_8615,N_8957);
xor U9445 (N_9445,N_8442,N_8803);
nor U9446 (N_9446,N_8660,N_8214);
nor U9447 (N_9447,N_8754,N_8039);
nor U9448 (N_9448,N_8251,N_8557);
and U9449 (N_9449,N_8470,N_8867);
or U9450 (N_9450,N_8091,N_8451);
nor U9451 (N_9451,N_8232,N_8116);
nor U9452 (N_9452,N_8249,N_8015);
nor U9453 (N_9453,N_8975,N_8295);
and U9454 (N_9454,N_8524,N_8842);
nor U9455 (N_9455,N_8311,N_8246);
nand U9456 (N_9456,N_8910,N_8791);
xnor U9457 (N_9457,N_8879,N_8021);
nor U9458 (N_9458,N_8054,N_8626);
nor U9459 (N_9459,N_8695,N_8812);
or U9460 (N_9460,N_8922,N_8968);
nor U9461 (N_9461,N_8042,N_8236);
or U9462 (N_9462,N_8502,N_8235);
nor U9463 (N_9463,N_8763,N_8379);
nand U9464 (N_9464,N_8793,N_8190);
or U9465 (N_9465,N_8832,N_8920);
nor U9466 (N_9466,N_8579,N_8861);
xnor U9467 (N_9467,N_8041,N_8290);
xor U9468 (N_9468,N_8022,N_8984);
or U9469 (N_9469,N_8134,N_8939);
nand U9470 (N_9470,N_8336,N_8415);
nand U9471 (N_9471,N_8580,N_8854);
and U9472 (N_9472,N_8769,N_8040);
nand U9473 (N_9473,N_8786,N_8289);
xor U9474 (N_9474,N_8211,N_8908);
nand U9475 (N_9475,N_8933,N_8165);
and U9476 (N_9476,N_8561,N_8497);
and U9477 (N_9477,N_8614,N_8209);
nor U9478 (N_9478,N_8440,N_8007);
xnor U9479 (N_9479,N_8059,N_8785);
nand U9480 (N_9480,N_8461,N_8361);
nand U9481 (N_9481,N_8837,N_8941);
nor U9482 (N_9482,N_8681,N_8112);
or U9483 (N_9483,N_8153,N_8273);
or U9484 (N_9484,N_8823,N_8086);
xnor U9485 (N_9485,N_8266,N_8362);
xnor U9486 (N_9486,N_8858,N_8575);
nand U9487 (N_9487,N_8591,N_8997);
xor U9488 (N_9488,N_8757,N_8293);
or U9489 (N_9489,N_8905,N_8481);
nand U9490 (N_9490,N_8197,N_8493);
nand U9491 (N_9491,N_8820,N_8101);
or U9492 (N_9492,N_8057,N_8460);
and U9493 (N_9493,N_8070,N_8096);
xnor U9494 (N_9494,N_8427,N_8877);
nor U9495 (N_9495,N_8940,N_8981);
nor U9496 (N_9496,N_8184,N_8234);
xnor U9497 (N_9497,N_8583,N_8966);
or U9498 (N_9498,N_8360,N_8504);
and U9499 (N_9499,N_8220,N_8329);
nand U9500 (N_9500,N_8966,N_8147);
xor U9501 (N_9501,N_8710,N_8899);
xnor U9502 (N_9502,N_8476,N_8531);
or U9503 (N_9503,N_8323,N_8892);
or U9504 (N_9504,N_8177,N_8901);
and U9505 (N_9505,N_8063,N_8779);
or U9506 (N_9506,N_8541,N_8283);
nor U9507 (N_9507,N_8430,N_8525);
xor U9508 (N_9508,N_8301,N_8580);
xnor U9509 (N_9509,N_8737,N_8531);
and U9510 (N_9510,N_8059,N_8651);
and U9511 (N_9511,N_8038,N_8128);
nor U9512 (N_9512,N_8390,N_8625);
and U9513 (N_9513,N_8888,N_8569);
or U9514 (N_9514,N_8934,N_8022);
and U9515 (N_9515,N_8453,N_8163);
xnor U9516 (N_9516,N_8141,N_8110);
and U9517 (N_9517,N_8160,N_8487);
xnor U9518 (N_9518,N_8691,N_8465);
xnor U9519 (N_9519,N_8778,N_8998);
nand U9520 (N_9520,N_8037,N_8562);
xnor U9521 (N_9521,N_8843,N_8201);
and U9522 (N_9522,N_8382,N_8218);
xor U9523 (N_9523,N_8629,N_8315);
nor U9524 (N_9524,N_8764,N_8318);
nand U9525 (N_9525,N_8870,N_8647);
xor U9526 (N_9526,N_8416,N_8476);
nor U9527 (N_9527,N_8050,N_8678);
xor U9528 (N_9528,N_8728,N_8276);
nor U9529 (N_9529,N_8493,N_8247);
nand U9530 (N_9530,N_8282,N_8368);
xnor U9531 (N_9531,N_8267,N_8399);
or U9532 (N_9532,N_8606,N_8380);
xnor U9533 (N_9533,N_8194,N_8349);
nor U9534 (N_9534,N_8925,N_8176);
or U9535 (N_9535,N_8528,N_8154);
nand U9536 (N_9536,N_8603,N_8260);
nand U9537 (N_9537,N_8335,N_8667);
and U9538 (N_9538,N_8221,N_8199);
or U9539 (N_9539,N_8929,N_8253);
or U9540 (N_9540,N_8661,N_8549);
nand U9541 (N_9541,N_8746,N_8174);
or U9542 (N_9542,N_8602,N_8425);
xor U9543 (N_9543,N_8293,N_8474);
xor U9544 (N_9544,N_8839,N_8234);
and U9545 (N_9545,N_8063,N_8409);
nand U9546 (N_9546,N_8798,N_8262);
or U9547 (N_9547,N_8056,N_8322);
nand U9548 (N_9548,N_8627,N_8007);
and U9549 (N_9549,N_8276,N_8655);
xor U9550 (N_9550,N_8229,N_8877);
nor U9551 (N_9551,N_8607,N_8363);
nand U9552 (N_9552,N_8866,N_8432);
nand U9553 (N_9553,N_8007,N_8108);
and U9554 (N_9554,N_8395,N_8107);
or U9555 (N_9555,N_8703,N_8335);
and U9556 (N_9556,N_8727,N_8647);
or U9557 (N_9557,N_8014,N_8250);
xnor U9558 (N_9558,N_8653,N_8929);
nand U9559 (N_9559,N_8624,N_8398);
nand U9560 (N_9560,N_8080,N_8776);
xnor U9561 (N_9561,N_8881,N_8201);
nor U9562 (N_9562,N_8424,N_8173);
and U9563 (N_9563,N_8991,N_8772);
nor U9564 (N_9564,N_8767,N_8827);
nand U9565 (N_9565,N_8440,N_8609);
nand U9566 (N_9566,N_8960,N_8775);
nor U9567 (N_9567,N_8358,N_8550);
xnor U9568 (N_9568,N_8946,N_8129);
or U9569 (N_9569,N_8611,N_8319);
nand U9570 (N_9570,N_8717,N_8048);
and U9571 (N_9571,N_8623,N_8078);
nand U9572 (N_9572,N_8925,N_8460);
nor U9573 (N_9573,N_8104,N_8168);
or U9574 (N_9574,N_8690,N_8939);
and U9575 (N_9575,N_8811,N_8488);
nand U9576 (N_9576,N_8039,N_8898);
nand U9577 (N_9577,N_8440,N_8407);
and U9578 (N_9578,N_8829,N_8637);
nand U9579 (N_9579,N_8522,N_8605);
or U9580 (N_9580,N_8202,N_8225);
nor U9581 (N_9581,N_8727,N_8331);
or U9582 (N_9582,N_8746,N_8665);
xnor U9583 (N_9583,N_8425,N_8434);
nor U9584 (N_9584,N_8323,N_8746);
or U9585 (N_9585,N_8024,N_8260);
xor U9586 (N_9586,N_8672,N_8241);
and U9587 (N_9587,N_8061,N_8658);
xnor U9588 (N_9588,N_8022,N_8571);
and U9589 (N_9589,N_8214,N_8551);
and U9590 (N_9590,N_8883,N_8740);
xor U9591 (N_9591,N_8860,N_8947);
nor U9592 (N_9592,N_8854,N_8695);
or U9593 (N_9593,N_8592,N_8785);
and U9594 (N_9594,N_8030,N_8270);
nand U9595 (N_9595,N_8181,N_8311);
nand U9596 (N_9596,N_8136,N_8763);
and U9597 (N_9597,N_8668,N_8587);
nand U9598 (N_9598,N_8553,N_8536);
nor U9599 (N_9599,N_8684,N_8097);
xnor U9600 (N_9600,N_8421,N_8311);
xor U9601 (N_9601,N_8253,N_8083);
nor U9602 (N_9602,N_8003,N_8021);
or U9603 (N_9603,N_8367,N_8293);
nand U9604 (N_9604,N_8085,N_8306);
xnor U9605 (N_9605,N_8919,N_8752);
and U9606 (N_9606,N_8771,N_8150);
and U9607 (N_9607,N_8513,N_8663);
or U9608 (N_9608,N_8527,N_8218);
or U9609 (N_9609,N_8261,N_8626);
and U9610 (N_9610,N_8024,N_8328);
xor U9611 (N_9611,N_8533,N_8509);
and U9612 (N_9612,N_8966,N_8537);
xor U9613 (N_9613,N_8427,N_8560);
and U9614 (N_9614,N_8079,N_8465);
or U9615 (N_9615,N_8687,N_8918);
nor U9616 (N_9616,N_8932,N_8553);
xnor U9617 (N_9617,N_8396,N_8921);
nor U9618 (N_9618,N_8012,N_8984);
and U9619 (N_9619,N_8569,N_8022);
and U9620 (N_9620,N_8452,N_8872);
nor U9621 (N_9621,N_8351,N_8746);
xor U9622 (N_9622,N_8651,N_8832);
nor U9623 (N_9623,N_8312,N_8462);
nor U9624 (N_9624,N_8771,N_8300);
or U9625 (N_9625,N_8174,N_8629);
and U9626 (N_9626,N_8328,N_8810);
nor U9627 (N_9627,N_8566,N_8678);
xnor U9628 (N_9628,N_8320,N_8764);
nor U9629 (N_9629,N_8303,N_8129);
and U9630 (N_9630,N_8051,N_8371);
or U9631 (N_9631,N_8123,N_8046);
nor U9632 (N_9632,N_8748,N_8603);
and U9633 (N_9633,N_8506,N_8083);
or U9634 (N_9634,N_8938,N_8733);
nor U9635 (N_9635,N_8362,N_8094);
nor U9636 (N_9636,N_8181,N_8280);
nor U9637 (N_9637,N_8376,N_8245);
nand U9638 (N_9638,N_8520,N_8602);
nand U9639 (N_9639,N_8538,N_8377);
nor U9640 (N_9640,N_8341,N_8210);
xor U9641 (N_9641,N_8504,N_8896);
nor U9642 (N_9642,N_8506,N_8776);
nand U9643 (N_9643,N_8605,N_8303);
and U9644 (N_9644,N_8307,N_8841);
or U9645 (N_9645,N_8746,N_8941);
or U9646 (N_9646,N_8004,N_8304);
nand U9647 (N_9647,N_8794,N_8693);
nor U9648 (N_9648,N_8952,N_8259);
xnor U9649 (N_9649,N_8450,N_8627);
nand U9650 (N_9650,N_8267,N_8798);
xnor U9651 (N_9651,N_8279,N_8215);
and U9652 (N_9652,N_8141,N_8550);
xnor U9653 (N_9653,N_8772,N_8300);
or U9654 (N_9654,N_8337,N_8020);
xor U9655 (N_9655,N_8045,N_8517);
nand U9656 (N_9656,N_8189,N_8385);
nor U9657 (N_9657,N_8424,N_8529);
or U9658 (N_9658,N_8222,N_8234);
or U9659 (N_9659,N_8336,N_8159);
or U9660 (N_9660,N_8154,N_8660);
nor U9661 (N_9661,N_8148,N_8816);
nand U9662 (N_9662,N_8929,N_8397);
nand U9663 (N_9663,N_8089,N_8688);
nor U9664 (N_9664,N_8910,N_8295);
nand U9665 (N_9665,N_8534,N_8458);
xnor U9666 (N_9666,N_8990,N_8108);
and U9667 (N_9667,N_8310,N_8789);
or U9668 (N_9668,N_8240,N_8079);
or U9669 (N_9669,N_8786,N_8705);
nand U9670 (N_9670,N_8613,N_8132);
xnor U9671 (N_9671,N_8465,N_8243);
nand U9672 (N_9672,N_8534,N_8463);
nand U9673 (N_9673,N_8909,N_8873);
or U9674 (N_9674,N_8773,N_8029);
xnor U9675 (N_9675,N_8723,N_8285);
or U9676 (N_9676,N_8133,N_8274);
nor U9677 (N_9677,N_8498,N_8430);
nand U9678 (N_9678,N_8966,N_8336);
and U9679 (N_9679,N_8755,N_8319);
nand U9680 (N_9680,N_8137,N_8183);
xor U9681 (N_9681,N_8816,N_8011);
nand U9682 (N_9682,N_8053,N_8356);
or U9683 (N_9683,N_8979,N_8207);
nand U9684 (N_9684,N_8246,N_8890);
and U9685 (N_9685,N_8951,N_8308);
xnor U9686 (N_9686,N_8918,N_8370);
nor U9687 (N_9687,N_8843,N_8978);
nand U9688 (N_9688,N_8437,N_8329);
xnor U9689 (N_9689,N_8557,N_8670);
nor U9690 (N_9690,N_8065,N_8859);
or U9691 (N_9691,N_8464,N_8708);
or U9692 (N_9692,N_8583,N_8515);
or U9693 (N_9693,N_8948,N_8405);
and U9694 (N_9694,N_8296,N_8352);
nand U9695 (N_9695,N_8939,N_8132);
nand U9696 (N_9696,N_8440,N_8848);
and U9697 (N_9697,N_8176,N_8516);
xor U9698 (N_9698,N_8978,N_8219);
nor U9699 (N_9699,N_8542,N_8032);
nand U9700 (N_9700,N_8133,N_8650);
and U9701 (N_9701,N_8758,N_8282);
xor U9702 (N_9702,N_8158,N_8134);
nand U9703 (N_9703,N_8828,N_8376);
or U9704 (N_9704,N_8143,N_8524);
or U9705 (N_9705,N_8028,N_8745);
or U9706 (N_9706,N_8584,N_8242);
xnor U9707 (N_9707,N_8360,N_8412);
nand U9708 (N_9708,N_8077,N_8120);
and U9709 (N_9709,N_8463,N_8826);
and U9710 (N_9710,N_8154,N_8423);
or U9711 (N_9711,N_8015,N_8652);
nor U9712 (N_9712,N_8315,N_8997);
and U9713 (N_9713,N_8730,N_8381);
nor U9714 (N_9714,N_8408,N_8596);
xor U9715 (N_9715,N_8158,N_8297);
and U9716 (N_9716,N_8756,N_8276);
or U9717 (N_9717,N_8119,N_8975);
nor U9718 (N_9718,N_8286,N_8915);
and U9719 (N_9719,N_8711,N_8415);
or U9720 (N_9720,N_8152,N_8419);
nand U9721 (N_9721,N_8619,N_8492);
nor U9722 (N_9722,N_8796,N_8070);
nand U9723 (N_9723,N_8843,N_8862);
nor U9724 (N_9724,N_8654,N_8006);
nand U9725 (N_9725,N_8609,N_8322);
xnor U9726 (N_9726,N_8513,N_8826);
nand U9727 (N_9727,N_8400,N_8027);
or U9728 (N_9728,N_8093,N_8715);
nor U9729 (N_9729,N_8427,N_8207);
nor U9730 (N_9730,N_8585,N_8415);
and U9731 (N_9731,N_8863,N_8039);
or U9732 (N_9732,N_8696,N_8239);
or U9733 (N_9733,N_8344,N_8204);
or U9734 (N_9734,N_8345,N_8445);
nor U9735 (N_9735,N_8950,N_8028);
nor U9736 (N_9736,N_8070,N_8346);
or U9737 (N_9737,N_8898,N_8174);
xnor U9738 (N_9738,N_8394,N_8263);
and U9739 (N_9739,N_8338,N_8536);
or U9740 (N_9740,N_8233,N_8445);
nor U9741 (N_9741,N_8349,N_8081);
and U9742 (N_9742,N_8460,N_8823);
nor U9743 (N_9743,N_8578,N_8620);
and U9744 (N_9744,N_8100,N_8931);
nor U9745 (N_9745,N_8660,N_8855);
and U9746 (N_9746,N_8308,N_8414);
xor U9747 (N_9747,N_8529,N_8098);
or U9748 (N_9748,N_8663,N_8849);
and U9749 (N_9749,N_8827,N_8499);
nand U9750 (N_9750,N_8669,N_8145);
xnor U9751 (N_9751,N_8585,N_8295);
nor U9752 (N_9752,N_8792,N_8694);
nand U9753 (N_9753,N_8961,N_8537);
and U9754 (N_9754,N_8285,N_8731);
or U9755 (N_9755,N_8211,N_8896);
nand U9756 (N_9756,N_8926,N_8217);
nand U9757 (N_9757,N_8804,N_8203);
or U9758 (N_9758,N_8489,N_8839);
or U9759 (N_9759,N_8557,N_8060);
nor U9760 (N_9760,N_8867,N_8993);
nand U9761 (N_9761,N_8444,N_8555);
xnor U9762 (N_9762,N_8600,N_8709);
xor U9763 (N_9763,N_8709,N_8264);
or U9764 (N_9764,N_8342,N_8464);
nand U9765 (N_9765,N_8264,N_8727);
and U9766 (N_9766,N_8188,N_8760);
or U9767 (N_9767,N_8129,N_8950);
or U9768 (N_9768,N_8605,N_8875);
or U9769 (N_9769,N_8134,N_8611);
nor U9770 (N_9770,N_8337,N_8487);
nor U9771 (N_9771,N_8621,N_8627);
xor U9772 (N_9772,N_8504,N_8665);
xnor U9773 (N_9773,N_8906,N_8432);
xnor U9774 (N_9774,N_8263,N_8086);
xor U9775 (N_9775,N_8308,N_8967);
xnor U9776 (N_9776,N_8511,N_8760);
nor U9777 (N_9777,N_8846,N_8397);
xor U9778 (N_9778,N_8759,N_8102);
or U9779 (N_9779,N_8630,N_8590);
nand U9780 (N_9780,N_8009,N_8656);
or U9781 (N_9781,N_8315,N_8394);
and U9782 (N_9782,N_8744,N_8373);
or U9783 (N_9783,N_8944,N_8640);
nand U9784 (N_9784,N_8035,N_8078);
nor U9785 (N_9785,N_8861,N_8648);
nor U9786 (N_9786,N_8052,N_8474);
or U9787 (N_9787,N_8432,N_8850);
and U9788 (N_9788,N_8370,N_8144);
nand U9789 (N_9789,N_8181,N_8541);
nor U9790 (N_9790,N_8116,N_8893);
nand U9791 (N_9791,N_8645,N_8198);
nand U9792 (N_9792,N_8527,N_8524);
and U9793 (N_9793,N_8355,N_8351);
and U9794 (N_9794,N_8355,N_8061);
and U9795 (N_9795,N_8684,N_8479);
nor U9796 (N_9796,N_8972,N_8357);
nor U9797 (N_9797,N_8054,N_8171);
and U9798 (N_9798,N_8720,N_8819);
and U9799 (N_9799,N_8871,N_8874);
nor U9800 (N_9800,N_8545,N_8535);
or U9801 (N_9801,N_8884,N_8880);
nor U9802 (N_9802,N_8952,N_8082);
xor U9803 (N_9803,N_8786,N_8374);
or U9804 (N_9804,N_8693,N_8045);
xor U9805 (N_9805,N_8680,N_8510);
xor U9806 (N_9806,N_8758,N_8054);
xnor U9807 (N_9807,N_8842,N_8513);
or U9808 (N_9808,N_8161,N_8900);
nor U9809 (N_9809,N_8865,N_8935);
nand U9810 (N_9810,N_8034,N_8928);
nand U9811 (N_9811,N_8314,N_8287);
and U9812 (N_9812,N_8743,N_8636);
nand U9813 (N_9813,N_8192,N_8776);
nor U9814 (N_9814,N_8576,N_8516);
and U9815 (N_9815,N_8276,N_8349);
xor U9816 (N_9816,N_8010,N_8942);
or U9817 (N_9817,N_8172,N_8126);
xnor U9818 (N_9818,N_8397,N_8598);
nor U9819 (N_9819,N_8345,N_8016);
and U9820 (N_9820,N_8429,N_8107);
or U9821 (N_9821,N_8515,N_8939);
xor U9822 (N_9822,N_8946,N_8475);
nand U9823 (N_9823,N_8283,N_8774);
nand U9824 (N_9824,N_8500,N_8998);
and U9825 (N_9825,N_8852,N_8495);
or U9826 (N_9826,N_8127,N_8930);
and U9827 (N_9827,N_8174,N_8828);
or U9828 (N_9828,N_8580,N_8544);
nor U9829 (N_9829,N_8216,N_8309);
nand U9830 (N_9830,N_8686,N_8595);
nor U9831 (N_9831,N_8499,N_8993);
nor U9832 (N_9832,N_8318,N_8423);
and U9833 (N_9833,N_8071,N_8438);
nand U9834 (N_9834,N_8983,N_8729);
and U9835 (N_9835,N_8829,N_8560);
nor U9836 (N_9836,N_8949,N_8487);
nor U9837 (N_9837,N_8228,N_8686);
nor U9838 (N_9838,N_8718,N_8101);
and U9839 (N_9839,N_8021,N_8274);
nand U9840 (N_9840,N_8695,N_8571);
or U9841 (N_9841,N_8852,N_8923);
nand U9842 (N_9842,N_8007,N_8211);
xor U9843 (N_9843,N_8875,N_8975);
xnor U9844 (N_9844,N_8708,N_8108);
and U9845 (N_9845,N_8159,N_8489);
and U9846 (N_9846,N_8602,N_8904);
or U9847 (N_9847,N_8513,N_8007);
xor U9848 (N_9848,N_8960,N_8176);
nand U9849 (N_9849,N_8050,N_8754);
and U9850 (N_9850,N_8286,N_8329);
xnor U9851 (N_9851,N_8149,N_8777);
xor U9852 (N_9852,N_8350,N_8977);
nand U9853 (N_9853,N_8877,N_8214);
nor U9854 (N_9854,N_8241,N_8447);
xnor U9855 (N_9855,N_8093,N_8265);
nand U9856 (N_9856,N_8670,N_8506);
xor U9857 (N_9857,N_8963,N_8271);
or U9858 (N_9858,N_8323,N_8685);
xnor U9859 (N_9859,N_8371,N_8171);
or U9860 (N_9860,N_8630,N_8785);
xor U9861 (N_9861,N_8850,N_8881);
and U9862 (N_9862,N_8412,N_8322);
nand U9863 (N_9863,N_8517,N_8672);
and U9864 (N_9864,N_8417,N_8944);
and U9865 (N_9865,N_8635,N_8244);
nand U9866 (N_9866,N_8264,N_8723);
nand U9867 (N_9867,N_8660,N_8810);
nand U9868 (N_9868,N_8710,N_8542);
xor U9869 (N_9869,N_8259,N_8017);
xor U9870 (N_9870,N_8444,N_8747);
xor U9871 (N_9871,N_8030,N_8095);
nor U9872 (N_9872,N_8010,N_8643);
nand U9873 (N_9873,N_8014,N_8948);
xor U9874 (N_9874,N_8262,N_8947);
nand U9875 (N_9875,N_8850,N_8908);
nand U9876 (N_9876,N_8826,N_8425);
nor U9877 (N_9877,N_8061,N_8830);
nor U9878 (N_9878,N_8406,N_8565);
and U9879 (N_9879,N_8830,N_8165);
and U9880 (N_9880,N_8967,N_8058);
nor U9881 (N_9881,N_8776,N_8455);
and U9882 (N_9882,N_8227,N_8927);
nand U9883 (N_9883,N_8530,N_8289);
and U9884 (N_9884,N_8572,N_8527);
nor U9885 (N_9885,N_8696,N_8701);
or U9886 (N_9886,N_8711,N_8330);
xor U9887 (N_9887,N_8302,N_8469);
or U9888 (N_9888,N_8584,N_8065);
or U9889 (N_9889,N_8554,N_8728);
or U9890 (N_9890,N_8761,N_8691);
or U9891 (N_9891,N_8088,N_8488);
nor U9892 (N_9892,N_8199,N_8125);
xnor U9893 (N_9893,N_8174,N_8250);
or U9894 (N_9894,N_8829,N_8721);
and U9895 (N_9895,N_8233,N_8311);
nor U9896 (N_9896,N_8460,N_8355);
and U9897 (N_9897,N_8329,N_8811);
xnor U9898 (N_9898,N_8389,N_8269);
nor U9899 (N_9899,N_8572,N_8885);
nand U9900 (N_9900,N_8721,N_8734);
and U9901 (N_9901,N_8736,N_8748);
nand U9902 (N_9902,N_8171,N_8922);
or U9903 (N_9903,N_8272,N_8601);
xnor U9904 (N_9904,N_8781,N_8899);
nor U9905 (N_9905,N_8828,N_8440);
xor U9906 (N_9906,N_8670,N_8904);
nand U9907 (N_9907,N_8931,N_8895);
and U9908 (N_9908,N_8653,N_8492);
nor U9909 (N_9909,N_8922,N_8990);
nand U9910 (N_9910,N_8241,N_8354);
xor U9911 (N_9911,N_8676,N_8659);
nand U9912 (N_9912,N_8805,N_8909);
xor U9913 (N_9913,N_8526,N_8951);
or U9914 (N_9914,N_8781,N_8732);
and U9915 (N_9915,N_8563,N_8922);
nand U9916 (N_9916,N_8371,N_8777);
nor U9917 (N_9917,N_8669,N_8654);
nor U9918 (N_9918,N_8562,N_8847);
and U9919 (N_9919,N_8889,N_8545);
nand U9920 (N_9920,N_8565,N_8647);
nand U9921 (N_9921,N_8639,N_8977);
xnor U9922 (N_9922,N_8235,N_8358);
nand U9923 (N_9923,N_8135,N_8915);
or U9924 (N_9924,N_8403,N_8762);
nand U9925 (N_9925,N_8226,N_8018);
or U9926 (N_9926,N_8762,N_8832);
nor U9927 (N_9927,N_8610,N_8306);
nand U9928 (N_9928,N_8552,N_8383);
and U9929 (N_9929,N_8825,N_8256);
nor U9930 (N_9930,N_8454,N_8208);
nor U9931 (N_9931,N_8065,N_8606);
xnor U9932 (N_9932,N_8620,N_8780);
nand U9933 (N_9933,N_8298,N_8199);
nor U9934 (N_9934,N_8048,N_8777);
nand U9935 (N_9935,N_8636,N_8247);
xor U9936 (N_9936,N_8452,N_8261);
nor U9937 (N_9937,N_8360,N_8259);
and U9938 (N_9938,N_8293,N_8032);
and U9939 (N_9939,N_8809,N_8616);
nor U9940 (N_9940,N_8566,N_8434);
xor U9941 (N_9941,N_8867,N_8712);
xor U9942 (N_9942,N_8985,N_8058);
and U9943 (N_9943,N_8277,N_8130);
xnor U9944 (N_9944,N_8231,N_8328);
nor U9945 (N_9945,N_8799,N_8050);
xnor U9946 (N_9946,N_8041,N_8338);
and U9947 (N_9947,N_8829,N_8545);
nand U9948 (N_9948,N_8125,N_8496);
or U9949 (N_9949,N_8782,N_8928);
nor U9950 (N_9950,N_8666,N_8031);
or U9951 (N_9951,N_8496,N_8948);
xor U9952 (N_9952,N_8218,N_8172);
or U9953 (N_9953,N_8858,N_8361);
or U9954 (N_9954,N_8161,N_8099);
nand U9955 (N_9955,N_8641,N_8958);
or U9956 (N_9956,N_8761,N_8322);
and U9957 (N_9957,N_8778,N_8031);
or U9958 (N_9958,N_8782,N_8198);
nor U9959 (N_9959,N_8048,N_8829);
or U9960 (N_9960,N_8246,N_8873);
nor U9961 (N_9961,N_8425,N_8630);
nand U9962 (N_9962,N_8490,N_8146);
or U9963 (N_9963,N_8261,N_8417);
nand U9964 (N_9964,N_8778,N_8212);
or U9965 (N_9965,N_8530,N_8051);
or U9966 (N_9966,N_8584,N_8424);
nor U9967 (N_9967,N_8407,N_8543);
nand U9968 (N_9968,N_8991,N_8670);
and U9969 (N_9969,N_8189,N_8489);
xor U9970 (N_9970,N_8825,N_8953);
or U9971 (N_9971,N_8634,N_8713);
or U9972 (N_9972,N_8004,N_8309);
and U9973 (N_9973,N_8677,N_8856);
or U9974 (N_9974,N_8159,N_8995);
nand U9975 (N_9975,N_8850,N_8091);
nand U9976 (N_9976,N_8656,N_8848);
xnor U9977 (N_9977,N_8268,N_8035);
or U9978 (N_9978,N_8101,N_8150);
xor U9979 (N_9979,N_8707,N_8133);
nand U9980 (N_9980,N_8903,N_8665);
and U9981 (N_9981,N_8794,N_8368);
xnor U9982 (N_9982,N_8094,N_8361);
and U9983 (N_9983,N_8929,N_8621);
nand U9984 (N_9984,N_8393,N_8724);
nor U9985 (N_9985,N_8943,N_8586);
nor U9986 (N_9986,N_8566,N_8476);
nor U9987 (N_9987,N_8307,N_8268);
nand U9988 (N_9988,N_8426,N_8830);
xnor U9989 (N_9989,N_8738,N_8991);
nor U9990 (N_9990,N_8132,N_8223);
xnor U9991 (N_9991,N_8138,N_8402);
nor U9992 (N_9992,N_8942,N_8480);
xor U9993 (N_9993,N_8208,N_8938);
and U9994 (N_9994,N_8568,N_8718);
xnor U9995 (N_9995,N_8699,N_8438);
and U9996 (N_9996,N_8370,N_8162);
nand U9997 (N_9997,N_8549,N_8365);
nand U9998 (N_9998,N_8421,N_8166);
or U9999 (N_9999,N_8474,N_8497);
or U10000 (N_10000,N_9481,N_9424);
xor U10001 (N_10001,N_9755,N_9610);
or U10002 (N_10002,N_9125,N_9508);
nor U10003 (N_10003,N_9007,N_9389);
and U10004 (N_10004,N_9153,N_9079);
nand U10005 (N_10005,N_9385,N_9824);
or U10006 (N_10006,N_9620,N_9047);
xnor U10007 (N_10007,N_9855,N_9783);
nor U10008 (N_10008,N_9842,N_9509);
nand U10009 (N_10009,N_9517,N_9780);
nor U10010 (N_10010,N_9694,N_9484);
or U10011 (N_10011,N_9496,N_9749);
nor U10012 (N_10012,N_9851,N_9272);
nor U10013 (N_10013,N_9378,N_9488);
xor U10014 (N_10014,N_9819,N_9564);
xnor U10015 (N_10015,N_9814,N_9663);
nor U10016 (N_10016,N_9394,N_9284);
and U10017 (N_10017,N_9067,N_9063);
nand U10018 (N_10018,N_9305,N_9585);
nor U10019 (N_10019,N_9023,N_9977);
xnor U10020 (N_10020,N_9471,N_9266);
xor U10021 (N_10021,N_9062,N_9836);
nand U10022 (N_10022,N_9794,N_9511);
xnor U10023 (N_10023,N_9562,N_9301);
nand U10024 (N_10024,N_9945,N_9539);
nor U10025 (N_10025,N_9691,N_9924);
nor U10026 (N_10026,N_9628,N_9269);
or U10027 (N_10027,N_9261,N_9144);
xor U10028 (N_10028,N_9798,N_9263);
and U10029 (N_10029,N_9561,N_9793);
xnor U10030 (N_10030,N_9558,N_9510);
nand U10031 (N_10031,N_9831,N_9392);
xnor U10032 (N_10032,N_9299,N_9138);
nor U10033 (N_10033,N_9766,N_9859);
xnor U10034 (N_10034,N_9887,N_9817);
xnor U10035 (N_10035,N_9487,N_9688);
nand U10036 (N_10036,N_9675,N_9160);
nor U10037 (N_10037,N_9233,N_9380);
nand U10038 (N_10038,N_9340,N_9122);
nand U10039 (N_10039,N_9148,N_9989);
xnor U10040 (N_10040,N_9974,N_9686);
and U10041 (N_10041,N_9210,N_9692);
and U10042 (N_10042,N_9698,N_9123);
and U10043 (N_10043,N_9024,N_9297);
and U10044 (N_10044,N_9529,N_9938);
or U10045 (N_10045,N_9760,N_9244);
or U10046 (N_10046,N_9041,N_9239);
nand U10047 (N_10047,N_9566,N_9942);
nor U10048 (N_10048,N_9782,N_9472);
xnor U10049 (N_10049,N_9020,N_9839);
nand U10050 (N_10050,N_9594,N_9386);
xnor U10051 (N_10051,N_9640,N_9161);
and U10052 (N_10052,N_9918,N_9255);
and U10053 (N_10053,N_9083,N_9056);
and U10054 (N_10054,N_9458,N_9711);
nor U10055 (N_10055,N_9554,N_9453);
or U10056 (N_10056,N_9913,N_9504);
and U10057 (N_10057,N_9136,N_9296);
nand U10058 (N_10058,N_9046,N_9601);
and U10059 (N_10059,N_9352,N_9682);
or U10060 (N_10060,N_9100,N_9571);
xnor U10061 (N_10061,N_9750,N_9057);
xor U10062 (N_10062,N_9823,N_9367);
xor U10063 (N_10063,N_9661,N_9575);
or U10064 (N_10064,N_9218,N_9507);
xnor U10065 (N_10065,N_9892,N_9770);
xnor U10066 (N_10066,N_9286,N_9528);
or U10067 (N_10067,N_9897,N_9489);
nand U10068 (N_10068,N_9486,N_9133);
and U10069 (N_10069,N_9593,N_9280);
or U10070 (N_10070,N_9717,N_9408);
and U10071 (N_10071,N_9442,N_9006);
xor U10072 (N_10072,N_9145,N_9420);
nand U10073 (N_10073,N_9664,N_9463);
nor U10074 (N_10074,N_9723,N_9372);
and U10075 (N_10075,N_9548,N_9492);
and U10076 (N_10076,N_9777,N_9583);
nor U10077 (N_10077,N_9344,N_9573);
or U10078 (N_10078,N_9584,N_9864);
or U10079 (N_10079,N_9095,N_9306);
or U10080 (N_10080,N_9812,N_9128);
or U10081 (N_10081,N_9633,N_9282);
nor U10082 (N_10082,N_9764,N_9448);
nor U10083 (N_10083,N_9973,N_9607);
nand U10084 (N_10084,N_9475,N_9910);
nand U10085 (N_10085,N_9157,N_9637);
and U10086 (N_10086,N_9337,N_9807);
nor U10087 (N_10087,N_9107,N_9165);
nor U10088 (N_10088,N_9333,N_9546);
xnor U10089 (N_10089,N_9235,N_9181);
and U10090 (N_10090,N_9848,N_9776);
or U10091 (N_10091,N_9746,N_9183);
nand U10092 (N_10092,N_9671,N_9615);
and U10093 (N_10093,N_9695,N_9479);
nor U10094 (N_10094,N_9844,N_9801);
xnor U10095 (N_10095,N_9240,N_9888);
nor U10096 (N_10096,N_9061,N_9689);
nand U10097 (N_10097,N_9912,N_9590);
and U10098 (N_10098,N_9478,N_9343);
nand U10099 (N_10099,N_9720,N_9099);
and U10100 (N_10100,N_9256,N_9310);
nor U10101 (N_10101,N_9000,N_9738);
nand U10102 (N_10102,N_9319,N_9495);
xor U10103 (N_10103,N_9792,N_9289);
xnor U10104 (N_10104,N_9521,N_9150);
nand U10105 (N_10105,N_9200,N_9719);
xor U10106 (N_10106,N_9121,N_9934);
and U10107 (N_10107,N_9645,N_9791);
nand U10108 (N_10108,N_9983,N_9098);
nor U10109 (N_10109,N_9903,N_9565);
xnor U10110 (N_10110,N_9763,N_9085);
nor U10111 (N_10111,N_9962,N_9984);
nand U10112 (N_10112,N_9440,N_9332);
or U10113 (N_10113,N_9568,N_9051);
or U10114 (N_10114,N_9541,N_9416);
nor U10115 (N_10115,N_9787,N_9435);
xnor U10116 (N_10116,N_9363,N_9952);
nand U10117 (N_10117,N_9781,N_9642);
nand U10118 (N_10118,N_9961,N_9089);
and U10119 (N_10119,N_9609,N_9957);
and U10120 (N_10120,N_9512,N_9908);
and U10121 (N_10121,N_9168,N_9230);
nand U10122 (N_10122,N_9731,N_9221);
nor U10123 (N_10123,N_9745,N_9674);
or U10124 (N_10124,N_9581,N_9676);
xor U10125 (N_10125,N_9335,N_9520);
and U10126 (N_10126,N_9011,N_9223);
nand U10127 (N_10127,N_9152,N_9081);
and U10128 (N_10128,N_9460,N_9025);
or U10129 (N_10129,N_9769,N_9874);
nand U10130 (N_10130,N_9834,N_9617);
xnor U10131 (N_10131,N_9369,N_9276);
and U10132 (N_10132,N_9660,N_9464);
xor U10133 (N_10133,N_9929,N_9368);
and U10134 (N_10134,N_9778,N_9680);
xnor U10135 (N_10135,N_9170,N_9841);
xnor U10136 (N_10136,N_9014,N_9253);
and U10137 (N_10137,N_9856,N_9326);
nor U10138 (N_10138,N_9298,N_9461);
nand U10139 (N_10139,N_9733,N_9423);
xnor U10140 (N_10140,N_9055,N_9375);
and U10141 (N_10141,N_9188,N_9709);
or U10142 (N_10142,N_9234,N_9884);
and U10143 (N_10143,N_9656,N_9515);
nand U10144 (N_10144,N_9533,N_9911);
nor U10145 (N_10145,N_9714,N_9936);
and U10146 (N_10146,N_9644,N_9053);
or U10147 (N_10147,N_9124,N_9197);
nor U10148 (N_10148,N_9390,N_9701);
and U10149 (N_10149,N_9456,N_9748);
nand U10150 (N_10150,N_9228,N_9909);
and U10151 (N_10151,N_9459,N_9741);
or U10152 (N_10152,N_9948,N_9670);
nor U10153 (N_10153,N_9825,N_9570);
nor U10154 (N_10154,N_9104,N_9826);
nand U10155 (N_10155,N_9870,N_9430);
or U10156 (N_10156,N_9699,N_9684);
or U10157 (N_10157,N_9574,N_9632);
xnor U10158 (N_10158,N_9623,N_9101);
nor U10159 (N_10159,N_9202,N_9470);
nand U10160 (N_10160,N_9074,N_9576);
xor U10161 (N_10161,N_9214,N_9904);
xor U10162 (N_10162,N_9606,N_9578);
and U10163 (N_10163,N_9252,N_9937);
or U10164 (N_10164,N_9796,N_9498);
and U10165 (N_10165,N_9679,N_9643);
and U10166 (N_10166,N_9873,N_9401);
and U10167 (N_10167,N_9920,N_9923);
or U10168 (N_10168,N_9681,N_9092);
and U10169 (N_10169,N_9991,N_9001);
xnor U10170 (N_10170,N_9027,N_9556);
nor U10171 (N_10171,N_9900,N_9706);
nand U10172 (N_10172,N_9330,N_9015);
and U10173 (N_10173,N_9111,N_9547);
and U10174 (N_10174,N_9754,N_9229);
nand U10175 (N_10175,N_9756,N_9032);
and U10176 (N_10176,N_9768,N_9209);
or U10177 (N_10177,N_9786,N_9894);
nor U10178 (N_10178,N_9166,N_9175);
and U10179 (N_10179,N_9550,N_9441);
nor U10180 (N_10180,N_9320,N_9968);
or U10181 (N_10181,N_9451,N_9905);
and U10182 (N_10182,N_9619,N_9143);
nor U10183 (N_10183,N_9759,N_9821);
xor U10184 (N_10184,N_9017,N_9052);
nor U10185 (N_10185,N_9321,N_9499);
or U10186 (N_10186,N_9480,N_9350);
nand U10187 (N_10187,N_9278,N_9523);
or U10188 (N_10188,N_9355,N_9975);
xor U10189 (N_10189,N_9673,N_9194);
nor U10190 (N_10190,N_9928,N_9260);
xor U10191 (N_10191,N_9611,N_9790);
and U10192 (N_10192,N_9088,N_9112);
nor U10193 (N_10193,N_9324,N_9718);
nand U10194 (N_10194,N_9603,N_9341);
nand U10195 (N_10195,N_9708,N_9653);
nor U10196 (N_10196,N_9932,N_9655);
nor U10197 (N_10197,N_9881,N_9012);
or U10198 (N_10198,N_9906,N_9516);
nand U10199 (N_10199,N_9518,N_9802);
and U10200 (N_10200,N_9428,N_9612);
nor U10201 (N_10201,N_9384,N_9201);
and U10202 (N_10202,N_9354,N_9858);
nand U10203 (N_10203,N_9846,N_9195);
nor U10204 (N_10204,N_9037,N_9734);
nor U10205 (N_10205,N_9028,N_9106);
xnor U10206 (N_10206,N_9947,N_9572);
and U10207 (N_10207,N_9608,N_9172);
and U10208 (N_10208,N_9677,N_9816);
nor U10209 (N_10209,N_9141,N_9018);
or U10210 (N_10210,N_9598,N_9494);
xnor U10211 (N_10211,N_9371,N_9361);
and U10212 (N_10212,N_9935,N_9334);
nor U10213 (N_10213,N_9449,N_9365);
xnor U10214 (N_10214,N_9293,N_9086);
nand U10215 (N_10215,N_9998,N_9752);
and U10216 (N_10216,N_9788,N_9290);
nand U10217 (N_10217,N_9277,N_9569);
nor U10218 (N_10218,N_9159,N_9105);
or U10219 (N_10219,N_9419,N_9308);
xnor U10220 (N_10220,N_9134,N_9462);
nor U10221 (N_10221,N_9431,N_9285);
nor U10222 (N_10222,N_9312,N_9466);
nor U10223 (N_10223,N_9281,N_9360);
or U10224 (N_10224,N_9065,N_9732);
or U10225 (N_10225,N_9251,N_9818);
xnor U10226 (N_10226,N_9662,N_9031);
or U10227 (N_10227,N_9432,N_9436);
or U10228 (N_10228,N_9995,N_9147);
or U10229 (N_10229,N_9454,N_9097);
nand U10230 (N_10230,N_9596,N_9485);
nor U10231 (N_10231,N_9059,N_9325);
nor U10232 (N_10232,N_9901,N_9762);
nor U10233 (N_10233,N_9693,N_9697);
and U10234 (N_10234,N_9477,N_9323);
or U10235 (N_10235,N_9589,N_9429);
xor U10236 (N_10236,N_9724,N_9930);
nor U10237 (N_10237,N_9403,N_9060);
or U10238 (N_10238,N_9852,N_9635);
or U10239 (N_10239,N_9503,N_9199);
xor U10240 (N_10240,N_9896,N_9311);
nand U10241 (N_10241,N_9127,N_9482);
and U10242 (N_10242,N_9117,N_9739);
nand U10243 (N_10243,N_9916,N_9810);
xor U10244 (N_10244,N_9189,N_9193);
nor U10245 (N_10245,N_9187,N_9502);
and U10246 (N_10246,N_9592,N_9019);
xnor U10247 (N_10247,N_9455,N_9652);
and U10248 (N_10248,N_9331,N_9907);
xnor U10249 (N_10249,N_9922,N_9156);
or U10250 (N_10250,N_9353,N_9054);
nor U10251 (N_10251,N_9009,N_9999);
xor U10252 (N_10252,N_9182,N_9066);
xor U10253 (N_10253,N_9070,N_9345);
or U10254 (N_10254,N_9207,N_9543);
xnor U10255 (N_10255,N_9618,N_9467);
xnor U10256 (N_10256,N_9316,N_9035);
xnor U10257 (N_10257,N_9026,N_9469);
or U10258 (N_10258,N_9191,N_9933);
nand U10259 (N_10259,N_9437,N_9877);
and U10260 (N_10260,N_9958,N_9291);
nand U10261 (N_10261,N_9672,N_9602);
nor U10262 (N_10262,N_9336,N_9154);
nor U10263 (N_10263,N_9624,N_9075);
or U10264 (N_10264,N_9967,N_9943);
and U10265 (N_10265,N_9555,N_9808);
nand U10266 (N_10266,N_9102,N_9542);
or U10267 (N_10267,N_9765,N_9010);
or U10268 (N_10268,N_9120,N_9730);
xor U10269 (N_10269,N_9950,N_9425);
nor U10270 (N_10270,N_9076,N_9580);
xor U10271 (N_10271,N_9667,N_9599);
or U10272 (N_10272,N_9418,N_9130);
or U10273 (N_10273,N_9500,N_9225);
nor U10274 (N_10274,N_9072,N_9833);
xor U10275 (N_10275,N_9109,N_9534);
xor U10276 (N_10276,N_9443,N_9315);
xnor U10277 (N_10277,N_9397,N_9295);
nor U10278 (N_10278,N_9275,N_9174);
xor U10279 (N_10279,N_9034,N_9946);
xnor U10280 (N_10280,N_9468,N_9177);
and U10281 (N_10281,N_9213,N_9728);
and U10282 (N_10282,N_9803,N_9422);
xnor U10283 (N_10283,N_9043,N_9996);
xor U10284 (N_10284,N_9445,N_9410);
and U10285 (N_10285,N_9268,N_9142);
nor U10286 (N_10286,N_9273,N_9951);
nand U10287 (N_10287,N_9891,N_9205);
xor U10288 (N_10288,N_9115,N_9283);
nand U10289 (N_10289,N_9358,N_9342);
nor U10290 (N_10290,N_9567,N_9224);
xor U10291 (N_10291,N_9530,N_9267);
and U10292 (N_10292,N_9309,N_9868);
nor U10293 (N_10293,N_9867,N_9753);
and U10294 (N_10294,N_9953,N_9069);
or U10295 (N_10295,N_9402,N_9257);
nor U10296 (N_10296,N_9862,N_9250);
and U10297 (N_10297,N_9044,N_9822);
and U10298 (N_10298,N_9346,N_9114);
nor U10299 (N_10299,N_9885,N_9433);
nor U10300 (N_10300,N_9162,N_9005);
nand U10301 (N_10301,N_9068,N_9743);
and U10302 (N_10302,N_9863,N_9004);
and U10303 (N_10303,N_9497,N_9190);
nand U10304 (N_10304,N_9356,N_9621);
nor U10305 (N_10305,N_9203,N_9158);
and U10306 (N_10306,N_9669,N_9016);
xor U10307 (N_10307,N_9806,N_9540);
or U10308 (N_10308,N_9129,N_9288);
or U10309 (N_10309,N_9217,N_9427);
nand U10310 (N_10310,N_9595,N_9860);
and U10311 (N_10311,N_9587,N_9634);
or U10312 (N_10312,N_9579,N_9215);
nand U10313 (N_10313,N_9990,N_9740);
xnor U10314 (N_10314,N_9625,N_9505);
and U10315 (N_10315,N_9292,N_9735);
xor U10316 (N_10316,N_9982,N_9220);
nand U10317 (N_10317,N_9374,N_9704);
xor U10318 (N_10318,N_9362,N_9399);
nand U10319 (N_10319,N_9837,N_9538);
or U10320 (N_10320,N_9779,N_9404);
nand U10321 (N_10321,N_9208,N_9600);
and U10322 (N_10322,N_9614,N_9767);
and U10323 (N_10323,N_9966,N_9994);
and U10324 (N_10324,N_9163,N_9048);
and U10325 (N_10325,N_9785,N_9744);
xnor U10326 (N_10326,N_9176,N_9872);
and U10327 (N_10327,N_9549,N_9997);
xor U10328 (N_10328,N_9560,N_9981);
nand U10329 (N_10329,N_9038,N_9631);
or U10330 (N_10330,N_9696,N_9113);
or U10331 (N_10331,N_9232,N_9829);
and U10332 (N_10332,N_9438,N_9514);
nand U10333 (N_10333,N_9939,N_9963);
and U10334 (N_10334,N_9917,N_9108);
nor U10335 (N_10335,N_9992,N_9532);
and U10336 (N_10336,N_9683,N_9364);
xnor U10337 (N_10337,N_9513,N_9751);
and U10338 (N_10338,N_9976,N_9042);
and U10339 (N_10339,N_9050,N_9525);
and U10340 (N_10340,N_9925,N_9204);
nor U10341 (N_10341,N_9164,N_9237);
and U10342 (N_10342,N_9828,N_9545);
and U10343 (N_10343,N_9940,N_9119);
xor U10344 (N_10344,N_9805,N_9902);
nor U10345 (N_10345,N_9096,N_9956);
nand U10346 (N_10346,N_9247,N_9775);
xnor U10347 (N_10347,N_9270,N_9536);
or U10348 (N_10348,N_9969,N_9407);
and U10349 (N_10349,N_9377,N_9021);
nor U10350 (N_10350,N_9591,N_9700);
xor U10351 (N_10351,N_9737,N_9970);
nand U10352 (N_10352,N_9830,N_9131);
or U10353 (N_10353,N_9029,N_9710);
nand U10354 (N_10354,N_9965,N_9639);
nand U10355 (N_10355,N_9294,N_9880);
nor U10356 (N_10356,N_9597,N_9093);
or U10357 (N_10357,N_9169,N_9003);
or U10358 (N_10358,N_9465,N_9702);
nand U10359 (N_10359,N_9627,N_9955);
and U10360 (N_10360,N_9211,N_9985);
or U10361 (N_10361,N_9827,N_9077);
xor U10362 (N_10362,N_9064,N_9577);
and U10363 (N_10363,N_9657,N_9231);
and U10364 (N_10364,N_9022,N_9426);
and U10365 (N_10365,N_9626,N_9960);
nand U10366 (N_10366,N_9915,N_9654);
xnor U10367 (N_10367,N_9307,N_9605);
and U10368 (N_10368,N_9993,N_9804);
nor U10369 (N_10369,N_9490,N_9789);
xnor U10370 (N_10370,N_9665,N_9649);
or U10371 (N_10371,N_9483,N_9721);
or U10372 (N_10372,N_9800,N_9450);
or U10373 (N_10373,N_9381,N_9238);
nor U10374 (N_10374,N_9893,N_9382);
nand U10375 (N_10375,N_9313,N_9444);
or U10376 (N_10376,N_9491,N_9373);
nor U10377 (N_10377,N_9388,N_9434);
nand U10378 (N_10378,N_9883,N_9987);
nor U10379 (N_10379,N_9651,N_9379);
or U10380 (N_10380,N_9348,N_9716);
nor U10381 (N_10381,N_9265,N_9359);
nand U10382 (N_10382,N_9033,N_9452);
and U10383 (N_10383,N_9964,N_9857);
xnor U10384 (N_10384,N_9198,N_9249);
and U10385 (N_10385,N_9087,N_9882);
nand U10386 (N_10386,N_9103,N_9411);
and U10387 (N_10387,N_9110,N_9302);
or U10388 (N_10388,N_9271,N_9522);
xnor U10389 (N_10389,N_9832,N_9091);
or U10390 (N_10390,N_9414,N_9002);
nor U10391 (N_10391,N_9537,N_9895);
nand U10392 (N_10392,N_9212,N_9135);
and U10393 (N_10393,N_9185,N_9889);
and U10394 (N_10394,N_9526,N_9685);
xnor U10395 (N_10395,N_9146,N_9049);
nand U10396 (N_10396,N_9853,N_9527);
and U10397 (N_10397,N_9866,N_9415);
nand U10398 (N_10398,N_9279,N_9126);
and U10399 (N_10399,N_9927,N_9391);
nor U10400 (N_10400,N_9186,N_9668);
or U10401 (N_10401,N_9811,N_9641);
nor U10402 (N_10402,N_9899,N_9328);
or U10403 (N_10403,N_9264,N_9588);
nor U10404 (N_10404,N_9073,N_9357);
xnor U10405 (N_10405,N_9322,N_9582);
xor U10406 (N_10406,N_9446,N_9687);
xnor U10407 (N_10407,N_9400,N_9551);
nor U10408 (N_10408,N_9725,N_9219);
nand U10409 (N_10409,N_9245,N_9493);
nor U10410 (N_10410,N_9604,N_9758);
and U10411 (N_10411,N_9300,N_9757);
nor U10412 (N_10412,N_9242,N_9222);
and U10413 (N_10413,N_9155,N_9835);
xor U10414 (N_10414,N_9854,N_9151);
and U10415 (N_10415,N_9613,N_9226);
or U10416 (N_10416,N_9406,N_9036);
or U10417 (N_10417,N_9678,N_9727);
or U10418 (N_10418,N_9557,N_9241);
xnor U10419 (N_10419,N_9008,N_9082);
nand U10420 (N_10420,N_9287,N_9729);
and U10421 (N_10421,N_9813,N_9393);
xnor U10422 (N_10422,N_9246,N_9616);
xnor U10423 (N_10423,N_9071,N_9742);
and U10424 (N_10424,N_9327,N_9959);
and U10425 (N_10425,N_9387,N_9931);
xor U10426 (N_10426,N_9647,N_9784);
nor U10427 (N_10427,N_9898,N_9838);
nand U10428 (N_10428,N_9712,N_9847);
or U10429 (N_10429,N_9771,N_9761);
or U10430 (N_10430,N_9876,N_9439);
nor U10431 (N_10431,N_9457,N_9949);
nor U10432 (N_10432,N_9366,N_9094);
and U10433 (N_10433,N_9843,N_9405);
and U10434 (N_10434,N_9879,N_9622);
nor U10435 (N_10435,N_9630,N_9173);
xor U10436 (N_10436,N_9886,N_9398);
nor U10437 (N_10437,N_9413,N_9317);
xor U10438 (N_10438,N_9988,N_9648);
and U10439 (N_10439,N_9347,N_9799);
xnor U10440 (N_10440,N_9919,N_9370);
and U10441 (N_10441,N_9149,N_9338);
nand U10442 (N_10442,N_9878,N_9412);
and U10443 (N_10443,N_9314,N_9132);
and U10444 (N_10444,N_9339,N_9206);
nor U10445 (N_10445,N_9795,N_9980);
or U10446 (N_10446,N_9262,N_9563);
and U10447 (N_10447,N_9180,N_9058);
nand U10448 (N_10448,N_9774,N_9329);
or U10449 (N_10449,N_9258,N_9040);
and U10450 (N_10450,N_9248,N_9476);
or U10451 (N_10451,N_9447,N_9629);
and U10452 (N_10452,N_9914,N_9986);
xor U10453 (N_10453,N_9736,N_9690);
nor U10454 (N_10454,N_9926,N_9944);
and U10455 (N_10455,N_9030,N_9658);
or U10456 (N_10456,N_9171,N_9179);
or U10457 (N_10457,N_9417,N_9318);
xor U10458 (N_10458,N_9845,N_9971);
xnor U10459 (N_10459,N_9921,N_9772);
nor U10460 (N_10460,N_9552,N_9524);
or U10461 (N_10461,N_9797,N_9840);
nor U10462 (N_10462,N_9713,N_9559);
nor U10463 (N_10463,N_9954,N_9553);
or U10464 (N_10464,N_9705,N_9167);
nand U10465 (N_10465,N_9116,N_9586);
nor U10466 (N_10466,N_9118,N_9090);
or U10467 (N_10467,N_9236,N_9303);
and U10468 (N_10468,N_9501,N_9715);
xnor U10469 (N_10469,N_9850,N_9137);
nand U10470 (N_10470,N_9544,N_9013);
or U10471 (N_10471,N_9216,N_9871);
nor U10472 (N_10472,N_9820,N_9045);
xnor U10473 (N_10473,N_9941,N_9726);
xnor U10474 (N_10474,N_9139,N_9636);
nand U10475 (N_10475,N_9861,N_9650);
xnor U10476 (N_10476,N_9383,N_9421);
and U10477 (N_10477,N_9815,N_9849);
and U10478 (N_10478,N_9473,N_9196);
xor U10479 (N_10479,N_9376,N_9809);
and U10480 (N_10480,N_9531,N_9349);
xor U10481 (N_10481,N_9396,N_9978);
nor U10482 (N_10482,N_9972,N_9395);
nor U10483 (N_10483,N_9869,N_9722);
xnor U10484 (N_10484,N_9184,N_9474);
and U10485 (N_10485,N_9084,N_9773);
nand U10486 (N_10486,N_9178,N_9703);
nand U10487 (N_10487,N_9646,N_9274);
and U10488 (N_10488,N_9409,N_9304);
and U10489 (N_10489,N_9875,N_9535);
and U10490 (N_10490,N_9890,N_9659);
and U10491 (N_10491,N_9519,N_9638);
nor U10492 (N_10492,N_9979,N_9078);
and U10493 (N_10493,N_9707,N_9140);
xnor U10494 (N_10494,N_9351,N_9259);
nor U10495 (N_10495,N_9747,N_9039);
xor U10496 (N_10496,N_9666,N_9192);
nand U10497 (N_10497,N_9506,N_9243);
and U10498 (N_10498,N_9227,N_9865);
nor U10499 (N_10499,N_9080,N_9254);
xnor U10500 (N_10500,N_9186,N_9922);
xnor U10501 (N_10501,N_9327,N_9623);
or U10502 (N_10502,N_9692,N_9551);
or U10503 (N_10503,N_9657,N_9073);
and U10504 (N_10504,N_9274,N_9016);
xor U10505 (N_10505,N_9074,N_9295);
or U10506 (N_10506,N_9403,N_9819);
nand U10507 (N_10507,N_9194,N_9022);
or U10508 (N_10508,N_9757,N_9340);
nor U10509 (N_10509,N_9885,N_9422);
and U10510 (N_10510,N_9462,N_9064);
nor U10511 (N_10511,N_9100,N_9243);
xor U10512 (N_10512,N_9885,N_9378);
nor U10513 (N_10513,N_9239,N_9739);
xnor U10514 (N_10514,N_9362,N_9291);
nor U10515 (N_10515,N_9001,N_9409);
nand U10516 (N_10516,N_9725,N_9798);
xor U10517 (N_10517,N_9991,N_9689);
or U10518 (N_10518,N_9688,N_9067);
nand U10519 (N_10519,N_9613,N_9758);
and U10520 (N_10520,N_9461,N_9506);
nor U10521 (N_10521,N_9232,N_9006);
and U10522 (N_10522,N_9504,N_9227);
xor U10523 (N_10523,N_9599,N_9067);
nand U10524 (N_10524,N_9041,N_9447);
nor U10525 (N_10525,N_9045,N_9453);
and U10526 (N_10526,N_9598,N_9622);
xor U10527 (N_10527,N_9671,N_9004);
xor U10528 (N_10528,N_9079,N_9867);
nand U10529 (N_10529,N_9380,N_9605);
nor U10530 (N_10530,N_9536,N_9022);
and U10531 (N_10531,N_9959,N_9418);
nand U10532 (N_10532,N_9096,N_9708);
nor U10533 (N_10533,N_9318,N_9450);
and U10534 (N_10534,N_9420,N_9664);
nor U10535 (N_10535,N_9149,N_9644);
nand U10536 (N_10536,N_9613,N_9325);
xor U10537 (N_10537,N_9886,N_9182);
nor U10538 (N_10538,N_9073,N_9519);
or U10539 (N_10539,N_9705,N_9232);
xor U10540 (N_10540,N_9861,N_9643);
nand U10541 (N_10541,N_9203,N_9923);
nor U10542 (N_10542,N_9260,N_9885);
or U10543 (N_10543,N_9338,N_9413);
xor U10544 (N_10544,N_9773,N_9302);
xor U10545 (N_10545,N_9757,N_9769);
and U10546 (N_10546,N_9328,N_9350);
and U10547 (N_10547,N_9948,N_9461);
nor U10548 (N_10548,N_9201,N_9020);
nor U10549 (N_10549,N_9330,N_9256);
nand U10550 (N_10550,N_9939,N_9040);
xnor U10551 (N_10551,N_9441,N_9396);
and U10552 (N_10552,N_9710,N_9220);
xnor U10553 (N_10553,N_9759,N_9170);
nand U10554 (N_10554,N_9618,N_9371);
and U10555 (N_10555,N_9005,N_9940);
nand U10556 (N_10556,N_9271,N_9235);
and U10557 (N_10557,N_9090,N_9142);
xnor U10558 (N_10558,N_9196,N_9283);
and U10559 (N_10559,N_9882,N_9598);
nor U10560 (N_10560,N_9123,N_9288);
nand U10561 (N_10561,N_9600,N_9517);
nand U10562 (N_10562,N_9202,N_9300);
or U10563 (N_10563,N_9835,N_9397);
and U10564 (N_10564,N_9306,N_9502);
or U10565 (N_10565,N_9262,N_9151);
nor U10566 (N_10566,N_9162,N_9691);
or U10567 (N_10567,N_9062,N_9417);
and U10568 (N_10568,N_9282,N_9647);
xnor U10569 (N_10569,N_9896,N_9743);
nor U10570 (N_10570,N_9852,N_9804);
nand U10571 (N_10571,N_9962,N_9749);
nand U10572 (N_10572,N_9722,N_9453);
nand U10573 (N_10573,N_9351,N_9296);
or U10574 (N_10574,N_9842,N_9947);
or U10575 (N_10575,N_9367,N_9986);
or U10576 (N_10576,N_9081,N_9809);
or U10577 (N_10577,N_9098,N_9722);
and U10578 (N_10578,N_9803,N_9951);
or U10579 (N_10579,N_9230,N_9145);
or U10580 (N_10580,N_9096,N_9012);
nand U10581 (N_10581,N_9318,N_9471);
or U10582 (N_10582,N_9657,N_9973);
xor U10583 (N_10583,N_9523,N_9820);
nand U10584 (N_10584,N_9717,N_9134);
xor U10585 (N_10585,N_9991,N_9236);
or U10586 (N_10586,N_9131,N_9858);
or U10587 (N_10587,N_9939,N_9777);
and U10588 (N_10588,N_9463,N_9314);
nor U10589 (N_10589,N_9266,N_9653);
nor U10590 (N_10590,N_9730,N_9607);
nor U10591 (N_10591,N_9789,N_9400);
nor U10592 (N_10592,N_9058,N_9032);
xnor U10593 (N_10593,N_9997,N_9596);
nor U10594 (N_10594,N_9148,N_9522);
xor U10595 (N_10595,N_9952,N_9048);
xor U10596 (N_10596,N_9913,N_9672);
nor U10597 (N_10597,N_9916,N_9582);
and U10598 (N_10598,N_9977,N_9028);
nand U10599 (N_10599,N_9884,N_9265);
and U10600 (N_10600,N_9913,N_9095);
and U10601 (N_10601,N_9681,N_9928);
or U10602 (N_10602,N_9512,N_9841);
xnor U10603 (N_10603,N_9369,N_9985);
nor U10604 (N_10604,N_9560,N_9387);
nor U10605 (N_10605,N_9495,N_9229);
xnor U10606 (N_10606,N_9465,N_9658);
xor U10607 (N_10607,N_9861,N_9818);
nor U10608 (N_10608,N_9461,N_9160);
or U10609 (N_10609,N_9495,N_9201);
nand U10610 (N_10610,N_9458,N_9159);
and U10611 (N_10611,N_9777,N_9769);
and U10612 (N_10612,N_9072,N_9864);
xor U10613 (N_10613,N_9654,N_9944);
xnor U10614 (N_10614,N_9723,N_9765);
or U10615 (N_10615,N_9945,N_9155);
and U10616 (N_10616,N_9693,N_9319);
and U10617 (N_10617,N_9157,N_9691);
and U10618 (N_10618,N_9896,N_9054);
or U10619 (N_10619,N_9814,N_9594);
nand U10620 (N_10620,N_9187,N_9055);
nor U10621 (N_10621,N_9863,N_9908);
xor U10622 (N_10622,N_9794,N_9780);
xnor U10623 (N_10623,N_9844,N_9102);
xnor U10624 (N_10624,N_9223,N_9746);
and U10625 (N_10625,N_9216,N_9135);
nor U10626 (N_10626,N_9639,N_9971);
or U10627 (N_10627,N_9181,N_9940);
nand U10628 (N_10628,N_9509,N_9899);
and U10629 (N_10629,N_9214,N_9245);
nand U10630 (N_10630,N_9565,N_9335);
and U10631 (N_10631,N_9039,N_9190);
and U10632 (N_10632,N_9367,N_9307);
xor U10633 (N_10633,N_9373,N_9410);
nor U10634 (N_10634,N_9527,N_9923);
xor U10635 (N_10635,N_9242,N_9155);
xnor U10636 (N_10636,N_9151,N_9478);
and U10637 (N_10637,N_9407,N_9813);
nor U10638 (N_10638,N_9465,N_9543);
nor U10639 (N_10639,N_9634,N_9283);
or U10640 (N_10640,N_9434,N_9378);
nor U10641 (N_10641,N_9417,N_9690);
and U10642 (N_10642,N_9313,N_9933);
and U10643 (N_10643,N_9112,N_9780);
xnor U10644 (N_10644,N_9525,N_9193);
xnor U10645 (N_10645,N_9151,N_9874);
or U10646 (N_10646,N_9034,N_9030);
and U10647 (N_10647,N_9003,N_9879);
nor U10648 (N_10648,N_9234,N_9982);
and U10649 (N_10649,N_9553,N_9195);
nor U10650 (N_10650,N_9098,N_9142);
nor U10651 (N_10651,N_9554,N_9570);
xor U10652 (N_10652,N_9886,N_9073);
nor U10653 (N_10653,N_9759,N_9508);
or U10654 (N_10654,N_9590,N_9433);
or U10655 (N_10655,N_9332,N_9583);
nand U10656 (N_10656,N_9068,N_9124);
xor U10657 (N_10657,N_9806,N_9318);
nor U10658 (N_10658,N_9668,N_9486);
xnor U10659 (N_10659,N_9951,N_9073);
xnor U10660 (N_10660,N_9270,N_9008);
xnor U10661 (N_10661,N_9601,N_9797);
and U10662 (N_10662,N_9571,N_9207);
nand U10663 (N_10663,N_9080,N_9887);
nor U10664 (N_10664,N_9841,N_9552);
nand U10665 (N_10665,N_9798,N_9133);
and U10666 (N_10666,N_9520,N_9067);
nor U10667 (N_10667,N_9266,N_9137);
nand U10668 (N_10668,N_9557,N_9387);
nor U10669 (N_10669,N_9355,N_9853);
or U10670 (N_10670,N_9382,N_9946);
nor U10671 (N_10671,N_9404,N_9726);
nor U10672 (N_10672,N_9698,N_9186);
nor U10673 (N_10673,N_9893,N_9294);
or U10674 (N_10674,N_9609,N_9213);
xor U10675 (N_10675,N_9506,N_9363);
xor U10676 (N_10676,N_9589,N_9077);
and U10677 (N_10677,N_9957,N_9644);
and U10678 (N_10678,N_9598,N_9506);
nand U10679 (N_10679,N_9540,N_9467);
xnor U10680 (N_10680,N_9176,N_9363);
nand U10681 (N_10681,N_9815,N_9023);
or U10682 (N_10682,N_9336,N_9374);
xor U10683 (N_10683,N_9285,N_9188);
nand U10684 (N_10684,N_9625,N_9617);
and U10685 (N_10685,N_9966,N_9042);
nor U10686 (N_10686,N_9159,N_9701);
nand U10687 (N_10687,N_9911,N_9233);
xnor U10688 (N_10688,N_9232,N_9174);
or U10689 (N_10689,N_9683,N_9869);
nor U10690 (N_10690,N_9986,N_9796);
nor U10691 (N_10691,N_9832,N_9025);
or U10692 (N_10692,N_9985,N_9832);
or U10693 (N_10693,N_9141,N_9215);
or U10694 (N_10694,N_9332,N_9611);
nor U10695 (N_10695,N_9166,N_9471);
xor U10696 (N_10696,N_9906,N_9533);
and U10697 (N_10697,N_9749,N_9321);
or U10698 (N_10698,N_9448,N_9489);
and U10699 (N_10699,N_9738,N_9107);
or U10700 (N_10700,N_9847,N_9376);
xor U10701 (N_10701,N_9592,N_9732);
and U10702 (N_10702,N_9077,N_9319);
or U10703 (N_10703,N_9917,N_9920);
or U10704 (N_10704,N_9475,N_9674);
or U10705 (N_10705,N_9541,N_9632);
or U10706 (N_10706,N_9013,N_9198);
xnor U10707 (N_10707,N_9737,N_9695);
or U10708 (N_10708,N_9639,N_9484);
nand U10709 (N_10709,N_9623,N_9280);
xnor U10710 (N_10710,N_9930,N_9575);
and U10711 (N_10711,N_9261,N_9502);
nor U10712 (N_10712,N_9046,N_9583);
xnor U10713 (N_10713,N_9508,N_9196);
xnor U10714 (N_10714,N_9815,N_9032);
nor U10715 (N_10715,N_9865,N_9500);
and U10716 (N_10716,N_9097,N_9518);
xnor U10717 (N_10717,N_9468,N_9294);
and U10718 (N_10718,N_9131,N_9917);
nor U10719 (N_10719,N_9756,N_9063);
xnor U10720 (N_10720,N_9563,N_9521);
and U10721 (N_10721,N_9929,N_9414);
and U10722 (N_10722,N_9772,N_9838);
nand U10723 (N_10723,N_9229,N_9728);
or U10724 (N_10724,N_9224,N_9029);
nand U10725 (N_10725,N_9337,N_9871);
or U10726 (N_10726,N_9719,N_9466);
nand U10727 (N_10727,N_9720,N_9016);
xnor U10728 (N_10728,N_9610,N_9656);
nand U10729 (N_10729,N_9892,N_9285);
nand U10730 (N_10730,N_9494,N_9617);
or U10731 (N_10731,N_9338,N_9465);
xnor U10732 (N_10732,N_9467,N_9985);
xor U10733 (N_10733,N_9184,N_9078);
nor U10734 (N_10734,N_9391,N_9392);
xnor U10735 (N_10735,N_9729,N_9709);
nand U10736 (N_10736,N_9281,N_9369);
nor U10737 (N_10737,N_9467,N_9128);
nand U10738 (N_10738,N_9050,N_9279);
nand U10739 (N_10739,N_9098,N_9501);
xor U10740 (N_10740,N_9466,N_9629);
xnor U10741 (N_10741,N_9445,N_9671);
xor U10742 (N_10742,N_9218,N_9991);
nand U10743 (N_10743,N_9378,N_9091);
xor U10744 (N_10744,N_9454,N_9009);
xor U10745 (N_10745,N_9633,N_9250);
or U10746 (N_10746,N_9956,N_9650);
and U10747 (N_10747,N_9471,N_9385);
nor U10748 (N_10748,N_9430,N_9564);
or U10749 (N_10749,N_9149,N_9146);
nor U10750 (N_10750,N_9576,N_9930);
nand U10751 (N_10751,N_9296,N_9311);
nand U10752 (N_10752,N_9384,N_9318);
and U10753 (N_10753,N_9489,N_9815);
nor U10754 (N_10754,N_9076,N_9313);
or U10755 (N_10755,N_9485,N_9520);
or U10756 (N_10756,N_9133,N_9233);
nand U10757 (N_10757,N_9518,N_9466);
nor U10758 (N_10758,N_9399,N_9820);
nor U10759 (N_10759,N_9887,N_9944);
nor U10760 (N_10760,N_9574,N_9722);
nor U10761 (N_10761,N_9054,N_9285);
and U10762 (N_10762,N_9676,N_9484);
nor U10763 (N_10763,N_9937,N_9256);
or U10764 (N_10764,N_9292,N_9061);
nand U10765 (N_10765,N_9297,N_9282);
nor U10766 (N_10766,N_9015,N_9197);
or U10767 (N_10767,N_9131,N_9892);
or U10768 (N_10768,N_9424,N_9618);
xor U10769 (N_10769,N_9116,N_9416);
nor U10770 (N_10770,N_9630,N_9683);
and U10771 (N_10771,N_9492,N_9506);
xnor U10772 (N_10772,N_9596,N_9155);
nand U10773 (N_10773,N_9323,N_9764);
xnor U10774 (N_10774,N_9358,N_9058);
nor U10775 (N_10775,N_9173,N_9925);
nand U10776 (N_10776,N_9443,N_9565);
and U10777 (N_10777,N_9807,N_9263);
or U10778 (N_10778,N_9037,N_9373);
or U10779 (N_10779,N_9026,N_9821);
and U10780 (N_10780,N_9222,N_9686);
and U10781 (N_10781,N_9909,N_9650);
xnor U10782 (N_10782,N_9962,N_9046);
or U10783 (N_10783,N_9214,N_9751);
xnor U10784 (N_10784,N_9151,N_9484);
nand U10785 (N_10785,N_9503,N_9000);
xor U10786 (N_10786,N_9409,N_9380);
nand U10787 (N_10787,N_9429,N_9260);
and U10788 (N_10788,N_9639,N_9272);
nor U10789 (N_10789,N_9586,N_9962);
nand U10790 (N_10790,N_9018,N_9963);
nor U10791 (N_10791,N_9028,N_9441);
or U10792 (N_10792,N_9717,N_9954);
and U10793 (N_10793,N_9397,N_9948);
nor U10794 (N_10794,N_9794,N_9908);
nand U10795 (N_10795,N_9282,N_9603);
xor U10796 (N_10796,N_9401,N_9591);
or U10797 (N_10797,N_9980,N_9975);
nand U10798 (N_10798,N_9828,N_9161);
or U10799 (N_10799,N_9446,N_9813);
xnor U10800 (N_10800,N_9215,N_9749);
nand U10801 (N_10801,N_9250,N_9030);
nor U10802 (N_10802,N_9304,N_9691);
xnor U10803 (N_10803,N_9096,N_9942);
xnor U10804 (N_10804,N_9475,N_9482);
xnor U10805 (N_10805,N_9535,N_9407);
and U10806 (N_10806,N_9383,N_9602);
nand U10807 (N_10807,N_9124,N_9016);
nand U10808 (N_10808,N_9531,N_9417);
nor U10809 (N_10809,N_9486,N_9546);
nor U10810 (N_10810,N_9272,N_9802);
nor U10811 (N_10811,N_9927,N_9137);
or U10812 (N_10812,N_9426,N_9559);
nand U10813 (N_10813,N_9325,N_9126);
nor U10814 (N_10814,N_9093,N_9690);
or U10815 (N_10815,N_9831,N_9489);
xnor U10816 (N_10816,N_9728,N_9483);
and U10817 (N_10817,N_9225,N_9920);
and U10818 (N_10818,N_9073,N_9708);
nand U10819 (N_10819,N_9084,N_9594);
nor U10820 (N_10820,N_9008,N_9880);
nand U10821 (N_10821,N_9715,N_9292);
nor U10822 (N_10822,N_9222,N_9156);
xnor U10823 (N_10823,N_9962,N_9640);
xnor U10824 (N_10824,N_9065,N_9521);
or U10825 (N_10825,N_9565,N_9667);
or U10826 (N_10826,N_9676,N_9252);
xnor U10827 (N_10827,N_9084,N_9810);
nor U10828 (N_10828,N_9498,N_9155);
nand U10829 (N_10829,N_9438,N_9932);
nor U10830 (N_10830,N_9480,N_9444);
and U10831 (N_10831,N_9394,N_9065);
xor U10832 (N_10832,N_9849,N_9829);
xor U10833 (N_10833,N_9870,N_9471);
and U10834 (N_10834,N_9630,N_9688);
and U10835 (N_10835,N_9247,N_9798);
and U10836 (N_10836,N_9806,N_9655);
or U10837 (N_10837,N_9141,N_9196);
and U10838 (N_10838,N_9452,N_9754);
or U10839 (N_10839,N_9293,N_9190);
and U10840 (N_10840,N_9106,N_9487);
xor U10841 (N_10841,N_9740,N_9500);
nor U10842 (N_10842,N_9843,N_9580);
nor U10843 (N_10843,N_9686,N_9445);
nor U10844 (N_10844,N_9202,N_9192);
and U10845 (N_10845,N_9155,N_9209);
nand U10846 (N_10846,N_9767,N_9453);
nand U10847 (N_10847,N_9512,N_9482);
nand U10848 (N_10848,N_9638,N_9619);
nand U10849 (N_10849,N_9889,N_9739);
and U10850 (N_10850,N_9689,N_9456);
nor U10851 (N_10851,N_9799,N_9864);
nand U10852 (N_10852,N_9712,N_9019);
nand U10853 (N_10853,N_9090,N_9430);
or U10854 (N_10854,N_9146,N_9284);
nand U10855 (N_10855,N_9898,N_9692);
xor U10856 (N_10856,N_9371,N_9258);
or U10857 (N_10857,N_9448,N_9264);
and U10858 (N_10858,N_9639,N_9254);
or U10859 (N_10859,N_9069,N_9779);
nand U10860 (N_10860,N_9747,N_9207);
xor U10861 (N_10861,N_9402,N_9136);
nand U10862 (N_10862,N_9837,N_9332);
nand U10863 (N_10863,N_9323,N_9605);
xor U10864 (N_10864,N_9436,N_9429);
and U10865 (N_10865,N_9953,N_9510);
xnor U10866 (N_10866,N_9205,N_9869);
or U10867 (N_10867,N_9562,N_9113);
nor U10868 (N_10868,N_9790,N_9821);
or U10869 (N_10869,N_9140,N_9129);
nand U10870 (N_10870,N_9081,N_9396);
nor U10871 (N_10871,N_9947,N_9665);
and U10872 (N_10872,N_9626,N_9519);
nand U10873 (N_10873,N_9515,N_9944);
xnor U10874 (N_10874,N_9521,N_9079);
nand U10875 (N_10875,N_9124,N_9892);
xor U10876 (N_10876,N_9947,N_9983);
or U10877 (N_10877,N_9234,N_9785);
and U10878 (N_10878,N_9309,N_9212);
xor U10879 (N_10879,N_9108,N_9928);
nand U10880 (N_10880,N_9133,N_9416);
or U10881 (N_10881,N_9684,N_9196);
nand U10882 (N_10882,N_9381,N_9386);
nand U10883 (N_10883,N_9776,N_9943);
nor U10884 (N_10884,N_9106,N_9898);
xnor U10885 (N_10885,N_9034,N_9740);
nor U10886 (N_10886,N_9581,N_9236);
or U10887 (N_10887,N_9268,N_9216);
nand U10888 (N_10888,N_9167,N_9540);
and U10889 (N_10889,N_9102,N_9604);
xor U10890 (N_10890,N_9137,N_9374);
nor U10891 (N_10891,N_9716,N_9831);
or U10892 (N_10892,N_9032,N_9178);
and U10893 (N_10893,N_9153,N_9606);
and U10894 (N_10894,N_9702,N_9511);
and U10895 (N_10895,N_9103,N_9782);
and U10896 (N_10896,N_9564,N_9044);
xnor U10897 (N_10897,N_9253,N_9194);
or U10898 (N_10898,N_9835,N_9025);
nand U10899 (N_10899,N_9227,N_9893);
nand U10900 (N_10900,N_9104,N_9429);
and U10901 (N_10901,N_9412,N_9416);
nand U10902 (N_10902,N_9512,N_9203);
or U10903 (N_10903,N_9200,N_9025);
xor U10904 (N_10904,N_9039,N_9077);
and U10905 (N_10905,N_9981,N_9025);
and U10906 (N_10906,N_9847,N_9308);
nand U10907 (N_10907,N_9046,N_9767);
xor U10908 (N_10908,N_9532,N_9283);
and U10909 (N_10909,N_9228,N_9883);
and U10910 (N_10910,N_9235,N_9382);
nor U10911 (N_10911,N_9369,N_9662);
xor U10912 (N_10912,N_9059,N_9475);
nand U10913 (N_10913,N_9185,N_9090);
nand U10914 (N_10914,N_9416,N_9651);
nor U10915 (N_10915,N_9492,N_9186);
nor U10916 (N_10916,N_9736,N_9023);
and U10917 (N_10917,N_9187,N_9348);
nor U10918 (N_10918,N_9946,N_9570);
nor U10919 (N_10919,N_9537,N_9089);
nor U10920 (N_10920,N_9853,N_9099);
and U10921 (N_10921,N_9625,N_9923);
or U10922 (N_10922,N_9131,N_9988);
xor U10923 (N_10923,N_9883,N_9617);
nor U10924 (N_10924,N_9494,N_9904);
and U10925 (N_10925,N_9304,N_9536);
xnor U10926 (N_10926,N_9472,N_9514);
nor U10927 (N_10927,N_9386,N_9618);
xor U10928 (N_10928,N_9126,N_9499);
nand U10929 (N_10929,N_9185,N_9952);
xor U10930 (N_10930,N_9776,N_9024);
xnor U10931 (N_10931,N_9052,N_9739);
or U10932 (N_10932,N_9794,N_9393);
xnor U10933 (N_10933,N_9019,N_9053);
xor U10934 (N_10934,N_9900,N_9332);
or U10935 (N_10935,N_9171,N_9945);
nor U10936 (N_10936,N_9511,N_9868);
and U10937 (N_10937,N_9153,N_9468);
nand U10938 (N_10938,N_9571,N_9852);
nor U10939 (N_10939,N_9219,N_9091);
nor U10940 (N_10940,N_9842,N_9389);
nor U10941 (N_10941,N_9878,N_9086);
xor U10942 (N_10942,N_9438,N_9876);
or U10943 (N_10943,N_9269,N_9225);
nor U10944 (N_10944,N_9032,N_9528);
nor U10945 (N_10945,N_9541,N_9683);
or U10946 (N_10946,N_9187,N_9737);
and U10947 (N_10947,N_9134,N_9786);
xnor U10948 (N_10948,N_9668,N_9021);
nand U10949 (N_10949,N_9970,N_9253);
nor U10950 (N_10950,N_9209,N_9827);
and U10951 (N_10951,N_9131,N_9307);
nor U10952 (N_10952,N_9006,N_9930);
xnor U10953 (N_10953,N_9828,N_9904);
xor U10954 (N_10954,N_9829,N_9617);
nand U10955 (N_10955,N_9893,N_9076);
nor U10956 (N_10956,N_9808,N_9366);
nand U10957 (N_10957,N_9881,N_9710);
or U10958 (N_10958,N_9853,N_9045);
nor U10959 (N_10959,N_9821,N_9960);
and U10960 (N_10960,N_9214,N_9326);
nor U10961 (N_10961,N_9534,N_9269);
or U10962 (N_10962,N_9075,N_9830);
nand U10963 (N_10963,N_9283,N_9806);
and U10964 (N_10964,N_9831,N_9496);
nor U10965 (N_10965,N_9171,N_9767);
xor U10966 (N_10966,N_9207,N_9777);
xor U10967 (N_10967,N_9346,N_9722);
or U10968 (N_10968,N_9295,N_9913);
nor U10969 (N_10969,N_9730,N_9702);
or U10970 (N_10970,N_9780,N_9515);
nor U10971 (N_10971,N_9177,N_9346);
nor U10972 (N_10972,N_9983,N_9321);
or U10973 (N_10973,N_9712,N_9068);
nor U10974 (N_10974,N_9950,N_9576);
or U10975 (N_10975,N_9640,N_9468);
nand U10976 (N_10976,N_9265,N_9196);
and U10977 (N_10977,N_9555,N_9421);
or U10978 (N_10978,N_9425,N_9215);
or U10979 (N_10979,N_9100,N_9336);
nand U10980 (N_10980,N_9841,N_9511);
and U10981 (N_10981,N_9221,N_9016);
nand U10982 (N_10982,N_9772,N_9667);
nor U10983 (N_10983,N_9192,N_9764);
xnor U10984 (N_10984,N_9078,N_9036);
or U10985 (N_10985,N_9990,N_9477);
and U10986 (N_10986,N_9999,N_9202);
nor U10987 (N_10987,N_9715,N_9124);
nand U10988 (N_10988,N_9848,N_9770);
nor U10989 (N_10989,N_9970,N_9641);
and U10990 (N_10990,N_9186,N_9325);
nand U10991 (N_10991,N_9616,N_9171);
or U10992 (N_10992,N_9299,N_9268);
xor U10993 (N_10993,N_9850,N_9445);
and U10994 (N_10994,N_9958,N_9906);
or U10995 (N_10995,N_9454,N_9347);
nand U10996 (N_10996,N_9783,N_9354);
or U10997 (N_10997,N_9095,N_9637);
xnor U10998 (N_10998,N_9198,N_9240);
and U10999 (N_10999,N_9322,N_9312);
and U11000 (N_11000,N_10356,N_10892);
nor U11001 (N_11001,N_10779,N_10435);
nand U11002 (N_11002,N_10776,N_10222);
nor U11003 (N_11003,N_10808,N_10104);
nor U11004 (N_11004,N_10291,N_10681);
and U11005 (N_11005,N_10741,N_10313);
nand U11006 (N_11006,N_10704,N_10031);
and U11007 (N_11007,N_10516,N_10372);
and U11008 (N_11008,N_10861,N_10765);
or U11009 (N_11009,N_10973,N_10209);
nand U11010 (N_11010,N_10803,N_10889);
xor U11011 (N_11011,N_10033,N_10826);
and U11012 (N_11012,N_10669,N_10598);
and U11013 (N_11013,N_10865,N_10307);
nor U11014 (N_11014,N_10950,N_10081);
xor U11015 (N_11015,N_10075,N_10205);
xnor U11016 (N_11016,N_10683,N_10721);
nand U11017 (N_11017,N_10623,N_10488);
and U11018 (N_11018,N_10627,N_10187);
xnor U11019 (N_11019,N_10891,N_10880);
nor U11020 (N_11020,N_10278,N_10596);
nor U11021 (N_11021,N_10367,N_10299);
nand U11022 (N_11022,N_10966,N_10628);
xnor U11023 (N_11023,N_10643,N_10399);
and U11024 (N_11024,N_10362,N_10662);
nor U11025 (N_11025,N_10847,N_10758);
or U11026 (N_11026,N_10613,N_10247);
and U11027 (N_11027,N_10170,N_10018);
or U11028 (N_11028,N_10505,N_10998);
nor U11029 (N_11029,N_10857,N_10084);
or U11030 (N_11030,N_10452,N_10798);
xnor U11031 (N_11031,N_10635,N_10941);
nand U11032 (N_11032,N_10746,N_10942);
or U11033 (N_11033,N_10058,N_10498);
and U11034 (N_11034,N_10897,N_10048);
and U11035 (N_11035,N_10640,N_10417);
nand U11036 (N_11036,N_10109,N_10925);
and U11037 (N_11037,N_10337,N_10771);
nand U11038 (N_11038,N_10426,N_10010);
or U11039 (N_11039,N_10896,N_10905);
and U11040 (N_11040,N_10605,N_10862);
nand U11041 (N_11041,N_10361,N_10547);
and U11042 (N_11042,N_10714,N_10402);
xnor U11043 (N_11043,N_10983,N_10873);
xnor U11044 (N_11044,N_10166,N_10700);
xnor U11045 (N_11045,N_10702,N_10445);
nand U11046 (N_11046,N_10607,N_10305);
xor U11047 (N_11047,N_10843,N_10701);
and U11048 (N_11048,N_10322,N_10929);
and U11049 (N_11049,N_10759,N_10988);
or U11050 (N_11050,N_10196,N_10118);
or U11051 (N_11051,N_10267,N_10347);
and U11052 (N_11052,N_10859,N_10723);
nand U11053 (N_11053,N_10316,N_10917);
nand U11054 (N_11054,N_10441,N_10673);
or U11055 (N_11055,N_10540,N_10154);
or U11056 (N_11056,N_10645,N_10436);
or U11057 (N_11057,N_10391,N_10223);
nand U11058 (N_11058,N_10342,N_10691);
nor U11059 (N_11059,N_10858,N_10649);
or U11060 (N_11060,N_10918,N_10215);
nand U11061 (N_11061,N_10920,N_10935);
or U11062 (N_11062,N_10056,N_10993);
nor U11063 (N_11063,N_10655,N_10024);
nor U11064 (N_11064,N_10901,N_10325);
or U11065 (N_11065,N_10801,N_10012);
nand U11066 (N_11066,N_10284,N_10338);
and U11067 (N_11067,N_10742,N_10087);
nor U11068 (N_11068,N_10981,N_10586);
xnor U11069 (N_11069,N_10424,N_10898);
nor U11070 (N_11070,N_10092,N_10448);
xor U11071 (N_11071,N_10921,N_10471);
and U11072 (N_11072,N_10678,N_10133);
xor U11073 (N_11073,N_10478,N_10997);
or U11074 (N_11074,N_10199,N_10616);
nand U11075 (N_11075,N_10239,N_10834);
nor U11076 (N_11076,N_10444,N_10829);
and U11077 (N_11077,N_10513,N_10579);
nor U11078 (N_11078,N_10725,N_10593);
nor U11079 (N_11079,N_10783,N_10972);
nor U11080 (N_11080,N_10396,N_10355);
or U11081 (N_11081,N_10962,N_10153);
nand U11082 (N_11082,N_10894,N_10615);
nor U11083 (N_11083,N_10777,N_10768);
or U11084 (N_11084,N_10549,N_10612);
or U11085 (N_11085,N_10289,N_10556);
or U11086 (N_11086,N_10413,N_10831);
nor U11087 (N_11087,N_10094,N_10242);
xnor U11088 (N_11088,N_10183,N_10521);
nor U11089 (N_11089,N_10403,N_10856);
nor U11090 (N_11090,N_10088,N_10955);
and U11091 (N_11091,N_10431,N_10482);
or U11092 (N_11092,N_10527,N_10314);
and U11093 (N_11093,N_10381,N_10667);
or U11094 (N_11094,N_10814,N_10161);
and U11095 (N_11095,N_10657,N_10158);
or U11096 (N_11096,N_10195,N_10766);
and U11097 (N_11097,N_10273,N_10308);
or U11098 (N_11098,N_10528,N_10047);
xnor U11099 (N_11099,N_10134,N_10648);
xor U11100 (N_11100,N_10440,N_10071);
nand U11101 (N_11101,N_10564,N_10220);
xor U11102 (N_11102,N_10975,N_10735);
xor U11103 (N_11103,N_10587,N_10760);
nand U11104 (N_11104,N_10739,N_10752);
nand U11105 (N_11105,N_10636,N_10016);
and U11106 (N_11106,N_10184,N_10690);
or U11107 (N_11107,N_10099,N_10585);
nor U11108 (N_11108,N_10511,N_10198);
xor U11109 (N_11109,N_10544,N_10588);
nand U11110 (N_11110,N_10869,N_10508);
and U11111 (N_11111,N_10959,N_10475);
and U11112 (N_11112,N_10692,N_10778);
and U11113 (N_11113,N_10619,N_10686);
xnor U11114 (N_11114,N_10874,N_10604);
xnor U11115 (N_11115,N_10825,N_10668);
nand U11116 (N_11116,N_10189,N_10115);
xnor U11117 (N_11117,N_10346,N_10583);
nor U11118 (N_11118,N_10025,N_10282);
nand U11119 (N_11119,N_10978,N_10989);
and U11120 (N_11120,N_10306,N_10866);
xor U11121 (N_11121,N_10083,N_10233);
xor U11122 (N_11122,N_10519,N_10698);
nor U11123 (N_11123,N_10117,N_10884);
nor U11124 (N_11124,N_10310,N_10332);
and U11125 (N_11125,N_10523,N_10204);
nand U11126 (N_11126,N_10947,N_10312);
or U11127 (N_11127,N_10142,N_10007);
nor U11128 (N_11128,N_10868,N_10823);
nand U11129 (N_11129,N_10731,N_10864);
nor U11130 (N_11130,N_10621,N_10703);
xnor U11131 (N_11131,N_10499,N_10026);
xor U11132 (N_11132,N_10952,N_10433);
nand U11133 (N_11133,N_10986,N_10437);
nand U11134 (N_11134,N_10096,N_10762);
or U11135 (N_11135,N_10535,N_10729);
xor U11136 (N_11136,N_10474,N_10639);
or U11137 (N_11137,N_10509,N_10589);
and U11138 (N_11138,N_10138,N_10990);
and U11139 (N_11139,N_10736,N_10984);
and U11140 (N_11140,N_10939,N_10178);
and U11141 (N_11141,N_10366,N_10524);
nand U11142 (N_11142,N_10795,N_10237);
and U11143 (N_11143,N_10781,N_10371);
xnor U11144 (N_11144,N_10129,N_10934);
nand U11145 (N_11145,N_10663,N_10713);
or U11146 (N_11146,N_10182,N_10875);
nor U11147 (N_11147,N_10911,N_10507);
nand U11148 (N_11148,N_10915,N_10961);
nor U11149 (N_11149,N_10270,N_10642);
xor U11150 (N_11150,N_10442,N_10542);
nand U11151 (N_11151,N_10852,N_10468);
xnor U11152 (N_11152,N_10622,N_10680);
and U11153 (N_11153,N_10201,N_10095);
xnor U11154 (N_11154,N_10343,N_10423);
and U11155 (N_11155,N_10971,N_10525);
or U11156 (N_11156,N_10149,N_10331);
and U11157 (N_11157,N_10531,N_10467);
nand U11158 (N_11158,N_10590,N_10878);
nor U11159 (N_11159,N_10719,N_10745);
nand U11160 (N_11160,N_10345,N_10545);
and U11161 (N_11161,N_10334,N_10839);
nor U11162 (N_11162,N_10206,N_10851);
and U11163 (N_11163,N_10926,N_10824);
nor U11164 (N_11164,N_10159,N_10999);
nand U11165 (N_11165,N_10463,N_10785);
and U11166 (N_11166,N_10877,N_10890);
nor U11167 (N_11167,N_10582,N_10994);
or U11168 (N_11168,N_10936,N_10810);
and U11169 (N_11169,N_10481,N_10430);
or U11170 (N_11170,N_10395,N_10541);
xnor U11171 (N_11171,N_10809,N_10753);
nand U11172 (N_11172,N_10539,N_10529);
nor U11173 (N_11173,N_10695,N_10817);
xnor U11174 (N_11174,N_10820,N_10318);
nand U11175 (N_11175,N_10283,N_10124);
nor U11176 (N_11176,N_10022,N_10098);
xor U11177 (N_11177,N_10451,N_10899);
nor U11178 (N_11178,N_10784,N_10571);
and U11179 (N_11179,N_10837,N_10110);
and U11180 (N_11180,N_10888,N_10949);
nand U11181 (N_11181,N_10344,N_10948);
and U11182 (N_11182,N_10756,N_10264);
and U11183 (N_11183,N_10211,N_10793);
nor U11184 (N_11184,N_10553,N_10062);
and U11185 (N_11185,N_10532,N_10718);
xnor U11186 (N_11186,N_10485,N_10418);
xor U11187 (N_11187,N_10606,N_10689);
and U11188 (N_11188,N_10560,N_10614);
xor U11189 (N_11189,N_10907,N_10840);
and U11190 (N_11190,N_10828,N_10080);
xnor U11191 (N_11191,N_10072,N_10646);
or U11192 (N_11192,N_10375,N_10536);
nor U11193 (N_11193,N_10450,N_10434);
or U11194 (N_11194,N_10594,N_10764);
and U11195 (N_11195,N_10102,N_10429);
and U11196 (N_11196,N_10015,N_10849);
and U11197 (N_11197,N_10956,N_10122);
and U11198 (N_11198,N_10459,N_10165);
and U11199 (N_11199,N_10716,N_10854);
or U11200 (N_11200,N_10044,N_10162);
and U11201 (N_11201,N_10664,N_10744);
or U11202 (N_11202,N_10548,N_10050);
xnor U11203 (N_11203,N_10288,N_10243);
xor U11204 (N_11204,N_10093,N_10512);
nor U11205 (N_11205,N_10155,N_10738);
nor U11206 (N_11206,N_10557,N_10086);
nand U11207 (N_11207,N_10169,N_10705);
and U11208 (N_11208,N_10136,N_10480);
xnor U11209 (N_11209,N_10913,N_10382);
nand U11210 (N_11210,N_10775,N_10597);
or U11211 (N_11211,N_10782,N_10401);
nand U11212 (N_11212,N_10991,N_10107);
xor U11213 (N_11213,N_10422,N_10797);
nand U11214 (N_11214,N_10324,N_10041);
nand U11215 (N_11215,N_10443,N_10937);
xnor U11216 (N_11216,N_10002,N_10833);
or U11217 (N_11217,N_10246,N_10131);
nand U11218 (N_11218,N_10600,N_10309);
and U11219 (N_11219,N_10301,N_10794);
nor U11220 (N_11220,N_10232,N_10295);
or U11221 (N_11221,N_10364,N_10427);
xnor U11222 (N_11222,N_10748,N_10023);
xor U11223 (N_11223,N_10303,N_10383);
and U11224 (N_11224,N_10287,N_10836);
and U11225 (N_11225,N_10787,N_10321);
xnor U11226 (N_11226,N_10171,N_10398);
and U11227 (N_11227,N_10626,N_10145);
and U11228 (N_11228,N_10221,N_10658);
nand U11229 (N_11229,N_10146,N_10039);
nor U11230 (N_11230,N_10518,N_10005);
nor U11231 (N_11231,N_10876,N_10326);
and U11232 (N_11232,N_10976,N_10908);
and U11233 (N_11233,N_10329,N_10164);
nor U11234 (N_11234,N_10057,N_10271);
and U11235 (N_11235,N_10176,N_10733);
or U11236 (N_11236,N_10009,N_10773);
or U11237 (N_11237,N_10500,N_10965);
and U11238 (N_11238,N_10281,N_10365);
and U11239 (N_11239,N_10051,N_10750);
nor U11240 (N_11240,N_10656,N_10200);
and U11241 (N_11241,N_10150,N_10708);
and U11242 (N_11242,N_10818,N_10101);
and U11243 (N_11243,N_10408,N_10315);
or U11244 (N_11244,N_10144,N_10453);
or U11245 (N_11245,N_10254,N_10035);
nor U11246 (N_11246,N_10757,N_10572);
nor U11247 (N_11247,N_10811,N_10252);
nand U11248 (N_11248,N_10327,N_10363);
xnor U11249 (N_11249,N_10727,N_10257);
nand U11250 (N_11250,N_10933,N_10774);
nand U11251 (N_11251,N_10938,N_10931);
nand U11252 (N_11252,N_10796,N_10819);
and U11253 (N_11253,N_10493,N_10052);
nor U11254 (N_11254,N_10106,N_10812);
xnor U11255 (N_11255,N_10791,N_10870);
xor U11256 (N_11256,N_10838,N_10651);
and U11257 (N_11257,N_10245,N_10620);
xor U11258 (N_11258,N_10230,N_10479);
nor U11259 (N_11259,N_10378,N_10624);
and U11260 (N_11260,N_10603,N_10294);
and U11261 (N_11261,N_10394,N_10379);
nand U11262 (N_11262,N_10419,N_10581);
and U11263 (N_11263,N_10555,N_10385);
nand U11264 (N_11264,N_10428,N_10489);
nand U11265 (N_11265,N_10097,N_10353);
nand U11266 (N_11266,N_10652,N_10190);
nand U11267 (N_11267,N_10415,N_10001);
and U11268 (N_11268,N_10567,N_10123);
xnor U11269 (N_11269,N_10064,N_10317);
xnor U11270 (N_11270,N_10932,N_10715);
or U11271 (N_11271,N_10261,N_10543);
or U11272 (N_11272,N_10188,N_10276);
and U11273 (N_11273,N_10660,N_10789);
and U11274 (N_11274,N_10711,N_10534);
and U11275 (N_11275,N_10611,N_10277);
nor U11276 (N_11276,N_10388,N_10494);
or U11277 (N_11277,N_10054,N_10397);
or U11278 (N_11278,N_10248,N_10883);
nand U11279 (N_11279,N_10767,N_10393);
xor U11280 (N_11280,N_10665,N_10653);
or U11281 (N_11281,N_10250,N_10004);
or U11282 (N_11282,N_10634,N_10706);
and U11283 (N_11283,N_10216,N_10006);
xor U11284 (N_11284,N_10595,N_10224);
nand U11285 (N_11285,N_10017,N_10732);
and U11286 (N_11286,N_10238,N_10465);
or U11287 (N_11287,N_10670,N_10377);
xnor U11288 (N_11288,N_10410,N_10279);
and U11289 (N_11289,N_10416,N_10800);
and U11290 (N_11290,N_10514,N_10568);
nand U11291 (N_11291,N_10501,N_10292);
xor U11292 (N_11292,N_10483,N_10061);
xor U11293 (N_11293,N_10761,N_10763);
nor U11294 (N_11294,N_10815,N_10684);
and U11295 (N_11295,N_10260,N_10964);
nand U11296 (N_11296,N_10747,N_10807);
nor U11297 (N_11297,N_10561,N_10091);
or U11298 (N_11298,N_10192,N_10404);
nor U11299 (N_11299,N_10042,N_10788);
nor U11300 (N_11300,N_10871,N_10349);
nand U11301 (N_11301,N_10040,N_10280);
nor U11302 (N_11302,N_10241,N_10996);
or U11303 (N_11303,N_10191,N_10546);
nand U11304 (N_11304,N_10637,N_10259);
nor U11305 (N_11305,N_10855,N_10275);
nand U11306 (N_11306,N_10618,N_10286);
xor U11307 (N_11307,N_10141,N_10882);
xor U11308 (N_11308,N_10341,N_10333);
and U11309 (N_11309,N_10258,N_10982);
xnor U11310 (N_11310,N_10910,N_10210);
nor U11311 (N_11311,N_10358,N_10181);
or U11312 (N_11312,N_10390,N_10699);
nand U11313 (N_11313,N_10940,N_10510);
nor U11314 (N_11314,N_10841,N_10272);
and U11315 (N_11315,N_10219,N_10687);
nand U11316 (N_11316,N_10520,N_10740);
nor U11317 (N_11317,N_10672,N_10806);
or U11318 (N_11318,N_10172,N_10887);
xnor U11319 (N_11319,N_10617,N_10522);
nor U11320 (N_11320,N_10231,N_10454);
xor U11321 (N_11321,N_10987,N_10339);
nand U11322 (N_11322,N_10486,N_10013);
nand U11323 (N_11323,N_10625,N_10772);
and U11324 (N_11324,N_10816,N_10458);
and U11325 (N_11325,N_10008,N_10256);
xor U11326 (N_11326,N_10848,N_10304);
or U11327 (N_11327,N_10786,N_10944);
and U11328 (N_11328,N_10710,N_10266);
nand U11329 (N_11329,N_10469,N_10405);
nand U11330 (N_11330,N_10923,N_10032);
nor U11331 (N_11331,N_10575,N_10174);
and U11332 (N_11332,N_10420,N_10328);
or U11333 (N_11333,N_10677,N_10111);
xnor U11334 (N_11334,N_10609,N_10078);
and U11335 (N_11335,N_10974,N_10592);
nand U11336 (N_11336,N_10969,N_10085);
and U11337 (N_11337,N_10226,N_10116);
xnor U11338 (N_11338,N_10335,N_10336);
nor U11339 (N_11339,N_10654,N_10455);
nand U11340 (N_11340,N_10157,N_10297);
xor U11341 (N_11341,N_10053,N_10886);
nand U11342 (N_11342,N_10409,N_10090);
nor U11343 (N_11343,N_10599,N_10067);
nand U11344 (N_11344,N_10065,N_10502);
nand U11345 (N_11345,N_10631,N_10068);
and U11346 (N_11346,N_10202,N_10160);
xnor U11347 (N_11347,N_10922,N_10707);
and U11348 (N_11348,N_10813,N_10574);
nor U11349 (N_11349,N_10506,N_10113);
nor U11350 (N_11350,N_10565,N_10135);
xnor U11351 (N_11351,N_10537,N_10927);
nor U11352 (N_11352,N_10967,N_10456);
xor U11353 (N_11353,N_10439,N_10844);
nor U11354 (N_11354,N_10446,N_10406);
or U11355 (N_11355,N_10311,N_10186);
nand U11356 (N_11356,N_10722,N_10960);
xnor U11357 (N_11357,N_10212,N_10608);
and U11358 (N_11358,N_10491,N_10951);
xnor U11359 (N_11359,N_10832,N_10082);
or U11360 (N_11360,N_10457,N_10676);
nor U11361 (N_11361,N_10487,N_10881);
nor U11362 (N_11362,N_10755,N_10156);
nand U11363 (N_11363,N_10029,N_10958);
nor U11364 (N_11364,N_10352,N_10591);
nand U11365 (N_11365,N_10728,N_10128);
and U11366 (N_11366,N_10197,N_10559);
nor U11367 (N_11367,N_10217,N_10464);
xnor U11368 (N_11368,N_10472,N_10139);
nor U11369 (N_11369,N_10830,N_10726);
or U11370 (N_11370,N_10515,N_10214);
or U11371 (N_11371,N_10251,N_10244);
xnor U11372 (N_11372,N_10126,N_10754);
or U11373 (N_11373,N_10235,N_10089);
nand U11374 (N_11374,N_10028,N_10517);
or U11375 (N_11375,N_10980,N_10447);
nand U11376 (N_11376,N_10953,N_10916);
xor U11377 (N_11377,N_10132,N_10885);
nor U11378 (N_11378,N_10253,N_10661);
xor U11379 (N_11379,N_10249,N_10063);
nor U11380 (N_11380,N_10985,N_10685);
and U11381 (N_11381,N_10380,N_10688);
nor U11382 (N_11382,N_10368,N_10140);
and U11383 (N_11383,N_10749,N_10957);
and U11384 (N_11384,N_10853,N_10632);
and U11385 (N_11385,N_10152,N_10225);
or U11386 (N_11386,N_10914,N_10148);
xnor U11387 (N_11387,N_10357,N_10100);
or U11388 (N_11388,N_10046,N_10376);
nand U11389 (N_11389,N_10822,N_10737);
and U11390 (N_11390,N_10979,N_10584);
or U11391 (N_11391,N_10895,N_10879);
or U11392 (N_11392,N_10438,N_10302);
nand U11393 (N_11393,N_10055,N_10717);
nor U11394 (N_11394,N_10943,N_10580);
nor U11395 (N_11395,N_10751,N_10400);
or U11396 (N_11396,N_10842,N_10769);
nor U11397 (N_11397,N_10340,N_10030);
or U11398 (N_11398,N_10629,N_10666);
nand U11399 (N_11399,N_10019,N_10867);
nor U11400 (N_11400,N_10633,N_10179);
xor U11401 (N_11401,N_10641,N_10108);
xor U11402 (N_11402,N_10790,N_10893);
or U11403 (N_11403,N_10079,N_10460);
nand U11404 (N_11404,N_10712,N_10240);
nand U11405 (N_11405,N_10076,N_10263);
or U11406 (N_11406,N_10647,N_10412);
and U11407 (N_11407,N_10180,N_10177);
nand U11408 (N_11408,N_10992,N_10168);
nor U11409 (N_11409,N_10504,N_10551);
xnor U11410 (N_11410,N_10709,N_10021);
nor U11411 (N_11411,N_10255,N_10954);
nor U11412 (N_11412,N_10462,N_10285);
or U11413 (N_11413,N_10218,N_10554);
xnor U11414 (N_11414,N_10425,N_10274);
nor U11415 (N_11415,N_10473,N_10034);
nor U11416 (N_11416,N_10414,N_10696);
nor U11417 (N_11417,N_10730,N_10373);
and U11418 (N_11418,N_10569,N_10003);
and U11419 (N_11419,N_10036,N_10120);
xnor U11420 (N_11420,N_10203,N_10675);
and U11421 (N_11421,N_10850,N_10492);
nor U11422 (N_11422,N_10213,N_10038);
xnor U11423 (N_11423,N_10821,N_10558);
and U11424 (N_11424,N_10384,N_10573);
nor U11425 (N_11425,N_10070,N_10900);
or U11426 (N_11426,N_10290,N_10490);
xnor U11427 (N_11427,N_10477,N_10112);
nand U11428 (N_11428,N_10578,N_10392);
and U11429 (N_11429,N_10930,N_10105);
xor U11430 (N_11430,N_10977,N_10293);
nand U11431 (N_11431,N_10027,N_10127);
nor U11432 (N_11432,N_10644,N_10300);
and U11433 (N_11433,N_10638,N_10296);
nor U11434 (N_11434,N_10682,N_10659);
and U11435 (N_11435,N_10137,N_10693);
and U11436 (N_11436,N_10835,N_10049);
nand U11437 (N_11437,N_10119,N_10562);
or U11438 (N_11438,N_10011,N_10073);
nor U11439 (N_11439,N_10043,N_10601);
or U11440 (N_11440,N_10208,N_10014);
or U11441 (N_11441,N_10602,N_10348);
and U11442 (N_11442,N_10130,N_10234);
nand U11443 (N_11443,N_10369,N_10946);
nor U11444 (N_11444,N_10432,N_10185);
nor U11445 (N_11445,N_10799,N_10163);
xnor U11446 (N_11446,N_10566,N_10470);
nor U11447 (N_11447,N_10912,N_10354);
or U11448 (N_11448,N_10194,N_10904);
nand U11449 (N_11449,N_10863,N_10526);
xor U11450 (N_11450,N_10674,N_10845);
nor U11451 (N_11451,N_10229,N_10963);
or U11452 (N_11452,N_10792,N_10533);
nand U11453 (N_11453,N_10147,N_10167);
nand U11454 (N_11454,N_10802,N_10805);
or U11455 (N_11455,N_10919,N_10968);
nand U11456 (N_11456,N_10538,N_10497);
nand U11457 (N_11457,N_10151,N_10630);
and U11458 (N_11458,N_10743,N_10476);
nand U11459 (N_11459,N_10370,N_10360);
nand U11460 (N_11460,N_10466,N_10449);
xnor U11461 (N_11461,N_10671,N_10679);
xor U11462 (N_11462,N_10359,N_10020);
and U11463 (N_11463,N_10909,N_10389);
nor U11464 (N_11464,N_10060,N_10970);
nand U11465 (N_11465,N_10804,N_10563);
nand U11466 (N_11466,N_10207,N_10386);
nand U11467 (N_11467,N_10236,N_10411);
and U11468 (N_11468,N_10262,N_10694);
nor U11469 (N_11469,N_10143,N_10577);
xor U11470 (N_11470,N_10265,N_10902);
xnor U11471 (N_11471,N_10484,N_10069);
and U11472 (N_11472,N_10374,N_10350);
nand U11473 (N_11473,N_10125,N_10720);
nor U11474 (N_11474,N_10114,N_10903);
xnor U11475 (N_11475,N_10103,N_10827);
xor U11476 (N_11476,N_10330,N_10724);
nand U11477 (N_11477,N_10066,N_10323);
nand U11478 (N_11478,N_10860,N_10037);
nor U11479 (N_11479,N_10530,N_10077);
or U11480 (N_11480,N_10461,N_10846);
xnor U11481 (N_11481,N_10495,N_10074);
and U11482 (N_11482,N_10610,N_10421);
nand U11483 (N_11483,N_10228,N_10503);
xnor U11484 (N_11484,N_10570,N_10121);
and U11485 (N_11485,N_10872,N_10387);
nor U11486 (N_11486,N_10059,N_10407);
nor U11487 (N_11487,N_10268,N_10924);
xnor U11488 (N_11488,N_10780,N_10298);
nand U11489 (N_11489,N_10650,N_10576);
or U11490 (N_11490,N_10928,N_10906);
xnor U11491 (N_11491,N_10175,N_10552);
nand U11492 (N_11492,N_10770,N_10045);
and U11493 (N_11493,N_10320,N_10496);
or U11494 (N_11494,N_10193,N_10995);
or U11495 (N_11495,N_10734,N_10000);
or U11496 (N_11496,N_10697,N_10550);
nor U11497 (N_11497,N_10945,N_10351);
nand U11498 (N_11498,N_10173,N_10227);
and U11499 (N_11499,N_10319,N_10269);
nor U11500 (N_11500,N_10558,N_10741);
nor U11501 (N_11501,N_10879,N_10555);
and U11502 (N_11502,N_10149,N_10733);
nand U11503 (N_11503,N_10427,N_10980);
nor U11504 (N_11504,N_10723,N_10799);
and U11505 (N_11505,N_10349,N_10380);
or U11506 (N_11506,N_10976,N_10426);
and U11507 (N_11507,N_10640,N_10050);
or U11508 (N_11508,N_10144,N_10129);
nor U11509 (N_11509,N_10594,N_10607);
or U11510 (N_11510,N_10183,N_10482);
xor U11511 (N_11511,N_10875,N_10472);
or U11512 (N_11512,N_10371,N_10531);
or U11513 (N_11513,N_10412,N_10778);
and U11514 (N_11514,N_10799,N_10589);
nand U11515 (N_11515,N_10459,N_10302);
nand U11516 (N_11516,N_10460,N_10450);
xor U11517 (N_11517,N_10508,N_10012);
or U11518 (N_11518,N_10082,N_10727);
nor U11519 (N_11519,N_10197,N_10443);
nor U11520 (N_11520,N_10989,N_10590);
xnor U11521 (N_11521,N_10940,N_10106);
nand U11522 (N_11522,N_10587,N_10726);
nor U11523 (N_11523,N_10087,N_10887);
nand U11524 (N_11524,N_10774,N_10443);
xnor U11525 (N_11525,N_10712,N_10838);
nor U11526 (N_11526,N_10136,N_10105);
nand U11527 (N_11527,N_10331,N_10827);
and U11528 (N_11528,N_10142,N_10037);
or U11529 (N_11529,N_10641,N_10295);
nand U11530 (N_11530,N_10069,N_10050);
nand U11531 (N_11531,N_10947,N_10713);
and U11532 (N_11532,N_10596,N_10886);
or U11533 (N_11533,N_10072,N_10215);
or U11534 (N_11534,N_10232,N_10723);
xor U11535 (N_11535,N_10613,N_10145);
xnor U11536 (N_11536,N_10620,N_10970);
nor U11537 (N_11537,N_10804,N_10075);
or U11538 (N_11538,N_10214,N_10862);
and U11539 (N_11539,N_10700,N_10720);
nor U11540 (N_11540,N_10880,N_10710);
and U11541 (N_11541,N_10683,N_10572);
nor U11542 (N_11542,N_10819,N_10179);
and U11543 (N_11543,N_10554,N_10881);
nor U11544 (N_11544,N_10707,N_10534);
nor U11545 (N_11545,N_10450,N_10363);
nor U11546 (N_11546,N_10968,N_10709);
nand U11547 (N_11547,N_10275,N_10653);
nor U11548 (N_11548,N_10506,N_10465);
or U11549 (N_11549,N_10874,N_10184);
xnor U11550 (N_11550,N_10565,N_10553);
and U11551 (N_11551,N_10616,N_10983);
or U11552 (N_11552,N_10484,N_10220);
or U11553 (N_11553,N_10701,N_10322);
and U11554 (N_11554,N_10376,N_10753);
or U11555 (N_11555,N_10275,N_10122);
or U11556 (N_11556,N_10260,N_10350);
or U11557 (N_11557,N_10238,N_10033);
and U11558 (N_11558,N_10315,N_10570);
and U11559 (N_11559,N_10931,N_10584);
and U11560 (N_11560,N_10287,N_10293);
nand U11561 (N_11561,N_10475,N_10061);
or U11562 (N_11562,N_10893,N_10236);
and U11563 (N_11563,N_10007,N_10054);
nand U11564 (N_11564,N_10648,N_10966);
nand U11565 (N_11565,N_10192,N_10248);
nand U11566 (N_11566,N_10835,N_10005);
xor U11567 (N_11567,N_10340,N_10111);
and U11568 (N_11568,N_10929,N_10757);
nor U11569 (N_11569,N_10884,N_10316);
xor U11570 (N_11570,N_10831,N_10609);
or U11571 (N_11571,N_10155,N_10943);
nand U11572 (N_11572,N_10620,N_10562);
xnor U11573 (N_11573,N_10990,N_10675);
xor U11574 (N_11574,N_10854,N_10548);
xnor U11575 (N_11575,N_10068,N_10454);
nor U11576 (N_11576,N_10628,N_10379);
or U11577 (N_11577,N_10057,N_10124);
xor U11578 (N_11578,N_10503,N_10944);
nand U11579 (N_11579,N_10318,N_10691);
nand U11580 (N_11580,N_10278,N_10365);
nor U11581 (N_11581,N_10888,N_10748);
nand U11582 (N_11582,N_10283,N_10099);
nor U11583 (N_11583,N_10797,N_10566);
xor U11584 (N_11584,N_10708,N_10594);
and U11585 (N_11585,N_10529,N_10844);
and U11586 (N_11586,N_10351,N_10308);
nand U11587 (N_11587,N_10978,N_10162);
xnor U11588 (N_11588,N_10014,N_10388);
nand U11589 (N_11589,N_10021,N_10044);
nand U11590 (N_11590,N_10773,N_10265);
nand U11591 (N_11591,N_10636,N_10138);
nor U11592 (N_11592,N_10587,N_10262);
nor U11593 (N_11593,N_10335,N_10074);
xnor U11594 (N_11594,N_10841,N_10355);
nand U11595 (N_11595,N_10499,N_10363);
or U11596 (N_11596,N_10001,N_10806);
nor U11597 (N_11597,N_10947,N_10213);
xor U11598 (N_11598,N_10780,N_10047);
xnor U11599 (N_11599,N_10097,N_10210);
nor U11600 (N_11600,N_10548,N_10468);
nand U11601 (N_11601,N_10406,N_10404);
and U11602 (N_11602,N_10443,N_10426);
or U11603 (N_11603,N_10223,N_10876);
xnor U11604 (N_11604,N_10636,N_10677);
xnor U11605 (N_11605,N_10227,N_10016);
or U11606 (N_11606,N_10828,N_10062);
xnor U11607 (N_11607,N_10487,N_10977);
and U11608 (N_11608,N_10108,N_10159);
nand U11609 (N_11609,N_10714,N_10397);
nand U11610 (N_11610,N_10612,N_10365);
and U11611 (N_11611,N_10577,N_10964);
or U11612 (N_11612,N_10061,N_10910);
and U11613 (N_11613,N_10330,N_10451);
nand U11614 (N_11614,N_10274,N_10542);
nor U11615 (N_11615,N_10583,N_10414);
nor U11616 (N_11616,N_10594,N_10042);
or U11617 (N_11617,N_10114,N_10588);
nand U11618 (N_11618,N_10159,N_10225);
nand U11619 (N_11619,N_10498,N_10500);
xnor U11620 (N_11620,N_10161,N_10323);
nand U11621 (N_11621,N_10589,N_10124);
nand U11622 (N_11622,N_10378,N_10530);
nand U11623 (N_11623,N_10440,N_10794);
and U11624 (N_11624,N_10489,N_10996);
nand U11625 (N_11625,N_10355,N_10444);
and U11626 (N_11626,N_10617,N_10327);
nor U11627 (N_11627,N_10038,N_10526);
xor U11628 (N_11628,N_10987,N_10107);
nand U11629 (N_11629,N_10901,N_10696);
nor U11630 (N_11630,N_10177,N_10774);
nand U11631 (N_11631,N_10652,N_10494);
or U11632 (N_11632,N_10745,N_10601);
nand U11633 (N_11633,N_10026,N_10382);
nand U11634 (N_11634,N_10447,N_10876);
and U11635 (N_11635,N_10400,N_10639);
nor U11636 (N_11636,N_10783,N_10651);
nor U11637 (N_11637,N_10727,N_10332);
xor U11638 (N_11638,N_10261,N_10968);
nand U11639 (N_11639,N_10397,N_10239);
nand U11640 (N_11640,N_10950,N_10369);
xnor U11641 (N_11641,N_10347,N_10696);
or U11642 (N_11642,N_10350,N_10795);
nor U11643 (N_11643,N_10859,N_10861);
nor U11644 (N_11644,N_10896,N_10713);
nor U11645 (N_11645,N_10704,N_10915);
nor U11646 (N_11646,N_10897,N_10832);
or U11647 (N_11647,N_10016,N_10719);
xor U11648 (N_11648,N_10408,N_10531);
xnor U11649 (N_11649,N_10787,N_10613);
xnor U11650 (N_11650,N_10593,N_10039);
or U11651 (N_11651,N_10389,N_10952);
and U11652 (N_11652,N_10850,N_10673);
xor U11653 (N_11653,N_10294,N_10043);
nor U11654 (N_11654,N_10771,N_10522);
nand U11655 (N_11655,N_10496,N_10974);
nor U11656 (N_11656,N_10454,N_10905);
or U11657 (N_11657,N_10044,N_10463);
and U11658 (N_11658,N_10646,N_10787);
or U11659 (N_11659,N_10906,N_10684);
nand U11660 (N_11660,N_10185,N_10728);
and U11661 (N_11661,N_10874,N_10478);
and U11662 (N_11662,N_10562,N_10349);
nor U11663 (N_11663,N_10595,N_10695);
nand U11664 (N_11664,N_10788,N_10103);
nand U11665 (N_11665,N_10028,N_10045);
and U11666 (N_11666,N_10872,N_10293);
or U11667 (N_11667,N_10026,N_10916);
and U11668 (N_11668,N_10471,N_10320);
and U11669 (N_11669,N_10701,N_10721);
xnor U11670 (N_11670,N_10922,N_10793);
or U11671 (N_11671,N_10819,N_10990);
xnor U11672 (N_11672,N_10616,N_10524);
or U11673 (N_11673,N_10283,N_10008);
xnor U11674 (N_11674,N_10118,N_10621);
xnor U11675 (N_11675,N_10076,N_10081);
or U11676 (N_11676,N_10231,N_10276);
and U11677 (N_11677,N_10771,N_10971);
and U11678 (N_11678,N_10948,N_10199);
nand U11679 (N_11679,N_10837,N_10360);
nor U11680 (N_11680,N_10484,N_10582);
xnor U11681 (N_11681,N_10975,N_10870);
or U11682 (N_11682,N_10033,N_10246);
nor U11683 (N_11683,N_10234,N_10394);
and U11684 (N_11684,N_10710,N_10409);
xnor U11685 (N_11685,N_10959,N_10666);
or U11686 (N_11686,N_10898,N_10947);
xnor U11687 (N_11687,N_10014,N_10138);
nor U11688 (N_11688,N_10516,N_10024);
xnor U11689 (N_11689,N_10594,N_10621);
and U11690 (N_11690,N_10128,N_10744);
or U11691 (N_11691,N_10720,N_10323);
xnor U11692 (N_11692,N_10859,N_10354);
nor U11693 (N_11693,N_10517,N_10813);
and U11694 (N_11694,N_10361,N_10574);
and U11695 (N_11695,N_10430,N_10639);
nand U11696 (N_11696,N_10830,N_10952);
xnor U11697 (N_11697,N_10050,N_10335);
nor U11698 (N_11698,N_10190,N_10687);
or U11699 (N_11699,N_10401,N_10102);
and U11700 (N_11700,N_10351,N_10177);
nand U11701 (N_11701,N_10214,N_10167);
xor U11702 (N_11702,N_10737,N_10612);
and U11703 (N_11703,N_10449,N_10367);
or U11704 (N_11704,N_10910,N_10309);
and U11705 (N_11705,N_10250,N_10900);
nor U11706 (N_11706,N_10055,N_10136);
and U11707 (N_11707,N_10040,N_10172);
nor U11708 (N_11708,N_10291,N_10908);
and U11709 (N_11709,N_10768,N_10179);
and U11710 (N_11710,N_10730,N_10385);
nor U11711 (N_11711,N_10914,N_10369);
nor U11712 (N_11712,N_10337,N_10630);
nand U11713 (N_11713,N_10311,N_10342);
and U11714 (N_11714,N_10517,N_10248);
and U11715 (N_11715,N_10217,N_10289);
and U11716 (N_11716,N_10835,N_10421);
xor U11717 (N_11717,N_10909,N_10816);
or U11718 (N_11718,N_10571,N_10879);
nand U11719 (N_11719,N_10654,N_10404);
nor U11720 (N_11720,N_10062,N_10034);
or U11721 (N_11721,N_10382,N_10027);
or U11722 (N_11722,N_10864,N_10738);
xor U11723 (N_11723,N_10083,N_10569);
xor U11724 (N_11724,N_10788,N_10884);
or U11725 (N_11725,N_10769,N_10070);
xnor U11726 (N_11726,N_10446,N_10690);
or U11727 (N_11727,N_10969,N_10740);
or U11728 (N_11728,N_10436,N_10784);
xor U11729 (N_11729,N_10214,N_10983);
and U11730 (N_11730,N_10446,N_10601);
and U11731 (N_11731,N_10539,N_10786);
or U11732 (N_11732,N_10580,N_10045);
nor U11733 (N_11733,N_10069,N_10249);
or U11734 (N_11734,N_10207,N_10526);
or U11735 (N_11735,N_10698,N_10394);
and U11736 (N_11736,N_10960,N_10922);
nand U11737 (N_11737,N_10275,N_10796);
or U11738 (N_11738,N_10999,N_10823);
xnor U11739 (N_11739,N_10374,N_10281);
xor U11740 (N_11740,N_10568,N_10204);
or U11741 (N_11741,N_10195,N_10845);
and U11742 (N_11742,N_10175,N_10892);
or U11743 (N_11743,N_10623,N_10454);
and U11744 (N_11744,N_10866,N_10496);
nand U11745 (N_11745,N_10538,N_10929);
or U11746 (N_11746,N_10566,N_10829);
or U11747 (N_11747,N_10608,N_10325);
and U11748 (N_11748,N_10037,N_10217);
nor U11749 (N_11749,N_10192,N_10980);
nand U11750 (N_11750,N_10306,N_10311);
xnor U11751 (N_11751,N_10542,N_10665);
nand U11752 (N_11752,N_10391,N_10176);
nor U11753 (N_11753,N_10874,N_10678);
or U11754 (N_11754,N_10041,N_10329);
nand U11755 (N_11755,N_10667,N_10513);
and U11756 (N_11756,N_10091,N_10852);
nor U11757 (N_11757,N_10169,N_10081);
or U11758 (N_11758,N_10684,N_10456);
or U11759 (N_11759,N_10527,N_10983);
and U11760 (N_11760,N_10180,N_10784);
and U11761 (N_11761,N_10194,N_10144);
and U11762 (N_11762,N_10053,N_10005);
xor U11763 (N_11763,N_10000,N_10256);
xor U11764 (N_11764,N_10360,N_10421);
xnor U11765 (N_11765,N_10744,N_10444);
xor U11766 (N_11766,N_10653,N_10075);
xor U11767 (N_11767,N_10819,N_10490);
and U11768 (N_11768,N_10125,N_10919);
nand U11769 (N_11769,N_10855,N_10284);
or U11770 (N_11770,N_10581,N_10315);
nand U11771 (N_11771,N_10500,N_10608);
xor U11772 (N_11772,N_10563,N_10163);
and U11773 (N_11773,N_10712,N_10587);
or U11774 (N_11774,N_10743,N_10770);
and U11775 (N_11775,N_10211,N_10633);
xnor U11776 (N_11776,N_10195,N_10921);
nor U11777 (N_11777,N_10972,N_10945);
and U11778 (N_11778,N_10883,N_10435);
nor U11779 (N_11779,N_10168,N_10085);
or U11780 (N_11780,N_10161,N_10125);
or U11781 (N_11781,N_10633,N_10436);
nor U11782 (N_11782,N_10827,N_10061);
xor U11783 (N_11783,N_10832,N_10582);
xnor U11784 (N_11784,N_10172,N_10577);
nor U11785 (N_11785,N_10361,N_10163);
and U11786 (N_11786,N_10054,N_10537);
and U11787 (N_11787,N_10244,N_10812);
xor U11788 (N_11788,N_10887,N_10277);
xnor U11789 (N_11789,N_10959,N_10138);
nand U11790 (N_11790,N_10831,N_10823);
and U11791 (N_11791,N_10797,N_10347);
nor U11792 (N_11792,N_10308,N_10649);
xor U11793 (N_11793,N_10422,N_10941);
xnor U11794 (N_11794,N_10329,N_10451);
or U11795 (N_11795,N_10904,N_10755);
and U11796 (N_11796,N_10460,N_10928);
nand U11797 (N_11797,N_10360,N_10975);
nand U11798 (N_11798,N_10623,N_10628);
xor U11799 (N_11799,N_10661,N_10612);
nand U11800 (N_11800,N_10042,N_10730);
nand U11801 (N_11801,N_10084,N_10512);
nand U11802 (N_11802,N_10878,N_10635);
nor U11803 (N_11803,N_10706,N_10217);
nand U11804 (N_11804,N_10378,N_10789);
xor U11805 (N_11805,N_10465,N_10177);
and U11806 (N_11806,N_10146,N_10791);
nand U11807 (N_11807,N_10923,N_10525);
xnor U11808 (N_11808,N_10122,N_10195);
nand U11809 (N_11809,N_10154,N_10027);
or U11810 (N_11810,N_10971,N_10361);
and U11811 (N_11811,N_10087,N_10762);
and U11812 (N_11812,N_10597,N_10104);
xnor U11813 (N_11813,N_10467,N_10687);
nand U11814 (N_11814,N_10283,N_10543);
nand U11815 (N_11815,N_10787,N_10589);
xor U11816 (N_11816,N_10486,N_10611);
nor U11817 (N_11817,N_10470,N_10751);
and U11818 (N_11818,N_10379,N_10322);
or U11819 (N_11819,N_10773,N_10790);
xnor U11820 (N_11820,N_10126,N_10368);
or U11821 (N_11821,N_10105,N_10340);
xnor U11822 (N_11822,N_10346,N_10087);
and U11823 (N_11823,N_10707,N_10980);
nor U11824 (N_11824,N_10812,N_10657);
or U11825 (N_11825,N_10739,N_10648);
xnor U11826 (N_11826,N_10714,N_10987);
and U11827 (N_11827,N_10506,N_10065);
or U11828 (N_11828,N_10096,N_10059);
nand U11829 (N_11829,N_10426,N_10293);
nor U11830 (N_11830,N_10839,N_10460);
nor U11831 (N_11831,N_10556,N_10285);
and U11832 (N_11832,N_10507,N_10398);
xor U11833 (N_11833,N_10893,N_10124);
nand U11834 (N_11834,N_10087,N_10091);
and U11835 (N_11835,N_10623,N_10617);
xnor U11836 (N_11836,N_10512,N_10677);
or U11837 (N_11837,N_10209,N_10011);
or U11838 (N_11838,N_10971,N_10175);
or U11839 (N_11839,N_10647,N_10413);
or U11840 (N_11840,N_10745,N_10981);
nand U11841 (N_11841,N_10930,N_10824);
and U11842 (N_11842,N_10768,N_10056);
or U11843 (N_11843,N_10904,N_10920);
xor U11844 (N_11844,N_10256,N_10857);
nand U11845 (N_11845,N_10028,N_10469);
nand U11846 (N_11846,N_10736,N_10487);
nand U11847 (N_11847,N_10478,N_10415);
and U11848 (N_11848,N_10807,N_10403);
or U11849 (N_11849,N_10872,N_10534);
nand U11850 (N_11850,N_10665,N_10857);
nand U11851 (N_11851,N_10562,N_10957);
nand U11852 (N_11852,N_10875,N_10997);
or U11853 (N_11853,N_10535,N_10139);
or U11854 (N_11854,N_10810,N_10398);
nand U11855 (N_11855,N_10362,N_10672);
or U11856 (N_11856,N_10278,N_10397);
nor U11857 (N_11857,N_10111,N_10103);
xnor U11858 (N_11858,N_10623,N_10726);
and U11859 (N_11859,N_10873,N_10329);
nor U11860 (N_11860,N_10591,N_10708);
nor U11861 (N_11861,N_10095,N_10137);
xnor U11862 (N_11862,N_10975,N_10145);
xor U11863 (N_11863,N_10462,N_10155);
or U11864 (N_11864,N_10901,N_10595);
nand U11865 (N_11865,N_10159,N_10626);
or U11866 (N_11866,N_10767,N_10215);
nand U11867 (N_11867,N_10905,N_10019);
nor U11868 (N_11868,N_10476,N_10157);
xor U11869 (N_11869,N_10548,N_10077);
xnor U11870 (N_11870,N_10007,N_10819);
and U11871 (N_11871,N_10617,N_10962);
or U11872 (N_11872,N_10019,N_10748);
and U11873 (N_11873,N_10114,N_10311);
and U11874 (N_11874,N_10814,N_10207);
xnor U11875 (N_11875,N_10929,N_10994);
and U11876 (N_11876,N_10301,N_10265);
or U11877 (N_11877,N_10590,N_10566);
nor U11878 (N_11878,N_10719,N_10453);
nand U11879 (N_11879,N_10144,N_10652);
nand U11880 (N_11880,N_10095,N_10212);
or U11881 (N_11881,N_10941,N_10425);
nand U11882 (N_11882,N_10778,N_10970);
nor U11883 (N_11883,N_10535,N_10624);
xnor U11884 (N_11884,N_10291,N_10897);
nand U11885 (N_11885,N_10972,N_10744);
xnor U11886 (N_11886,N_10933,N_10359);
and U11887 (N_11887,N_10539,N_10912);
xnor U11888 (N_11888,N_10366,N_10399);
xnor U11889 (N_11889,N_10361,N_10260);
or U11890 (N_11890,N_10659,N_10937);
and U11891 (N_11891,N_10527,N_10298);
nand U11892 (N_11892,N_10263,N_10751);
xnor U11893 (N_11893,N_10452,N_10858);
or U11894 (N_11894,N_10168,N_10697);
nor U11895 (N_11895,N_10027,N_10711);
nand U11896 (N_11896,N_10376,N_10105);
xor U11897 (N_11897,N_10601,N_10154);
xor U11898 (N_11898,N_10822,N_10600);
nor U11899 (N_11899,N_10744,N_10408);
nand U11900 (N_11900,N_10111,N_10098);
nand U11901 (N_11901,N_10081,N_10818);
or U11902 (N_11902,N_10773,N_10004);
nand U11903 (N_11903,N_10525,N_10962);
xor U11904 (N_11904,N_10148,N_10013);
nor U11905 (N_11905,N_10308,N_10061);
nor U11906 (N_11906,N_10832,N_10849);
or U11907 (N_11907,N_10371,N_10964);
xor U11908 (N_11908,N_10484,N_10933);
xor U11909 (N_11909,N_10592,N_10201);
xor U11910 (N_11910,N_10995,N_10150);
and U11911 (N_11911,N_10425,N_10340);
and U11912 (N_11912,N_10611,N_10896);
and U11913 (N_11913,N_10422,N_10712);
nor U11914 (N_11914,N_10121,N_10514);
nand U11915 (N_11915,N_10749,N_10161);
nor U11916 (N_11916,N_10130,N_10499);
nand U11917 (N_11917,N_10855,N_10796);
nor U11918 (N_11918,N_10294,N_10528);
and U11919 (N_11919,N_10739,N_10088);
and U11920 (N_11920,N_10584,N_10340);
nand U11921 (N_11921,N_10965,N_10708);
xnor U11922 (N_11922,N_10939,N_10424);
or U11923 (N_11923,N_10755,N_10443);
nor U11924 (N_11924,N_10568,N_10323);
nand U11925 (N_11925,N_10425,N_10946);
nor U11926 (N_11926,N_10180,N_10328);
nand U11927 (N_11927,N_10437,N_10053);
xor U11928 (N_11928,N_10787,N_10355);
and U11929 (N_11929,N_10952,N_10509);
xnor U11930 (N_11930,N_10030,N_10254);
xnor U11931 (N_11931,N_10472,N_10692);
and U11932 (N_11932,N_10056,N_10608);
xor U11933 (N_11933,N_10228,N_10294);
and U11934 (N_11934,N_10387,N_10321);
and U11935 (N_11935,N_10661,N_10466);
xnor U11936 (N_11936,N_10835,N_10519);
xor U11937 (N_11937,N_10135,N_10517);
or U11938 (N_11938,N_10633,N_10651);
and U11939 (N_11939,N_10220,N_10980);
xnor U11940 (N_11940,N_10279,N_10317);
and U11941 (N_11941,N_10795,N_10622);
nand U11942 (N_11942,N_10463,N_10000);
nand U11943 (N_11943,N_10754,N_10230);
and U11944 (N_11944,N_10614,N_10999);
xnor U11945 (N_11945,N_10063,N_10603);
or U11946 (N_11946,N_10129,N_10988);
and U11947 (N_11947,N_10151,N_10959);
nand U11948 (N_11948,N_10368,N_10383);
nor U11949 (N_11949,N_10716,N_10606);
and U11950 (N_11950,N_10041,N_10219);
or U11951 (N_11951,N_10120,N_10313);
xnor U11952 (N_11952,N_10886,N_10576);
and U11953 (N_11953,N_10582,N_10339);
xor U11954 (N_11954,N_10770,N_10718);
and U11955 (N_11955,N_10332,N_10131);
or U11956 (N_11956,N_10241,N_10045);
xnor U11957 (N_11957,N_10822,N_10466);
nand U11958 (N_11958,N_10957,N_10092);
and U11959 (N_11959,N_10696,N_10904);
and U11960 (N_11960,N_10596,N_10318);
or U11961 (N_11961,N_10400,N_10125);
nand U11962 (N_11962,N_10103,N_10090);
nor U11963 (N_11963,N_10085,N_10821);
nand U11964 (N_11964,N_10612,N_10466);
xnor U11965 (N_11965,N_10908,N_10356);
or U11966 (N_11966,N_10971,N_10929);
nor U11967 (N_11967,N_10919,N_10357);
xor U11968 (N_11968,N_10983,N_10171);
and U11969 (N_11969,N_10374,N_10250);
nand U11970 (N_11970,N_10606,N_10236);
and U11971 (N_11971,N_10600,N_10517);
nor U11972 (N_11972,N_10411,N_10741);
or U11973 (N_11973,N_10278,N_10230);
nand U11974 (N_11974,N_10692,N_10096);
or U11975 (N_11975,N_10987,N_10164);
and U11976 (N_11976,N_10619,N_10570);
nand U11977 (N_11977,N_10529,N_10400);
nand U11978 (N_11978,N_10839,N_10384);
or U11979 (N_11979,N_10108,N_10334);
and U11980 (N_11980,N_10091,N_10276);
nand U11981 (N_11981,N_10990,N_10696);
xor U11982 (N_11982,N_10841,N_10395);
or U11983 (N_11983,N_10349,N_10352);
or U11984 (N_11984,N_10911,N_10406);
or U11985 (N_11985,N_10967,N_10944);
nor U11986 (N_11986,N_10472,N_10928);
nand U11987 (N_11987,N_10032,N_10263);
xnor U11988 (N_11988,N_10989,N_10503);
xnor U11989 (N_11989,N_10012,N_10562);
xor U11990 (N_11990,N_10336,N_10681);
or U11991 (N_11991,N_10680,N_10141);
or U11992 (N_11992,N_10498,N_10652);
and U11993 (N_11993,N_10320,N_10888);
and U11994 (N_11994,N_10753,N_10200);
nor U11995 (N_11995,N_10538,N_10229);
or U11996 (N_11996,N_10636,N_10279);
nor U11997 (N_11997,N_10000,N_10855);
xnor U11998 (N_11998,N_10438,N_10103);
nand U11999 (N_11999,N_10439,N_10992);
and U12000 (N_12000,N_11452,N_11781);
and U12001 (N_12001,N_11690,N_11117);
nand U12002 (N_12002,N_11614,N_11983);
nor U12003 (N_12003,N_11047,N_11887);
nor U12004 (N_12004,N_11605,N_11577);
xor U12005 (N_12005,N_11782,N_11809);
or U12006 (N_12006,N_11975,N_11790);
xor U12007 (N_12007,N_11071,N_11817);
xor U12008 (N_12008,N_11113,N_11133);
nand U12009 (N_12009,N_11920,N_11188);
xnor U12010 (N_12010,N_11742,N_11974);
nor U12011 (N_12011,N_11526,N_11357);
nor U12012 (N_12012,N_11321,N_11602);
or U12013 (N_12013,N_11565,N_11396);
nor U12014 (N_12014,N_11640,N_11165);
nand U12015 (N_12015,N_11240,N_11827);
nor U12016 (N_12016,N_11997,N_11302);
and U12017 (N_12017,N_11941,N_11462);
nor U12018 (N_12018,N_11898,N_11391);
and U12019 (N_12019,N_11804,N_11493);
nor U12020 (N_12020,N_11433,N_11627);
nand U12021 (N_12021,N_11509,N_11850);
nand U12022 (N_12022,N_11623,N_11807);
or U12023 (N_12023,N_11888,N_11193);
and U12024 (N_12024,N_11119,N_11931);
and U12025 (N_12025,N_11649,N_11678);
nand U12026 (N_12026,N_11100,N_11570);
and U12027 (N_12027,N_11057,N_11751);
xnor U12028 (N_12028,N_11022,N_11533);
xor U12029 (N_12029,N_11486,N_11154);
nand U12030 (N_12030,N_11599,N_11358);
xor U12031 (N_12031,N_11097,N_11989);
or U12032 (N_12032,N_11428,N_11234);
xnor U12033 (N_12033,N_11684,N_11716);
or U12034 (N_12034,N_11663,N_11143);
and U12035 (N_12035,N_11819,N_11949);
and U12036 (N_12036,N_11339,N_11040);
and U12037 (N_12037,N_11399,N_11021);
nand U12038 (N_12038,N_11194,N_11140);
nand U12039 (N_12039,N_11511,N_11685);
nor U12040 (N_12040,N_11648,N_11156);
and U12041 (N_12041,N_11192,N_11408);
xor U12042 (N_12042,N_11908,N_11767);
and U12043 (N_12043,N_11544,N_11904);
nand U12044 (N_12044,N_11185,N_11628);
nand U12045 (N_12045,N_11786,N_11764);
nor U12046 (N_12046,N_11271,N_11971);
and U12047 (N_12047,N_11775,N_11993);
nor U12048 (N_12048,N_11128,N_11814);
nor U12049 (N_12049,N_11499,N_11876);
xor U12050 (N_12050,N_11946,N_11741);
xor U12051 (N_12051,N_11555,N_11168);
nor U12052 (N_12052,N_11110,N_11851);
nor U12053 (N_12053,N_11992,N_11913);
nor U12054 (N_12054,N_11410,N_11447);
or U12055 (N_12055,N_11300,N_11183);
nand U12056 (N_12056,N_11771,N_11725);
xnor U12057 (N_12057,N_11650,N_11472);
or U12058 (N_12058,N_11539,N_11413);
or U12059 (N_12059,N_11629,N_11116);
and U12060 (N_12060,N_11086,N_11606);
nand U12061 (N_12061,N_11982,N_11066);
and U12062 (N_12062,N_11593,N_11865);
nand U12063 (N_12063,N_11743,N_11615);
nand U12064 (N_12064,N_11497,N_11564);
xor U12065 (N_12065,N_11646,N_11456);
nor U12066 (N_12066,N_11706,N_11845);
nor U12067 (N_12067,N_11507,N_11502);
nand U12068 (N_12068,N_11444,N_11265);
or U12069 (N_12069,N_11607,N_11379);
and U12070 (N_12070,N_11074,N_11651);
nand U12071 (N_12071,N_11981,N_11422);
nor U12072 (N_12072,N_11642,N_11315);
and U12073 (N_12073,N_11225,N_11704);
and U12074 (N_12074,N_11178,N_11858);
xor U12075 (N_12075,N_11122,N_11988);
nor U12076 (N_12076,N_11813,N_11214);
nor U12077 (N_12077,N_11779,N_11293);
and U12078 (N_12078,N_11977,N_11731);
xor U12079 (N_12079,N_11255,N_11177);
and U12080 (N_12080,N_11039,N_11763);
nand U12081 (N_12081,N_11619,N_11187);
or U12082 (N_12082,N_11206,N_11392);
or U12083 (N_12083,N_11377,N_11231);
xor U12084 (N_12084,N_11869,N_11144);
or U12085 (N_12085,N_11191,N_11266);
and U12086 (N_12086,N_11528,N_11137);
nor U12087 (N_12087,N_11621,N_11959);
and U12088 (N_12088,N_11211,N_11317);
and U12089 (N_12089,N_11175,N_11670);
nand U12090 (N_12090,N_11045,N_11414);
nand U12091 (N_12091,N_11776,N_11603);
nand U12092 (N_12092,N_11912,N_11833);
nand U12093 (N_12093,N_11760,N_11003);
nor U12094 (N_12094,N_11868,N_11340);
or U12095 (N_12095,N_11109,N_11279);
and U12096 (N_12096,N_11824,N_11223);
xnor U12097 (N_12097,N_11314,N_11159);
or U12098 (N_12098,N_11987,N_11553);
nor U12099 (N_12099,N_11361,N_11346);
and U12100 (N_12100,N_11735,N_11364);
or U12101 (N_12101,N_11440,N_11072);
xor U12102 (N_12102,N_11837,N_11515);
nand U12103 (N_12103,N_11718,N_11802);
and U12104 (N_12104,N_11381,N_11506);
or U12105 (N_12105,N_11765,N_11008);
or U12106 (N_12106,N_11123,N_11350);
nand U12107 (N_12107,N_11939,N_11504);
xnor U12108 (N_12108,N_11873,N_11367);
and U12109 (N_12109,N_11220,N_11169);
nand U12110 (N_12110,N_11487,N_11471);
nand U12111 (N_12111,N_11483,N_11758);
xnor U12112 (N_12112,N_11469,N_11429);
nor U12113 (N_12113,N_11463,N_11980);
or U12114 (N_12114,N_11705,N_11141);
nand U12115 (N_12115,N_11519,N_11843);
xor U12116 (N_12116,N_11149,N_11454);
nor U12117 (N_12117,N_11816,N_11249);
or U12118 (N_12118,N_11874,N_11148);
or U12119 (N_12119,N_11347,N_11612);
and U12120 (N_12120,N_11571,N_11382);
or U12121 (N_12121,N_11235,N_11905);
nand U12122 (N_12122,N_11721,N_11679);
or U12123 (N_12123,N_11563,N_11942);
nor U12124 (N_12124,N_11581,N_11228);
or U12125 (N_12125,N_11277,N_11229);
xnor U12126 (N_12126,N_11625,N_11859);
nor U12127 (N_12127,N_11585,N_11488);
nor U12128 (N_12128,N_11891,N_11065);
nor U12129 (N_12129,N_11466,N_11274);
and U12130 (N_12130,N_11004,N_11963);
nor U12131 (N_12131,N_11543,N_11023);
xor U12132 (N_12132,N_11815,N_11958);
xor U12133 (N_12133,N_11923,N_11761);
nand U12134 (N_12134,N_11425,N_11991);
and U12135 (N_12135,N_11268,N_11070);
nor U12136 (N_12136,N_11616,N_11139);
nor U12137 (N_12137,N_11655,N_11884);
nor U12138 (N_12138,N_11600,N_11681);
or U12139 (N_12139,N_11821,N_11842);
nor U12140 (N_12140,N_11880,N_11592);
and U12141 (N_12141,N_11395,N_11967);
nor U12142 (N_12142,N_11244,N_11723);
or U12143 (N_12143,N_11459,N_11443);
or U12144 (N_12144,N_11245,N_11883);
nor U12145 (N_12145,N_11703,N_11479);
nor U12146 (N_12146,N_11831,N_11928);
and U12147 (N_12147,N_11841,N_11531);
or U12148 (N_12148,N_11107,N_11405);
or U12149 (N_12149,N_11675,N_11287);
or U12150 (N_12150,N_11029,N_11846);
xnor U12151 (N_12151,N_11730,N_11124);
nor U12152 (N_12152,N_11298,N_11664);
nand U12153 (N_12153,N_11952,N_11199);
or U12154 (N_12154,N_11714,N_11702);
and U12155 (N_12155,N_11369,N_11441);
and U12156 (N_12156,N_11101,N_11984);
or U12157 (N_12157,N_11748,N_11432);
and U12158 (N_12158,N_11182,N_11125);
nor U12159 (N_12159,N_11792,N_11516);
and U12160 (N_12160,N_11032,N_11344);
nor U12161 (N_12161,N_11305,N_11503);
xor U12162 (N_12162,N_11789,N_11374);
and U12163 (N_12163,N_11849,N_11878);
nand U12164 (N_12164,N_11046,N_11517);
and U12165 (N_12165,N_11586,N_11836);
and U12166 (N_12166,N_11083,N_11701);
nand U12167 (N_12167,N_11351,N_11800);
nor U12168 (N_12168,N_11398,N_11407);
and U12169 (N_12169,N_11067,N_11342);
xor U12170 (N_12170,N_11104,N_11631);
and U12171 (N_12171,N_11477,N_11412);
nor U12172 (N_12172,N_11728,N_11246);
xor U12173 (N_12173,N_11464,N_11383);
xnor U12174 (N_12174,N_11366,N_11334);
or U12175 (N_12175,N_11514,N_11881);
nand U12176 (N_12176,N_11024,N_11525);
nor U12177 (N_12177,N_11090,N_11500);
and U12178 (N_12178,N_11142,N_11009);
nor U12179 (N_12179,N_11947,N_11696);
xor U12180 (N_12180,N_11068,N_11930);
xor U12181 (N_12181,N_11442,N_11686);
nor U12182 (N_12182,N_11152,N_11257);
or U12183 (N_12183,N_11394,N_11677);
or U12184 (N_12184,N_11190,N_11167);
or U12185 (N_12185,N_11372,N_11950);
or U12186 (N_12186,N_11825,N_11840);
nand U12187 (N_12187,N_11584,N_11164);
and U12188 (N_12188,N_11508,N_11759);
and U12189 (N_12189,N_11058,N_11734);
nand U12190 (N_12190,N_11676,N_11510);
nor U12191 (N_12191,N_11915,N_11532);
nor U12192 (N_12192,N_11138,N_11711);
xor U12193 (N_12193,N_11601,N_11115);
xnor U12194 (N_12194,N_11470,N_11798);
xnor U12195 (N_12195,N_11420,N_11870);
nand U12196 (N_12196,N_11547,N_11198);
xnor U12197 (N_12197,N_11455,N_11864);
nand U12198 (N_12198,N_11360,N_11091);
nor U12199 (N_12199,N_11427,N_11201);
and U12200 (N_12200,N_11672,N_11378);
nor U12201 (N_12201,N_11285,N_11404);
nand U12202 (N_12202,N_11031,N_11536);
nor U12203 (N_12203,N_11294,N_11697);
nand U12204 (N_12204,N_11476,N_11691);
nor U12205 (N_12205,N_11892,N_11926);
nand U12206 (N_12206,N_11961,N_11400);
xor U12207 (N_12207,N_11227,N_11740);
and U12208 (N_12208,N_11431,N_11203);
nor U12209 (N_12209,N_11830,N_11535);
nand U12210 (N_12210,N_11693,N_11558);
and U12211 (N_12211,N_11386,N_11699);
and U12212 (N_12212,N_11248,N_11527);
nand U12213 (N_12213,N_11215,N_11575);
nor U12214 (N_12214,N_11017,N_11368);
or U12215 (N_12215,N_11911,N_11973);
nand U12216 (N_12216,N_11254,N_11799);
nand U12217 (N_12217,N_11902,N_11747);
or U12218 (N_12218,N_11262,N_11376);
and U12219 (N_12219,N_11630,N_11944);
or U12220 (N_12220,N_11922,N_11822);
xor U12221 (N_12221,N_11200,N_11919);
xnor U12222 (N_12222,N_11595,N_11885);
or U12223 (N_12223,N_11180,N_11823);
or U12224 (N_12224,N_11371,N_11756);
and U12225 (N_12225,N_11794,N_11251);
nor U12226 (N_12226,N_11695,N_11166);
or U12227 (N_12227,N_11299,N_11098);
xor U12228 (N_12228,N_11120,N_11269);
and U12229 (N_12229,N_11273,N_11998);
or U12230 (N_12230,N_11863,N_11540);
nor U12231 (N_12231,N_11838,N_11491);
and U12232 (N_12232,N_11524,N_11475);
and U12233 (N_12233,N_11917,N_11238);
or U12234 (N_12234,N_11309,N_11738);
and U12235 (N_12235,N_11076,N_11953);
and U12236 (N_12236,N_11498,N_11176);
and U12237 (N_12237,N_11292,N_11118);
xor U12238 (N_12238,N_11501,N_11899);
or U12239 (N_12239,N_11801,N_11457);
or U12240 (N_12240,N_11416,N_11624);
xor U12241 (N_12241,N_11943,N_11549);
nand U12242 (N_12242,N_11620,N_11935);
and U12243 (N_12243,N_11312,N_11256);
nor U12244 (N_12244,N_11202,N_11247);
nand U12245 (N_12245,N_11014,N_11095);
nand U12246 (N_12246,N_11644,N_11184);
or U12247 (N_12247,N_11985,N_11929);
xnor U12248 (N_12248,N_11925,N_11860);
and U12249 (N_12249,N_11411,N_11446);
and U12250 (N_12250,N_11772,N_11803);
xor U12251 (N_12251,N_11242,N_11662);
nand U12252 (N_12252,N_11847,N_11770);
nand U12253 (N_12253,N_11688,N_11363);
nand U12254 (N_12254,N_11250,N_11979);
nor U12255 (N_12255,N_11523,N_11330);
xnor U12256 (N_12256,N_11810,N_11522);
nand U12257 (N_12257,N_11529,N_11936);
xnor U12258 (N_12258,N_11538,N_11795);
nor U12259 (N_12259,N_11753,N_11766);
or U12260 (N_12260,N_11594,N_11064);
nor U12261 (N_12261,N_11755,N_11667);
and U12262 (N_12262,N_11557,N_11724);
or U12263 (N_12263,N_11496,N_11430);
and U12264 (N_12264,N_11559,N_11435);
nor U12265 (N_12265,N_11957,N_11835);
or U12266 (N_12266,N_11715,N_11481);
nand U12267 (N_12267,N_11236,N_11316);
nor U12268 (N_12268,N_11088,N_11060);
nor U12269 (N_12269,N_11806,N_11436);
xor U12270 (N_12270,N_11518,N_11019);
or U12271 (N_12271,N_11729,N_11886);
nor U12272 (N_12272,N_11005,N_11787);
xor U12273 (N_12273,N_11951,N_11566);
and U12274 (N_12274,N_11112,N_11204);
and U12275 (N_12275,N_11537,N_11857);
or U12276 (N_12276,N_11970,N_11181);
nor U12277 (N_12277,N_11355,N_11002);
xor U12278 (N_12278,N_11263,N_11818);
nor U12279 (N_12279,N_11468,N_11896);
xor U12280 (N_12280,N_11530,N_11207);
or U12281 (N_12281,N_11828,N_11015);
xnor U12282 (N_12282,N_11362,N_11622);
nand U12283 (N_12283,N_11707,N_11893);
and U12284 (N_12284,N_11375,N_11232);
nor U12285 (N_12285,N_11839,N_11856);
or U12286 (N_12286,N_11965,N_11296);
and U12287 (N_12287,N_11635,N_11327);
nor U12288 (N_12288,N_11658,N_11749);
xor U12289 (N_12289,N_11996,N_11134);
and U12290 (N_12290,N_11322,N_11438);
and U12291 (N_12291,N_11073,N_11576);
and U12292 (N_12292,N_11713,N_11778);
nor U12293 (N_12293,N_11796,N_11011);
nor U12294 (N_12294,N_11871,N_11954);
xnor U12295 (N_12295,N_11877,N_11030);
nor U12296 (N_12296,N_11439,N_11276);
nand U12297 (N_12297,N_11638,N_11639);
nand U12298 (N_12298,N_11937,N_11224);
or U12299 (N_12299,N_11545,N_11709);
xor U12300 (N_12300,N_11660,N_11791);
nand U12301 (N_12301,N_11708,N_11574);
nor U12302 (N_12302,N_11310,N_11567);
nor U12303 (N_12303,N_11582,N_11727);
or U12304 (N_12304,N_11932,N_11028);
and U12305 (N_12305,N_11473,N_11938);
nor U12306 (N_12306,N_11990,N_11258);
xor U12307 (N_12307,N_11048,N_11356);
and U12308 (N_12308,N_11171,N_11053);
or U12309 (N_12309,N_11520,N_11862);
xor U12310 (N_12310,N_11805,N_11853);
and U12311 (N_12311,N_11757,N_11490);
nand U12312 (N_12312,N_11001,N_11580);
xor U12313 (N_12313,N_11633,N_11389);
and U12314 (N_12314,N_11637,N_11270);
nand U12315 (N_12315,N_11035,N_11419);
nand U12316 (N_12316,N_11041,N_11513);
nor U12317 (N_12317,N_11209,N_11554);
or U12318 (N_12318,N_11163,N_11222);
or U12319 (N_12319,N_11777,N_11415);
xnor U12320 (N_12320,N_11085,N_11082);
and U12321 (N_12321,N_11084,N_11050);
or U12322 (N_12322,N_11812,N_11548);
nand U12323 (N_12323,N_11788,N_11426);
nand U12324 (N_12324,N_11754,N_11855);
and U12325 (N_12325,N_11034,N_11210);
nor U12326 (N_12326,N_11556,N_11059);
nand U12327 (N_12327,N_11306,N_11618);
xor U12328 (N_12328,N_11647,N_11056);
and U12329 (N_12329,N_11720,N_11505);
nor U12330 (N_12330,N_11080,N_11955);
or U12331 (N_12331,N_11026,N_11866);
xnor U12332 (N_12332,N_11611,N_11485);
and U12333 (N_12333,N_11089,N_11722);
and U12334 (N_12334,N_11569,N_11495);
xnor U12335 (N_12335,N_11978,N_11657);
or U12336 (N_12336,N_11634,N_11608);
xor U12337 (N_12337,N_11325,N_11283);
nand U12338 (N_12338,N_11698,N_11694);
nand U12339 (N_12339,N_11132,N_11205);
nor U12340 (N_12340,N_11352,N_11458);
nand U12341 (N_12341,N_11492,N_11746);
nand U12342 (N_12342,N_11424,N_11617);
xnor U12343 (N_12343,N_11195,N_11094);
xnor U12344 (N_12344,N_11656,N_11474);
nor U12345 (N_12345,N_11077,N_11264);
nor U12346 (N_12346,N_11719,N_11861);
or U12347 (N_12347,N_11671,N_11384);
nand U12348 (N_12348,N_11578,N_11659);
xnor U12349 (N_12349,N_11037,N_11189);
nor U12350 (N_12350,N_11587,N_11288);
and U12351 (N_12351,N_11551,N_11906);
or U12352 (N_12352,N_11093,N_11380);
or U12353 (N_12353,N_11826,N_11653);
nor U12354 (N_12354,N_11291,N_11669);
and U12355 (N_12355,N_11882,N_11387);
and U12356 (N_12356,N_11301,N_11710);
and U12357 (N_12357,N_11489,N_11272);
or U12358 (N_12358,N_11216,N_11682);
nor U12359 (N_12359,N_11598,N_11010);
and U12360 (N_12360,N_11042,N_11289);
and U12361 (N_12361,N_11999,N_11969);
and U12362 (N_12362,N_11158,N_11393);
and U12363 (N_12363,N_11145,N_11461);
nand U12364 (N_12364,N_11096,N_11945);
xor U12365 (N_12365,N_11610,N_11226);
and U12366 (N_12366,N_11894,N_11793);
xor U12367 (N_12367,N_11995,N_11829);
nor U12368 (N_12368,N_11259,N_11160);
or U12369 (N_12369,N_11962,N_11307);
nor U12370 (N_12370,N_11051,N_11927);
xnor U12371 (N_12371,N_11910,N_11036);
and U12372 (N_12372,N_11972,N_11092);
nand U12373 (N_12373,N_11897,N_11319);
or U12374 (N_12374,N_11924,N_11717);
xnor U12375 (N_12375,N_11572,N_11583);
or U12376 (N_12376,N_11121,N_11282);
nand U12377 (N_12377,N_11221,N_11534);
nor U12378 (N_12378,N_11127,N_11852);
nand U12379 (N_12379,N_11308,N_11636);
nor U12380 (N_12380,N_11780,N_11337);
nor U12381 (N_12381,N_11797,N_11909);
or U12382 (N_12382,N_11783,N_11903);
and U12383 (N_12383,N_11895,N_11752);
nor U12384 (N_12384,N_11589,N_11196);
xnor U12385 (N_12385,N_11049,N_11129);
xor U12386 (N_12386,N_11403,N_11318);
xor U12387 (N_12387,N_11541,N_11018);
nor U12388 (N_12388,N_11230,N_11683);
xnor U12389 (N_12389,N_11774,N_11512);
and U12390 (N_12390,N_11964,N_11114);
xor U12391 (N_12391,N_11645,N_11712);
or U12392 (N_12392,N_11521,N_11460);
nand U12393 (N_12393,N_11237,N_11733);
or U12394 (N_12394,N_11590,N_11437);
nor U12395 (N_12395,N_11641,N_11007);
or U12396 (N_12396,N_11153,N_11006);
nor U12397 (N_12397,N_11079,N_11162);
xnor U12398 (N_12398,N_11561,N_11324);
and U12399 (N_12399,N_11668,N_11373);
and U12400 (N_12400,N_11820,N_11260);
nand U12401 (N_12401,N_11478,N_11700);
nand U12402 (N_12402,N_11013,N_11170);
nand U12403 (N_12403,N_11654,N_11808);
and U12404 (N_12404,N_11147,N_11406);
or U12405 (N_12405,N_11768,N_11033);
and U12406 (N_12406,N_11890,N_11421);
nand U12407 (N_12407,N_11020,N_11130);
nand U12408 (N_12408,N_11243,N_11157);
nor U12409 (N_12409,N_11054,N_11773);
nor U12410 (N_12410,N_11632,N_11451);
nor U12411 (N_12411,N_11689,N_11025);
nand U12412 (N_12412,N_11241,N_11297);
or U12413 (N_12413,N_11326,N_11673);
or U12414 (N_12414,N_11854,N_11434);
or U12415 (N_12415,N_11666,N_11354);
and U12416 (N_12416,N_11313,N_11609);
and U12417 (N_12417,N_11409,N_11901);
nand U12418 (N_12418,N_11345,N_11562);
or U12419 (N_12419,N_11875,N_11343);
nand U12420 (N_12420,N_11365,N_11044);
nand U12421 (N_12421,N_11359,N_11311);
nand U12422 (N_12422,N_11484,N_11063);
nor U12423 (N_12423,N_11994,N_11450);
xor U12424 (N_12424,N_11161,N_11323);
nor U12425 (N_12425,N_11736,N_11052);
nand U12426 (N_12426,N_11626,N_11131);
nand U12427 (N_12427,N_11568,N_11331);
xor U12428 (N_12428,N_11043,N_11550);
xnor U12429 (N_12429,N_11151,N_11219);
xnor U12430 (N_12430,N_11136,N_11069);
nand U12431 (N_12431,N_11332,N_11016);
or U12432 (N_12432,N_11055,N_11081);
xnor U12433 (N_12433,N_11546,N_11267);
or U12434 (N_12434,N_11286,N_11328);
nand U12435 (N_12435,N_11834,N_11062);
nand U12436 (N_12436,N_11832,N_11333);
nand U12437 (N_12437,N_11150,N_11811);
nor U12438 (N_12438,N_11349,N_11872);
xor U12439 (N_12439,N_11239,N_11579);
nand U12440 (N_12440,N_11986,N_11916);
nand U12441 (N_12441,N_11652,N_11105);
or U12442 (N_12442,N_11106,N_11338);
or U12443 (N_12443,N_11948,N_11370);
xor U12444 (N_12444,N_11336,N_11465);
or U12445 (N_12445,N_11111,N_11745);
or U12446 (N_12446,N_11934,N_11665);
nor U12447 (N_12447,N_11208,N_11341);
and U12448 (N_12448,N_11000,N_11687);
or U12449 (N_12449,N_11867,N_11402);
nor U12450 (N_12450,N_11275,N_11921);
or U12451 (N_12451,N_11290,N_11785);
nor U12452 (N_12452,N_11844,N_11417);
nand U12453 (N_12453,N_11284,N_11335);
xor U12454 (N_12454,N_11960,N_11281);
nor U12455 (N_12455,N_11956,N_11726);
nor U12456 (N_12456,N_11692,N_11918);
and U12457 (N_12457,N_11212,N_11613);
nor U12458 (N_12458,N_11732,N_11217);
or U12459 (N_12459,N_11233,N_11108);
nand U12460 (N_12460,N_11329,N_11588);
nor U12461 (N_12461,N_11966,N_11103);
and U12462 (N_12462,N_11744,N_11900);
and U12463 (N_12463,N_11889,N_11769);
or U12464 (N_12464,N_11038,N_11186);
and U12465 (N_12465,N_11353,N_11552);
or U12466 (N_12466,N_11449,N_11012);
nor U12467 (N_12467,N_11596,N_11643);
nor U12468 (N_12468,N_11218,N_11303);
xor U12469 (N_12469,N_11494,N_11401);
or U12470 (N_12470,N_11453,N_11591);
or U12471 (N_12471,N_11252,N_11280);
xor U12472 (N_12472,N_11914,N_11907);
or U12473 (N_12473,N_11135,N_11423);
xnor U12474 (N_12474,N_11968,N_11197);
xnor U12475 (N_12475,N_11674,N_11390);
and U12476 (N_12476,N_11750,N_11179);
or U12477 (N_12477,N_11261,N_11542);
and U12478 (N_12478,N_11680,N_11604);
nor U12479 (N_12479,N_11739,N_11448);
and U12480 (N_12480,N_11467,N_11174);
and U12481 (N_12481,N_11087,N_11976);
and U12482 (N_12482,N_11172,N_11295);
nand U12483 (N_12483,N_11661,N_11445);
xor U12484 (N_12484,N_11027,N_11173);
and U12485 (N_12485,N_11480,N_11560);
and U12486 (N_12486,N_11304,N_11278);
nand U12487 (N_12487,N_11213,N_11078);
or U12488 (N_12488,N_11418,N_11573);
xor U12489 (N_12489,N_11762,N_11075);
or U12490 (N_12490,N_11061,N_11397);
or U12491 (N_12491,N_11253,N_11388);
or U12492 (N_12492,N_11848,N_11933);
xnor U12493 (N_12493,N_11099,N_11879);
nand U12494 (N_12494,N_11102,N_11126);
and U12495 (N_12495,N_11146,N_11784);
or U12496 (N_12496,N_11348,N_11155);
nor U12497 (N_12497,N_11940,N_11597);
and U12498 (N_12498,N_11320,N_11385);
and U12499 (N_12499,N_11482,N_11737);
and U12500 (N_12500,N_11224,N_11661);
nand U12501 (N_12501,N_11338,N_11460);
nand U12502 (N_12502,N_11197,N_11167);
nor U12503 (N_12503,N_11751,N_11046);
or U12504 (N_12504,N_11261,N_11133);
nor U12505 (N_12505,N_11373,N_11289);
xor U12506 (N_12506,N_11288,N_11773);
or U12507 (N_12507,N_11930,N_11105);
and U12508 (N_12508,N_11667,N_11739);
or U12509 (N_12509,N_11074,N_11256);
xnor U12510 (N_12510,N_11166,N_11457);
and U12511 (N_12511,N_11237,N_11032);
or U12512 (N_12512,N_11967,N_11754);
or U12513 (N_12513,N_11574,N_11188);
nand U12514 (N_12514,N_11691,N_11179);
and U12515 (N_12515,N_11724,N_11013);
nand U12516 (N_12516,N_11251,N_11192);
nand U12517 (N_12517,N_11972,N_11884);
and U12518 (N_12518,N_11393,N_11914);
xnor U12519 (N_12519,N_11529,N_11293);
or U12520 (N_12520,N_11487,N_11966);
xnor U12521 (N_12521,N_11858,N_11426);
nor U12522 (N_12522,N_11642,N_11344);
and U12523 (N_12523,N_11369,N_11487);
xnor U12524 (N_12524,N_11100,N_11195);
xnor U12525 (N_12525,N_11323,N_11090);
and U12526 (N_12526,N_11033,N_11478);
nor U12527 (N_12527,N_11156,N_11953);
or U12528 (N_12528,N_11312,N_11696);
and U12529 (N_12529,N_11263,N_11840);
and U12530 (N_12530,N_11899,N_11287);
or U12531 (N_12531,N_11103,N_11173);
nor U12532 (N_12532,N_11163,N_11125);
and U12533 (N_12533,N_11447,N_11310);
or U12534 (N_12534,N_11930,N_11891);
nand U12535 (N_12535,N_11215,N_11529);
or U12536 (N_12536,N_11715,N_11911);
and U12537 (N_12537,N_11998,N_11382);
nand U12538 (N_12538,N_11529,N_11018);
nor U12539 (N_12539,N_11189,N_11279);
xor U12540 (N_12540,N_11578,N_11588);
and U12541 (N_12541,N_11627,N_11369);
or U12542 (N_12542,N_11895,N_11616);
nand U12543 (N_12543,N_11791,N_11064);
xnor U12544 (N_12544,N_11952,N_11972);
or U12545 (N_12545,N_11893,N_11786);
nor U12546 (N_12546,N_11134,N_11014);
nor U12547 (N_12547,N_11942,N_11620);
nand U12548 (N_12548,N_11776,N_11705);
and U12549 (N_12549,N_11233,N_11554);
nand U12550 (N_12550,N_11652,N_11409);
and U12551 (N_12551,N_11199,N_11413);
and U12552 (N_12552,N_11400,N_11084);
xor U12553 (N_12553,N_11408,N_11425);
xnor U12554 (N_12554,N_11458,N_11445);
xor U12555 (N_12555,N_11202,N_11177);
xnor U12556 (N_12556,N_11502,N_11809);
or U12557 (N_12557,N_11471,N_11419);
nand U12558 (N_12558,N_11323,N_11634);
or U12559 (N_12559,N_11305,N_11392);
xnor U12560 (N_12560,N_11972,N_11574);
and U12561 (N_12561,N_11574,N_11144);
xor U12562 (N_12562,N_11338,N_11068);
nand U12563 (N_12563,N_11793,N_11137);
xor U12564 (N_12564,N_11710,N_11234);
xor U12565 (N_12565,N_11097,N_11680);
and U12566 (N_12566,N_11301,N_11193);
nor U12567 (N_12567,N_11424,N_11843);
nand U12568 (N_12568,N_11971,N_11010);
xnor U12569 (N_12569,N_11070,N_11473);
xnor U12570 (N_12570,N_11245,N_11406);
nand U12571 (N_12571,N_11561,N_11212);
or U12572 (N_12572,N_11320,N_11607);
nand U12573 (N_12573,N_11033,N_11302);
nor U12574 (N_12574,N_11744,N_11507);
xnor U12575 (N_12575,N_11050,N_11007);
and U12576 (N_12576,N_11666,N_11575);
and U12577 (N_12577,N_11944,N_11818);
nor U12578 (N_12578,N_11822,N_11032);
or U12579 (N_12579,N_11868,N_11824);
and U12580 (N_12580,N_11660,N_11475);
and U12581 (N_12581,N_11532,N_11450);
nand U12582 (N_12582,N_11510,N_11333);
or U12583 (N_12583,N_11091,N_11937);
nor U12584 (N_12584,N_11186,N_11223);
nand U12585 (N_12585,N_11291,N_11921);
nor U12586 (N_12586,N_11198,N_11891);
or U12587 (N_12587,N_11775,N_11096);
nand U12588 (N_12588,N_11286,N_11132);
or U12589 (N_12589,N_11134,N_11294);
or U12590 (N_12590,N_11805,N_11781);
xnor U12591 (N_12591,N_11806,N_11054);
nand U12592 (N_12592,N_11629,N_11165);
or U12593 (N_12593,N_11579,N_11947);
nor U12594 (N_12594,N_11668,N_11298);
xor U12595 (N_12595,N_11831,N_11374);
xor U12596 (N_12596,N_11218,N_11328);
xnor U12597 (N_12597,N_11670,N_11529);
nand U12598 (N_12598,N_11051,N_11855);
or U12599 (N_12599,N_11007,N_11205);
or U12600 (N_12600,N_11231,N_11553);
and U12601 (N_12601,N_11240,N_11032);
nor U12602 (N_12602,N_11479,N_11101);
nand U12603 (N_12603,N_11945,N_11761);
or U12604 (N_12604,N_11564,N_11078);
and U12605 (N_12605,N_11810,N_11458);
xnor U12606 (N_12606,N_11036,N_11951);
xor U12607 (N_12607,N_11853,N_11481);
nor U12608 (N_12608,N_11203,N_11902);
nand U12609 (N_12609,N_11028,N_11279);
and U12610 (N_12610,N_11047,N_11637);
nor U12611 (N_12611,N_11546,N_11694);
xor U12612 (N_12612,N_11445,N_11810);
xor U12613 (N_12613,N_11315,N_11028);
and U12614 (N_12614,N_11707,N_11703);
nand U12615 (N_12615,N_11906,N_11380);
or U12616 (N_12616,N_11661,N_11793);
xor U12617 (N_12617,N_11836,N_11489);
nand U12618 (N_12618,N_11129,N_11760);
or U12619 (N_12619,N_11341,N_11300);
nand U12620 (N_12620,N_11056,N_11510);
or U12621 (N_12621,N_11784,N_11695);
or U12622 (N_12622,N_11535,N_11753);
xor U12623 (N_12623,N_11270,N_11916);
nor U12624 (N_12624,N_11915,N_11749);
or U12625 (N_12625,N_11117,N_11509);
nor U12626 (N_12626,N_11377,N_11370);
xor U12627 (N_12627,N_11627,N_11705);
nor U12628 (N_12628,N_11981,N_11019);
or U12629 (N_12629,N_11125,N_11982);
or U12630 (N_12630,N_11074,N_11842);
nor U12631 (N_12631,N_11843,N_11742);
xnor U12632 (N_12632,N_11329,N_11920);
and U12633 (N_12633,N_11576,N_11986);
nand U12634 (N_12634,N_11815,N_11205);
xnor U12635 (N_12635,N_11597,N_11738);
or U12636 (N_12636,N_11487,N_11093);
or U12637 (N_12637,N_11682,N_11200);
nand U12638 (N_12638,N_11205,N_11966);
xor U12639 (N_12639,N_11186,N_11591);
nor U12640 (N_12640,N_11732,N_11355);
nand U12641 (N_12641,N_11739,N_11453);
or U12642 (N_12642,N_11411,N_11741);
nor U12643 (N_12643,N_11351,N_11031);
or U12644 (N_12644,N_11102,N_11544);
and U12645 (N_12645,N_11203,N_11848);
and U12646 (N_12646,N_11229,N_11831);
nand U12647 (N_12647,N_11289,N_11741);
xnor U12648 (N_12648,N_11388,N_11160);
nor U12649 (N_12649,N_11433,N_11259);
xnor U12650 (N_12650,N_11057,N_11831);
or U12651 (N_12651,N_11046,N_11960);
or U12652 (N_12652,N_11551,N_11528);
or U12653 (N_12653,N_11625,N_11135);
or U12654 (N_12654,N_11815,N_11725);
xor U12655 (N_12655,N_11252,N_11971);
nor U12656 (N_12656,N_11877,N_11701);
nand U12657 (N_12657,N_11631,N_11525);
xor U12658 (N_12658,N_11967,N_11694);
or U12659 (N_12659,N_11703,N_11416);
nor U12660 (N_12660,N_11937,N_11137);
or U12661 (N_12661,N_11417,N_11880);
and U12662 (N_12662,N_11590,N_11489);
nand U12663 (N_12663,N_11340,N_11414);
and U12664 (N_12664,N_11691,N_11709);
nand U12665 (N_12665,N_11435,N_11163);
or U12666 (N_12666,N_11086,N_11685);
nand U12667 (N_12667,N_11805,N_11831);
nor U12668 (N_12668,N_11734,N_11751);
and U12669 (N_12669,N_11009,N_11081);
nor U12670 (N_12670,N_11777,N_11362);
xnor U12671 (N_12671,N_11633,N_11933);
or U12672 (N_12672,N_11198,N_11893);
and U12673 (N_12673,N_11096,N_11731);
nand U12674 (N_12674,N_11651,N_11129);
nor U12675 (N_12675,N_11371,N_11730);
nor U12676 (N_12676,N_11656,N_11746);
nand U12677 (N_12677,N_11793,N_11696);
nand U12678 (N_12678,N_11048,N_11281);
or U12679 (N_12679,N_11141,N_11642);
and U12680 (N_12680,N_11674,N_11324);
and U12681 (N_12681,N_11204,N_11517);
or U12682 (N_12682,N_11439,N_11797);
nor U12683 (N_12683,N_11491,N_11183);
nand U12684 (N_12684,N_11769,N_11107);
xor U12685 (N_12685,N_11760,N_11047);
nand U12686 (N_12686,N_11712,N_11691);
nor U12687 (N_12687,N_11166,N_11117);
xor U12688 (N_12688,N_11518,N_11259);
nand U12689 (N_12689,N_11992,N_11111);
nor U12690 (N_12690,N_11444,N_11756);
xor U12691 (N_12691,N_11761,N_11291);
nand U12692 (N_12692,N_11729,N_11887);
nor U12693 (N_12693,N_11576,N_11405);
nor U12694 (N_12694,N_11424,N_11192);
or U12695 (N_12695,N_11747,N_11904);
or U12696 (N_12696,N_11341,N_11778);
nor U12697 (N_12697,N_11073,N_11662);
nor U12698 (N_12698,N_11394,N_11306);
nor U12699 (N_12699,N_11063,N_11245);
nand U12700 (N_12700,N_11501,N_11427);
nand U12701 (N_12701,N_11726,N_11994);
xnor U12702 (N_12702,N_11228,N_11753);
and U12703 (N_12703,N_11452,N_11585);
xor U12704 (N_12704,N_11467,N_11659);
xor U12705 (N_12705,N_11356,N_11287);
nand U12706 (N_12706,N_11099,N_11570);
nand U12707 (N_12707,N_11501,N_11375);
and U12708 (N_12708,N_11082,N_11349);
or U12709 (N_12709,N_11874,N_11833);
nand U12710 (N_12710,N_11632,N_11741);
xor U12711 (N_12711,N_11799,N_11882);
or U12712 (N_12712,N_11270,N_11402);
nor U12713 (N_12713,N_11561,N_11867);
nor U12714 (N_12714,N_11874,N_11945);
nand U12715 (N_12715,N_11885,N_11162);
nor U12716 (N_12716,N_11998,N_11963);
nand U12717 (N_12717,N_11725,N_11792);
nand U12718 (N_12718,N_11802,N_11175);
or U12719 (N_12719,N_11872,N_11266);
nor U12720 (N_12720,N_11520,N_11245);
or U12721 (N_12721,N_11759,N_11545);
nor U12722 (N_12722,N_11290,N_11621);
and U12723 (N_12723,N_11274,N_11675);
nor U12724 (N_12724,N_11122,N_11962);
nand U12725 (N_12725,N_11445,N_11420);
and U12726 (N_12726,N_11381,N_11370);
nor U12727 (N_12727,N_11855,N_11808);
or U12728 (N_12728,N_11596,N_11044);
or U12729 (N_12729,N_11323,N_11466);
nor U12730 (N_12730,N_11372,N_11145);
and U12731 (N_12731,N_11752,N_11008);
or U12732 (N_12732,N_11889,N_11962);
and U12733 (N_12733,N_11763,N_11268);
or U12734 (N_12734,N_11660,N_11410);
and U12735 (N_12735,N_11724,N_11016);
xnor U12736 (N_12736,N_11492,N_11964);
and U12737 (N_12737,N_11949,N_11222);
nand U12738 (N_12738,N_11576,N_11436);
or U12739 (N_12739,N_11828,N_11911);
nor U12740 (N_12740,N_11672,N_11613);
or U12741 (N_12741,N_11568,N_11697);
and U12742 (N_12742,N_11248,N_11648);
nand U12743 (N_12743,N_11309,N_11074);
xor U12744 (N_12744,N_11972,N_11900);
xnor U12745 (N_12745,N_11090,N_11739);
nor U12746 (N_12746,N_11019,N_11230);
nor U12747 (N_12747,N_11901,N_11325);
or U12748 (N_12748,N_11879,N_11147);
and U12749 (N_12749,N_11613,N_11804);
or U12750 (N_12750,N_11763,N_11294);
nor U12751 (N_12751,N_11530,N_11772);
xor U12752 (N_12752,N_11664,N_11090);
and U12753 (N_12753,N_11793,N_11070);
xnor U12754 (N_12754,N_11691,N_11149);
and U12755 (N_12755,N_11288,N_11434);
and U12756 (N_12756,N_11925,N_11584);
nand U12757 (N_12757,N_11093,N_11662);
nor U12758 (N_12758,N_11824,N_11053);
nand U12759 (N_12759,N_11463,N_11139);
or U12760 (N_12760,N_11325,N_11701);
nor U12761 (N_12761,N_11769,N_11885);
and U12762 (N_12762,N_11342,N_11518);
nor U12763 (N_12763,N_11248,N_11262);
xnor U12764 (N_12764,N_11856,N_11158);
and U12765 (N_12765,N_11313,N_11727);
nor U12766 (N_12766,N_11016,N_11127);
or U12767 (N_12767,N_11819,N_11971);
and U12768 (N_12768,N_11113,N_11287);
nand U12769 (N_12769,N_11521,N_11271);
or U12770 (N_12770,N_11307,N_11101);
nand U12771 (N_12771,N_11572,N_11386);
nand U12772 (N_12772,N_11422,N_11631);
nand U12773 (N_12773,N_11677,N_11647);
and U12774 (N_12774,N_11605,N_11696);
nand U12775 (N_12775,N_11653,N_11946);
xor U12776 (N_12776,N_11286,N_11491);
nand U12777 (N_12777,N_11769,N_11098);
xor U12778 (N_12778,N_11983,N_11455);
xor U12779 (N_12779,N_11702,N_11732);
nand U12780 (N_12780,N_11730,N_11751);
nand U12781 (N_12781,N_11803,N_11291);
nand U12782 (N_12782,N_11471,N_11327);
nor U12783 (N_12783,N_11231,N_11300);
xor U12784 (N_12784,N_11098,N_11922);
nor U12785 (N_12785,N_11389,N_11337);
xnor U12786 (N_12786,N_11453,N_11336);
or U12787 (N_12787,N_11861,N_11359);
nand U12788 (N_12788,N_11824,N_11300);
nor U12789 (N_12789,N_11495,N_11263);
xnor U12790 (N_12790,N_11725,N_11879);
nand U12791 (N_12791,N_11087,N_11560);
or U12792 (N_12792,N_11229,N_11573);
and U12793 (N_12793,N_11458,N_11193);
nor U12794 (N_12794,N_11052,N_11985);
xnor U12795 (N_12795,N_11746,N_11302);
or U12796 (N_12796,N_11263,N_11597);
xnor U12797 (N_12797,N_11248,N_11132);
and U12798 (N_12798,N_11235,N_11961);
nand U12799 (N_12799,N_11739,N_11674);
xnor U12800 (N_12800,N_11775,N_11206);
and U12801 (N_12801,N_11909,N_11066);
or U12802 (N_12802,N_11238,N_11001);
or U12803 (N_12803,N_11166,N_11734);
nor U12804 (N_12804,N_11481,N_11435);
nand U12805 (N_12805,N_11629,N_11046);
nor U12806 (N_12806,N_11592,N_11071);
nor U12807 (N_12807,N_11734,N_11864);
xor U12808 (N_12808,N_11794,N_11125);
or U12809 (N_12809,N_11728,N_11308);
xor U12810 (N_12810,N_11382,N_11647);
and U12811 (N_12811,N_11520,N_11716);
nand U12812 (N_12812,N_11783,N_11256);
or U12813 (N_12813,N_11931,N_11584);
and U12814 (N_12814,N_11767,N_11268);
nor U12815 (N_12815,N_11967,N_11537);
and U12816 (N_12816,N_11047,N_11382);
or U12817 (N_12817,N_11834,N_11082);
or U12818 (N_12818,N_11055,N_11167);
nand U12819 (N_12819,N_11591,N_11397);
or U12820 (N_12820,N_11049,N_11995);
and U12821 (N_12821,N_11525,N_11610);
nand U12822 (N_12822,N_11959,N_11636);
xnor U12823 (N_12823,N_11789,N_11345);
nand U12824 (N_12824,N_11948,N_11228);
or U12825 (N_12825,N_11916,N_11307);
or U12826 (N_12826,N_11197,N_11377);
xnor U12827 (N_12827,N_11275,N_11833);
nor U12828 (N_12828,N_11953,N_11560);
and U12829 (N_12829,N_11899,N_11078);
xnor U12830 (N_12830,N_11450,N_11397);
or U12831 (N_12831,N_11579,N_11965);
xnor U12832 (N_12832,N_11643,N_11522);
nand U12833 (N_12833,N_11239,N_11524);
and U12834 (N_12834,N_11723,N_11056);
or U12835 (N_12835,N_11631,N_11092);
nor U12836 (N_12836,N_11158,N_11887);
nor U12837 (N_12837,N_11537,N_11994);
nor U12838 (N_12838,N_11334,N_11916);
xnor U12839 (N_12839,N_11900,N_11037);
nand U12840 (N_12840,N_11404,N_11760);
or U12841 (N_12841,N_11149,N_11690);
xor U12842 (N_12842,N_11388,N_11401);
or U12843 (N_12843,N_11104,N_11384);
xor U12844 (N_12844,N_11260,N_11803);
nand U12845 (N_12845,N_11119,N_11915);
and U12846 (N_12846,N_11916,N_11811);
nand U12847 (N_12847,N_11752,N_11361);
nand U12848 (N_12848,N_11011,N_11008);
xor U12849 (N_12849,N_11634,N_11774);
xnor U12850 (N_12850,N_11188,N_11947);
and U12851 (N_12851,N_11576,N_11802);
xnor U12852 (N_12852,N_11802,N_11309);
or U12853 (N_12853,N_11135,N_11111);
nor U12854 (N_12854,N_11394,N_11009);
nand U12855 (N_12855,N_11917,N_11466);
or U12856 (N_12856,N_11225,N_11618);
xor U12857 (N_12857,N_11236,N_11866);
nor U12858 (N_12858,N_11278,N_11461);
or U12859 (N_12859,N_11938,N_11579);
and U12860 (N_12860,N_11451,N_11490);
xnor U12861 (N_12861,N_11680,N_11509);
or U12862 (N_12862,N_11109,N_11619);
xnor U12863 (N_12863,N_11688,N_11012);
or U12864 (N_12864,N_11209,N_11116);
and U12865 (N_12865,N_11661,N_11607);
xor U12866 (N_12866,N_11276,N_11357);
xnor U12867 (N_12867,N_11298,N_11158);
or U12868 (N_12868,N_11492,N_11805);
xnor U12869 (N_12869,N_11611,N_11333);
nor U12870 (N_12870,N_11941,N_11010);
nor U12871 (N_12871,N_11584,N_11535);
xor U12872 (N_12872,N_11781,N_11819);
xnor U12873 (N_12873,N_11405,N_11841);
nor U12874 (N_12874,N_11214,N_11030);
nand U12875 (N_12875,N_11037,N_11573);
xor U12876 (N_12876,N_11021,N_11674);
or U12877 (N_12877,N_11989,N_11059);
xor U12878 (N_12878,N_11918,N_11521);
or U12879 (N_12879,N_11681,N_11570);
nor U12880 (N_12880,N_11122,N_11574);
or U12881 (N_12881,N_11686,N_11433);
nand U12882 (N_12882,N_11573,N_11578);
nand U12883 (N_12883,N_11765,N_11125);
nor U12884 (N_12884,N_11744,N_11430);
nor U12885 (N_12885,N_11241,N_11482);
or U12886 (N_12886,N_11546,N_11475);
nand U12887 (N_12887,N_11695,N_11071);
xor U12888 (N_12888,N_11587,N_11922);
nor U12889 (N_12889,N_11560,N_11769);
nand U12890 (N_12890,N_11310,N_11667);
or U12891 (N_12891,N_11739,N_11841);
nand U12892 (N_12892,N_11956,N_11901);
and U12893 (N_12893,N_11679,N_11572);
nand U12894 (N_12894,N_11943,N_11772);
nand U12895 (N_12895,N_11012,N_11096);
or U12896 (N_12896,N_11410,N_11010);
nor U12897 (N_12897,N_11689,N_11671);
nand U12898 (N_12898,N_11020,N_11445);
nand U12899 (N_12899,N_11095,N_11366);
and U12900 (N_12900,N_11570,N_11843);
or U12901 (N_12901,N_11981,N_11264);
or U12902 (N_12902,N_11980,N_11747);
nand U12903 (N_12903,N_11198,N_11372);
or U12904 (N_12904,N_11581,N_11926);
or U12905 (N_12905,N_11814,N_11848);
or U12906 (N_12906,N_11382,N_11543);
nand U12907 (N_12907,N_11756,N_11041);
nand U12908 (N_12908,N_11496,N_11945);
xnor U12909 (N_12909,N_11578,N_11876);
xor U12910 (N_12910,N_11597,N_11805);
or U12911 (N_12911,N_11599,N_11504);
and U12912 (N_12912,N_11728,N_11241);
or U12913 (N_12913,N_11472,N_11800);
and U12914 (N_12914,N_11824,N_11104);
or U12915 (N_12915,N_11388,N_11231);
and U12916 (N_12916,N_11376,N_11404);
or U12917 (N_12917,N_11530,N_11990);
nand U12918 (N_12918,N_11374,N_11375);
nor U12919 (N_12919,N_11962,N_11815);
nand U12920 (N_12920,N_11189,N_11689);
or U12921 (N_12921,N_11532,N_11571);
nand U12922 (N_12922,N_11767,N_11313);
or U12923 (N_12923,N_11801,N_11945);
nor U12924 (N_12924,N_11214,N_11095);
and U12925 (N_12925,N_11785,N_11056);
or U12926 (N_12926,N_11219,N_11664);
and U12927 (N_12927,N_11911,N_11410);
nand U12928 (N_12928,N_11168,N_11317);
and U12929 (N_12929,N_11848,N_11377);
or U12930 (N_12930,N_11104,N_11369);
or U12931 (N_12931,N_11004,N_11090);
and U12932 (N_12932,N_11871,N_11600);
nand U12933 (N_12933,N_11065,N_11407);
xor U12934 (N_12934,N_11225,N_11735);
xnor U12935 (N_12935,N_11329,N_11440);
nor U12936 (N_12936,N_11527,N_11205);
nor U12937 (N_12937,N_11922,N_11193);
or U12938 (N_12938,N_11216,N_11322);
and U12939 (N_12939,N_11532,N_11889);
or U12940 (N_12940,N_11194,N_11037);
nand U12941 (N_12941,N_11105,N_11015);
nor U12942 (N_12942,N_11761,N_11566);
and U12943 (N_12943,N_11933,N_11162);
xor U12944 (N_12944,N_11400,N_11412);
nor U12945 (N_12945,N_11974,N_11882);
nand U12946 (N_12946,N_11419,N_11820);
or U12947 (N_12947,N_11124,N_11450);
xnor U12948 (N_12948,N_11951,N_11403);
or U12949 (N_12949,N_11545,N_11939);
and U12950 (N_12950,N_11919,N_11292);
nand U12951 (N_12951,N_11139,N_11000);
or U12952 (N_12952,N_11681,N_11324);
nor U12953 (N_12953,N_11113,N_11254);
and U12954 (N_12954,N_11185,N_11882);
and U12955 (N_12955,N_11911,N_11822);
nand U12956 (N_12956,N_11688,N_11767);
and U12957 (N_12957,N_11810,N_11330);
and U12958 (N_12958,N_11877,N_11674);
or U12959 (N_12959,N_11079,N_11150);
or U12960 (N_12960,N_11371,N_11631);
nand U12961 (N_12961,N_11825,N_11433);
and U12962 (N_12962,N_11412,N_11872);
or U12963 (N_12963,N_11099,N_11192);
xor U12964 (N_12964,N_11546,N_11985);
nor U12965 (N_12965,N_11597,N_11475);
nor U12966 (N_12966,N_11395,N_11089);
or U12967 (N_12967,N_11704,N_11135);
nand U12968 (N_12968,N_11832,N_11826);
and U12969 (N_12969,N_11690,N_11893);
xnor U12970 (N_12970,N_11266,N_11016);
nor U12971 (N_12971,N_11511,N_11380);
nor U12972 (N_12972,N_11387,N_11714);
nand U12973 (N_12973,N_11817,N_11755);
nor U12974 (N_12974,N_11413,N_11999);
and U12975 (N_12975,N_11843,N_11449);
or U12976 (N_12976,N_11089,N_11052);
nor U12977 (N_12977,N_11259,N_11426);
or U12978 (N_12978,N_11318,N_11142);
xor U12979 (N_12979,N_11177,N_11903);
xnor U12980 (N_12980,N_11321,N_11855);
nor U12981 (N_12981,N_11616,N_11642);
xor U12982 (N_12982,N_11246,N_11523);
or U12983 (N_12983,N_11699,N_11318);
or U12984 (N_12984,N_11253,N_11519);
or U12985 (N_12985,N_11453,N_11766);
or U12986 (N_12986,N_11212,N_11963);
xor U12987 (N_12987,N_11829,N_11726);
or U12988 (N_12988,N_11538,N_11275);
and U12989 (N_12989,N_11652,N_11005);
nand U12990 (N_12990,N_11169,N_11777);
nand U12991 (N_12991,N_11513,N_11370);
or U12992 (N_12992,N_11712,N_11253);
nor U12993 (N_12993,N_11953,N_11569);
and U12994 (N_12994,N_11495,N_11243);
nor U12995 (N_12995,N_11132,N_11880);
nor U12996 (N_12996,N_11286,N_11767);
xnor U12997 (N_12997,N_11551,N_11031);
nand U12998 (N_12998,N_11389,N_11883);
and U12999 (N_12999,N_11353,N_11564);
nand U13000 (N_13000,N_12921,N_12629);
xor U13001 (N_13001,N_12498,N_12485);
nor U13002 (N_13002,N_12997,N_12819);
or U13003 (N_13003,N_12540,N_12324);
or U13004 (N_13004,N_12019,N_12685);
nand U13005 (N_13005,N_12695,N_12200);
or U13006 (N_13006,N_12349,N_12398);
and U13007 (N_13007,N_12592,N_12919);
nand U13008 (N_13008,N_12242,N_12886);
and U13009 (N_13009,N_12007,N_12317);
nor U13010 (N_13010,N_12751,N_12191);
or U13011 (N_13011,N_12437,N_12616);
xor U13012 (N_13012,N_12532,N_12712);
and U13013 (N_13013,N_12418,N_12541);
xnor U13014 (N_13014,N_12406,N_12464);
nor U13015 (N_13015,N_12284,N_12419);
nand U13016 (N_13016,N_12421,N_12246);
nand U13017 (N_13017,N_12615,N_12223);
or U13018 (N_13018,N_12624,N_12841);
or U13019 (N_13019,N_12034,N_12272);
and U13020 (N_13020,N_12333,N_12756);
or U13021 (N_13021,N_12292,N_12551);
xnor U13022 (N_13022,N_12101,N_12516);
and U13023 (N_13023,N_12724,N_12062);
or U13024 (N_13024,N_12987,N_12608);
xor U13025 (N_13025,N_12230,N_12832);
or U13026 (N_13026,N_12689,N_12879);
and U13027 (N_13027,N_12298,N_12894);
or U13028 (N_13028,N_12203,N_12664);
nor U13029 (N_13029,N_12008,N_12507);
or U13030 (N_13030,N_12563,N_12341);
or U13031 (N_13031,N_12305,N_12108);
xnor U13032 (N_13032,N_12026,N_12829);
nand U13033 (N_13033,N_12387,N_12121);
or U13034 (N_13034,N_12802,N_12095);
nor U13035 (N_13035,N_12836,N_12210);
nand U13036 (N_13036,N_12887,N_12959);
and U13037 (N_13037,N_12767,N_12479);
nor U13038 (N_13038,N_12499,N_12786);
xor U13039 (N_13039,N_12127,N_12198);
xor U13040 (N_13040,N_12031,N_12974);
or U13041 (N_13041,N_12816,N_12533);
nor U13042 (N_13042,N_12545,N_12484);
nand U13043 (N_13043,N_12377,N_12981);
nor U13044 (N_13044,N_12681,N_12784);
nor U13045 (N_13045,N_12726,N_12221);
xnor U13046 (N_13046,N_12104,N_12414);
or U13047 (N_13047,N_12061,N_12639);
xor U13048 (N_13048,N_12408,N_12877);
or U13049 (N_13049,N_12232,N_12171);
nand U13050 (N_13050,N_12474,N_12407);
nand U13051 (N_13051,N_12260,N_12658);
nand U13052 (N_13052,N_12081,N_12389);
nor U13053 (N_13053,N_12452,N_12092);
xor U13054 (N_13054,N_12701,N_12287);
and U13055 (N_13055,N_12274,N_12021);
xnor U13056 (N_13056,N_12134,N_12370);
nor U13057 (N_13057,N_12614,N_12483);
and U13058 (N_13058,N_12299,N_12590);
nor U13059 (N_13059,N_12692,N_12674);
xnor U13060 (N_13060,N_12466,N_12462);
and U13061 (N_13061,N_12023,N_12873);
nand U13062 (N_13062,N_12720,N_12989);
and U13063 (N_13063,N_12451,N_12025);
nand U13064 (N_13064,N_12293,N_12968);
and U13065 (N_13065,N_12368,N_12005);
and U13066 (N_13066,N_12691,N_12672);
and U13067 (N_13067,N_12991,N_12717);
nand U13068 (N_13068,N_12938,N_12177);
xnor U13069 (N_13069,N_12503,N_12901);
xnor U13070 (N_13070,N_12326,N_12337);
and U13071 (N_13071,N_12404,N_12702);
nand U13072 (N_13072,N_12772,N_12831);
xnor U13073 (N_13073,N_12911,N_12983);
xnor U13074 (N_13074,N_12956,N_12666);
and U13075 (N_13075,N_12363,N_12209);
and U13076 (N_13076,N_12584,N_12146);
or U13077 (N_13077,N_12971,N_12319);
nor U13078 (N_13078,N_12494,N_12753);
xor U13079 (N_13079,N_12160,N_12677);
or U13080 (N_13080,N_12824,N_12055);
nor U13081 (N_13081,N_12830,N_12914);
nor U13082 (N_13082,N_12890,N_12301);
and U13083 (N_13083,N_12520,N_12892);
and U13084 (N_13084,N_12910,N_12935);
xor U13085 (N_13085,N_12028,N_12510);
or U13086 (N_13086,N_12295,N_12996);
nor U13087 (N_13087,N_12626,N_12711);
and U13088 (N_13088,N_12680,N_12382);
or U13089 (N_13089,N_12509,N_12847);
or U13090 (N_13090,N_12164,N_12132);
nand U13091 (N_13091,N_12535,N_12226);
or U13092 (N_13092,N_12630,N_12058);
nor U13093 (N_13093,N_12920,N_12874);
and U13094 (N_13094,N_12436,N_12011);
and U13095 (N_13095,N_12605,N_12794);
nor U13096 (N_13096,N_12385,N_12265);
xor U13097 (N_13097,N_12978,N_12856);
xor U13098 (N_13098,N_12995,N_12641);
and U13099 (N_13099,N_12447,N_12506);
xor U13100 (N_13100,N_12827,N_12777);
or U13101 (N_13101,N_12620,N_12947);
nand U13102 (N_13102,N_12053,N_12942);
xor U13103 (N_13103,N_12788,N_12825);
or U13104 (N_13104,N_12849,N_12490);
or U13105 (N_13105,N_12477,N_12826);
nand U13106 (N_13106,N_12951,N_12040);
nor U13107 (N_13107,N_12098,N_12416);
xnor U13108 (N_13108,N_12975,N_12163);
and U13109 (N_13109,N_12000,N_12236);
nand U13110 (N_13110,N_12627,N_12478);
or U13111 (N_13111,N_12763,N_12637);
and U13112 (N_13112,N_12846,N_12603);
and U13113 (N_13113,N_12460,N_12621);
or U13114 (N_13114,N_12313,N_12747);
xor U13115 (N_13115,N_12077,N_12923);
and U13116 (N_13116,N_12315,N_12683);
and U13117 (N_13117,N_12076,N_12610);
nor U13118 (N_13118,N_12687,N_12821);
and U13119 (N_13119,N_12852,N_12165);
xnor U13120 (N_13120,N_12340,N_12530);
xnor U13121 (N_13121,N_12056,N_12515);
nor U13122 (N_13122,N_12190,N_12231);
nand U13123 (N_13123,N_12949,N_12310);
xor U13124 (N_13124,N_12379,N_12227);
and U13125 (N_13125,N_12769,N_12539);
nor U13126 (N_13126,N_12848,N_12833);
and U13127 (N_13127,N_12933,N_12659);
nor U13128 (N_13128,N_12193,N_12905);
and U13129 (N_13129,N_12517,N_12344);
and U13130 (N_13130,N_12338,N_12609);
xnor U13131 (N_13131,N_12524,N_12162);
nand U13132 (N_13132,N_12554,N_12367);
xnor U13133 (N_13133,N_12760,N_12676);
nand U13134 (N_13134,N_12569,N_12793);
nand U13135 (N_13135,N_12931,N_12789);
nor U13136 (N_13136,N_12537,N_12239);
or U13137 (N_13137,N_12454,N_12854);
or U13138 (N_13138,N_12441,N_12813);
xor U13139 (N_13139,N_12930,N_12251);
and U13140 (N_13140,N_12775,N_12449);
nor U13141 (N_13141,N_12380,N_12967);
nand U13142 (N_13142,N_12514,N_12334);
or U13143 (N_13143,N_12252,N_12270);
and U13144 (N_13144,N_12667,N_12402);
nand U13145 (N_13145,N_12668,N_12065);
and U13146 (N_13146,N_12138,N_12208);
or U13147 (N_13147,N_12762,N_12154);
xnor U13148 (N_13148,N_12858,N_12766);
nand U13149 (N_13149,N_12822,N_12534);
and U13150 (N_13150,N_12508,N_12222);
nand U13151 (N_13151,N_12851,N_12869);
and U13152 (N_13152,N_12745,N_12803);
xnor U13153 (N_13153,N_12391,N_12792);
nand U13154 (N_13154,N_12531,N_12128);
or U13155 (N_13155,N_12646,N_12078);
xnor U13156 (N_13156,N_12752,N_12502);
or U13157 (N_13157,N_12586,N_12487);
nor U13158 (N_13158,N_12913,N_12290);
nor U13159 (N_13159,N_12625,N_12107);
or U13160 (N_13160,N_12918,N_12185);
nand U13161 (N_13161,N_12872,N_12307);
xor U13162 (N_13162,N_12732,N_12882);
nand U13163 (N_13163,N_12593,N_12030);
nand U13164 (N_13164,N_12355,N_12562);
nand U13165 (N_13165,N_12424,N_12657);
xnor U13166 (N_13166,N_12728,N_12897);
xnor U13167 (N_13167,N_12100,N_12366);
nand U13168 (N_13168,N_12268,N_12468);
or U13169 (N_13169,N_12577,N_12840);
and U13170 (N_13170,N_12799,N_12597);
and U13171 (N_13171,N_12471,N_12184);
xnor U13172 (N_13172,N_12582,N_12915);
nor U13173 (N_13173,N_12348,N_12051);
nor U13174 (N_13174,N_12282,N_12392);
or U13175 (N_13175,N_12352,N_12277);
xnor U13176 (N_13176,N_12156,N_12097);
and U13177 (N_13177,N_12663,N_12926);
or U13178 (N_13178,N_12750,N_12388);
xnor U13179 (N_13179,N_12180,N_12707);
nand U13180 (N_13180,N_12445,N_12175);
nor U13181 (N_13181,N_12512,N_12511);
nor U13182 (N_13182,N_12652,N_12998);
xor U13183 (N_13183,N_12122,N_12309);
nor U13184 (N_13184,N_12264,N_12457);
nand U13185 (N_13185,N_12795,N_12757);
xnor U13186 (N_13186,N_12700,N_12089);
xor U13187 (N_13187,N_12286,N_12119);
xnor U13188 (N_13188,N_12150,N_12373);
xor U13189 (N_13189,N_12488,N_12966);
nor U13190 (N_13190,N_12188,N_12288);
xnor U13191 (N_13191,N_12126,N_12048);
nand U13192 (N_13192,N_12662,N_12759);
nor U13193 (N_13193,N_12893,N_12546);
and U13194 (N_13194,N_12665,N_12710);
nand U13195 (N_13195,N_12014,N_12013);
nand U13196 (N_13196,N_12381,N_12613);
nor U13197 (N_13197,N_12401,N_12261);
nor U13198 (N_13198,N_12331,N_12046);
and U13199 (N_13199,N_12924,N_12925);
or U13200 (N_13200,N_12525,N_12705);
and U13201 (N_13201,N_12179,N_12470);
nor U13202 (N_13202,N_12722,N_12085);
and U13203 (N_13203,N_12770,N_12741);
nand U13204 (N_13204,N_12578,N_12801);
or U13205 (N_13205,N_12623,N_12716);
nor U13206 (N_13206,N_12992,N_12505);
or U13207 (N_13207,N_12174,N_12785);
nand U13208 (N_13208,N_12999,N_12573);
nor U13209 (N_13209,N_12891,N_12853);
nand U13210 (N_13210,N_12360,N_12675);
xnor U13211 (N_13211,N_12601,N_12906);
or U13212 (N_13212,N_12304,N_12631);
nor U13213 (N_13213,N_12697,N_12482);
or U13214 (N_13214,N_12907,N_12976);
or U13215 (N_13215,N_12022,N_12117);
nor U13216 (N_13216,N_12946,N_12815);
nor U13217 (N_13217,N_12245,N_12771);
nor U13218 (N_13218,N_12839,N_12279);
or U13219 (N_13219,N_12944,N_12111);
nand U13220 (N_13220,N_12715,N_12088);
xor U13221 (N_13221,N_12467,N_12576);
or U13222 (N_13222,N_12247,N_12047);
and U13223 (N_13223,N_12489,N_12276);
nor U13224 (N_13224,N_12583,N_12280);
nand U13225 (N_13225,N_12837,N_12057);
xnor U13226 (N_13226,N_12560,N_12773);
nand U13227 (N_13227,N_12908,N_12797);
xor U13228 (N_13228,N_12860,N_12425);
or U13229 (N_13229,N_12783,N_12552);
nand U13230 (N_13230,N_12383,N_12086);
xnor U13231 (N_13231,N_12220,N_12571);
or U13232 (N_13232,N_12543,N_12725);
xor U13233 (N_13233,N_12281,N_12863);
and U13234 (N_13234,N_12339,N_12187);
and U13235 (N_13235,N_12139,N_12806);
nor U13236 (N_13236,N_12114,N_12842);
nor U13237 (N_13237,N_12730,N_12342);
xor U13238 (N_13238,N_12063,N_12384);
xnor U13239 (N_13239,N_12708,N_12776);
xnor U13240 (N_13240,N_12812,N_12589);
nor U13241 (N_13241,N_12990,N_12250);
xor U13242 (N_13242,N_12472,N_12744);
nand U13243 (N_13243,N_12645,N_12594);
and U13244 (N_13244,N_12491,N_12884);
and U13245 (N_13245,N_12258,N_12544);
xor U13246 (N_13246,N_12060,N_12001);
nand U13247 (N_13247,N_12015,N_12269);
or U13248 (N_13248,N_12575,N_12954);
nor U13249 (N_13249,N_12343,N_12176);
or U13250 (N_13250,N_12988,N_12588);
xnor U13251 (N_13251,N_12256,N_12428);
and U13252 (N_13252,N_12740,N_12093);
nand U13253 (N_13253,N_12952,N_12415);
xnor U13254 (N_13254,N_12357,N_12798);
xor U13255 (N_13255,N_12557,N_12902);
nor U13256 (N_13256,N_12818,N_12861);
nand U13257 (N_13257,N_12318,N_12066);
or U13258 (N_13258,N_12393,N_12526);
nand U13259 (N_13259,N_12410,N_12074);
nor U13260 (N_13260,N_12320,N_12653);
and U13261 (N_13261,N_12144,N_12713);
nand U13262 (N_13262,N_12969,N_12916);
nor U13263 (N_13263,N_12958,N_12591);
xor U13264 (N_13264,N_12196,N_12755);
nand U13265 (N_13265,N_12492,N_12403);
or U13266 (N_13266,N_12120,N_12754);
xnor U13267 (N_13267,N_12037,N_12585);
xor U13268 (N_13268,N_12378,N_12706);
nand U13269 (N_13269,N_12137,N_12297);
nor U13270 (N_13270,N_12810,N_12109);
and U13271 (N_13271,N_12638,N_12643);
and U13272 (N_13272,N_12400,N_12555);
xor U13273 (N_13273,N_12774,N_12033);
nand U13274 (N_13274,N_12064,N_12895);
nand U13275 (N_13275,N_12096,N_12012);
nor U13276 (N_13276,N_12746,N_12204);
xnor U13277 (N_13277,N_12296,N_12475);
and U13278 (N_13278,N_12431,N_12345);
and U13279 (N_13279,N_12473,N_12670);
xor U13280 (N_13280,N_12444,N_12070);
and U13281 (N_13281,N_12604,N_12796);
and U13282 (N_13282,N_12955,N_12729);
or U13283 (N_13283,N_12644,N_12648);
nor U13284 (N_13284,N_12413,N_12455);
and U13285 (N_13285,N_12719,N_12192);
xnor U13286 (N_13286,N_12820,N_12632);
nor U13287 (N_13287,N_12993,N_12376);
xor U13288 (N_13288,N_12386,N_12855);
xnor U13289 (N_13289,N_12237,N_12984);
nand U13290 (N_13290,N_12679,N_12587);
xnor U13291 (N_13291,N_12275,N_12718);
nand U13292 (N_13292,N_12880,N_12075);
xnor U13293 (N_13293,N_12116,N_12228);
xor U13294 (N_13294,N_12123,N_12035);
or U13295 (N_13295,N_12432,N_12496);
nand U13296 (N_13296,N_12314,N_12328);
or U13297 (N_13297,N_12636,N_12024);
or U13298 (N_13298,N_12103,N_12347);
nand U13299 (N_13299,N_12327,N_12607);
xor U13300 (N_13300,N_12422,N_12655);
xnor U13301 (N_13301,N_12405,N_12864);
xnor U13302 (N_13302,N_12397,N_12216);
nor U13303 (N_13303,N_12536,N_12936);
and U13304 (N_13304,N_12650,N_12390);
xnor U13305 (N_13305,N_12172,N_12145);
nand U13306 (N_13306,N_12838,N_12749);
nor U13307 (N_13307,N_12922,N_12500);
and U13308 (N_13308,N_12940,N_12580);
xnor U13309 (N_13309,N_12504,N_12004);
nand U13310 (N_13310,N_12278,N_12238);
nor U13311 (N_13311,N_12084,N_12302);
nand U13312 (N_13312,N_12734,N_12857);
xor U13313 (N_13313,N_12157,N_12943);
or U13314 (N_13314,N_12042,N_12291);
or U13315 (N_13315,N_12110,N_12721);
and U13316 (N_13316,N_12358,N_12090);
nor U13317 (N_13317,N_12758,N_12426);
or U13318 (N_13318,N_12254,N_12748);
or U13319 (N_13319,N_12738,N_12263);
xor U13320 (N_13320,N_12612,N_12303);
and U13321 (N_13321,N_12189,N_12029);
and U13322 (N_13322,N_12244,N_12395);
nand U13323 (N_13323,N_12495,N_12443);
or U13324 (N_13324,N_12927,N_12130);
nor U13325 (N_13325,N_12142,N_12283);
xnor U13326 (N_13326,N_12602,N_12182);
and U13327 (N_13327,N_12963,N_12972);
or U13328 (N_13328,N_12359,N_12538);
or U13329 (N_13329,N_12964,N_12235);
nor U13330 (N_13330,N_12434,N_12159);
xor U13331 (N_13331,N_12945,N_12423);
or U13332 (N_13332,N_12115,N_12181);
nor U13333 (N_13333,N_12939,N_12202);
nand U13334 (N_13334,N_12308,N_12131);
and U13335 (N_13335,N_12240,N_12871);
and U13336 (N_13336,N_12069,N_12899);
nand U13337 (N_13337,N_12417,N_12948);
and U13338 (N_13338,N_12448,N_12497);
xor U13339 (N_13339,N_12986,N_12364);
or U13340 (N_13340,N_12206,N_12805);
nand U13341 (N_13341,N_12412,N_12082);
nor U13342 (N_13342,N_12929,N_12125);
nor U13343 (N_13343,N_12017,N_12735);
or U13344 (N_13344,N_12501,N_12669);
nand U13345 (N_13345,N_12883,N_12982);
or U13346 (N_13346,N_12565,N_12465);
xnor U13347 (N_13347,N_12522,N_12962);
nor U13348 (N_13348,N_12080,N_12950);
or U13349 (N_13349,N_12259,N_12294);
nand U13350 (N_13350,N_12173,N_12731);
or U13351 (N_13351,N_12960,N_12054);
or U13352 (N_13352,N_12218,N_12018);
nor U13353 (N_13353,N_12481,N_12493);
xor U13354 (N_13354,N_12778,N_12654);
xnor U13355 (N_13355,N_12129,N_12743);
nand U13356 (N_13356,N_12814,N_12660);
xnor U13357 (N_13357,N_12889,N_12598);
xnor U13358 (N_13358,N_12225,N_12912);
xor U13359 (N_13359,N_12266,N_12709);
nor U13360 (N_13360,N_12059,N_12152);
or U13361 (N_13361,N_12678,N_12782);
xnor U13362 (N_13362,N_12486,N_12881);
or U13363 (N_13363,N_12862,N_12878);
xor U13364 (N_13364,N_12970,N_12693);
xor U13365 (N_13365,N_12106,N_12010);
nand U13366 (N_13366,N_12703,N_12723);
and U13367 (N_13367,N_12020,N_12330);
and U13368 (N_13368,N_12888,N_12273);
and U13369 (N_13369,N_12323,N_12727);
or U13370 (N_13370,N_12411,N_12306);
xor U13371 (N_13371,N_12321,N_12332);
and U13372 (N_13372,N_12807,N_12346);
and U13373 (N_13373,N_12079,N_12828);
nand U13374 (N_13374,N_12312,N_12765);
nand U13375 (N_13375,N_12934,N_12135);
xor U13376 (N_13376,N_12809,N_12568);
nor U13377 (N_13377,N_12518,N_12704);
xnor U13378 (N_13378,N_12566,N_12041);
or U13379 (N_13379,N_12197,N_12595);
nor U13380 (N_13380,N_12038,N_12761);
nand U13381 (N_13381,N_12673,N_12147);
nand U13382 (N_13382,N_12804,N_12141);
or U13383 (N_13383,N_12651,N_12438);
and U13384 (N_13384,N_12194,N_12006);
or U13385 (N_13385,N_12570,N_12205);
and U13386 (N_13386,N_12800,N_12635);
and U13387 (N_13387,N_12835,N_12480);
xnor U13388 (N_13388,N_12937,N_12325);
and U13389 (N_13389,N_12153,N_12476);
xnor U13390 (N_13390,N_12214,N_12696);
xor U13391 (N_13391,N_12167,N_12071);
nand U13392 (N_13392,N_12361,N_12979);
nor U13393 (N_13393,N_12656,N_12241);
nand U13394 (N_13394,N_12219,N_12742);
and U13395 (N_13395,N_12050,N_12567);
nand U13396 (N_13396,N_12350,N_12736);
nand U13397 (N_13397,N_12435,N_12178);
nor U13398 (N_13398,N_12087,N_12043);
and U13399 (N_13399,N_12149,N_12596);
nor U13400 (N_13400,N_12002,N_12161);
nand U13401 (N_13401,N_12542,N_12371);
or U13402 (N_13402,N_12255,N_12859);
or U13403 (N_13403,N_12211,N_12083);
and U13404 (N_13404,N_12091,N_12427);
nand U13405 (N_13405,N_12229,N_12528);
or U13406 (N_13406,N_12170,N_12136);
nor U13407 (N_13407,N_12617,N_12845);
xnor U13408 (N_13408,N_12694,N_12779);
nand U13409 (N_13409,N_12354,N_12399);
xor U13410 (N_13410,N_12550,N_12737);
or U13411 (N_13411,N_12574,N_12102);
and U13412 (N_13412,N_12875,N_12420);
xnor U13413 (N_13413,N_12985,N_12618);
or U13414 (N_13414,N_12600,N_12036);
nor U13415 (N_13415,N_12661,N_12843);
nand U13416 (N_13416,N_12699,N_12866);
nand U13417 (N_13417,N_12909,N_12634);
nor U13418 (N_13418,N_12642,N_12039);
nand U13419 (N_13419,N_12248,N_12155);
xor U13420 (N_13420,N_12356,N_12215);
xor U13421 (N_13421,N_12365,N_12876);
or U13422 (N_13422,N_12199,N_12409);
or U13423 (N_13423,N_12994,N_12168);
or U13424 (N_13424,N_12808,N_12791);
xor U13425 (N_13425,N_12374,N_12073);
nor U13426 (N_13426,N_12686,N_12553);
nor U13427 (N_13427,N_12353,N_12682);
nor U13428 (N_13428,N_12072,N_12105);
and U13429 (N_13429,N_12394,N_12739);
or U13430 (N_13430,N_12977,N_12099);
nor U13431 (N_13431,N_12823,N_12456);
or U13432 (N_13432,N_12556,N_12044);
and U13433 (N_13433,N_12885,N_12271);
and U13434 (N_13434,N_12458,N_12519);
nand U13435 (N_13435,N_12781,N_12764);
nor U13436 (N_13436,N_12207,N_12698);
xnor U13437 (N_13437,N_12581,N_12549);
xnor U13438 (N_13438,N_12440,N_12671);
or U13439 (N_13439,N_12003,N_12186);
xor U13440 (N_13440,N_12140,N_12790);
xnor U13441 (N_13441,N_12068,N_12868);
xor U13442 (N_13442,N_12817,N_12527);
nor U13443 (N_13443,N_12606,N_12300);
nor U13444 (N_13444,N_12233,N_12733);
nor U13445 (N_13445,N_12714,N_12844);
nor U13446 (N_13446,N_12558,N_12133);
and U13447 (N_13447,N_12311,N_12124);
nand U13448 (N_13448,N_12067,N_12973);
xor U13449 (N_13449,N_12253,N_12094);
nand U13450 (N_13450,N_12768,N_12684);
nand U13451 (N_13451,N_12224,N_12195);
or U13452 (N_13452,N_12523,N_12027);
xnor U13453 (N_13453,N_12961,N_12513);
nor U13454 (N_13454,N_12118,N_12201);
nor U13455 (N_13455,N_12113,N_12599);
nor U13456 (N_13456,N_12647,N_12262);
or U13457 (N_13457,N_12351,N_12249);
xor U13458 (N_13458,N_12372,N_12463);
xor U13459 (N_13459,N_12234,N_12903);
nor U13460 (N_13460,N_12561,N_12369);
nand U13461 (N_13461,N_12953,N_12941);
or U13462 (N_13462,N_12433,N_12469);
nand U13463 (N_13463,N_12362,N_12257);
nand U13464 (N_13464,N_12169,N_12316);
or U13465 (N_13465,N_12430,N_12622);
or U13466 (N_13466,N_12980,N_12439);
and U13467 (N_13467,N_12212,N_12285);
xnor U13468 (N_13468,N_12243,N_12429);
or U13469 (N_13469,N_12850,N_12112);
nand U13470 (N_13470,N_12932,N_12045);
or U13471 (N_13471,N_12965,N_12572);
or U13472 (N_13472,N_12148,N_12529);
and U13473 (N_13473,N_12865,N_12867);
or U13474 (N_13474,N_12442,N_12183);
or U13475 (N_13475,N_12217,N_12690);
xor U13476 (N_13476,N_12780,N_12151);
nand U13477 (N_13477,N_12016,N_12213);
nor U13478 (N_13478,N_12928,N_12453);
or U13479 (N_13479,N_12166,N_12521);
nand U13480 (N_13480,N_12896,N_12267);
or U13481 (N_13481,N_12336,N_12787);
or U13482 (N_13482,N_12811,N_12628);
or U13483 (N_13483,N_12032,N_12898);
nand U13484 (N_13484,N_12564,N_12957);
xnor U13485 (N_13485,N_12049,N_12009);
and U13486 (N_13486,N_12559,N_12611);
nor U13487 (N_13487,N_12547,N_12461);
nor U13488 (N_13488,N_12870,N_12329);
and U13489 (N_13489,N_12579,N_12619);
xnor U13490 (N_13490,N_12396,N_12052);
xnor U13491 (N_13491,N_12375,N_12143);
xnor U13492 (N_13492,N_12900,N_12335);
nor U13493 (N_13493,N_12322,N_12649);
nand U13494 (N_13494,N_12459,N_12904);
xor U13495 (N_13495,N_12640,N_12289);
nor U13496 (N_13496,N_12158,N_12688);
xnor U13497 (N_13497,N_12834,N_12917);
xnor U13498 (N_13498,N_12450,N_12446);
xor U13499 (N_13499,N_12548,N_12633);
xor U13500 (N_13500,N_12750,N_12089);
or U13501 (N_13501,N_12533,N_12837);
xor U13502 (N_13502,N_12490,N_12360);
or U13503 (N_13503,N_12847,N_12962);
and U13504 (N_13504,N_12815,N_12911);
and U13505 (N_13505,N_12725,N_12917);
nand U13506 (N_13506,N_12545,N_12699);
or U13507 (N_13507,N_12194,N_12839);
and U13508 (N_13508,N_12865,N_12487);
and U13509 (N_13509,N_12126,N_12854);
nor U13510 (N_13510,N_12507,N_12891);
or U13511 (N_13511,N_12442,N_12098);
xor U13512 (N_13512,N_12109,N_12993);
or U13513 (N_13513,N_12092,N_12520);
nor U13514 (N_13514,N_12949,N_12914);
xor U13515 (N_13515,N_12816,N_12333);
or U13516 (N_13516,N_12434,N_12569);
xnor U13517 (N_13517,N_12126,N_12304);
nor U13518 (N_13518,N_12003,N_12837);
or U13519 (N_13519,N_12692,N_12745);
nor U13520 (N_13520,N_12369,N_12989);
nor U13521 (N_13521,N_12330,N_12354);
xor U13522 (N_13522,N_12205,N_12705);
nor U13523 (N_13523,N_12880,N_12602);
nand U13524 (N_13524,N_12584,N_12104);
nand U13525 (N_13525,N_12025,N_12978);
nor U13526 (N_13526,N_12814,N_12883);
nand U13527 (N_13527,N_12192,N_12275);
xnor U13528 (N_13528,N_12748,N_12102);
and U13529 (N_13529,N_12546,N_12217);
nand U13530 (N_13530,N_12833,N_12502);
nor U13531 (N_13531,N_12310,N_12342);
nor U13532 (N_13532,N_12156,N_12744);
nor U13533 (N_13533,N_12295,N_12497);
xor U13534 (N_13534,N_12913,N_12229);
xnor U13535 (N_13535,N_12506,N_12925);
nor U13536 (N_13536,N_12610,N_12728);
xor U13537 (N_13537,N_12248,N_12495);
and U13538 (N_13538,N_12813,N_12068);
nand U13539 (N_13539,N_12897,N_12620);
or U13540 (N_13540,N_12528,N_12160);
or U13541 (N_13541,N_12048,N_12115);
or U13542 (N_13542,N_12686,N_12065);
nor U13543 (N_13543,N_12909,N_12229);
or U13544 (N_13544,N_12919,N_12917);
xnor U13545 (N_13545,N_12338,N_12900);
and U13546 (N_13546,N_12776,N_12238);
and U13547 (N_13547,N_12674,N_12683);
nand U13548 (N_13548,N_12615,N_12609);
or U13549 (N_13549,N_12515,N_12046);
nor U13550 (N_13550,N_12871,N_12301);
nand U13551 (N_13551,N_12715,N_12672);
or U13552 (N_13552,N_12891,N_12345);
xnor U13553 (N_13553,N_12406,N_12288);
and U13554 (N_13554,N_12592,N_12129);
nor U13555 (N_13555,N_12891,N_12644);
xor U13556 (N_13556,N_12691,N_12263);
and U13557 (N_13557,N_12367,N_12643);
nand U13558 (N_13558,N_12076,N_12356);
and U13559 (N_13559,N_12220,N_12831);
nor U13560 (N_13560,N_12679,N_12961);
xnor U13561 (N_13561,N_12768,N_12664);
and U13562 (N_13562,N_12673,N_12622);
nand U13563 (N_13563,N_12131,N_12677);
xnor U13564 (N_13564,N_12779,N_12598);
xnor U13565 (N_13565,N_12636,N_12301);
nor U13566 (N_13566,N_12025,N_12357);
or U13567 (N_13567,N_12307,N_12609);
or U13568 (N_13568,N_12285,N_12224);
nand U13569 (N_13569,N_12415,N_12224);
nand U13570 (N_13570,N_12863,N_12929);
and U13571 (N_13571,N_12955,N_12029);
or U13572 (N_13572,N_12923,N_12782);
xor U13573 (N_13573,N_12111,N_12560);
and U13574 (N_13574,N_12848,N_12783);
or U13575 (N_13575,N_12420,N_12336);
nor U13576 (N_13576,N_12588,N_12951);
or U13577 (N_13577,N_12833,N_12462);
nor U13578 (N_13578,N_12022,N_12046);
or U13579 (N_13579,N_12399,N_12967);
and U13580 (N_13580,N_12213,N_12152);
or U13581 (N_13581,N_12936,N_12784);
nand U13582 (N_13582,N_12684,N_12233);
nand U13583 (N_13583,N_12936,N_12302);
xnor U13584 (N_13584,N_12986,N_12215);
nand U13585 (N_13585,N_12929,N_12670);
and U13586 (N_13586,N_12220,N_12983);
nor U13587 (N_13587,N_12145,N_12556);
nand U13588 (N_13588,N_12027,N_12197);
or U13589 (N_13589,N_12706,N_12415);
and U13590 (N_13590,N_12860,N_12654);
and U13591 (N_13591,N_12837,N_12662);
nor U13592 (N_13592,N_12798,N_12259);
or U13593 (N_13593,N_12176,N_12813);
nand U13594 (N_13594,N_12167,N_12950);
nand U13595 (N_13595,N_12324,N_12728);
or U13596 (N_13596,N_12015,N_12571);
xor U13597 (N_13597,N_12256,N_12692);
xor U13598 (N_13598,N_12686,N_12311);
nand U13599 (N_13599,N_12578,N_12474);
or U13600 (N_13600,N_12728,N_12737);
xor U13601 (N_13601,N_12409,N_12081);
xnor U13602 (N_13602,N_12459,N_12347);
nand U13603 (N_13603,N_12442,N_12070);
nor U13604 (N_13604,N_12362,N_12661);
xnor U13605 (N_13605,N_12394,N_12017);
nor U13606 (N_13606,N_12959,N_12955);
xnor U13607 (N_13607,N_12515,N_12419);
nand U13608 (N_13608,N_12219,N_12280);
and U13609 (N_13609,N_12667,N_12108);
xnor U13610 (N_13610,N_12065,N_12389);
xnor U13611 (N_13611,N_12441,N_12910);
xor U13612 (N_13612,N_12443,N_12942);
xor U13613 (N_13613,N_12704,N_12218);
nor U13614 (N_13614,N_12459,N_12161);
and U13615 (N_13615,N_12815,N_12093);
nand U13616 (N_13616,N_12318,N_12607);
nor U13617 (N_13617,N_12551,N_12234);
nand U13618 (N_13618,N_12451,N_12488);
nor U13619 (N_13619,N_12382,N_12569);
xor U13620 (N_13620,N_12269,N_12119);
nor U13621 (N_13621,N_12735,N_12577);
nor U13622 (N_13622,N_12181,N_12547);
nand U13623 (N_13623,N_12226,N_12188);
and U13624 (N_13624,N_12190,N_12536);
and U13625 (N_13625,N_12547,N_12893);
and U13626 (N_13626,N_12192,N_12641);
xor U13627 (N_13627,N_12127,N_12578);
and U13628 (N_13628,N_12608,N_12602);
or U13629 (N_13629,N_12427,N_12189);
nor U13630 (N_13630,N_12566,N_12440);
nor U13631 (N_13631,N_12447,N_12941);
or U13632 (N_13632,N_12091,N_12596);
nand U13633 (N_13633,N_12080,N_12265);
xor U13634 (N_13634,N_12895,N_12827);
and U13635 (N_13635,N_12993,N_12076);
nand U13636 (N_13636,N_12893,N_12757);
or U13637 (N_13637,N_12931,N_12983);
xor U13638 (N_13638,N_12524,N_12986);
nand U13639 (N_13639,N_12680,N_12990);
or U13640 (N_13640,N_12193,N_12526);
xor U13641 (N_13641,N_12850,N_12422);
nand U13642 (N_13642,N_12443,N_12018);
or U13643 (N_13643,N_12327,N_12063);
nor U13644 (N_13644,N_12515,N_12623);
nor U13645 (N_13645,N_12482,N_12003);
nor U13646 (N_13646,N_12332,N_12051);
nand U13647 (N_13647,N_12676,N_12632);
xnor U13648 (N_13648,N_12538,N_12970);
nor U13649 (N_13649,N_12416,N_12693);
nor U13650 (N_13650,N_12945,N_12464);
and U13651 (N_13651,N_12689,N_12227);
xor U13652 (N_13652,N_12173,N_12400);
xnor U13653 (N_13653,N_12372,N_12469);
nand U13654 (N_13654,N_12188,N_12854);
or U13655 (N_13655,N_12271,N_12008);
or U13656 (N_13656,N_12783,N_12255);
nor U13657 (N_13657,N_12231,N_12058);
or U13658 (N_13658,N_12152,N_12159);
or U13659 (N_13659,N_12719,N_12811);
xnor U13660 (N_13660,N_12988,N_12224);
and U13661 (N_13661,N_12870,N_12323);
nor U13662 (N_13662,N_12452,N_12342);
nor U13663 (N_13663,N_12386,N_12169);
nand U13664 (N_13664,N_12957,N_12867);
and U13665 (N_13665,N_12882,N_12311);
and U13666 (N_13666,N_12757,N_12924);
nor U13667 (N_13667,N_12737,N_12587);
nor U13668 (N_13668,N_12941,N_12828);
nand U13669 (N_13669,N_12406,N_12012);
nand U13670 (N_13670,N_12726,N_12170);
or U13671 (N_13671,N_12593,N_12186);
nand U13672 (N_13672,N_12341,N_12926);
nand U13673 (N_13673,N_12010,N_12334);
and U13674 (N_13674,N_12298,N_12908);
xnor U13675 (N_13675,N_12314,N_12212);
nand U13676 (N_13676,N_12095,N_12151);
nor U13677 (N_13677,N_12663,N_12997);
xnor U13678 (N_13678,N_12515,N_12144);
nor U13679 (N_13679,N_12550,N_12640);
nand U13680 (N_13680,N_12014,N_12620);
xor U13681 (N_13681,N_12254,N_12222);
nand U13682 (N_13682,N_12684,N_12777);
nor U13683 (N_13683,N_12913,N_12982);
xor U13684 (N_13684,N_12735,N_12265);
or U13685 (N_13685,N_12435,N_12128);
and U13686 (N_13686,N_12001,N_12678);
nor U13687 (N_13687,N_12123,N_12599);
or U13688 (N_13688,N_12055,N_12520);
or U13689 (N_13689,N_12137,N_12123);
nor U13690 (N_13690,N_12184,N_12108);
and U13691 (N_13691,N_12296,N_12512);
nor U13692 (N_13692,N_12435,N_12517);
xnor U13693 (N_13693,N_12303,N_12484);
nor U13694 (N_13694,N_12000,N_12771);
and U13695 (N_13695,N_12979,N_12311);
and U13696 (N_13696,N_12284,N_12154);
nand U13697 (N_13697,N_12486,N_12284);
or U13698 (N_13698,N_12968,N_12067);
nor U13699 (N_13699,N_12994,N_12466);
or U13700 (N_13700,N_12032,N_12005);
nand U13701 (N_13701,N_12833,N_12832);
nor U13702 (N_13702,N_12157,N_12836);
xnor U13703 (N_13703,N_12052,N_12392);
and U13704 (N_13704,N_12051,N_12887);
nand U13705 (N_13705,N_12403,N_12848);
or U13706 (N_13706,N_12360,N_12732);
or U13707 (N_13707,N_12902,N_12466);
or U13708 (N_13708,N_12863,N_12162);
nor U13709 (N_13709,N_12463,N_12111);
nand U13710 (N_13710,N_12294,N_12543);
or U13711 (N_13711,N_12058,N_12802);
nand U13712 (N_13712,N_12428,N_12390);
xnor U13713 (N_13713,N_12177,N_12807);
nand U13714 (N_13714,N_12548,N_12726);
xnor U13715 (N_13715,N_12623,N_12020);
xor U13716 (N_13716,N_12204,N_12611);
and U13717 (N_13717,N_12895,N_12975);
and U13718 (N_13718,N_12700,N_12308);
xnor U13719 (N_13719,N_12020,N_12880);
or U13720 (N_13720,N_12035,N_12424);
nor U13721 (N_13721,N_12554,N_12070);
xor U13722 (N_13722,N_12313,N_12959);
xnor U13723 (N_13723,N_12437,N_12353);
nand U13724 (N_13724,N_12163,N_12277);
nor U13725 (N_13725,N_12640,N_12468);
and U13726 (N_13726,N_12012,N_12933);
nor U13727 (N_13727,N_12438,N_12213);
nand U13728 (N_13728,N_12092,N_12430);
nor U13729 (N_13729,N_12238,N_12910);
xor U13730 (N_13730,N_12542,N_12922);
nor U13731 (N_13731,N_12411,N_12272);
or U13732 (N_13732,N_12403,N_12579);
nand U13733 (N_13733,N_12975,N_12529);
or U13734 (N_13734,N_12998,N_12352);
or U13735 (N_13735,N_12261,N_12569);
xor U13736 (N_13736,N_12583,N_12498);
or U13737 (N_13737,N_12584,N_12367);
and U13738 (N_13738,N_12101,N_12124);
xnor U13739 (N_13739,N_12026,N_12038);
or U13740 (N_13740,N_12765,N_12334);
or U13741 (N_13741,N_12775,N_12013);
and U13742 (N_13742,N_12696,N_12886);
nand U13743 (N_13743,N_12895,N_12929);
nor U13744 (N_13744,N_12220,N_12363);
xnor U13745 (N_13745,N_12855,N_12782);
xnor U13746 (N_13746,N_12664,N_12420);
nor U13747 (N_13747,N_12052,N_12926);
and U13748 (N_13748,N_12008,N_12261);
or U13749 (N_13749,N_12692,N_12349);
and U13750 (N_13750,N_12855,N_12173);
nor U13751 (N_13751,N_12330,N_12297);
and U13752 (N_13752,N_12240,N_12309);
nor U13753 (N_13753,N_12919,N_12123);
nand U13754 (N_13754,N_12755,N_12271);
xnor U13755 (N_13755,N_12232,N_12788);
and U13756 (N_13756,N_12053,N_12287);
or U13757 (N_13757,N_12445,N_12583);
nor U13758 (N_13758,N_12238,N_12851);
xnor U13759 (N_13759,N_12627,N_12544);
xor U13760 (N_13760,N_12065,N_12255);
or U13761 (N_13761,N_12391,N_12052);
xor U13762 (N_13762,N_12308,N_12946);
nor U13763 (N_13763,N_12837,N_12537);
or U13764 (N_13764,N_12344,N_12133);
nand U13765 (N_13765,N_12788,N_12906);
xnor U13766 (N_13766,N_12758,N_12006);
or U13767 (N_13767,N_12091,N_12956);
or U13768 (N_13768,N_12964,N_12254);
and U13769 (N_13769,N_12996,N_12208);
and U13770 (N_13770,N_12711,N_12803);
xor U13771 (N_13771,N_12900,N_12366);
nor U13772 (N_13772,N_12647,N_12978);
xor U13773 (N_13773,N_12211,N_12263);
xor U13774 (N_13774,N_12905,N_12391);
nand U13775 (N_13775,N_12723,N_12488);
xnor U13776 (N_13776,N_12846,N_12384);
nor U13777 (N_13777,N_12068,N_12953);
nor U13778 (N_13778,N_12557,N_12702);
nor U13779 (N_13779,N_12978,N_12709);
and U13780 (N_13780,N_12481,N_12698);
and U13781 (N_13781,N_12178,N_12127);
nand U13782 (N_13782,N_12238,N_12862);
nand U13783 (N_13783,N_12578,N_12167);
and U13784 (N_13784,N_12380,N_12713);
nand U13785 (N_13785,N_12668,N_12930);
nor U13786 (N_13786,N_12509,N_12366);
xor U13787 (N_13787,N_12808,N_12794);
nor U13788 (N_13788,N_12626,N_12093);
nand U13789 (N_13789,N_12350,N_12765);
nor U13790 (N_13790,N_12818,N_12614);
nand U13791 (N_13791,N_12508,N_12051);
xnor U13792 (N_13792,N_12426,N_12604);
nor U13793 (N_13793,N_12850,N_12827);
and U13794 (N_13794,N_12830,N_12282);
or U13795 (N_13795,N_12809,N_12628);
nand U13796 (N_13796,N_12721,N_12366);
xor U13797 (N_13797,N_12232,N_12569);
and U13798 (N_13798,N_12016,N_12237);
or U13799 (N_13799,N_12113,N_12829);
nor U13800 (N_13800,N_12670,N_12910);
or U13801 (N_13801,N_12953,N_12636);
or U13802 (N_13802,N_12366,N_12803);
and U13803 (N_13803,N_12900,N_12607);
nor U13804 (N_13804,N_12030,N_12950);
or U13805 (N_13805,N_12485,N_12060);
or U13806 (N_13806,N_12826,N_12533);
or U13807 (N_13807,N_12353,N_12689);
and U13808 (N_13808,N_12474,N_12275);
nand U13809 (N_13809,N_12773,N_12569);
and U13810 (N_13810,N_12014,N_12342);
nand U13811 (N_13811,N_12885,N_12862);
nor U13812 (N_13812,N_12544,N_12976);
nand U13813 (N_13813,N_12239,N_12775);
or U13814 (N_13814,N_12929,N_12748);
xnor U13815 (N_13815,N_12255,N_12609);
or U13816 (N_13816,N_12566,N_12729);
or U13817 (N_13817,N_12785,N_12114);
nand U13818 (N_13818,N_12682,N_12814);
and U13819 (N_13819,N_12658,N_12390);
xor U13820 (N_13820,N_12748,N_12281);
or U13821 (N_13821,N_12498,N_12059);
or U13822 (N_13822,N_12053,N_12984);
nand U13823 (N_13823,N_12691,N_12950);
nand U13824 (N_13824,N_12726,N_12824);
nand U13825 (N_13825,N_12539,N_12345);
or U13826 (N_13826,N_12405,N_12743);
nor U13827 (N_13827,N_12509,N_12148);
nand U13828 (N_13828,N_12060,N_12136);
nor U13829 (N_13829,N_12734,N_12690);
xnor U13830 (N_13830,N_12541,N_12188);
nor U13831 (N_13831,N_12539,N_12618);
or U13832 (N_13832,N_12189,N_12333);
and U13833 (N_13833,N_12345,N_12081);
or U13834 (N_13834,N_12147,N_12328);
nor U13835 (N_13835,N_12348,N_12487);
or U13836 (N_13836,N_12475,N_12324);
nor U13837 (N_13837,N_12455,N_12170);
nand U13838 (N_13838,N_12335,N_12123);
and U13839 (N_13839,N_12814,N_12493);
or U13840 (N_13840,N_12894,N_12882);
and U13841 (N_13841,N_12224,N_12546);
or U13842 (N_13842,N_12897,N_12810);
xor U13843 (N_13843,N_12460,N_12976);
nand U13844 (N_13844,N_12094,N_12699);
and U13845 (N_13845,N_12250,N_12129);
nand U13846 (N_13846,N_12642,N_12779);
or U13847 (N_13847,N_12008,N_12200);
and U13848 (N_13848,N_12887,N_12910);
and U13849 (N_13849,N_12478,N_12760);
nor U13850 (N_13850,N_12396,N_12599);
nand U13851 (N_13851,N_12431,N_12089);
nand U13852 (N_13852,N_12908,N_12399);
xnor U13853 (N_13853,N_12447,N_12138);
xor U13854 (N_13854,N_12392,N_12624);
and U13855 (N_13855,N_12488,N_12199);
xnor U13856 (N_13856,N_12451,N_12288);
or U13857 (N_13857,N_12848,N_12644);
nor U13858 (N_13858,N_12111,N_12867);
xnor U13859 (N_13859,N_12121,N_12593);
nor U13860 (N_13860,N_12552,N_12239);
nand U13861 (N_13861,N_12580,N_12120);
xor U13862 (N_13862,N_12159,N_12706);
nand U13863 (N_13863,N_12198,N_12798);
xor U13864 (N_13864,N_12284,N_12046);
nor U13865 (N_13865,N_12119,N_12059);
nor U13866 (N_13866,N_12158,N_12200);
nor U13867 (N_13867,N_12294,N_12278);
and U13868 (N_13868,N_12694,N_12663);
or U13869 (N_13869,N_12966,N_12332);
and U13870 (N_13870,N_12306,N_12271);
and U13871 (N_13871,N_12268,N_12059);
nand U13872 (N_13872,N_12419,N_12851);
nor U13873 (N_13873,N_12703,N_12037);
nand U13874 (N_13874,N_12102,N_12966);
or U13875 (N_13875,N_12371,N_12895);
nor U13876 (N_13876,N_12704,N_12230);
nand U13877 (N_13877,N_12067,N_12217);
and U13878 (N_13878,N_12232,N_12371);
and U13879 (N_13879,N_12207,N_12958);
nand U13880 (N_13880,N_12315,N_12220);
or U13881 (N_13881,N_12479,N_12135);
or U13882 (N_13882,N_12025,N_12413);
nor U13883 (N_13883,N_12847,N_12720);
nor U13884 (N_13884,N_12677,N_12009);
xor U13885 (N_13885,N_12186,N_12209);
and U13886 (N_13886,N_12062,N_12387);
nor U13887 (N_13887,N_12672,N_12105);
xnor U13888 (N_13888,N_12832,N_12208);
or U13889 (N_13889,N_12364,N_12794);
or U13890 (N_13890,N_12216,N_12472);
nor U13891 (N_13891,N_12571,N_12888);
xor U13892 (N_13892,N_12688,N_12930);
nand U13893 (N_13893,N_12127,N_12358);
xor U13894 (N_13894,N_12511,N_12826);
xor U13895 (N_13895,N_12678,N_12604);
nor U13896 (N_13896,N_12180,N_12077);
or U13897 (N_13897,N_12048,N_12961);
xor U13898 (N_13898,N_12548,N_12454);
xnor U13899 (N_13899,N_12889,N_12469);
and U13900 (N_13900,N_12294,N_12613);
nor U13901 (N_13901,N_12059,N_12846);
xnor U13902 (N_13902,N_12585,N_12332);
nand U13903 (N_13903,N_12813,N_12400);
and U13904 (N_13904,N_12079,N_12204);
nand U13905 (N_13905,N_12362,N_12265);
xor U13906 (N_13906,N_12257,N_12421);
nor U13907 (N_13907,N_12179,N_12124);
xnor U13908 (N_13908,N_12171,N_12800);
and U13909 (N_13909,N_12107,N_12416);
nand U13910 (N_13910,N_12550,N_12314);
or U13911 (N_13911,N_12602,N_12635);
or U13912 (N_13912,N_12909,N_12953);
nor U13913 (N_13913,N_12828,N_12920);
and U13914 (N_13914,N_12880,N_12803);
or U13915 (N_13915,N_12476,N_12911);
nor U13916 (N_13916,N_12655,N_12222);
xnor U13917 (N_13917,N_12062,N_12265);
nand U13918 (N_13918,N_12878,N_12405);
or U13919 (N_13919,N_12966,N_12642);
or U13920 (N_13920,N_12577,N_12818);
xor U13921 (N_13921,N_12424,N_12134);
and U13922 (N_13922,N_12177,N_12225);
and U13923 (N_13923,N_12068,N_12264);
nand U13924 (N_13924,N_12420,N_12161);
nor U13925 (N_13925,N_12777,N_12357);
nor U13926 (N_13926,N_12615,N_12751);
nand U13927 (N_13927,N_12251,N_12055);
nor U13928 (N_13928,N_12031,N_12752);
and U13929 (N_13929,N_12401,N_12973);
and U13930 (N_13930,N_12658,N_12724);
xnor U13931 (N_13931,N_12560,N_12193);
nand U13932 (N_13932,N_12878,N_12796);
or U13933 (N_13933,N_12887,N_12029);
nor U13934 (N_13934,N_12843,N_12650);
nor U13935 (N_13935,N_12976,N_12513);
or U13936 (N_13936,N_12949,N_12322);
nor U13937 (N_13937,N_12007,N_12076);
and U13938 (N_13938,N_12289,N_12383);
nor U13939 (N_13939,N_12793,N_12576);
and U13940 (N_13940,N_12118,N_12657);
nand U13941 (N_13941,N_12438,N_12768);
nand U13942 (N_13942,N_12908,N_12747);
nand U13943 (N_13943,N_12896,N_12934);
or U13944 (N_13944,N_12968,N_12901);
or U13945 (N_13945,N_12855,N_12649);
or U13946 (N_13946,N_12053,N_12052);
or U13947 (N_13947,N_12327,N_12206);
and U13948 (N_13948,N_12890,N_12368);
nor U13949 (N_13949,N_12130,N_12211);
xnor U13950 (N_13950,N_12942,N_12492);
or U13951 (N_13951,N_12740,N_12945);
xnor U13952 (N_13952,N_12516,N_12410);
nor U13953 (N_13953,N_12441,N_12917);
xnor U13954 (N_13954,N_12553,N_12446);
nor U13955 (N_13955,N_12557,N_12155);
nor U13956 (N_13956,N_12659,N_12191);
or U13957 (N_13957,N_12583,N_12310);
nand U13958 (N_13958,N_12291,N_12206);
and U13959 (N_13959,N_12487,N_12223);
or U13960 (N_13960,N_12561,N_12217);
or U13961 (N_13961,N_12893,N_12705);
and U13962 (N_13962,N_12503,N_12102);
nand U13963 (N_13963,N_12430,N_12640);
or U13964 (N_13964,N_12870,N_12627);
nor U13965 (N_13965,N_12698,N_12178);
or U13966 (N_13966,N_12016,N_12192);
nand U13967 (N_13967,N_12433,N_12952);
or U13968 (N_13968,N_12900,N_12425);
xor U13969 (N_13969,N_12810,N_12691);
nor U13970 (N_13970,N_12320,N_12970);
nor U13971 (N_13971,N_12499,N_12921);
nand U13972 (N_13972,N_12687,N_12970);
and U13973 (N_13973,N_12254,N_12939);
nand U13974 (N_13974,N_12943,N_12077);
xnor U13975 (N_13975,N_12777,N_12497);
xor U13976 (N_13976,N_12992,N_12506);
nand U13977 (N_13977,N_12315,N_12897);
nand U13978 (N_13978,N_12657,N_12417);
xor U13979 (N_13979,N_12011,N_12368);
or U13980 (N_13980,N_12862,N_12192);
nand U13981 (N_13981,N_12437,N_12219);
and U13982 (N_13982,N_12932,N_12122);
nand U13983 (N_13983,N_12650,N_12488);
and U13984 (N_13984,N_12919,N_12518);
xor U13985 (N_13985,N_12154,N_12013);
nor U13986 (N_13986,N_12749,N_12310);
or U13987 (N_13987,N_12000,N_12811);
nor U13988 (N_13988,N_12502,N_12672);
or U13989 (N_13989,N_12682,N_12607);
xor U13990 (N_13990,N_12470,N_12398);
xnor U13991 (N_13991,N_12481,N_12185);
xnor U13992 (N_13992,N_12898,N_12655);
and U13993 (N_13993,N_12977,N_12925);
nor U13994 (N_13994,N_12883,N_12964);
nor U13995 (N_13995,N_12326,N_12673);
or U13996 (N_13996,N_12573,N_12129);
or U13997 (N_13997,N_12914,N_12769);
and U13998 (N_13998,N_12841,N_12296);
nor U13999 (N_13999,N_12905,N_12377);
or U14000 (N_14000,N_13788,N_13635);
and U14001 (N_14001,N_13947,N_13114);
nand U14002 (N_14002,N_13809,N_13026);
nor U14003 (N_14003,N_13608,N_13410);
nor U14004 (N_14004,N_13983,N_13991);
xor U14005 (N_14005,N_13133,N_13127);
xor U14006 (N_14006,N_13209,N_13703);
or U14007 (N_14007,N_13370,N_13261);
and U14008 (N_14008,N_13413,N_13101);
and U14009 (N_14009,N_13585,N_13920);
nor U14010 (N_14010,N_13633,N_13817);
nand U14011 (N_14011,N_13134,N_13303);
nand U14012 (N_14012,N_13486,N_13362);
nand U14013 (N_14013,N_13769,N_13269);
nor U14014 (N_14014,N_13218,N_13859);
nand U14015 (N_14015,N_13091,N_13989);
nor U14016 (N_14016,N_13067,N_13847);
nor U14017 (N_14017,N_13924,N_13137);
and U14018 (N_14018,N_13524,N_13036);
xnor U14019 (N_14019,N_13008,N_13699);
and U14020 (N_14020,N_13141,N_13746);
nand U14021 (N_14021,N_13429,N_13874);
or U14022 (N_14022,N_13994,N_13182);
nor U14023 (N_14023,N_13157,N_13088);
and U14024 (N_14024,N_13241,N_13946);
nand U14025 (N_14025,N_13339,N_13588);
nor U14026 (N_14026,N_13568,N_13822);
nand U14027 (N_14027,N_13276,N_13499);
nor U14028 (N_14028,N_13371,N_13293);
and U14029 (N_14029,N_13461,N_13501);
nand U14030 (N_14030,N_13135,N_13298);
xnor U14031 (N_14031,N_13318,N_13709);
xor U14032 (N_14032,N_13054,N_13727);
and U14033 (N_14033,N_13735,N_13476);
xor U14034 (N_14034,N_13776,N_13651);
and U14035 (N_14035,N_13684,N_13708);
xnor U14036 (N_14036,N_13502,N_13344);
or U14037 (N_14037,N_13216,N_13985);
nand U14038 (N_14038,N_13129,N_13556);
xor U14039 (N_14039,N_13740,N_13849);
nor U14040 (N_14040,N_13372,N_13052);
nand U14041 (N_14041,N_13995,N_13836);
nand U14042 (N_14042,N_13056,N_13870);
and U14043 (N_14043,N_13470,N_13719);
nand U14044 (N_14044,N_13662,N_13104);
or U14045 (N_14045,N_13522,N_13926);
nor U14046 (N_14046,N_13916,N_13966);
nor U14047 (N_14047,N_13123,N_13225);
xnor U14048 (N_14048,N_13488,N_13144);
and U14049 (N_14049,N_13627,N_13017);
and U14050 (N_14050,N_13047,N_13971);
nor U14051 (N_14051,N_13235,N_13059);
nor U14052 (N_14052,N_13265,N_13640);
or U14053 (N_14053,N_13351,N_13748);
and U14054 (N_14054,N_13866,N_13935);
and U14055 (N_14055,N_13083,N_13458);
or U14056 (N_14056,N_13644,N_13698);
xor U14057 (N_14057,N_13508,N_13271);
nand U14058 (N_14058,N_13234,N_13661);
xor U14059 (N_14059,N_13530,N_13595);
or U14060 (N_14060,N_13469,N_13162);
xor U14061 (N_14061,N_13944,N_13405);
or U14062 (N_14062,N_13035,N_13259);
nand U14063 (N_14063,N_13593,N_13895);
xor U14064 (N_14064,N_13840,N_13291);
or U14065 (N_14065,N_13041,N_13366);
and U14066 (N_14066,N_13664,N_13007);
xnor U14067 (N_14067,N_13672,N_13602);
or U14068 (N_14068,N_13093,N_13065);
nor U14069 (N_14069,N_13215,N_13019);
xor U14070 (N_14070,N_13519,N_13030);
nand U14071 (N_14071,N_13306,N_13714);
or U14072 (N_14072,N_13782,N_13625);
xor U14073 (N_14073,N_13029,N_13611);
nor U14074 (N_14074,N_13579,N_13004);
xnor U14075 (N_14075,N_13732,N_13489);
xor U14076 (N_14076,N_13348,N_13089);
and U14077 (N_14077,N_13353,N_13069);
or U14078 (N_14078,N_13781,N_13108);
xnor U14079 (N_14079,N_13958,N_13024);
and U14080 (N_14080,N_13598,N_13242);
or U14081 (N_14081,N_13592,N_13365);
or U14082 (N_14082,N_13987,N_13941);
or U14083 (N_14083,N_13409,N_13221);
or U14084 (N_14084,N_13542,N_13424);
xnor U14085 (N_14085,N_13045,N_13889);
nand U14086 (N_14086,N_13620,N_13773);
nor U14087 (N_14087,N_13658,N_13667);
or U14088 (N_14088,N_13175,N_13465);
nor U14089 (N_14089,N_13331,N_13569);
and U14090 (N_14090,N_13867,N_13034);
and U14091 (N_14091,N_13752,N_13285);
nor U14092 (N_14092,N_13578,N_13712);
or U14093 (N_14093,N_13884,N_13444);
xnor U14094 (N_14094,N_13280,N_13184);
or U14095 (N_14095,N_13388,N_13220);
xnor U14096 (N_14096,N_13233,N_13070);
nand U14097 (N_14097,N_13230,N_13566);
nor U14098 (N_14098,N_13287,N_13976);
or U14099 (N_14099,N_13132,N_13915);
xnor U14100 (N_14100,N_13784,N_13309);
nor U14101 (N_14101,N_13440,N_13140);
or U14102 (N_14102,N_13479,N_13606);
nor U14103 (N_14103,N_13316,N_13142);
or U14104 (N_14104,N_13828,N_13996);
and U14105 (N_14105,N_13415,N_13350);
or U14106 (N_14106,N_13616,N_13912);
nor U14107 (N_14107,N_13167,N_13484);
nor U14108 (N_14108,N_13443,N_13990);
and U14109 (N_14109,N_13016,N_13503);
or U14110 (N_14110,N_13552,N_13792);
nor U14111 (N_14111,N_13838,N_13072);
nor U14112 (N_14112,N_13613,N_13927);
and U14113 (N_14113,N_13624,N_13222);
and U14114 (N_14114,N_13082,N_13441);
nand U14115 (N_14115,N_13892,N_13675);
nand U14116 (N_14116,N_13655,N_13452);
and U14117 (N_14117,N_13487,N_13948);
nand U14118 (N_14118,N_13749,N_13124);
and U14119 (N_14119,N_13610,N_13189);
or U14120 (N_14120,N_13361,N_13978);
and U14121 (N_14121,N_13492,N_13854);
nand U14122 (N_14122,N_13956,N_13724);
or U14123 (N_14123,N_13904,N_13374);
nor U14124 (N_14124,N_13205,N_13320);
or U14125 (N_14125,N_13071,N_13737);
or U14126 (N_14126,N_13553,N_13097);
nand U14127 (N_14127,N_13964,N_13571);
nor U14128 (N_14128,N_13637,N_13360);
nor U14129 (N_14129,N_13422,N_13993);
and U14130 (N_14130,N_13536,N_13560);
or U14131 (N_14131,N_13621,N_13177);
nand U14132 (N_14132,N_13497,N_13587);
nor U14133 (N_14133,N_13880,N_13378);
xnor U14134 (N_14134,N_13063,N_13206);
and U14135 (N_14135,N_13283,N_13393);
or U14136 (N_14136,N_13406,N_13831);
or U14137 (N_14137,N_13934,N_13011);
or U14138 (N_14138,N_13367,N_13921);
xor U14139 (N_14139,N_13025,N_13918);
xor U14140 (N_14140,N_13818,N_13686);
and U14141 (N_14141,N_13023,N_13357);
nor U14142 (N_14142,N_13582,N_13952);
and U14143 (N_14143,N_13473,N_13173);
and U14144 (N_14144,N_13901,N_13191);
or U14145 (N_14145,N_13323,N_13474);
or U14146 (N_14146,N_13053,N_13228);
nor U14147 (N_14147,N_13196,N_13005);
or U14148 (N_14148,N_13329,N_13418);
xor U14149 (N_14149,N_13211,N_13647);
nand U14150 (N_14150,N_13538,N_13103);
xnor U14151 (N_14151,N_13594,N_13885);
xnor U14152 (N_14152,N_13738,N_13389);
or U14153 (N_14153,N_13080,N_13893);
or U14154 (N_14154,N_13660,N_13801);
and U14155 (N_14155,N_13117,N_13403);
nand U14156 (N_14156,N_13858,N_13012);
nor U14157 (N_14157,N_13882,N_13970);
and U14158 (N_14158,N_13439,N_13273);
nand U14159 (N_14159,N_13693,N_13210);
nand U14160 (N_14160,N_13645,N_13256);
nand U14161 (N_14161,N_13744,N_13813);
nand U14162 (N_14162,N_13623,N_13028);
xnor U14163 (N_14163,N_13301,N_13617);
xnor U14164 (N_14164,N_13176,N_13187);
or U14165 (N_14165,N_13515,N_13500);
nor U14166 (N_14166,N_13816,N_13546);
and U14167 (N_14167,N_13003,N_13148);
or U14168 (N_14168,N_13495,N_13972);
or U14169 (N_14169,N_13800,N_13251);
and U14170 (N_14170,N_13919,N_13482);
nor U14171 (N_14171,N_13857,N_13827);
nand U14172 (N_14172,N_13512,N_13670);
nand U14173 (N_14173,N_13483,N_13346);
nand U14174 (N_14174,N_13426,N_13853);
nand U14175 (N_14175,N_13720,N_13668);
xnor U14176 (N_14176,N_13887,N_13201);
nand U14177 (N_14177,N_13094,N_13757);
and U14178 (N_14178,N_13058,N_13965);
or U14179 (N_14179,N_13669,N_13150);
nor U14180 (N_14180,N_13730,N_13710);
and U14181 (N_14181,N_13758,N_13706);
nor U14182 (N_14182,N_13506,N_13629);
and U14183 (N_14183,N_13020,N_13636);
nand U14184 (N_14184,N_13525,N_13729);
nor U14185 (N_14185,N_13061,N_13183);
nand U14186 (N_14186,N_13288,N_13986);
xnor U14187 (N_14187,N_13363,N_13478);
nor U14188 (N_14188,N_13257,N_13463);
xnor U14189 (N_14189,N_13604,N_13988);
or U14190 (N_14190,N_13618,N_13208);
nor U14191 (N_14191,N_13244,N_13181);
nand U14192 (N_14192,N_13281,N_13355);
nor U14193 (N_14193,N_13060,N_13615);
nor U14194 (N_14194,N_13475,N_13819);
nor U14195 (N_14195,N_13879,N_13711);
or U14196 (N_14196,N_13352,N_13953);
nor U14197 (N_14197,N_13431,N_13833);
or U14198 (N_14198,N_13539,N_13683);
nand U14199 (N_14199,N_13928,N_13899);
xnor U14200 (N_14200,N_13428,N_13731);
nor U14201 (N_14201,N_13286,N_13632);
and U14202 (N_14202,N_13421,N_13505);
nor U14203 (N_14203,N_13697,N_13881);
nand U14204 (N_14204,N_13120,N_13414);
and U14205 (N_14205,N_13159,N_13382);
nand U14206 (N_14206,N_13938,N_13435);
xnor U14207 (N_14207,N_13340,N_13681);
nand U14208 (N_14208,N_13464,N_13533);
and U14209 (N_14209,N_13314,N_13704);
or U14210 (N_14210,N_13835,N_13638);
and U14211 (N_14211,N_13619,N_13518);
or U14212 (N_14212,N_13573,N_13095);
or U14213 (N_14213,N_13839,N_13315);
and U14214 (N_14214,N_13564,N_13805);
or U14215 (N_14215,N_13407,N_13334);
nand U14216 (N_14216,N_13513,N_13327);
or U14217 (N_14217,N_13420,N_13128);
and U14218 (N_14218,N_13923,N_13364);
nand U14219 (N_14219,N_13937,N_13649);
and U14220 (N_14220,N_13375,N_13680);
and U14221 (N_14221,N_13785,N_13961);
or U14222 (N_14222,N_13547,N_13846);
xor U14223 (N_14223,N_13674,N_13778);
and U14224 (N_14224,N_13570,N_13814);
or U14225 (N_14225,N_13434,N_13600);
xor U14226 (N_14226,N_13736,N_13721);
and U14227 (N_14227,N_13417,N_13490);
nor U14228 (N_14228,N_13678,N_13010);
or U14229 (N_14229,N_13147,N_13081);
nand U14230 (N_14230,N_13018,N_13102);
or U14231 (N_14231,N_13368,N_13641);
nor U14232 (N_14232,N_13027,N_13380);
nor U14233 (N_14233,N_13759,N_13349);
or U14234 (N_14234,N_13305,N_13888);
xnor U14235 (N_14235,N_13743,N_13969);
nand U14236 (N_14236,N_13171,N_13541);
xnor U14237 (N_14237,N_13158,N_13180);
and U14238 (N_14238,N_13436,N_13931);
nand U14239 (N_14239,N_13260,N_13116);
xnor U14240 (N_14240,N_13913,N_13009);
nor U14241 (N_14241,N_13718,N_13526);
and U14242 (N_14242,N_13454,N_13110);
nor U14243 (N_14243,N_13877,N_13717);
nand U14244 (N_14244,N_13197,N_13358);
or U14245 (N_14245,N_13455,N_13385);
nor U14246 (N_14246,N_13219,N_13255);
nand U14247 (N_14247,N_13015,N_13654);
nand U14248 (N_14248,N_13467,N_13466);
or U14249 (N_14249,N_13107,N_13832);
nor U14250 (N_14250,N_13540,N_13902);
nor U14251 (N_14251,N_13238,N_13263);
or U14252 (N_14252,N_13307,N_13317);
xor U14253 (N_14253,N_13622,N_13087);
xor U14254 (N_14254,N_13278,N_13325);
or U14255 (N_14255,N_13580,N_13377);
xnor U14256 (N_14256,N_13328,N_13745);
nor U14257 (N_14257,N_13558,N_13726);
and U14258 (N_14258,N_13125,N_13174);
or U14259 (N_14259,N_13830,N_13237);
or U14260 (N_14260,N_13170,N_13433);
nor U14261 (N_14261,N_13359,N_13051);
and U14262 (N_14262,N_13868,N_13311);
nor U14263 (N_14263,N_13815,N_13064);
nand U14264 (N_14264,N_13650,N_13543);
and U14265 (N_14265,N_13974,N_13797);
and U14266 (N_14266,N_13762,N_13930);
or U14267 (N_14267,N_13396,N_13576);
or U14268 (N_14268,N_13666,N_13826);
or U14269 (N_14269,N_13341,N_13481);
xnor U14270 (N_14270,N_13875,N_13977);
or U14271 (N_14271,N_13825,N_13723);
xor U14272 (N_14272,N_13925,N_13354);
nand U14273 (N_14273,N_13262,N_13224);
xnor U14274 (N_14274,N_13696,N_13922);
and U14275 (N_14275,N_13545,N_13472);
nand U14276 (N_14276,N_13450,N_13949);
and U14277 (N_14277,N_13430,N_13936);
nor U14278 (N_14278,N_13597,N_13863);
xnor U14279 (N_14279,N_13575,N_13105);
nand U14280 (N_14280,N_13692,N_13628);
or U14281 (N_14281,N_13783,N_13014);
nand U14282 (N_14282,N_13551,N_13292);
xnor U14283 (N_14283,N_13214,N_13549);
xnor U14284 (N_14284,N_13240,N_13510);
xnor U14285 (N_14285,N_13079,N_13336);
nor U14286 (N_14286,N_13663,N_13734);
or U14287 (N_14287,N_13185,N_13299);
or U14288 (N_14288,N_13894,N_13939);
xor U14289 (N_14289,N_13485,N_13462);
nand U14290 (N_14290,N_13775,N_13728);
and U14291 (N_14291,N_13810,N_13852);
xor U14292 (N_14292,N_13639,N_13153);
nand U14293 (N_14293,N_13954,N_13445);
or U14294 (N_14294,N_13275,N_13856);
xor U14295 (N_14295,N_13790,N_13038);
and U14296 (N_14296,N_13226,N_13249);
and U14297 (N_14297,N_13824,N_13400);
xnor U14298 (N_14298,N_13131,N_13691);
xor U14299 (N_14299,N_13685,N_13152);
xnor U14300 (N_14300,N_13277,N_13399);
nor U14301 (N_14301,N_13033,N_13607);
nor U14302 (N_14302,N_13121,N_13213);
nor U14303 (N_14303,N_13767,N_13077);
and U14304 (N_14304,N_13113,N_13779);
nor U14305 (N_14305,N_13166,N_13160);
and U14306 (N_14306,N_13761,N_13246);
and U14307 (N_14307,N_13957,N_13119);
nand U14308 (N_14308,N_13855,N_13006);
or U14309 (N_14309,N_13715,N_13448);
or U14310 (N_14310,N_13254,N_13044);
nor U14311 (N_14311,N_13284,N_13890);
xor U14312 (N_14312,N_13872,N_13126);
nor U14313 (N_14313,N_13338,N_13544);
and U14314 (N_14314,N_13747,N_13772);
or U14315 (N_14315,N_13653,N_13626);
and U14316 (N_14316,N_13907,N_13155);
or U14317 (N_14317,N_13862,N_13751);
nand U14318 (N_14318,N_13139,N_13771);
or U14319 (N_14319,N_13130,N_13217);
nand U14320 (N_14320,N_13270,N_13193);
and U14321 (N_14321,N_13308,N_13973);
xnor U14322 (N_14322,N_13085,N_13803);
xor U14323 (N_14323,N_13195,N_13701);
nor U14324 (N_14324,N_13416,N_13532);
or U14325 (N_14325,N_13457,N_13178);
xor U14326 (N_14326,N_13192,N_13106);
xor U14327 (N_14327,N_13268,N_13982);
xnor U14328 (N_14328,N_13212,N_13200);
nand U14329 (N_14329,N_13310,N_13387);
xnor U14330 (N_14330,N_13459,N_13172);
or U14331 (N_14331,N_13203,N_13031);
nor U14332 (N_14332,N_13820,N_13806);
and U14333 (N_14333,N_13911,N_13092);
xnor U14334 (N_14334,N_13793,N_13202);
nor U14335 (N_14335,N_13204,N_13343);
nor U14336 (N_14336,N_13282,N_13634);
xnor U14337 (N_14337,N_13313,N_13860);
nor U14338 (N_14338,N_13401,N_13295);
or U14339 (N_14339,N_13046,N_13766);
nand U14340 (N_14340,N_13562,N_13848);
and U14341 (N_14341,N_13040,N_13086);
nand U14342 (N_14342,N_13909,N_13245);
or U14343 (N_14343,N_13565,N_13402);
nor U14344 (N_14344,N_13321,N_13186);
and U14345 (N_14345,N_13446,N_13770);
nor U14346 (N_14346,N_13886,N_13154);
or U14347 (N_14347,N_13665,N_13567);
and U14348 (N_14348,N_13391,N_13851);
nand U14349 (N_14349,N_13707,N_13844);
nor U14350 (N_14350,N_13962,N_13646);
xnor U14351 (N_14351,N_13039,N_13021);
xor U14352 (N_14352,N_13190,N_13821);
and U14353 (N_14353,N_13574,N_13774);
xnor U14354 (N_14354,N_13705,N_13763);
nand U14355 (N_14355,N_13850,N_13764);
nand U14356 (N_14356,N_13643,N_13427);
xnor U14357 (N_14357,N_13369,N_13337);
nor U14358 (N_14358,N_13531,N_13753);
and U14359 (N_14359,N_13100,N_13161);
xor U14360 (N_14360,N_13968,N_13933);
and U14361 (N_14361,N_13768,N_13940);
and U14362 (N_14362,N_13236,N_13043);
xor U14363 (N_14363,N_13975,N_13605);
or U14364 (N_14364,N_13168,N_13842);
or U14365 (N_14365,N_13905,N_13980);
xor U14366 (N_14366,N_13294,N_13062);
xnor U14367 (N_14367,N_13789,N_13312);
nor U14368 (N_14368,N_13381,N_13798);
nor U14369 (N_14369,N_13090,N_13164);
nand U14370 (N_14370,N_13165,N_13612);
xor U14371 (N_14371,N_13676,N_13347);
xor U14372 (N_14372,N_13013,N_13794);
or U14373 (N_14373,N_13599,N_13279);
or U14374 (N_14374,N_13050,N_13335);
nand U14375 (N_14375,N_13873,N_13412);
and U14376 (N_14376,N_13432,N_13841);
and U14377 (N_14377,N_13494,N_13042);
and U14378 (N_14378,N_13741,N_13900);
nor U14379 (N_14379,N_13419,N_13871);
and U14380 (N_14380,N_13659,N_13967);
or U14381 (N_14381,N_13504,N_13631);
and U14382 (N_14382,N_13322,N_13002);
and U14383 (N_14383,N_13345,N_13796);
or U14384 (N_14384,N_13442,N_13390);
nor U14385 (N_14385,N_13861,N_13138);
and U14386 (N_14386,N_13845,N_13514);
or U14387 (N_14387,N_13603,N_13507);
xnor U14388 (N_14388,N_13756,N_13955);
or U14389 (N_14389,N_13266,N_13332);
nand U14390 (N_14390,N_13929,N_13523);
or U14391 (N_14391,N_13520,N_13289);
or U14392 (N_14392,N_13906,N_13397);
xnor U14393 (N_14393,N_13229,N_13297);
nor U14394 (N_14394,N_13992,N_13075);
and U14395 (N_14395,N_13657,N_13115);
nor U14396 (N_14396,N_13823,N_13146);
or U14397 (N_14397,N_13959,N_13267);
nor U14398 (N_14398,N_13795,N_13437);
and U14399 (N_14399,N_13496,N_13725);
or U14400 (N_14400,N_13979,N_13787);
and U14401 (N_14401,N_13791,N_13066);
nor U14402 (N_14402,N_13742,N_13000);
nand U14403 (N_14403,N_13807,N_13098);
nor U14404 (N_14404,N_13780,N_13702);
or U14405 (N_14405,N_13865,N_13917);
xor U14406 (N_14406,N_13843,N_13074);
and U14407 (N_14407,N_13384,N_13755);
nand U14408 (N_14408,N_13557,N_13689);
nand U14409 (N_14409,N_13333,N_13057);
xor U14410 (N_14410,N_13648,N_13754);
xor U14411 (N_14411,N_13760,N_13583);
and U14412 (N_14412,N_13527,N_13883);
xor U14413 (N_14413,N_13156,N_13682);
or U14414 (N_14414,N_13777,N_13837);
xnor U14415 (N_14415,N_13687,N_13572);
nand U14416 (N_14416,N_13690,N_13078);
and U14417 (N_14417,N_13163,N_13324);
nand U14418 (N_14418,N_13136,N_13111);
and U14419 (N_14419,N_13404,N_13897);
xnor U14420 (N_14420,N_13480,N_13194);
or U14421 (N_14421,N_13555,N_13561);
or U14422 (N_14422,N_13739,N_13491);
or U14423 (N_14423,N_13581,N_13232);
nand U14424 (N_14424,N_13910,N_13673);
nor U14425 (N_14425,N_13614,N_13149);
and U14426 (N_14426,N_13584,N_13438);
nor U14427 (N_14427,N_13394,N_13250);
or U14428 (N_14428,N_13356,N_13534);
and U14429 (N_14429,N_13722,N_13804);
xnor U14430 (N_14430,N_13477,N_13383);
or U14431 (N_14431,N_13589,N_13932);
nor U14432 (N_14432,N_13786,N_13373);
or U14433 (N_14433,N_13528,N_13498);
and U14434 (N_14434,N_13652,N_13049);
or U14435 (N_14435,N_13223,N_13151);
and U14436 (N_14436,N_13945,N_13898);
xnor U14437 (N_14437,N_13342,N_13908);
nor U14438 (N_14438,N_13960,N_13521);
and U14439 (N_14439,N_13876,N_13290);
or U14440 (N_14440,N_13272,N_13516);
xnor U14441 (N_14441,N_13984,N_13529);
and U14442 (N_14442,N_13963,N_13379);
and U14443 (N_14443,N_13330,N_13799);
nor U14444 (N_14444,N_13981,N_13998);
xnor U14445 (N_14445,N_13112,N_13022);
nor U14446 (N_14446,N_13447,N_13109);
and U14447 (N_14447,N_13037,N_13577);
or U14448 (N_14448,N_13942,N_13207);
nand U14449 (N_14449,N_13231,N_13386);
nand U14450 (N_14450,N_13864,N_13453);
nand U14451 (N_14451,N_13713,N_13188);
and U14452 (N_14452,N_13449,N_13198);
or U14453 (N_14453,N_13914,N_13609);
xnor U14454 (N_14454,N_13411,N_13300);
nand U14455 (N_14455,N_13563,N_13559);
and U14456 (N_14456,N_13048,N_13997);
nor U14457 (N_14457,N_13258,N_13550);
xnor U14458 (N_14458,N_13055,N_13099);
xor U14459 (N_14459,N_13319,N_13765);
nor U14460 (N_14460,N_13951,N_13239);
nor U14461 (N_14461,N_13252,N_13468);
and U14462 (N_14462,N_13247,N_13392);
nand U14463 (N_14463,N_13829,N_13802);
nor U14464 (N_14464,N_13096,N_13517);
nand U14465 (N_14465,N_13834,N_13811);
and U14466 (N_14466,N_13145,N_13423);
nand U14467 (N_14467,N_13642,N_13591);
nand U14468 (N_14468,N_13999,N_13535);
or U14469 (N_14469,N_13199,N_13700);
nand U14470 (N_14470,N_13425,N_13253);
nor U14471 (N_14471,N_13326,N_13032);
nand U14472 (N_14472,N_13903,N_13671);
nand U14473 (N_14473,N_13073,N_13896);
xnor U14474 (N_14474,N_13076,N_13227);
nor U14475 (N_14475,N_13398,N_13274);
nand U14476 (N_14476,N_13586,N_13304);
nand U14477 (N_14477,N_13068,N_13296);
nand U14478 (N_14478,N_13302,N_13812);
xnor U14479 (N_14479,N_13590,N_13716);
nor U14480 (N_14480,N_13084,N_13001);
and U14481 (N_14481,N_13118,N_13733);
xnor U14482 (N_14482,N_13679,N_13248);
or U14483 (N_14483,N_13630,N_13891);
and U14484 (N_14484,N_13869,N_13548);
nor U14485 (N_14485,N_13808,N_13376);
nor U14486 (N_14486,N_13656,N_13471);
or U14487 (N_14487,N_13601,N_13596);
or U14488 (N_14488,N_13456,N_13169);
or U14489 (N_14489,N_13694,N_13179);
and U14490 (N_14490,N_13677,N_13408);
or U14491 (N_14491,N_13243,N_13460);
or U14492 (N_14492,N_13950,N_13493);
nor U14493 (N_14493,N_13395,N_13537);
nor U14494 (N_14494,N_13695,N_13143);
or U14495 (N_14495,N_13688,N_13511);
nand U14496 (N_14496,N_13943,N_13122);
or U14497 (N_14497,N_13264,N_13554);
and U14498 (N_14498,N_13878,N_13451);
or U14499 (N_14499,N_13750,N_13509);
and U14500 (N_14500,N_13361,N_13695);
nand U14501 (N_14501,N_13546,N_13065);
xor U14502 (N_14502,N_13103,N_13709);
and U14503 (N_14503,N_13149,N_13021);
and U14504 (N_14504,N_13085,N_13135);
nor U14505 (N_14505,N_13380,N_13079);
xor U14506 (N_14506,N_13473,N_13464);
nor U14507 (N_14507,N_13611,N_13443);
xnor U14508 (N_14508,N_13859,N_13488);
xnor U14509 (N_14509,N_13430,N_13738);
nor U14510 (N_14510,N_13823,N_13878);
nor U14511 (N_14511,N_13988,N_13398);
nand U14512 (N_14512,N_13704,N_13750);
nor U14513 (N_14513,N_13457,N_13301);
or U14514 (N_14514,N_13324,N_13944);
xor U14515 (N_14515,N_13861,N_13291);
xnor U14516 (N_14516,N_13727,N_13534);
xnor U14517 (N_14517,N_13952,N_13318);
and U14518 (N_14518,N_13867,N_13816);
or U14519 (N_14519,N_13613,N_13700);
nand U14520 (N_14520,N_13784,N_13700);
nor U14521 (N_14521,N_13707,N_13022);
or U14522 (N_14522,N_13393,N_13840);
nor U14523 (N_14523,N_13892,N_13149);
and U14524 (N_14524,N_13752,N_13851);
or U14525 (N_14525,N_13937,N_13272);
and U14526 (N_14526,N_13059,N_13654);
or U14527 (N_14527,N_13684,N_13565);
nor U14528 (N_14528,N_13531,N_13885);
nand U14529 (N_14529,N_13523,N_13118);
or U14530 (N_14530,N_13906,N_13430);
or U14531 (N_14531,N_13380,N_13875);
xnor U14532 (N_14532,N_13930,N_13075);
xor U14533 (N_14533,N_13234,N_13169);
nand U14534 (N_14534,N_13794,N_13619);
nor U14535 (N_14535,N_13356,N_13532);
or U14536 (N_14536,N_13825,N_13861);
and U14537 (N_14537,N_13833,N_13170);
and U14538 (N_14538,N_13562,N_13093);
nor U14539 (N_14539,N_13937,N_13725);
nor U14540 (N_14540,N_13109,N_13735);
or U14541 (N_14541,N_13557,N_13551);
nand U14542 (N_14542,N_13049,N_13391);
or U14543 (N_14543,N_13924,N_13835);
xnor U14544 (N_14544,N_13581,N_13042);
nor U14545 (N_14545,N_13016,N_13331);
nor U14546 (N_14546,N_13177,N_13692);
or U14547 (N_14547,N_13941,N_13382);
nand U14548 (N_14548,N_13163,N_13229);
and U14549 (N_14549,N_13295,N_13044);
nand U14550 (N_14550,N_13889,N_13103);
nand U14551 (N_14551,N_13511,N_13193);
and U14552 (N_14552,N_13372,N_13378);
and U14553 (N_14553,N_13577,N_13575);
nand U14554 (N_14554,N_13345,N_13405);
nor U14555 (N_14555,N_13463,N_13610);
nor U14556 (N_14556,N_13455,N_13468);
nand U14557 (N_14557,N_13230,N_13636);
xor U14558 (N_14558,N_13215,N_13516);
nor U14559 (N_14559,N_13263,N_13166);
xor U14560 (N_14560,N_13821,N_13237);
or U14561 (N_14561,N_13793,N_13657);
nand U14562 (N_14562,N_13996,N_13177);
nor U14563 (N_14563,N_13268,N_13862);
nand U14564 (N_14564,N_13871,N_13691);
nand U14565 (N_14565,N_13358,N_13714);
and U14566 (N_14566,N_13566,N_13973);
nor U14567 (N_14567,N_13045,N_13957);
nand U14568 (N_14568,N_13044,N_13346);
or U14569 (N_14569,N_13695,N_13152);
xnor U14570 (N_14570,N_13576,N_13031);
nand U14571 (N_14571,N_13734,N_13454);
nand U14572 (N_14572,N_13914,N_13932);
xor U14573 (N_14573,N_13650,N_13751);
nor U14574 (N_14574,N_13582,N_13425);
xnor U14575 (N_14575,N_13418,N_13182);
or U14576 (N_14576,N_13520,N_13531);
nor U14577 (N_14577,N_13749,N_13668);
or U14578 (N_14578,N_13613,N_13068);
and U14579 (N_14579,N_13772,N_13636);
xor U14580 (N_14580,N_13096,N_13437);
nor U14581 (N_14581,N_13969,N_13764);
nand U14582 (N_14582,N_13884,N_13528);
nand U14583 (N_14583,N_13044,N_13088);
nand U14584 (N_14584,N_13439,N_13354);
and U14585 (N_14585,N_13037,N_13954);
and U14586 (N_14586,N_13809,N_13172);
nand U14587 (N_14587,N_13145,N_13996);
and U14588 (N_14588,N_13979,N_13471);
and U14589 (N_14589,N_13747,N_13949);
or U14590 (N_14590,N_13456,N_13462);
and U14591 (N_14591,N_13616,N_13174);
xnor U14592 (N_14592,N_13228,N_13064);
nor U14593 (N_14593,N_13149,N_13576);
xnor U14594 (N_14594,N_13433,N_13128);
or U14595 (N_14595,N_13510,N_13276);
nand U14596 (N_14596,N_13981,N_13638);
nor U14597 (N_14597,N_13666,N_13790);
nand U14598 (N_14598,N_13138,N_13373);
and U14599 (N_14599,N_13630,N_13561);
xnor U14600 (N_14600,N_13454,N_13386);
nor U14601 (N_14601,N_13861,N_13559);
or U14602 (N_14602,N_13109,N_13252);
nor U14603 (N_14603,N_13759,N_13061);
nor U14604 (N_14604,N_13008,N_13275);
nor U14605 (N_14605,N_13268,N_13828);
or U14606 (N_14606,N_13723,N_13567);
or U14607 (N_14607,N_13178,N_13889);
xor U14608 (N_14608,N_13791,N_13888);
and U14609 (N_14609,N_13236,N_13257);
or U14610 (N_14610,N_13709,N_13180);
nor U14611 (N_14611,N_13918,N_13534);
and U14612 (N_14612,N_13706,N_13243);
nand U14613 (N_14613,N_13997,N_13829);
and U14614 (N_14614,N_13094,N_13770);
xnor U14615 (N_14615,N_13869,N_13799);
nor U14616 (N_14616,N_13780,N_13949);
nand U14617 (N_14617,N_13283,N_13473);
xnor U14618 (N_14618,N_13481,N_13282);
nand U14619 (N_14619,N_13156,N_13240);
nand U14620 (N_14620,N_13863,N_13670);
and U14621 (N_14621,N_13235,N_13031);
or U14622 (N_14622,N_13644,N_13957);
xor U14623 (N_14623,N_13895,N_13784);
xor U14624 (N_14624,N_13901,N_13903);
and U14625 (N_14625,N_13143,N_13674);
and U14626 (N_14626,N_13005,N_13865);
nor U14627 (N_14627,N_13486,N_13974);
and U14628 (N_14628,N_13291,N_13977);
and U14629 (N_14629,N_13943,N_13251);
nand U14630 (N_14630,N_13259,N_13189);
nor U14631 (N_14631,N_13162,N_13555);
xor U14632 (N_14632,N_13977,N_13127);
xnor U14633 (N_14633,N_13942,N_13384);
nor U14634 (N_14634,N_13426,N_13099);
xnor U14635 (N_14635,N_13630,N_13523);
and U14636 (N_14636,N_13520,N_13024);
nand U14637 (N_14637,N_13437,N_13397);
xnor U14638 (N_14638,N_13617,N_13703);
nor U14639 (N_14639,N_13230,N_13223);
xnor U14640 (N_14640,N_13712,N_13925);
xor U14641 (N_14641,N_13854,N_13868);
nand U14642 (N_14642,N_13757,N_13814);
or U14643 (N_14643,N_13005,N_13746);
and U14644 (N_14644,N_13455,N_13291);
or U14645 (N_14645,N_13726,N_13293);
nand U14646 (N_14646,N_13876,N_13366);
or U14647 (N_14647,N_13007,N_13851);
nor U14648 (N_14648,N_13514,N_13167);
nand U14649 (N_14649,N_13990,N_13069);
and U14650 (N_14650,N_13783,N_13596);
and U14651 (N_14651,N_13272,N_13849);
nand U14652 (N_14652,N_13605,N_13071);
nand U14653 (N_14653,N_13569,N_13937);
xnor U14654 (N_14654,N_13956,N_13506);
or U14655 (N_14655,N_13364,N_13740);
nand U14656 (N_14656,N_13612,N_13016);
nor U14657 (N_14657,N_13482,N_13767);
nand U14658 (N_14658,N_13647,N_13272);
or U14659 (N_14659,N_13827,N_13148);
or U14660 (N_14660,N_13496,N_13655);
xnor U14661 (N_14661,N_13646,N_13164);
or U14662 (N_14662,N_13619,N_13104);
nand U14663 (N_14663,N_13732,N_13169);
nor U14664 (N_14664,N_13342,N_13845);
and U14665 (N_14665,N_13742,N_13880);
nor U14666 (N_14666,N_13977,N_13178);
and U14667 (N_14667,N_13326,N_13597);
nand U14668 (N_14668,N_13060,N_13809);
nor U14669 (N_14669,N_13263,N_13394);
nand U14670 (N_14670,N_13640,N_13308);
or U14671 (N_14671,N_13675,N_13836);
and U14672 (N_14672,N_13415,N_13086);
nand U14673 (N_14673,N_13876,N_13951);
nor U14674 (N_14674,N_13089,N_13771);
nand U14675 (N_14675,N_13416,N_13822);
or U14676 (N_14676,N_13374,N_13545);
xor U14677 (N_14677,N_13986,N_13672);
and U14678 (N_14678,N_13853,N_13773);
and U14679 (N_14679,N_13144,N_13191);
nand U14680 (N_14680,N_13993,N_13961);
nand U14681 (N_14681,N_13497,N_13235);
or U14682 (N_14682,N_13752,N_13315);
nor U14683 (N_14683,N_13594,N_13591);
nor U14684 (N_14684,N_13776,N_13147);
and U14685 (N_14685,N_13595,N_13541);
nand U14686 (N_14686,N_13813,N_13305);
xnor U14687 (N_14687,N_13609,N_13312);
and U14688 (N_14688,N_13771,N_13661);
nand U14689 (N_14689,N_13649,N_13119);
nor U14690 (N_14690,N_13372,N_13155);
and U14691 (N_14691,N_13763,N_13759);
xor U14692 (N_14692,N_13248,N_13875);
nand U14693 (N_14693,N_13130,N_13092);
or U14694 (N_14694,N_13969,N_13904);
nand U14695 (N_14695,N_13808,N_13382);
xor U14696 (N_14696,N_13928,N_13404);
xor U14697 (N_14697,N_13755,N_13115);
or U14698 (N_14698,N_13984,N_13092);
xor U14699 (N_14699,N_13573,N_13704);
nor U14700 (N_14700,N_13693,N_13885);
xnor U14701 (N_14701,N_13409,N_13894);
or U14702 (N_14702,N_13243,N_13999);
and U14703 (N_14703,N_13302,N_13006);
and U14704 (N_14704,N_13491,N_13020);
nand U14705 (N_14705,N_13893,N_13985);
xnor U14706 (N_14706,N_13105,N_13127);
xnor U14707 (N_14707,N_13852,N_13691);
or U14708 (N_14708,N_13562,N_13769);
nor U14709 (N_14709,N_13962,N_13031);
and U14710 (N_14710,N_13592,N_13131);
nor U14711 (N_14711,N_13880,N_13506);
and U14712 (N_14712,N_13858,N_13718);
nand U14713 (N_14713,N_13741,N_13698);
or U14714 (N_14714,N_13696,N_13018);
nand U14715 (N_14715,N_13330,N_13543);
xnor U14716 (N_14716,N_13937,N_13955);
xor U14717 (N_14717,N_13179,N_13479);
nand U14718 (N_14718,N_13230,N_13983);
and U14719 (N_14719,N_13456,N_13432);
xnor U14720 (N_14720,N_13047,N_13544);
or U14721 (N_14721,N_13943,N_13801);
nor U14722 (N_14722,N_13119,N_13843);
and U14723 (N_14723,N_13515,N_13583);
xor U14724 (N_14724,N_13076,N_13493);
xnor U14725 (N_14725,N_13887,N_13873);
and U14726 (N_14726,N_13596,N_13071);
nand U14727 (N_14727,N_13930,N_13619);
and U14728 (N_14728,N_13373,N_13689);
nand U14729 (N_14729,N_13313,N_13804);
xnor U14730 (N_14730,N_13989,N_13946);
xnor U14731 (N_14731,N_13590,N_13571);
and U14732 (N_14732,N_13918,N_13118);
nand U14733 (N_14733,N_13380,N_13810);
or U14734 (N_14734,N_13791,N_13337);
nor U14735 (N_14735,N_13233,N_13503);
nor U14736 (N_14736,N_13748,N_13039);
nand U14737 (N_14737,N_13407,N_13379);
and U14738 (N_14738,N_13308,N_13951);
xor U14739 (N_14739,N_13648,N_13876);
xnor U14740 (N_14740,N_13123,N_13005);
nand U14741 (N_14741,N_13742,N_13285);
nand U14742 (N_14742,N_13983,N_13338);
xor U14743 (N_14743,N_13617,N_13139);
xor U14744 (N_14744,N_13885,N_13936);
nand U14745 (N_14745,N_13624,N_13036);
or U14746 (N_14746,N_13226,N_13291);
nand U14747 (N_14747,N_13933,N_13853);
and U14748 (N_14748,N_13114,N_13490);
nand U14749 (N_14749,N_13039,N_13484);
or U14750 (N_14750,N_13736,N_13150);
xnor U14751 (N_14751,N_13424,N_13734);
xnor U14752 (N_14752,N_13817,N_13493);
and U14753 (N_14753,N_13686,N_13937);
or U14754 (N_14754,N_13348,N_13140);
nand U14755 (N_14755,N_13940,N_13262);
nand U14756 (N_14756,N_13924,N_13708);
xor U14757 (N_14757,N_13203,N_13735);
or U14758 (N_14758,N_13632,N_13027);
nand U14759 (N_14759,N_13035,N_13735);
nor U14760 (N_14760,N_13648,N_13481);
or U14761 (N_14761,N_13805,N_13319);
and U14762 (N_14762,N_13626,N_13464);
xnor U14763 (N_14763,N_13312,N_13679);
nand U14764 (N_14764,N_13435,N_13349);
nor U14765 (N_14765,N_13193,N_13825);
and U14766 (N_14766,N_13832,N_13064);
nand U14767 (N_14767,N_13379,N_13828);
and U14768 (N_14768,N_13010,N_13654);
nand U14769 (N_14769,N_13324,N_13129);
nor U14770 (N_14770,N_13958,N_13159);
or U14771 (N_14771,N_13524,N_13576);
xor U14772 (N_14772,N_13779,N_13662);
nor U14773 (N_14773,N_13338,N_13805);
xnor U14774 (N_14774,N_13771,N_13065);
and U14775 (N_14775,N_13456,N_13793);
xor U14776 (N_14776,N_13343,N_13353);
nor U14777 (N_14777,N_13149,N_13467);
xnor U14778 (N_14778,N_13245,N_13417);
xnor U14779 (N_14779,N_13609,N_13999);
nor U14780 (N_14780,N_13216,N_13484);
or U14781 (N_14781,N_13923,N_13163);
nand U14782 (N_14782,N_13408,N_13051);
nand U14783 (N_14783,N_13723,N_13460);
nor U14784 (N_14784,N_13327,N_13506);
nand U14785 (N_14785,N_13484,N_13741);
and U14786 (N_14786,N_13996,N_13201);
and U14787 (N_14787,N_13215,N_13862);
and U14788 (N_14788,N_13650,N_13829);
nand U14789 (N_14789,N_13639,N_13511);
nand U14790 (N_14790,N_13676,N_13917);
xor U14791 (N_14791,N_13487,N_13508);
or U14792 (N_14792,N_13354,N_13992);
xor U14793 (N_14793,N_13359,N_13071);
and U14794 (N_14794,N_13526,N_13579);
nor U14795 (N_14795,N_13991,N_13385);
nand U14796 (N_14796,N_13299,N_13007);
nor U14797 (N_14797,N_13751,N_13359);
nand U14798 (N_14798,N_13052,N_13098);
nand U14799 (N_14799,N_13370,N_13218);
xnor U14800 (N_14800,N_13759,N_13305);
and U14801 (N_14801,N_13036,N_13855);
nor U14802 (N_14802,N_13406,N_13275);
or U14803 (N_14803,N_13619,N_13324);
nand U14804 (N_14804,N_13657,N_13959);
or U14805 (N_14805,N_13928,N_13299);
and U14806 (N_14806,N_13683,N_13074);
nand U14807 (N_14807,N_13436,N_13572);
nand U14808 (N_14808,N_13861,N_13858);
nand U14809 (N_14809,N_13369,N_13956);
nor U14810 (N_14810,N_13586,N_13488);
nor U14811 (N_14811,N_13346,N_13457);
nand U14812 (N_14812,N_13025,N_13223);
and U14813 (N_14813,N_13560,N_13548);
nor U14814 (N_14814,N_13552,N_13798);
and U14815 (N_14815,N_13091,N_13715);
or U14816 (N_14816,N_13270,N_13795);
or U14817 (N_14817,N_13799,N_13214);
and U14818 (N_14818,N_13807,N_13293);
xor U14819 (N_14819,N_13021,N_13477);
nand U14820 (N_14820,N_13406,N_13434);
xor U14821 (N_14821,N_13387,N_13377);
and U14822 (N_14822,N_13511,N_13632);
or U14823 (N_14823,N_13046,N_13758);
nor U14824 (N_14824,N_13054,N_13649);
nor U14825 (N_14825,N_13060,N_13223);
and U14826 (N_14826,N_13046,N_13274);
and U14827 (N_14827,N_13614,N_13275);
nor U14828 (N_14828,N_13350,N_13559);
nand U14829 (N_14829,N_13399,N_13101);
nor U14830 (N_14830,N_13920,N_13570);
xnor U14831 (N_14831,N_13001,N_13945);
and U14832 (N_14832,N_13550,N_13646);
nand U14833 (N_14833,N_13788,N_13398);
or U14834 (N_14834,N_13263,N_13758);
or U14835 (N_14835,N_13510,N_13935);
nand U14836 (N_14836,N_13607,N_13450);
nand U14837 (N_14837,N_13805,N_13342);
xor U14838 (N_14838,N_13213,N_13666);
and U14839 (N_14839,N_13082,N_13710);
nand U14840 (N_14840,N_13160,N_13508);
or U14841 (N_14841,N_13077,N_13543);
xnor U14842 (N_14842,N_13466,N_13095);
or U14843 (N_14843,N_13552,N_13157);
or U14844 (N_14844,N_13365,N_13304);
nand U14845 (N_14845,N_13527,N_13391);
xor U14846 (N_14846,N_13408,N_13558);
nor U14847 (N_14847,N_13664,N_13856);
nand U14848 (N_14848,N_13632,N_13205);
and U14849 (N_14849,N_13464,N_13325);
xnor U14850 (N_14850,N_13979,N_13162);
xnor U14851 (N_14851,N_13364,N_13951);
or U14852 (N_14852,N_13164,N_13914);
xnor U14853 (N_14853,N_13956,N_13091);
or U14854 (N_14854,N_13633,N_13978);
xnor U14855 (N_14855,N_13110,N_13614);
xnor U14856 (N_14856,N_13813,N_13233);
or U14857 (N_14857,N_13339,N_13733);
xnor U14858 (N_14858,N_13791,N_13641);
nand U14859 (N_14859,N_13889,N_13373);
or U14860 (N_14860,N_13691,N_13575);
nor U14861 (N_14861,N_13237,N_13530);
and U14862 (N_14862,N_13208,N_13533);
nor U14863 (N_14863,N_13203,N_13354);
nor U14864 (N_14864,N_13873,N_13043);
and U14865 (N_14865,N_13054,N_13489);
or U14866 (N_14866,N_13690,N_13592);
xor U14867 (N_14867,N_13010,N_13053);
and U14868 (N_14868,N_13329,N_13812);
or U14869 (N_14869,N_13057,N_13923);
and U14870 (N_14870,N_13540,N_13626);
or U14871 (N_14871,N_13976,N_13395);
nor U14872 (N_14872,N_13992,N_13699);
nor U14873 (N_14873,N_13623,N_13936);
nand U14874 (N_14874,N_13466,N_13012);
nor U14875 (N_14875,N_13262,N_13994);
nand U14876 (N_14876,N_13330,N_13672);
and U14877 (N_14877,N_13404,N_13248);
nor U14878 (N_14878,N_13662,N_13210);
or U14879 (N_14879,N_13318,N_13243);
xor U14880 (N_14880,N_13483,N_13156);
or U14881 (N_14881,N_13452,N_13071);
or U14882 (N_14882,N_13125,N_13483);
or U14883 (N_14883,N_13481,N_13925);
and U14884 (N_14884,N_13200,N_13081);
nor U14885 (N_14885,N_13653,N_13437);
and U14886 (N_14886,N_13005,N_13675);
or U14887 (N_14887,N_13693,N_13334);
nand U14888 (N_14888,N_13008,N_13842);
xor U14889 (N_14889,N_13044,N_13438);
and U14890 (N_14890,N_13623,N_13265);
nor U14891 (N_14891,N_13243,N_13070);
nor U14892 (N_14892,N_13588,N_13334);
nor U14893 (N_14893,N_13583,N_13216);
and U14894 (N_14894,N_13999,N_13150);
xnor U14895 (N_14895,N_13280,N_13889);
nor U14896 (N_14896,N_13523,N_13762);
nand U14897 (N_14897,N_13186,N_13118);
nand U14898 (N_14898,N_13727,N_13502);
nor U14899 (N_14899,N_13324,N_13011);
xnor U14900 (N_14900,N_13139,N_13297);
nand U14901 (N_14901,N_13700,N_13127);
xor U14902 (N_14902,N_13922,N_13491);
nand U14903 (N_14903,N_13336,N_13241);
nor U14904 (N_14904,N_13849,N_13696);
nor U14905 (N_14905,N_13656,N_13318);
or U14906 (N_14906,N_13025,N_13809);
or U14907 (N_14907,N_13082,N_13170);
and U14908 (N_14908,N_13026,N_13960);
or U14909 (N_14909,N_13150,N_13095);
nor U14910 (N_14910,N_13729,N_13889);
or U14911 (N_14911,N_13645,N_13760);
nor U14912 (N_14912,N_13328,N_13256);
nor U14913 (N_14913,N_13815,N_13676);
or U14914 (N_14914,N_13538,N_13371);
or U14915 (N_14915,N_13271,N_13340);
nor U14916 (N_14916,N_13825,N_13875);
xor U14917 (N_14917,N_13721,N_13723);
nor U14918 (N_14918,N_13258,N_13909);
nor U14919 (N_14919,N_13517,N_13961);
nand U14920 (N_14920,N_13115,N_13687);
and U14921 (N_14921,N_13361,N_13782);
and U14922 (N_14922,N_13287,N_13699);
nand U14923 (N_14923,N_13954,N_13665);
nor U14924 (N_14924,N_13958,N_13411);
nor U14925 (N_14925,N_13720,N_13714);
nand U14926 (N_14926,N_13661,N_13156);
or U14927 (N_14927,N_13523,N_13742);
nand U14928 (N_14928,N_13135,N_13419);
xnor U14929 (N_14929,N_13365,N_13416);
nand U14930 (N_14930,N_13985,N_13503);
and U14931 (N_14931,N_13343,N_13244);
nand U14932 (N_14932,N_13097,N_13394);
nor U14933 (N_14933,N_13241,N_13762);
xnor U14934 (N_14934,N_13762,N_13431);
nor U14935 (N_14935,N_13893,N_13271);
xnor U14936 (N_14936,N_13224,N_13996);
xor U14937 (N_14937,N_13908,N_13152);
or U14938 (N_14938,N_13370,N_13008);
nand U14939 (N_14939,N_13857,N_13850);
nor U14940 (N_14940,N_13548,N_13143);
xnor U14941 (N_14941,N_13415,N_13220);
xor U14942 (N_14942,N_13506,N_13250);
xor U14943 (N_14943,N_13014,N_13123);
nand U14944 (N_14944,N_13493,N_13129);
nor U14945 (N_14945,N_13093,N_13388);
and U14946 (N_14946,N_13420,N_13262);
nor U14947 (N_14947,N_13908,N_13264);
nor U14948 (N_14948,N_13291,N_13721);
and U14949 (N_14949,N_13187,N_13799);
nor U14950 (N_14950,N_13787,N_13700);
xnor U14951 (N_14951,N_13688,N_13105);
and U14952 (N_14952,N_13493,N_13847);
xor U14953 (N_14953,N_13541,N_13854);
nor U14954 (N_14954,N_13718,N_13213);
nand U14955 (N_14955,N_13502,N_13844);
or U14956 (N_14956,N_13776,N_13901);
xnor U14957 (N_14957,N_13889,N_13908);
nand U14958 (N_14958,N_13193,N_13005);
xor U14959 (N_14959,N_13699,N_13339);
nor U14960 (N_14960,N_13334,N_13692);
or U14961 (N_14961,N_13455,N_13224);
or U14962 (N_14962,N_13393,N_13223);
nand U14963 (N_14963,N_13437,N_13291);
or U14964 (N_14964,N_13192,N_13055);
nor U14965 (N_14965,N_13265,N_13599);
or U14966 (N_14966,N_13121,N_13830);
nor U14967 (N_14967,N_13504,N_13560);
or U14968 (N_14968,N_13559,N_13865);
nand U14969 (N_14969,N_13865,N_13992);
nor U14970 (N_14970,N_13132,N_13619);
or U14971 (N_14971,N_13868,N_13560);
or U14972 (N_14972,N_13385,N_13724);
xnor U14973 (N_14973,N_13250,N_13210);
and U14974 (N_14974,N_13930,N_13717);
xnor U14975 (N_14975,N_13565,N_13077);
nand U14976 (N_14976,N_13176,N_13537);
xor U14977 (N_14977,N_13783,N_13599);
and U14978 (N_14978,N_13826,N_13246);
and U14979 (N_14979,N_13080,N_13662);
nor U14980 (N_14980,N_13122,N_13212);
and U14981 (N_14981,N_13337,N_13984);
xnor U14982 (N_14982,N_13944,N_13969);
nor U14983 (N_14983,N_13456,N_13883);
nand U14984 (N_14984,N_13013,N_13632);
xor U14985 (N_14985,N_13226,N_13478);
nand U14986 (N_14986,N_13468,N_13591);
xor U14987 (N_14987,N_13428,N_13408);
and U14988 (N_14988,N_13587,N_13172);
nand U14989 (N_14989,N_13559,N_13620);
and U14990 (N_14990,N_13917,N_13722);
and U14991 (N_14991,N_13951,N_13998);
and U14992 (N_14992,N_13758,N_13940);
and U14993 (N_14993,N_13479,N_13381);
and U14994 (N_14994,N_13811,N_13178);
xnor U14995 (N_14995,N_13109,N_13335);
and U14996 (N_14996,N_13102,N_13764);
xor U14997 (N_14997,N_13083,N_13459);
or U14998 (N_14998,N_13244,N_13495);
xor U14999 (N_14999,N_13788,N_13063);
xnor U15000 (N_15000,N_14103,N_14084);
nand U15001 (N_15001,N_14726,N_14698);
and U15002 (N_15002,N_14023,N_14685);
nor U15003 (N_15003,N_14937,N_14274);
and U15004 (N_15004,N_14936,N_14615);
or U15005 (N_15005,N_14846,N_14580);
xnor U15006 (N_15006,N_14840,N_14695);
xor U15007 (N_15007,N_14659,N_14096);
or U15008 (N_15008,N_14683,N_14102);
nor U15009 (N_15009,N_14110,N_14073);
xor U15010 (N_15010,N_14980,N_14199);
and U15011 (N_15011,N_14884,N_14144);
nand U15012 (N_15012,N_14140,N_14829);
nand U15013 (N_15013,N_14126,N_14043);
nor U15014 (N_15014,N_14155,N_14069);
or U15015 (N_15015,N_14582,N_14774);
nor U15016 (N_15016,N_14879,N_14215);
nor U15017 (N_15017,N_14762,N_14117);
and U15018 (N_15018,N_14721,N_14598);
or U15019 (N_15019,N_14260,N_14709);
and U15020 (N_15020,N_14636,N_14836);
xor U15021 (N_15021,N_14597,N_14730);
nand U15022 (N_15022,N_14862,N_14603);
nand U15023 (N_15023,N_14401,N_14910);
nand U15024 (N_15024,N_14358,N_14923);
or U15025 (N_15025,N_14429,N_14901);
xor U15026 (N_15026,N_14185,N_14254);
and U15027 (N_15027,N_14444,N_14978);
or U15028 (N_15028,N_14784,N_14166);
nor U15029 (N_15029,N_14236,N_14844);
and U15030 (N_15030,N_14228,N_14875);
nand U15031 (N_15031,N_14489,N_14543);
or U15032 (N_15032,N_14684,N_14523);
and U15033 (N_15033,N_14116,N_14336);
or U15034 (N_15034,N_14115,N_14176);
xor U15035 (N_15035,N_14055,N_14586);
xor U15036 (N_15036,N_14499,N_14389);
xor U15037 (N_15037,N_14682,N_14864);
nor U15038 (N_15038,N_14807,N_14677);
nand U15039 (N_15039,N_14061,N_14893);
nand U15040 (N_15040,N_14371,N_14468);
and U15041 (N_15041,N_14241,N_14922);
or U15042 (N_15042,N_14259,N_14793);
and U15043 (N_15043,N_14307,N_14814);
nand U15044 (N_15044,N_14510,N_14347);
xor U15045 (N_15045,N_14273,N_14506);
or U15046 (N_15046,N_14609,N_14189);
nand U15047 (N_15047,N_14781,N_14817);
and U15048 (N_15048,N_14513,N_14294);
nand U15049 (N_15049,N_14338,N_14042);
xor U15050 (N_15050,N_14000,N_14383);
nor U15051 (N_15051,N_14153,N_14789);
or U15052 (N_15052,N_14127,N_14146);
or U15053 (N_15053,N_14595,N_14749);
nand U15054 (N_15054,N_14617,N_14822);
nand U15055 (N_15055,N_14594,N_14778);
and U15056 (N_15056,N_14145,N_14492);
nand U15057 (N_15057,N_14183,N_14812);
nor U15058 (N_15058,N_14442,N_14613);
nand U15059 (N_15059,N_14452,N_14841);
or U15060 (N_15060,N_14987,N_14099);
nor U15061 (N_15061,N_14856,N_14415);
and U15062 (N_15062,N_14370,N_14995);
or U15063 (N_15063,N_14854,N_14293);
or U15064 (N_15064,N_14960,N_14471);
xor U15065 (N_15065,N_14038,N_14083);
nor U15066 (N_15066,N_14093,N_14625);
xor U15067 (N_15067,N_14971,N_14122);
nand U15068 (N_15068,N_14138,N_14006);
and U15069 (N_15069,N_14114,N_14249);
nand U15070 (N_15070,N_14424,N_14328);
nand U15071 (N_15071,N_14342,N_14426);
nor U15072 (N_15072,N_14213,N_14818);
nor U15073 (N_15073,N_14515,N_14410);
or U15074 (N_15074,N_14802,N_14877);
or U15075 (N_15075,N_14903,N_14712);
or U15076 (N_15076,N_14128,N_14390);
nor U15077 (N_15077,N_14231,N_14160);
or U15078 (N_15078,N_14958,N_14962);
xor U15079 (N_15079,N_14795,N_14212);
or U15080 (N_15080,N_14743,N_14137);
nor U15081 (N_15081,N_14378,N_14188);
nor U15082 (N_15082,N_14197,N_14640);
xnor U15083 (N_15083,N_14696,N_14425);
nor U15084 (N_15084,N_14981,N_14039);
nor U15085 (N_15085,N_14885,N_14238);
nor U15086 (N_15086,N_14407,N_14644);
xnor U15087 (N_15087,N_14041,N_14275);
and U15088 (N_15088,N_14505,N_14806);
xor U15089 (N_15089,N_14654,N_14939);
xor U15090 (N_15090,N_14965,N_14159);
nor U15091 (N_15091,N_14728,N_14217);
nor U15092 (N_15092,N_14230,N_14917);
xor U15093 (N_15093,N_14930,N_14690);
and U15094 (N_15094,N_14905,N_14966);
and U15095 (N_15095,N_14037,N_14310);
nand U15096 (N_15096,N_14150,N_14758);
xnor U15097 (N_15097,N_14869,N_14356);
nor U15098 (N_15098,N_14895,N_14926);
and U15099 (N_15099,N_14266,N_14060);
and U15100 (N_15100,N_14797,N_14693);
nand U15101 (N_15101,N_14196,N_14141);
nor U15102 (N_15102,N_14479,N_14279);
and U15103 (N_15103,N_14172,N_14202);
or U15104 (N_15104,N_14898,N_14081);
and U15105 (N_15105,N_14193,N_14337);
xor U15106 (N_15106,N_14933,N_14999);
xnor U15107 (N_15107,N_14450,N_14020);
nand U15108 (N_15108,N_14349,N_14932);
nand U15109 (N_15109,N_14831,N_14894);
xnor U15110 (N_15110,N_14092,N_14950);
nand U15111 (N_15111,N_14400,N_14803);
or U15112 (N_15112,N_14233,N_14628);
nor U15113 (N_15113,N_14972,N_14245);
or U15114 (N_15114,N_14470,N_14437);
nand U15115 (N_15115,N_14427,N_14668);
nor U15116 (N_15116,N_14641,N_14514);
nand U15117 (N_15117,N_14168,N_14255);
nor U15118 (N_15118,N_14573,N_14610);
nand U15119 (N_15119,N_14123,N_14033);
nor U15120 (N_15120,N_14148,N_14462);
nand U15121 (N_15121,N_14970,N_14624);
or U15122 (N_15122,N_14741,N_14568);
or U15123 (N_15123,N_14344,N_14572);
or U15124 (N_15124,N_14301,N_14171);
xnor U15125 (N_15125,N_14843,N_14333);
xnor U15126 (N_15126,N_14334,N_14482);
or U15127 (N_15127,N_14395,N_14511);
and U15128 (N_15128,N_14820,N_14634);
nor U15129 (N_15129,N_14710,N_14291);
nor U15130 (N_15130,N_14873,N_14512);
or U15131 (N_15131,N_14441,N_14085);
xnor U15132 (N_15132,N_14218,N_14821);
nor U15133 (N_15133,N_14056,N_14621);
or U15134 (N_15134,N_14453,N_14780);
and U15135 (N_15135,N_14527,N_14439);
nor U15136 (N_15136,N_14203,N_14941);
and U15137 (N_15137,N_14012,N_14318);
nand U15138 (N_15138,N_14013,N_14044);
nand U15139 (N_15139,N_14054,N_14147);
nor U15140 (N_15140,N_14554,N_14475);
nor U15141 (N_15141,N_14469,N_14714);
and U15142 (N_15142,N_14626,N_14742);
nand U15143 (N_15143,N_14062,N_14913);
xor U15144 (N_15144,N_14379,N_14849);
xnor U15145 (N_15145,N_14436,N_14773);
and U15146 (N_15146,N_14216,N_14352);
nand U15147 (N_15147,N_14911,N_14267);
and U15148 (N_15148,N_14772,N_14645);
or U15149 (N_15149,N_14558,N_14067);
nand U15150 (N_15150,N_14767,N_14974);
nand U15151 (N_15151,N_14252,N_14919);
xnor U15152 (N_15152,N_14248,N_14385);
nand U15153 (N_15153,N_14018,N_14764);
xor U15154 (N_15154,N_14495,N_14285);
nand U15155 (N_15155,N_14048,N_14057);
nand U15156 (N_15156,N_14483,N_14465);
xor U15157 (N_15157,N_14906,N_14459);
and U15158 (N_15158,N_14244,N_14736);
nand U15159 (N_15159,N_14566,N_14364);
or U15160 (N_15160,N_14768,N_14237);
and U15161 (N_15161,N_14559,N_14718);
or U15162 (N_15162,N_14263,N_14480);
xnor U15163 (N_15163,N_14232,N_14394);
xnor U15164 (N_15164,N_14181,N_14766);
or U15165 (N_15165,N_14763,N_14107);
nand U15166 (N_15166,N_14221,N_14297);
xnor U15167 (N_15167,N_14963,N_14642);
and U15168 (N_15168,N_14614,N_14946);
or U15169 (N_15169,N_14493,N_14143);
xor U15170 (N_15170,N_14417,N_14320);
nor U15171 (N_15171,N_14920,N_14687);
or U15172 (N_15172,N_14791,N_14019);
nand U15173 (N_15173,N_14516,N_14757);
or U15174 (N_15174,N_14992,N_14694);
xnor U15175 (N_15175,N_14938,N_14487);
and U15176 (N_15176,N_14868,N_14375);
and U15177 (N_15177,N_14646,N_14440);
nor U15178 (N_15178,N_14957,N_14961);
and U15179 (N_15179,N_14177,N_14296);
nor U15180 (N_15180,N_14653,N_14111);
nor U15181 (N_15181,N_14080,N_14940);
and U15182 (N_15182,N_14403,N_14173);
and U15183 (N_15183,N_14076,N_14079);
xor U15184 (N_15184,N_14881,N_14416);
xor U15185 (N_15185,N_14719,N_14315);
or U15186 (N_15186,N_14544,N_14388);
nor U15187 (N_15187,N_14577,N_14478);
nor U15188 (N_15188,N_14049,N_14548);
nand U15189 (N_15189,N_14090,N_14207);
or U15190 (N_15190,N_14369,N_14071);
and U15191 (N_15191,N_14815,N_14725);
xnor U15192 (N_15192,N_14521,N_14051);
nor U15193 (N_15193,N_14498,N_14392);
xor U15194 (N_15194,N_14376,N_14545);
or U15195 (N_15195,N_14540,N_14072);
nor U15196 (N_15196,N_14538,N_14731);
and U15197 (N_15197,N_14954,N_14823);
xnor U15198 (N_15198,N_14261,N_14637);
nand U15199 (N_15199,N_14876,N_14874);
nand U15200 (N_15200,N_14567,N_14086);
xnor U15201 (N_15201,N_14271,N_14063);
and U15202 (N_15202,N_14317,N_14309);
or U15203 (N_15203,N_14656,N_14201);
xnor U15204 (N_15204,N_14182,N_14446);
or U15205 (N_15205,N_14065,N_14702);
and U15206 (N_15206,N_14502,N_14286);
or U15207 (N_15207,N_14570,N_14748);
nor U15208 (N_15208,N_14847,N_14484);
and U15209 (N_15209,N_14346,N_14619);
xnor U15210 (N_15210,N_14890,N_14727);
or U15211 (N_15211,N_14976,N_14325);
or U15212 (N_15212,N_14855,N_14027);
nand U15213 (N_15213,N_14703,N_14120);
nor U15214 (N_15214,N_14998,N_14030);
nand U15215 (N_15215,N_14760,N_14681);
nor U15216 (N_15216,N_14672,N_14016);
nand U15217 (N_15217,N_14574,N_14750);
and U15218 (N_15218,N_14880,N_14889);
xnor U15219 (N_15219,N_14871,N_14638);
or U15220 (N_15220,N_14341,N_14135);
nand U15221 (N_15221,N_14372,N_14985);
nand U15222 (N_15222,N_14878,N_14386);
nand U15223 (N_15223,N_14863,N_14800);
or U15224 (N_15224,N_14539,N_14993);
and U15225 (N_15225,N_14283,N_14204);
nor U15226 (N_15226,N_14496,N_14973);
xnor U15227 (N_15227,N_14220,N_14737);
and U15228 (N_15228,N_14679,N_14227);
or U15229 (N_15229,N_14104,N_14125);
and U15230 (N_15230,N_14024,N_14472);
and U15231 (N_15231,N_14332,N_14311);
or U15232 (N_15232,N_14205,N_14052);
nand U15233 (N_15233,N_14848,N_14948);
or U15234 (N_15234,N_14732,N_14553);
nor U15235 (N_15235,N_14433,N_14959);
xor U15236 (N_15236,N_14156,N_14191);
or U15237 (N_15237,N_14374,N_14657);
nand U15238 (N_15238,N_14537,N_14918);
and U15239 (N_15239,N_14295,N_14139);
and U15240 (N_15240,N_14733,N_14734);
or U15241 (N_15241,N_14989,N_14397);
and U15242 (N_15242,N_14556,N_14331);
xnor U15243 (N_15243,N_14852,N_14008);
and U15244 (N_15244,N_14790,N_14546);
nor U15245 (N_15245,N_14720,N_14953);
and U15246 (N_15246,N_14108,N_14130);
or U15247 (N_15247,N_14671,N_14557);
nand U15248 (N_15248,N_14287,N_14330);
and U15249 (N_15249,N_14124,N_14828);
nor U15250 (N_15250,N_14381,N_14488);
nand U15251 (N_15251,N_14997,N_14777);
and U15252 (N_15252,N_14639,N_14792);
nand U15253 (N_15253,N_14359,N_14620);
and U15254 (N_15254,N_14017,N_14715);
and U15255 (N_15255,N_14711,N_14581);
or U15256 (N_15256,N_14225,N_14529);
nor U15257 (N_15257,N_14535,N_14082);
xor U15258 (N_15258,N_14280,N_14387);
xor U15259 (N_15259,N_14326,N_14314);
xor U15260 (N_15260,N_14602,N_14943);
and U15261 (N_15261,N_14208,N_14755);
nand U15262 (N_15262,N_14312,N_14655);
and U15263 (N_15263,N_14988,N_14666);
xor U15264 (N_15264,N_14078,N_14968);
and U15265 (N_15265,N_14779,N_14701);
and U15266 (N_15266,N_14652,N_14662);
nor U15267 (N_15267,N_14087,N_14588);
or U15268 (N_15268,N_14786,N_14045);
nand U15269 (N_15269,N_14658,N_14050);
and U15270 (N_15270,N_14327,N_14925);
nor U15271 (N_15271,N_14700,N_14738);
and U15272 (N_15272,N_14665,N_14996);
and U15273 (N_15273,N_14040,N_14706);
and U15274 (N_15274,N_14161,N_14412);
nor U15275 (N_15275,N_14321,N_14632);
nor U15276 (N_15276,N_14771,N_14924);
nand U15277 (N_15277,N_14837,N_14670);
nand U15278 (N_15278,N_14827,N_14430);
and U15279 (N_15279,N_14678,N_14363);
xor U15280 (N_15280,N_14481,N_14770);
nand U15281 (N_15281,N_14302,N_14747);
nor U15282 (N_15282,N_14431,N_14782);
nor U15283 (N_15283,N_14979,N_14222);
and U15284 (N_15284,N_14691,N_14503);
or U15285 (N_15285,N_14522,N_14819);
xor U15286 (N_15286,N_14454,N_14799);
xnor U15287 (N_15287,N_14629,N_14490);
nor U15288 (N_15288,N_14457,N_14585);
nor U15289 (N_15289,N_14304,N_14377);
nor U15290 (N_15290,N_14754,N_14004);
or U15291 (N_15291,N_14319,N_14579);
nor U15292 (N_15292,N_14268,N_14097);
nor U15293 (N_15293,N_14262,N_14206);
and U15294 (N_15294,N_14313,N_14449);
or U15295 (N_15295,N_14179,N_14835);
xnor U15296 (N_15296,N_14927,N_14075);
and U15297 (N_15297,N_14801,N_14360);
nor U15298 (N_15298,N_14674,N_14154);
nor U15299 (N_15299,N_14547,N_14845);
nand U15300 (N_15300,N_14010,N_14354);
xor U15301 (N_15301,N_14590,N_14853);
or U15302 (N_15302,N_14983,N_14109);
xnor U15303 (N_15303,N_14896,N_14826);
xnor U15304 (N_15304,N_14021,N_14345);
xnor U15305 (N_15305,N_14811,N_14046);
nor U15306 (N_15306,N_14167,N_14929);
nor U15307 (N_15307,N_14643,N_14428);
nand U15308 (N_15308,N_14680,N_14034);
nor U15309 (N_15309,N_14775,N_14612);
xnor U15310 (N_15310,N_14870,N_14184);
or U15311 (N_15311,N_14361,N_14589);
and U15312 (N_15312,N_14900,N_14098);
nor U15313 (N_15313,N_14170,N_14340);
nor U15314 (N_15314,N_14025,N_14902);
nor U15315 (N_15315,N_14005,N_14243);
or U15316 (N_15316,N_14676,N_14707);
nor U15317 (N_15317,N_14367,N_14456);
nor U15318 (N_15318,N_14907,N_14435);
or U15319 (N_15319,N_14494,N_14509);
nand U15320 (N_15320,N_14651,N_14669);
or U15321 (N_15321,N_14794,N_14947);
or U15322 (N_15322,N_14157,N_14607);
and U15323 (N_15323,N_14292,N_14788);
nand U15324 (N_15324,N_14745,N_14861);
nor U15325 (N_15325,N_14969,N_14282);
and U15326 (N_15326,N_14288,N_14716);
or U15327 (N_15327,N_14887,N_14583);
or U15328 (N_15328,N_14362,N_14165);
xnor U15329 (N_15329,N_14928,N_14813);
nand U15330 (N_15330,N_14178,N_14563);
nor U15331 (N_15331,N_14839,N_14421);
xnor U15332 (N_15332,N_14247,N_14990);
and U15333 (N_15333,N_14270,N_14611);
or U15334 (N_15334,N_14106,N_14631);
xnor U15335 (N_15335,N_14525,N_14562);
nand U15336 (N_15336,N_14647,N_14031);
or U15337 (N_15337,N_14575,N_14904);
xor U15338 (N_15338,N_14408,N_14158);
nand U15339 (N_15339,N_14131,N_14074);
or U15340 (N_15340,N_14284,N_14002);
nor U15341 (N_15341,N_14524,N_14785);
xor U15342 (N_15342,N_14136,N_14169);
xnor U15343 (N_15343,N_14278,N_14445);
xnor U15344 (N_15344,N_14411,N_14501);
or U15345 (N_15345,N_14192,N_14761);
or U15346 (N_15346,N_14648,N_14047);
and U15347 (N_15347,N_14373,N_14466);
nor U15348 (N_15348,N_14622,N_14219);
nand U15349 (N_15349,N_14623,N_14195);
or U15350 (N_15350,N_14414,N_14277);
and U15351 (N_15351,N_14432,N_14740);
nand U15352 (N_15352,N_14649,N_14576);
xnor U15353 (N_15353,N_14824,N_14001);
and U15354 (N_15354,N_14604,N_14564);
and U15355 (N_15355,N_14982,N_14186);
xor U15356 (N_15356,N_14420,N_14265);
nor U15357 (N_15357,N_14704,N_14235);
or U15358 (N_15358,N_14289,N_14447);
nand U15359 (N_15359,N_14269,N_14486);
or U15360 (N_15360,N_14210,N_14485);
nor U15361 (N_15361,N_14816,N_14633);
or U15362 (N_15362,N_14601,N_14423);
or U15363 (N_15363,N_14094,N_14867);
and U15364 (N_15364,N_14351,N_14162);
xor U15365 (N_15365,N_14467,N_14324);
nand U15366 (N_15366,N_14542,N_14977);
and U15367 (N_15367,N_14549,N_14630);
and U15368 (N_15368,N_14029,N_14664);
and U15369 (N_15369,N_14765,N_14650);
and U15370 (N_15370,N_14365,N_14956);
nor U15371 (N_15371,N_14246,N_14118);
nor U15372 (N_15372,N_14739,N_14842);
nor U15373 (N_15373,N_14627,N_14476);
or U15374 (N_15374,N_14914,N_14329);
or U15375 (N_15375,N_14384,N_14149);
nand U15376 (N_15376,N_14708,N_14717);
xnor U15377 (N_15377,N_14555,N_14759);
nand U15378 (N_15378,N_14009,N_14473);
xor U15379 (N_15379,N_14951,N_14565);
nand U15380 (N_15380,N_14688,N_14909);
and U15381 (N_15381,N_14660,N_14306);
and U15382 (N_15382,N_14175,N_14883);
nand U15383 (N_15383,N_14339,N_14300);
and U15384 (N_15384,N_14606,N_14460);
nand U15385 (N_15385,N_14011,N_14944);
nand U15386 (N_15386,N_14723,N_14015);
xnor U15387 (N_15387,N_14226,N_14722);
xnor U15388 (N_15388,N_14151,N_14587);
or U15389 (N_15389,N_14105,N_14942);
nor U15390 (N_15390,N_14100,N_14134);
nor U15391 (N_15391,N_14809,N_14497);
and U15392 (N_15392,N_14519,N_14593);
or U15393 (N_15393,N_14393,N_14366);
xnor U15394 (N_15394,N_14035,N_14380);
or U15395 (N_15395,N_14455,N_14808);
and U15396 (N_15396,N_14967,N_14234);
xnor U15397 (N_15397,N_14253,N_14975);
or U15398 (N_15398,N_14507,N_14077);
or U15399 (N_15399,N_14121,N_14251);
nand U15400 (N_15400,N_14406,N_14571);
and U15401 (N_15401,N_14152,N_14303);
xor U15402 (N_15402,N_14705,N_14908);
xnor U15403 (N_15403,N_14551,N_14014);
xor U15404 (N_15404,N_14070,N_14751);
nor U15405 (N_15405,N_14194,N_14834);
nor U15406 (N_15406,N_14798,N_14783);
and U15407 (N_15407,N_14964,N_14686);
nand U15408 (N_15408,N_14675,N_14089);
or U15409 (N_15409,N_14443,N_14689);
and U15410 (N_15410,N_14769,N_14934);
nand U15411 (N_15411,N_14224,N_14991);
xnor U15412 (N_15412,N_14599,N_14348);
or U15413 (N_15413,N_14886,N_14290);
nor U15414 (N_15414,N_14825,N_14560);
nor U15415 (N_15415,N_14434,N_14541);
nand U15416 (N_15416,N_14596,N_14888);
nand U15417 (N_15417,N_14592,N_14350);
nand U15418 (N_15418,N_14399,N_14214);
or U15419 (N_15419,N_14461,N_14699);
xor U15420 (N_15420,N_14744,N_14591);
nor U15421 (N_15421,N_14198,N_14112);
and U15422 (N_15422,N_14463,N_14242);
and U15423 (N_15423,N_14858,N_14316);
and U15424 (N_15424,N_14101,N_14859);
or U15425 (N_15425,N_14787,N_14458);
or U15426 (N_15426,N_14133,N_14600);
xnor U15427 (N_15427,N_14343,N_14355);
nand U15428 (N_15428,N_14713,N_14756);
and U15429 (N_15429,N_14882,N_14796);
or U15430 (N_15430,N_14994,N_14091);
nor U15431 (N_15431,N_14119,N_14448);
xnor U15432 (N_15432,N_14438,N_14673);
or U15433 (N_15433,N_14984,N_14892);
xor U15434 (N_15434,N_14955,N_14528);
or U15435 (N_15435,N_14810,N_14724);
nand U15436 (N_15436,N_14391,N_14850);
and U15437 (N_15437,N_14211,N_14552);
nor U15438 (N_15438,N_14451,N_14059);
nand U15439 (N_15439,N_14857,N_14418);
xor U15440 (N_15440,N_14419,N_14028);
nor U15441 (N_15441,N_14663,N_14229);
nand U15442 (N_15442,N_14323,N_14986);
or U15443 (N_15443,N_14464,N_14526);
xnor U15444 (N_15444,N_14353,N_14661);
nand U15445 (N_15445,N_14550,N_14872);
and U15446 (N_15446,N_14163,N_14534);
or U15447 (N_15447,N_14095,N_14240);
nor U15448 (N_15448,N_14899,N_14533);
or U15449 (N_15449,N_14305,N_14322);
and U15450 (N_15450,N_14264,N_14935);
xnor U15451 (N_15451,N_14382,N_14931);
and U15452 (N_15452,N_14256,N_14357);
or U15453 (N_15453,N_14504,N_14174);
or U15454 (N_15454,N_14003,N_14912);
xor U15455 (N_15455,N_14239,N_14865);
xnor U15456 (N_15456,N_14860,N_14518);
or U15457 (N_15457,N_14833,N_14053);
nor U15458 (N_15458,N_14805,N_14578);
nand U15459 (N_15459,N_14584,N_14404);
nand U15460 (N_15460,N_14409,N_14032);
or U15461 (N_15461,N_14405,N_14735);
nand U15462 (N_15462,N_14368,N_14299);
or U15463 (N_15463,N_14258,N_14608);
and U15464 (N_15464,N_14530,N_14088);
xnor U15465 (N_15465,N_14187,N_14422);
and U15466 (N_15466,N_14064,N_14752);
or U15467 (N_15467,N_14335,N_14916);
nand U15468 (N_15468,N_14520,N_14729);
nand U15469 (N_15469,N_14697,N_14508);
xor U15470 (N_15470,N_14949,N_14298);
xnor U15471 (N_15471,N_14007,N_14616);
or U15472 (N_15472,N_14952,N_14113);
xnor U15473 (N_15473,N_14500,N_14396);
nor U15474 (N_15474,N_14491,N_14838);
xor U15475 (N_15475,N_14753,N_14129);
xnor U15476 (N_15476,N_14891,N_14897);
nand U15477 (N_15477,N_14036,N_14921);
nor U15478 (N_15478,N_14635,N_14536);
or U15479 (N_15479,N_14474,N_14132);
or U15480 (N_15480,N_14746,N_14058);
nor U15481 (N_15481,N_14142,N_14308);
nand U15482 (N_15482,N_14851,N_14281);
or U15483 (N_15483,N_14413,N_14209);
nand U15484 (N_15484,N_14532,N_14945);
or U15485 (N_15485,N_14066,N_14223);
or U15486 (N_15486,N_14026,N_14022);
or U15487 (N_15487,N_14164,N_14804);
and U15488 (N_15488,N_14276,N_14618);
and U15489 (N_15489,N_14832,N_14866);
or U15490 (N_15490,N_14561,N_14776);
and U15491 (N_15491,N_14667,N_14180);
nand U15492 (N_15492,N_14272,N_14190);
nor U15493 (N_15493,N_14915,N_14068);
nor U15494 (N_15494,N_14402,N_14830);
nand U15495 (N_15495,N_14517,N_14200);
nor U15496 (N_15496,N_14257,N_14605);
and U15497 (N_15497,N_14569,N_14692);
nor U15498 (N_15498,N_14398,N_14477);
nor U15499 (N_15499,N_14250,N_14531);
nand U15500 (N_15500,N_14613,N_14068);
or U15501 (N_15501,N_14678,N_14869);
xor U15502 (N_15502,N_14549,N_14995);
or U15503 (N_15503,N_14102,N_14879);
and U15504 (N_15504,N_14886,N_14059);
nor U15505 (N_15505,N_14525,N_14702);
xor U15506 (N_15506,N_14249,N_14108);
and U15507 (N_15507,N_14605,N_14033);
and U15508 (N_15508,N_14404,N_14291);
or U15509 (N_15509,N_14634,N_14289);
nand U15510 (N_15510,N_14191,N_14736);
nand U15511 (N_15511,N_14011,N_14371);
xnor U15512 (N_15512,N_14079,N_14691);
or U15513 (N_15513,N_14377,N_14968);
nor U15514 (N_15514,N_14497,N_14838);
xor U15515 (N_15515,N_14232,N_14192);
or U15516 (N_15516,N_14993,N_14452);
or U15517 (N_15517,N_14589,N_14578);
or U15518 (N_15518,N_14389,N_14373);
nor U15519 (N_15519,N_14950,N_14659);
nor U15520 (N_15520,N_14643,N_14767);
or U15521 (N_15521,N_14136,N_14157);
or U15522 (N_15522,N_14738,N_14619);
and U15523 (N_15523,N_14503,N_14677);
and U15524 (N_15524,N_14332,N_14670);
xnor U15525 (N_15525,N_14023,N_14900);
xnor U15526 (N_15526,N_14963,N_14341);
xnor U15527 (N_15527,N_14017,N_14273);
xor U15528 (N_15528,N_14772,N_14095);
xnor U15529 (N_15529,N_14523,N_14912);
or U15530 (N_15530,N_14166,N_14516);
xnor U15531 (N_15531,N_14666,N_14640);
xnor U15532 (N_15532,N_14018,N_14347);
nor U15533 (N_15533,N_14374,N_14234);
and U15534 (N_15534,N_14264,N_14967);
nor U15535 (N_15535,N_14480,N_14098);
and U15536 (N_15536,N_14039,N_14774);
nand U15537 (N_15537,N_14432,N_14828);
or U15538 (N_15538,N_14081,N_14749);
or U15539 (N_15539,N_14174,N_14208);
and U15540 (N_15540,N_14745,N_14539);
or U15541 (N_15541,N_14187,N_14080);
or U15542 (N_15542,N_14074,N_14262);
xnor U15543 (N_15543,N_14037,N_14596);
or U15544 (N_15544,N_14811,N_14959);
or U15545 (N_15545,N_14680,N_14619);
xor U15546 (N_15546,N_14499,N_14140);
or U15547 (N_15547,N_14378,N_14464);
or U15548 (N_15548,N_14504,N_14490);
and U15549 (N_15549,N_14059,N_14266);
nor U15550 (N_15550,N_14692,N_14746);
or U15551 (N_15551,N_14299,N_14119);
nor U15552 (N_15552,N_14897,N_14026);
or U15553 (N_15553,N_14730,N_14721);
or U15554 (N_15554,N_14896,N_14592);
xnor U15555 (N_15555,N_14699,N_14626);
nor U15556 (N_15556,N_14108,N_14149);
nand U15557 (N_15557,N_14323,N_14209);
xnor U15558 (N_15558,N_14542,N_14381);
nand U15559 (N_15559,N_14447,N_14281);
nor U15560 (N_15560,N_14687,N_14805);
xnor U15561 (N_15561,N_14257,N_14626);
nor U15562 (N_15562,N_14147,N_14644);
or U15563 (N_15563,N_14393,N_14440);
nor U15564 (N_15564,N_14912,N_14410);
and U15565 (N_15565,N_14191,N_14694);
nand U15566 (N_15566,N_14413,N_14949);
xnor U15567 (N_15567,N_14267,N_14567);
or U15568 (N_15568,N_14142,N_14154);
nand U15569 (N_15569,N_14875,N_14027);
nor U15570 (N_15570,N_14479,N_14854);
xor U15571 (N_15571,N_14324,N_14065);
nand U15572 (N_15572,N_14506,N_14026);
or U15573 (N_15573,N_14434,N_14376);
nand U15574 (N_15574,N_14529,N_14523);
xor U15575 (N_15575,N_14357,N_14290);
or U15576 (N_15576,N_14578,N_14391);
xnor U15577 (N_15577,N_14227,N_14942);
or U15578 (N_15578,N_14417,N_14177);
nor U15579 (N_15579,N_14011,N_14048);
or U15580 (N_15580,N_14063,N_14627);
or U15581 (N_15581,N_14005,N_14290);
nor U15582 (N_15582,N_14565,N_14078);
or U15583 (N_15583,N_14138,N_14262);
and U15584 (N_15584,N_14146,N_14068);
and U15585 (N_15585,N_14694,N_14976);
and U15586 (N_15586,N_14539,N_14576);
and U15587 (N_15587,N_14874,N_14836);
xor U15588 (N_15588,N_14915,N_14301);
xnor U15589 (N_15589,N_14566,N_14780);
nor U15590 (N_15590,N_14733,N_14850);
nand U15591 (N_15591,N_14868,N_14815);
or U15592 (N_15592,N_14955,N_14313);
xnor U15593 (N_15593,N_14196,N_14893);
nor U15594 (N_15594,N_14938,N_14427);
and U15595 (N_15595,N_14111,N_14210);
or U15596 (N_15596,N_14065,N_14189);
nand U15597 (N_15597,N_14689,N_14287);
nand U15598 (N_15598,N_14502,N_14676);
nor U15599 (N_15599,N_14073,N_14271);
nor U15600 (N_15600,N_14037,N_14881);
and U15601 (N_15601,N_14512,N_14217);
and U15602 (N_15602,N_14081,N_14115);
and U15603 (N_15603,N_14178,N_14188);
xnor U15604 (N_15604,N_14509,N_14891);
xor U15605 (N_15605,N_14162,N_14801);
nand U15606 (N_15606,N_14530,N_14393);
nor U15607 (N_15607,N_14892,N_14276);
and U15608 (N_15608,N_14439,N_14771);
or U15609 (N_15609,N_14168,N_14136);
nand U15610 (N_15610,N_14922,N_14272);
and U15611 (N_15611,N_14952,N_14037);
and U15612 (N_15612,N_14454,N_14055);
nor U15613 (N_15613,N_14716,N_14877);
nor U15614 (N_15614,N_14823,N_14769);
nor U15615 (N_15615,N_14292,N_14081);
nand U15616 (N_15616,N_14097,N_14112);
xnor U15617 (N_15617,N_14723,N_14491);
nand U15618 (N_15618,N_14880,N_14170);
nor U15619 (N_15619,N_14301,N_14011);
nand U15620 (N_15620,N_14924,N_14897);
and U15621 (N_15621,N_14812,N_14109);
nand U15622 (N_15622,N_14138,N_14726);
xnor U15623 (N_15623,N_14364,N_14748);
or U15624 (N_15624,N_14855,N_14568);
nand U15625 (N_15625,N_14691,N_14084);
xnor U15626 (N_15626,N_14721,N_14642);
nand U15627 (N_15627,N_14127,N_14550);
or U15628 (N_15628,N_14093,N_14038);
or U15629 (N_15629,N_14569,N_14577);
nand U15630 (N_15630,N_14637,N_14528);
nor U15631 (N_15631,N_14000,N_14684);
xor U15632 (N_15632,N_14424,N_14434);
or U15633 (N_15633,N_14887,N_14791);
nor U15634 (N_15634,N_14745,N_14540);
and U15635 (N_15635,N_14567,N_14989);
nor U15636 (N_15636,N_14528,N_14513);
or U15637 (N_15637,N_14696,N_14570);
nand U15638 (N_15638,N_14773,N_14209);
and U15639 (N_15639,N_14562,N_14430);
and U15640 (N_15640,N_14798,N_14022);
nand U15641 (N_15641,N_14751,N_14060);
xor U15642 (N_15642,N_14884,N_14392);
nor U15643 (N_15643,N_14584,N_14913);
or U15644 (N_15644,N_14578,N_14874);
and U15645 (N_15645,N_14696,N_14439);
xor U15646 (N_15646,N_14429,N_14609);
or U15647 (N_15647,N_14133,N_14518);
nor U15648 (N_15648,N_14983,N_14364);
xor U15649 (N_15649,N_14300,N_14902);
or U15650 (N_15650,N_14367,N_14493);
or U15651 (N_15651,N_14492,N_14252);
nor U15652 (N_15652,N_14916,N_14287);
and U15653 (N_15653,N_14954,N_14718);
nor U15654 (N_15654,N_14880,N_14882);
and U15655 (N_15655,N_14819,N_14429);
or U15656 (N_15656,N_14401,N_14118);
and U15657 (N_15657,N_14493,N_14653);
and U15658 (N_15658,N_14493,N_14902);
nand U15659 (N_15659,N_14745,N_14085);
nand U15660 (N_15660,N_14881,N_14712);
xor U15661 (N_15661,N_14310,N_14188);
and U15662 (N_15662,N_14160,N_14135);
or U15663 (N_15663,N_14809,N_14168);
nor U15664 (N_15664,N_14625,N_14904);
nor U15665 (N_15665,N_14463,N_14481);
nor U15666 (N_15666,N_14398,N_14029);
nor U15667 (N_15667,N_14475,N_14903);
or U15668 (N_15668,N_14510,N_14350);
and U15669 (N_15669,N_14370,N_14558);
and U15670 (N_15670,N_14219,N_14547);
and U15671 (N_15671,N_14848,N_14758);
xor U15672 (N_15672,N_14105,N_14402);
xnor U15673 (N_15673,N_14732,N_14448);
xor U15674 (N_15674,N_14439,N_14955);
and U15675 (N_15675,N_14785,N_14091);
or U15676 (N_15676,N_14249,N_14201);
nand U15677 (N_15677,N_14562,N_14228);
or U15678 (N_15678,N_14056,N_14021);
nand U15679 (N_15679,N_14560,N_14808);
nand U15680 (N_15680,N_14839,N_14658);
xor U15681 (N_15681,N_14431,N_14202);
nand U15682 (N_15682,N_14433,N_14058);
and U15683 (N_15683,N_14075,N_14014);
nand U15684 (N_15684,N_14409,N_14721);
xor U15685 (N_15685,N_14928,N_14800);
nor U15686 (N_15686,N_14521,N_14911);
nand U15687 (N_15687,N_14482,N_14380);
and U15688 (N_15688,N_14938,N_14294);
nand U15689 (N_15689,N_14277,N_14875);
xor U15690 (N_15690,N_14046,N_14688);
and U15691 (N_15691,N_14607,N_14546);
or U15692 (N_15692,N_14368,N_14715);
and U15693 (N_15693,N_14774,N_14138);
nand U15694 (N_15694,N_14475,N_14145);
xnor U15695 (N_15695,N_14313,N_14887);
nand U15696 (N_15696,N_14134,N_14849);
nor U15697 (N_15697,N_14355,N_14741);
nand U15698 (N_15698,N_14482,N_14600);
or U15699 (N_15699,N_14573,N_14077);
nor U15700 (N_15700,N_14407,N_14198);
xnor U15701 (N_15701,N_14392,N_14684);
nand U15702 (N_15702,N_14566,N_14090);
or U15703 (N_15703,N_14805,N_14496);
nor U15704 (N_15704,N_14701,N_14830);
nor U15705 (N_15705,N_14918,N_14155);
or U15706 (N_15706,N_14311,N_14790);
xnor U15707 (N_15707,N_14887,N_14316);
xnor U15708 (N_15708,N_14600,N_14978);
or U15709 (N_15709,N_14796,N_14757);
and U15710 (N_15710,N_14735,N_14681);
nand U15711 (N_15711,N_14076,N_14182);
and U15712 (N_15712,N_14538,N_14572);
nand U15713 (N_15713,N_14670,N_14263);
xnor U15714 (N_15714,N_14617,N_14583);
and U15715 (N_15715,N_14801,N_14559);
or U15716 (N_15716,N_14833,N_14524);
and U15717 (N_15717,N_14525,N_14383);
xnor U15718 (N_15718,N_14580,N_14512);
or U15719 (N_15719,N_14263,N_14378);
nor U15720 (N_15720,N_14876,N_14646);
xor U15721 (N_15721,N_14836,N_14731);
nand U15722 (N_15722,N_14996,N_14483);
nor U15723 (N_15723,N_14048,N_14354);
nand U15724 (N_15724,N_14196,N_14536);
nor U15725 (N_15725,N_14260,N_14239);
nor U15726 (N_15726,N_14040,N_14505);
nand U15727 (N_15727,N_14114,N_14472);
and U15728 (N_15728,N_14224,N_14834);
nand U15729 (N_15729,N_14193,N_14181);
nand U15730 (N_15730,N_14608,N_14145);
nand U15731 (N_15731,N_14741,N_14727);
nor U15732 (N_15732,N_14748,N_14541);
nand U15733 (N_15733,N_14450,N_14134);
nor U15734 (N_15734,N_14910,N_14475);
nand U15735 (N_15735,N_14178,N_14086);
and U15736 (N_15736,N_14287,N_14664);
nor U15737 (N_15737,N_14241,N_14410);
and U15738 (N_15738,N_14678,N_14688);
or U15739 (N_15739,N_14844,N_14109);
xor U15740 (N_15740,N_14218,N_14909);
nor U15741 (N_15741,N_14651,N_14697);
nor U15742 (N_15742,N_14037,N_14669);
nor U15743 (N_15743,N_14519,N_14260);
and U15744 (N_15744,N_14965,N_14151);
nor U15745 (N_15745,N_14873,N_14590);
nor U15746 (N_15746,N_14030,N_14928);
nor U15747 (N_15747,N_14294,N_14799);
xor U15748 (N_15748,N_14434,N_14781);
nand U15749 (N_15749,N_14456,N_14458);
nor U15750 (N_15750,N_14435,N_14737);
and U15751 (N_15751,N_14111,N_14182);
and U15752 (N_15752,N_14304,N_14470);
nor U15753 (N_15753,N_14327,N_14088);
nor U15754 (N_15754,N_14099,N_14058);
or U15755 (N_15755,N_14899,N_14551);
or U15756 (N_15756,N_14261,N_14870);
nand U15757 (N_15757,N_14414,N_14451);
nand U15758 (N_15758,N_14436,N_14472);
nor U15759 (N_15759,N_14509,N_14073);
or U15760 (N_15760,N_14267,N_14602);
and U15761 (N_15761,N_14515,N_14191);
nor U15762 (N_15762,N_14369,N_14365);
or U15763 (N_15763,N_14883,N_14511);
xor U15764 (N_15764,N_14574,N_14641);
xnor U15765 (N_15765,N_14919,N_14257);
nand U15766 (N_15766,N_14266,N_14785);
and U15767 (N_15767,N_14480,N_14786);
nor U15768 (N_15768,N_14708,N_14399);
or U15769 (N_15769,N_14304,N_14013);
nand U15770 (N_15770,N_14504,N_14994);
and U15771 (N_15771,N_14406,N_14171);
and U15772 (N_15772,N_14566,N_14221);
or U15773 (N_15773,N_14986,N_14328);
nor U15774 (N_15774,N_14644,N_14183);
nor U15775 (N_15775,N_14803,N_14799);
and U15776 (N_15776,N_14253,N_14195);
nor U15777 (N_15777,N_14913,N_14709);
nand U15778 (N_15778,N_14580,N_14861);
and U15779 (N_15779,N_14664,N_14508);
or U15780 (N_15780,N_14795,N_14240);
nor U15781 (N_15781,N_14944,N_14821);
nand U15782 (N_15782,N_14102,N_14598);
nor U15783 (N_15783,N_14594,N_14370);
xor U15784 (N_15784,N_14398,N_14515);
and U15785 (N_15785,N_14251,N_14095);
and U15786 (N_15786,N_14201,N_14719);
nor U15787 (N_15787,N_14931,N_14348);
nand U15788 (N_15788,N_14574,N_14188);
nand U15789 (N_15789,N_14788,N_14110);
xor U15790 (N_15790,N_14681,N_14378);
and U15791 (N_15791,N_14102,N_14435);
nor U15792 (N_15792,N_14418,N_14299);
or U15793 (N_15793,N_14284,N_14694);
xnor U15794 (N_15794,N_14128,N_14000);
and U15795 (N_15795,N_14693,N_14932);
and U15796 (N_15796,N_14878,N_14187);
xor U15797 (N_15797,N_14265,N_14088);
nor U15798 (N_15798,N_14485,N_14818);
or U15799 (N_15799,N_14624,N_14070);
xnor U15800 (N_15800,N_14412,N_14430);
or U15801 (N_15801,N_14367,N_14313);
nand U15802 (N_15802,N_14698,N_14155);
or U15803 (N_15803,N_14414,N_14509);
nor U15804 (N_15804,N_14199,N_14858);
nand U15805 (N_15805,N_14611,N_14693);
xor U15806 (N_15806,N_14570,N_14408);
nand U15807 (N_15807,N_14558,N_14569);
nor U15808 (N_15808,N_14105,N_14815);
nand U15809 (N_15809,N_14818,N_14594);
nor U15810 (N_15810,N_14710,N_14518);
nand U15811 (N_15811,N_14998,N_14930);
and U15812 (N_15812,N_14599,N_14301);
xnor U15813 (N_15813,N_14378,N_14237);
nand U15814 (N_15814,N_14421,N_14848);
nand U15815 (N_15815,N_14370,N_14204);
or U15816 (N_15816,N_14428,N_14003);
nor U15817 (N_15817,N_14223,N_14410);
xor U15818 (N_15818,N_14219,N_14446);
and U15819 (N_15819,N_14435,N_14105);
or U15820 (N_15820,N_14645,N_14413);
and U15821 (N_15821,N_14316,N_14441);
nand U15822 (N_15822,N_14379,N_14162);
or U15823 (N_15823,N_14941,N_14056);
and U15824 (N_15824,N_14502,N_14832);
nor U15825 (N_15825,N_14228,N_14755);
xnor U15826 (N_15826,N_14464,N_14919);
nand U15827 (N_15827,N_14981,N_14959);
xor U15828 (N_15828,N_14894,N_14566);
xor U15829 (N_15829,N_14830,N_14994);
nor U15830 (N_15830,N_14978,N_14660);
xnor U15831 (N_15831,N_14736,N_14838);
nor U15832 (N_15832,N_14999,N_14753);
nand U15833 (N_15833,N_14587,N_14174);
and U15834 (N_15834,N_14887,N_14687);
nor U15835 (N_15835,N_14520,N_14715);
and U15836 (N_15836,N_14902,N_14738);
xor U15837 (N_15837,N_14765,N_14526);
nand U15838 (N_15838,N_14370,N_14051);
nand U15839 (N_15839,N_14779,N_14397);
nor U15840 (N_15840,N_14938,N_14637);
or U15841 (N_15841,N_14178,N_14834);
and U15842 (N_15842,N_14727,N_14097);
xnor U15843 (N_15843,N_14916,N_14672);
nor U15844 (N_15844,N_14586,N_14700);
nor U15845 (N_15845,N_14031,N_14916);
or U15846 (N_15846,N_14620,N_14559);
and U15847 (N_15847,N_14990,N_14302);
or U15848 (N_15848,N_14955,N_14126);
and U15849 (N_15849,N_14260,N_14058);
and U15850 (N_15850,N_14878,N_14272);
nand U15851 (N_15851,N_14244,N_14319);
nor U15852 (N_15852,N_14144,N_14399);
nor U15853 (N_15853,N_14587,N_14502);
or U15854 (N_15854,N_14111,N_14194);
nand U15855 (N_15855,N_14493,N_14296);
and U15856 (N_15856,N_14116,N_14325);
xor U15857 (N_15857,N_14919,N_14522);
nor U15858 (N_15858,N_14799,N_14027);
or U15859 (N_15859,N_14108,N_14835);
xnor U15860 (N_15860,N_14087,N_14115);
and U15861 (N_15861,N_14329,N_14599);
or U15862 (N_15862,N_14623,N_14720);
xor U15863 (N_15863,N_14098,N_14599);
xnor U15864 (N_15864,N_14747,N_14298);
nand U15865 (N_15865,N_14913,N_14220);
or U15866 (N_15866,N_14679,N_14716);
or U15867 (N_15867,N_14717,N_14839);
or U15868 (N_15868,N_14638,N_14316);
nor U15869 (N_15869,N_14819,N_14506);
or U15870 (N_15870,N_14590,N_14046);
or U15871 (N_15871,N_14044,N_14356);
or U15872 (N_15872,N_14872,N_14099);
nand U15873 (N_15873,N_14160,N_14951);
nand U15874 (N_15874,N_14234,N_14497);
nand U15875 (N_15875,N_14363,N_14042);
and U15876 (N_15876,N_14664,N_14281);
or U15877 (N_15877,N_14073,N_14175);
nand U15878 (N_15878,N_14022,N_14968);
nor U15879 (N_15879,N_14268,N_14888);
nor U15880 (N_15880,N_14599,N_14562);
xnor U15881 (N_15881,N_14163,N_14216);
nor U15882 (N_15882,N_14437,N_14640);
nor U15883 (N_15883,N_14124,N_14590);
nand U15884 (N_15884,N_14635,N_14035);
or U15885 (N_15885,N_14521,N_14052);
xnor U15886 (N_15886,N_14238,N_14764);
nand U15887 (N_15887,N_14887,N_14694);
nand U15888 (N_15888,N_14240,N_14709);
xnor U15889 (N_15889,N_14121,N_14492);
and U15890 (N_15890,N_14417,N_14961);
or U15891 (N_15891,N_14463,N_14819);
nand U15892 (N_15892,N_14753,N_14216);
xor U15893 (N_15893,N_14082,N_14842);
nor U15894 (N_15894,N_14728,N_14743);
or U15895 (N_15895,N_14850,N_14911);
nor U15896 (N_15896,N_14642,N_14229);
or U15897 (N_15897,N_14744,N_14033);
xnor U15898 (N_15898,N_14845,N_14489);
nor U15899 (N_15899,N_14161,N_14457);
or U15900 (N_15900,N_14988,N_14887);
and U15901 (N_15901,N_14357,N_14397);
or U15902 (N_15902,N_14437,N_14819);
nand U15903 (N_15903,N_14925,N_14159);
and U15904 (N_15904,N_14174,N_14591);
and U15905 (N_15905,N_14273,N_14208);
xnor U15906 (N_15906,N_14845,N_14996);
and U15907 (N_15907,N_14985,N_14651);
and U15908 (N_15908,N_14248,N_14073);
nor U15909 (N_15909,N_14564,N_14473);
nor U15910 (N_15910,N_14708,N_14564);
and U15911 (N_15911,N_14077,N_14255);
nor U15912 (N_15912,N_14526,N_14580);
and U15913 (N_15913,N_14262,N_14388);
or U15914 (N_15914,N_14564,N_14787);
and U15915 (N_15915,N_14813,N_14811);
or U15916 (N_15916,N_14444,N_14190);
nor U15917 (N_15917,N_14298,N_14022);
xnor U15918 (N_15918,N_14218,N_14685);
and U15919 (N_15919,N_14240,N_14369);
or U15920 (N_15920,N_14174,N_14477);
xnor U15921 (N_15921,N_14267,N_14507);
nor U15922 (N_15922,N_14295,N_14779);
or U15923 (N_15923,N_14621,N_14557);
xor U15924 (N_15924,N_14167,N_14881);
or U15925 (N_15925,N_14425,N_14563);
nand U15926 (N_15926,N_14852,N_14105);
or U15927 (N_15927,N_14710,N_14391);
nand U15928 (N_15928,N_14063,N_14953);
xnor U15929 (N_15929,N_14560,N_14259);
nand U15930 (N_15930,N_14133,N_14916);
and U15931 (N_15931,N_14052,N_14395);
xnor U15932 (N_15932,N_14810,N_14901);
xnor U15933 (N_15933,N_14056,N_14451);
or U15934 (N_15934,N_14845,N_14874);
nor U15935 (N_15935,N_14079,N_14186);
or U15936 (N_15936,N_14022,N_14147);
nand U15937 (N_15937,N_14785,N_14743);
and U15938 (N_15938,N_14176,N_14711);
nor U15939 (N_15939,N_14662,N_14464);
nand U15940 (N_15940,N_14381,N_14252);
or U15941 (N_15941,N_14792,N_14224);
and U15942 (N_15942,N_14809,N_14101);
nand U15943 (N_15943,N_14329,N_14140);
or U15944 (N_15944,N_14659,N_14078);
nor U15945 (N_15945,N_14192,N_14336);
nand U15946 (N_15946,N_14768,N_14101);
nor U15947 (N_15947,N_14993,N_14726);
and U15948 (N_15948,N_14774,N_14113);
nand U15949 (N_15949,N_14821,N_14596);
nand U15950 (N_15950,N_14130,N_14403);
nand U15951 (N_15951,N_14437,N_14684);
xnor U15952 (N_15952,N_14505,N_14668);
nand U15953 (N_15953,N_14103,N_14013);
and U15954 (N_15954,N_14724,N_14682);
or U15955 (N_15955,N_14799,N_14147);
nand U15956 (N_15956,N_14144,N_14021);
or U15957 (N_15957,N_14681,N_14481);
nand U15958 (N_15958,N_14782,N_14715);
nand U15959 (N_15959,N_14586,N_14311);
or U15960 (N_15960,N_14475,N_14032);
xor U15961 (N_15961,N_14432,N_14820);
xor U15962 (N_15962,N_14073,N_14898);
nand U15963 (N_15963,N_14963,N_14299);
nor U15964 (N_15964,N_14409,N_14474);
xor U15965 (N_15965,N_14903,N_14202);
and U15966 (N_15966,N_14963,N_14879);
or U15967 (N_15967,N_14882,N_14689);
nor U15968 (N_15968,N_14598,N_14196);
and U15969 (N_15969,N_14908,N_14928);
nor U15970 (N_15970,N_14691,N_14637);
nand U15971 (N_15971,N_14756,N_14053);
nor U15972 (N_15972,N_14204,N_14035);
nand U15973 (N_15973,N_14570,N_14327);
nand U15974 (N_15974,N_14287,N_14532);
or U15975 (N_15975,N_14783,N_14937);
xor U15976 (N_15976,N_14532,N_14384);
nor U15977 (N_15977,N_14433,N_14864);
nor U15978 (N_15978,N_14033,N_14387);
nand U15979 (N_15979,N_14759,N_14812);
nand U15980 (N_15980,N_14990,N_14079);
or U15981 (N_15981,N_14148,N_14536);
and U15982 (N_15982,N_14356,N_14452);
nor U15983 (N_15983,N_14182,N_14853);
nor U15984 (N_15984,N_14333,N_14577);
nand U15985 (N_15985,N_14562,N_14730);
and U15986 (N_15986,N_14152,N_14287);
xnor U15987 (N_15987,N_14469,N_14535);
nor U15988 (N_15988,N_14957,N_14095);
nand U15989 (N_15989,N_14679,N_14979);
xnor U15990 (N_15990,N_14419,N_14062);
nor U15991 (N_15991,N_14894,N_14879);
xnor U15992 (N_15992,N_14785,N_14726);
xnor U15993 (N_15993,N_14586,N_14333);
and U15994 (N_15994,N_14264,N_14266);
xnor U15995 (N_15995,N_14272,N_14348);
xnor U15996 (N_15996,N_14145,N_14177);
nand U15997 (N_15997,N_14241,N_14148);
and U15998 (N_15998,N_14603,N_14811);
nor U15999 (N_15999,N_14889,N_14997);
nor U16000 (N_16000,N_15692,N_15142);
xnor U16001 (N_16001,N_15824,N_15305);
or U16002 (N_16002,N_15197,N_15149);
nand U16003 (N_16003,N_15826,N_15586);
or U16004 (N_16004,N_15465,N_15929);
nand U16005 (N_16005,N_15712,N_15118);
and U16006 (N_16006,N_15440,N_15090);
and U16007 (N_16007,N_15265,N_15287);
nand U16008 (N_16008,N_15718,N_15040);
and U16009 (N_16009,N_15639,N_15626);
or U16010 (N_16010,N_15927,N_15207);
or U16011 (N_16011,N_15426,N_15582);
or U16012 (N_16012,N_15466,N_15263);
nor U16013 (N_16013,N_15389,N_15600);
nand U16014 (N_16014,N_15760,N_15926);
nor U16015 (N_16015,N_15752,N_15993);
nand U16016 (N_16016,N_15917,N_15780);
or U16017 (N_16017,N_15449,N_15219);
xnor U16018 (N_16018,N_15884,N_15827);
and U16019 (N_16019,N_15975,N_15416);
nor U16020 (N_16020,N_15001,N_15778);
nand U16021 (N_16021,N_15279,N_15052);
nand U16022 (N_16022,N_15156,N_15401);
and U16023 (N_16023,N_15837,N_15105);
nand U16024 (N_16024,N_15842,N_15821);
and U16025 (N_16025,N_15218,N_15977);
nand U16026 (N_16026,N_15301,N_15269);
xnor U16027 (N_16027,N_15098,N_15103);
xnor U16028 (N_16028,N_15008,N_15336);
nor U16029 (N_16029,N_15041,N_15633);
nand U16030 (N_16030,N_15726,N_15770);
xnor U16031 (N_16031,N_15550,N_15392);
and U16032 (N_16032,N_15019,N_15189);
or U16033 (N_16033,N_15755,N_15194);
nor U16034 (N_16034,N_15622,N_15454);
xnor U16035 (N_16035,N_15237,N_15832);
or U16036 (N_16036,N_15610,N_15963);
and U16037 (N_16037,N_15529,N_15082);
or U16038 (N_16038,N_15397,N_15025);
and U16039 (N_16039,N_15614,N_15996);
xnor U16040 (N_16040,N_15545,N_15185);
nor U16041 (N_16041,N_15522,N_15300);
or U16042 (N_16042,N_15871,N_15839);
nand U16043 (N_16043,N_15875,N_15234);
and U16044 (N_16044,N_15569,N_15461);
or U16045 (N_16045,N_15646,N_15914);
nor U16046 (N_16046,N_15519,N_15276);
nor U16047 (N_16047,N_15378,N_15972);
and U16048 (N_16048,N_15169,N_15321);
xnor U16049 (N_16049,N_15304,N_15618);
nor U16050 (N_16050,N_15964,N_15326);
nand U16051 (N_16051,N_15874,N_15734);
nor U16052 (N_16052,N_15223,N_15362);
and U16053 (N_16053,N_15377,N_15989);
and U16054 (N_16054,N_15611,N_15604);
or U16055 (N_16055,N_15257,N_15126);
or U16056 (N_16056,N_15111,N_15616);
or U16057 (N_16057,N_15107,N_15475);
xnor U16058 (N_16058,N_15933,N_15596);
and U16059 (N_16059,N_15408,N_15763);
nand U16060 (N_16060,N_15724,N_15779);
nand U16061 (N_16061,N_15016,N_15312);
or U16062 (N_16062,N_15442,N_15801);
or U16063 (N_16063,N_15405,N_15645);
or U16064 (N_16064,N_15201,N_15697);
nor U16065 (N_16065,N_15655,N_15864);
and U16066 (N_16066,N_15608,N_15141);
nor U16067 (N_16067,N_15491,N_15089);
or U16068 (N_16068,N_15367,N_15364);
and U16069 (N_16069,N_15895,N_15383);
nor U16070 (N_16070,N_15418,N_15709);
xnor U16071 (N_16071,N_15000,N_15854);
xor U16072 (N_16072,N_15341,N_15590);
and U16073 (N_16073,N_15115,N_15547);
nor U16074 (N_16074,N_15479,N_15490);
nor U16075 (N_16075,N_15317,N_15469);
nand U16076 (N_16076,N_15177,N_15632);
and U16077 (N_16077,N_15518,N_15096);
xor U16078 (N_16078,N_15244,N_15249);
xor U16079 (N_16079,N_15831,N_15046);
nand U16080 (N_16080,N_15277,N_15638);
nor U16081 (N_16081,N_15686,N_15468);
and U16082 (N_16082,N_15206,N_15805);
nand U16083 (N_16083,N_15662,N_15121);
and U16084 (N_16084,N_15051,N_15698);
nand U16085 (N_16085,N_15495,N_15771);
and U16086 (N_16086,N_15908,N_15371);
nand U16087 (N_16087,N_15815,N_15850);
and U16088 (N_16088,N_15966,N_15564);
or U16089 (N_16089,N_15982,N_15446);
xor U16090 (N_16090,N_15332,N_15938);
nor U16091 (N_16091,N_15236,N_15151);
nor U16092 (N_16092,N_15375,N_15880);
nand U16093 (N_16093,N_15044,N_15535);
or U16094 (N_16094,N_15109,N_15047);
or U16095 (N_16095,N_15765,N_15147);
and U16096 (N_16096,N_15634,N_15039);
and U16097 (N_16097,N_15767,N_15602);
nand U16098 (N_16098,N_15949,N_15330);
and U16099 (N_16099,N_15087,N_15427);
nor U16100 (N_16100,N_15736,N_15737);
and U16101 (N_16101,N_15685,N_15642);
nand U16102 (N_16102,N_15555,N_15102);
and U16103 (N_16103,N_15097,N_15138);
nand U16104 (N_16104,N_15811,N_15203);
nor U16105 (N_16105,N_15443,N_15084);
xnor U16106 (N_16106,N_15879,N_15117);
and U16107 (N_16107,N_15623,N_15882);
or U16108 (N_16108,N_15352,N_15599);
xor U16109 (N_16109,N_15369,N_15159);
nand U16110 (N_16110,N_15387,N_15857);
nand U16111 (N_16111,N_15504,N_15055);
nand U16112 (N_16112,N_15943,N_15015);
nor U16113 (N_16113,N_15132,N_15784);
or U16114 (N_16114,N_15687,N_15013);
and U16115 (N_16115,N_15431,N_15669);
nand U16116 (N_16116,N_15554,N_15009);
and U16117 (N_16117,N_15259,N_15222);
and U16118 (N_16118,N_15987,N_15979);
or U16119 (N_16119,N_15790,N_15937);
nand U16120 (N_16120,N_15834,N_15166);
xnor U16121 (N_16121,N_15588,N_15225);
nand U16122 (N_16122,N_15877,N_15509);
xor U16123 (N_16123,N_15487,N_15829);
xnor U16124 (N_16124,N_15565,N_15192);
nand U16125 (N_16125,N_15088,N_15460);
nor U16126 (N_16126,N_15474,N_15160);
or U16127 (N_16127,N_15548,N_15229);
nand U16128 (N_16128,N_15212,N_15906);
nand U16129 (N_16129,N_15940,N_15756);
nand U16130 (N_16130,N_15394,N_15316);
nor U16131 (N_16131,N_15947,N_15417);
and U16132 (N_16132,N_15061,N_15543);
nor U16133 (N_16133,N_15310,N_15258);
xnor U16134 (N_16134,N_15447,N_15580);
nand U16135 (N_16135,N_15386,N_15080);
or U16136 (N_16136,N_15407,N_15546);
nor U16137 (N_16137,N_15643,N_15761);
and U16138 (N_16138,N_15788,N_15007);
and U16139 (N_16139,N_15808,N_15021);
nor U16140 (N_16140,N_15445,N_15482);
or U16141 (N_16141,N_15925,N_15050);
or U16142 (N_16142,N_15022,N_15794);
or U16143 (N_16143,N_15146,N_15216);
nand U16144 (N_16144,N_15422,N_15356);
nor U16145 (N_16145,N_15250,N_15085);
or U16146 (N_16146,N_15713,N_15343);
nor U16147 (N_16147,N_15211,N_15665);
or U16148 (N_16148,N_15911,N_15744);
nor U16149 (N_16149,N_15594,N_15045);
or U16150 (N_16150,N_15553,N_15335);
or U16151 (N_16151,N_15031,N_15570);
and U16152 (N_16152,N_15601,N_15999);
nor U16153 (N_16153,N_15360,N_15795);
nand U16154 (N_16154,N_15836,N_15253);
nand U16155 (N_16155,N_15372,N_15951);
and U16156 (N_16156,N_15666,N_15847);
xnor U16157 (N_16157,N_15042,N_15799);
nand U16158 (N_16158,N_15533,N_15345);
nand U16159 (N_16159,N_15302,N_15524);
nand U16160 (N_16160,N_15133,N_15284);
or U16161 (N_16161,N_15406,N_15520);
or U16162 (N_16162,N_15581,N_15484);
xnor U16163 (N_16163,N_15749,N_15433);
xor U16164 (N_16164,N_15254,N_15672);
or U16165 (N_16165,N_15036,N_15204);
nor U16166 (N_16166,N_15043,N_15458);
xnor U16167 (N_16167,N_15423,N_15932);
nand U16168 (N_16168,N_15477,N_15521);
or U16169 (N_16169,N_15507,N_15324);
and U16170 (N_16170,N_15057,N_15293);
nand U16171 (N_16171,N_15956,N_15283);
or U16172 (N_16172,N_15694,N_15180);
or U16173 (N_16173,N_15199,N_15514);
nand U16174 (N_16174,N_15591,N_15186);
and U16175 (N_16175,N_15359,N_15278);
or U16176 (N_16176,N_15948,N_15910);
xor U16177 (N_16177,N_15577,N_15656);
xnor U16178 (N_16178,N_15235,N_15231);
nor U16179 (N_16179,N_15074,N_15980);
and U16180 (N_16180,N_15573,N_15391);
nor U16181 (N_16181,N_15171,N_15322);
nor U16182 (N_16182,N_15158,N_15624);
or U16183 (N_16183,N_15717,N_15029);
and U16184 (N_16184,N_15900,N_15523);
or U16185 (N_16185,N_15455,N_15973);
nor U16186 (N_16186,N_15093,N_15497);
xnor U16187 (N_16187,N_15451,N_15885);
or U16188 (N_16188,N_15696,N_15512);
xor U16189 (N_16189,N_15680,N_15769);
nand U16190 (N_16190,N_15167,N_15266);
and U16191 (N_16191,N_15489,N_15721);
and U16192 (N_16192,N_15309,N_15774);
or U16193 (N_16193,N_15628,N_15114);
or U16194 (N_16194,N_15888,N_15851);
and U16195 (N_16195,N_15246,N_15150);
nand U16196 (N_16196,N_15747,N_15153);
nor U16197 (N_16197,N_15384,N_15593);
and U16198 (N_16198,N_15541,N_15403);
and U16199 (N_16199,N_15786,N_15873);
or U16200 (N_16200,N_15483,N_15382);
and U16201 (N_16201,N_15308,N_15318);
nor U16202 (N_16202,N_15240,N_15511);
or U16203 (N_16203,N_15499,N_15969);
and U16204 (N_16204,N_15400,N_15135);
nand U16205 (N_16205,N_15034,N_15746);
nor U16206 (N_16206,N_15571,N_15331);
xnor U16207 (N_16207,N_15463,N_15974);
or U16208 (N_16208,N_15540,N_15781);
nor U16209 (N_16209,N_15075,N_15228);
nor U16210 (N_16210,N_15603,N_15700);
nand U16211 (N_16211,N_15561,N_15239);
nor U16212 (N_16212,N_15673,N_15459);
nand U16213 (N_16213,N_15961,N_15393);
nand U16214 (N_16214,N_15741,N_15732);
nor U16215 (N_16215,N_15373,N_15315);
xor U16216 (N_16216,N_15255,N_15684);
xnor U16217 (N_16217,N_15486,N_15701);
nor U16218 (N_16218,N_15689,N_15967);
or U16219 (N_16219,N_15165,N_15707);
and U16220 (N_16220,N_15131,N_15915);
nand U16221 (N_16221,N_15506,N_15004);
and U16222 (N_16222,N_15453,N_15472);
and U16223 (N_16223,N_15068,N_15347);
xnor U16224 (N_16224,N_15783,N_15889);
and U16225 (N_16225,N_15681,N_15652);
xnor U16226 (N_16226,N_15396,N_15606);
and U16227 (N_16227,N_15714,N_15325);
nor U16228 (N_16228,N_15739,N_15730);
and U16229 (N_16229,N_15187,N_15711);
xnor U16230 (N_16230,N_15992,N_15501);
xor U16231 (N_16231,N_15860,N_15429);
and U16232 (N_16232,N_15728,N_15441);
and U16233 (N_16233,N_15720,N_15764);
xor U16234 (N_16234,N_15539,N_15868);
xnor U16235 (N_16235,N_15527,N_15395);
or U16236 (N_16236,N_15478,N_15448);
nand U16237 (N_16237,N_15748,N_15605);
nand U16238 (N_16238,N_15220,N_15411);
xor U16239 (N_16239,N_15759,N_15476);
and U16240 (N_16240,N_15464,N_15766);
xnor U16241 (N_16241,N_15072,N_15542);
or U16242 (N_16242,N_15462,N_15575);
xor U16243 (N_16243,N_15157,N_15178);
xor U16244 (N_16244,N_15682,N_15430);
and U16245 (N_16245,N_15667,N_15968);
xnor U16246 (N_16246,N_15905,N_15134);
or U16247 (N_16247,N_15835,N_15221);
nor U16248 (N_16248,N_15232,N_15957);
and U16249 (N_16249,N_15731,N_15500);
or U16250 (N_16250,N_15584,N_15496);
and U16251 (N_16251,N_15776,N_15439);
xnor U16252 (N_16252,N_15858,N_15248);
or U16253 (N_16253,N_15168,N_15688);
nor U16254 (N_16254,N_15091,N_15725);
nand U16255 (N_16255,N_15894,N_15777);
nor U16256 (N_16256,N_15334,N_15904);
xor U16257 (N_16257,N_15872,N_15559);
or U16258 (N_16258,N_15358,N_15558);
nand U16259 (N_16259,N_15876,N_15674);
nor U16260 (N_16260,N_15027,N_15179);
or U16261 (N_16261,N_15054,N_15637);
and U16262 (N_16262,N_15648,N_15438);
and U16263 (N_16263,N_15653,N_15313);
nand U16264 (N_16264,N_15399,N_15161);
nor U16265 (N_16265,N_15892,N_15916);
xor U16266 (N_16266,N_15994,N_15838);
nor U16267 (N_16267,N_15307,N_15883);
nor U16268 (N_16268,N_15657,N_15902);
and U16269 (N_16269,N_15921,N_15671);
nand U16270 (N_16270,N_15390,N_15798);
nor U16271 (N_16271,N_15502,N_15076);
and U16272 (N_16272,N_15812,N_15480);
or U16273 (N_16273,N_15067,N_15374);
nand U16274 (N_16274,N_15078,N_15704);
or U16275 (N_16275,N_15370,N_15128);
xor U16276 (N_16276,N_15557,N_15958);
xor U16277 (N_16277,N_15579,N_15410);
nand U16278 (N_16278,N_15970,N_15053);
xnor U16279 (N_16279,N_15243,N_15845);
and U16280 (N_16280,N_15750,N_15702);
and U16281 (N_16281,N_15768,N_15175);
nor U16282 (N_16282,N_15471,N_15260);
or U16283 (N_16283,N_15402,N_15470);
or U16284 (N_16284,N_15789,N_15174);
xnor U16285 (N_16285,N_15722,N_15679);
or U16286 (N_16286,N_15340,N_15421);
nor U16287 (N_16287,N_15213,N_15620);
xnor U16288 (N_16288,N_15856,N_15913);
nor U16289 (N_16289,N_15844,N_15242);
or U16290 (N_16290,N_15154,N_15797);
nand U16291 (N_16291,N_15339,N_15297);
or U16292 (N_16292,N_15552,N_15754);
or U16293 (N_16293,N_15849,N_15807);
or U16294 (N_16294,N_15881,N_15855);
or U16295 (N_16295,N_15960,N_15006);
or U16296 (N_16296,N_15544,N_15986);
xnor U16297 (N_16297,N_15215,N_15162);
nor U16298 (N_16298,N_15152,N_15621);
nand U16299 (N_16299,N_15145,N_15955);
or U16300 (N_16300,N_15077,N_15574);
nor U16301 (N_16301,N_15742,N_15428);
nand U16302 (N_16302,N_15023,N_15791);
xnor U16303 (N_16303,N_15981,N_15531);
xnor U16304 (N_16304,N_15120,N_15272);
nor U16305 (N_16305,N_15144,N_15320);
nand U16306 (N_16306,N_15513,N_15890);
xnor U16307 (N_16307,N_15743,N_15003);
nor U16308 (N_16308,N_15944,N_15976);
nor U16309 (N_16309,N_15945,N_15530);
and U16310 (N_16310,N_15172,N_15083);
nand U16311 (N_16311,N_15058,N_15631);
and U16312 (N_16312,N_15715,N_15899);
xnor U16313 (N_16313,N_15668,N_15063);
nand U16314 (N_16314,N_15492,N_15110);
nand U16315 (N_16315,N_15424,N_15290);
or U16316 (N_16316,N_15990,N_15663);
or U16317 (N_16317,N_15281,N_15256);
nor U16318 (N_16318,N_15456,N_15337);
and U16319 (N_16319,N_15738,N_15912);
xor U16320 (N_16320,N_15901,N_15677);
nand U16321 (N_16321,N_15946,N_15935);
and U16322 (N_16322,N_15164,N_15923);
xor U16323 (N_16323,N_15415,N_15033);
and U16324 (N_16324,N_15139,N_15488);
and U16325 (N_16325,N_15238,N_15723);
nand U16326 (N_16326,N_15866,N_15285);
nor U16327 (N_16327,N_15585,N_15226);
nand U16328 (N_16328,N_15069,N_15971);
or U16329 (N_16329,N_15419,N_15716);
and U16330 (N_16330,N_15810,N_15804);
nor U16331 (N_16331,N_15931,N_15583);
or U16332 (N_16332,N_15525,N_15607);
nand U16333 (N_16333,N_15772,N_15368);
and U16334 (N_16334,N_15988,N_15011);
xor U16335 (N_16335,N_15567,N_15409);
xor U16336 (N_16336,N_15209,N_15435);
nand U16337 (N_16337,N_15205,N_15640);
and U16338 (N_16338,N_15163,N_15745);
nor U16339 (N_16339,N_15630,N_15028);
nand U16340 (N_16340,N_15355,N_15998);
nor U16341 (N_16341,N_15843,N_15846);
and U16342 (N_16342,N_15361,N_15329);
xor U16343 (N_16343,N_15196,N_15129);
xnor U16344 (N_16344,N_15978,N_15349);
xnor U16345 (N_16345,N_15612,N_15896);
xnor U16346 (N_16346,N_15404,N_15985);
nand U16347 (N_16347,N_15597,N_15170);
xnor U16348 (N_16348,N_15298,N_15647);
or U16349 (N_16349,N_15928,N_15233);
or U16350 (N_16350,N_15809,N_15127);
or U16351 (N_16351,N_15173,N_15753);
nand U16352 (N_16352,N_15959,N_15878);
xor U16353 (N_16353,N_15823,N_15002);
nand U16354 (N_16354,N_15820,N_15056);
or U16355 (N_16355,N_15193,N_15282);
and U16356 (N_16356,N_15942,N_15936);
and U16357 (N_16357,N_15920,N_15813);
and U16358 (N_16358,N_15289,N_15534);
or U16359 (N_16359,N_15690,N_15342);
and U16360 (N_16360,N_15636,N_15261);
or U16361 (N_16361,N_15560,N_15859);
or U16362 (N_16362,N_15566,N_15247);
nand U16363 (N_16363,N_15344,N_15155);
nor U16364 (N_16364,N_15800,N_15609);
nand U16365 (N_16365,N_15751,N_15274);
and U16366 (N_16366,N_15997,N_15675);
nand U16367 (N_16367,N_15869,N_15292);
nor U16368 (N_16368,N_15676,N_15841);
nor U16369 (N_16369,N_15327,N_15271);
or U16370 (N_16370,N_15014,N_15862);
nor U16371 (N_16371,N_15840,N_15909);
or U16372 (N_16372,N_15587,N_15357);
or U16373 (N_16373,N_15012,N_15104);
xor U16374 (N_16374,N_15227,N_15048);
nor U16375 (N_16375,N_15100,N_15934);
nand U16376 (N_16376,N_15140,N_15727);
and U16377 (N_16377,N_15020,N_15962);
xor U16378 (N_16378,N_15870,N_15886);
nand U16379 (N_16379,N_15005,N_15062);
or U16380 (N_16380,N_15024,N_15398);
or U16381 (N_16381,N_15264,N_15346);
nor U16382 (N_16382,N_15617,N_15644);
and U16383 (N_16383,N_15113,N_15286);
and U16384 (N_16384,N_15651,N_15549);
nand U16385 (N_16385,N_15683,N_15641);
nor U16386 (N_16386,N_15493,N_15516);
and U16387 (N_16387,N_15625,N_15195);
or U16388 (N_16388,N_15863,N_15528);
or U16389 (N_16389,N_15143,N_15434);
xnor U16390 (N_16390,N_15825,N_15354);
nor U16391 (N_16391,N_15729,N_15314);
and U16392 (N_16392,N_15288,N_15299);
and U16393 (N_16393,N_15853,N_15830);
or U16394 (N_16394,N_15444,N_15619);
and U16395 (N_16395,N_15852,N_15661);
or U16396 (N_16396,N_15572,N_15952);
or U16397 (N_16397,N_15592,N_15119);
and U16398 (N_16398,N_15536,N_15941);
and U16399 (N_16399,N_15245,N_15295);
nor U16400 (N_16400,N_15388,N_15818);
nand U16401 (N_16401,N_15510,N_15338);
nand U16402 (N_16402,N_15066,N_15241);
nor U16403 (N_16403,N_15867,N_15210);
nand U16404 (N_16404,N_15699,N_15414);
and U16405 (N_16405,N_15136,N_15353);
xnor U16406 (N_16406,N_15664,N_15202);
nor U16407 (N_16407,N_15413,N_15613);
nor U16408 (N_16408,N_15635,N_15412);
and U16409 (N_16409,N_15814,N_15079);
and U16410 (N_16410,N_15563,N_15073);
and U16411 (N_16411,N_15538,N_15551);
xnor U16412 (N_16412,N_15030,N_15939);
xnor U16413 (N_16413,N_15311,N_15757);
xor U16414 (N_16414,N_15773,N_15148);
nand U16415 (N_16415,N_15893,N_15190);
nor U16416 (N_16416,N_15268,N_15762);
nor U16417 (N_16417,N_15116,N_15984);
nor U16418 (N_16418,N_15891,N_15740);
and U16419 (N_16419,N_15275,N_15517);
nand U16420 (N_16420,N_15833,N_15775);
nor U16421 (N_16421,N_15010,N_15865);
xor U16422 (N_16422,N_15710,N_15328);
xnor U16423 (N_16423,N_15695,N_15954);
nor U16424 (N_16424,N_15576,N_15191);
and U16425 (N_16425,N_15071,N_15294);
and U16426 (N_16426,N_15562,N_15064);
nor U16427 (N_16427,N_15595,N_15670);
nand U16428 (N_16428,N_15363,N_15306);
and U16429 (N_16429,N_15924,N_15296);
and U16430 (N_16430,N_15659,N_15348);
nand U16431 (N_16431,N_15816,N_15450);
xnor U16432 (N_16432,N_15494,N_15017);
and U16433 (N_16433,N_15568,N_15919);
and U16434 (N_16434,N_15200,N_15705);
nor U16435 (N_16435,N_15660,N_15930);
and U16436 (N_16436,N_15086,N_15991);
nand U16437 (N_16437,N_15983,N_15262);
xor U16438 (N_16438,N_15198,N_15035);
nor U16439 (N_16439,N_15230,N_15099);
nor U16440 (N_16440,N_15124,N_15803);
nand U16441 (N_16441,N_15385,N_15319);
nand U16442 (N_16442,N_15267,N_15782);
nor U16443 (N_16443,N_15649,N_15351);
nor U16444 (N_16444,N_15787,N_15184);
nor U16445 (N_16445,N_15059,N_15183);
nand U16446 (N_16446,N_15995,N_15270);
and U16447 (N_16447,N_15556,N_15578);
xor U16448 (N_16448,N_15526,N_15081);
or U16449 (N_16449,N_15965,N_15379);
nor U16450 (N_16450,N_15708,N_15112);
and U16451 (N_16451,N_15101,N_15252);
xor U16452 (N_16452,N_15208,N_15654);
nor U16453 (N_16453,N_15432,N_15457);
nand U16454 (N_16454,N_15792,N_15922);
xnor U16455 (N_16455,N_15323,N_15503);
or U16456 (N_16456,N_15130,N_15785);
nor U16457 (N_16457,N_15366,N_15381);
nor U16458 (N_16458,N_15303,N_15907);
nor U16459 (N_16459,N_15026,N_15802);
xnor U16460 (N_16460,N_15481,N_15251);
nor U16461 (N_16461,N_15049,N_15094);
nor U16462 (N_16462,N_15018,N_15106);
or U16463 (N_16463,N_15537,N_15532);
and U16464 (N_16464,N_15897,N_15598);
and U16465 (N_16465,N_15380,N_15224);
and U16466 (N_16466,N_15793,N_15365);
xor U16467 (N_16467,N_15070,N_15796);
and U16468 (N_16468,N_15038,N_15065);
xnor U16469 (N_16469,N_15629,N_15032);
and U16470 (N_16470,N_15806,N_15452);
nand U16471 (N_16471,N_15848,N_15650);
and U16472 (N_16472,N_15508,N_15060);
or U16473 (N_16473,N_15627,N_15350);
or U16474 (N_16474,N_15123,N_15898);
nor U16475 (N_16475,N_15515,N_15817);
or U16476 (N_16476,N_15953,N_15473);
or U16477 (N_16477,N_15467,N_15436);
nor U16478 (N_16478,N_15693,N_15095);
nor U16479 (N_16479,N_15333,N_15485);
or U16480 (N_16480,N_15273,N_15658);
nor U16481 (N_16481,N_15376,N_15108);
nor U16482 (N_16482,N_15903,N_15887);
xnor U16483 (N_16483,N_15037,N_15615);
or U16484 (N_16484,N_15589,N_15703);
nand U16485 (N_16485,N_15733,N_15214);
xor U16486 (N_16486,N_15828,N_15498);
and U16487 (N_16487,N_15691,N_15735);
nand U16488 (N_16488,N_15758,N_15182);
and U16489 (N_16489,N_15950,N_15176);
nand U16490 (N_16490,N_15822,N_15819);
and U16491 (N_16491,N_15122,N_15291);
nor U16492 (N_16492,N_15861,N_15505);
nand U16493 (N_16493,N_15719,N_15420);
nor U16494 (N_16494,N_15137,N_15280);
xor U16495 (N_16495,N_15678,N_15092);
or U16496 (N_16496,N_15217,N_15425);
or U16497 (N_16497,N_15437,N_15125);
nand U16498 (N_16498,N_15918,N_15181);
xnor U16499 (N_16499,N_15188,N_15706);
xor U16500 (N_16500,N_15467,N_15716);
nor U16501 (N_16501,N_15142,N_15122);
xor U16502 (N_16502,N_15881,N_15725);
nand U16503 (N_16503,N_15332,N_15579);
and U16504 (N_16504,N_15916,N_15944);
xor U16505 (N_16505,N_15880,N_15106);
xor U16506 (N_16506,N_15433,N_15018);
and U16507 (N_16507,N_15602,N_15069);
nor U16508 (N_16508,N_15550,N_15001);
and U16509 (N_16509,N_15275,N_15681);
xnor U16510 (N_16510,N_15982,N_15242);
or U16511 (N_16511,N_15909,N_15815);
nor U16512 (N_16512,N_15850,N_15346);
nand U16513 (N_16513,N_15861,N_15338);
nor U16514 (N_16514,N_15635,N_15216);
and U16515 (N_16515,N_15801,N_15259);
xor U16516 (N_16516,N_15515,N_15840);
and U16517 (N_16517,N_15809,N_15600);
xnor U16518 (N_16518,N_15525,N_15830);
and U16519 (N_16519,N_15077,N_15393);
nor U16520 (N_16520,N_15401,N_15818);
nor U16521 (N_16521,N_15886,N_15792);
nand U16522 (N_16522,N_15639,N_15942);
or U16523 (N_16523,N_15111,N_15862);
or U16524 (N_16524,N_15048,N_15680);
and U16525 (N_16525,N_15323,N_15406);
nor U16526 (N_16526,N_15072,N_15299);
xnor U16527 (N_16527,N_15392,N_15586);
nand U16528 (N_16528,N_15650,N_15756);
nand U16529 (N_16529,N_15811,N_15415);
xnor U16530 (N_16530,N_15524,N_15098);
and U16531 (N_16531,N_15161,N_15723);
nand U16532 (N_16532,N_15733,N_15333);
nor U16533 (N_16533,N_15799,N_15133);
nor U16534 (N_16534,N_15478,N_15041);
nand U16535 (N_16535,N_15698,N_15882);
xnor U16536 (N_16536,N_15644,N_15037);
and U16537 (N_16537,N_15261,N_15643);
and U16538 (N_16538,N_15418,N_15517);
or U16539 (N_16539,N_15672,N_15692);
nor U16540 (N_16540,N_15579,N_15244);
or U16541 (N_16541,N_15528,N_15891);
nor U16542 (N_16542,N_15980,N_15259);
nor U16543 (N_16543,N_15289,N_15187);
xnor U16544 (N_16544,N_15275,N_15818);
xor U16545 (N_16545,N_15636,N_15040);
nand U16546 (N_16546,N_15909,N_15108);
xnor U16547 (N_16547,N_15280,N_15202);
nand U16548 (N_16548,N_15538,N_15360);
or U16549 (N_16549,N_15153,N_15699);
nand U16550 (N_16550,N_15049,N_15423);
nand U16551 (N_16551,N_15739,N_15320);
xnor U16552 (N_16552,N_15174,N_15032);
and U16553 (N_16553,N_15768,N_15340);
nor U16554 (N_16554,N_15990,N_15411);
nor U16555 (N_16555,N_15253,N_15311);
or U16556 (N_16556,N_15889,N_15391);
nor U16557 (N_16557,N_15827,N_15002);
or U16558 (N_16558,N_15259,N_15036);
and U16559 (N_16559,N_15300,N_15544);
or U16560 (N_16560,N_15600,N_15301);
nand U16561 (N_16561,N_15364,N_15705);
nand U16562 (N_16562,N_15720,N_15749);
xor U16563 (N_16563,N_15735,N_15345);
nor U16564 (N_16564,N_15159,N_15174);
and U16565 (N_16565,N_15522,N_15846);
or U16566 (N_16566,N_15564,N_15178);
xor U16567 (N_16567,N_15830,N_15749);
and U16568 (N_16568,N_15079,N_15406);
nand U16569 (N_16569,N_15654,N_15375);
nor U16570 (N_16570,N_15783,N_15194);
or U16571 (N_16571,N_15135,N_15202);
xnor U16572 (N_16572,N_15911,N_15103);
or U16573 (N_16573,N_15087,N_15985);
nand U16574 (N_16574,N_15806,N_15761);
xnor U16575 (N_16575,N_15443,N_15117);
nand U16576 (N_16576,N_15939,N_15922);
nor U16577 (N_16577,N_15819,N_15329);
and U16578 (N_16578,N_15728,N_15724);
xor U16579 (N_16579,N_15840,N_15128);
xnor U16580 (N_16580,N_15364,N_15281);
and U16581 (N_16581,N_15641,N_15061);
and U16582 (N_16582,N_15196,N_15627);
or U16583 (N_16583,N_15943,N_15750);
xor U16584 (N_16584,N_15702,N_15600);
nand U16585 (N_16585,N_15331,N_15289);
nor U16586 (N_16586,N_15460,N_15092);
xnor U16587 (N_16587,N_15034,N_15227);
or U16588 (N_16588,N_15440,N_15909);
and U16589 (N_16589,N_15117,N_15778);
and U16590 (N_16590,N_15455,N_15294);
and U16591 (N_16591,N_15173,N_15727);
nand U16592 (N_16592,N_15049,N_15296);
nand U16593 (N_16593,N_15653,N_15009);
and U16594 (N_16594,N_15205,N_15896);
xnor U16595 (N_16595,N_15135,N_15684);
nor U16596 (N_16596,N_15771,N_15910);
or U16597 (N_16597,N_15377,N_15225);
nand U16598 (N_16598,N_15764,N_15481);
xnor U16599 (N_16599,N_15066,N_15283);
and U16600 (N_16600,N_15103,N_15327);
and U16601 (N_16601,N_15727,N_15541);
nand U16602 (N_16602,N_15256,N_15247);
xnor U16603 (N_16603,N_15376,N_15823);
and U16604 (N_16604,N_15267,N_15126);
or U16605 (N_16605,N_15969,N_15201);
and U16606 (N_16606,N_15269,N_15733);
nor U16607 (N_16607,N_15733,N_15629);
or U16608 (N_16608,N_15881,N_15433);
xor U16609 (N_16609,N_15304,N_15953);
and U16610 (N_16610,N_15072,N_15550);
and U16611 (N_16611,N_15775,N_15056);
and U16612 (N_16612,N_15372,N_15629);
xnor U16613 (N_16613,N_15417,N_15513);
or U16614 (N_16614,N_15388,N_15110);
xnor U16615 (N_16615,N_15617,N_15408);
nand U16616 (N_16616,N_15419,N_15880);
nand U16617 (N_16617,N_15539,N_15657);
or U16618 (N_16618,N_15197,N_15612);
and U16619 (N_16619,N_15462,N_15288);
xnor U16620 (N_16620,N_15473,N_15780);
xor U16621 (N_16621,N_15828,N_15638);
nor U16622 (N_16622,N_15289,N_15406);
xnor U16623 (N_16623,N_15137,N_15265);
xor U16624 (N_16624,N_15704,N_15490);
and U16625 (N_16625,N_15620,N_15438);
xnor U16626 (N_16626,N_15164,N_15666);
nand U16627 (N_16627,N_15419,N_15669);
and U16628 (N_16628,N_15020,N_15400);
or U16629 (N_16629,N_15433,N_15172);
or U16630 (N_16630,N_15100,N_15083);
or U16631 (N_16631,N_15983,N_15738);
and U16632 (N_16632,N_15238,N_15573);
xor U16633 (N_16633,N_15122,N_15738);
nor U16634 (N_16634,N_15368,N_15885);
or U16635 (N_16635,N_15414,N_15627);
and U16636 (N_16636,N_15479,N_15656);
nand U16637 (N_16637,N_15722,N_15409);
nor U16638 (N_16638,N_15055,N_15270);
or U16639 (N_16639,N_15317,N_15494);
nand U16640 (N_16640,N_15909,N_15532);
and U16641 (N_16641,N_15014,N_15487);
xor U16642 (N_16642,N_15354,N_15785);
and U16643 (N_16643,N_15076,N_15388);
nand U16644 (N_16644,N_15825,N_15975);
nor U16645 (N_16645,N_15797,N_15564);
nor U16646 (N_16646,N_15796,N_15109);
and U16647 (N_16647,N_15034,N_15039);
nand U16648 (N_16648,N_15670,N_15520);
and U16649 (N_16649,N_15342,N_15562);
nor U16650 (N_16650,N_15187,N_15069);
xor U16651 (N_16651,N_15305,N_15437);
nand U16652 (N_16652,N_15480,N_15982);
nand U16653 (N_16653,N_15487,N_15229);
or U16654 (N_16654,N_15832,N_15887);
xor U16655 (N_16655,N_15036,N_15387);
nor U16656 (N_16656,N_15178,N_15545);
or U16657 (N_16657,N_15623,N_15540);
or U16658 (N_16658,N_15159,N_15545);
or U16659 (N_16659,N_15886,N_15131);
and U16660 (N_16660,N_15584,N_15544);
nor U16661 (N_16661,N_15928,N_15865);
xnor U16662 (N_16662,N_15756,N_15501);
xnor U16663 (N_16663,N_15944,N_15206);
nor U16664 (N_16664,N_15059,N_15877);
or U16665 (N_16665,N_15015,N_15166);
xor U16666 (N_16666,N_15626,N_15776);
and U16667 (N_16667,N_15257,N_15265);
xnor U16668 (N_16668,N_15184,N_15243);
nand U16669 (N_16669,N_15830,N_15297);
or U16670 (N_16670,N_15188,N_15146);
or U16671 (N_16671,N_15124,N_15333);
xnor U16672 (N_16672,N_15102,N_15044);
nand U16673 (N_16673,N_15742,N_15006);
nand U16674 (N_16674,N_15762,N_15538);
and U16675 (N_16675,N_15255,N_15522);
and U16676 (N_16676,N_15480,N_15648);
and U16677 (N_16677,N_15652,N_15651);
nand U16678 (N_16678,N_15711,N_15300);
and U16679 (N_16679,N_15792,N_15131);
xor U16680 (N_16680,N_15596,N_15022);
and U16681 (N_16681,N_15566,N_15545);
nor U16682 (N_16682,N_15699,N_15606);
and U16683 (N_16683,N_15958,N_15677);
nand U16684 (N_16684,N_15389,N_15575);
nand U16685 (N_16685,N_15117,N_15212);
xnor U16686 (N_16686,N_15903,N_15608);
and U16687 (N_16687,N_15872,N_15181);
nand U16688 (N_16688,N_15830,N_15461);
nand U16689 (N_16689,N_15076,N_15505);
or U16690 (N_16690,N_15008,N_15875);
nor U16691 (N_16691,N_15837,N_15614);
or U16692 (N_16692,N_15162,N_15877);
and U16693 (N_16693,N_15088,N_15731);
nand U16694 (N_16694,N_15954,N_15161);
and U16695 (N_16695,N_15163,N_15447);
and U16696 (N_16696,N_15985,N_15480);
and U16697 (N_16697,N_15170,N_15646);
or U16698 (N_16698,N_15308,N_15742);
or U16699 (N_16699,N_15392,N_15173);
nand U16700 (N_16700,N_15705,N_15140);
nor U16701 (N_16701,N_15379,N_15307);
and U16702 (N_16702,N_15319,N_15369);
xnor U16703 (N_16703,N_15038,N_15355);
nor U16704 (N_16704,N_15720,N_15965);
and U16705 (N_16705,N_15525,N_15445);
or U16706 (N_16706,N_15845,N_15247);
nand U16707 (N_16707,N_15909,N_15082);
or U16708 (N_16708,N_15550,N_15350);
nor U16709 (N_16709,N_15655,N_15720);
xnor U16710 (N_16710,N_15681,N_15839);
or U16711 (N_16711,N_15722,N_15673);
nand U16712 (N_16712,N_15732,N_15245);
nor U16713 (N_16713,N_15270,N_15567);
xnor U16714 (N_16714,N_15986,N_15566);
nand U16715 (N_16715,N_15448,N_15291);
and U16716 (N_16716,N_15575,N_15829);
or U16717 (N_16717,N_15856,N_15971);
xor U16718 (N_16718,N_15449,N_15428);
nand U16719 (N_16719,N_15318,N_15822);
nor U16720 (N_16720,N_15931,N_15539);
nor U16721 (N_16721,N_15570,N_15124);
or U16722 (N_16722,N_15469,N_15164);
or U16723 (N_16723,N_15915,N_15657);
xnor U16724 (N_16724,N_15683,N_15105);
nor U16725 (N_16725,N_15508,N_15325);
nand U16726 (N_16726,N_15444,N_15886);
nand U16727 (N_16727,N_15076,N_15765);
and U16728 (N_16728,N_15848,N_15249);
or U16729 (N_16729,N_15207,N_15998);
nand U16730 (N_16730,N_15855,N_15023);
nand U16731 (N_16731,N_15584,N_15083);
nand U16732 (N_16732,N_15625,N_15692);
xnor U16733 (N_16733,N_15792,N_15742);
or U16734 (N_16734,N_15388,N_15300);
xor U16735 (N_16735,N_15788,N_15490);
nor U16736 (N_16736,N_15564,N_15217);
xnor U16737 (N_16737,N_15099,N_15819);
nand U16738 (N_16738,N_15731,N_15937);
nand U16739 (N_16739,N_15036,N_15533);
or U16740 (N_16740,N_15106,N_15008);
nand U16741 (N_16741,N_15521,N_15998);
and U16742 (N_16742,N_15242,N_15814);
nor U16743 (N_16743,N_15698,N_15015);
and U16744 (N_16744,N_15773,N_15550);
or U16745 (N_16745,N_15480,N_15727);
and U16746 (N_16746,N_15925,N_15628);
nand U16747 (N_16747,N_15449,N_15274);
xnor U16748 (N_16748,N_15100,N_15721);
nand U16749 (N_16749,N_15241,N_15176);
and U16750 (N_16750,N_15298,N_15560);
xnor U16751 (N_16751,N_15773,N_15232);
nand U16752 (N_16752,N_15875,N_15533);
or U16753 (N_16753,N_15592,N_15191);
xor U16754 (N_16754,N_15519,N_15873);
nand U16755 (N_16755,N_15971,N_15733);
nand U16756 (N_16756,N_15805,N_15719);
xnor U16757 (N_16757,N_15078,N_15246);
nand U16758 (N_16758,N_15353,N_15289);
and U16759 (N_16759,N_15613,N_15068);
xor U16760 (N_16760,N_15623,N_15121);
xor U16761 (N_16761,N_15494,N_15955);
nor U16762 (N_16762,N_15481,N_15336);
nand U16763 (N_16763,N_15376,N_15739);
nand U16764 (N_16764,N_15238,N_15684);
xnor U16765 (N_16765,N_15521,N_15924);
and U16766 (N_16766,N_15860,N_15287);
xnor U16767 (N_16767,N_15303,N_15694);
or U16768 (N_16768,N_15685,N_15564);
nor U16769 (N_16769,N_15416,N_15919);
and U16770 (N_16770,N_15120,N_15689);
and U16771 (N_16771,N_15569,N_15372);
nor U16772 (N_16772,N_15503,N_15622);
xnor U16773 (N_16773,N_15521,N_15440);
or U16774 (N_16774,N_15642,N_15573);
xnor U16775 (N_16775,N_15665,N_15467);
and U16776 (N_16776,N_15873,N_15234);
or U16777 (N_16777,N_15145,N_15422);
or U16778 (N_16778,N_15338,N_15526);
nand U16779 (N_16779,N_15701,N_15926);
or U16780 (N_16780,N_15510,N_15284);
and U16781 (N_16781,N_15915,N_15351);
nand U16782 (N_16782,N_15971,N_15497);
or U16783 (N_16783,N_15413,N_15155);
nand U16784 (N_16784,N_15841,N_15498);
and U16785 (N_16785,N_15324,N_15538);
xnor U16786 (N_16786,N_15083,N_15317);
nor U16787 (N_16787,N_15665,N_15216);
xor U16788 (N_16788,N_15758,N_15224);
nand U16789 (N_16789,N_15015,N_15726);
nor U16790 (N_16790,N_15237,N_15709);
xnor U16791 (N_16791,N_15847,N_15612);
and U16792 (N_16792,N_15896,N_15370);
xnor U16793 (N_16793,N_15138,N_15287);
nand U16794 (N_16794,N_15160,N_15480);
nor U16795 (N_16795,N_15186,N_15959);
or U16796 (N_16796,N_15180,N_15296);
xnor U16797 (N_16797,N_15458,N_15854);
and U16798 (N_16798,N_15782,N_15018);
nor U16799 (N_16799,N_15891,N_15244);
nor U16800 (N_16800,N_15344,N_15244);
or U16801 (N_16801,N_15562,N_15203);
and U16802 (N_16802,N_15209,N_15155);
nor U16803 (N_16803,N_15085,N_15980);
nand U16804 (N_16804,N_15517,N_15087);
nand U16805 (N_16805,N_15013,N_15094);
and U16806 (N_16806,N_15375,N_15902);
and U16807 (N_16807,N_15476,N_15730);
or U16808 (N_16808,N_15663,N_15013);
xnor U16809 (N_16809,N_15650,N_15598);
or U16810 (N_16810,N_15386,N_15090);
nand U16811 (N_16811,N_15818,N_15506);
or U16812 (N_16812,N_15436,N_15710);
or U16813 (N_16813,N_15749,N_15014);
and U16814 (N_16814,N_15018,N_15673);
and U16815 (N_16815,N_15021,N_15018);
or U16816 (N_16816,N_15599,N_15140);
or U16817 (N_16817,N_15667,N_15741);
nor U16818 (N_16818,N_15261,N_15064);
or U16819 (N_16819,N_15125,N_15734);
nand U16820 (N_16820,N_15095,N_15727);
or U16821 (N_16821,N_15502,N_15967);
or U16822 (N_16822,N_15696,N_15170);
nand U16823 (N_16823,N_15491,N_15099);
and U16824 (N_16824,N_15212,N_15655);
and U16825 (N_16825,N_15685,N_15321);
xnor U16826 (N_16826,N_15544,N_15239);
xor U16827 (N_16827,N_15217,N_15369);
nor U16828 (N_16828,N_15323,N_15728);
xnor U16829 (N_16829,N_15713,N_15833);
or U16830 (N_16830,N_15980,N_15881);
or U16831 (N_16831,N_15286,N_15214);
nor U16832 (N_16832,N_15681,N_15762);
nor U16833 (N_16833,N_15434,N_15773);
or U16834 (N_16834,N_15566,N_15073);
nor U16835 (N_16835,N_15035,N_15465);
nand U16836 (N_16836,N_15823,N_15790);
nor U16837 (N_16837,N_15202,N_15357);
and U16838 (N_16838,N_15500,N_15868);
xor U16839 (N_16839,N_15433,N_15904);
nor U16840 (N_16840,N_15968,N_15013);
nand U16841 (N_16841,N_15426,N_15596);
nand U16842 (N_16842,N_15139,N_15383);
and U16843 (N_16843,N_15341,N_15395);
nand U16844 (N_16844,N_15343,N_15214);
and U16845 (N_16845,N_15928,N_15746);
xnor U16846 (N_16846,N_15335,N_15263);
and U16847 (N_16847,N_15401,N_15281);
xor U16848 (N_16848,N_15057,N_15520);
and U16849 (N_16849,N_15732,N_15044);
nor U16850 (N_16850,N_15722,N_15856);
nand U16851 (N_16851,N_15224,N_15617);
and U16852 (N_16852,N_15863,N_15556);
nand U16853 (N_16853,N_15616,N_15028);
and U16854 (N_16854,N_15508,N_15951);
nor U16855 (N_16855,N_15136,N_15345);
or U16856 (N_16856,N_15890,N_15538);
nor U16857 (N_16857,N_15747,N_15469);
or U16858 (N_16858,N_15671,N_15399);
xor U16859 (N_16859,N_15698,N_15281);
nor U16860 (N_16860,N_15152,N_15562);
xor U16861 (N_16861,N_15145,N_15751);
or U16862 (N_16862,N_15249,N_15100);
nand U16863 (N_16863,N_15117,N_15354);
and U16864 (N_16864,N_15931,N_15733);
or U16865 (N_16865,N_15165,N_15532);
nor U16866 (N_16866,N_15666,N_15090);
or U16867 (N_16867,N_15026,N_15976);
nor U16868 (N_16868,N_15193,N_15856);
or U16869 (N_16869,N_15273,N_15794);
xor U16870 (N_16870,N_15462,N_15092);
and U16871 (N_16871,N_15171,N_15509);
and U16872 (N_16872,N_15168,N_15884);
and U16873 (N_16873,N_15915,N_15790);
and U16874 (N_16874,N_15814,N_15843);
xor U16875 (N_16875,N_15474,N_15103);
xnor U16876 (N_16876,N_15580,N_15648);
xnor U16877 (N_16877,N_15433,N_15772);
xnor U16878 (N_16878,N_15101,N_15939);
or U16879 (N_16879,N_15461,N_15548);
xnor U16880 (N_16880,N_15240,N_15018);
or U16881 (N_16881,N_15597,N_15355);
nor U16882 (N_16882,N_15881,N_15565);
or U16883 (N_16883,N_15180,N_15746);
xnor U16884 (N_16884,N_15710,N_15039);
nor U16885 (N_16885,N_15760,N_15274);
or U16886 (N_16886,N_15780,N_15027);
and U16887 (N_16887,N_15625,N_15082);
nor U16888 (N_16888,N_15214,N_15013);
nor U16889 (N_16889,N_15604,N_15007);
xor U16890 (N_16890,N_15991,N_15217);
nor U16891 (N_16891,N_15838,N_15549);
nor U16892 (N_16892,N_15996,N_15401);
xor U16893 (N_16893,N_15052,N_15111);
xnor U16894 (N_16894,N_15994,N_15507);
and U16895 (N_16895,N_15922,N_15765);
or U16896 (N_16896,N_15890,N_15015);
nand U16897 (N_16897,N_15304,N_15737);
and U16898 (N_16898,N_15053,N_15743);
nor U16899 (N_16899,N_15801,N_15325);
xor U16900 (N_16900,N_15058,N_15033);
nand U16901 (N_16901,N_15782,N_15774);
xnor U16902 (N_16902,N_15539,N_15823);
or U16903 (N_16903,N_15879,N_15781);
nor U16904 (N_16904,N_15913,N_15165);
nand U16905 (N_16905,N_15831,N_15658);
or U16906 (N_16906,N_15721,N_15108);
nand U16907 (N_16907,N_15939,N_15274);
xor U16908 (N_16908,N_15824,N_15907);
nand U16909 (N_16909,N_15415,N_15797);
and U16910 (N_16910,N_15834,N_15029);
nor U16911 (N_16911,N_15021,N_15672);
nor U16912 (N_16912,N_15524,N_15067);
nor U16913 (N_16913,N_15000,N_15490);
or U16914 (N_16914,N_15476,N_15167);
nor U16915 (N_16915,N_15286,N_15174);
nand U16916 (N_16916,N_15555,N_15442);
or U16917 (N_16917,N_15033,N_15506);
or U16918 (N_16918,N_15634,N_15247);
nor U16919 (N_16919,N_15570,N_15709);
or U16920 (N_16920,N_15246,N_15297);
nor U16921 (N_16921,N_15221,N_15279);
nor U16922 (N_16922,N_15351,N_15941);
and U16923 (N_16923,N_15330,N_15944);
xnor U16924 (N_16924,N_15284,N_15458);
nand U16925 (N_16925,N_15655,N_15067);
and U16926 (N_16926,N_15045,N_15439);
and U16927 (N_16927,N_15229,N_15998);
nand U16928 (N_16928,N_15798,N_15235);
xor U16929 (N_16929,N_15521,N_15603);
nand U16930 (N_16930,N_15308,N_15003);
or U16931 (N_16931,N_15059,N_15815);
or U16932 (N_16932,N_15290,N_15796);
nand U16933 (N_16933,N_15537,N_15495);
or U16934 (N_16934,N_15622,N_15563);
or U16935 (N_16935,N_15395,N_15834);
nand U16936 (N_16936,N_15499,N_15142);
nand U16937 (N_16937,N_15668,N_15671);
nor U16938 (N_16938,N_15284,N_15978);
xor U16939 (N_16939,N_15055,N_15487);
nor U16940 (N_16940,N_15842,N_15575);
and U16941 (N_16941,N_15317,N_15004);
xor U16942 (N_16942,N_15467,N_15262);
xor U16943 (N_16943,N_15166,N_15704);
nand U16944 (N_16944,N_15149,N_15250);
and U16945 (N_16945,N_15475,N_15881);
xnor U16946 (N_16946,N_15602,N_15423);
xnor U16947 (N_16947,N_15600,N_15123);
or U16948 (N_16948,N_15103,N_15219);
nand U16949 (N_16949,N_15897,N_15010);
nand U16950 (N_16950,N_15207,N_15544);
xnor U16951 (N_16951,N_15576,N_15030);
nand U16952 (N_16952,N_15781,N_15021);
nand U16953 (N_16953,N_15996,N_15865);
nand U16954 (N_16954,N_15090,N_15162);
nor U16955 (N_16955,N_15341,N_15122);
nand U16956 (N_16956,N_15065,N_15432);
xnor U16957 (N_16957,N_15643,N_15578);
nor U16958 (N_16958,N_15068,N_15861);
and U16959 (N_16959,N_15524,N_15279);
xor U16960 (N_16960,N_15999,N_15891);
or U16961 (N_16961,N_15632,N_15352);
nand U16962 (N_16962,N_15812,N_15864);
nor U16963 (N_16963,N_15964,N_15648);
and U16964 (N_16964,N_15195,N_15895);
nand U16965 (N_16965,N_15904,N_15579);
nand U16966 (N_16966,N_15401,N_15710);
nand U16967 (N_16967,N_15880,N_15617);
xnor U16968 (N_16968,N_15807,N_15468);
xor U16969 (N_16969,N_15819,N_15416);
or U16970 (N_16970,N_15031,N_15127);
or U16971 (N_16971,N_15801,N_15148);
and U16972 (N_16972,N_15171,N_15726);
nand U16973 (N_16973,N_15289,N_15015);
and U16974 (N_16974,N_15843,N_15956);
and U16975 (N_16975,N_15103,N_15136);
and U16976 (N_16976,N_15051,N_15221);
nand U16977 (N_16977,N_15157,N_15118);
nand U16978 (N_16978,N_15688,N_15199);
xor U16979 (N_16979,N_15537,N_15728);
and U16980 (N_16980,N_15251,N_15448);
nand U16981 (N_16981,N_15752,N_15393);
nand U16982 (N_16982,N_15788,N_15977);
nand U16983 (N_16983,N_15375,N_15775);
nand U16984 (N_16984,N_15220,N_15951);
nor U16985 (N_16985,N_15496,N_15497);
xnor U16986 (N_16986,N_15615,N_15862);
nand U16987 (N_16987,N_15546,N_15779);
xor U16988 (N_16988,N_15084,N_15273);
nand U16989 (N_16989,N_15809,N_15484);
xnor U16990 (N_16990,N_15577,N_15211);
nand U16991 (N_16991,N_15155,N_15702);
and U16992 (N_16992,N_15156,N_15039);
xor U16993 (N_16993,N_15568,N_15063);
or U16994 (N_16994,N_15156,N_15403);
nand U16995 (N_16995,N_15818,N_15094);
nand U16996 (N_16996,N_15473,N_15116);
or U16997 (N_16997,N_15261,N_15364);
xor U16998 (N_16998,N_15617,N_15194);
xnor U16999 (N_16999,N_15955,N_15223);
nand U17000 (N_17000,N_16359,N_16596);
nand U17001 (N_17001,N_16431,N_16999);
nor U17002 (N_17002,N_16973,N_16003);
and U17003 (N_17003,N_16201,N_16702);
nand U17004 (N_17004,N_16471,N_16270);
nor U17005 (N_17005,N_16054,N_16375);
nand U17006 (N_17006,N_16949,N_16229);
nor U17007 (N_17007,N_16879,N_16724);
nand U17008 (N_17008,N_16539,N_16391);
nor U17009 (N_17009,N_16437,N_16110);
nor U17010 (N_17010,N_16068,N_16062);
nor U17011 (N_17011,N_16900,N_16590);
xnor U17012 (N_17012,N_16822,N_16851);
xnor U17013 (N_17013,N_16259,N_16899);
nand U17014 (N_17014,N_16395,N_16502);
xnor U17015 (N_17015,N_16563,N_16117);
nor U17016 (N_17016,N_16135,N_16407);
xor U17017 (N_17017,N_16745,N_16027);
nand U17018 (N_17018,N_16241,N_16782);
xor U17019 (N_17019,N_16690,N_16882);
or U17020 (N_17020,N_16878,N_16527);
or U17021 (N_17021,N_16756,N_16328);
and U17022 (N_17022,N_16072,N_16569);
or U17023 (N_17023,N_16653,N_16111);
nand U17024 (N_17024,N_16573,N_16846);
nand U17025 (N_17025,N_16630,N_16393);
nand U17026 (N_17026,N_16513,N_16808);
nor U17027 (N_17027,N_16585,N_16044);
xor U17028 (N_17028,N_16752,N_16872);
nand U17029 (N_17029,N_16277,N_16108);
nor U17030 (N_17030,N_16193,N_16762);
nor U17031 (N_17031,N_16491,N_16689);
nor U17032 (N_17032,N_16048,N_16746);
nor U17033 (N_17033,N_16633,N_16459);
xor U17034 (N_17034,N_16858,N_16795);
or U17035 (N_17035,N_16097,N_16183);
nor U17036 (N_17036,N_16285,N_16673);
nor U17037 (N_17037,N_16521,N_16837);
xnor U17038 (N_17038,N_16280,N_16397);
xor U17039 (N_17039,N_16028,N_16890);
or U17040 (N_17040,N_16042,N_16192);
nor U17041 (N_17041,N_16610,N_16550);
nor U17042 (N_17042,N_16251,N_16123);
xnor U17043 (N_17043,N_16071,N_16312);
and U17044 (N_17044,N_16368,N_16707);
nand U17045 (N_17045,N_16379,N_16972);
and U17046 (N_17046,N_16852,N_16616);
xnor U17047 (N_17047,N_16926,N_16834);
xor U17048 (N_17048,N_16001,N_16939);
nand U17049 (N_17049,N_16578,N_16528);
and U17050 (N_17050,N_16242,N_16996);
xor U17051 (N_17051,N_16284,N_16056);
xor U17052 (N_17052,N_16642,N_16225);
and U17053 (N_17053,N_16418,N_16091);
nor U17054 (N_17054,N_16820,N_16092);
nand U17055 (N_17055,N_16211,N_16420);
xor U17056 (N_17056,N_16703,N_16230);
nor U17057 (N_17057,N_16560,N_16166);
and U17058 (N_17058,N_16295,N_16726);
nand U17059 (N_17059,N_16322,N_16419);
xnor U17060 (N_17060,N_16207,N_16069);
and U17061 (N_17061,N_16853,N_16957);
and U17062 (N_17062,N_16611,N_16990);
nor U17063 (N_17063,N_16351,N_16264);
or U17064 (N_17064,N_16916,N_16980);
or U17065 (N_17065,N_16389,N_16576);
and U17066 (N_17066,N_16710,N_16920);
or U17067 (N_17067,N_16704,N_16780);
nand U17068 (N_17068,N_16338,N_16716);
xor U17069 (N_17069,N_16064,N_16382);
or U17070 (N_17070,N_16544,N_16961);
nand U17071 (N_17071,N_16315,N_16260);
and U17072 (N_17072,N_16529,N_16682);
or U17073 (N_17073,N_16517,N_16336);
nor U17074 (N_17074,N_16962,N_16128);
or U17075 (N_17075,N_16605,N_16153);
and U17076 (N_17076,N_16798,N_16742);
nor U17077 (N_17077,N_16771,N_16253);
or U17078 (N_17078,N_16905,N_16250);
or U17079 (N_17079,N_16779,N_16927);
nand U17080 (N_17080,N_16602,N_16791);
xor U17081 (N_17081,N_16744,N_16023);
nor U17082 (N_17082,N_16469,N_16405);
or U17083 (N_17083,N_16969,N_16354);
nor U17084 (N_17084,N_16627,N_16532);
nand U17085 (N_17085,N_16214,N_16383);
and U17086 (N_17086,N_16334,N_16786);
nand U17087 (N_17087,N_16505,N_16674);
or U17088 (N_17088,N_16217,N_16538);
xor U17089 (N_17089,N_16258,N_16272);
xnor U17090 (N_17090,N_16432,N_16688);
xnor U17091 (N_17091,N_16620,N_16361);
or U17092 (N_17092,N_16483,N_16457);
and U17093 (N_17093,N_16235,N_16219);
and U17094 (N_17094,N_16612,N_16970);
and U17095 (N_17095,N_16227,N_16933);
and U17096 (N_17096,N_16765,N_16271);
or U17097 (N_17097,N_16187,N_16324);
xnor U17098 (N_17098,N_16384,N_16617);
nor U17099 (N_17099,N_16317,N_16196);
nor U17100 (N_17100,N_16588,N_16516);
and U17101 (N_17101,N_16120,N_16238);
and U17102 (N_17102,N_16824,N_16014);
nor U17103 (N_17103,N_16755,N_16931);
nor U17104 (N_17104,N_16377,N_16306);
and U17105 (N_17105,N_16794,N_16537);
or U17106 (N_17106,N_16190,N_16850);
nor U17107 (N_17107,N_16113,N_16199);
xnor U17108 (N_17108,N_16252,N_16959);
nor U17109 (N_17109,N_16904,N_16448);
xor U17110 (N_17110,N_16353,N_16276);
nor U17111 (N_17111,N_16813,N_16341);
nor U17112 (N_17112,N_16936,N_16706);
nand U17113 (N_17113,N_16995,N_16655);
and U17114 (N_17114,N_16168,N_16347);
and U17115 (N_17115,N_16447,N_16760);
and U17116 (N_17116,N_16945,N_16803);
nand U17117 (N_17117,N_16533,N_16650);
or U17118 (N_17118,N_16868,N_16019);
and U17119 (N_17119,N_16006,N_16938);
nor U17120 (N_17120,N_16589,N_16895);
xor U17121 (N_17121,N_16835,N_16804);
xnor U17122 (N_17122,N_16137,N_16016);
nor U17123 (N_17123,N_16138,N_16993);
and U17124 (N_17124,N_16793,N_16671);
and U17125 (N_17125,N_16554,N_16018);
xor U17126 (N_17126,N_16387,N_16313);
nand U17127 (N_17127,N_16208,N_16281);
or U17128 (N_17128,N_16928,N_16649);
or U17129 (N_17129,N_16442,N_16519);
and U17130 (N_17130,N_16778,N_16444);
nor U17131 (N_17131,N_16925,N_16005);
or U17132 (N_17132,N_16559,N_16712);
or U17133 (N_17133,N_16883,N_16240);
nor U17134 (N_17134,N_16035,N_16609);
and U17135 (N_17135,N_16220,N_16713);
nand U17136 (N_17136,N_16600,N_16860);
nand U17137 (N_17137,N_16039,N_16133);
or U17138 (N_17138,N_16719,N_16479);
nand U17139 (N_17139,N_16848,N_16063);
or U17140 (N_17140,N_16057,N_16263);
nor U17141 (N_17141,N_16735,N_16049);
nor U17142 (N_17142,N_16294,N_16046);
nand U17143 (N_17143,N_16823,N_16681);
and U17144 (N_17144,N_16663,N_16864);
and U17145 (N_17145,N_16549,N_16484);
nand U17146 (N_17146,N_16174,N_16090);
xor U17147 (N_17147,N_16767,N_16401);
and U17148 (N_17148,N_16412,N_16162);
nand U17149 (N_17149,N_16314,N_16374);
and U17150 (N_17150,N_16917,N_16818);
or U17151 (N_17151,N_16182,N_16426);
nor U17152 (N_17152,N_16591,N_16723);
nor U17153 (N_17153,N_16662,N_16159);
xor U17154 (N_17154,N_16380,N_16698);
xor U17155 (N_17155,N_16526,N_16799);
nor U17156 (N_17156,N_16262,N_16751);
and U17157 (N_17157,N_16098,N_16077);
nor U17158 (N_17158,N_16366,N_16950);
xnor U17159 (N_17159,N_16392,N_16825);
xor U17160 (N_17160,N_16845,N_16919);
and U17161 (N_17161,N_16148,N_16634);
nand U17162 (N_17162,N_16222,N_16523);
or U17163 (N_17163,N_16507,N_16810);
or U17164 (N_17164,N_16093,N_16855);
and U17165 (N_17165,N_16540,N_16126);
and U17166 (N_17166,N_16886,N_16816);
or U17167 (N_17167,N_16819,N_16370);
or U17168 (N_17168,N_16989,N_16884);
nor U17169 (N_17169,N_16496,N_16267);
or U17170 (N_17170,N_16555,N_16177);
and U17171 (N_17171,N_16398,N_16246);
xnor U17172 (N_17172,N_16856,N_16893);
nor U17173 (N_17173,N_16223,N_16923);
xnor U17174 (N_17174,N_16988,N_16299);
nor U17175 (N_17175,N_16814,N_16955);
or U17176 (N_17176,N_16525,N_16124);
xnor U17177 (N_17177,N_16621,N_16141);
and U17178 (N_17178,N_16115,N_16968);
xor U17179 (N_17179,N_16435,N_16311);
nand U17180 (N_17180,N_16200,N_16015);
nor U17181 (N_17181,N_16871,N_16558);
or U17182 (N_17182,N_16075,N_16282);
or U17183 (N_17183,N_16058,N_16105);
xor U17184 (N_17184,N_16415,N_16708);
and U17185 (N_17185,N_16880,N_16759);
xnor U17186 (N_17186,N_16358,N_16360);
nand U17187 (N_17187,N_16041,N_16615);
nand U17188 (N_17188,N_16583,N_16140);
or U17189 (N_17189,N_16644,N_16709);
or U17190 (N_17190,N_16189,N_16943);
or U17191 (N_17191,N_16215,N_16720);
and U17192 (N_17192,N_16971,N_16065);
and U17193 (N_17193,N_16008,N_16036);
nand U17194 (N_17194,N_16781,N_16302);
or U17195 (N_17195,N_16535,N_16757);
xnor U17196 (N_17196,N_16821,N_16078);
xor U17197 (N_17197,N_16118,N_16462);
nor U17198 (N_17198,N_16982,N_16503);
nand U17199 (N_17199,N_16572,N_16287);
nand U17200 (N_17200,N_16386,N_16290);
nor U17201 (N_17201,N_16186,N_16547);
nand U17202 (N_17202,N_16577,N_16331);
xor U17203 (N_17203,N_16838,N_16458);
and U17204 (N_17204,N_16908,N_16425);
and U17205 (N_17205,N_16656,N_16929);
xor U17206 (N_17206,N_16030,N_16658);
and U17207 (N_17207,N_16348,N_16408);
nand U17208 (N_17208,N_16342,N_16866);
and U17209 (N_17209,N_16983,N_16870);
and U17210 (N_17210,N_16226,N_16343);
xor U17211 (N_17211,N_16815,N_16842);
xnor U17212 (N_17212,N_16461,N_16307);
nand U17213 (N_17213,N_16902,N_16326);
or U17214 (N_17214,N_16731,N_16512);
xnor U17215 (N_17215,N_16520,N_16244);
and U17216 (N_17216,N_16404,N_16715);
nor U17217 (N_17217,N_16668,N_16754);
nor U17218 (N_17218,N_16472,N_16500);
nor U17219 (N_17219,N_16511,N_16732);
or U17220 (N_17220,N_16439,N_16032);
and U17221 (N_17221,N_16454,N_16085);
xor U17222 (N_17222,N_16665,N_16443);
xnor U17223 (N_17223,N_16954,N_16865);
nand U17224 (N_17224,N_16099,N_16721);
or U17225 (N_17225,N_16729,N_16020);
nand U17226 (N_17226,N_16965,N_16421);
or U17227 (N_17227,N_16994,N_16785);
nor U17228 (N_17228,N_16792,N_16188);
or U17229 (N_17229,N_16243,N_16985);
or U17230 (N_17230,N_16089,N_16566);
nand U17231 (N_17231,N_16501,N_16021);
xor U17232 (N_17232,N_16467,N_16891);
and U17233 (N_17233,N_16086,N_16385);
nand U17234 (N_17234,N_16034,N_16691);
or U17235 (N_17235,N_16869,N_16770);
xor U17236 (N_17236,N_16722,N_16390);
nand U17237 (N_17237,N_16847,N_16981);
nand U17238 (N_17238,N_16998,N_16743);
nand U17239 (N_17239,N_16645,N_16209);
nand U17240 (N_17240,N_16495,N_16509);
and U17241 (N_17241,N_16273,N_16934);
nor U17242 (N_17242,N_16127,N_16234);
xor U17243 (N_17243,N_16010,N_16414);
and U17244 (N_17244,N_16007,N_16073);
xnor U17245 (N_17245,N_16158,N_16918);
and U17246 (N_17246,N_16897,N_16599);
xor U17247 (N_17247,N_16876,N_16130);
nand U17248 (N_17248,N_16967,N_16172);
xnor U17249 (N_17249,N_16912,N_16739);
and U17250 (N_17250,N_16693,N_16333);
or U17251 (N_17251,N_16449,N_16275);
xor U17252 (N_17252,N_16508,N_16321);
nand U17253 (N_17253,N_16473,N_16930);
xor U17254 (N_17254,N_16861,N_16146);
xnor U17255 (N_17255,N_16608,N_16403);
or U17256 (N_17256,N_16635,N_16080);
nor U17257 (N_17257,N_16687,N_16921);
xnor U17258 (N_17258,N_16678,N_16074);
xor U17259 (N_17259,N_16518,N_16051);
nand U17260 (N_17260,N_16647,N_16316);
nand U17261 (N_17261,N_16436,N_16987);
nor U17262 (N_17262,N_16265,N_16178);
xnor U17263 (N_17263,N_16817,N_16216);
nand U17264 (N_17264,N_16797,N_16632);
nand U17265 (N_17265,N_16867,N_16011);
nor U17266 (N_17266,N_16670,N_16300);
nand U17267 (N_17267,N_16329,N_16429);
nand U17268 (N_17268,N_16849,N_16323);
and U17269 (N_17269,N_16801,N_16593);
nand U17270 (N_17270,N_16037,N_16740);
nor U17271 (N_17271,N_16788,N_16237);
and U17272 (N_17272,N_16292,N_16543);
or U17273 (N_17273,N_16613,N_16571);
nand U17274 (N_17274,N_16686,N_16601);
xnor U17275 (N_17275,N_16409,N_16974);
nor U17276 (N_17276,N_16477,N_16664);
or U17277 (N_17277,N_16318,N_16734);
and U17278 (N_17278,N_16083,N_16154);
nand U17279 (N_17279,N_16109,N_16411);
nor U17280 (N_17280,N_16807,N_16000);
and U17281 (N_17281,N_16701,N_16832);
nor U17282 (N_17282,N_16881,N_16909);
nand U17283 (N_17283,N_16356,N_16646);
nand U17284 (N_17284,N_16013,N_16233);
nand U17285 (N_17285,N_16595,N_16198);
and U17286 (N_17286,N_16004,N_16684);
nand U17287 (N_17287,N_16119,N_16935);
or U17288 (N_17288,N_16789,N_16705);
xor U17289 (N_17289,N_16924,N_16450);
or U17290 (N_17290,N_16986,N_16297);
nor U17291 (N_17291,N_16696,N_16660);
xor U17292 (N_17292,N_16308,N_16066);
nor U17293 (N_17293,N_16344,N_16677);
xor U17294 (N_17294,N_16622,N_16197);
or U17295 (N_17295,N_16640,N_16661);
nand U17296 (N_17296,N_16906,N_16176);
xor U17297 (N_17297,N_16433,N_16654);
xnor U17298 (N_17298,N_16094,N_16561);
and U17299 (N_17299,N_16106,N_16232);
nor U17300 (N_17300,N_16301,N_16337);
xnor U17301 (N_17301,N_16303,N_16733);
and U17302 (N_17302,N_16125,N_16603);
and U17303 (N_17303,N_16641,N_16941);
and U17304 (N_17304,N_16180,N_16598);
and U17305 (N_17305,N_16060,N_16371);
and U17306 (N_17306,N_16874,N_16592);
xor U17307 (N_17307,N_16156,N_16749);
nand U17308 (N_17308,N_16460,N_16052);
nor U17309 (N_17309,N_16185,N_16914);
nor U17310 (N_17310,N_16506,N_16475);
and U17311 (N_17311,N_16012,N_16680);
or U17312 (N_17312,N_16485,N_16424);
and U17313 (N_17313,N_16570,N_16061);
nand U17314 (N_17314,N_16402,N_16164);
and U17315 (N_17315,N_16221,N_16470);
and U17316 (N_17316,N_16753,N_16149);
nor U17317 (N_17317,N_16910,N_16624);
and U17318 (N_17318,N_16963,N_16979);
xor U17319 (N_17319,N_16776,N_16553);
nor U17320 (N_17320,N_16376,N_16255);
or U17321 (N_17321,N_16026,N_16956);
nand U17322 (N_17322,N_16515,N_16400);
xnor U17323 (N_17323,N_16638,N_16150);
or U17324 (N_17324,N_16932,N_16697);
xnor U17325 (N_17325,N_16427,N_16875);
xor U17326 (N_17326,N_16584,N_16278);
nor U17327 (N_17327,N_16545,N_16958);
nor U17328 (N_17328,N_16946,N_16121);
xnor U17329 (N_17329,N_16679,N_16648);
or U17330 (N_17330,N_16766,N_16350);
nand U17331 (N_17331,N_16873,N_16488);
xnor U17332 (N_17332,N_16254,N_16107);
nand U17333 (N_17333,N_16877,N_16181);
or U17334 (N_17334,N_16717,N_16132);
xnor U17335 (N_17335,N_16806,N_16800);
and U17336 (N_17336,N_16628,N_16487);
and U17337 (N_17337,N_16446,N_16095);
or U17338 (N_17338,N_16490,N_16279);
xnor U17339 (N_17339,N_16976,N_16257);
and U17340 (N_17340,N_16606,N_16079);
and U17341 (N_17341,N_16076,N_16631);
nor U17342 (N_17342,N_16453,N_16579);
xnor U17343 (N_17343,N_16977,N_16204);
xnor U17344 (N_17344,N_16896,N_16143);
or U17345 (N_17345,N_16040,N_16184);
or U17346 (N_17346,N_16349,N_16619);
xnor U17347 (N_17347,N_16388,N_16396);
or U17348 (N_17348,N_16038,N_16964);
and U17349 (N_17349,N_16055,N_16827);
or U17350 (N_17350,N_16694,N_16289);
and U17351 (N_17351,N_16552,N_16784);
nor U17352 (N_17352,N_16145,N_16340);
and U17353 (N_17353,N_16777,N_16594);
and U17354 (N_17354,N_16659,N_16478);
or U17355 (N_17355,N_16541,N_16228);
and U17356 (N_17356,N_16464,N_16607);
or U17357 (N_17357,N_16937,N_16524);
xnor U17358 (N_17358,N_16017,N_16102);
xor U17359 (N_17359,N_16768,N_16155);
nor U17360 (N_17360,N_16718,N_16497);
xnor U17361 (N_17361,N_16542,N_16492);
nand U17362 (N_17362,N_16288,N_16944);
nor U17363 (N_17363,N_16476,N_16167);
and U17364 (N_17364,N_16643,N_16548);
nand U17365 (N_17365,N_16675,N_16562);
nor U17366 (N_17366,N_16352,N_16836);
and U17367 (N_17367,N_16669,N_16863);
or U17368 (N_17368,N_16901,N_16984);
nor U17369 (N_17369,N_16564,N_16493);
or U17370 (N_17370,N_16714,N_16747);
nor U17371 (N_17371,N_16179,N_16966);
nor U17372 (N_17372,N_16463,N_16088);
nor U17373 (N_17373,N_16738,N_16327);
or U17374 (N_17374,N_16103,N_16367);
nor U17375 (N_17375,N_16430,N_16728);
and U17376 (N_17376,N_16203,N_16268);
or U17377 (N_17377,N_16504,N_16748);
xnor U17378 (N_17378,N_16975,N_16758);
xor U17379 (N_17379,N_16339,N_16486);
xnor U17380 (N_17380,N_16831,N_16657);
and U17381 (N_17381,N_16885,N_16911);
nand U17382 (N_17382,N_16951,N_16205);
nor U17383 (N_17383,N_16695,N_16378);
or U17384 (N_17384,N_16913,N_16830);
or U17385 (N_17385,N_16399,N_16889);
nor U17386 (N_17386,N_16261,N_16811);
nand U17387 (N_17387,N_16084,N_16031);
or U17388 (N_17388,N_16854,N_16531);
or U17389 (N_17389,N_16833,N_16626);
nor U17390 (N_17390,N_16171,N_16319);
or U17391 (N_17391,N_16169,N_16978);
nand U17392 (N_17392,N_16614,N_16991);
nor U17393 (N_17393,N_16456,N_16922);
xor U17394 (N_17394,N_16047,N_16355);
or U17395 (N_17395,N_16618,N_16296);
xor U17396 (N_17396,N_16489,N_16249);
nand U17397 (N_17397,N_16774,N_16100);
nor U17398 (N_17398,N_16139,N_16332);
xnor U17399 (N_17399,N_16050,N_16286);
or U17400 (N_17400,N_16152,N_16775);
nand U17401 (N_17401,N_16033,N_16769);
and U17402 (N_17402,N_16330,N_16499);
or U17403 (N_17403,N_16423,N_16116);
xnor U17404 (N_17404,N_16451,N_16212);
and U17405 (N_17405,N_16494,N_16960);
and U17406 (N_17406,N_16997,N_16269);
and U17407 (N_17407,N_16248,N_16373);
xnor U17408 (N_17408,N_16637,N_16580);
nand U17409 (N_17409,N_16346,N_16683);
nor U17410 (N_17410,N_16218,N_16365);
xnor U17411 (N_17411,N_16438,N_16676);
or U17412 (N_17412,N_16236,N_16581);
and U17413 (N_17413,N_16840,N_16231);
xor U17414 (N_17414,N_16029,N_16764);
xnor U17415 (N_17415,N_16692,N_16070);
nor U17416 (N_17416,N_16888,N_16362);
or U17417 (N_17417,N_16841,N_16809);
and U17418 (N_17418,N_16802,N_16134);
nor U17419 (N_17419,N_16522,N_16160);
nor U17420 (N_17420,N_16942,N_16002);
nor U17421 (N_17421,N_16053,N_16952);
nor U17422 (N_17422,N_16163,N_16575);
nand U17423 (N_17423,N_16812,N_16805);
nand U17424 (N_17424,N_16565,N_16586);
nor U17425 (N_17425,N_16067,N_16514);
nor U17426 (N_17426,N_16283,N_16953);
nor U17427 (N_17427,N_16857,N_16700);
nand U17428 (N_17428,N_16245,N_16157);
and U17429 (N_17429,N_16466,N_16843);
nor U17430 (N_17430,N_16325,N_16907);
or U17431 (N_17431,N_16510,N_16557);
or U17432 (N_17432,N_16202,N_16761);
and U17433 (N_17433,N_16101,N_16574);
and U17434 (N_17434,N_16381,N_16947);
and U17435 (N_17435,N_16727,N_16940);
and U17436 (N_17436,N_16112,N_16597);
nand U17437 (N_17437,N_16372,N_16364);
nand U17438 (N_17438,N_16144,N_16266);
nor U17439 (N_17439,N_16892,N_16194);
xnor U17440 (N_17440,N_16195,N_16045);
and U17441 (N_17441,N_16666,N_16711);
xor U17442 (N_17442,N_16498,N_16887);
nand U17443 (N_17443,N_16024,N_16773);
and U17444 (N_17444,N_16191,N_16081);
or U17445 (N_17445,N_16468,N_16667);
xor U17446 (N_17446,N_16465,N_16898);
nor U17447 (N_17447,N_16417,N_16915);
nand U17448 (N_17448,N_16122,N_16894);
or U17449 (N_17449,N_16293,N_16556);
nor U17450 (N_17450,N_16298,N_16416);
and U17451 (N_17451,N_16059,N_16587);
nand U17452 (N_17452,N_16750,N_16536);
xnor U17453 (N_17453,N_16828,N_16839);
and U17454 (N_17454,N_16844,N_16104);
and U17455 (N_17455,N_16672,N_16625);
xnor U17456 (N_17456,N_16165,N_16310);
nor U17457 (N_17457,N_16434,N_16859);
and U17458 (N_17458,N_16741,N_16948);
nor U17459 (N_17459,N_16175,N_16441);
or U17460 (N_17460,N_16410,N_16025);
xor U17461 (N_17461,N_16452,N_16129);
nand U17462 (N_17462,N_16736,N_16206);
or U17463 (N_17463,N_16534,N_16096);
xor U17464 (N_17464,N_16763,N_16730);
nor U17465 (N_17465,N_16567,N_16582);
xor U17466 (N_17466,N_16413,N_16787);
nor U17467 (N_17467,N_16151,N_16480);
or U17468 (N_17468,N_16826,N_16481);
nand U17469 (N_17469,N_16428,N_16445);
nand U17470 (N_17470,N_16639,N_16142);
xor U17471 (N_17471,N_16320,N_16213);
and U17472 (N_17472,N_16304,N_16161);
or U17473 (N_17473,N_16291,N_16147);
nand U17474 (N_17474,N_16903,N_16256);
or U17475 (N_17475,N_16992,N_16546);
or U17476 (N_17476,N_16783,N_16043);
and U17477 (N_17477,N_16239,N_16455);
nor U17478 (N_17478,N_16725,N_16224);
and U17479 (N_17479,N_16082,N_16651);
nor U17480 (N_17480,N_16862,N_16699);
or U17481 (N_17481,N_16136,N_16482);
and U17482 (N_17482,N_16274,N_16406);
nand U17483 (N_17483,N_16247,N_16394);
nor U17484 (N_17484,N_16440,N_16345);
nand U17485 (N_17485,N_16369,N_16309);
nor U17486 (N_17486,N_16305,N_16685);
nand U17487 (N_17487,N_16790,N_16652);
nand U17488 (N_17488,N_16551,N_16422);
nand U17489 (N_17489,N_16829,N_16335);
and U17490 (N_17490,N_16131,N_16363);
nand U17491 (N_17491,N_16796,N_16772);
and U17492 (N_17492,N_16737,N_16022);
nor U17493 (N_17493,N_16636,N_16530);
or U17494 (N_17494,N_16009,N_16087);
and U17495 (N_17495,N_16623,N_16357);
or U17496 (N_17496,N_16629,N_16114);
and U17497 (N_17497,N_16474,N_16604);
and U17498 (N_17498,N_16173,N_16210);
and U17499 (N_17499,N_16170,N_16568);
and U17500 (N_17500,N_16162,N_16349);
or U17501 (N_17501,N_16647,N_16245);
or U17502 (N_17502,N_16264,N_16941);
nor U17503 (N_17503,N_16088,N_16589);
and U17504 (N_17504,N_16591,N_16527);
xnor U17505 (N_17505,N_16961,N_16626);
nand U17506 (N_17506,N_16405,N_16615);
nand U17507 (N_17507,N_16011,N_16596);
nand U17508 (N_17508,N_16199,N_16258);
or U17509 (N_17509,N_16736,N_16251);
nand U17510 (N_17510,N_16537,N_16826);
nor U17511 (N_17511,N_16639,N_16525);
or U17512 (N_17512,N_16792,N_16530);
or U17513 (N_17513,N_16278,N_16495);
nand U17514 (N_17514,N_16454,N_16051);
nand U17515 (N_17515,N_16444,N_16892);
and U17516 (N_17516,N_16498,N_16410);
nand U17517 (N_17517,N_16677,N_16857);
xor U17518 (N_17518,N_16636,N_16670);
nand U17519 (N_17519,N_16449,N_16277);
xnor U17520 (N_17520,N_16298,N_16294);
xor U17521 (N_17521,N_16564,N_16032);
and U17522 (N_17522,N_16321,N_16736);
xnor U17523 (N_17523,N_16399,N_16434);
or U17524 (N_17524,N_16964,N_16337);
nand U17525 (N_17525,N_16359,N_16666);
nor U17526 (N_17526,N_16575,N_16103);
xor U17527 (N_17527,N_16617,N_16904);
nor U17528 (N_17528,N_16627,N_16353);
xor U17529 (N_17529,N_16989,N_16476);
or U17530 (N_17530,N_16305,N_16824);
nor U17531 (N_17531,N_16775,N_16235);
and U17532 (N_17532,N_16132,N_16210);
and U17533 (N_17533,N_16000,N_16588);
and U17534 (N_17534,N_16411,N_16050);
and U17535 (N_17535,N_16078,N_16921);
or U17536 (N_17536,N_16123,N_16669);
or U17537 (N_17537,N_16765,N_16933);
nand U17538 (N_17538,N_16552,N_16935);
nor U17539 (N_17539,N_16166,N_16526);
or U17540 (N_17540,N_16460,N_16141);
nand U17541 (N_17541,N_16466,N_16195);
and U17542 (N_17542,N_16559,N_16599);
and U17543 (N_17543,N_16896,N_16677);
nor U17544 (N_17544,N_16929,N_16788);
and U17545 (N_17545,N_16725,N_16193);
nand U17546 (N_17546,N_16863,N_16651);
and U17547 (N_17547,N_16775,N_16014);
xnor U17548 (N_17548,N_16350,N_16785);
nor U17549 (N_17549,N_16966,N_16881);
xnor U17550 (N_17550,N_16600,N_16451);
xor U17551 (N_17551,N_16228,N_16503);
or U17552 (N_17552,N_16625,N_16344);
or U17553 (N_17553,N_16803,N_16248);
nor U17554 (N_17554,N_16393,N_16267);
nand U17555 (N_17555,N_16940,N_16087);
nand U17556 (N_17556,N_16417,N_16770);
and U17557 (N_17557,N_16170,N_16663);
nand U17558 (N_17558,N_16078,N_16516);
nand U17559 (N_17559,N_16547,N_16189);
nand U17560 (N_17560,N_16654,N_16841);
and U17561 (N_17561,N_16910,N_16921);
nand U17562 (N_17562,N_16818,N_16694);
nand U17563 (N_17563,N_16107,N_16601);
and U17564 (N_17564,N_16426,N_16712);
nand U17565 (N_17565,N_16498,N_16642);
nor U17566 (N_17566,N_16311,N_16006);
xnor U17567 (N_17567,N_16090,N_16139);
nor U17568 (N_17568,N_16263,N_16480);
nor U17569 (N_17569,N_16065,N_16441);
nand U17570 (N_17570,N_16592,N_16196);
nand U17571 (N_17571,N_16092,N_16530);
nand U17572 (N_17572,N_16770,N_16060);
and U17573 (N_17573,N_16385,N_16242);
nand U17574 (N_17574,N_16410,N_16142);
nor U17575 (N_17575,N_16945,N_16659);
nor U17576 (N_17576,N_16072,N_16143);
nor U17577 (N_17577,N_16378,N_16931);
nand U17578 (N_17578,N_16970,N_16107);
and U17579 (N_17579,N_16182,N_16254);
nand U17580 (N_17580,N_16864,N_16473);
nor U17581 (N_17581,N_16895,N_16834);
nand U17582 (N_17582,N_16115,N_16776);
nand U17583 (N_17583,N_16957,N_16252);
or U17584 (N_17584,N_16992,N_16304);
xnor U17585 (N_17585,N_16337,N_16122);
and U17586 (N_17586,N_16262,N_16146);
nand U17587 (N_17587,N_16618,N_16227);
and U17588 (N_17588,N_16413,N_16074);
nand U17589 (N_17589,N_16776,N_16456);
nor U17590 (N_17590,N_16538,N_16155);
or U17591 (N_17591,N_16233,N_16475);
nand U17592 (N_17592,N_16841,N_16430);
or U17593 (N_17593,N_16069,N_16967);
and U17594 (N_17594,N_16203,N_16524);
nand U17595 (N_17595,N_16118,N_16051);
and U17596 (N_17596,N_16693,N_16642);
nand U17597 (N_17597,N_16732,N_16834);
and U17598 (N_17598,N_16037,N_16558);
xor U17599 (N_17599,N_16252,N_16121);
and U17600 (N_17600,N_16906,N_16345);
and U17601 (N_17601,N_16065,N_16231);
nor U17602 (N_17602,N_16035,N_16415);
nand U17603 (N_17603,N_16263,N_16997);
or U17604 (N_17604,N_16491,N_16249);
and U17605 (N_17605,N_16113,N_16642);
and U17606 (N_17606,N_16045,N_16661);
or U17607 (N_17607,N_16419,N_16446);
nand U17608 (N_17608,N_16507,N_16777);
or U17609 (N_17609,N_16911,N_16439);
nand U17610 (N_17610,N_16681,N_16644);
or U17611 (N_17611,N_16291,N_16158);
and U17612 (N_17612,N_16214,N_16853);
and U17613 (N_17613,N_16981,N_16329);
xnor U17614 (N_17614,N_16615,N_16378);
nor U17615 (N_17615,N_16738,N_16662);
or U17616 (N_17616,N_16853,N_16315);
or U17617 (N_17617,N_16103,N_16096);
and U17618 (N_17618,N_16022,N_16497);
xnor U17619 (N_17619,N_16793,N_16903);
nor U17620 (N_17620,N_16771,N_16898);
nor U17621 (N_17621,N_16403,N_16465);
or U17622 (N_17622,N_16495,N_16506);
nand U17623 (N_17623,N_16194,N_16632);
and U17624 (N_17624,N_16845,N_16211);
and U17625 (N_17625,N_16977,N_16574);
nand U17626 (N_17626,N_16747,N_16120);
nand U17627 (N_17627,N_16601,N_16912);
and U17628 (N_17628,N_16428,N_16936);
nand U17629 (N_17629,N_16311,N_16420);
nand U17630 (N_17630,N_16412,N_16059);
nor U17631 (N_17631,N_16480,N_16131);
nand U17632 (N_17632,N_16859,N_16375);
or U17633 (N_17633,N_16781,N_16755);
nand U17634 (N_17634,N_16105,N_16563);
xnor U17635 (N_17635,N_16947,N_16215);
nor U17636 (N_17636,N_16902,N_16363);
or U17637 (N_17637,N_16957,N_16427);
xor U17638 (N_17638,N_16853,N_16155);
nor U17639 (N_17639,N_16982,N_16071);
and U17640 (N_17640,N_16965,N_16540);
nand U17641 (N_17641,N_16018,N_16332);
xor U17642 (N_17642,N_16474,N_16361);
nor U17643 (N_17643,N_16292,N_16375);
xnor U17644 (N_17644,N_16620,N_16658);
nor U17645 (N_17645,N_16301,N_16424);
nand U17646 (N_17646,N_16390,N_16230);
or U17647 (N_17647,N_16702,N_16299);
and U17648 (N_17648,N_16034,N_16421);
and U17649 (N_17649,N_16744,N_16156);
and U17650 (N_17650,N_16761,N_16745);
nor U17651 (N_17651,N_16841,N_16925);
and U17652 (N_17652,N_16146,N_16167);
and U17653 (N_17653,N_16845,N_16788);
or U17654 (N_17654,N_16755,N_16768);
xor U17655 (N_17655,N_16747,N_16281);
nand U17656 (N_17656,N_16800,N_16386);
nand U17657 (N_17657,N_16335,N_16370);
or U17658 (N_17658,N_16980,N_16204);
or U17659 (N_17659,N_16583,N_16754);
and U17660 (N_17660,N_16024,N_16589);
nand U17661 (N_17661,N_16583,N_16653);
nand U17662 (N_17662,N_16096,N_16476);
xnor U17663 (N_17663,N_16317,N_16074);
nor U17664 (N_17664,N_16819,N_16805);
and U17665 (N_17665,N_16129,N_16569);
xor U17666 (N_17666,N_16360,N_16042);
xor U17667 (N_17667,N_16951,N_16758);
nand U17668 (N_17668,N_16038,N_16192);
nand U17669 (N_17669,N_16697,N_16729);
and U17670 (N_17670,N_16191,N_16667);
nand U17671 (N_17671,N_16018,N_16521);
or U17672 (N_17672,N_16848,N_16048);
or U17673 (N_17673,N_16187,N_16737);
and U17674 (N_17674,N_16803,N_16828);
and U17675 (N_17675,N_16980,N_16362);
nand U17676 (N_17676,N_16935,N_16022);
nand U17677 (N_17677,N_16930,N_16956);
or U17678 (N_17678,N_16305,N_16779);
nand U17679 (N_17679,N_16192,N_16136);
or U17680 (N_17680,N_16286,N_16393);
nor U17681 (N_17681,N_16562,N_16210);
or U17682 (N_17682,N_16298,N_16841);
or U17683 (N_17683,N_16182,N_16054);
xor U17684 (N_17684,N_16553,N_16663);
nand U17685 (N_17685,N_16026,N_16797);
and U17686 (N_17686,N_16768,N_16889);
xor U17687 (N_17687,N_16427,N_16853);
nand U17688 (N_17688,N_16173,N_16765);
and U17689 (N_17689,N_16078,N_16068);
and U17690 (N_17690,N_16390,N_16468);
nand U17691 (N_17691,N_16178,N_16767);
nor U17692 (N_17692,N_16214,N_16887);
and U17693 (N_17693,N_16553,N_16417);
nor U17694 (N_17694,N_16203,N_16267);
and U17695 (N_17695,N_16369,N_16478);
xnor U17696 (N_17696,N_16844,N_16684);
xnor U17697 (N_17697,N_16782,N_16829);
nand U17698 (N_17698,N_16632,N_16005);
and U17699 (N_17699,N_16438,N_16624);
nand U17700 (N_17700,N_16790,N_16572);
nand U17701 (N_17701,N_16907,N_16521);
and U17702 (N_17702,N_16682,N_16092);
nand U17703 (N_17703,N_16754,N_16052);
nand U17704 (N_17704,N_16718,N_16962);
nor U17705 (N_17705,N_16876,N_16803);
nor U17706 (N_17706,N_16121,N_16235);
nand U17707 (N_17707,N_16310,N_16388);
xor U17708 (N_17708,N_16486,N_16424);
xnor U17709 (N_17709,N_16440,N_16937);
xnor U17710 (N_17710,N_16905,N_16280);
nand U17711 (N_17711,N_16510,N_16781);
or U17712 (N_17712,N_16081,N_16190);
nor U17713 (N_17713,N_16851,N_16018);
nor U17714 (N_17714,N_16579,N_16874);
nor U17715 (N_17715,N_16570,N_16343);
or U17716 (N_17716,N_16117,N_16660);
xnor U17717 (N_17717,N_16254,N_16463);
nand U17718 (N_17718,N_16517,N_16717);
and U17719 (N_17719,N_16947,N_16459);
and U17720 (N_17720,N_16809,N_16548);
nand U17721 (N_17721,N_16226,N_16693);
nor U17722 (N_17722,N_16706,N_16349);
xor U17723 (N_17723,N_16167,N_16679);
xor U17724 (N_17724,N_16420,N_16320);
or U17725 (N_17725,N_16640,N_16929);
nor U17726 (N_17726,N_16325,N_16518);
nor U17727 (N_17727,N_16001,N_16765);
xnor U17728 (N_17728,N_16974,N_16772);
or U17729 (N_17729,N_16741,N_16023);
xor U17730 (N_17730,N_16983,N_16277);
xnor U17731 (N_17731,N_16249,N_16457);
nand U17732 (N_17732,N_16360,N_16381);
nor U17733 (N_17733,N_16713,N_16894);
or U17734 (N_17734,N_16647,N_16613);
nand U17735 (N_17735,N_16769,N_16836);
and U17736 (N_17736,N_16910,N_16503);
and U17737 (N_17737,N_16145,N_16574);
nand U17738 (N_17738,N_16319,N_16614);
xnor U17739 (N_17739,N_16616,N_16868);
xor U17740 (N_17740,N_16787,N_16063);
xnor U17741 (N_17741,N_16754,N_16765);
nand U17742 (N_17742,N_16185,N_16152);
xor U17743 (N_17743,N_16092,N_16284);
xnor U17744 (N_17744,N_16047,N_16514);
nand U17745 (N_17745,N_16826,N_16197);
and U17746 (N_17746,N_16054,N_16948);
and U17747 (N_17747,N_16086,N_16886);
or U17748 (N_17748,N_16676,N_16407);
xnor U17749 (N_17749,N_16360,N_16131);
xnor U17750 (N_17750,N_16581,N_16584);
nor U17751 (N_17751,N_16534,N_16982);
nand U17752 (N_17752,N_16185,N_16826);
nand U17753 (N_17753,N_16120,N_16194);
and U17754 (N_17754,N_16820,N_16922);
and U17755 (N_17755,N_16275,N_16667);
nand U17756 (N_17756,N_16108,N_16020);
nor U17757 (N_17757,N_16173,N_16679);
nand U17758 (N_17758,N_16067,N_16533);
xnor U17759 (N_17759,N_16778,N_16244);
nor U17760 (N_17760,N_16436,N_16398);
xnor U17761 (N_17761,N_16434,N_16146);
nor U17762 (N_17762,N_16542,N_16375);
nor U17763 (N_17763,N_16370,N_16006);
xnor U17764 (N_17764,N_16211,N_16725);
nand U17765 (N_17765,N_16276,N_16518);
or U17766 (N_17766,N_16151,N_16269);
nand U17767 (N_17767,N_16395,N_16478);
nor U17768 (N_17768,N_16047,N_16885);
or U17769 (N_17769,N_16138,N_16691);
xnor U17770 (N_17770,N_16181,N_16298);
xor U17771 (N_17771,N_16447,N_16554);
nand U17772 (N_17772,N_16061,N_16745);
xor U17773 (N_17773,N_16076,N_16380);
nand U17774 (N_17774,N_16954,N_16171);
or U17775 (N_17775,N_16366,N_16222);
nand U17776 (N_17776,N_16975,N_16969);
nor U17777 (N_17777,N_16843,N_16695);
nand U17778 (N_17778,N_16719,N_16586);
or U17779 (N_17779,N_16013,N_16781);
or U17780 (N_17780,N_16905,N_16126);
and U17781 (N_17781,N_16328,N_16144);
and U17782 (N_17782,N_16134,N_16431);
nor U17783 (N_17783,N_16882,N_16936);
or U17784 (N_17784,N_16800,N_16873);
xor U17785 (N_17785,N_16563,N_16525);
nor U17786 (N_17786,N_16636,N_16753);
or U17787 (N_17787,N_16569,N_16654);
or U17788 (N_17788,N_16828,N_16445);
xor U17789 (N_17789,N_16791,N_16056);
xnor U17790 (N_17790,N_16682,N_16541);
nand U17791 (N_17791,N_16153,N_16577);
and U17792 (N_17792,N_16796,N_16497);
or U17793 (N_17793,N_16898,N_16228);
or U17794 (N_17794,N_16710,N_16779);
or U17795 (N_17795,N_16823,N_16558);
and U17796 (N_17796,N_16706,N_16608);
nor U17797 (N_17797,N_16726,N_16957);
xor U17798 (N_17798,N_16200,N_16273);
or U17799 (N_17799,N_16851,N_16542);
or U17800 (N_17800,N_16898,N_16275);
or U17801 (N_17801,N_16602,N_16954);
nand U17802 (N_17802,N_16983,N_16114);
nand U17803 (N_17803,N_16488,N_16804);
or U17804 (N_17804,N_16527,N_16135);
nand U17805 (N_17805,N_16766,N_16850);
or U17806 (N_17806,N_16764,N_16991);
or U17807 (N_17807,N_16654,N_16272);
or U17808 (N_17808,N_16941,N_16568);
and U17809 (N_17809,N_16906,N_16130);
and U17810 (N_17810,N_16524,N_16306);
xor U17811 (N_17811,N_16505,N_16616);
nand U17812 (N_17812,N_16736,N_16851);
nand U17813 (N_17813,N_16223,N_16568);
or U17814 (N_17814,N_16307,N_16502);
and U17815 (N_17815,N_16209,N_16050);
nand U17816 (N_17816,N_16824,N_16328);
xnor U17817 (N_17817,N_16730,N_16228);
or U17818 (N_17818,N_16750,N_16282);
or U17819 (N_17819,N_16691,N_16732);
xnor U17820 (N_17820,N_16129,N_16936);
or U17821 (N_17821,N_16041,N_16167);
and U17822 (N_17822,N_16518,N_16435);
and U17823 (N_17823,N_16791,N_16352);
nand U17824 (N_17824,N_16640,N_16031);
and U17825 (N_17825,N_16023,N_16576);
and U17826 (N_17826,N_16401,N_16656);
nor U17827 (N_17827,N_16516,N_16404);
nor U17828 (N_17828,N_16240,N_16139);
nand U17829 (N_17829,N_16203,N_16432);
xnor U17830 (N_17830,N_16415,N_16400);
or U17831 (N_17831,N_16179,N_16529);
nor U17832 (N_17832,N_16673,N_16626);
nor U17833 (N_17833,N_16528,N_16437);
and U17834 (N_17834,N_16957,N_16623);
nor U17835 (N_17835,N_16856,N_16503);
nand U17836 (N_17836,N_16290,N_16585);
nand U17837 (N_17837,N_16472,N_16328);
xor U17838 (N_17838,N_16735,N_16809);
nor U17839 (N_17839,N_16251,N_16850);
nor U17840 (N_17840,N_16340,N_16541);
or U17841 (N_17841,N_16909,N_16341);
or U17842 (N_17842,N_16912,N_16044);
xor U17843 (N_17843,N_16444,N_16684);
and U17844 (N_17844,N_16013,N_16642);
nand U17845 (N_17845,N_16473,N_16191);
nor U17846 (N_17846,N_16297,N_16554);
and U17847 (N_17847,N_16107,N_16620);
nand U17848 (N_17848,N_16964,N_16305);
or U17849 (N_17849,N_16719,N_16495);
nor U17850 (N_17850,N_16922,N_16660);
and U17851 (N_17851,N_16510,N_16966);
nor U17852 (N_17852,N_16741,N_16877);
nor U17853 (N_17853,N_16547,N_16845);
nand U17854 (N_17854,N_16331,N_16169);
nor U17855 (N_17855,N_16298,N_16413);
xor U17856 (N_17856,N_16574,N_16619);
and U17857 (N_17857,N_16404,N_16218);
nand U17858 (N_17858,N_16085,N_16510);
nand U17859 (N_17859,N_16098,N_16936);
xor U17860 (N_17860,N_16633,N_16914);
nor U17861 (N_17861,N_16273,N_16307);
and U17862 (N_17862,N_16668,N_16504);
nor U17863 (N_17863,N_16339,N_16026);
or U17864 (N_17864,N_16135,N_16050);
or U17865 (N_17865,N_16473,N_16485);
nor U17866 (N_17866,N_16678,N_16091);
nand U17867 (N_17867,N_16342,N_16294);
and U17868 (N_17868,N_16782,N_16413);
xor U17869 (N_17869,N_16823,N_16712);
xor U17870 (N_17870,N_16324,N_16519);
nor U17871 (N_17871,N_16033,N_16342);
nor U17872 (N_17872,N_16015,N_16889);
or U17873 (N_17873,N_16810,N_16621);
nor U17874 (N_17874,N_16927,N_16591);
nor U17875 (N_17875,N_16930,N_16907);
and U17876 (N_17876,N_16342,N_16552);
or U17877 (N_17877,N_16452,N_16121);
nand U17878 (N_17878,N_16832,N_16727);
and U17879 (N_17879,N_16328,N_16096);
nand U17880 (N_17880,N_16309,N_16263);
nor U17881 (N_17881,N_16397,N_16630);
nand U17882 (N_17882,N_16639,N_16004);
xor U17883 (N_17883,N_16108,N_16432);
nand U17884 (N_17884,N_16953,N_16794);
nand U17885 (N_17885,N_16330,N_16039);
and U17886 (N_17886,N_16420,N_16441);
or U17887 (N_17887,N_16130,N_16904);
nand U17888 (N_17888,N_16819,N_16542);
and U17889 (N_17889,N_16950,N_16625);
nor U17890 (N_17890,N_16807,N_16952);
or U17891 (N_17891,N_16252,N_16199);
xnor U17892 (N_17892,N_16188,N_16391);
nand U17893 (N_17893,N_16958,N_16136);
xor U17894 (N_17894,N_16069,N_16072);
and U17895 (N_17895,N_16673,N_16447);
nor U17896 (N_17896,N_16081,N_16612);
xnor U17897 (N_17897,N_16116,N_16133);
nand U17898 (N_17898,N_16772,N_16650);
xor U17899 (N_17899,N_16175,N_16779);
xnor U17900 (N_17900,N_16228,N_16607);
and U17901 (N_17901,N_16205,N_16840);
xor U17902 (N_17902,N_16569,N_16547);
and U17903 (N_17903,N_16474,N_16005);
nand U17904 (N_17904,N_16157,N_16277);
or U17905 (N_17905,N_16513,N_16712);
nand U17906 (N_17906,N_16009,N_16341);
or U17907 (N_17907,N_16527,N_16495);
or U17908 (N_17908,N_16786,N_16397);
or U17909 (N_17909,N_16823,N_16795);
nor U17910 (N_17910,N_16837,N_16274);
and U17911 (N_17911,N_16470,N_16339);
xor U17912 (N_17912,N_16764,N_16036);
or U17913 (N_17913,N_16159,N_16772);
nor U17914 (N_17914,N_16771,N_16999);
and U17915 (N_17915,N_16757,N_16918);
or U17916 (N_17916,N_16225,N_16262);
nand U17917 (N_17917,N_16021,N_16448);
or U17918 (N_17918,N_16174,N_16186);
xor U17919 (N_17919,N_16574,N_16387);
and U17920 (N_17920,N_16677,N_16142);
and U17921 (N_17921,N_16200,N_16971);
and U17922 (N_17922,N_16568,N_16816);
nor U17923 (N_17923,N_16400,N_16661);
nand U17924 (N_17924,N_16636,N_16500);
or U17925 (N_17925,N_16190,N_16354);
nor U17926 (N_17926,N_16388,N_16959);
xor U17927 (N_17927,N_16853,N_16081);
nand U17928 (N_17928,N_16341,N_16699);
or U17929 (N_17929,N_16720,N_16704);
and U17930 (N_17930,N_16006,N_16549);
xor U17931 (N_17931,N_16848,N_16169);
nand U17932 (N_17932,N_16629,N_16066);
xor U17933 (N_17933,N_16984,N_16565);
xnor U17934 (N_17934,N_16039,N_16523);
nand U17935 (N_17935,N_16337,N_16199);
xnor U17936 (N_17936,N_16021,N_16778);
or U17937 (N_17937,N_16197,N_16181);
xor U17938 (N_17938,N_16155,N_16219);
or U17939 (N_17939,N_16477,N_16228);
or U17940 (N_17940,N_16800,N_16282);
nand U17941 (N_17941,N_16911,N_16777);
xor U17942 (N_17942,N_16355,N_16816);
xor U17943 (N_17943,N_16363,N_16528);
and U17944 (N_17944,N_16546,N_16111);
nand U17945 (N_17945,N_16803,N_16802);
nor U17946 (N_17946,N_16171,N_16660);
and U17947 (N_17947,N_16543,N_16915);
nor U17948 (N_17948,N_16687,N_16652);
nor U17949 (N_17949,N_16999,N_16930);
xor U17950 (N_17950,N_16252,N_16736);
xor U17951 (N_17951,N_16534,N_16780);
xnor U17952 (N_17952,N_16092,N_16234);
or U17953 (N_17953,N_16263,N_16040);
nor U17954 (N_17954,N_16606,N_16284);
nand U17955 (N_17955,N_16294,N_16087);
xnor U17956 (N_17956,N_16709,N_16706);
nand U17957 (N_17957,N_16032,N_16982);
or U17958 (N_17958,N_16963,N_16388);
and U17959 (N_17959,N_16603,N_16471);
nand U17960 (N_17960,N_16816,N_16976);
nand U17961 (N_17961,N_16456,N_16430);
or U17962 (N_17962,N_16723,N_16681);
and U17963 (N_17963,N_16238,N_16059);
or U17964 (N_17964,N_16227,N_16335);
nor U17965 (N_17965,N_16662,N_16322);
xor U17966 (N_17966,N_16565,N_16665);
nor U17967 (N_17967,N_16995,N_16452);
or U17968 (N_17968,N_16684,N_16005);
nand U17969 (N_17969,N_16636,N_16495);
xnor U17970 (N_17970,N_16847,N_16437);
xor U17971 (N_17971,N_16014,N_16180);
nand U17972 (N_17972,N_16355,N_16191);
nand U17973 (N_17973,N_16090,N_16689);
or U17974 (N_17974,N_16759,N_16574);
nor U17975 (N_17975,N_16386,N_16390);
nand U17976 (N_17976,N_16376,N_16762);
nand U17977 (N_17977,N_16632,N_16481);
and U17978 (N_17978,N_16290,N_16874);
or U17979 (N_17979,N_16101,N_16285);
xor U17980 (N_17980,N_16606,N_16340);
nor U17981 (N_17981,N_16549,N_16321);
and U17982 (N_17982,N_16136,N_16214);
nor U17983 (N_17983,N_16623,N_16182);
xor U17984 (N_17984,N_16872,N_16439);
and U17985 (N_17985,N_16884,N_16939);
nand U17986 (N_17986,N_16131,N_16444);
or U17987 (N_17987,N_16764,N_16973);
xor U17988 (N_17988,N_16649,N_16447);
or U17989 (N_17989,N_16737,N_16993);
nor U17990 (N_17990,N_16117,N_16902);
nor U17991 (N_17991,N_16013,N_16957);
xor U17992 (N_17992,N_16947,N_16635);
nor U17993 (N_17993,N_16601,N_16882);
nand U17994 (N_17994,N_16444,N_16496);
or U17995 (N_17995,N_16710,N_16009);
xnor U17996 (N_17996,N_16543,N_16794);
xor U17997 (N_17997,N_16360,N_16125);
xnor U17998 (N_17998,N_16571,N_16387);
or U17999 (N_17999,N_16630,N_16350);
xor U18000 (N_18000,N_17266,N_17735);
or U18001 (N_18001,N_17200,N_17288);
or U18002 (N_18002,N_17438,N_17111);
and U18003 (N_18003,N_17561,N_17258);
or U18004 (N_18004,N_17477,N_17282);
xnor U18005 (N_18005,N_17113,N_17248);
nor U18006 (N_18006,N_17413,N_17498);
xnor U18007 (N_18007,N_17660,N_17900);
nor U18008 (N_18008,N_17131,N_17965);
nand U18009 (N_18009,N_17488,N_17124);
nand U18010 (N_18010,N_17220,N_17336);
nor U18011 (N_18011,N_17354,N_17208);
xor U18012 (N_18012,N_17516,N_17351);
or U18013 (N_18013,N_17221,N_17217);
nand U18014 (N_18014,N_17355,N_17983);
xor U18015 (N_18015,N_17261,N_17385);
or U18016 (N_18016,N_17320,N_17633);
or U18017 (N_18017,N_17155,N_17985);
nand U18018 (N_18018,N_17144,N_17140);
nand U18019 (N_18019,N_17218,N_17193);
nor U18020 (N_18020,N_17453,N_17305);
xnor U18021 (N_18021,N_17340,N_17089);
xor U18022 (N_18022,N_17970,N_17606);
and U18023 (N_18023,N_17007,N_17454);
and U18024 (N_18024,N_17800,N_17790);
xor U18025 (N_18025,N_17923,N_17115);
and U18026 (N_18026,N_17005,N_17520);
and U18027 (N_18027,N_17695,N_17298);
and U18028 (N_18028,N_17246,N_17887);
or U18029 (N_18029,N_17977,N_17074);
and U18030 (N_18030,N_17646,N_17830);
nor U18031 (N_18031,N_17540,N_17511);
xnor U18032 (N_18032,N_17749,N_17651);
or U18033 (N_18033,N_17460,N_17592);
nand U18034 (N_18034,N_17291,N_17116);
xnor U18035 (N_18035,N_17570,N_17507);
or U18036 (N_18036,N_17079,N_17768);
or U18037 (N_18037,N_17035,N_17058);
nand U18038 (N_18038,N_17741,N_17049);
or U18039 (N_18039,N_17294,N_17710);
or U18040 (N_18040,N_17988,N_17734);
or U18041 (N_18041,N_17743,N_17024);
nor U18042 (N_18042,N_17350,N_17362);
or U18043 (N_18043,N_17941,N_17833);
and U18044 (N_18044,N_17521,N_17622);
or U18045 (N_18045,N_17764,N_17630);
xor U18046 (N_18046,N_17730,N_17102);
xnor U18047 (N_18047,N_17014,N_17077);
or U18048 (N_18048,N_17605,N_17034);
and U18049 (N_18049,N_17067,N_17657);
and U18050 (N_18050,N_17012,N_17348);
nand U18051 (N_18051,N_17062,N_17231);
xnor U18052 (N_18052,N_17125,N_17372);
nand U18053 (N_18053,N_17636,N_17788);
and U18054 (N_18054,N_17100,N_17553);
and U18055 (N_18055,N_17127,N_17342);
or U18056 (N_18056,N_17653,N_17022);
and U18057 (N_18057,N_17037,N_17275);
and U18058 (N_18058,N_17552,N_17006);
xnor U18059 (N_18059,N_17823,N_17137);
nor U18060 (N_18060,N_17361,N_17237);
xnor U18061 (N_18061,N_17821,N_17724);
or U18062 (N_18062,N_17343,N_17652);
xor U18063 (N_18063,N_17108,N_17283);
nor U18064 (N_18064,N_17370,N_17047);
or U18065 (N_18065,N_17338,N_17090);
xor U18066 (N_18066,N_17055,N_17199);
or U18067 (N_18067,N_17324,N_17304);
nand U18068 (N_18068,N_17335,N_17213);
xor U18069 (N_18069,N_17591,N_17228);
xnor U18070 (N_18070,N_17222,N_17164);
xnor U18071 (N_18071,N_17295,N_17718);
xor U18072 (N_18072,N_17419,N_17549);
or U18073 (N_18073,N_17416,N_17325);
nor U18074 (N_18074,N_17502,N_17410);
and U18075 (N_18075,N_17271,N_17243);
nand U18076 (N_18076,N_17112,N_17776);
and U18077 (N_18077,N_17711,N_17545);
nor U18078 (N_18078,N_17713,N_17472);
or U18079 (N_18079,N_17281,N_17471);
or U18080 (N_18080,N_17063,N_17647);
nand U18081 (N_18081,N_17420,N_17693);
nand U18082 (N_18082,N_17028,N_17942);
and U18083 (N_18083,N_17110,N_17932);
nand U18084 (N_18084,N_17292,N_17329);
or U18085 (N_18085,N_17601,N_17596);
or U18086 (N_18086,N_17474,N_17945);
and U18087 (N_18087,N_17754,N_17991);
nand U18088 (N_18088,N_17949,N_17412);
nand U18089 (N_18089,N_17639,N_17302);
and U18090 (N_18090,N_17106,N_17019);
xor U18091 (N_18091,N_17427,N_17689);
nor U18092 (N_18092,N_17026,N_17848);
nand U18093 (N_18093,N_17202,N_17499);
or U18094 (N_18094,N_17838,N_17859);
xor U18095 (N_18095,N_17389,N_17986);
xnor U18096 (N_18096,N_17892,N_17742);
nor U18097 (N_18097,N_17748,N_17797);
or U18098 (N_18098,N_17969,N_17216);
nor U18099 (N_18099,N_17714,N_17170);
nor U18100 (N_18100,N_17645,N_17947);
nand U18101 (N_18101,N_17840,N_17688);
nand U18102 (N_18102,N_17725,N_17539);
xnor U18103 (N_18103,N_17478,N_17436);
xnor U18104 (N_18104,N_17344,N_17421);
or U18105 (N_18105,N_17924,N_17886);
xnor U18106 (N_18106,N_17721,N_17306);
xnor U18107 (N_18107,N_17697,N_17223);
or U18108 (N_18108,N_17978,N_17444);
nand U18109 (N_18109,N_17383,N_17893);
nor U18110 (N_18110,N_17824,N_17629);
and U18111 (N_18111,N_17230,N_17259);
nor U18112 (N_18112,N_17896,N_17321);
or U18113 (N_18113,N_17066,N_17121);
xnor U18114 (N_18114,N_17434,N_17274);
xnor U18115 (N_18115,N_17015,N_17835);
nor U18116 (N_18116,N_17229,N_17882);
xnor U18117 (N_18117,N_17240,N_17611);
and U18118 (N_18118,N_17560,N_17148);
nand U18119 (N_18119,N_17804,N_17273);
nand U18120 (N_18120,N_17384,N_17569);
or U18121 (N_18121,N_17204,N_17819);
nand U18122 (N_18122,N_17709,N_17674);
and U18123 (N_18123,N_17732,N_17373);
or U18124 (N_18124,N_17578,N_17371);
nand U18125 (N_18125,N_17235,N_17141);
xnor U18126 (N_18126,N_17209,N_17875);
xnor U18127 (N_18127,N_17686,N_17534);
nor U18128 (N_18128,N_17481,N_17154);
or U18129 (N_18129,N_17849,N_17084);
xnor U18130 (N_18130,N_17088,N_17326);
or U18131 (N_18131,N_17755,N_17435);
and U18132 (N_18132,N_17512,N_17334);
nor U18133 (N_18133,N_17907,N_17175);
xor U18134 (N_18134,N_17812,N_17571);
nor U18135 (N_18135,N_17930,N_17514);
nor U18136 (N_18136,N_17786,N_17577);
nand U18137 (N_18137,N_17146,N_17117);
xnor U18138 (N_18138,N_17491,N_17670);
xor U18139 (N_18139,N_17699,N_17162);
nand U18140 (N_18140,N_17360,N_17964);
xnor U18141 (N_18141,N_17065,N_17150);
nand U18142 (N_18142,N_17814,N_17604);
xor U18143 (N_18143,N_17618,N_17729);
xor U18144 (N_18144,N_17309,N_17249);
nor U18145 (N_18145,N_17315,N_17929);
and U18146 (N_18146,N_17497,N_17857);
and U18147 (N_18147,N_17861,N_17803);
or U18148 (N_18148,N_17039,N_17264);
nand U18149 (N_18149,N_17704,N_17917);
xnor U18150 (N_18150,N_17186,N_17212);
or U18151 (N_18151,N_17738,N_17739);
nand U18152 (N_18152,N_17980,N_17020);
and U18153 (N_18153,N_17610,N_17939);
xnor U18154 (N_18154,N_17375,N_17388);
nor U18155 (N_18155,N_17505,N_17504);
xnor U18156 (N_18156,N_17897,N_17133);
nor U18157 (N_18157,N_17008,N_17912);
xnor U18158 (N_18158,N_17702,N_17537);
nand U18159 (N_18159,N_17779,N_17692);
or U18160 (N_18160,N_17556,N_17029);
and U18161 (N_18161,N_17094,N_17157);
nor U18162 (N_18162,N_17046,N_17432);
nor U18163 (N_18163,N_17717,N_17548);
and U18164 (N_18164,N_17581,N_17927);
or U18165 (N_18165,N_17147,N_17813);
nor U18166 (N_18166,N_17443,N_17962);
nor U18167 (N_18167,N_17214,N_17177);
and U18168 (N_18168,N_17314,N_17098);
and U18169 (N_18169,N_17789,N_17902);
nor U18170 (N_18170,N_17048,N_17682);
nor U18171 (N_18171,N_17774,N_17706);
and U18172 (N_18172,N_17936,N_17627);
nor U18173 (N_18173,N_17045,N_17270);
nand U18174 (N_18174,N_17946,N_17871);
and U18175 (N_18175,N_17903,N_17183);
and U18176 (N_18176,N_17531,N_17793);
nand U18177 (N_18177,N_17075,N_17428);
nand U18178 (N_18178,N_17854,N_17683);
or U18179 (N_18179,N_17673,N_17938);
nand U18180 (N_18180,N_17817,N_17846);
and U18181 (N_18181,N_17064,N_17994);
xor U18182 (N_18182,N_17114,N_17104);
nor U18183 (N_18183,N_17358,N_17449);
xnor U18184 (N_18184,N_17700,N_17527);
xnor U18185 (N_18185,N_17393,N_17013);
nor U18186 (N_18186,N_17873,N_17874);
nor U18187 (N_18187,N_17836,N_17463);
nand U18188 (N_18188,N_17973,N_17715);
nor U18189 (N_18189,N_17415,N_17832);
nand U18190 (N_18190,N_17036,N_17226);
or U18191 (N_18191,N_17620,N_17784);
nor U18192 (N_18192,N_17349,N_17911);
xnor U18193 (N_18193,N_17862,N_17303);
and U18194 (N_18194,N_17203,N_17669);
nor U18195 (N_18195,N_17042,N_17906);
and U18196 (N_18196,N_17759,N_17285);
xnor U18197 (N_18197,N_17244,N_17944);
nand U18198 (N_18198,N_17086,N_17771);
nor U18199 (N_18199,N_17992,N_17572);
nor U18200 (N_18200,N_17658,N_17659);
xor U18201 (N_18201,N_17441,N_17720);
nand U18202 (N_18202,N_17473,N_17407);
xnor U18203 (N_18203,N_17613,N_17395);
xnor U18204 (N_18204,N_17009,N_17870);
or U18205 (N_18205,N_17559,N_17967);
and U18206 (N_18206,N_17424,N_17447);
and U18207 (N_18207,N_17327,N_17323);
and U18208 (N_18208,N_17595,N_17847);
nand U18209 (N_18209,N_17557,N_17322);
nand U18210 (N_18210,N_17189,N_17958);
or U18211 (N_18211,N_17585,N_17227);
or U18212 (N_18212,N_17455,N_17635);
nand U18213 (N_18213,N_17642,N_17798);
nor U18214 (N_18214,N_17173,N_17417);
or U18215 (N_18215,N_17957,N_17215);
and U18216 (N_18216,N_17777,N_17656);
nand U18217 (N_18217,N_17763,N_17464);
xnor U18218 (N_18218,N_17661,N_17097);
or U18219 (N_18219,N_17542,N_17950);
nor U18220 (N_18220,N_17567,N_17486);
nor U18221 (N_18221,N_17403,N_17095);
nor U18222 (N_18222,N_17864,N_17071);
nor U18223 (N_18223,N_17439,N_17339);
nand U18224 (N_18224,N_17767,N_17564);
or U18225 (N_18225,N_17233,N_17241);
xor U18226 (N_18226,N_17582,N_17663);
nand U18227 (N_18227,N_17990,N_17301);
nand U18228 (N_18228,N_17489,N_17960);
or U18229 (N_18229,N_17268,N_17378);
xor U18230 (N_18230,N_17668,N_17152);
and U18231 (N_18231,N_17877,N_17404);
or U18232 (N_18232,N_17580,N_17644);
nor U18233 (N_18233,N_17607,N_17129);
or U18234 (N_18234,N_17982,N_17895);
nand U18235 (N_18235,N_17551,N_17852);
nand U18236 (N_18236,N_17418,N_17728);
and U18237 (N_18237,N_17820,N_17568);
or U18238 (N_18238,N_17465,N_17746);
or U18239 (N_18239,N_17206,N_17313);
nor U18240 (N_18240,N_17654,N_17032);
nor U18241 (N_18241,N_17054,N_17554);
and U18242 (N_18242,N_17369,N_17562);
xnor U18243 (N_18243,N_17558,N_17758);
or U18244 (N_18244,N_17425,N_17541);
nor U18245 (N_18245,N_17025,N_17575);
and U18246 (N_18246,N_17782,N_17040);
and U18247 (N_18247,N_17188,N_17769);
nand U18248 (N_18248,N_17251,N_17602);
and U18249 (N_18249,N_17130,N_17138);
and U18250 (N_18250,N_17898,N_17480);
or U18251 (N_18251,N_17860,N_17002);
or U18252 (N_18252,N_17081,N_17289);
nor U18253 (N_18253,N_17440,N_17153);
and U18254 (N_18254,N_17523,N_17536);
nand U18255 (N_18255,N_17915,N_17802);
or U18256 (N_18256,N_17479,N_17747);
and U18257 (N_18257,N_17003,N_17070);
xnor U18258 (N_18258,N_17617,N_17555);
nor U18259 (N_18259,N_17400,N_17676);
or U18260 (N_18260,N_17011,N_17853);
and U18261 (N_18261,N_17346,N_17311);
xnor U18262 (N_18262,N_17884,N_17448);
xnor U18263 (N_18263,N_17219,N_17422);
nand U18264 (N_18264,N_17809,N_17307);
xnor U18265 (N_18265,N_17356,N_17999);
or U18266 (N_18266,N_17414,N_17484);
and U18267 (N_18267,N_17855,N_17722);
and U18268 (N_18268,N_17331,N_17856);
xor U18269 (N_18269,N_17143,N_17837);
nand U18270 (N_18270,N_17723,N_17299);
or U18271 (N_18271,N_17059,N_17495);
nand U18272 (N_18272,N_17799,N_17816);
xnor U18273 (N_18273,N_17919,N_17158);
and U18274 (N_18274,N_17593,N_17773);
and U18275 (N_18275,N_17031,N_17910);
and U18276 (N_18276,N_17211,N_17000);
nor U18277 (N_18277,N_17135,N_17194);
nand U18278 (N_18278,N_17476,N_17918);
nand U18279 (N_18279,N_17631,N_17648);
nor U18280 (N_18280,N_17638,N_17057);
and U18281 (N_18281,N_17377,N_17083);
or U18282 (N_18282,N_17966,N_17082);
or U18283 (N_18283,N_17072,N_17408);
or U18284 (N_18284,N_17878,N_17667);
nor U18285 (N_18285,N_17528,N_17801);
nor U18286 (N_18286,N_17120,N_17250);
or U18287 (N_18287,N_17701,N_17885);
nor U18288 (N_18288,N_17858,N_17452);
and U18289 (N_18289,N_17201,N_17600);
nor U18290 (N_18290,N_17968,N_17376);
and U18291 (N_18291,N_17889,N_17665);
or U18292 (N_18292,N_17238,N_17679);
and U18293 (N_18293,N_17312,N_17016);
nand U18294 (N_18294,N_17640,N_17625);
and U18295 (N_18295,N_17257,N_17494);
nand U18296 (N_18296,N_17386,N_17989);
xnor U18297 (N_18297,N_17445,N_17263);
xor U18298 (N_18298,N_17513,N_17056);
and U18299 (N_18299,N_17598,N_17550);
or U18300 (N_18300,N_17650,N_17736);
and U18301 (N_18301,N_17382,N_17995);
nand U18302 (N_18302,N_17363,N_17822);
xor U18303 (N_18303,N_17756,N_17156);
nand U18304 (N_18304,N_17526,N_17051);
xnor U18305 (N_18305,N_17500,N_17664);
and U18306 (N_18306,N_17159,N_17778);
and U18307 (N_18307,N_17954,N_17196);
nor U18308 (N_18308,N_17808,N_17546);
xnor U18309 (N_18309,N_17904,N_17456);
and U18310 (N_18310,N_17905,N_17041);
xnor U18311 (N_18311,N_17492,N_17247);
nor U18312 (N_18312,N_17766,N_17643);
or U18313 (N_18313,N_17296,N_17485);
nand U18314 (N_18314,N_17353,N_17139);
or U18315 (N_18315,N_17879,N_17818);
or U18316 (N_18316,N_17888,N_17566);
or U18317 (N_18317,N_17252,N_17765);
and U18318 (N_18318,N_17624,N_17399);
nand U18319 (N_18319,N_17431,N_17010);
or U18320 (N_18320,N_17851,N_17178);
nand U18321 (N_18321,N_17163,N_17179);
or U18322 (N_18322,N_17165,N_17187);
nand U18323 (N_18323,N_17844,N_17805);
nor U18324 (N_18324,N_17265,N_17811);
nor U18325 (N_18325,N_17828,N_17781);
xor U18326 (N_18326,N_17023,N_17951);
and U18327 (N_18327,N_17843,N_17925);
nand U18328 (N_18328,N_17719,N_17330);
xor U18329 (N_18329,N_17396,N_17182);
and U18330 (N_18330,N_17757,N_17053);
and U18331 (N_18331,N_17696,N_17694);
or U18332 (N_18332,N_17677,N_17641);
nor U18333 (N_18333,N_17791,N_17328);
nor U18334 (N_18334,N_17914,N_17080);
and U18335 (N_18335,N_17959,N_17087);
nor U18336 (N_18336,N_17615,N_17197);
nor U18337 (N_18337,N_17745,N_17744);
or U18338 (N_18338,N_17190,N_17181);
nand U18339 (N_18339,N_17894,N_17921);
xnor U18340 (N_18340,N_17457,N_17933);
and U18341 (N_18341,N_17195,N_17359);
and U18342 (N_18342,N_17775,N_17787);
or U18343 (N_18343,N_17128,N_17207);
nor U18344 (N_18344,N_17050,N_17269);
or U18345 (N_18345,N_17381,N_17300);
nand U18346 (N_18346,N_17681,N_17626);
nand U18347 (N_18347,N_17690,N_17519);
nand U18348 (N_18348,N_17628,N_17038);
nor U18349 (N_18349,N_17357,N_17260);
nand U18350 (N_18350,N_17167,N_17532);
nor U18351 (N_18351,N_17374,N_17880);
xor U18352 (N_18352,N_17971,N_17069);
xnor U18353 (N_18353,N_17573,N_17733);
xnor U18354 (N_18354,N_17176,N_17594);
or U18355 (N_18355,N_17272,N_17956);
and U18356 (N_18356,N_17928,N_17621);
or U18357 (N_18357,N_17174,N_17872);
xnor U18358 (N_18358,N_17398,N_17831);
xnor U18359 (N_18359,N_17563,N_17671);
nand U18360 (N_18360,N_17469,N_17490);
or U18361 (N_18361,N_17483,N_17948);
nand U18362 (N_18362,N_17698,N_17337);
nand U18363 (N_18363,N_17565,N_17883);
and U18364 (N_18364,N_17185,N_17783);
xnor U18365 (N_18365,N_17772,N_17678);
or U18366 (N_18366,N_17390,N_17401);
xor U18367 (N_18367,N_17751,N_17614);
nand U18368 (N_18368,N_17365,N_17780);
and U18369 (N_18369,N_17332,N_17623);
xnor U18370 (N_18370,N_17825,N_17101);
or U18371 (N_18371,N_17409,N_17792);
xnor U18372 (N_18372,N_17934,N_17810);
nor U18373 (N_18373,N_17017,N_17865);
nand U18374 (N_18374,N_17518,N_17517);
or U18375 (N_18375,N_17450,N_17675);
nor U18376 (N_18376,N_17587,N_17429);
xor U18377 (N_18377,N_17169,N_17392);
xnor U18378 (N_18378,N_17459,N_17030);
nand U18379 (N_18379,N_17118,N_17397);
nand U18380 (N_18380,N_17891,N_17402);
or U18381 (N_18381,N_17367,N_17493);
xor U18382 (N_18382,N_17926,N_17796);
nor U18383 (N_18383,N_17524,N_17462);
nor U18384 (N_18384,N_17943,N_17119);
xnor U18385 (N_18385,N_17496,N_17508);
xnor U18386 (N_18386,N_17262,N_17426);
nand U18387 (N_18387,N_17609,N_17916);
nand U18388 (N_18388,N_17379,N_17616);
or U18389 (N_18389,N_17411,N_17149);
xor U18390 (N_18390,N_17279,N_17806);
or U18391 (N_18391,N_17380,N_17850);
and U18392 (N_18392,N_17649,N_17705);
or U18393 (N_18393,N_17795,N_17109);
and U18394 (N_18394,N_17466,N_17961);
nand U18395 (N_18395,N_17085,N_17975);
nor U18396 (N_18396,N_17078,N_17276);
xor U18397 (N_18397,N_17515,N_17287);
nand U18398 (N_18398,N_17845,N_17953);
nor U18399 (N_18399,N_17612,N_17770);
or U18400 (N_18400,N_17107,N_17245);
nand U18401 (N_18401,N_17881,N_17437);
or U18402 (N_18402,N_17506,N_17922);
and U18403 (N_18403,N_17073,N_17487);
or U18404 (N_18404,N_17530,N_17703);
nor U18405 (N_18405,N_17239,N_17762);
nor U18406 (N_18406,N_17184,N_17060);
nor U18407 (N_18407,N_17091,N_17869);
nand U18408 (N_18408,N_17205,N_17666);
nand U18409 (N_18409,N_17655,N_17868);
or U18410 (N_18410,N_17021,N_17433);
and U18411 (N_18411,N_17333,N_17052);
nand U18412 (N_18412,N_17815,N_17256);
or U18413 (N_18413,N_17841,N_17752);
and U18414 (N_18414,N_17785,N_17685);
xor U18415 (N_18415,N_17632,N_17972);
or U18416 (N_18416,N_17761,N_17543);
xor U18417 (N_18417,N_17027,N_17935);
and U18418 (N_18418,N_17863,N_17308);
nor U18419 (N_18419,N_17267,N_17901);
xnor U18420 (N_18420,N_17920,N_17867);
xnor U18421 (N_18421,N_17993,N_17242);
xnor U18422 (N_18422,N_17225,N_17192);
or U18423 (N_18423,N_17727,N_17347);
and U18424 (N_18424,N_17908,N_17716);
and U18425 (N_18425,N_17001,N_17984);
and U18426 (N_18426,N_17004,N_17366);
nand U18427 (N_18427,N_17405,N_17255);
and U18428 (N_18428,N_17684,N_17317);
and U18429 (N_18429,N_17501,N_17451);
and U18430 (N_18430,N_17955,N_17364);
nand U18431 (N_18431,N_17544,N_17461);
nand U18432 (N_18432,N_17123,N_17105);
xor U18433 (N_18433,N_17297,N_17160);
and U18434 (N_18434,N_17589,N_17103);
and U18435 (N_18435,N_17310,N_17583);
nor U18436 (N_18436,N_17076,N_17232);
and U18437 (N_18437,N_17981,N_17890);
and U18438 (N_18438,N_17168,N_17253);
and U18439 (N_18439,N_17423,N_17277);
xor U18440 (N_18440,N_17753,N_17286);
nand U18441 (N_18441,N_17482,N_17937);
and U18442 (N_18442,N_17092,N_17707);
nand U18443 (N_18443,N_17406,N_17750);
xor U18444 (N_18444,N_17368,N_17234);
nor U18445 (N_18445,N_17191,N_17987);
nor U18446 (N_18446,N_17899,N_17018);
nand U18447 (N_18447,N_17807,N_17533);
nand U18448 (N_18448,N_17740,N_17525);
nor U18449 (N_18449,N_17603,N_17134);
nor U18450 (N_18450,N_17458,N_17619);
or U18451 (N_18451,N_17608,N_17093);
nor U18452 (N_18452,N_17293,N_17737);
xor U18453 (N_18453,N_17166,N_17597);
nor U18454 (N_18454,N_17180,N_17997);
nand U18455 (N_18455,N_17254,N_17278);
or U18456 (N_18456,N_17584,N_17979);
xor U18457 (N_18457,N_17061,N_17827);
xnor U18458 (N_18458,N_17198,N_17503);
and U18459 (N_18459,N_17132,N_17547);
xor U18460 (N_18460,N_17913,N_17931);
nand U18461 (N_18461,N_17974,N_17522);
nor U18462 (N_18462,N_17712,N_17099);
nor U18463 (N_18463,N_17319,N_17909);
or U18464 (N_18464,N_17963,N_17126);
nor U18465 (N_18465,N_17579,N_17826);
nor U18466 (N_18466,N_17687,N_17352);
nor U18467 (N_18467,N_17136,N_17866);
nor U18468 (N_18468,N_17976,N_17345);
and U18469 (N_18469,N_17236,N_17708);
and U18470 (N_18470,N_17122,N_17876);
nand U18471 (N_18471,N_17430,N_17680);
or U18472 (N_18472,N_17535,N_17996);
and U18473 (N_18473,N_17952,N_17142);
nand U18474 (N_18474,N_17224,N_17391);
or U18475 (N_18475,N_17794,N_17387);
or U18476 (N_18476,N_17210,N_17662);
xor U18477 (N_18477,N_17839,N_17280);
nand U18478 (N_18478,N_17691,N_17442);
nor U18479 (N_18479,N_17634,N_17068);
nand U18480 (N_18480,N_17467,N_17145);
nor U18481 (N_18481,N_17574,N_17284);
and U18482 (N_18482,N_17470,N_17161);
xor U18483 (N_18483,N_17290,N_17726);
xor U18484 (N_18484,N_17151,N_17510);
xnor U18485 (N_18485,N_17318,N_17394);
or U18486 (N_18486,N_17044,N_17468);
nand U18487 (N_18487,N_17538,N_17672);
nand U18488 (N_18488,N_17599,N_17172);
nand U18489 (N_18489,N_17475,N_17760);
nor U18490 (N_18490,N_17576,N_17316);
nor U18491 (N_18491,N_17446,N_17529);
xor U18492 (N_18492,N_17731,N_17829);
nor U18493 (N_18493,N_17590,N_17637);
nor U18494 (N_18494,N_17940,N_17588);
and U18495 (N_18495,N_17834,N_17509);
or U18496 (N_18496,N_17171,N_17842);
xnor U18497 (N_18497,N_17033,N_17043);
or U18498 (N_18498,N_17096,N_17998);
and U18499 (N_18499,N_17586,N_17341);
nor U18500 (N_18500,N_17830,N_17988);
xnor U18501 (N_18501,N_17771,N_17977);
nand U18502 (N_18502,N_17467,N_17591);
or U18503 (N_18503,N_17950,N_17332);
and U18504 (N_18504,N_17149,N_17136);
nand U18505 (N_18505,N_17838,N_17315);
nand U18506 (N_18506,N_17276,N_17086);
nor U18507 (N_18507,N_17906,N_17524);
nor U18508 (N_18508,N_17505,N_17953);
or U18509 (N_18509,N_17275,N_17770);
or U18510 (N_18510,N_17060,N_17102);
nand U18511 (N_18511,N_17737,N_17256);
and U18512 (N_18512,N_17822,N_17455);
and U18513 (N_18513,N_17830,N_17266);
xor U18514 (N_18514,N_17351,N_17629);
and U18515 (N_18515,N_17506,N_17211);
and U18516 (N_18516,N_17754,N_17335);
nor U18517 (N_18517,N_17018,N_17399);
or U18518 (N_18518,N_17651,N_17419);
xor U18519 (N_18519,N_17335,N_17729);
xor U18520 (N_18520,N_17446,N_17205);
nand U18521 (N_18521,N_17010,N_17196);
nor U18522 (N_18522,N_17026,N_17623);
or U18523 (N_18523,N_17211,N_17198);
nand U18524 (N_18524,N_17880,N_17915);
and U18525 (N_18525,N_17208,N_17146);
xor U18526 (N_18526,N_17692,N_17725);
and U18527 (N_18527,N_17900,N_17018);
xnor U18528 (N_18528,N_17234,N_17831);
nand U18529 (N_18529,N_17629,N_17126);
and U18530 (N_18530,N_17003,N_17049);
or U18531 (N_18531,N_17450,N_17229);
and U18532 (N_18532,N_17214,N_17791);
nand U18533 (N_18533,N_17189,N_17097);
or U18534 (N_18534,N_17814,N_17495);
and U18535 (N_18535,N_17108,N_17128);
nor U18536 (N_18536,N_17502,N_17375);
and U18537 (N_18537,N_17586,N_17027);
nand U18538 (N_18538,N_17837,N_17533);
or U18539 (N_18539,N_17096,N_17005);
nor U18540 (N_18540,N_17818,N_17180);
and U18541 (N_18541,N_17327,N_17349);
nand U18542 (N_18542,N_17219,N_17623);
xor U18543 (N_18543,N_17691,N_17531);
or U18544 (N_18544,N_17309,N_17215);
and U18545 (N_18545,N_17841,N_17678);
nor U18546 (N_18546,N_17169,N_17140);
nor U18547 (N_18547,N_17962,N_17005);
or U18548 (N_18548,N_17486,N_17879);
or U18549 (N_18549,N_17279,N_17437);
and U18550 (N_18550,N_17836,N_17002);
nor U18551 (N_18551,N_17468,N_17419);
nor U18552 (N_18552,N_17541,N_17996);
nor U18553 (N_18553,N_17950,N_17536);
nand U18554 (N_18554,N_17937,N_17133);
nor U18555 (N_18555,N_17074,N_17854);
xor U18556 (N_18556,N_17726,N_17216);
xor U18557 (N_18557,N_17803,N_17771);
nand U18558 (N_18558,N_17667,N_17274);
xnor U18559 (N_18559,N_17102,N_17124);
xor U18560 (N_18560,N_17010,N_17715);
xor U18561 (N_18561,N_17866,N_17778);
nor U18562 (N_18562,N_17065,N_17280);
nand U18563 (N_18563,N_17499,N_17067);
or U18564 (N_18564,N_17484,N_17346);
and U18565 (N_18565,N_17183,N_17829);
nand U18566 (N_18566,N_17651,N_17360);
nand U18567 (N_18567,N_17227,N_17170);
nor U18568 (N_18568,N_17450,N_17056);
xnor U18569 (N_18569,N_17776,N_17342);
or U18570 (N_18570,N_17500,N_17132);
or U18571 (N_18571,N_17158,N_17007);
nand U18572 (N_18572,N_17773,N_17883);
nor U18573 (N_18573,N_17914,N_17443);
nand U18574 (N_18574,N_17032,N_17749);
and U18575 (N_18575,N_17483,N_17681);
nand U18576 (N_18576,N_17653,N_17815);
nor U18577 (N_18577,N_17476,N_17270);
nand U18578 (N_18578,N_17512,N_17388);
nand U18579 (N_18579,N_17403,N_17508);
xor U18580 (N_18580,N_17698,N_17603);
nor U18581 (N_18581,N_17166,N_17561);
nand U18582 (N_18582,N_17342,N_17389);
and U18583 (N_18583,N_17549,N_17196);
nor U18584 (N_18584,N_17926,N_17285);
nand U18585 (N_18585,N_17110,N_17054);
nand U18586 (N_18586,N_17116,N_17737);
nand U18587 (N_18587,N_17649,N_17708);
and U18588 (N_18588,N_17441,N_17236);
and U18589 (N_18589,N_17106,N_17055);
and U18590 (N_18590,N_17965,N_17006);
and U18591 (N_18591,N_17475,N_17828);
nand U18592 (N_18592,N_17601,N_17916);
or U18593 (N_18593,N_17892,N_17442);
nor U18594 (N_18594,N_17221,N_17737);
nand U18595 (N_18595,N_17442,N_17830);
and U18596 (N_18596,N_17150,N_17488);
nand U18597 (N_18597,N_17038,N_17534);
xnor U18598 (N_18598,N_17692,N_17574);
nor U18599 (N_18599,N_17129,N_17841);
nand U18600 (N_18600,N_17207,N_17936);
or U18601 (N_18601,N_17744,N_17021);
and U18602 (N_18602,N_17064,N_17612);
xor U18603 (N_18603,N_17809,N_17136);
xnor U18604 (N_18604,N_17309,N_17592);
xnor U18605 (N_18605,N_17048,N_17287);
nor U18606 (N_18606,N_17224,N_17645);
nor U18607 (N_18607,N_17981,N_17345);
or U18608 (N_18608,N_17141,N_17072);
nor U18609 (N_18609,N_17289,N_17469);
and U18610 (N_18610,N_17280,N_17087);
or U18611 (N_18611,N_17411,N_17105);
or U18612 (N_18612,N_17182,N_17521);
nand U18613 (N_18613,N_17652,N_17033);
nor U18614 (N_18614,N_17718,N_17937);
and U18615 (N_18615,N_17289,N_17327);
xnor U18616 (N_18616,N_17367,N_17052);
nand U18617 (N_18617,N_17075,N_17542);
nor U18618 (N_18618,N_17915,N_17709);
and U18619 (N_18619,N_17991,N_17606);
xnor U18620 (N_18620,N_17225,N_17113);
nor U18621 (N_18621,N_17845,N_17789);
xor U18622 (N_18622,N_17606,N_17212);
nor U18623 (N_18623,N_17341,N_17572);
nand U18624 (N_18624,N_17903,N_17812);
nand U18625 (N_18625,N_17320,N_17754);
nand U18626 (N_18626,N_17899,N_17655);
nor U18627 (N_18627,N_17762,N_17411);
nor U18628 (N_18628,N_17208,N_17855);
and U18629 (N_18629,N_17218,N_17496);
nor U18630 (N_18630,N_17683,N_17965);
nand U18631 (N_18631,N_17893,N_17878);
xnor U18632 (N_18632,N_17334,N_17449);
xnor U18633 (N_18633,N_17530,N_17904);
and U18634 (N_18634,N_17378,N_17984);
and U18635 (N_18635,N_17619,N_17648);
and U18636 (N_18636,N_17245,N_17362);
xor U18637 (N_18637,N_17224,N_17092);
or U18638 (N_18638,N_17826,N_17974);
or U18639 (N_18639,N_17884,N_17569);
nand U18640 (N_18640,N_17032,N_17622);
nand U18641 (N_18641,N_17174,N_17010);
xor U18642 (N_18642,N_17867,N_17433);
or U18643 (N_18643,N_17573,N_17210);
nand U18644 (N_18644,N_17712,N_17206);
xor U18645 (N_18645,N_17156,N_17762);
nor U18646 (N_18646,N_17266,N_17446);
and U18647 (N_18647,N_17555,N_17861);
nand U18648 (N_18648,N_17480,N_17458);
nand U18649 (N_18649,N_17813,N_17255);
nor U18650 (N_18650,N_17584,N_17102);
nor U18651 (N_18651,N_17125,N_17118);
and U18652 (N_18652,N_17487,N_17799);
xnor U18653 (N_18653,N_17638,N_17840);
xor U18654 (N_18654,N_17245,N_17274);
nand U18655 (N_18655,N_17773,N_17993);
nor U18656 (N_18656,N_17782,N_17801);
and U18657 (N_18657,N_17830,N_17236);
nor U18658 (N_18658,N_17056,N_17856);
xnor U18659 (N_18659,N_17866,N_17526);
nand U18660 (N_18660,N_17308,N_17517);
nor U18661 (N_18661,N_17579,N_17854);
and U18662 (N_18662,N_17707,N_17785);
or U18663 (N_18663,N_17533,N_17121);
and U18664 (N_18664,N_17733,N_17221);
and U18665 (N_18665,N_17936,N_17821);
nand U18666 (N_18666,N_17423,N_17188);
xnor U18667 (N_18667,N_17249,N_17944);
or U18668 (N_18668,N_17952,N_17446);
nor U18669 (N_18669,N_17564,N_17252);
or U18670 (N_18670,N_17581,N_17422);
nor U18671 (N_18671,N_17424,N_17394);
nor U18672 (N_18672,N_17349,N_17753);
nor U18673 (N_18673,N_17895,N_17584);
and U18674 (N_18674,N_17257,N_17118);
nand U18675 (N_18675,N_17557,N_17559);
nor U18676 (N_18676,N_17353,N_17439);
or U18677 (N_18677,N_17186,N_17264);
xnor U18678 (N_18678,N_17897,N_17851);
or U18679 (N_18679,N_17771,N_17217);
nor U18680 (N_18680,N_17831,N_17432);
nand U18681 (N_18681,N_17866,N_17312);
and U18682 (N_18682,N_17425,N_17590);
nor U18683 (N_18683,N_17786,N_17653);
or U18684 (N_18684,N_17446,N_17944);
or U18685 (N_18685,N_17352,N_17237);
nor U18686 (N_18686,N_17265,N_17872);
or U18687 (N_18687,N_17855,N_17162);
nor U18688 (N_18688,N_17050,N_17275);
and U18689 (N_18689,N_17033,N_17167);
xnor U18690 (N_18690,N_17391,N_17596);
xor U18691 (N_18691,N_17241,N_17450);
nor U18692 (N_18692,N_17620,N_17824);
or U18693 (N_18693,N_17270,N_17325);
or U18694 (N_18694,N_17200,N_17457);
or U18695 (N_18695,N_17258,N_17394);
xnor U18696 (N_18696,N_17155,N_17546);
and U18697 (N_18697,N_17059,N_17904);
xor U18698 (N_18698,N_17532,N_17781);
or U18699 (N_18699,N_17563,N_17404);
or U18700 (N_18700,N_17257,N_17469);
nand U18701 (N_18701,N_17338,N_17346);
xnor U18702 (N_18702,N_17410,N_17927);
nand U18703 (N_18703,N_17791,N_17577);
nor U18704 (N_18704,N_17357,N_17818);
nor U18705 (N_18705,N_17245,N_17184);
and U18706 (N_18706,N_17469,N_17958);
nand U18707 (N_18707,N_17288,N_17891);
nor U18708 (N_18708,N_17604,N_17350);
nand U18709 (N_18709,N_17672,N_17770);
nand U18710 (N_18710,N_17621,N_17271);
nor U18711 (N_18711,N_17001,N_17736);
nand U18712 (N_18712,N_17452,N_17499);
and U18713 (N_18713,N_17233,N_17968);
nor U18714 (N_18714,N_17822,N_17020);
nand U18715 (N_18715,N_17116,N_17128);
or U18716 (N_18716,N_17963,N_17961);
nor U18717 (N_18717,N_17530,N_17080);
xor U18718 (N_18718,N_17332,N_17057);
and U18719 (N_18719,N_17166,N_17488);
xor U18720 (N_18720,N_17700,N_17913);
and U18721 (N_18721,N_17323,N_17517);
nand U18722 (N_18722,N_17760,N_17243);
nor U18723 (N_18723,N_17354,N_17855);
or U18724 (N_18724,N_17767,N_17443);
nand U18725 (N_18725,N_17019,N_17483);
and U18726 (N_18726,N_17536,N_17208);
xnor U18727 (N_18727,N_17481,N_17496);
and U18728 (N_18728,N_17829,N_17757);
xnor U18729 (N_18729,N_17183,N_17707);
nand U18730 (N_18730,N_17273,N_17543);
or U18731 (N_18731,N_17916,N_17682);
nor U18732 (N_18732,N_17378,N_17552);
nand U18733 (N_18733,N_17833,N_17377);
nor U18734 (N_18734,N_17203,N_17072);
or U18735 (N_18735,N_17747,N_17699);
or U18736 (N_18736,N_17037,N_17077);
and U18737 (N_18737,N_17075,N_17298);
or U18738 (N_18738,N_17976,N_17824);
nor U18739 (N_18739,N_17985,N_17111);
nand U18740 (N_18740,N_17146,N_17749);
xor U18741 (N_18741,N_17184,N_17423);
nand U18742 (N_18742,N_17603,N_17352);
xnor U18743 (N_18743,N_17344,N_17157);
nand U18744 (N_18744,N_17714,N_17431);
nor U18745 (N_18745,N_17352,N_17711);
or U18746 (N_18746,N_17411,N_17542);
or U18747 (N_18747,N_17963,N_17575);
nor U18748 (N_18748,N_17337,N_17248);
nor U18749 (N_18749,N_17012,N_17919);
and U18750 (N_18750,N_17235,N_17481);
xnor U18751 (N_18751,N_17163,N_17290);
xnor U18752 (N_18752,N_17106,N_17763);
nand U18753 (N_18753,N_17895,N_17237);
nand U18754 (N_18754,N_17397,N_17998);
nand U18755 (N_18755,N_17082,N_17580);
or U18756 (N_18756,N_17074,N_17033);
xor U18757 (N_18757,N_17699,N_17531);
and U18758 (N_18758,N_17790,N_17431);
and U18759 (N_18759,N_17594,N_17268);
nor U18760 (N_18760,N_17285,N_17305);
and U18761 (N_18761,N_17876,N_17314);
nor U18762 (N_18762,N_17305,N_17297);
nand U18763 (N_18763,N_17007,N_17778);
nand U18764 (N_18764,N_17570,N_17459);
xnor U18765 (N_18765,N_17618,N_17004);
or U18766 (N_18766,N_17813,N_17710);
nand U18767 (N_18767,N_17246,N_17292);
nor U18768 (N_18768,N_17919,N_17257);
or U18769 (N_18769,N_17664,N_17062);
or U18770 (N_18770,N_17331,N_17869);
xor U18771 (N_18771,N_17853,N_17052);
and U18772 (N_18772,N_17413,N_17044);
nand U18773 (N_18773,N_17948,N_17473);
and U18774 (N_18774,N_17382,N_17558);
and U18775 (N_18775,N_17527,N_17837);
and U18776 (N_18776,N_17494,N_17442);
or U18777 (N_18777,N_17047,N_17214);
nand U18778 (N_18778,N_17967,N_17844);
nand U18779 (N_18779,N_17605,N_17275);
or U18780 (N_18780,N_17637,N_17140);
nand U18781 (N_18781,N_17731,N_17283);
nor U18782 (N_18782,N_17550,N_17022);
or U18783 (N_18783,N_17930,N_17298);
nand U18784 (N_18784,N_17054,N_17359);
nand U18785 (N_18785,N_17587,N_17955);
xnor U18786 (N_18786,N_17022,N_17158);
nand U18787 (N_18787,N_17901,N_17194);
and U18788 (N_18788,N_17064,N_17079);
and U18789 (N_18789,N_17807,N_17693);
nand U18790 (N_18790,N_17088,N_17978);
or U18791 (N_18791,N_17430,N_17615);
and U18792 (N_18792,N_17841,N_17627);
xnor U18793 (N_18793,N_17982,N_17523);
nor U18794 (N_18794,N_17334,N_17811);
nand U18795 (N_18795,N_17905,N_17885);
nand U18796 (N_18796,N_17147,N_17444);
xor U18797 (N_18797,N_17713,N_17477);
and U18798 (N_18798,N_17038,N_17153);
nand U18799 (N_18799,N_17318,N_17988);
or U18800 (N_18800,N_17939,N_17053);
or U18801 (N_18801,N_17122,N_17724);
and U18802 (N_18802,N_17090,N_17862);
nor U18803 (N_18803,N_17666,N_17923);
or U18804 (N_18804,N_17772,N_17981);
and U18805 (N_18805,N_17059,N_17108);
nand U18806 (N_18806,N_17572,N_17478);
nand U18807 (N_18807,N_17726,N_17810);
nor U18808 (N_18808,N_17945,N_17691);
and U18809 (N_18809,N_17285,N_17398);
or U18810 (N_18810,N_17501,N_17439);
xnor U18811 (N_18811,N_17733,N_17249);
or U18812 (N_18812,N_17913,N_17782);
xnor U18813 (N_18813,N_17172,N_17427);
nor U18814 (N_18814,N_17551,N_17579);
nand U18815 (N_18815,N_17646,N_17453);
nand U18816 (N_18816,N_17084,N_17461);
nor U18817 (N_18817,N_17804,N_17802);
and U18818 (N_18818,N_17954,N_17031);
nand U18819 (N_18819,N_17287,N_17289);
nand U18820 (N_18820,N_17827,N_17870);
or U18821 (N_18821,N_17879,N_17567);
and U18822 (N_18822,N_17153,N_17574);
and U18823 (N_18823,N_17809,N_17677);
nand U18824 (N_18824,N_17259,N_17165);
or U18825 (N_18825,N_17914,N_17536);
nor U18826 (N_18826,N_17980,N_17817);
nand U18827 (N_18827,N_17940,N_17718);
and U18828 (N_18828,N_17740,N_17179);
nor U18829 (N_18829,N_17348,N_17791);
xnor U18830 (N_18830,N_17271,N_17463);
nor U18831 (N_18831,N_17561,N_17222);
xnor U18832 (N_18832,N_17884,N_17101);
and U18833 (N_18833,N_17877,N_17136);
nor U18834 (N_18834,N_17639,N_17802);
nor U18835 (N_18835,N_17954,N_17913);
nor U18836 (N_18836,N_17397,N_17918);
nor U18837 (N_18837,N_17898,N_17539);
and U18838 (N_18838,N_17064,N_17418);
and U18839 (N_18839,N_17251,N_17183);
xor U18840 (N_18840,N_17390,N_17035);
xor U18841 (N_18841,N_17664,N_17310);
or U18842 (N_18842,N_17923,N_17091);
and U18843 (N_18843,N_17244,N_17489);
nor U18844 (N_18844,N_17025,N_17820);
xnor U18845 (N_18845,N_17572,N_17385);
xor U18846 (N_18846,N_17557,N_17062);
nand U18847 (N_18847,N_17713,N_17061);
nand U18848 (N_18848,N_17105,N_17460);
and U18849 (N_18849,N_17408,N_17959);
and U18850 (N_18850,N_17894,N_17509);
xor U18851 (N_18851,N_17698,N_17656);
and U18852 (N_18852,N_17887,N_17470);
nand U18853 (N_18853,N_17361,N_17555);
nor U18854 (N_18854,N_17135,N_17482);
and U18855 (N_18855,N_17015,N_17237);
or U18856 (N_18856,N_17662,N_17150);
nand U18857 (N_18857,N_17301,N_17006);
nor U18858 (N_18858,N_17759,N_17580);
xor U18859 (N_18859,N_17568,N_17171);
or U18860 (N_18860,N_17006,N_17028);
or U18861 (N_18861,N_17516,N_17623);
nor U18862 (N_18862,N_17042,N_17049);
nand U18863 (N_18863,N_17046,N_17303);
nand U18864 (N_18864,N_17344,N_17226);
nor U18865 (N_18865,N_17312,N_17764);
and U18866 (N_18866,N_17825,N_17759);
nor U18867 (N_18867,N_17202,N_17698);
and U18868 (N_18868,N_17681,N_17412);
and U18869 (N_18869,N_17810,N_17146);
nor U18870 (N_18870,N_17246,N_17868);
nand U18871 (N_18871,N_17108,N_17783);
and U18872 (N_18872,N_17999,N_17488);
xnor U18873 (N_18873,N_17817,N_17765);
or U18874 (N_18874,N_17739,N_17236);
and U18875 (N_18875,N_17885,N_17801);
nor U18876 (N_18876,N_17412,N_17436);
or U18877 (N_18877,N_17923,N_17187);
nor U18878 (N_18878,N_17009,N_17828);
nand U18879 (N_18879,N_17114,N_17504);
nor U18880 (N_18880,N_17639,N_17512);
and U18881 (N_18881,N_17104,N_17374);
xnor U18882 (N_18882,N_17909,N_17756);
nand U18883 (N_18883,N_17567,N_17611);
xor U18884 (N_18884,N_17848,N_17609);
or U18885 (N_18885,N_17789,N_17884);
xnor U18886 (N_18886,N_17370,N_17033);
and U18887 (N_18887,N_17569,N_17090);
and U18888 (N_18888,N_17090,N_17335);
nand U18889 (N_18889,N_17017,N_17293);
nor U18890 (N_18890,N_17006,N_17235);
and U18891 (N_18891,N_17442,N_17374);
or U18892 (N_18892,N_17169,N_17754);
nor U18893 (N_18893,N_17283,N_17023);
and U18894 (N_18894,N_17002,N_17291);
or U18895 (N_18895,N_17934,N_17076);
nor U18896 (N_18896,N_17071,N_17944);
or U18897 (N_18897,N_17934,N_17888);
nor U18898 (N_18898,N_17663,N_17859);
xor U18899 (N_18899,N_17868,N_17729);
nor U18900 (N_18900,N_17349,N_17547);
xnor U18901 (N_18901,N_17282,N_17340);
xnor U18902 (N_18902,N_17654,N_17850);
nand U18903 (N_18903,N_17107,N_17509);
xor U18904 (N_18904,N_17048,N_17662);
xor U18905 (N_18905,N_17979,N_17603);
xor U18906 (N_18906,N_17190,N_17809);
or U18907 (N_18907,N_17734,N_17110);
nor U18908 (N_18908,N_17220,N_17667);
xnor U18909 (N_18909,N_17271,N_17581);
nand U18910 (N_18910,N_17257,N_17365);
and U18911 (N_18911,N_17818,N_17542);
or U18912 (N_18912,N_17209,N_17836);
xor U18913 (N_18913,N_17192,N_17830);
nor U18914 (N_18914,N_17019,N_17484);
or U18915 (N_18915,N_17628,N_17596);
nand U18916 (N_18916,N_17416,N_17674);
nand U18917 (N_18917,N_17027,N_17213);
nor U18918 (N_18918,N_17982,N_17864);
nand U18919 (N_18919,N_17805,N_17109);
xor U18920 (N_18920,N_17703,N_17577);
nor U18921 (N_18921,N_17678,N_17116);
xnor U18922 (N_18922,N_17935,N_17129);
nor U18923 (N_18923,N_17777,N_17658);
nor U18924 (N_18924,N_17210,N_17780);
xnor U18925 (N_18925,N_17714,N_17814);
or U18926 (N_18926,N_17260,N_17196);
nor U18927 (N_18927,N_17608,N_17464);
nand U18928 (N_18928,N_17465,N_17066);
nor U18929 (N_18929,N_17804,N_17174);
or U18930 (N_18930,N_17196,N_17308);
nor U18931 (N_18931,N_17162,N_17603);
or U18932 (N_18932,N_17583,N_17917);
xor U18933 (N_18933,N_17367,N_17599);
xor U18934 (N_18934,N_17292,N_17021);
or U18935 (N_18935,N_17143,N_17116);
nor U18936 (N_18936,N_17897,N_17217);
or U18937 (N_18937,N_17223,N_17256);
and U18938 (N_18938,N_17862,N_17951);
nor U18939 (N_18939,N_17086,N_17884);
and U18940 (N_18940,N_17683,N_17292);
and U18941 (N_18941,N_17495,N_17320);
and U18942 (N_18942,N_17447,N_17847);
nor U18943 (N_18943,N_17985,N_17104);
nor U18944 (N_18944,N_17948,N_17165);
xnor U18945 (N_18945,N_17904,N_17241);
nor U18946 (N_18946,N_17779,N_17594);
and U18947 (N_18947,N_17319,N_17981);
and U18948 (N_18948,N_17130,N_17614);
nand U18949 (N_18949,N_17694,N_17821);
or U18950 (N_18950,N_17571,N_17017);
or U18951 (N_18951,N_17321,N_17464);
and U18952 (N_18952,N_17758,N_17320);
nor U18953 (N_18953,N_17841,N_17053);
or U18954 (N_18954,N_17895,N_17497);
nand U18955 (N_18955,N_17715,N_17226);
or U18956 (N_18956,N_17246,N_17217);
or U18957 (N_18957,N_17606,N_17805);
and U18958 (N_18958,N_17102,N_17019);
nor U18959 (N_18959,N_17930,N_17751);
or U18960 (N_18960,N_17649,N_17757);
nor U18961 (N_18961,N_17495,N_17371);
xnor U18962 (N_18962,N_17449,N_17437);
xnor U18963 (N_18963,N_17521,N_17825);
nor U18964 (N_18964,N_17765,N_17375);
nor U18965 (N_18965,N_17525,N_17156);
xor U18966 (N_18966,N_17137,N_17442);
and U18967 (N_18967,N_17587,N_17993);
xor U18968 (N_18968,N_17981,N_17847);
or U18969 (N_18969,N_17865,N_17193);
and U18970 (N_18970,N_17489,N_17847);
nand U18971 (N_18971,N_17833,N_17138);
and U18972 (N_18972,N_17266,N_17238);
and U18973 (N_18973,N_17993,N_17356);
xor U18974 (N_18974,N_17474,N_17961);
xor U18975 (N_18975,N_17077,N_17728);
or U18976 (N_18976,N_17292,N_17071);
and U18977 (N_18977,N_17766,N_17052);
or U18978 (N_18978,N_17275,N_17230);
and U18979 (N_18979,N_17608,N_17026);
nor U18980 (N_18980,N_17802,N_17459);
and U18981 (N_18981,N_17377,N_17932);
and U18982 (N_18982,N_17208,N_17293);
and U18983 (N_18983,N_17052,N_17366);
or U18984 (N_18984,N_17613,N_17253);
nor U18985 (N_18985,N_17852,N_17826);
or U18986 (N_18986,N_17429,N_17329);
or U18987 (N_18987,N_17902,N_17920);
nand U18988 (N_18988,N_17001,N_17891);
nand U18989 (N_18989,N_17707,N_17900);
nor U18990 (N_18990,N_17271,N_17563);
and U18991 (N_18991,N_17913,N_17538);
xor U18992 (N_18992,N_17220,N_17457);
or U18993 (N_18993,N_17331,N_17338);
nor U18994 (N_18994,N_17768,N_17765);
xnor U18995 (N_18995,N_17426,N_17122);
nand U18996 (N_18996,N_17594,N_17802);
or U18997 (N_18997,N_17681,N_17553);
or U18998 (N_18998,N_17921,N_17875);
nand U18999 (N_18999,N_17276,N_17785);
and U19000 (N_19000,N_18673,N_18482);
xor U19001 (N_19001,N_18729,N_18273);
xor U19002 (N_19002,N_18466,N_18281);
and U19003 (N_19003,N_18340,N_18839);
nand U19004 (N_19004,N_18980,N_18381);
and U19005 (N_19005,N_18688,N_18593);
nand U19006 (N_19006,N_18266,N_18797);
nor U19007 (N_19007,N_18385,N_18452);
nand U19008 (N_19008,N_18424,N_18081);
xor U19009 (N_19009,N_18988,N_18224);
xor U19010 (N_19010,N_18061,N_18199);
nor U19011 (N_19011,N_18551,N_18989);
nor U19012 (N_19012,N_18763,N_18136);
and U19013 (N_19013,N_18478,N_18389);
nor U19014 (N_19014,N_18781,N_18263);
nand U19015 (N_19015,N_18074,N_18086);
xor U19016 (N_19016,N_18695,N_18615);
nor U19017 (N_19017,N_18993,N_18473);
or U19018 (N_19018,N_18446,N_18701);
nor U19019 (N_19019,N_18543,N_18335);
nand U19020 (N_19020,N_18840,N_18184);
nor U19021 (N_19021,N_18142,N_18139);
xnor U19022 (N_19022,N_18994,N_18612);
or U19023 (N_19023,N_18878,N_18757);
nand U19024 (N_19024,N_18157,N_18745);
xnor U19025 (N_19025,N_18905,N_18349);
nor U19026 (N_19026,N_18454,N_18893);
nand U19027 (N_19027,N_18703,N_18880);
or U19028 (N_19028,N_18087,N_18548);
or U19029 (N_19029,N_18238,N_18949);
or U19030 (N_19030,N_18773,N_18276);
xor U19031 (N_19031,N_18896,N_18176);
or U19032 (N_19032,N_18277,N_18479);
nand U19033 (N_19033,N_18249,N_18736);
nor U19034 (N_19034,N_18258,N_18637);
nor U19035 (N_19035,N_18354,N_18747);
and U19036 (N_19036,N_18068,N_18721);
nand U19037 (N_19037,N_18187,N_18861);
nor U19038 (N_19038,N_18391,N_18941);
and U19039 (N_19039,N_18906,N_18483);
or U19040 (N_19040,N_18304,N_18230);
nand U19041 (N_19041,N_18958,N_18328);
and U19042 (N_19042,N_18293,N_18926);
and U19043 (N_19043,N_18928,N_18241);
nand U19044 (N_19044,N_18642,N_18645);
and U19045 (N_19045,N_18749,N_18559);
xor U19046 (N_19046,N_18170,N_18890);
xnor U19047 (N_19047,N_18754,N_18985);
xor U19048 (N_19048,N_18217,N_18373);
nand U19049 (N_19049,N_18298,N_18716);
xnor U19050 (N_19050,N_18755,N_18674);
xor U19051 (N_19051,N_18843,N_18795);
or U19052 (N_19052,N_18297,N_18892);
nand U19053 (N_19053,N_18966,N_18678);
or U19054 (N_19054,N_18290,N_18041);
xnor U19055 (N_19055,N_18664,N_18095);
nand U19056 (N_19056,N_18540,N_18007);
nor U19057 (N_19057,N_18618,N_18414);
nor U19058 (N_19058,N_18789,N_18022);
xor U19059 (N_19059,N_18455,N_18228);
or U19060 (N_19060,N_18072,N_18753);
or U19061 (N_19061,N_18623,N_18243);
or U19062 (N_19062,N_18393,N_18964);
and U19063 (N_19063,N_18576,N_18937);
and U19064 (N_19064,N_18425,N_18535);
nand U19065 (N_19065,N_18711,N_18047);
xor U19066 (N_19066,N_18215,N_18311);
and U19067 (N_19067,N_18287,N_18338);
nand U19068 (N_19068,N_18271,N_18324);
nor U19069 (N_19069,N_18613,N_18529);
nand U19070 (N_19070,N_18206,N_18846);
and U19071 (N_19071,N_18520,N_18501);
and U19072 (N_19072,N_18185,N_18894);
and U19073 (N_19073,N_18620,N_18648);
nor U19074 (N_19074,N_18734,N_18025);
xor U19075 (N_19075,N_18428,N_18938);
and U19076 (N_19076,N_18411,N_18953);
nand U19077 (N_19077,N_18126,N_18093);
xor U19078 (N_19078,N_18869,N_18852);
xnor U19079 (N_19079,N_18715,N_18141);
or U19080 (N_19080,N_18621,N_18762);
or U19081 (N_19081,N_18550,N_18485);
and U19082 (N_19082,N_18592,N_18499);
nand U19083 (N_19083,N_18200,N_18310);
xnor U19084 (N_19084,N_18440,N_18607);
xnor U19085 (N_19085,N_18223,N_18497);
or U19086 (N_19086,N_18313,N_18983);
and U19087 (N_19087,N_18806,N_18033);
nand U19088 (N_19088,N_18288,N_18788);
and U19089 (N_19089,N_18687,N_18653);
nor U19090 (N_19090,N_18756,N_18252);
or U19091 (N_19091,N_18769,N_18089);
nor U19092 (N_19092,N_18009,N_18114);
nand U19093 (N_19093,N_18805,N_18303);
nor U19094 (N_19094,N_18831,N_18737);
nand U19095 (N_19095,N_18740,N_18524);
and U19096 (N_19096,N_18541,N_18321);
nand U19097 (N_19097,N_18069,N_18608);
or U19098 (N_19098,N_18117,N_18682);
xor U19099 (N_19099,N_18563,N_18132);
or U19100 (N_19100,N_18334,N_18870);
nor U19101 (N_19101,N_18060,N_18475);
xor U19102 (N_19102,N_18987,N_18094);
nand U19103 (N_19103,N_18821,N_18359);
xnor U19104 (N_19104,N_18219,N_18783);
and U19105 (N_19105,N_18034,N_18911);
xnor U19106 (N_19106,N_18873,N_18690);
or U19107 (N_19107,N_18560,N_18636);
and U19108 (N_19108,N_18166,N_18325);
or U19109 (N_19109,N_18662,N_18884);
and U19110 (N_19110,N_18979,N_18946);
or U19111 (N_19111,N_18901,N_18706);
xor U19112 (N_19112,N_18488,N_18188);
xnor U19113 (N_19113,N_18956,N_18037);
nor U19114 (N_19114,N_18426,N_18649);
nand U19115 (N_19115,N_18363,N_18309);
nand U19116 (N_19116,N_18886,N_18810);
xor U19117 (N_19117,N_18793,N_18405);
and U19118 (N_19118,N_18262,N_18766);
or U19119 (N_19119,N_18748,N_18777);
or U19120 (N_19120,N_18380,N_18464);
and U19121 (N_19121,N_18472,N_18545);
or U19122 (N_19122,N_18713,N_18056);
or U19123 (N_19123,N_18169,N_18168);
or U19124 (N_19124,N_18190,N_18511);
and U19125 (N_19125,N_18018,N_18730);
or U19126 (N_19126,N_18704,N_18841);
xnor U19127 (N_19127,N_18237,N_18218);
xnor U19128 (N_19128,N_18598,N_18796);
xnor U19129 (N_19129,N_18016,N_18879);
or U19130 (N_19130,N_18570,N_18400);
xor U19131 (N_19131,N_18194,N_18539);
nor U19132 (N_19132,N_18635,N_18952);
and U19133 (N_19133,N_18855,N_18689);
nand U19134 (N_19134,N_18656,N_18907);
or U19135 (N_19135,N_18165,N_18981);
and U19136 (N_19136,N_18995,N_18633);
xor U19137 (N_19137,N_18547,N_18684);
xnor U19138 (N_19138,N_18948,N_18278);
nor U19139 (N_19139,N_18523,N_18759);
nand U19140 (N_19140,N_18480,N_18883);
and U19141 (N_19141,N_18144,N_18434);
and U19142 (N_19142,N_18161,N_18172);
or U19143 (N_19143,N_18344,N_18566);
nor U19144 (N_19144,N_18897,N_18863);
nor U19145 (N_19145,N_18546,N_18179);
nand U19146 (N_19146,N_18513,N_18449);
or U19147 (N_19147,N_18931,N_18986);
and U19148 (N_19148,N_18407,N_18386);
and U19149 (N_19149,N_18600,N_18315);
and U19150 (N_19150,N_18284,N_18031);
nor U19151 (N_19151,N_18020,N_18395);
xnor U19152 (N_19152,N_18435,N_18666);
or U19153 (N_19153,N_18040,N_18357);
and U19154 (N_19154,N_18229,N_18437);
and U19155 (N_19155,N_18279,N_18629);
or U19156 (N_19156,N_18854,N_18851);
or U19157 (N_19157,N_18105,N_18858);
and U19158 (N_19158,N_18776,N_18671);
nand U19159 (N_19159,N_18201,N_18017);
nor U19160 (N_19160,N_18705,N_18264);
xnor U19161 (N_19161,N_18619,N_18103);
nor U19162 (N_19162,N_18152,N_18580);
xnor U19163 (N_19163,N_18801,N_18991);
and U19164 (N_19164,N_18146,N_18719);
xnor U19165 (N_19165,N_18564,N_18397);
nand U19166 (N_19166,N_18453,N_18787);
or U19167 (N_19167,N_18151,N_18147);
xor U19168 (N_19168,N_18382,N_18680);
or U19169 (N_19169,N_18676,N_18503);
nand U19170 (N_19170,N_18790,N_18046);
and U19171 (N_19171,N_18495,N_18764);
and U19172 (N_19172,N_18235,N_18771);
nand U19173 (N_19173,N_18052,N_18812);
xor U19174 (N_19174,N_18915,N_18871);
and U19175 (N_19175,N_18207,N_18401);
xor U19176 (N_19176,N_18834,N_18646);
and U19177 (N_19177,N_18532,N_18246);
or U19178 (N_19178,N_18491,N_18631);
nand U19179 (N_19179,N_18250,N_18387);
xnor U19180 (N_19180,N_18536,N_18330);
nand U19181 (N_19181,N_18617,N_18461);
and U19182 (N_19182,N_18392,N_18416);
nand U19183 (N_19183,N_18352,N_18417);
and U19184 (N_19184,N_18578,N_18735);
nand U19185 (N_19185,N_18558,N_18700);
nor U19186 (N_19186,N_18679,N_18245);
nand U19187 (N_19187,N_18782,N_18202);
or U19188 (N_19188,N_18794,N_18244);
nand U19189 (N_19189,N_18236,N_18572);
nand U19190 (N_19190,N_18088,N_18112);
nor U19191 (N_19191,N_18289,N_18195);
and U19192 (N_19192,N_18317,N_18167);
xor U19193 (N_19193,N_18082,N_18850);
or U19194 (N_19194,N_18992,N_18542);
and U19195 (N_19195,N_18837,N_18492);
and U19196 (N_19196,N_18128,N_18582);
xnor U19197 (N_19197,N_18413,N_18439);
nor U19198 (N_19198,N_18534,N_18921);
nand U19199 (N_19199,N_18933,N_18127);
xnor U19200 (N_19200,N_18509,N_18376);
nor U19201 (N_19201,N_18832,N_18909);
nand U19202 (N_19202,N_18857,N_18961);
nor U19203 (N_19203,N_18050,N_18396);
nand U19204 (N_19204,N_18875,N_18398);
and U19205 (N_19205,N_18450,N_18902);
xnor U19206 (N_19206,N_18419,N_18922);
nand U19207 (N_19207,N_18800,N_18486);
nor U19208 (N_19208,N_18549,N_18345);
or U19209 (N_19209,N_18573,N_18442);
xor U19210 (N_19210,N_18927,N_18192);
xor U19211 (N_19211,N_18436,N_18302);
nor U19212 (N_19212,N_18145,N_18675);
and U19213 (N_19213,N_18226,N_18256);
nand U19214 (N_19214,N_18375,N_18191);
and U19215 (N_19215,N_18942,N_18447);
and U19216 (N_19216,N_18581,N_18028);
xor U19217 (N_19217,N_18067,N_18346);
nor U19218 (N_19218,N_18143,N_18347);
nand U19219 (N_19219,N_18725,N_18859);
nor U19220 (N_19220,N_18350,N_18247);
and U19221 (N_19221,N_18242,N_18294);
nand U19222 (N_19222,N_18738,N_18300);
or U19223 (N_19223,N_18283,N_18012);
and U19224 (N_19224,N_18282,N_18930);
xnor U19225 (N_19225,N_18544,N_18835);
nand U19226 (N_19226,N_18484,N_18099);
nand U19227 (N_19227,N_18370,N_18098);
nand U19228 (N_19228,N_18221,N_18552);
and U19229 (N_19229,N_18842,N_18934);
xor U19230 (N_19230,N_18515,N_18514);
xnor U19231 (N_19231,N_18292,N_18336);
nand U19232 (N_19232,N_18422,N_18887);
nand U19233 (N_19233,N_18665,N_18954);
xor U19234 (N_19234,N_18973,N_18365);
nor U19235 (N_19235,N_18799,N_18808);
xnor U19236 (N_19236,N_18845,N_18778);
nor U19237 (N_19237,N_18148,N_18744);
nor U19238 (N_19238,N_18063,N_18997);
nand U19239 (N_19239,N_18658,N_18822);
nand U19240 (N_19240,N_18654,N_18914);
nand U19241 (N_19241,N_18388,N_18746);
nand U19242 (N_19242,N_18770,N_18603);
xnor U19243 (N_19243,N_18468,N_18120);
nand U19244 (N_19244,N_18272,N_18912);
or U19245 (N_19245,N_18183,N_18978);
nor U19246 (N_19246,N_18358,N_18722);
or U19247 (N_19247,N_18962,N_18943);
and U19248 (N_19248,N_18083,N_18423);
nor U19249 (N_19249,N_18220,N_18355);
and U19250 (N_19250,N_18006,N_18364);
or U19251 (N_19251,N_18159,N_18360);
nor U19252 (N_19252,N_18819,N_18882);
xnor U19253 (N_19253,N_18670,N_18005);
xnor U19254 (N_19254,N_18402,N_18590);
xnor U19255 (N_19255,N_18611,N_18699);
xor U19256 (N_19256,N_18240,N_18830);
and U19257 (N_19257,N_18204,N_18518);
nand U19258 (N_19258,N_18369,N_18096);
xnor U19259 (N_19259,N_18124,N_18433);
xnor U19260 (N_19260,N_18521,N_18295);
xnor U19261 (N_19261,N_18057,N_18599);
nand U19262 (N_19262,N_18691,N_18925);
or U19263 (N_19263,N_18091,N_18326);
and U19264 (N_19264,N_18955,N_18174);
nor U19265 (N_19265,N_18751,N_18100);
nor U19266 (N_19266,N_18038,N_18048);
nand U19267 (N_19267,N_18222,N_18571);
nand U19268 (N_19268,N_18577,N_18774);
or U19269 (N_19269,N_18640,N_18667);
nor U19270 (N_19270,N_18959,N_18008);
and U19271 (N_19271,N_18075,N_18610);
nand U19272 (N_19272,N_18138,N_18366);
xnor U19273 (N_19273,N_18384,N_18556);
xnor U19274 (N_19274,N_18092,N_18918);
and U19275 (N_19275,N_18917,N_18775);
xnor U19276 (N_19276,N_18066,N_18601);
or U19277 (N_19277,N_18996,N_18677);
xor U19278 (N_19278,N_18418,N_18490);
nor U19279 (N_19279,N_18628,N_18936);
nor U19280 (N_19280,N_18348,N_18865);
nand U19281 (N_19281,N_18940,N_18779);
or U19282 (N_19282,N_18817,N_18898);
or U19283 (N_19283,N_18826,N_18339);
or U19284 (N_19284,N_18833,N_18614);
nand U19285 (N_19285,N_18332,N_18367);
nor U19286 (N_19286,N_18874,N_18605);
or U19287 (N_19287,N_18742,N_18196);
xor U19288 (N_19288,N_18561,N_18254);
nand U19289 (N_19289,N_18049,N_18862);
nor U19290 (N_19290,N_18255,N_18286);
and U19291 (N_19291,N_18210,N_18071);
or U19292 (N_19292,N_18162,N_18351);
or U19293 (N_19293,N_18761,N_18441);
xnor U19294 (N_19294,N_18584,N_18399);
and U19295 (N_19295,N_18101,N_18693);
and U19296 (N_19296,N_18527,N_18720);
or U19297 (N_19297,N_18280,N_18661);
nor U19298 (N_19298,N_18697,N_18158);
nand U19299 (N_19299,N_18624,N_18371);
and U19300 (N_19300,N_18853,N_18950);
and U19301 (N_19301,N_18408,N_18908);
xor U19302 (N_19302,N_18567,N_18155);
xor U19303 (N_19303,N_18231,N_18314);
nand U19304 (N_19304,N_18638,N_18504);
or U19305 (N_19305,N_18724,N_18516);
or U19306 (N_19306,N_18984,N_18059);
nor U19307 (N_19307,N_18299,N_18923);
or U19308 (N_19308,N_18043,N_18026);
xnor U19309 (N_19309,N_18844,N_18924);
xor U19310 (N_19310,N_18458,N_18957);
nand U19311 (N_19311,N_18239,N_18108);
or U19312 (N_19312,N_18595,N_18825);
xor U19313 (N_19313,N_18463,N_18814);
nor U19314 (N_19314,N_18644,N_18084);
xnor U19315 (N_19315,N_18824,N_18750);
and U19316 (N_19316,N_18487,N_18974);
nand U19317 (N_19317,N_18506,N_18232);
xor U19318 (N_19318,N_18919,N_18752);
or U19319 (N_19319,N_18070,N_18717);
nor U19320 (N_19320,N_18013,N_18731);
or U19321 (N_19321,N_18733,N_18916);
or U19322 (N_19322,N_18327,N_18895);
or U19323 (N_19323,N_18838,N_18248);
nor U19324 (N_19324,N_18260,N_18198);
or U19325 (N_19325,N_18456,N_18626);
xnor U19326 (N_19326,N_18214,N_18259);
nand U19327 (N_19327,N_18171,N_18225);
xor U19328 (N_19328,N_18651,N_18627);
xnor U19329 (N_19329,N_18998,N_18150);
xnor U19330 (N_19330,N_18153,N_18641);
or U19331 (N_19331,N_18982,N_18073);
xor U19332 (N_19332,N_18910,N_18517);
and U19333 (N_19333,N_18650,N_18780);
xor U19334 (N_19334,N_18390,N_18133);
xnor U19335 (N_19335,N_18786,N_18507);
or U19336 (N_19336,N_18947,N_18421);
or U19337 (N_19337,N_18029,N_18669);
or U19338 (N_19338,N_18211,N_18045);
nor U19339 (N_19339,N_18876,N_18696);
nand U19340 (N_19340,N_18102,N_18445);
nor U19341 (N_19341,N_18493,N_18616);
nand U19342 (N_19342,N_18791,N_18011);
or U19343 (N_19343,N_18356,N_18591);
or U19344 (N_19344,N_18209,N_18929);
nor U19345 (N_19345,N_18530,N_18574);
xnor U19346 (N_19346,N_18156,N_18866);
or U19347 (N_19347,N_18444,N_18412);
or U19348 (N_19348,N_18537,N_18233);
and U19349 (N_19349,N_18270,N_18622);
nor U19350 (N_19350,N_18714,N_18427);
nand U19351 (N_19351,N_18076,N_18476);
and U19352 (N_19352,N_18913,N_18053);
nor U19353 (N_19353,N_18632,N_18975);
nor U19354 (N_19354,N_18798,N_18265);
xor U19355 (N_19355,N_18708,N_18976);
nor U19356 (N_19356,N_18960,N_18430);
and U19357 (N_19357,N_18003,N_18469);
or U19358 (N_19358,N_18368,N_18014);
xor U19359 (N_19359,N_18362,N_18307);
or U19360 (N_19360,N_18121,N_18505);
or U19361 (N_19361,N_18760,N_18881);
and U19362 (N_19362,N_18587,N_18969);
nand U19363 (N_19363,N_18379,N_18268);
nand U19364 (N_19364,N_18465,N_18149);
and U19365 (N_19365,N_18415,N_18180);
xor U19366 (N_19366,N_18589,N_18110);
nor U19367 (N_19367,N_18032,N_18602);
xor U19368 (N_19368,N_18885,N_18267);
xnor U19369 (N_19369,N_18802,N_18331);
nor U19370 (N_19370,N_18939,N_18409);
or U19371 (N_19371,N_18498,N_18154);
nor U19372 (N_19372,N_18030,N_18285);
nor U19373 (N_19373,N_18058,N_18015);
xnor U19374 (N_19374,N_18119,N_18448);
xnor U19375 (N_19375,N_18106,N_18035);
nor U19376 (N_19376,N_18945,N_18652);
or U19377 (N_19377,N_18718,N_18227);
xor U19378 (N_19378,N_18829,N_18019);
nand U19379 (N_19379,N_18361,N_18588);
xor U19380 (N_19380,N_18630,N_18508);
nor U19381 (N_19381,N_18432,N_18732);
or U19382 (N_19382,N_18163,N_18594);
xnor U19383 (N_19383,N_18410,N_18039);
nor U19384 (N_19384,N_18604,N_18337);
or U19385 (N_19385,N_18116,N_18027);
xor U19386 (N_19386,N_18109,N_18702);
xor U19387 (N_19387,N_18462,N_18178);
and U19388 (N_19388,N_18062,N_18054);
nor U19389 (N_19389,N_18555,N_18660);
nor U19390 (N_19390,N_18329,N_18522);
or U19391 (N_19391,N_18301,N_18494);
nor U19392 (N_19392,N_18177,N_18848);
nand U19393 (N_19393,N_18586,N_18768);
or U19394 (N_19394,N_18296,N_18021);
nand U19395 (N_19395,N_18308,N_18212);
nand U19396 (N_19396,N_18597,N_18374);
or U19397 (N_19397,N_18213,N_18077);
nor U19398 (N_19398,N_18443,N_18668);
nand U19399 (N_19399,N_18500,N_18944);
and U19400 (N_19400,N_18140,N_18130);
nand U19401 (N_19401,N_18803,N_18864);
or U19402 (N_19402,N_18765,N_18333);
or U19403 (N_19403,N_18305,N_18000);
nand U19404 (N_19404,N_18868,N_18291);
nor U19405 (N_19405,N_18554,N_18583);
nor U19406 (N_19406,N_18526,N_18968);
nor U19407 (N_19407,N_18686,N_18122);
xor U19408 (N_19408,N_18173,N_18261);
or U19409 (N_19409,N_18342,N_18809);
or U19410 (N_19410,N_18010,N_18111);
nor U19411 (N_19411,N_18078,N_18269);
nand U19412 (N_19412,N_18569,N_18951);
nand U19413 (N_19413,N_18900,N_18538);
nor U19414 (N_19414,N_18967,N_18477);
nor U19415 (N_19415,N_18643,N_18519);
nor U19416 (N_19416,N_18181,N_18051);
or U19417 (N_19417,N_18899,N_18727);
and U19418 (N_19418,N_18085,N_18275);
and U19419 (N_19419,N_18460,N_18977);
nor U19420 (N_19420,N_18525,N_18903);
nand U19421 (N_19421,N_18306,N_18377);
nand U19422 (N_19422,N_18891,N_18097);
nand U19423 (N_19423,N_18889,N_18672);
or U19424 (N_19424,N_18625,N_18197);
and U19425 (N_19425,N_18234,N_18420);
nand U19426 (N_19426,N_18856,N_18553);
nor U19427 (N_19427,N_18135,N_18080);
or U19428 (N_19428,N_18406,N_18065);
or U19429 (N_19429,N_18562,N_18320);
nor U19430 (N_19430,N_18685,N_18710);
and U19431 (N_19431,N_18728,N_18319);
xnor U19432 (N_19432,N_18655,N_18849);
nand U19433 (N_19433,N_18739,N_18470);
or U19434 (N_19434,N_18596,N_18403);
xnor U19435 (N_19435,N_18251,N_18182);
or U19436 (N_19436,N_18160,N_18807);
nor U19437 (N_19437,N_18123,N_18129);
nor U19438 (N_19438,N_18510,N_18253);
nand U19439 (N_19439,N_18785,N_18001);
and U19440 (N_19440,N_18175,N_18257);
and U19441 (N_19441,N_18932,N_18481);
xnor U19442 (N_19442,N_18847,N_18828);
nand U19443 (N_19443,N_18531,N_18216);
xnor U19444 (N_19444,N_18107,N_18818);
or U19445 (N_19445,N_18990,N_18042);
or U19446 (N_19446,N_18681,N_18431);
nor U19447 (N_19447,N_18634,N_18811);
nor U19448 (N_19448,N_18712,N_18659);
nor U19449 (N_19449,N_18372,N_18823);
and U19450 (N_19450,N_18471,N_18827);
nand U19451 (N_19451,N_18164,N_18118);
or U19452 (N_19452,N_18723,N_18044);
nor U19453 (N_19453,N_18137,N_18208);
and U19454 (N_19454,N_18378,N_18457);
or U19455 (N_19455,N_18575,N_18205);
nor U19456 (N_19456,N_18502,N_18767);
or U19457 (N_19457,N_18533,N_18024);
and U19458 (N_19458,N_18758,N_18726);
or U19459 (N_19459,N_18663,N_18404);
nor U19460 (N_19460,N_18528,N_18467);
or U19461 (N_19461,N_18316,N_18312);
nor U19462 (N_19462,N_18353,N_18341);
nor U19463 (N_19463,N_18104,N_18090);
xnor U19464 (N_19464,N_18860,N_18784);
or U19465 (N_19465,N_18867,N_18322);
and U19466 (N_19466,N_18512,N_18394);
xnor U19467 (N_19467,N_18568,N_18707);
and U19468 (N_19468,N_18036,N_18970);
and U19469 (N_19469,N_18023,N_18002);
nand U19470 (N_19470,N_18557,N_18872);
and U19471 (N_19471,N_18429,N_18134);
nand U19472 (N_19472,N_18203,N_18474);
and U19473 (N_19473,N_18189,N_18965);
nand U19474 (N_19474,N_18274,N_18999);
and U19475 (N_19475,N_18877,N_18972);
or U19476 (N_19476,N_18694,N_18496);
nor U19477 (N_19477,N_18489,N_18115);
nand U19478 (N_19478,N_18813,N_18743);
and U19479 (N_19479,N_18804,N_18815);
or U19480 (N_19480,N_18565,N_18318);
and U19481 (N_19481,N_18459,N_18963);
and U19482 (N_19482,N_18079,N_18816);
nor U19483 (N_19483,N_18579,N_18438);
or U19484 (N_19484,N_18451,N_18683);
xor U19485 (N_19485,N_18657,N_18323);
xor U19486 (N_19486,N_18971,N_18692);
nand U19487 (N_19487,N_18585,N_18383);
xnor U19488 (N_19488,N_18888,N_18820);
nor U19489 (N_19489,N_18647,N_18193);
xor U19490 (N_19490,N_18055,N_18343);
nand U19491 (N_19491,N_18772,N_18004);
xor U19492 (N_19492,N_18698,N_18709);
xnor U19493 (N_19493,N_18904,N_18131);
nor U19494 (N_19494,N_18186,N_18113);
nor U19495 (N_19495,N_18125,N_18920);
xor U19496 (N_19496,N_18639,N_18064);
nor U19497 (N_19497,N_18606,N_18792);
and U19498 (N_19498,N_18935,N_18741);
or U19499 (N_19499,N_18609,N_18836);
or U19500 (N_19500,N_18329,N_18990);
nor U19501 (N_19501,N_18276,N_18372);
and U19502 (N_19502,N_18768,N_18941);
and U19503 (N_19503,N_18714,N_18247);
xnor U19504 (N_19504,N_18754,N_18044);
xnor U19505 (N_19505,N_18662,N_18078);
nand U19506 (N_19506,N_18760,N_18582);
or U19507 (N_19507,N_18382,N_18237);
or U19508 (N_19508,N_18122,N_18726);
or U19509 (N_19509,N_18630,N_18444);
xnor U19510 (N_19510,N_18679,N_18405);
nor U19511 (N_19511,N_18214,N_18966);
nor U19512 (N_19512,N_18009,N_18390);
nor U19513 (N_19513,N_18401,N_18024);
nor U19514 (N_19514,N_18208,N_18631);
xor U19515 (N_19515,N_18688,N_18067);
nor U19516 (N_19516,N_18621,N_18021);
nor U19517 (N_19517,N_18279,N_18331);
or U19518 (N_19518,N_18174,N_18476);
nand U19519 (N_19519,N_18940,N_18484);
and U19520 (N_19520,N_18611,N_18427);
nand U19521 (N_19521,N_18983,N_18267);
or U19522 (N_19522,N_18922,N_18321);
xor U19523 (N_19523,N_18361,N_18378);
or U19524 (N_19524,N_18058,N_18223);
nor U19525 (N_19525,N_18577,N_18941);
nand U19526 (N_19526,N_18993,N_18654);
xnor U19527 (N_19527,N_18389,N_18002);
or U19528 (N_19528,N_18485,N_18441);
or U19529 (N_19529,N_18074,N_18225);
and U19530 (N_19530,N_18079,N_18410);
xor U19531 (N_19531,N_18249,N_18523);
or U19532 (N_19532,N_18720,N_18920);
nor U19533 (N_19533,N_18952,N_18149);
nor U19534 (N_19534,N_18232,N_18241);
and U19535 (N_19535,N_18647,N_18969);
nor U19536 (N_19536,N_18366,N_18369);
or U19537 (N_19537,N_18754,N_18946);
nand U19538 (N_19538,N_18960,N_18084);
or U19539 (N_19539,N_18339,N_18523);
xor U19540 (N_19540,N_18614,N_18732);
nor U19541 (N_19541,N_18375,N_18597);
xnor U19542 (N_19542,N_18921,N_18021);
xor U19543 (N_19543,N_18655,N_18041);
nand U19544 (N_19544,N_18054,N_18595);
and U19545 (N_19545,N_18442,N_18718);
nand U19546 (N_19546,N_18643,N_18428);
or U19547 (N_19547,N_18578,N_18501);
or U19548 (N_19548,N_18455,N_18212);
xnor U19549 (N_19549,N_18956,N_18320);
xor U19550 (N_19550,N_18990,N_18452);
nand U19551 (N_19551,N_18759,N_18897);
nand U19552 (N_19552,N_18652,N_18998);
or U19553 (N_19553,N_18236,N_18400);
nor U19554 (N_19554,N_18442,N_18572);
nand U19555 (N_19555,N_18173,N_18142);
or U19556 (N_19556,N_18045,N_18487);
nand U19557 (N_19557,N_18474,N_18209);
or U19558 (N_19558,N_18931,N_18836);
and U19559 (N_19559,N_18045,N_18978);
nor U19560 (N_19560,N_18688,N_18371);
nor U19561 (N_19561,N_18295,N_18093);
xnor U19562 (N_19562,N_18871,N_18393);
and U19563 (N_19563,N_18726,N_18044);
xnor U19564 (N_19564,N_18469,N_18344);
and U19565 (N_19565,N_18943,N_18735);
nand U19566 (N_19566,N_18154,N_18469);
xor U19567 (N_19567,N_18440,N_18307);
or U19568 (N_19568,N_18788,N_18320);
xor U19569 (N_19569,N_18700,N_18462);
nand U19570 (N_19570,N_18339,N_18350);
and U19571 (N_19571,N_18819,N_18157);
nor U19572 (N_19572,N_18534,N_18619);
nor U19573 (N_19573,N_18482,N_18655);
nand U19574 (N_19574,N_18283,N_18568);
nand U19575 (N_19575,N_18849,N_18434);
nand U19576 (N_19576,N_18857,N_18567);
and U19577 (N_19577,N_18888,N_18384);
nand U19578 (N_19578,N_18352,N_18095);
xnor U19579 (N_19579,N_18131,N_18757);
nand U19580 (N_19580,N_18084,N_18501);
nor U19581 (N_19581,N_18607,N_18969);
nor U19582 (N_19582,N_18924,N_18854);
nand U19583 (N_19583,N_18211,N_18210);
nor U19584 (N_19584,N_18176,N_18106);
or U19585 (N_19585,N_18341,N_18852);
nand U19586 (N_19586,N_18023,N_18719);
and U19587 (N_19587,N_18713,N_18708);
nand U19588 (N_19588,N_18778,N_18111);
nand U19589 (N_19589,N_18633,N_18218);
xnor U19590 (N_19590,N_18835,N_18996);
nand U19591 (N_19591,N_18176,N_18812);
and U19592 (N_19592,N_18247,N_18726);
nand U19593 (N_19593,N_18096,N_18499);
or U19594 (N_19594,N_18487,N_18080);
nand U19595 (N_19595,N_18471,N_18664);
xor U19596 (N_19596,N_18779,N_18182);
or U19597 (N_19597,N_18232,N_18657);
nor U19598 (N_19598,N_18847,N_18923);
and U19599 (N_19599,N_18584,N_18930);
nand U19600 (N_19600,N_18157,N_18303);
nand U19601 (N_19601,N_18282,N_18482);
nor U19602 (N_19602,N_18141,N_18302);
xor U19603 (N_19603,N_18597,N_18495);
or U19604 (N_19604,N_18875,N_18745);
and U19605 (N_19605,N_18413,N_18324);
nor U19606 (N_19606,N_18856,N_18800);
and U19607 (N_19607,N_18207,N_18426);
nor U19608 (N_19608,N_18155,N_18936);
nor U19609 (N_19609,N_18410,N_18188);
xor U19610 (N_19610,N_18190,N_18057);
xor U19611 (N_19611,N_18742,N_18067);
or U19612 (N_19612,N_18026,N_18441);
or U19613 (N_19613,N_18198,N_18104);
xnor U19614 (N_19614,N_18110,N_18511);
nand U19615 (N_19615,N_18935,N_18980);
nand U19616 (N_19616,N_18167,N_18726);
xor U19617 (N_19617,N_18019,N_18934);
or U19618 (N_19618,N_18724,N_18223);
nor U19619 (N_19619,N_18018,N_18477);
nand U19620 (N_19620,N_18378,N_18349);
nor U19621 (N_19621,N_18217,N_18781);
nor U19622 (N_19622,N_18741,N_18624);
or U19623 (N_19623,N_18089,N_18680);
or U19624 (N_19624,N_18786,N_18212);
or U19625 (N_19625,N_18608,N_18953);
and U19626 (N_19626,N_18015,N_18351);
nand U19627 (N_19627,N_18480,N_18254);
and U19628 (N_19628,N_18784,N_18166);
nand U19629 (N_19629,N_18213,N_18058);
or U19630 (N_19630,N_18487,N_18839);
and U19631 (N_19631,N_18855,N_18668);
nor U19632 (N_19632,N_18875,N_18782);
or U19633 (N_19633,N_18387,N_18252);
nor U19634 (N_19634,N_18531,N_18986);
or U19635 (N_19635,N_18116,N_18818);
nor U19636 (N_19636,N_18392,N_18448);
xnor U19637 (N_19637,N_18554,N_18406);
nor U19638 (N_19638,N_18283,N_18597);
nor U19639 (N_19639,N_18493,N_18436);
nand U19640 (N_19640,N_18511,N_18946);
or U19641 (N_19641,N_18645,N_18699);
xor U19642 (N_19642,N_18282,N_18974);
nor U19643 (N_19643,N_18768,N_18997);
nor U19644 (N_19644,N_18103,N_18946);
nand U19645 (N_19645,N_18675,N_18937);
nor U19646 (N_19646,N_18478,N_18068);
and U19647 (N_19647,N_18751,N_18759);
and U19648 (N_19648,N_18923,N_18937);
nand U19649 (N_19649,N_18300,N_18939);
xor U19650 (N_19650,N_18241,N_18276);
xnor U19651 (N_19651,N_18535,N_18350);
nor U19652 (N_19652,N_18950,N_18247);
nor U19653 (N_19653,N_18051,N_18708);
or U19654 (N_19654,N_18284,N_18940);
nor U19655 (N_19655,N_18076,N_18904);
xnor U19656 (N_19656,N_18735,N_18750);
xnor U19657 (N_19657,N_18738,N_18351);
xnor U19658 (N_19658,N_18971,N_18178);
xor U19659 (N_19659,N_18632,N_18721);
nand U19660 (N_19660,N_18634,N_18974);
nor U19661 (N_19661,N_18400,N_18893);
nand U19662 (N_19662,N_18716,N_18610);
nor U19663 (N_19663,N_18104,N_18293);
or U19664 (N_19664,N_18114,N_18458);
nand U19665 (N_19665,N_18330,N_18679);
nand U19666 (N_19666,N_18636,N_18914);
nand U19667 (N_19667,N_18168,N_18199);
or U19668 (N_19668,N_18406,N_18208);
nor U19669 (N_19669,N_18502,N_18696);
nand U19670 (N_19670,N_18886,N_18912);
xnor U19671 (N_19671,N_18712,N_18563);
nor U19672 (N_19672,N_18453,N_18495);
and U19673 (N_19673,N_18020,N_18814);
xnor U19674 (N_19674,N_18681,N_18123);
nand U19675 (N_19675,N_18954,N_18077);
nor U19676 (N_19676,N_18796,N_18348);
xnor U19677 (N_19677,N_18072,N_18184);
nor U19678 (N_19678,N_18793,N_18248);
nor U19679 (N_19679,N_18245,N_18668);
or U19680 (N_19680,N_18788,N_18988);
nand U19681 (N_19681,N_18478,N_18955);
and U19682 (N_19682,N_18495,N_18199);
xnor U19683 (N_19683,N_18369,N_18808);
nor U19684 (N_19684,N_18011,N_18663);
xnor U19685 (N_19685,N_18630,N_18251);
nand U19686 (N_19686,N_18399,N_18821);
or U19687 (N_19687,N_18414,N_18750);
nor U19688 (N_19688,N_18670,N_18474);
xnor U19689 (N_19689,N_18750,N_18475);
xnor U19690 (N_19690,N_18363,N_18268);
nor U19691 (N_19691,N_18660,N_18689);
and U19692 (N_19692,N_18402,N_18255);
nor U19693 (N_19693,N_18018,N_18021);
xor U19694 (N_19694,N_18152,N_18369);
xor U19695 (N_19695,N_18274,N_18607);
and U19696 (N_19696,N_18140,N_18193);
and U19697 (N_19697,N_18910,N_18157);
nand U19698 (N_19698,N_18977,N_18933);
or U19699 (N_19699,N_18351,N_18625);
or U19700 (N_19700,N_18218,N_18682);
or U19701 (N_19701,N_18445,N_18326);
nor U19702 (N_19702,N_18436,N_18787);
xnor U19703 (N_19703,N_18455,N_18536);
or U19704 (N_19704,N_18319,N_18125);
or U19705 (N_19705,N_18241,N_18686);
nand U19706 (N_19706,N_18552,N_18337);
nand U19707 (N_19707,N_18160,N_18994);
nand U19708 (N_19708,N_18726,N_18549);
or U19709 (N_19709,N_18740,N_18370);
nand U19710 (N_19710,N_18006,N_18102);
nand U19711 (N_19711,N_18524,N_18386);
or U19712 (N_19712,N_18496,N_18345);
nor U19713 (N_19713,N_18110,N_18558);
nand U19714 (N_19714,N_18141,N_18478);
or U19715 (N_19715,N_18064,N_18856);
nor U19716 (N_19716,N_18413,N_18351);
nor U19717 (N_19717,N_18953,N_18312);
or U19718 (N_19718,N_18838,N_18825);
nor U19719 (N_19719,N_18214,N_18816);
and U19720 (N_19720,N_18679,N_18743);
nor U19721 (N_19721,N_18676,N_18621);
and U19722 (N_19722,N_18082,N_18597);
or U19723 (N_19723,N_18853,N_18298);
nand U19724 (N_19724,N_18515,N_18574);
xor U19725 (N_19725,N_18946,N_18357);
nand U19726 (N_19726,N_18935,N_18004);
nor U19727 (N_19727,N_18614,N_18876);
nor U19728 (N_19728,N_18514,N_18976);
or U19729 (N_19729,N_18640,N_18365);
xnor U19730 (N_19730,N_18826,N_18197);
xnor U19731 (N_19731,N_18876,N_18628);
nand U19732 (N_19732,N_18874,N_18509);
xnor U19733 (N_19733,N_18611,N_18076);
nand U19734 (N_19734,N_18316,N_18566);
nand U19735 (N_19735,N_18457,N_18446);
xnor U19736 (N_19736,N_18591,N_18651);
and U19737 (N_19737,N_18794,N_18263);
and U19738 (N_19738,N_18752,N_18989);
nor U19739 (N_19739,N_18266,N_18130);
and U19740 (N_19740,N_18414,N_18326);
or U19741 (N_19741,N_18568,N_18998);
nand U19742 (N_19742,N_18440,N_18377);
and U19743 (N_19743,N_18702,N_18322);
nand U19744 (N_19744,N_18137,N_18960);
nor U19745 (N_19745,N_18118,N_18609);
xnor U19746 (N_19746,N_18408,N_18434);
nor U19747 (N_19747,N_18475,N_18710);
or U19748 (N_19748,N_18674,N_18811);
or U19749 (N_19749,N_18071,N_18548);
xnor U19750 (N_19750,N_18646,N_18988);
and U19751 (N_19751,N_18670,N_18859);
nand U19752 (N_19752,N_18616,N_18402);
or U19753 (N_19753,N_18431,N_18271);
or U19754 (N_19754,N_18345,N_18908);
nor U19755 (N_19755,N_18288,N_18533);
and U19756 (N_19756,N_18908,N_18552);
or U19757 (N_19757,N_18924,N_18677);
nor U19758 (N_19758,N_18785,N_18409);
nand U19759 (N_19759,N_18726,N_18825);
nor U19760 (N_19760,N_18636,N_18143);
nor U19761 (N_19761,N_18924,N_18194);
or U19762 (N_19762,N_18565,N_18420);
and U19763 (N_19763,N_18432,N_18693);
nor U19764 (N_19764,N_18996,N_18362);
nor U19765 (N_19765,N_18664,N_18079);
and U19766 (N_19766,N_18287,N_18102);
or U19767 (N_19767,N_18354,N_18432);
or U19768 (N_19768,N_18424,N_18601);
or U19769 (N_19769,N_18403,N_18565);
nand U19770 (N_19770,N_18898,N_18114);
and U19771 (N_19771,N_18597,N_18363);
nand U19772 (N_19772,N_18981,N_18477);
nand U19773 (N_19773,N_18088,N_18791);
nor U19774 (N_19774,N_18638,N_18239);
and U19775 (N_19775,N_18162,N_18881);
nand U19776 (N_19776,N_18184,N_18801);
or U19777 (N_19777,N_18781,N_18116);
or U19778 (N_19778,N_18911,N_18025);
nor U19779 (N_19779,N_18946,N_18740);
nor U19780 (N_19780,N_18541,N_18991);
nand U19781 (N_19781,N_18605,N_18236);
or U19782 (N_19782,N_18728,N_18977);
xor U19783 (N_19783,N_18953,N_18665);
or U19784 (N_19784,N_18010,N_18148);
nand U19785 (N_19785,N_18545,N_18134);
nor U19786 (N_19786,N_18421,N_18216);
and U19787 (N_19787,N_18077,N_18504);
nand U19788 (N_19788,N_18529,N_18623);
and U19789 (N_19789,N_18279,N_18026);
and U19790 (N_19790,N_18401,N_18072);
nor U19791 (N_19791,N_18419,N_18978);
and U19792 (N_19792,N_18127,N_18401);
nor U19793 (N_19793,N_18935,N_18217);
and U19794 (N_19794,N_18733,N_18470);
xor U19795 (N_19795,N_18418,N_18542);
or U19796 (N_19796,N_18752,N_18341);
or U19797 (N_19797,N_18230,N_18386);
nand U19798 (N_19798,N_18329,N_18485);
xor U19799 (N_19799,N_18454,N_18599);
nand U19800 (N_19800,N_18757,N_18990);
nor U19801 (N_19801,N_18653,N_18490);
nand U19802 (N_19802,N_18063,N_18059);
or U19803 (N_19803,N_18967,N_18596);
xnor U19804 (N_19804,N_18919,N_18578);
xnor U19805 (N_19805,N_18824,N_18945);
and U19806 (N_19806,N_18772,N_18030);
or U19807 (N_19807,N_18653,N_18549);
and U19808 (N_19808,N_18250,N_18304);
xor U19809 (N_19809,N_18789,N_18727);
or U19810 (N_19810,N_18214,N_18954);
xor U19811 (N_19811,N_18629,N_18246);
and U19812 (N_19812,N_18481,N_18102);
xor U19813 (N_19813,N_18687,N_18106);
or U19814 (N_19814,N_18863,N_18948);
nand U19815 (N_19815,N_18642,N_18040);
and U19816 (N_19816,N_18529,N_18307);
and U19817 (N_19817,N_18215,N_18638);
xnor U19818 (N_19818,N_18552,N_18255);
and U19819 (N_19819,N_18529,N_18884);
nand U19820 (N_19820,N_18870,N_18499);
or U19821 (N_19821,N_18475,N_18348);
nor U19822 (N_19822,N_18110,N_18871);
nand U19823 (N_19823,N_18196,N_18782);
nand U19824 (N_19824,N_18346,N_18138);
xnor U19825 (N_19825,N_18807,N_18444);
xnor U19826 (N_19826,N_18097,N_18876);
and U19827 (N_19827,N_18216,N_18205);
or U19828 (N_19828,N_18635,N_18760);
or U19829 (N_19829,N_18712,N_18141);
xor U19830 (N_19830,N_18143,N_18751);
nand U19831 (N_19831,N_18097,N_18259);
nand U19832 (N_19832,N_18860,N_18896);
and U19833 (N_19833,N_18881,N_18415);
xnor U19834 (N_19834,N_18340,N_18030);
and U19835 (N_19835,N_18974,N_18329);
and U19836 (N_19836,N_18472,N_18761);
or U19837 (N_19837,N_18454,N_18302);
nor U19838 (N_19838,N_18899,N_18323);
nor U19839 (N_19839,N_18239,N_18376);
nor U19840 (N_19840,N_18576,N_18543);
nor U19841 (N_19841,N_18374,N_18167);
or U19842 (N_19842,N_18279,N_18491);
nand U19843 (N_19843,N_18390,N_18283);
or U19844 (N_19844,N_18726,N_18717);
nand U19845 (N_19845,N_18522,N_18131);
and U19846 (N_19846,N_18407,N_18771);
nor U19847 (N_19847,N_18303,N_18922);
nor U19848 (N_19848,N_18487,N_18428);
nor U19849 (N_19849,N_18634,N_18578);
or U19850 (N_19850,N_18128,N_18911);
xor U19851 (N_19851,N_18877,N_18649);
nor U19852 (N_19852,N_18589,N_18906);
nand U19853 (N_19853,N_18892,N_18029);
xnor U19854 (N_19854,N_18115,N_18450);
nor U19855 (N_19855,N_18117,N_18974);
or U19856 (N_19856,N_18635,N_18488);
and U19857 (N_19857,N_18032,N_18708);
and U19858 (N_19858,N_18378,N_18252);
nand U19859 (N_19859,N_18793,N_18481);
nand U19860 (N_19860,N_18206,N_18895);
nand U19861 (N_19861,N_18472,N_18446);
or U19862 (N_19862,N_18336,N_18195);
nor U19863 (N_19863,N_18833,N_18026);
and U19864 (N_19864,N_18586,N_18916);
and U19865 (N_19865,N_18396,N_18265);
and U19866 (N_19866,N_18480,N_18565);
nor U19867 (N_19867,N_18930,N_18222);
and U19868 (N_19868,N_18408,N_18001);
nand U19869 (N_19869,N_18472,N_18996);
and U19870 (N_19870,N_18837,N_18207);
xnor U19871 (N_19871,N_18030,N_18663);
and U19872 (N_19872,N_18937,N_18436);
and U19873 (N_19873,N_18903,N_18185);
xnor U19874 (N_19874,N_18416,N_18151);
nand U19875 (N_19875,N_18814,N_18410);
and U19876 (N_19876,N_18311,N_18356);
xor U19877 (N_19877,N_18939,N_18442);
nand U19878 (N_19878,N_18714,N_18261);
xor U19879 (N_19879,N_18925,N_18328);
and U19880 (N_19880,N_18624,N_18199);
xor U19881 (N_19881,N_18043,N_18227);
nor U19882 (N_19882,N_18011,N_18200);
nor U19883 (N_19883,N_18897,N_18431);
or U19884 (N_19884,N_18273,N_18554);
and U19885 (N_19885,N_18706,N_18907);
or U19886 (N_19886,N_18456,N_18217);
nand U19887 (N_19887,N_18081,N_18325);
and U19888 (N_19888,N_18840,N_18566);
xnor U19889 (N_19889,N_18676,N_18661);
nand U19890 (N_19890,N_18097,N_18810);
xnor U19891 (N_19891,N_18656,N_18286);
nor U19892 (N_19892,N_18909,N_18922);
or U19893 (N_19893,N_18342,N_18767);
xor U19894 (N_19894,N_18266,N_18023);
and U19895 (N_19895,N_18575,N_18532);
nor U19896 (N_19896,N_18316,N_18812);
nand U19897 (N_19897,N_18780,N_18505);
nor U19898 (N_19898,N_18912,N_18101);
and U19899 (N_19899,N_18675,N_18421);
or U19900 (N_19900,N_18044,N_18993);
nor U19901 (N_19901,N_18510,N_18656);
nor U19902 (N_19902,N_18506,N_18531);
nand U19903 (N_19903,N_18592,N_18509);
nand U19904 (N_19904,N_18407,N_18769);
nand U19905 (N_19905,N_18556,N_18526);
nand U19906 (N_19906,N_18737,N_18990);
nand U19907 (N_19907,N_18939,N_18988);
nand U19908 (N_19908,N_18765,N_18517);
xor U19909 (N_19909,N_18759,N_18244);
and U19910 (N_19910,N_18546,N_18912);
and U19911 (N_19911,N_18986,N_18037);
xnor U19912 (N_19912,N_18857,N_18593);
nor U19913 (N_19913,N_18554,N_18781);
nand U19914 (N_19914,N_18768,N_18431);
and U19915 (N_19915,N_18968,N_18802);
nor U19916 (N_19916,N_18306,N_18718);
nor U19917 (N_19917,N_18508,N_18796);
or U19918 (N_19918,N_18880,N_18889);
nand U19919 (N_19919,N_18806,N_18567);
xor U19920 (N_19920,N_18510,N_18559);
or U19921 (N_19921,N_18845,N_18635);
or U19922 (N_19922,N_18452,N_18360);
nor U19923 (N_19923,N_18571,N_18553);
or U19924 (N_19924,N_18832,N_18459);
nor U19925 (N_19925,N_18106,N_18865);
or U19926 (N_19926,N_18544,N_18749);
or U19927 (N_19927,N_18326,N_18310);
nand U19928 (N_19928,N_18936,N_18127);
and U19929 (N_19929,N_18766,N_18475);
and U19930 (N_19930,N_18925,N_18483);
nand U19931 (N_19931,N_18616,N_18268);
nor U19932 (N_19932,N_18193,N_18150);
nand U19933 (N_19933,N_18076,N_18468);
and U19934 (N_19934,N_18081,N_18507);
nor U19935 (N_19935,N_18238,N_18192);
nor U19936 (N_19936,N_18271,N_18777);
xor U19937 (N_19937,N_18183,N_18242);
and U19938 (N_19938,N_18502,N_18479);
xor U19939 (N_19939,N_18010,N_18572);
or U19940 (N_19940,N_18557,N_18658);
nor U19941 (N_19941,N_18222,N_18012);
nand U19942 (N_19942,N_18304,N_18613);
or U19943 (N_19943,N_18256,N_18118);
xor U19944 (N_19944,N_18068,N_18357);
nor U19945 (N_19945,N_18082,N_18998);
xnor U19946 (N_19946,N_18678,N_18834);
nor U19947 (N_19947,N_18420,N_18992);
nor U19948 (N_19948,N_18322,N_18054);
nand U19949 (N_19949,N_18333,N_18578);
nor U19950 (N_19950,N_18584,N_18659);
xnor U19951 (N_19951,N_18860,N_18585);
nand U19952 (N_19952,N_18390,N_18371);
xor U19953 (N_19953,N_18674,N_18975);
or U19954 (N_19954,N_18321,N_18121);
nand U19955 (N_19955,N_18565,N_18691);
nor U19956 (N_19956,N_18738,N_18181);
xor U19957 (N_19957,N_18886,N_18761);
xnor U19958 (N_19958,N_18553,N_18100);
and U19959 (N_19959,N_18592,N_18061);
xnor U19960 (N_19960,N_18427,N_18228);
nand U19961 (N_19961,N_18677,N_18800);
or U19962 (N_19962,N_18244,N_18226);
and U19963 (N_19963,N_18302,N_18690);
nand U19964 (N_19964,N_18301,N_18695);
nand U19965 (N_19965,N_18060,N_18773);
nor U19966 (N_19966,N_18847,N_18349);
and U19967 (N_19967,N_18224,N_18890);
xnor U19968 (N_19968,N_18478,N_18464);
or U19969 (N_19969,N_18271,N_18849);
xnor U19970 (N_19970,N_18733,N_18227);
and U19971 (N_19971,N_18895,N_18518);
xor U19972 (N_19972,N_18493,N_18400);
or U19973 (N_19973,N_18861,N_18911);
xnor U19974 (N_19974,N_18289,N_18435);
and U19975 (N_19975,N_18338,N_18446);
nor U19976 (N_19976,N_18813,N_18944);
or U19977 (N_19977,N_18889,N_18683);
and U19978 (N_19978,N_18500,N_18130);
xor U19979 (N_19979,N_18809,N_18061);
and U19980 (N_19980,N_18783,N_18714);
or U19981 (N_19981,N_18215,N_18624);
xnor U19982 (N_19982,N_18165,N_18239);
nand U19983 (N_19983,N_18497,N_18876);
and U19984 (N_19984,N_18226,N_18306);
nor U19985 (N_19985,N_18654,N_18922);
nor U19986 (N_19986,N_18328,N_18754);
and U19987 (N_19987,N_18830,N_18918);
and U19988 (N_19988,N_18178,N_18572);
nor U19989 (N_19989,N_18322,N_18993);
xor U19990 (N_19990,N_18858,N_18831);
or U19991 (N_19991,N_18909,N_18821);
or U19992 (N_19992,N_18401,N_18822);
or U19993 (N_19993,N_18088,N_18398);
nor U19994 (N_19994,N_18897,N_18856);
or U19995 (N_19995,N_18269,N_18151);
and U19996 (N_19996,N_18830,N_18840);
xnor U19997 (N_19997,N_18478,N_18546);
xor U19998 (N_19998,N_18592,N_18094);
and U19999 (N_19999,N_18780,N_18030);
or U20000 (N_20000,N_19422,N_19997);
xnor U20001 (N_20001,N_19489,N_19419);
or U20002 (N_20002,N_19095,N_19412);
nor U20003 (N_20003,N_19856,N_19801);
nor U20004 (N_20004,N_19667,N_19459);
nand U20005 (N_20005,N_19590,N_19164);
or U20006 (N_20006,N_19349,N_19955);
nand U20007 (N_20007,N_19872,N_19094);
and U20008 (N_20008,N_19807,N_19682);
and U20009 (N_20009,N_19987,N_19659);
nand U20010 (N_20010,N_19298,N_19012);
and U20011 (N_20011,N_19711,N_19900);
and U20012 (N_20012,N_19362,N_19072);
xnor U20013 (N_20013,N_19731,N_19415);
or U20014 (N_20014,N_19594,N_19342);
and U20015 (N_20015,N_19396,N_19181);
xnor U20016 (N_20016,N_19283,N_19739);
nor U20017 (N_20017,N_19702,N_19668);
and U20018 (N_20018,N_19388,N_19505);
nor U20019 (N_20019,N_19448,N_19496);
nand U20020 (N_20020,N_19624,N_19832);
and U20021 (N_20021,N_19289,N_19554);
or U20022 (N_20022,N_19228,N_19381);
nand U20023 (N_20023,N_19983,N_19134);
and U20024 (N_20024,N_19339,N_19100);
xnor U20025 (N_20025,N_19102,N_19860);
or U20026 (N_20026,N_19636,N_19450);
nand U20027 (N_20027,N_19613,N_19064);
xnor U20028 (N_20028,N_19897,N_19548);
nand U20029 (N_20029,N_19846,N_19272);
or U20030 (N_20030,N_19268,N_19082);
and U20031 (N_20031,N_19165,N_19648);
nor U20032 (N_20032,N_19942,N_19681);
nand U20033 (N_20033,N_19603,N_19537);
and U20034 (N_20034,N_19553,N_19794);
xor U20035 (N_20035,N_19720,N_19823);
or U20036 (N_20036,N_19107,N_19136);
or U20037 (N_20037,N_19741,N_19157);
nand U20038 (N_20038,N_19347,N_19340);
nor U20039 (N_20039,N_19247,N_19067);
nor U20040 (N_20040,N_19189,N_19217);
nand U20041 (N_20041,N_19299,N_19059);
nand U20042 (N_20042,N_19907,N_19356);
xor U20043 (N_20043,N_19203,N_19457);
nor U20044 (N_20044,N_19111,N_19454);
nand U20045 (N_20045,N_19025,N_19416);
and U20046 (N_20046,N_19243,N_19526);
xor U20047 (N_20047,N_19529,N_19176);
nand U20048 (N_20048,N_19475,N_19658);
nand U20049 (N_20049,N_19894,N_19026);
nor U20050 (N_20050,N_19953,N_19976);
nand U20051 (N_20051,N_19015,N_19940);
nor U20052 (N_20052,N_19568,N_19782);
and U20053 (N_20053,N_19112,N_19844);
xnor U20054 (N_20054,N_19225,N_19132);
nor U20055 (N_20055,N_19487,N_19127);
or U20056 (N_20056,N_19979,N_19319);
or U20057 (N_20057,N_19871,N_19401);
or U20058 (N_20058,N_19742,N_19806);
nand U20059 (N_20059,N_19790,N_19210);
or U20060 (N_20060,N_19331,N_19128);
xnor U20061 (N_20061,N_19383,N_19106);
nand U20062 (N_20062,N_19758,N_19022);
nor U20063 (N_20063,N_19508,N_19586);
or U20064 (N_20064,N_19382,N_19995);
and U20065 (N_20065,N_19889,N_19617);
and U20066 (N_20066,N_19596,N_19558);
nor U20067 (N_20067,N_19536,N_19560);
nand U20068 (N_20068,N_19484,N_19476);
nand U20069 (N_20069,N_19559,N_19192);
xor U20070 (N_20070,N_19267,N_19923);
nand U20071 (N_20071,N_19928,N_19737);
xor U20072 (N_20072,N_19992,N_19566);
xnor U20073 (N_20073,N_19110,N_19108);
and U20074 (N_20074,N_19611,N_19389);
nor U20075 (N_20075,N_19302,N_19926);
nor U20076 (N_20076,N_19716,N_19839);
and U20077 (N_20077,N_19543,N_19732);
or U20078 (N_20078,N_19403,N_19241);
xnor U20079 (N_20079,N_19501,N_19320);
and U20080 (N_20080,N_19744,N_19514);
nand U20081 (N_20081,N_19104,N_19088);
nor U20082 (N_20082,N_19982,N_19256);
and U20083 (N_20083,N_19723,N_19993);
and U20084 (N_20084,N_19056,N_19701);
and U20085 (N_20085,N_19273,N_19162);
nor U20086 (N_20086,N_19375,N_19809);
nor U20087 (N_20087,N_19713,N_19142);
nor U20088 (N_20088,N_19138,N_19936);
and U20089 (N_20089,N_19421,N_19405);
and U20090 (N_20090,N_19527,N_19290);
or U20091 (N_20091,N_19666,N_19369);
or U20092 (N_20092,N_19639,N_19277);
or U20093 (N_20093,N_19146,N_19291);
and U20094 (N_20094,N_19266,N_19365);
nand U20095 (N_20095,N_19540,N_19891);
xnor U20096 (N_20096,N_19318,N_19530);
xnor U20097 (N_20097,N_19629,N_19929);
and U20098 (N_20098,N_19214,N_19429);
nor U20099 (N_20099,N_19721,N_19893);
nand U20100 (N_20100,N_19948,N_19444);
xnor U20101 (N_20101,N_19949,N_19002);
and U20102 (N_20102,N_19439,N_19227);
nand U20103 (N_20103,N_19129,N_19812);
nand U20104 (N_20104,N_19981,N_19951);
nand U20105 (N_20105,N_19335,N_19646);
nor U20106 (N_20106,N_19877,N_19883);
nor U20107 (N_20107,N_19061,N_19557);
nor U20108 (N_20108,N_19715,N_19441);
nand U20109 (N_20109,N_19627,N_19467);
nor U20110 (N_20110,N_19609,N_19148);
nand U20111 (N_20111,N_19588,N_19163);
and U20112 (N_20112,N_19699,N_19610);
nand U20113 (N_20113,N_19927,N_19509);
xor U20114 (N_20114,N_19519,N_19688);
and U20115 (N_20115,N_19654,N_19240);
and U20116 (N_20116,N_19262,N_19756);
nor U20117 (N_20117,N_19994,N_19925);
nand U20118 (N_20118,N_19888,N_19235);
nor U20119 (N_20119,N_19763,N_19269);
xor U20120 (N_20120,N_19196,N_19524);
or U20121 (N_20121,N_19647,N_19151);
and U20122 (N_20122,N_19873,N_19140);
nand U20123 (N_20123,N_19550,N_19071);
or U20124 (N_20124,N_19348,N_19954);
or U20125 (N_20125,N_19886,N_19885);
xor U20126 (N_20126,N_19602,N_19865);
and U20127 (N_20127,N_19297,N_19895);
or U20128 (N_20128,N_19820,N_19119);
nor U20129 (N_20129,N_19686,N_19292);
nor U20130 (N_20130,N_19676,N_19915);
nor U20131 (N_20131,N_19837,N_19670);
nand U20132 (N_20132,N_19693,N_19638);
and U20133 (N_20133,N_19921,N_19169);
and U20134 (N_20134,N_19117,N_19447);
and U20135 (N_20135,N_19551,N_19202);
nor U20136 (N_20136,N_19781,N_19041);
nor U20137 (N_20137,N_19314,N_19188);
xor U20138 (N_20138,N_19078,N_19472);
nand U20139 (N_20139,N_19653,N_19433);
and U20140 (N_20140,N_19764,N_19321);
and U20141 (N_20141,N_19248,N_19974);
and U20142 (N_20142,N_19743,N_19988);
nor U20143 (N_20143,N_19174,N_19958);
xnor U20144 (N_20144,N_19735,N_19710);
and U20145 (N_20145,N_19555,N_19947);
and U20146 (N_20146,N_19355,N_19101);
xnor U20147 (N_20147,N_19473,N_19480);
nor U20148 (N_20148,N_19400,N_19696);
or U20149 (N_20149,N_19135,N_19506);
xnor U20150 (N_20150,N_19023,N_19191);
or U20151 (N_20151,N_19058,N_19284);
and U20152 (N_20152,N_19991,N_19694);
and U20153 (N_20153,N_19168,N_19734);
nor U20154 (N_20154,N_19036,N_19068);
nand U20155 (N_20155,N_19680,N_19034);
nor U20156 (N_20156,N_19249,N_19295);
nor U20157 (N_20157,N_19829,N_19231);
and U20158 (N_20158,N_19391,N_19154);
or U20159 (N_20159,N_19255,N_19152);
xor U20160 (N_20160,N_19600,N_19999);
nor U20161 (N_20161,N_19470,N_19166);
nor U20162 (N_20162,N_19673,N_19826);
nor U20163 (N_20163,N_19697,N_19625);
nand U20164 (N_20164,N_19853,N_19591);
and U20165 (N_20165,N_19069,N_19322);
and U20166 (N_20166,N_19155,N_19493);
or U20167 (N_20167,N_19063,N_19941);
nor U20168 (N_20168,N_19963,N_19229);
xor U20169 (N_20169,N_19533,N_19324);
and U20170 (N_20170,N_19308,N_19413);
xnor U20171 (N_20171,N_19222,N_19521);
and U20172 (N_20172,N_19316,N_19462);
or U20173 (N_20173,N_19011,N_19628);
nor U20174 (N_20174,N_19193,N_19035);
nand U20175 (N_20175,N_19516,N_19884);
nor U20176 (N_20176,N_19712,N_19817);
nand U20177 (N_20177,N_19728,N_19455);
nor U20178 (N_20178,N_19150,N_19153);
and U20179 (N_20179,N_19626,N_19642);
and U20180 (N_20180,N_19254,N_19286);
or U20181 (N_20181,N_19213,N_19180);
and U20182 (N_20182,N_19705,N_19387);
xnor U20183 (N_20183,N_19097,N_19523);
xor U20184 (N_20184,N_19931,N_19131);
nand U20185 (N_20185,N_19280,N_19589);
or U20186 (N_20186,N_19683,N_19838);
and U20187 (N_20187,N_19440,N_19869);
or U20188 (N_20188,N_19851,N_19330);
nand U20189 (N_20189,N_19386,N_19468);
nand U20190 (N_20190,N_19261,N_19799);
nand U20191 (N_20191,N_19260,N_19512);
xor U20192 (N_20192,N_19460,N_19664);
nand U20193 (N_20193,N_19236,N_19679);
nand U20194 (N_20194,N_19288,N_19998);
nor U20195 (N_20195,N_19704,N_19973);
xnor U20196 (N_20196,N_19209,N_19752);
xnor U20197 (N_20197,N_19504,N_19377);
xor U20198 (N_20198,N_19394,N_19099);
xnor U20199 (N_20199,N_19374,N_19479);
or U20200 (N_20200,N_19436,N_19096);
nand U20201 (N_20201,N_19488,N_19113);
nor U20202 (N_20202,N_19633,N_19881);
nand U20203 (N_20203,N_19825,N_19417);
or U20204 (N_20204,N_19546,N_19730);
and U20205 (N_20205,N_19592,N_19390);
nor U20206 (N_20206,N_19380,N_19147);
xnor U20207 (N_20207,N_19052,N_19677);
or U20208 (N_20208,N_19919,N_19170);
and U20209 (N_20209,N_19087,N_19569);
nor U20210 (N_20210,N_19746,N_19379);
and U20211 (N_20211,N_19378,N_19587);
nand U20212 (N_20212,N_19778,N_19616);
or U20213 (N_20213,N_19896,N_19274);
and U20214 (N_20214,N_19327,N_19874);
or U20215 (N_20215,N_19828,N_19840);
and U20216 (N_20216,N_19779,N_19552);
xnor U20217 (N_20217,N_19221,N_19021);
xor U20218 (N_20218,N_19054,N_19599);
xnor U20219 (N_20219,N_19336,N_19880);
nor U20220 (N_20220,N_19797,N_19738);
and U20221 (N_20221,N_19309,N_19343);
or U20222 (N_20222,N_19768,N_19703);
or U20223 (N_20223,N_19250,N_19430);
xnor U20224 (N_20224,N_19195,N_19033);
nand U20225 (N_20225,N_19252,N_19464);
and U20226 (N_20226,N_19952,N_19622);
nand U20227 (N_20227,N_19845,N_19232);
xor U20228 (N_20228,N_19120,N_19811);
xor U20229 (N_20229,N_19143,N_19350);
nor U20230 (N_20230,N_19967,N_19352);
xnor U20231 (N_20231,N_19635,N_19545);
or U20232 (N_20232,N_19939,N_19172);
and U20233 (N_20233,N_19632,N_19815);
or U20234 (N_20234,N_19990,N_19452);
nand U20235 (N_20235,N_19597,N_19215);
or U20236 (N_20236,N_19507,N_19774);
xnor U20237 (N_20237,N_19373,N_19497);
nand U20238 (N_20238,N_19050,N_19714);
and U20239 (N_20239,N_19208,N_19086);
nand U20240 (N_20240,N_19736,N_19282);
xnor U20241 (N_20241,N_19822,N_19031);
and U20242 (N_20242,N_19899,N_19834);
nor U20243 (N_20243,N_19565,N_19698);
and U20244 (N_20244,N_19511,N_19662);
or U20245 (N_20245,N_19233,N_19017);
or U20246 (N_20246,N_19158,N_19357);
nand U20247 (N_20247,N_19466,N_19385);
or U20248 (N_20248,N_19027,N_19259);
or U20249 (N_20249,N_19751,N_19079);
xnor U20250 (N_20250,N_19438,N_19453);
nand U20251 (N_20251,N_19244,N_19014);
nor U20252 (N_20252,N_19902,N_19315);
nand U20253 (N_20253,N_19171,N_19606);
or U20254 (N_20254,N_19787,N_19426);
nor U20255 (N_20255,N_19841,N_19006);
nor U20256 (N_20256,N_19125,N_19098);
or U20257 (N_20257,N_19449,N_19264);
nor U20258 (N_20258,N_19862,N_19062);
and U20259 (N_20259,N_19561,N_19223);
nor U20260 (N_20260,N_19788,N_19535);
or U20261 (N_20261,N_19525,N_19490);
nor U20262 (N_20262,N_19855,N_19605);
nor U20263 (N_20263,N_19910,N_19753);
and U20264 (N_20264,N_19904,N_19916);
and U20265 (N_20265,N_19325,N_19534);
nand U20266 (N_20266,N_19937,N_19692);
and U20267 (N_20267,N_19858,N_19968);
nor U20268 (N_20268,N_19372,N_19531);
and U20269 (N_20269,N_19984,N_19371);
xor U20270 (N_20270,N_19177,N_19532);
xnor U20271 (N_20271,N_19908,N_19695);
or U20272 (N_20272,N_19528,N_19366);
nor U20273 (N_20273,N_19133,N_19866);
xor U20274 (N_20274,N_19124,N_19760);
xor U20275 (N_20275,N_19691,N_19344);
or U20276 (N_20276,N_19404,N_19007);
or U20277 (N_20277,N_19930,N_19934);
nand U20278 (N_20278,N_19144,N_19123);
nand U20279 (N_20279,N_19541,N_19492);
or U20280 (N_20280,N_19685,N_19199);
or U20281 (N_20281,N_19257,N_19337);
and U20282 (N_20282,N_19796,N_19271);
nor U20283 (N_20283,N_19542,N_19969);
xnor U20284 (N_20284,N_19009,N_19620);
xor U20285 (N_20285,N_19769,N_19808);
xor U20286 (N_20286,N_19878,N_19194);
xnor U20287 (N_20287,N_19573,N_19848);
and U20288 (N_20288,N_19043,N_19200);
or U20289 (N_20289,N_19234,N_19707);
xnor U20290 (N_20290,N_19898,N_19019);
and U20291 (N_20291,N_19503,N_19367);
or U20292 (N_20292,N_19065,N_19598);
or U20293 (N_20293,N_19329,N_19206);
nand U20294 (N_20294,N_19918,N_19748);
xor U20295 (N_20295,N_19328,N_19402);
xor U20296 (N_20296,N_19471,N_19296);
and U20297 (N_20297,N_19092,N_19965);
nand U20298 (N_20298,N_19219,N_19080);
nor U20299 (N_20299,N_19793,N_19830);
and U20300 (N_20300,N_19184,N_19463);
nand U20301 (N_20301,N_19049,N_19724);
and U20302 (N_20302,N_19814,N_19018);
nor U20303 (N_20303,N_19323,N_19118);
and U20304 (N_20304,N_19957,N_19777);
nor U20305 (N_20305,N_19601,N_19945);
or U20306 (N_20306,N_19414,N_19474);
or U20307 (N_20307,N_19001,N_19085);
nor U20308 (N_20308,N_19305,N_19420);
or U20309 (N_20309,N_19495,N_19310);
or U20310 (N_20310,N_19428,N_19105);
or U20311 (N_20311,N_19513,N_19813);
nand U20312 (N_20312,N_19985,N_19418);
nor U20313 (N_20313,N_19042,N_19115);
nor U20314 (N_20314,N_19595,N_19334);
xor U20315 (N_20315,N_19640,N_19795);
nor U20316 (N_20316,N_19376,N_19384);
and U20317 (N_20317,N_19037,N_19689);
nor U20318 (N_20318,N_19810,N_19766);
and U20319 (N_20319,N_19996,N_19109);
nand U20320 (N_20320,N_19564,N_19913);
and U20321 (N_20321,N_19649,N_19581);
xnor U20322 (N_20322,N_19634,N_19585);
and U20323 (N_20323,N_19345,N_19719);
nand U20324 (N_20324,N_19656,N_19665);
nand U20325 (N_20325,N_19178,N_19024);
xor U20326 (N_20326,N_19045,N_19427);
and U20327 (N_20327,N_19368,N_19580);
or U20328 (N_20328,N_19563,N_19451);
and U20329 (N_20329,N_19425,N_19818);
nand U20330 (N_20330,N_19197,N_19126);
nand U20331 (N_20331,N_19246,N_19749);
xor U20332 (N_20332,N_19040,N_19663);
nor U20333 (N_20333,N_19819,N_19767);
nand U20334 (N_20334,N_19762,N_19167);
nand U20335 (N_20335,N_19909,N_19776);
nand U20336 (N_20336,N_19944,N_19986);
or U20337 (N_20337,N_19718,N_19631);
xnor U20338 (N_20338,N_19226,N_19161);
nand U20339 (N_20339,N_19149,N_19847);
nand U20340 (N_20340,N_19029,N_19179);
or U20341 (N_20341,N_19090,N_19623);
nor U20342 (N_20342,N_19081,N_19783);
nand U20343 (N_20343,N_19674,N_19575);
nand U20344 (N_20344,N_19791,N_19446);
xnor U20345 (N_20345,N_19160,N_19057);
or U20346 (N_20346,N_19786,N_19461);
nand U20347 (N_20347,N_19313,N_19970);
and U20348 (N_20348,N_19351,N_19130);
nand U20349 (N_20349,N_19905,N_19630);
nand U20350 (N_20350,N_19518,N_19835);
or U20351 (N_20351,N_19864,N_19827);
and U20352 (N_20352,N_19083,N_19964);
and U20353 (N_20353,N_19842,N_19423);
xor U20354 (N_20354,N_19747,N_19353);
nand U20355 (N_20355,N_19091,N_19145);
and U20356 (N_20356,N_19047,N_19684);
and U20357 (N_20357,N_19879,N_19977);
xnor U20358 (N_20358,N_19887,N_19854);
xor U20359 (N_20359,N_19914,N_19116);
or U20360 (N_20360,N_19486,N_19122);
nor U20361 (N_20361,N_19075,N_19556);
xor U20362 (N_20362,N_19185,N_19481);
or U20363 (N_20363,N_19579,N_19643);
nand U20364 (N_20364,N_19392,N_19645);
or U20365 (N_20365,N_19359,N_19700);
nor U20366 (N_20366,N_19275,N_19771);
and U20367 (N_20367,N_19139,N_19708);
and U20368 (N_20368,N_19103,N_19070);
xor U20369 (N_20369,N_19584,N_19201);
and U20370 (N_20370,N_19445,N_19077);
xnor U20371 (N_20371,N_19867,N_19943);
and U20372 (N_20372,N_19972,N_19615);
or U20373 (N_20373,N_19824,N_19831);
and U20374 (N_20374,N_19607,N_19912);
and U20375 (N_20375,N_19477,N_19121);
and U20376 (N_20376,N_19836,N_19303);
and U20377 (N_20377,N_19230,N_19499);
xnor U20378 (N_20378,N_19770,N_19924);
nor U20379 (N_20379,N_19044,N_19725);
nand U20380 (N_20380,N_19204,N_19652);
and U20381 (N_20381,N_19935,N_19661);
or U20382 (N_20382,N_19861,N_19570);
and U20383 (N_20383,N_19784,N_19619);
and U20384 (N_20384,N_19046,N_19458);
and U20385 (N_20385,N_19242,N_19522);
or U20386 (N_20386,N_19706,N_19003);
and U20387 (N_20387,N_19265,N_19572);
nor U20388 (N_20388,N_19276,N_19859);
and U20389 (N_20389,N_19432,N_19051);
nor U20390 (N_20390,N_19443,N_19510);
nor U20391 (N_20391,N_19053,N_19821);
nor U20392 (N_20392,N_19870,N_19114);
nor U20393 (N_20393,N_19759,N_19055);
xor U20394 (N_20394,N_19141,N_19346);
nor U20395 (N_20395,N_19773,N_19901);
and U20396 (N_20396,N_19358,N_19364);
nor U20397 (N_20397,N_19338,N_19576);
nand U20398 (N_20398,N_19772,N_19205);
or U20399 (N_20399,N_19956,N_19326);
and U20400 (N_20400,N_19482,N_19483);
nor U20401 (N_20401,N_19198,N_19032);
and U20402 (N_20402,N_19363,N_19220);
xnor U20403 (N_20403,N_19816,N_19183);
nor U20404 (N_20404,N_19175,N_19669);
and U20405 (N_20405,N_19442,N_19173);
xor U20406 (N_20406,N_19843,N_19675);
and U20407 (N_20407,N_19549,N_19360);
nand U20408 (N_20408,N_19013,N_19039);
and U20409 (N_20409,N_19048,N_19727);
nand U20410 (N_20410,N_19644,N_19574);
nand U20411 (N_20411,N_19301,N_19798);
or U20412 (N_20412,N_19938,N_19437);
or U20413 (N_20413,N_19745,N_19410);
or U20414 (N_20414,N_19000,N_19137);
xor U20415 (N_20415,N_19270,N_19008);
and U20416 (N_20416,N_19792,N_19186);
xnor U20417 (N_20417,N_19539,N_19399);
nor U20418 (N_20418,N_19785,N_19370);
or U20419 (N_20419,N_19805,N_19754);
nor U20420 (N_20420,N_19671,N_19655);
and U20421 (N_20421,N_19239,N_19946);
xnor U20422 (N_20422,N_19515,N_19397);
nand U20423 (N_20423,N_19621,N_19311);
nor U20424 (N_20424,N_19030,N_19517);
nand U20425 (N_20425,N_19038,N_19567);
nand U20426 (N_20426,N_19975,N_19190);
xor U20427 (N_20427,N_19074,N_19593);
and U20428 (N_20428,N_19850,N_19717);
or U20429 (N_20429,N_19398,N_19978);
nand U20430 (N_20430,N_19852,N_19278);
or U20431 (N_20431,N_19361,N_19612);
nor U20432 (N_20432,N_19775,N_19757);
or U20433 (N_20433,N_19538,N_19733);
or U20434 (N_20434,N_19604,N_19804);
or U20435 (N_20435,N_19657,N_19089);
nor U20436 (N_20436,N_19395,N_19803);
and U20437 (N_20437,N_19156,N_19212);
nor U20438 (N_20438,N_19906,N_19312);
nand U20439 (N_20439,N_19980,N_19755);
xnor U20440 (N_20440,N_19187,N_19224);
xor U20441 (N_20441,N_19618,N_19740);
nand U20442 (N_20442,N_19258,N_19253);
nand U20443 (N_20443,N_19304,N_19608);
and U20444 (N_20444,N_19502,N_19424);
nor U20445 (N_20445,N_19285,N_19307);
or U20446 (N_20446,N_19076,N_19294);
xor U20447 (N_20447,N_19498,N_19409);
nand U20448 (N_20448,N_19933,N_19494);
and U20449 (N_20449,N_19571,N_19849);
xnor U20450 (N_20450,N_19500,N_19911);
nand U20451 (N_20451,N_19060,N_19750);
nand U20452 (N_20452,N_19182,N_19004);
nand U20453 (N_20453,N_19465,N_19435);
nand U20454 (N_20454,N_19800,N_19614);
and U20455 (N_20455,N_19010,N_19456);
nor U20456 (N_20456,N_19237,N_19651);
and U20457 (N_20457,N_19582,N_19765);
or U20458 (N_20458,N_19020,N_19341);
or U20459 (N_20459,N_19962,N_19971);
nand U20460 (N_20460,N_19729,N_19577);
and U20461 (N_20461,N_19868,N_19961);
or U20462 (N_20462,N_19761,N_19709);
xor U20463 (N_20463,N_19917,N_19317);
nor U20464 (N_20464,N_19238,N_19245);
nor U20465 (N_20465,N_19722,N_19028);
nand U20466 (N_20466,N_19005,N_19875);
or U20467 (N_20467,N_19332,N_19084);
xnor U20468 (N_20468,N_19406,N_19251);
or U20469 (N_20469,N_19890,N_19411);
nand U20470 (N_20470,N_19922,N_19892);
or U20471 (N_20471,N_19690,N_19279);
nor U20472 (N_20472,N_19687,N_19434);
and U20473 (N_20473,N_19354,N_19520);
xor U20474 (N_20474,N_19780,N_19263);
nor U20475 (N_20475,N_19547,N_19960);
xor U20476 (N_20476,N_19583,N_19431);
xnor U20477 (N_20477,N_19073,N_19408);
nand U20478 (N_20478,N_19966,N_19469);
nand U20479 (N_20479,N_19066,N_19578);
xnor U20480 (N_20480,N_19407,N_19989);
nand U20481 (N_20481,N_19950,N_19650);
xor U20482 (N_20482,N_19544,N_19882);
xor U20483 (N_20483,N_19789,N_19491);
and U20484 (N_20484,N_19287,N_19932);
xor U20485 (N_20485,N_19876,N_19959);
nand U20486 (N_20486,N_19207,N_19293);
nand U20487 (N_20487,N_19281,N_19093);
xor U20488 (N_20488,N_19211,N_19306);
or U20489 (N_20489,N_19562,N_19478);
and U20490 (N_20490,N_19726,N_19920);
and U20491 (N_20491,N_19637,N_19903);
nor U20492 (N_20492,N_19218,N_19216);
nand U20493 (N_20493,N_19857,N_19802);
and U20494 (N_20494,N_19641,N_19300);
xnor U20495 (N_20495,N_19833,N_19678);
or U20496 (N_20496,N_19159,N_19393);
and U20497 (N_20497,N_19485,N_19333);
nor U20498 (N_20498,N_19863,N_19660);
nor U20499 (N_20499,N_19672,N_19016);
nor U20500 (N_20500,N_19894,N_19867);
or U20501 (N_20501,N_19239,N_19268);
or U20502 (N_20502,N_19294,N_19318);
and U20503 (N_20503,N_19606,N_19582);
and U20504 (N_20504,N_19850,N_19422);
nor U20505 (N_20505,N_19320,N_19427);
nor U20506 (N_20506,N_19518,N_19326);
or U20507 (N_20507,N_19816,N_19227);
xnor U20508 (N_20508,N_19871,N_19648);
nor U20509 (N_20509,N_19095,N_19634);
nand U20510 (N_20510,N_19583,N_19444);
xnor U20511 (N_20511,N_19849,N_19397);
or U20512 (N_20512,N_19773,N_19116);
nand U20513 (N_20513,N_19859,N_19485);
or U20514 (N_20514,N_19605,N_19347);
nor U20515 (N_20515,N_19105,N_19336);
xor U20516 (N_20516,N_19312,N_19099);
nand U20517 (N_20517,N_19028,N_19288);
xnor U20518 (N_20518,N_19080,N_19918);
nand U20519 (N_20519,N_19140,N_19938);
xnor U20520 (N_20520,N_19522,N_19382);
and U20521 (N_20521,N_19374,N_19888);
nor U20522 (N_20522,N_19959,N_19556);
nand U20523 (N_20523,N_19944,N_19102);
xnor U20524 (N_20524,N_19604,N_19320);
nor U20525 (N_20525,N_19787,N_19969);
or U20526 (N_20526,N_19056,N_19434);
xor U20527 (N_20527,N_19678,N_19399);
or U20528 (N_20528,N_19932,N_19455);
and U20529 (N_20529,N_19125,N_19604);
nor U20530 (N_20530,N_19747,N_19612);
xor U20531 (N_20531,N_19939,N_19993);
or U20532 (N_20532,N_19479,N_19197);
xnor U20533 (N_20533,N_19684,N_19731);
xnor U20534 (N_20534,N_19656,N_19892);
or U20535 (N_20535,N_19785,N_19163);
and U20536 (N_20536,N_19211,N_19453);
xor U20537 (N_20537,N_19104,N_19879);
nor U20538 (N_20538,N_19513,N_19038);
xor U20539 (N_20539,N_19675,N_19022);
nand U20540 (N_20540,N_19115,N_19665);
or U20541 (N_20541,N_19929,N_19899);
xor U20542 (N_20542,N_19215,N_19466);
nand U20543 (N_20543,N_19997,N_19790);
or U20544 (N_20544,N_19359,N_19609);
nor U20545 (N_20545,N_19048,N_19338);
nand U20546 (N_20546,N_19126,N_19694);
xnor U20547 (N_20547,N_19340,N_19221);
or U20548 (N_20548,N_19182,N_19864);
nand U20549 (N_20549,N_19919,N_19913);
nand U20550 (N_20550,N_19126,N_19215);
nor U20551 (N_20551,N_19518,N_19551);
nand U20552 (N_20552,N_19196,N_19890);
xnor U20553 (N_20553,N_19114,N_19123);
xor U20554 (N_20554,N_19912,N_19815);
nand U20555 (N_20555,N_19570,N_19886);
or U20556 (N_20556,N_19908,N_19655);
xnor U20557 (N_20557,N_19571,N_19479);
and U20558 (N_20558,N_19630,N_19316);
nor U20559 (N_20559,N_19699,N_19379);
nand U20560 (N_20560,N_19093,N_19820);
nand U20561 (N_20561,N_19877,N_19344);
nand U20562 (N_20562,N_19638,N_19980);
xnor U20563 (N_20563,N_19103,N_19334);
and U20564 (N_20564,N_19403,N_19842);
xnor U20565 (N_20565,N_19697,N_19270);
nand U20566 (N_20566,N_19736,N_19776);
or U20567 (N_20567,N_19511,N_19430);
or U20568 (N_20568,N_19013,N_19327);
or U20569 (N_20569,N_19854,N_19676);
nor U20570 (N_20570,N_19719,N_19931);
nand U20571 (N_20571,N_19102,N_19728);
and U20572 (N_20572,N_19402,N_19764);
nor U20573 (N_20573,N_19485,N_19647);
and U20574 (N_20574,N_19337,N_19325);
and U20575 (N_20575,N_19372,N_19625);
nor U20576 (N_20576,N_19503,N_19768);
nand U20577 (N_20577,N_19718,N_19323);
xnor U20578 (N_20578,N_19823,N_19416);
nand U20579 (N_20579,N_19275,N_19356);
or U20580 (N_20580,N_19338,N_19876);
nor U20581 (N_20581,N_19152,N_19545);
and U20582 (N_20582,N_19881,N_19832);
nand U20583 (N_20583,N_19194,N_19382);
or U20584 (N_20584,N_19192,N_19744);
nor U20585 (N_20585,N_19130,N_19898);
and U20586 (N_20586,N_19629,N_19974);
xnor U20587 (N_20587,N_19426,N_19148);
xor U20588 (N_20588,N_19170,N_19009);
and U20589 (N_20589,N_19333,N_19501);
or U20590 (N_20590,N_19529,N_19847);
nand U20591 (N_20591,N_19226,N_19112);
xnor U20592 (N_20592,N_19001,N_19843);
and U20593 (N_20593,N_19860,N_19226);
nor U20594 (N_20594,N_19208,N_19966);
or U20595 (N_20595,N_19989,N_19789);
or U20596 (N_20596,N_19509,N_19483);
xnor U20597 (N_20597,N_19892,N_19513);
nor U20598 (N_20598,N_19545,N_19281);
xnor U20599 (N_20599,N_19499,N_19031);
and U20600 (N_20600,N_19651,N_19467);
nand U20601 (N_20601,N_19019,N_19775);
xnor U20602 (N_20602,N_19409,N_19386);
or U20603 (N_20603,N_19814,N_19181);
nand U20604 (N_20604,N_19104,N_19270);
nand U20605 (N_20605,N_19347,N_19198);
nor U20606 (N_20606,N_19812,N_19596);
xnor U20607 (N_20607,N_19664,N_19170);
and U20608 (N_20608,N_19475,N_19886);
and U20609 (N_20609,N_19524,N_19205);
xor U20610 (N_20610,N_19261,N_19768);
xor U20611 (N_20611,N_19180,N_19118);
nand U20612 (N_20612,N_19170,N_19781);
xor U20613 (N_20613,N_19473,N_19277);
xor U20614 (N_20614,N_19483,N_19417);
xor U20615 (N_20615,N_19651,N_19158);
nor U20616 (N_20616,N_19116,N_19892);
nand U20617 (N_20617,N_19315,N_19006);
nor U20618 (N_20618,N_19057,N_19844);
or U20619 (N_20619,N_19988,N_19070);
or U20620 (N_20620,N_19778,N_19914);
nand U20621 (N_20621,N_19535,N_19635);
or U20622 (N_20622,N_19563,N_19195);
nand U20623 (N_20623,N_19389,N_19713);
or U20624 (N_20624,N_19177,N_19570);
nand U20625 (N_20625,N_19860,N_19372);
nand U20626 (N_20626,N_19997,N_19394);
nand U20627 (N_20627,N_19779,N_19382);
nor U20628 (N_20628,N_19759,N_19033);
nor U20629 (N_20629,N_19675,N_19201);
xor U20630 (N_20630,N_19392,N_19277);
and U20631 (N_20631,N_19120,N_19861);
and U20632 (N_20632,N_19096,N_19064);
nand U20633 (N_20633,N_19769,N_19658);
nand U20634 (N_20634,N_19589,N_19234);
or U20635 (N_20635,N_19154,N_19755);
xor U20636 (N_20636,N_19875,N_19174);
or U20637 (N_20637,N_19353,N_19577);
nor U20638 (N_20638,N_19673,N_19044);
nor U20639 (N_20639,N_19484,N_19863);
and U20640 (N_20640,N_19993,N_19558);
and U20641 (N_20641,N_19295,N_19632);
xor U20642 (N_20642,N_19945,N_19870);
or U20643 (N_20643,N_19799,N_19327);
and U20644 (N_20644,N_19555,N_19538);
xnor U20645 (N_20645,N_19974,N_19261);
or U20646 (N_20646,N_19619,N_19285);
nor U20647 (N_20647,N_19909,N_19084);
nor U20648 (N_20648,N_19344,N_19597);
nand U20649 (N_20649,N_19549,N_19035);
nor U20650 (N_20650,N_19161,N_19151);
xnor U20651 (N_20651,N_19892,N_19697);
or U20652 (N_20652,N_19531,N_19020);
nor U20653 (N_20653,N_19059,N_19270);
nor U20654 (N_20654,N_19046,N_19597);
or U20655 (N_20655,N_19447,N_19938);
and U20656 (N_20656,N_19749,N_19551);
nor U20657 (N_20657,N_19818,N_19501);
nor U20658 (N_20658,N_19938,N_19579);
and U20659 (N_20659,N_19911,N_19964);
or U20660 (N_20660,N_19926,N_19709);
nor U20661 (N_20661,N_19973,N_19920);
nand U20662 (N_20662,N_19958,N_19035);
or U20663 (N_20663,N_19841,N_19592);
nand U20664 (N_20664,N_19499,N_19223);
and U20665 (N_20665,N_19064,N_19460);
xor U20666 (N_20666,N_19723,N_19880);
nor U20667 (N_20667,N_19977,N_19694);
nand U20668 (N_20668,N_19672,N_19703);
nor U20669 (N_20669,N_19295,N_19485);
nand U20670 (N_20670,N_19458,N_19400);
xnor U20671 (N_20671,N_19807,N_19384);
nand U20672 (N_20672,N_19138,N_19671);
or U20673 (N_20673,N_19259,N_19093);
and U20674 (N_20674,N_19488,N_19889);
nor U20675 (N_20675,N_19260,N_19714);
nor U20676 (N_20676,N_19807,N_19023);
nor U20677 (N_20677,N_19173,N_19684);
nor U20678 (N_20678,N_19669,N_19412);
nor U20679 (N_20679,N_19642,N_19077);
and U20680 (N_20680,N_19818,N_19701);
or U20681 (N_20681,N_19763,N_19254);
or U20682 (N_20682,N_19348,N_19658);
or U20683 (N_20683,N_19818,N_19823);
and U20684 (N_20684,N_19703,N_19029);
nor U20685 (N_20685,N_19767,N_19021);
nand U20686 (N_20686,N_19256,N_19949);
nor U20687 (N_20687,N_19352,N_19581);
nor U20688 (N_20688,N_19535,N_19163);
nor U20689 (N_20689,N_19455,N_19038);
nor U20690 (N_20690,N_19212,N_19199);
nand U20691 (N_20691,N_19235,N_19393);
nand U20692 (N_20692,N_19279,N_19455);
nand U20693 (N_20693,N_19524,N_19134);
or U20694 (N_20694,N_19492,N_19448);
and U20695 (N_20695,N_19506,N_19564);
and U20696 (N_20696,N_19457,N_19789);
xor U20697 (N_20697,N_19302,N_19951);
or U20698 (N_20698,N_19877,N_19479);
nor U20699 (N_20699,N_19481,N_19877);
or U20700 (N_20700,N_19109,N_19074);
and U20701 (N_20701,N_19841,N_19333);
or U20702 (N_20702,N_19100,N_19568);
xor U20703 (N_20703,N_19333,N_19405);
nand U20704 (N_20704,N_19901,N_19019);
nand U20705 (N_20705,N_19356,N_19461);
nand U20706 (N_20706,N_19582,N_19179);
and U20707 (N_20707,N_19514,N_19446);
xor U20708 (N_20708,N_19110,N_19298);
nor U20709 (N_20709,N_19632,N_19547);
or U20710 (N_20710,N_19370,N_19718);
nor U20711 (N_20711,N_19346,N_19146);
xnor U20712 (N_20712,N_19360,N_19641);
nor U20713 (N_20713,N_19857,N_19787);
or U20714 (N_20714,N_19281,N_19237);
or U20715 (N_20715,N_19877,N_19060);
nand U20716 (N_20716,N_19320,N_19035);
or U20717 (N_20717,N_19743,N_19932);
xnor U20718 (N_20718,N_19669,N_19129);
or U20719 (N_20719,N_19827,N_19464);
xor U20720 (N_20720,N_19920,N_19680);
nand U20721 (N_20721,N_19075,N_19601);
nand U20722 (N_20722,N_19304,N_19015);
nand U20723 (N_20723,N_19977,N_19347);
nand U20724 (N_20724,N_19509,N_19527);
nand U20725 (N_20725,N_19327,N_19255);
xor U20726 (N_20726,N_19950,N_19500);
or U20727 (N_20727,N_19689,N_19245);
and U20728 (N_20728,N_19193,N_19925);
xor U20729 (N_20729,N_19590,N_19929);
or U20730 (N_20730,N_19045,N_19192);
xnor U20731 (N_20731,N_19743,N_19873);
nor U20732 (N_20732,N_19979,N_19698);
xor U20733 (N_20733,N_19961,N_19166);
xnor U20734 (N_20734,N_19037,N_19112);
xnor U20735 (N_20735,N_19166,N_19763);
and U20736 (N_20736,N_19507,N_19668);
or U20737 (N_20737,N_19785,N_19383);
and U20738 (N_20738,N_19440,N_19664);
xor U20739 (N_20739,N_19110,N_19531);
nand U20740 (N_20740,N_19589,N_19107);
xor U20741 (N_20741,N_19319,N_19887);
or U20742 (N_20742,N_19820,N_19647);
xnor U20743 (N_20743,N_19044,N_19022);
xnor U20744 (N_20744,N_19508,N_19262);
nand U20745 (N_20745,N_19797,N_19393);
nand U20746 (N_20746,N_19025,N_19016);
nand U20747 (N_20747,N_19518,N_19720);
nand U20748 (N_20748,N_19317,N_19181);
and U20749 (N_20749,N_19200,N_19593);
nand U20750 (N_20750,N_19860,N_19832);
nor U20751 (N_20751,N_19495,N_19368);
nor U20752 (N_20752,N_19679,N_19619);
or U20753 (N_20753,N_19530,N_19472);
nor U20754 (N_20754,N_19635,N_19936);
or U20755 (N_20755,N_19192,N_19939);
nor U20756 (N_20756,N_19824,N_19715);
or U20757 (N_20757,N_19675,N_19818);
and U20758 (N_20758,N_19717,N_19877);
nand U20759 (N_20759,N_19471,N_19142);
nor U20760 (N_20760,N_19965,N_19484);
and U20761 (N_20761,N_19796,N_19090);
or U20762 (N_20762,N_19968,N_19726);
or U20763 (N_20763,N_19190,N_19221);
or U20764 (N_20764,N_19194,N_19778);
nor U20765 (N_20765,N_19823,N_19455);
xor U20766 (N_20766,N_19500,N_19536);
and U20767 (N_20767,N_19360,N_19401);
and U20768 (N_20768,N_19885,N_19724);
nor U20769 (N_20769,N_19647,N_19558);
xor U20770 (N_20770,N_19945,N_19636);
or U20771 (N_20771,N_19096,N_19019);
and U20772 (N_20772,N_19611,N_19180);
nand U20773 (N_20773,N_19252,N_19194);
and U20774 (N_20774,N_19222,N_19148);
xnor U20775 (N_20775,N_19150,N_19434);
nor U20776 (N_20776,N_19998,N_19873);
and U20777 (N_20777,N_19087,N_19883);
nor U20778 (N_20778,N_19517,N_19496);
or U20779 (N_20779,N_19478,N_19188);
nand U20780 (N_20780,N_19181,N_19360);
nor U20781 (N_20781,N_19515,N_19616);
nor U20782 (N_20782,N_19655,N_19590);
or U20783 (N_20783,N_19172,N_19804);
nor U20784 (N_20784,N_19092,N_19811);
nand U20785 (N_20785,N_19799,N_19525);
and U20786 (N_20786,N_19226,N_19018);
nand U20787 (N_20787,N_19530,N_19225);
nor U20788 (N_20788,N_19474,N_19944);
or U20789 (N_20789,N_19719,N_19922);
nor U20790 (N_20790,N_19924,N_19330);
nor U20791 (N_20791,N_19972,N_19878);
or U20792 (N_20792,N_19639,N_19099);
nor U20793 (N_20793,N_19995,N_19913);
and U20794 (N_20794,N_19945,N_19926);
and U20795 (N_20795,N_19307,N_19277);
and U20796 (N_20796,N_19795,N_19399);
nor U20797 (N_20797,N_19257,N_19052);
or U20798 (N_20798,N_19055,N_19135);
or U20799 (N_20799,N_19537,N_19995);
nor U20800 (N_20800,N_19476,N_19991);
xor U20801 (N_20801,N_19439,N_19880);
or U20802 (N_20802,N_19369,N_19416);
nand U20803 (N_20803,N_19942,N_19935);
nor U20804 (N_20804,N_19436,N_19028);
xnor U20805 (N_20805,N_19402,N_19641);
nand U20806 (N_20806,N_19562,N_19500);
xor U20807 (N_20807,N_19226,N_19485);
xor U20808 (N_20808,N_19696,N_19038);
nand U20809 (N_20809,N_19366,N_19444);
nor U20810 (N_20810,N_19611,N_19515);
and U20811 (N_20811,N_19521,N_19313);
or U20812 (N_20812,N_19994,N_19447);
xor U20813 (N_20813,N_19023,N_19702);
xnor U20814 (N_20814,N_19286,N_19222);
and U20815 (N_20815,N_19240,N_19772);
and U20816 (N_20816,N_19495,N_19827);
xor U20817 (N_20817,N_19255,N_19258);
xor U20818 (N_20818,N_19762,N_19950);
and U20819 (N_20819,N_19806,N_19070);
and U20820 (N_20820,N_19845,N_19037);
xnor U20821 (N_20821,N_19719,N_19304);
and U20822 (N_20822,N_19478,N_19313);
nand U20823 (N_20823,N_19326,N_19591);
and U20824 (N_20824,N_19595,N_19375);
nor U20825 (N_20825,N_19959,N_19310);
or U20826 (N_20826,N_19258,N_19452);
nand U20827 (N_20827,N_19781,N_19378);
xnor U20828 (N_20828,N_19120,N_19913);
nor U20829 (N_20829,N_19895,N_19744);
nand U20830 (N_20830,N_19816,N_19622);
nor U20831 (N_20831,N_19076,N_19249);
nor U20832 (N_20832,N_19113,N_19377);
and U20833 (N_20833,N_19273,N_19244);
or U20834 (N_20834,N_19428,N_19540);
nor U20835 (N_20835,N_19680,N_19590);
xnor U20836 (N_20836,N_19160,N_19714);
nand U20837 (N_20837,N_19686,N_19182);
xor U20838 (N_20838,N_19476,N_19893);
nor U20839 (N_20839,N_19899,N_19549);
nor U20840 (N_20840,N_19693,N_19214);
nand U20841 (N_20841,N_19738,N_19998);
or U20842 (N_20842,N_19477,N_19158);
or U20843 (N_20843,N_19859,N_19051);
xnor U20844 (N_20844,N_19589,N_19151);
or U20845 (N_20845,N_19220,N_19342);
xor U20846 (N_20846,N_19389,N_19865);
xnor U20847 (N_20847,N_19705,N_19141);
xnor U20848 (N_20848,N_19435,N_19045);
nand U20849 (N_20849,N_19228,N_19276);
nand U20850 (N_20850,N_19614,N_19936);
xnor U20851 (N_20851,N_19357,N_19071);
nor U20852 (N_20852,N_19783,N_19477);
xnor U20853 (N_20853,N_19290,N_19829);
nor U20854 (N_20854,N_19265,N_19992);
and U20855 (N_20855,N_19482,N_19429);
and U20856 (N_20856,N_19507,N_19370);
nand U20857 (N_20857,N_19185,N_19067);
nand U20858 (N_20858,N_19559,N_19379);
xnor U20859 (N_20859,N_19649,N_19246);
and U20860 (N_20860,N_19238,N_19955);
and U20861 (N_20861,N_19321,N_19290);
nor U20862 (N_20862,N_19354,N_19187);
xor U20863 (N_20863,N_19666,N_19936);
nor U20864 (N_20864,N_19566,N_19458);
and U20865 (N_20865,N_19466,N_19233);
or U20866 (N_20866,N_19927,N_19588);
or U20867 (N_20867,N_19854,N_19418);
nand U20868 (N_20868,N_19049,N_19834);
and U20869 (N_20869,N_19677,N_19636);
xnor U20870 (N_20870,N_19982,N_19796);
nand U20871 (N_20871,N_19877,N_19675);
nand U20872 (N_20872,N_19743,N_19603);
nand U20873 (N_20873,N_19507,N_19963);
xnor U20874 (N_20874,N_19161,N_19374);
nand U20875 (N_20875,N_19524,N_19496);
and U20876 (N_20876,N_19083,N_19455);
nand U20877 (N_20877,N_19462,N_19489);
nor U20878 (N_20878,N_19265,N_19311);
xor U20879 (N_20879,N_19874,N_19413);
nor U20880 (N_20880,N_19208,N_19128);
nor U20881 (N_20881,N_19722,N_19557);
and U20882 (N_20882,N_19029,N_19175);
nor U20883 (N_20883,N_19823,N_19380);
or U20884 (N_20884,N_19579,N_19826);
nand U20885 (N_20885,N_19148,N_19321);
xnor U20886 (N_20886,N_19961,N_19716);
nor U20887 (N_20887,N_19907,N_19251);
xor U20888 (N_20888,N_19176,N_19765);
and U20889 (N_20889,N_19671,N_19963);
xor U20890 (N_20890,N_19222,N_19532);
nor U20891 (N_20891,N_19995,N_19700);
nand U20892 (N_20892,N_19064,N_19963);
or U20893 (N_20893,N_19356,N_19392);
or U20894 (N_20894,N_19504,N_19706);
and U20895 (N_20895,N_19473,N_19283);
nand U20896 (N_20896,N_19874,N_19522);
or U20897 (N_20897,N_19840,N_19245);
nand U20898 (N_20898,N_19517,N_19788);
nor U20899 (N_20899,N_19218,N_19393);
and U20900 (N_20900,N_19693,N_19299);
and U20901 (N_20901,N_19207,N_19632);
or U20902 (N_20902,N_19801,N_19235);
nor U20903 (N_20903,N_19999,N_19801);
and U20904 (N_20904,N_19259,N_19452);
nand U20905 (N_20905,N_19878,N_19182);
nand U20906 (N_20906,N_19985,N_19304);
xor U20907 (N_20907,N_19155,N_19339);
and U20908 (N_20908,N_19170,N_19510);
nand U20909 (N_20909,N_19499,N_19493);
xnor U20910 (N_20910,N_19305,N_19515);
nor U20911 (N_20911,N_19885,N_19128);
nor U20912 (N_20912,N_19157,N_19790);
nor U20913 (N_20913,N_19307,N_19227);
and U20914 (N_20914,N_19882,N_19196);
and U20915 (N_20915,N_19958,N_19241);
nand U20916 (N_20916,N_19756,N_19238);
nor U20917 (N_20917,N_19971,N_19226);
or U20918 (N_20918,N_19992,N_19488);
xnor U20919 (N_20919,N_19143,N_19560);
xor U20920 (N_20920,N_19917,N_19183);
nand U20921 (N_20921,N_19405,N_19877);
xor U20922 (N_20922,N_19265,N_19471);
nand U20923 (N_20923,N_19641,N_19878);
or U20924 (N_20924,N_19040,N_19931);
nand U20925 (N_20925,N_19330,N_19963);
nand U20926 (N_20926,N_19545,N_19466);
nor U20927 (N_20927,N_19425,N_19247);
nand U20928 (N_20928,N_19117,N_19515);
and U20929 (N_20929,N_19822,N_19963);
xor U20930 (N_20930,N_19550,N_19726);
xnor U20931 (N_20931,N_19616,N_19392);
xnor U20932 (N_20932,N_19300,N_19169);
or U20933 (N_20933,N_19217,N_19364);
and U20934 (N_20934,N_19142,N_19073);
xor U20935 (N_20935,N_19956,N_19923);
or U20936 (N_20936,N_19669,N_19992);
nor U20937 (N_20937,N_19684,N_19086);
or U20938 (N_20938,N_19900,N_19120);
xnor U20939 (N_20939,N_19425,N_19341);
nor U20940 (N_20940,N_19563,N_19371);
nor U20941 (N_20941,N_19182,N_19720);
or U20942 (N_20942,N_19380,N_19698);
nand U20943 (N_20943,N_19503,N_19335);
nor U20944 (N_20944,N_19772,N_19705);
nor U20945 (N_20945,N_19870,N_19715);
or U20946 (N_20946,N_19905,N_19183);
nand U20947 (N_20947,N_19196,N_19104);
nand U20948 (N_20948,N_19355,N_19047);
xnor U20949 (N_20949,N_19130,N_19965);
nand U20950 (N_20950,N_19187,N_19666);
or U20951 (N_20951,N_19768,N_19639);
nand U20952 (N_20952,N_19774,N_19476);
xor U20953 (N_20953,N_19997,N_19097);
and U20954 (N_20954,N_19888,N_19865);
nand U20955 (N_20955,N_19665,N_19091);
nand U20956 (N_20956,N_19951,N_19256);
nand U20957 (N_20957,N_19772,N_19091);
or U20958 (N_20958,N_19832,N_19044);
nand U20959 (N_20959,N_19332,N_19672);
xor U20960 (N_20960,N_19130,N_19539);
nor U20961 (N_20961,N_19714,N_19705);
xnor U20962 (N_20962,N_19828,N_19528);
nor U20963 (N_20963,N_19803,N_19843);
xnor U20964 (N_20964,N_19415,N_19735);
nand U20965 (N_20965,N_19395,N_19986);
and U20966 (N_20966,N_19050,N_19803);
and U20967 (N_20967,N_19032,N_19690);
xnor U20968 (N_20968,N_19076,N_19292);
and U20969 (N_20969,N_19092,N_19873);
xor U20970 (N_20970,N_19355,N_19614);
and U20971 (N_20971,N_19537,N_19189);
or U20972 (N_20972,N_19610,N_19614);
or U20973 (N_20973,N_19728,N_19511);
nor U20974 (N_20974,N_19115,N_19830);
nor U20975 (N_20975,N_19155,N_19212);
xnor U20976 (N_20976,N_19875,N_19428);
or U20977 (N_20977,N_19203,N_19255);
or U20978 (N_20978,N_19175,N_19667);
xnor U20979 (N_20979,N_19892,N_19976);
and U20980 (N_20980,N_19109,N_19079);
nor U20981 (N_20981,N_19337,N_19487);
and U20982 (N_20982,N_19442,N_19257);
xnor U20983 (N_20983,N_19504,N_19006);
or U20984 (N_20984,N_19337,N_19020);
and U20985 (N_20985,N_19706,N_19229);
nor U20986 (N_20986,N_19852,N_19388);
nand U20987 (N_20987,N_19577,N_19059);
xnor U20988 (N_20988,N_19688,N_19114);
and U20989 (N_20989,N_19805,N_19106);
or U20990 (N_20990,N_19358,N_19679);
nand U20991 (N_20991,N_19657,N_19478);
nand U20992 (N_20992,N_19786,N_19608);
xnor U20993 (N_20993,N_19060,N_19819);
and U20994 (N_20994,N_19589,N_19374);
nand U20995 (N_20995,N_19806,N_19298);
or U20996 (N_20996,N_19225,N_19131);
xnor U20997 (N_20997,N_19474,N_19145);
and U20998 (N_20998,N_19731,N_19675);
and U20999 (N_20999,N_19167,N_19579);
nor U21000 (N_21000,N_20453,N_20510);
nand U21001 (N_21001,N_20605,N_20688);
nor U21002 (N_21002,N_20342,N_20365);
and U21003 (N_21003,N_20777,N_20463);
or U21004 (N_21004,N_20962,N_20149);
nand U21005 (N_21005,N_20237,N_20960);
and U21006 (N_21006,N_20611,N_20207);
xor U21007 (N_21007,N_20056,N_20895);
and U21008 (N_21008,N_20241,N_20886);
nor U21009 (N_21009,N_20200,N_20528);
nor U21010 (N_21010,N_20825,N_20088);
xor U21011 (N_21011,N_20987,N_20862);
or U21012 (N_21012,N_20107,N_20867);
nand U21013 (N_21013,N_20831,N_20262);
or U21014 (N_21014,N_20730,N_20722);
or U21015 (N_21015,N_20236,N_20058);
and U21016 (N_21016,N_20803,N_20440);
nor U21017 (N_21017,N_20340,N_20026);
xnor U21018 (N_21018,N_20087,N_20823);
nand U21019 (N_21019,N_20721,N_20285);
xor U21020 (N_21020,N_20143,N_20238);
xor U21021 (N_21021,N_20907,N_20197);
nand U21022 (N_21022,N_20979,N_20530);
nor U21023 (N_21023,N_20290,N_20656);
nor U21024 (N_21024,N_20851,N_20917);
or U21025 (N_21025,N_20063,N_20927);
xnor U21026 (N_21026,N_20188,N_20269);
and U21027 (N_21027,N_20943,N_20403);
nand U21028 (N_21028,N_20925,N_20921);
xnor U21029 (N_21029,N_20360,N_20167);
and U21030 (N_21030,N_20083,N_20878);
nor U21031 (N_21031,N_20859,N_20002);
nor U21032 (N_21032,N_20334,N_20909);
nand U21033 (N_21033,N_20701,N_20601);
nand U21034 (N_21034,N_20216,N_20915);
xor U21035 (N_21035,N_20336,N_20935);
and U21036 (N_21036,N_20792,N_20355);
nor U21037 (N_21037,N_20848,N_20116);
nand U21038 (N_21038,N_20180,N_20743);
or U21039 (N_21039,N_20281,N_20413);
xor U21040 (N_21040,N_20538,N_20304);
or U21041 (N_21041,N_20379,N_20890);
or U21042 (N_21042,N_20193,N_20748);
and U21043 (N_21043,N_20571,N_20888);
nand U21044 (N_21044,N_20104,N_20028);
nor U21045 (N_21045,N_20489,N_20439);
nor U21046 (N_21046,N_20785,N_20273);
nor U21047 (N_21047,N_20306,N_20723);
nand U21048 (N_21048,N_20132,N_20959);
xnor U21049 (N_21049,N_20141,N_20551);
or U21050 (N_21050,N_20337,N_20583);
nor U21051 (N_21051,N_20364,N_20993);
nor U21052 (N_21052,N_20557,N_20980);
or U21053 (N_21053,N_20402,N_20647);
or U21054 (N_21054,N_20398,N_20870);
and U21055 (N_21055,N_20247,N_20584);
or U21056 (N_21056,N_20173,N_20469);
or U21057 (N_21057,N_20989,N_20901);
and U21058 (N_21058,N_20122,N_20084);
nor U21059 (N_21059,N_20427,N_20120);
and U21060 (N_21060,N_20081,N_20997);
xnor U21061 (N_21061,N_20539,N_20800);
nor U21062 (N_21062,N_20487,N_20418);
or U21063 (N_21063,N_20508,N_20258);
and U21064 (N_21064,N_20010,N_20838);
xnor U21065 (N_21065,N_20559,N_20872);
nor U21066 (N_21066,N_20079,N_20251);
xnor U21067 (N_21067,N_20986,N_20380);
xnor U21068 (N_21068,N_20902,N_20178);
nor U21069 (N_21069,N_20225,N_20674);
and U21070 (N_21070,N_20804,N_20694);
and U21071 (N_21071,N_20593,N_20548);
and U21072 (N_21072,N_20125,N_20531);
or U21073 (N_21073,N_20267,N_20345);
and U21074 (N_21074,N_20108,N_20455);
nand U21075 (N_21075,N_20617,N_20343);
or U21076 (N_21076,N_20335,N_20372);
nand U21077 (N_21077,N_20763,N_20856);
or U21078 (N_21078,N_20199,N_20492);
xnor U21079 (N_21079,N_20071,N_20272);
or U21080 (N_21080,N_20212,N_20136);
nor U21081 (N_21081,N_20388,N_20810);
and U21082 (N_21082,N_20672,N_20154);
and U21083 (N_21083,N_20261,N_20406);
nor U21084 (N_21084,N_20201,N_20051);
or U21085 (N_21085,N_20327,N_20483);
nand U21086 (N_21086,N_20462,N_20952);
or U21087 (N_21087,N_20266,N_20348);
nand U21088 (N_21088,N_20973,N_20930);
nand U21089 (N_21089,N_20985,N_20495);
and U21090 (N_21090,N_20958,N_20347);
xnor U21091 (N_21091,N_20760,N_20466);
or U21092 (N_21092,N_20170,N_20752);
nand U21093 (N_21093,N_20519,N_20160);
or U21094 (N_21094,N_20322,N_20875);
or U21095 (N_21095,N_20908,N_20727);
and U21096 (N_21096,N_20183,N_20203);
nor U21097 (N_21097,N_20246,N_20771);
nand U21098 (N_21098,N_20494,N_20702);
nor U21099 (N_21099,N_20227,N_20544);
or U21100 (N_21100,N_20249,N_20186);
or U21101 (N_21101,N_20817,N_20184);
and U21102 (N_21102,N_20061,N_20728);
and U21103 (N_21103,N_20351,N_20503);
or U21104 (N_21104,N_20357,N_20585);
and U21105 (N_21105,N_20371,N_20014);
nor U21106 (N_21106,N_20929,N_20138);
or U21107 (N_21107,N_20550,N_20198);
nor U21108 (N_21108,N_20067,N_20277);
nor U21109 (N_21109,N_20738,N_20594);
or U21110 (N_21110,N_20021,N_20471);
nand U21111 (N_21111,N_20712,N_20928);
xnor U21112 (N_21112,N_20680,N_20295);
and U21113 (N_21113,N_20181,N_20474);
and U21114 (N_21114,N_20595,N_20911);
xnor U21115 (N_21115,N_20946,N_20782);
or U21116 (N_21116,N_20622,N_20918);
and U21117 (N_21117,N_20298,N_20709);
xnor U21118 (N_21118,N_20103,N_20953);
nor U21119 (N_21119,N_20383,N_20852);
nand U21120 (N_21120,N_20232,N_20592);
and U21121 (N_21121,N_20317,N_20366);
xnor U21122 (N_21122,N_20844,N_20751);
nand U21123 (N_21123,N_20377,N_20369);
nand U21124 (N_21124,N_20243,N_20969);
and U21125 (N_21125,N_20003,N_20770);
nand U21126 (N_21126,N_20038,N_20478);
and U21127 (N_21127,N_20954,N_20824);
or U21128 (N_21128,N_20210,N_20678);
nand U21129 (N_21129,N_20430,N_20786);
nor U21130 (N_21130,N_20265,N_20644);
nor U21131 (N_21131,N_20972,N_20789);
nor U21132 (N_21132,N_20704,N_20846);
nand U21133 (N_21133,N_20699,N_20080);
or U21134 (N_21134,N_20042,N_20527);
and U21135 (N_21135,N_20049,N_20260);
or U21136 (N_21136,N_20553,N_20191);
xor U21137 (N_21137,N_20448,N_20681);
or U21138 (N_21138,N_20773,N_20395);
nor U21139 (N_21139,N_20577,N_20637);
and U21140 (N_21140,N_20431,N_20580);
nor U21141 (N_21141,N_20609,N_20239);
and U21142 (N_21142,N_20164,N_20172);
xor U21143 (N_21143,N_20613,N_20725);
nor U21144 (N_21144,N_20912,N_20816);
and U21145 (N_21145,N_20421,N_20209);
nor U21146 (N_21146,N_20683,N_20603);
xnor U21147 (N_21147,N_20756,N_20323);
nand U21148 (N_21148,N_20697,N_20023);
xor U21149 (N_21149,N_20964,N_20903);
xor U21150 (N_21150,N_20939,N_20898);
and U21151 (N_21151,N_20843,N_20500);
and U21152 (N_21152,N_20022,N_20479);
nand U21153 (N_21153,N_20994,N_20155);
or U21154 (N_21154,N_20151,N_20668);
nor U21155 (N_21155,N_20971,N_20480);
nor U21156 (N_21156,N_20967,N_20196);
or U21157 (N_21157,N_20558,N_20339);
nor U21158 (N_21158,N_20338,N_20161);
nor U21159 (N_21159,N_20050,N_20124);
nor U21160 (N_21160,N_20441,N_20625);
or U21161 (N_21161,N_20133,N_20407);
nor U21162 (N_21162,N_20409,N_20213);
nand U21163 (N_21163,N_20110,N_20546);
or U21164 (N_21164,N_20127,N_20233);
and U21165 (N_21165,N_20025,N_20333);
nand U21166 (N_21166,N_20205,N_20001);
nor U21167 (N_21167,N_20904,N_20828);
or U21168 (N_21168,N_20621,N_20673);
nand U21169 (N_21169,N_20948,N_20600);
and U21170 (N_21170,N_20436,N_20072);
nor U21171 (N_21171,N_20653,N_20192);
or U21172 (N_21172,N_20381,N_20477);
xnor U21173 (N_21173,N_20498,N_20586);
xor U21174 (N_21174,N_20714,N_20642);
nand U21175 (N_21175,N_20849,N_20419);
or U21176 (N_21176,N_20030,N_20982);
xnor U21177 (N_21177,N_20045,N_20762);
or U21178 (N_21178,N_20535,N_20385);
xor U21179 (N_21179,N_20187,N_20597);
and U21180 (N_21180,N_20717,N_20111);
nor U21181 (N_21181,N_20115,N_20534);
nand U21182 (N_21182,N_20879,N_20537);
nor U21183 (N_21183,N_20949,N_20386);
nor U21184 (N_21184,N_20796,N_20596);
nand U21185 (N_21185,N_20975,N_20623);
nor U21186 (N_21186,N_20005,N_20288);
or U21187 (N_21187,N_20486,N_20018);
xor U21188 (N_21188,N_20944,N_20361);
nor U21189 (N_21189,N_20812,N_20437);
nand U21190 (N_21190,N_20344,N_20995);
xor U21191 (N_21191,N_20991,N_20839);
nand U21192 (N_21192,N_20822,N_20420);
and U21193 (N_21193,N_20685,N_20788);
nand U21194 (N_21194,N_20556,N_20957);
nor U21195 (N_21195,N_20208,N_20194);
or U21196 (N_21196,N_20842,N_20502);
and U21197 (N_21197,N_20378,N_20602);
xnor U21198 (N_21198,N_20891,N_20873);
and U21199 (N_21199,N_20860,N_20117);
nor U21200 (N_21200,N_20029,N_20914);
nand U21201 (N_21201,N_20497,N_20341);
and U21202 (N_21202,N_20148,N_20765);
and U21203 (N_21203,N_20449,N_20565);
or U21204 (N_21204,N_20526,N_20607);
nand U21205 (N_21205,N_20865,N_20636);
or U21206 (N_21206,N_20428,N_20065);
nor U21207 (N_21207,N_20068,N_20169);
nor U21208 (N_21208,N_20629,N_20650);
and U21209 (N_21209,N_20139,N_20640);
nor U21210 (N_21210,N_20082,N_20073);
nor U21211 (N_21211,N_20518,N_20687);
xor U21212 (N_21212,N_20819,N_20657);
and U21213 (N_21213,N_20706,N_20326);
and U21214 (N_21214,N_20228,N_20159);
xnor U21215 (N_21215,N_20696,N_20411);
nor U21216 (N_21216,N_20708,N_20575);
nor U21217 (N_21217,N_20443,N_20086);
xor U21218 (N_21218,N_20620,N_20264);
nor U21219 (N_21219,N_20999,N_20204);
nor U21220 (N_21220,N_20561,N_20833);
nand U21221 (N_21221,N_20099,N_20889);
xor U21222 (N_21222,N_20313,N_20598);
nor U21223 (N_21223,N_20147,N_20162);
nand U21224 (N_21224,N_20452,N_20686);
nor U21225 (N_21225,N_20118,N_20638);
xnor U21226 (N_21226,N_20434,N_20009);
and U21227 (N_21227,N_20863,N_20280);
xor U21228 (N_21228,N_20887,N_20809);
nand U21229 (N_21229,N_20924,N_20077);
and U21230 (N_21230,N_20276,N_20066);
nor U21231 (N_21231,N_20900,N_20716);
xor U21232 (N_21232,N_20224,N_20695);
and U21233 (N_21233,N_20855,N_20362);
and U21234 (N_21234,N_20412,N_20813);
xor U21235 (N_21235,N_20129,N_20284);
xor U21236 (N_21236,N_20984,N_20504);
nor U21237 (N_21237,N_20632,N_20263);
nor U21238 (N_21238,N_20608,N_20031);
and U21239 (N_21239,N_20299,N_20736);
and U21240 (N_21240,N_20746,N_20660);
and U21241 (N_21241,N_20564,N_20222);
and U21242 (N_21242,N_20710,N_20775);
xnor U21243 (N_21243,N_20798,N_20916);
nand U21244 (N_21244,N_20591,N_20737);
or U21245 (N_21245,N_20433,N_20218);
nor U21246 (N_21246,N_20257,N_20303);
xor U21247 (N_21247,N_20974,N_20445);
or U21248 (N_21248,N_20389,N_20324);
nand U21249 (N_21249,N_20845,N_20932);
nand U21250 (N_21250,N_20017,N_20589);
nor U21251 (N_21251,N_20325,N_20020);
xnor U21252 (N_21252,N_20000,N_20783);
or U21253 (N_21253,N_20998,N_20074);
or U21254 (N_21254,N_20007,N_20349);
or U21255 (N_21255,N_20158,N_20793);
and U21256 (N_21256,N_20945,N_20542);
nor U21257 (N_21257,N_20415,N_20215);
or U21258 (N_21258,N_20835,N_20392);
xor U21259 (N_21259,N_20882,N_20075);
nor U21260 (N_21260,N_20245,N_20599);
and U21261 (N_21261,N_20226,N_20572);
nand U21262 (N_21262,N_20757,N_20829);
xnor U21263 (N_21263,N_20297,N_20085);
xnor U21264 (N_21264,N_20032,N_20741);
xor U21265 (N_21265,N_20936,N_20432);
nand U21266 (N_21266,N_20676,N_20460);
xnor U21267 (N_21267,N_20871,N_20536);
xnor U21268 (N_21268,N_20664,N_20938);
or U21269 (N_21269,N_20836,N_20950);
xor U21270 (N_21270,N_20098,N_20689);
and U21271 (N_21271,N_20052,N_20970);
or U21272 (N_21272,N_20758,N_20753);
nor U21273 (N_21273,N_20626,N_20093);
xor U21274 (N_21274,N_20543,N_20511);
or U21275 (N_21275,N_20787,N_20404);
and U21276 (N_21276,N_20978,N_20874);
nor U21277 (N_21277,N_20624,N_20552);
and U21278 (N_21278,N_20861,N_20229);
nor U21279 (N_21279,N_20923,N_20648);
nor U21280 (N_21280,N_20137,N_20457);
xnor U21281 (N_21281,N_20293,N_20521);
and U21282 (N_21282,N_20509,N_20353);
nor U21283 (N_21283,N_20618,N_20157);
nor U21284 (N_21284,N_20214,N_20316);
nand U21285 (N_21285,N_20422,N_20896);
nand U21286 (N_21286,N_20897,N_20016);
nor U21287 (N_21287,N_20641,N_20726);
nor U21288 (N_21288,N_20646,N_20152);
or U21289 (N_21289,N_20275,N_20482);
and U21290 (N_21290,N_20514,N_20513);
and U21291 (N_21291,N_20314,N_20966);
xor U21292 (N_21292,N_20145,N_20034);
nor U21293 (N_21293,N_20576,N_20036);
nor U21294 (N_21294,N_20095,N_20130);
or U21295 (N_21295,N_20554,N_20300);
nand U21296 (N_21296,N_20818,N_20253);
and U21297 (N_21297,N_20866,N_20069);
xnor U21298 (N_21298,N_20296,N_20240);
nand U21299 (N_21299,N_20567,N_20105);
nor U21300 (N_21300,N_20382,N_20794);
nor U21301 (N_21301,N_20910,N_20675);
and U21302 (N_21302,N_20220,N_20101);
xnor U21303 (N_21303,N_20135,N_20078);
nor U21304 (N_21304,N_20713,N_20040);
and U21305 (N_21305,N_20501,N_20894);
or U21306 (N_21306,N_20619,N_20573);
or U21307 (N_21307,N_20146,N_20308);
nor U21308 (N_21308,N_20857,N_20955);
or U21309 (N_21309,N_20144,N_20057);
nand U21310 (N_21310,N_20268,N_20354);
nand U21311 (N_21311,N_20291,N_20035);
and U21312 (N_21312,N_20830,N_20332);
nor U21313 (N_21313,N_20456,N_20174);
and U21314 (N_21314,N_20096,N_20307);
or U21315 (N_21315,N_20490,N_20292);
nand U21316 (N_21316,N_20705,N_20754);
or U21317 (N_21317,N_20278,N_20808);
xor U21318 (N_21318,N_20634,N_20677);
or U21319 (N_21319,N_20691,N_20750);
or U21320 (N_21320,N_20540,N_20176);
or U21321 (N_21321,N_20506,N_20426);
xor U21322 (N_21322,N_20358,N_20799);
or U21323 (N_21323,N_20318,N_20662);
and U21324 (N_21324,N_20013,N_20892);
and U21325 (N_21325,N_20610,N_20252);
or U21326 (N_21326,N_20522,N_20881);
nand U21327 (N_21327,N_20834,N_20363);
nand U21328 (N_21328,N_20126,N_20346);
or U21329 (N_21329,N_20821,N_20475);
xor U21330 (N_21330,N_20692,N_20217);
or U21331 (N_21331,N_20202,N_20092);
or U21332 (N_21332,N_20190,N_20850);
xor U21333 (N_21333,N_20759,N_20123);
xor U21334 (N_21334,N_20114,N_20163);
nand U21335 (N_21335,N_20920,N_20715);
xnor U21336 (N_21336,N_20195,N_20992);
nor U21337 (N_21337,N_20242,N_20905);
nor U21338 (N_21338,N_20488,N_20711);
or U21339 (N_21339,N_20840,N_20230);
or U21340 (N_21340,N_20179,N_20811);
xor U21341 (N_21341,N_20397,N_20739);
nand U21342 (N_21342,N_20767,N_20033);
and U21343 (N_21343,N_20569,N_20484);
nand U21344 (N_21344,N_20832,N_20700);
or U21345 (N_21345,N_20880,N_20669);
or U21346 (N_21346,N_20545,N_20121);
and U21347 (N_21347,N_20352,N_20628);
nand U21348 (N_21348,N_20951,N_20019);
nand U21349 (N_21349,N_20631,N_20493);
nand U21350 (N_21350,N_20934,N_20464);
and U21351 (N_21351,N_20532,N_20271);
xor U21352 (N_21352,N_20054,N_20359);
or U21353 (N_21353,N_20279,N_20919);
or U21354 (N_21354,N_20405,N_20931);
nor U21355 (N_21355,N_20259,N_20731);
nor U21356 (N_21356,N_20070,N_20523);
xor U21357 (N_21357,N_20106,N_20447);
xor U21358 (N_21358,N_20250,N_20734);
nand U21359 (N_21359,N_20761,N_20368);
or U21360 (N_21360,N_20424,N_20320);
and U21361 (N_21361,N_20076,N_20206);
xnor U21362 (N_21362,N_20899,N_20091);
xor U21363 (N_21363,N_20826,N_20956);
nor U21364 (N_21364,N_20394,N_20315);
or U21365 (N_21365,N_20373,N_20254);
nand U21366 (N_21366,N_20667,N_20517);
nor U21367 (N_21367,N_20302,N_20578);
nor U21368 (N_21368,N_20961,N_20166);
xor U21369 (N_21369,N_20582,N_20707);
nor U21370 (N_21370,N_20563,N_20541);
or U21371 (N_21371,N_20735,N_20330);
nor U21372 (N_21372,N_20053,N_20131);
xnor U21373 (N_21373,N_20779,N_20516);
or U21374 (N_21374,N_20549,N_20283);
nand U21375 (N_21375,N_20574,N_20732);
or U21376 (N_21376,N_20312,N_20684);
nor U21377 (N_21377,N_20733,N_20451);
nor U21378 (N_21378,N_20854,N_20047);
nor U21379 (N_21379,N_20755,N_20864);
and U21380 (N_21380,N_20645,N_20442);
nor U21381 (N_21381,N_20524,N_20940);
or U21382 (N_21382,N_20491,N_20046);
and U21383 (N_21383,N_20024,N_20976);
nand U21384 (N_21384,N_20496,N_20791);
nor U21385 (N_21385,N_20234,N_20877);
or U21386 (N_21386,N_20112,N_20375);
xnor U21387 (N_21387,N_20612,N_20893);
or U21388 (N_21388,N_20627,N_20505);
or U21389 (N_21389,N_20814,N_20795);
nand U21390 (N_21390,N_20113,N_20807);
and U21391 (N_21391,N_20665,N_20168);
nor U21392 (N_21392,N_20512,N_20635);
nand U21393 (N_21393,N_20282,N_20408);
xor U21394 (N_21394,N_20011,N_20438);
xor U21395 (N_21395,N_20778,N_20768);
xor U21396 (N_21396,N_20467,N_20868);
nor U21397 (N_21397,N_20719,N_20965);
nor U21398 (N_21398,N_20094,N_20328);
or U21399 (N_21399,N_20776,N_20802);
or U21400 (N_21400,N_20764,N_20703);
xnor U21401 (N_21401,N_20801,N_20044);
nand U21402 (N_21402,N_20309,N_20461);
nor U21403 (N_21403,N_20926,N_20185);
or U21404 (N_21404,N_20659,N_20745);
and U21405 (N_21405,N_20097,N_20682);
xor U21406 (N_21406,N_20922,N_20481);
and U21407 (N_21407,N_20064,N_20287);
nor U21408 (N_21408,N_20289,N_20235);
xor U21409 (N_21409,N_20219,N_20876);
or U21410 (N_21410,N_20128,N_20742);
xnor U21411 (N_21411,N_20156,N_20633);
or U21412 (N_21412,N_20853,N_20189);
nor U21413 (N_21413,N_20401,N_20244);
or U21414 (N_21414,N_20400,N_20331);
nor U21415 (N_21415,N_20465,N_20520);
nand U21416 (N_21416,N_20906,N_20454);
and U21417 (N_21417,N_20350,N_20039);
nor U21418 (N_21418,N_20140,N_20529);
nor U21419 (N_21419,N_20294,N_20525);
and U21420 (N_21420,N_20869,N_20004);
xor U21421 (N_21421,N_20305,N_20396);
nand U21422 (N_21422,N_20274,N_20153);
and U21423 (N_21423,N_20150,N_20827);
xnor U21424 (N_21424,N_20231,N_20740);
or U21425 (N_21425,N_20416,N_20485);
and U21426 (N_21426,N_20615,N_20671);
nand U21427 (N_21427,N_20604,N_20473);
and U21428 (N_21428,N_20841,N_20724);
nand U21429 (N_21429,N_20560,N_20109);
and U21430 (N_21430,N_20270,N_20175);
nand U21431 (N_21431,N_20988,N_20643);
xor U21432 (N_21432,N_20568,N_20815);
and U21433 (N_21433,N_20367,N_20037);
nor U21434 (N_21434,N_20165,N_20774);
or U21435 (N_21435,N_20060,N_20384);
xnor U21436 (N_21436,N_20444,N_20679);
and U21437 (N_21437,N_20171,N_20102);
and U21438 (N_21438,N_20820,N_20566);
nand U21439 (N_21439,N_20781,N_20654);
nor U21440 (N_21440,N_20606,N_20790);
xor U21441 (N_21441,N_20211,N_20256);
and U21442 (N_21442,N_20425,N_20470);
nor U21443 (N_21443,N_20720,N_20616);
and U21444 (N_21444,N_20649,N_20947);
xnor U21445 (N_21445,N_20006,N_20806);
and U21446 (N_21446,N_20570,N_20374);
nand U21447 (N_21447,N_20885,N_20744);
nor U21448 (N_21448,N_20329,N_20614);
xnor U21449 (N_21449,N_20499,N_20446);
or U21450 (N_21450,N_20387,N_20937);
nor U21451 (N_21451,N_20090,N_20766);
xor U21452 (N_21452,N_20507,N_20652);
and U21453 (N_21453,N_20391,N_20968);
nand U21454 (N_21454,N_20579,N_20015);
or U21455 (N_21455,N_20658,N_20772);
xnor U21456 (N_21456,N_20301,N_20942);
nor U21457 (N_21457,N_20913,N_20749);
nand U21458 (N_21458,N_20459,N_20769);
xor U21459 (N_21459,N_20562,N_20729);
nor U21460 (N_21460,N_20693,N_20515);
nand U21461 (N_21461,N_20670,N_20780);
nand U21462 (N_21462,N_20399,N_20472);
xor U21463 (N_21463,N_20718,N_20784);
xnor U21464 (N_21464,N_20255,N_20883);
nor U21465 (N_21465,N_20698,N_20248);
nor U21466 (N_21466,N_20376,N_20533);
nand U21467 (N_21467,N_20356,N_20414);
xnor U21468 (N_21468,N_20321,N_20996);
xor U21469 (N_21469,N_20119,N_20048);
or U21470 (N_21470,N_20012,N_20555);
xor U21471 (N_21471,N_20310,N_20933);
or U21472 (N_21472,N_20100,N_20429);
xor U21473 (N_21473,N_20588,N_20221);
and U21474 (N_21474,N_20142,N_20027);
xnor U21475 (N_21475,N_20458,N_20590);
nand U21476 (N_21476,N_20663,N_20884);
nor U21477 (N_21477,N_20547,N_20805);
nand U21478 (N_21478,N_20059,N_20690);
nand U21479 (N_21479,N_20651,N_20223);
or U21480 (N_21480,N_20587,N_20630);
nand U21481 (N_21481,N_20476,N_20941);
xor U21482 (N_21482,N_20043,N_20311);
and U21483 (N_21483,N_20981,N_20008);
nand U21484 (N_21484,N_20666,N_20858);
and U21485 (N_21485,N_20435,N_20055);
xor U21486 (N_21486,N_20977,N_20286);
nand U21487 (N_21487,N_20062,N_20655);
nand U21488 (N_21488,N_20041,N_20417);
nand U21489 (N_21489,N_20393,N_20423);
or U21490 (N_21490,N_20639,N_20990);
and U21491 (N_21491,N_20661,N_20370);
xnor U21492 (N_21492,N_20319,N_20983);
nand U21493 (N_21493,N_20963,N_20450);
or U21494 (N_21494,N_20134,N_20837);
xor U21495 (N_21495,N_20468,N_20747);
nand U21496 (N_21496,N_20089,N_20847);
xnor U21497 (N_21497,N_20182,N_20797);
and U21498 (N_21498,N_20177,N_20581);
or U21499 (N_21499,N_20390,N_20410);
xnor U21500 (N_21500,N_20594,N_20716);
xor U21501 (N_21501,N_20434,N_20721);
or U21502 (N_21502,N_20328,N_20574);
nand U21503 (N_21503,N_20781,N_20491);
nand U21504 (N_21504,N_20760,N_20126);
nor U21505 (N_21505,N_20342,N_20473);
xor U21506 (N_21506,N_20057,N_20805);
nand U21507 (N_21507,N_20141,N_20588);
and U21508 (N_21508,N_20482,N_20417);
nand U21509 (N_21509,N_20090,N_20488);
and U21510 (N_21510,N_20987,N_20870);
nand U21511 (N_21511,N_20938,N_20775);
and U21512 (N_21512,N_20424,N_20654);
nand U21513 (N_21513,N_20781,N_20075);
and U21514 (N_21514,N_20938,N_20462);
xor U21515 (N_21515,N_20754,N_20055);
nand U21516 (N_21516,N_20780,N_20323);
xor U21517 (N_21517,N_20517,N_20330);
nor U21518 (N_21518,N_20673,N_20576);
and U21519 (N_21519,N_20140,N_20334);
nand U21520 (N_21520,N_20523,N_20313);
nor U21521 (N_21521,N_20284,N_20983);
xor U21522 (N_21522,N_20418,N_20333);
nand U21523 (N_21523,N_20193,N_20258);
nor U21524 (N_21524,N_20386,N_20933);
xnor U21525 (N_21525,N_20697,N_20610);
nand U21526 (N_21526,N_20020,N_20049);
and U21527 (N_21527,N_20687,N_20112);
and U21528 (N_21528,N_20035,N_20799);
nand U21529 (N_21529,N_20275,N_20819);
nand U21530 (N_21530,N_20257,N_20351);
nor U21531 (N_21531,N_20169,N_20041);
nand U21532 (N_21532,N_20455,N_20049);
nand U21533 (N_21533,N_20472,N_20332);
or U21534 (N_21534,N_20944,N_20206);
and U21535 (N_21535,N_20431,N_20890);
and U21536 (N_21536,N_20046,N_20247);
and U21537 (N_21537,N_20726,N_20801);
nand U21538 (N_21538,N_20080,N_20563);
or U21539 (N_21539,N_20075,N_20660);
xnor U21540 (N_21540,N_20193,N_20787);
nor U21541 (N_21541,N_20420,N_20830);
xor U21542 (N_21542,N_20688,N_20324);
nand U21543 (N_21543,N_20745,N_20183);
nor U21544 (N_21544,N_20340,N_20760);
xnor U21545 (N_21545,N_20753,N_20124);
nor U21546 (N_21546,N_20736,N_20098);
and U21547 (N_21547,N_20435,N_20873);
or U21548 (N_21548,N_20520,N_20519);
nand U21549 (N_21549,N_20231,N_20279);
nand U21550 (N_21550,N_20120,N_20392);
xnor U21551 (N_21551,N_20446,N_20438);
xnor U21552 (N_21552,N_20979,N_20570);
and U21553 (N_21553,N_20999,N_20636);
nor U21554 (N_21554,N_20049,N_20299);
xor U21555 (N_21555,N_20746,N_20341);
and U21556 (N_21556,N_20889,N_20282);
xnor U21557 (N_21557,N_20921,N_20569);
and U21558 (N_21558,N_20201,N_20449);
and U21559 (N_21559,N_20785,N_20015);
nor U21560 (N_21560,N_20114,N_20229);
or U21561 (N_21561,N_20005,N_20874);
xnor U21562 (N_21562,N_20232,N_20942);
or U21563 (N_21563,N_20615,N_20272);
nor U21564 (N_21564,N_20522,N_20757);
and U21565 (N_21565,N_20479,N_20487);
xor U21566 (N_21566,N_20486,N_20911);
nand U21567 (N_21567,N_20244,N_20989);
and U21568 (N_21568,N_20354,N_20139);
and U21569 (N_21569,N_20888,N_20214);
xor U21570 (N_21570,N_20035,N_20944);
nand U21571 (N_21571,N_20149,N_20533);
and U21572 (N_21572,N_20805,N_20570);
and U21573 (N_21573,N_20948,N_20771);
nor U21574 (N_21574,N_20508,N_20875);
xor U21575 (N_21575,N_20342,N_20347);
nor U21576 (N_21576,N_20846,N_20384);
nand U21577 (N_21577,N_20728,N_20682);
or U21578 (N_21578,N_20195,N_20793);
and U21579 (N_21579,N_20956,N_20540);
nand U21580 (N_21580,N_20793,N_20322);
or U21581 (N_21581,N_20136,N_20897);
and U21582 (N_21582,N_20487,N_20941);
and U21583 (N_21583,N_20661,N_20493);
nand U21584 (N_21584,N_20180,N_20309);
or U21585 (N_21585,N_20305,N_20862);
xnor U21586 (N_21586,N_20956,N_20147);
nor U21587 (N_21587,N_20988,N_20279);
nand U21588 (N_21588,N_20424,N_20312);
or U21589 (N_21589,N_20149,N_20794);
xnor U21590 (N_21590,N_20786,N_20344);
nor U21591 (N_21591,N_20751,N_20946);
nand U21592 (N_21592,N_20764,N_20358);
and U21593 (N_21593,N_20956,N_20264);
nand U21594 (N_21594,N_20790,N_20344);
nand U21595 (N_21595,N_20084,N_20263);
nand U21596 (N_21596,N_20038,N_20225);
or U21597 (N_21597,N_20948,N_20912);
or U21598 (N_21598,N_20494,N_20423);
or U21599 (N_21599,N_20129,N_20844);
nor U21600 (N_21600,N_20450,N_20697);
xor U21601 (N_21601,N_20637,N_20398);
nor U21602 (N_21602,N_20078,N_20819);
nand U21603 (N_21603,N_20062,N_20729);
xnor U21604 (N_21604,N_20983,N_20046);
nand U21605 (N_21605,N_20871,N_20532);
nand U21606 (N_21606,N_20835,N_20939);
nand U21607 (N_21607,N_20964,N_20009);
or U21608 (N_21608,N_20373,N_20867);
or U21609 (N_21609,N_20316,N_20217);
nand U21610 (N_21610,N_20005,N_20891);
or U21611 (N_21611,N_20415,N_20095);
nor U21612 (N_21612,N_20516,N_20664);
nor U21613 (N_21613,N_20803,N_20433);
nand U21614 (N_21614,N_20602,N_20406);
nand U21615 (N_21615,N_20524,N_20679);
or U21616 (N_21616,N_20225,N_20289);
and U21617 (N_21617,N_20656,N_20172);
xor U21618 (N_21618,N_20124,N_20364);
and U21619 (N_21619,N_20540,N_20091);
and U21620 (N_21620,N_20432,N_20110);
nor U21621 (N_21621,N_20279,N_20879);
xor U21622 (N_21622,N_20943,N_20818);
nor U21623 (N_21623,N_20239,N_20229);
or U21624 (N_21624,N_20182,N_20477);
xor U21625 (N_21625,N_20652,N_20578);
nor U21626 (N_21626,N_20672,N_20958);
and U21627 (N_21627,N_20768,N_20947);
xor U21628 (N_21628,N_20356,N_20008);
xnor U21629 (N_21629,N_20921,N_20291);
nand U21630 (N_21630,N_20412,N_20199);
or U21631 (N_21631,N_20579,N_20693);
nand U21632 (N_21632,N_20533,N_20164);
or U21633 (N_21633,N_20691,N_20974);
or U21634 (N_21634,N_20459,N_20766);
nor U21635 (N_21635,N_20281,N_20795);
xnor U21636 (N_21636,N_20571,N_20119);
xnor U21637 (N_21637,N_20491,N_20493);
xnor U21638 (N_21638,N_20369,N_20485);
xor U21639 (N_21639,N_20610,N_20506);
xnor U21640 (N_21640,N_20065,N_20701);
nand U21641 (N_21641,N_20341,N_20802);
and U21642 (N_21642,N_20868,N_20044);
and U21643 (N_21643,N_20633,N_20382);
xor U21644 (N_21644,N_20250,N_20202);
or U21645 (N_21645,N_20606,N_20099);
or U21646 (N_21646,N_20053,N_20849);
nor U21647 (N_21647,N_20845,N_20905);
nor U21648 (N_21648,N_20119,N_20634);
nand U21649 (N_21649,N_20478,N_20766);
nand U21650 (N_21650,N_20578,N_20293);
or U21651 (N_21651,N_20353,N_20421);
and U21652 (N_21652,N_20716,N_20783);
nand U21653 (N_21653,N_20834,N_20278);
or U21654 (N_21654,N_20258,N_20721);
nand U21655 (N_21655,N_20656,N_20210);
nand U21656 (N_21656,N_20458,N_20735);
nand U21657 (N_21657,N_20659,N_20915);
nor U21658 (N_21658,N_20487,N_20131);
and U21659 (N_21659,N_20957,N_20565);
xor U21660 (N_21660,N_20489,N_20197);
or U21661 (N_21661,N_20044,N_20724);
or U21662 (N_21662,N_20856,N_20441);
nand U21663 (N_21663,N_20163,N_20918);
xnor U21664 (N_21664,N_20954,N_20769);
nor U21665 (N_21665,N_20142,N_20855);
nand U21666 (N_21666,N_20306,N_20752);
xnor U21667 (N_21667,N_20255,N_20906);
nor U21668 (N_21668,N_20006,N_20294);
xnor U21669 (N_21669,N_20965,N_20731);
nor U21670 (N_21670,N_20134,N_20344);
or U21671 (N_21671,N_20307,N_20475);
nand U21672 (N_21672,N_20069,N_20114);
or U21673 (N_21673,N_20178,N_20187);
and U21674 (N_21674,N_20798,N_20723);
and U21675 (N_21675,N_20409,N_20240);
nand U21676 (N_21676,N_20173,N_20495);
xor U21677 (N_21677,N_20104,N_20194);
and U21678 (N_21678,N_20509,N_20779);
xor U21679 (N_21679,N_20532,N_20897);
and U21680 (N_21680,N_20110,N_20658);
xnor U21681 (N_21681,N_20387,N_20720);
and U21682 (N_21682,N_20028,N_20461);
or U21683 (N_21683,N_20289,N_20540);
nand U21684 (N_21684,N_20279,N_20146);
nand U21685 (N_21685,N_20640,N_20036);
and U21686 (N_21686,N_20927,N_20596);
nor U21687 (N_21687,N_20501,N_20918);
nor U21688 (N_21688,N_20332,N_20319);
and U21689 (N_21689,N_20153,N_20185);
nor U21690 (N_21690,N_20117,N_20595);
nor U21691 (N_21691,N_20804,N_20961);
nor U21692 (N_21692,N_20261,N_20756);
xor U21693 (N_21693,N_20999,N_20759);
xnor U21694 (N_21694,N_20669,N_20997);
nor U21695 (N_21695,N_20803,N_20655);
nand U21696 (N_21696,N_20719,N_20403);
and U21697 (N_21697,N_20728,N_20828);
nand U21698 (N_21698,N_20686,N_20068);
or U21699 (N_21699,N_20508,N_20611);
nand U21700 (N_21700,N_20180,N_20252);
xor U21701 (N_21701,N_20141,N_20802);
nor U21702 (N_21702,N_20243,N_20321);
or U21703 (N_21703,N_20756,N_20203);
and U21704 (N_21704,N_20494,N_20947);
and U21705 (N_21705,N_20579,N_20517);
xnor U21706 (N_21706,N_20122,N_20990);
or U21707 (N_21707,N_20653,N_20186);
xor U21708 (N_21708,N_20629,N_20512);
nor U21709 (N_21709,N_20385,N_20025);
and U21710 (N_21710,N_20987,N_20590);
xor U21711 (N_21711,N_20135,N_20029);
nor U21712 (N_21712,N_20216,N_20549);
or U21713 (N_21713,N_20573,N_20052);
or U21714 (N_21714,N_20601,N_20835);
nor U21715 (N_21715,N_20143,N_20670);
nor U21716 (N_21716,N_20717,N_20515);
xor U21717 (N_21717,N_20992,N_20666);
and U21718 (N_21718,N_20110,N_20217);
or U21719 (N_21719,N_20409,N_20505);
or U21720 (N_21720,N_20570,N_20660);
or U21721 (N_21721,N_20556,N_20904);
nor U21722 (N_21722,N_20270,N_20639);
xnor U21723 (N_21723,N_20395,N_20994);
or U21724 (N_21724,N_20671,N_20606);
nand U21725 (N_21725,N_20804,N_20077);
and U21726 (N_21726,N_20781,N_20215);
nor U21727 (N_21727,N_20693,N_20586);
and U21728 (N_21728,N_20878,N_20451);
xor U21729 (N_21729,N_20997,N_20373);
and U21730 (N_21730,N_20066,N_20126);
xnor U21731 (N_21731,N_20487,N_20402);
or U21732 (N_21732,N_20989,N_20157);
xnor U21733 (N_21733,N_20595,N_20300);
xor U21734 (N_21734,N_20099,N_20128);
nor U21735 (N_21735,N_20736,N_20071);
or U21736 (N_21736,N_20459,N_20087);
and U21737 (N_21737,N_20180,N_20963);
and U21738 (N_21738,N_20267,N_20840);
and U21739 (N_21739,N_20389,N_20591);
nor U21740 (N_21740,N_20658,N_20646);
xnor U21741 (N_21741,N_20119,N_20829);
nand U21742 (N_21742,N_20641,N_20671);
and U21743 (N_21743,N_20239,N_20773);
nand U21744 (N_21744,N_20362,N_20327);
and U21745 (N_21745,N_20322,N_20578);
and U21746 (N_21746,N_20949,N_20533);
and U21747 (N_21747,N_20046,N_20456);
nor U21748 (N_21748,N_20707,N_20540);
and U21749 (N_21749,N_20771,N_20720);
xnor U21750 (N_21750,N_20006,N_20756);
and U21751 (N_21751,N_20703,N_20215);
and U21752 (N_21752,N_20205,N_20433);
nand U21753 (N_21753,N_20807,N_20451);
or U21754 (N_21754,N_20370,N_20771);
or U21755 (N_21755,N_20946,N_20076);
nor U21756 (N_21756,N_20682,N_20566);
and U21757 (N_21757,N_20781,N_20823);
xor U21758 (N_21758,N_20291,N_20828);
nand U21759 (N_21759,N_20983,N_20498);
nand U21760 (N_21760,N_20355,N_20556);
or U21761 (N_21761,N_20395,N_20105);
nand U21762 (N_21762,N_20452,N_20705);
nor U21763 (N_21763,N_20795,N_20214);
nand U21764 (N_21764,N_20196,N_20401);
xor U21765 (N_21765,N_20421,N_20489);
nor U21766 (N_21766,N_20176,N_20661);
nor U21767 (N_21767,N_20570,N_20693);
xor U21768 (N_21768,N_20859,N_20011);
nor U21769 (N_21769,N_20472,N_20620);
xor U21770 (N_21770,N_20539,N_20100);
nor U21771 (N_21771,N_20538,N_20741);
xnor U21772 (N_21772,N_20745,N_20919);
and U21773 (N_21773,N_20028,N_20298);
nand U21774 (N_21774,N_20903,N_20010);
xor U21775 (N_21775,N_20117,N_20453);
nor U21776 (N_21776,N_20037,N_20226);
nor U21777 (N_21777,N_20890,N_20738);
or U21778 (N_21778,N_20453,N_20885);
xnor U21779 (N_21779,N_20555,N_20048);
nand U21780 (N_21780,N_20548,N_20256);
nor U21781 (N_21781,N_20262,N_20658);
xor U21782 (N_21782,N_20736,N_20638);
xnor U21783 (N_21783,N_20510,N_20780);
or U21784 (N_21784,N_20376,N_20456);
or U21785 (N_21785,N_20529,N_20254);
nand U21786 (N_21786,N_20790,N_20091);
nand U21787 (N_21787,N_20611,N_20655);
nand U21788 (N_21788,N_20610,N_20278);
or U21789 (N_21789,N_20551,N_20342);
nor U21790 (N_21790,N_20796,N_20967);
or U21791 (N_21791,N_20534,N_20886);
nand U21792 (N_21792,N_20536,N_20403);
xor U21793 (N_21793,N_20711,N_20678);
and U21794 (N_21794,N_20461,N_20296);
xnor U21795 (N_21795,N_20203,N_20857);
nand U21796 (N_21796,N_20924,N_20892);
nor U21797 (N_21797,N_20434,N_20501);
and U21798 (N_21798,N_20945,N_20191);
and U21799 (N_21799,N_20515,N_20449);
and U21800 (N_21800,N_20450,N_20310);
or U21801 (N_21801,N_20814,N_20587);
xnor U21802 (N_21802,N_20237,N_20949);
nor U21803 (N_21803,N_20867,N_20802);
and U21804 (N_21804,N_20318,N_20042);
or U21805 (N_21805,N_20768,N_20203);
xor U21806 (N_21806,N_20040,N_20117);
or U21807 (N_21807,N_20593,N_20560);
xor U21808 (N_21808,N_20431,N_20167);
nor U21809 (N_21809,N_20319,N_20549);
nor U21810 (N_21810,N_20121,N_20447);
and U21811 (N_21811,N_20853,N_20431);
nand U21812 (N_21812,N_20300,N_20889);
nor U21813 (N_21813,N_20356,N_20211);
and U21814 (N_21814,N_20133,N_20317);
nor U21815 (N_21815,N_20412,N_20236);
and U21816 (N_21816,N_20571,N_20296);
nor U21817 (N_21817,N_20272,N_20972);
or U21818 (N_21818,N_20649,N_20146);
nor U21819 (N_21819,N_20234,N_20311);
or U21820 (N_21820,N_20269,N_20466);
and U21821 (N_21821,N_20276,N_20526);
nor U21822 (N_21822,N_20416,N_20672);
nor U21823 (N_21823,N_20966,N_20528);
nand U21824 (N_21824,N_20512,N_20356);
and U21825 (N_21825,N_20823,N_20204);
xnor U21826 (N_21826,N_20396,N_20505);
nor U21827 (N_21827,N_20304,N_20239);
and U21828 (N_21828,N_20366,N_20025);
xnor U21829 (N_21829,N_20293,N_20755);
nor U21830 (N_21830,N_20810,N_20974);
xnor U21831 (N_21831,N_20563,N_20626);
nor U21832 (N_21832,N_20708,N_20894);
nor U21833 (N_21833,N_20441,N_20619);
xor U21834 (N_21834,N_20572,N_20222);
or U21835 (N_21835,N_20016,N_20039);
and U21836 (N_21836,N_20347,N_20454);
or U21837 (N_21837,N_20953,N_20303);
and U21838 (N_21838,N_20466,N_20817);
nor U21839 (N_21839,N_20424,N_20601);
nor U21840 (N_21840,N_20421,N_20601);
nand U21841 (N_21841,N_20953,N_20570);
nand U21842 (N_21842,N_20343,N_20790);
nor U21843 (N_21843,N_20583,N_20454);
xnor U21844 (N_21844,N_20245,N_20327);
nor U21845 (N_21845,N_20139,N_20811);
and U21846 (N_21846,N_20223,N_20395);
and U21847 (N_21847,N_20319,N_20740);
and U21848 (N_21848,N_20537,N_20855);
nand U21849 (N_21849,N_20860,N_20603);
nand U21850 (N_21850,N_20487,N_20730);
nor U21851 (N_21851,N_20822,N_20727);
or U21852 (N_21852,N_20912,N_20969);
nor U21853 (N_21853,N_20715,N_20631);
nand U21854 (N_21854,N_20156,N_20421);
and U21855 (N_21855,N_20877,N_20792);
and U21856 (N_21856,N_20027,N_20669);
and U21857 (N_21857,N_20177,N_20579);
and U21858 (N_21858,N_20046,N_20344);
xnor U21859 (N_21859,N_20095,N_20048);
xor U21860 (N_21860,N_20690,N_20383);
xor U21861 (N_21861,N_20397,N_20348);
and U21862 (N_21862,N_20360,N_20635);
xnor U21863 (N_21863,N_20168,N_20610);
nand U21864 (N_21864,N_20626,N_20694);
nand U21865 (N_21865,N_20129,N_20695);
nor U21866 (N_21866,N_20254,N_20956);
nand U21867 (N_21867,N_20919,N_20288);
or U21868 (N_21868,N_20450,N_20480);
nor U21869 (N_21869,N_20017,N_20009);
nor U21870 (N_21870,N_20808,N_20154);
and U21871 (N_21871,N_20217,N_20350);
nand U21872 (N_21872,N_20858,N_20793);
and U21873 (N_21873,N_20980,N_20405);
and U21874 (N_21874,N_20992,N_20127);
or U21875 (N_21875,N_20349,N_20724);
xor U21876 (N_21876,N_20070,N_20919);
and U21877 (N_21877,N_20904,N_20985);
nand U21878 (N_21878,N_20319,N_20352);
xor U21879 (N_21879,N_20228,N_20975);
and U21880 (N_21880,N_20588,N_20456);
and U21881 (N_21881,N_20945,N_20405);
nor U21882 (N_21882,N_20720,N_20607);
nor U21883 (N_21883,N_20803,N_20760);
and U21884 (N_21884,N_20851,N_20743);
and U21885 (N_21885,N_20822,N_20142);
nand U21886 (N_21886,N_20668,N_20238);
and U21887 (N_21887,N_20097,N_20915);
nand U21888 (N_21888,N_20623,N_20547);
nor U21889 (N_21889,N_20912,N_20607);
or U21890 (N_21890,N_20688,N_20834);
nor U21891 (N_21891,N_20327,N_20281);
nor U21892 (N_21892,N_20365,N_20352);
and U21893 (N_21893,N_20882,N_20062);
xor U21894 (N_21894,N_20859,N_20247);
nor U21895 (N_21895,N_20761,N_20096);
and U21896 (N_21896,N_20514,N_20212);
or U21897 (N_21897,N_20864,N_20407);
nor U21898 (N_21898,N_20988,N_20167);
and U21899 (N_21899,N_20999,N_20718);
or U21900 (N_21900,N_20577,N_20826);
nor U21901 (N_21901,N_20161,N_20157);
nand U21902 (N_21902,N_20556,N_20256);
nand U21903 (N_21903,N_20573,N_20448);
or U21904 (N_21904,N_20108,N_20465);
nor U21905 (N_21905,N_20288,N_20531);
and U21906 (N_21906,N_20756,N_20990);
and U21907 (N_21907,N_20943,N_20723);
nand U21908 (N_21908,N_20296,N_20964);
or U21909 (N_21909,N_20173,N_20185);
nor U21910 (N_21910,N_20895,N_20050);
xnor U21911 (N_21911,N_20870,N_20073);
and U21912 (N_21912,N_20522,N_20977);
nand U21913 (N_21913,N_20528,N_20319);
nand U21914 (N_21914,N_20582,N_20811);
or U21915 (N_21915,N_20292,N_20534);
xor U21916 (N_21916,N_20634,N_20833);
or U21917 (N_21917,N_20851,N_20002);
xor U21918 (N_21918,N_20229,N_20465);
xor U21919 (N_21919,N_20005,N_20125);
and U21920 (N_21920,N_20413,N_20663);
or U21921 (N_21921,N_20453,N_20700);
xor U21922 (N_21922,N_20089,N_20291);
nor U21923 (N_21923,N_20478,N_20578);
and U21924 (N_21924,N_20811,N_20322);
xnor U21925 (N_21925,N_20776,N_20033);
nor U21926 (N_21926,N_20621,N_20097);
or U21927 (N_21927,N_20855,N_20230);
nand U21928 (N_21928,N_20893,N_20744);
or U21929 (N_21929,N_20717,N_20179);
nor U21930 (N_21930,N_20941,N_20417);
nor U21931 (N_21931,N_20420,N_20551);
nor U21932 (N_21932,N_20416,N_20458);
or U21933 (N_21933,N_20340,N_20920);
nand U21934 (N_21934,N_20666,N_20527);
nor U21935 (N_21935,N_20441,N_20394);
nand U21936 (N_21936,N_20034,N_20007);
nand U21937 (N_21937,N_20202,N_20435);
nor U21938 (N_21938,N_20321,N_20435);
or U21939 (N_21939,N_20206,N_20272);
xor U21940 (N_21940,N_20480,N_20257);
xnor U21941 (N_21941,N_20379,N_20941);
xor U21942 (N_21942,N_20365,N_20067);
or U21943 (N_21943,N_20846,N_20433);
nor U21944 (N_21944,N_20173,N_20102);
nor U21945 (N_21945,N_20289,N_20402);
nor U21946 (N_21946,N_20503,N_20907);
and U21947 (N_21947,N_20817,N_20585);
nor U21948 (N_21948,N_20273,N_20354);
nor U21949 (N_21949,N_20344,N_20719);
nand U21950 (N_21950,N_20096,N_20403);
and U21951 (N_21951,N_20345,N_20172);
nand U21952 (N_21952,N_20080,N_20732);
or U21953 (N_21953,N_20577,N_20904);
xnor U21954 (N_21954,N_20320,N_20352);
and U21955 (N_21955,N_20825,N_20261);
or U21956 (N_21956,N_20024,N_20912);
or U21957 (N_21957,N_20743,N_20938);
or U21958 (N_21958,N_20836,N_20763);
xor U21959 (N_21959,N_20611,N_20496);
or U21960 (N_21960,N_20452,N_20054);
or U21961 (N_21961,N_20494,N_20729);
nor U21962 (N_21962,N_20536,N_20313);
xor U21963 (N_21963,N_20106,N_20658);
nor U21964 (N_21964,N_20374,N_20679);
and U21965 (N_21965,N_20789,N_20287);
and U21966 (N_21966,N_20111,N_20603);
and U21967 (N_21967,N_20546,N_20409);
or U21968 (N_21968,N_20448,N_20873);
nand U21969 (N_21969,N_20794,N_20564);
and U21970 (N_21970,N_20404,N_20711);
nor U21971 (N_21971,N_20475,N_20139);
or U21972 (N_21972,N_20725,N_20383);
nand U21973 (N_21973,N_20112,N_20862);
nor U21974 (N_21974,N_20578,N_20936);
xnor U21975 (N_21975,N_20598,N_20249);
xnor U21976 (N_21976,N_20496,N_20561);
or U21977 (N_21977,N_20421,N_20847);
or U21978 (N_21978,N_20419,N_20338);
nand U21979 (N_21979,N_20417,N_20048);
or U21980 (N_21980,N_20769,N_20260);
nand U21981 (N_21981,N_20960,N_20834);
xnor U21982 (N_21982,N_20019,N_20358);
nand U21983 (N_21983,N_20723,N_20318);
nand U21984 (N_21984,N_20021,N_20081);
or U21985 (N_21985,N_20605,N_20986);
nor U21986 (N_21986,N_20570,N_20802);
xnor U21987 (N_21987,N_20204,N_20100);
nor U21988 (N_21988,N_20579,N_20246);
xnor U21989 (N_21989,N_20485,N_20346);
and U21990 (N_21990,N_20717,N_20849);
nand U21991 (N_21991,N_20009,N_20561);
nand U21992 (N_21992,N_20885,N_20149);
and U21993 (N_21993,N_20953,N_20007);
nand U21994 (N_21994,N_20131,N_20268);
and U21995 (N_21995,N_20346,N_20540);
nand U21996 (N_21996,N_20759,N_20937);
nor U21997 (N_21997,N_20456,N_20758);
nor U21998 (N_21998,N_20380,N_20780);
nor U21999 (N_21999,N_20534,N_20477);
nor U22000 (N_22000,N_21519,N_21827);
xnor U22001 (N_22001,N_21132,N_21478);
or U22002 (N_22002,N_21240,N_21420);
or U22003 (N_22003,N_21379,N_21003);
and U22004 (N_22004,N_21826,N_21388);
nor U22005 (N_22005,N_21100,N_21216);
nand U22006 (N_22006,N_21207,N_21764);
or U22007 (N_22007,N_21244,N_21626);
xor U22008 (N_22008,N_21792,N_21503);
xnor U22009 (N_22009,N_21635,N_21424);
and U22010 (N_22010,N_21303,N_21265);
nor U22011 (N_22011,N_21884,N_21599);
nor U22012 (N_22012,N_21177,N_21540);
or U22013 (N_22013,N_21958,N_21256);
or U22014 (N_22014,N_21849,N_21895);
nand U22015 (N_22015,N_21086,N_21889);
and U22016 (N_22016,N_21128,N_21171);
and U22017 (N_22017,N_21660,N_21162);
nand U22018 (N_22018,N_21771,N_21515);
nand U22019 (N_22019,N_21910,N_21701);
and U22020 (N_22020,N_21316,N_21641);
and U22021 (N_22021,N_21880,N_21102);
nor U22022 (N_22022,N_21000,N_21600);
nor U22023 (N_22023,N_21984,N_21899);
or U22024 (N_22024,N_21746,N_21042);
nor U22025 (N_22025,N_21470,N_21422);
nand U22026 (N_22026,N_21124,N_21770);
nor U22027 (N_22027,N_21924,N_21345);
nand U22028 (N_22028,N_21304,N_21935);
nand U22029 (N_22029,N_21752,N_21725);
nor U22030 (N_22030,N_21759,N_21509);
or U22031 (N_22031,N_21134,N_21987);
and U22032 (N_22032,N_21625,N_21065);
and U22033 (N_22033,N_21313,N_21718);
and U22034 (N_22034,N_21264,N_21914);
and U22035 (N_22035,N_21765,N_21290);
nand U22036 (N_22036,N_21549,N_21988);
and U22037 (N_22037,N_21367,N_21385);
or U22038 (N_22038,N_21961,N_21663);
and U22039 (N_22039,N_21824,N_21412);
nand U22040 (N_22040,N_21782,N_21566);
or U22041 (N_22041,N_21804,N_21917);
nand U22042 (N_22042,N_21278,N_21706);
nor U22043 (N_22043,N_21037,N_21029);
and U22044 (N_22044,N_21273,N_21002);
nand U22045 (N_22045,N_21896,N_21722);
and U22046 (N_22046,N_21212,N_21596);
or U22047 (N_22047,N_21109,N_21327);
nor U22048 (N_22048,N_21035,N_21435);
xor U22049 (N_22049,N_21983,N_21793);
and U22050 (N_22050,N_21032,N_21461);
and U22051 (N_22051,N_21862,N_21514);
or U22052 (N_22052,N_21500,N_21659);
and U22053 (N_22053,N_21059,N_21350);
or U22054 (N_22054,N_21950,N_21730);
xor U22055 (N_22055,N_21133,N_21913);
nor U22056 (N_22056,N_21919,N_21607);
or U22057 (N_22057,N_21881,N_21400);
xnor U22058 (N_22058,N_21015,N_21450);
xor U22059 (N_22059,N_21370,N_21932);
nor U22060 (N_22060,N_21221,N_21834);
xor U22061 (N_22061,N_21794,N_21837);
xor U22062 (N_22062,N_21806,N_21994);
or U22063 (N_22063,N_21639,N_21518);
nand U22064 (N_22064,N_21473,N_21358);
nand U22065 (N_22065,N_21254,N_21172);
nand U22066 (N_22066,N_21406,N_21044);
xor U22067 (N_22067,N_21326,N_21148);
nand U22068 (N_22068,N_21920,N_21971);
nor U22069 (N_22069,N_21159,N_21903);
xnor U22070 (N_22070,N_21665,N_21760);
nor U22071 (N_22071,N_21481,N_21650);
or U22072 (N_22072,N_21947,N_21944);
and U22073 (N_22073,N_21018,N_21452);
or U22074 (N_22074,N_21047,N_21449);
nand U22075 (N_22075,N_21399,N_21209);
xnor U22076 (N_22076,N_21191,N_21643);
xor U22077 (N_22077,N_21407,N_21351);
nand U22078 (N_22078,N_21799,N_21397);
or U22079 (N_22079,N_21292,N_21439);
and U22080 (N_22080,N_21743,N_21858);
or U22081 (N_22081,N_21977,N_21820);
or U22082 (N_22082,N_21550,N_21624);
xnor U22083 (N_22083,N_21538,N_21081);
xor U22084 (N_22084,N_21866,N_21393);
nor U22085 (N_22085,N_21085,N_21025);
or U22086 (N_22086,N_21161,N_21027);
and U22087 (N_22087,N_21705,N_21306);
and U22088 (N_22088,N_21269,N_21170);
or U22089 (N_22089,N_21845,N_21411);
xnor U22090 (N_22090,N_21619,N_21425);
or U22091 (N_22091,N_21401,N_21548);
or U22092 (N_22092,N_21176,N_21480);
or U22093 (N_22093,N_21646,N_21680);
and U22094 (N_22094,N_21854,N_21976);
or U22095 (N_22095,N_21231,N_21729);
nor U22096 (N_22096,N_21459,N_21689);
and U22097 (N_22097,N_21048,N_21555);
nand U22098 (N_22098,N_21954,N_21078);
nor U22099 (N_22099,N_21955,N_21590);
and U22100 (N_22100,N_21959,N_21603);
xor U22101 (N_22101,N_21617,N_21783);
and U22102 (N_22102,N_21011,N_21569);
nand U22103 (N_22103,N_21797,N_21576);
and U22104 (N_22104,N_21922,N_21627);
or U22105 (N_22105,N_21267,N_21588);
nand U22106 (N_22106,N_21777,N_21986);
nand U22107 (N_22107,N_21749,N_21953);
or U22108 (N_22108,N_21876,N_21146);
nor U22109 (N_22109,N_21507,N_21384);
xnor U22110 (N_22110,N_21853,N_21529);
or U22111 (N_22111,N_21214,N_21688);
or U22112 (N_22112,N_21758,N_21785);
nand U22113 (N_22113,N_21638,N_21113);
nor U22114 (N_22114,N_21735,N_21761);
or U22115 (N_22115,N_21152,N_21423);
or U22116 (N_22116,N_21030,N_21522);
xnor U22117 (N_22117,N_21318,N_21182);
xnor U22118 (N_22118,N_21387,N_21070);
nand U22119 (N_22119,N_21186,N_21447);
xor U22120 (N_22120,N_21242,N_21852);
nor U22121 (N_22121,N_21578,N_21380);
or U22122 (N_22122,N_21587,N_21929);
or U22123 (N_22123,N_21960,N_21392);
nand U22124 (N_22124,N_21674,N_21941);
nor U22125 (N_22125,N_21754,N_21690);
nand U22126 (N_22126,N_21312,N_21652);
nand U22127 (N_22127,N_21655,N_21045);
nand U22128 (N_22128,N_21163,N_21181);
nor U22129 (N_22129,N_21293,N_21488);
and U22130 (N_22130,N_21831,N_21877);
xor U22131 (N_22131,N_21322,N_21609);
xnor U22132 (N_22132,N_21651,N_21252);
or U22133 (N_22133,N_21230,N_21506);
and U22134 (N_22134,N_21714,N_21592);
or U22135 (N_22135,N_21942,N_21539);
nand U22136 (N_22136,N_21331,N_21199);
and U22137 (N_22137,N_21137,N_21696);
xor U22138 (N_22138,N_21838,N_21426);
xor U22139 (N_22139,N_21250,N_21004);
nand U22140 (N_22140,N_21263,N_21697);
xor U22141 (N_22141,N_21757,N_21742);
nand U22142 (N_22142,N_21456,N_21012);
xnor U22143 (N_22143,N_21427,N_21939);
nand U22144 (N_22144,N_21679,N_21280);
nor U22145 (N_22145,N_21021,N_21106);
xnor U22146 (N_22146,N_21046,N_21973);
nor U22147 (N_22147,N_21830,N_21258);
and U22148 (N_22148,N_21937,N_21251);
nor U22149 (N_22149,N_21574,N_21239);
nand U22150 (N_22150,N_21325,N_21378);
or U22151 (N_22151,N_21860,N_21693);
and U22152 (N_22152,N_21995,N_21369);
xor U22153 (N_22153,N_21658,N_21395);
and U22154 (N_22154,N_21287,N_21512);
or U22155 (N_22155,N_21098,N_21972);
or U22156 (N_22156,N_21872,N_21339);
xnor U22157 (N_22157,N_21888,N_21766);
nor U22158 (N_22158,N_21798,N_21049);
or U22159 (N_22159,N_21062,N_21173);
nor U22160 (N_22160,N_21008,N_21043);
xnor U22161 (N_22161,N_21362,N_21090);
nor U22162 (N_22162,N_21923,N_21778);
nand U22163 (N_22163,N_21074,N_21390);
nand U22164 (N_22164,N_21433,N_21598);
xor U22165 (N_22165,N_21623,N_21464);
and U22166 (N_22166,N_21408,N_21748);
or U22167 (N_22167,N_21904,N_21238);
nor U22168 (N_22168,N_21482,N_21383);
nor U22169 (N_22169,N_21839,N_21918);
xor U22170 (N_22170,N_21476,N_21466);
nand U22171 (N_22171,N_21374,N_21200);
nand U22172 (N_22172,N_21057,N_21443);
or U22173 (N_22173,N_21165,N_21964);
or U22174 (N_22174,N_21286,N_21898);
or U22175 (N_22175,N_21386,N_21381);
nor U22176 (N_22176,N_21906,N_21121);
or U22177 (N_22177,N_21968,N_21436);
or U22178 (N_22178,N_21192,N_21786);
and U22179 (N_22179,N_21213,N_21299);
or U22180 (N_22180,N_21907,N_21520);
nor U22181 (N_22181,N_21755,N_21962);
nand U22182 (N_22182,N_21204,N_21281);
nor U22183 (N_22183,N_21802,N_21572);
nand U22184 (N_22184,N_21135,N_21727);
xnor U22185 (N_22185,N_21205,N_21353);
or U22186 (N_22186,N_21394,N_21870);
or U22187 (N_22187,N_21026,N_21324);
and U22188 (N_22188,N_21809,N_21801);
or U22189 (N_22189,N_21259,N_21279);
and U22190 (N_22190,N_21933,N_21563);
or U22191 (N_22191,N_21483,N_21175);
or U22192 (N_22192,N_21185,N_21850);
or U22193 (N_22193,N_21726,N_21371);
or U22194 (N_22194,N_21410,N_21716);
nand U22195 (N_22195,N_21763,N_21229);
xnor U22196 (N_22196,N_21431,N_21458);
xnor U22197 (N_22197,N_21808,N_21266);
nor U22198 (N_22198,N_21900,N_21608);
or U22199 (N_22199,N_21979,N_21684);
nand U22200 (N_22200,N_21807,N_21811);
and U22201 (N_22201,N_21111,N_21274);
or U22202 (N_22202,N_21141,N_21298);
and U22203 (N_22203,N_21277,N_21195);
or U22204 (N_22204,N_21149,N_21096);
or U22205 (N_22205,N_21521,N_21320);
nand U22206 (N_22206,N_21467,N_21661);
nand U22207 (N_22207,N_21855,N_21982);
xor U22208 (N_22208,N_21558,N_21672);
nor U22209 (N_22209,N_21041,N_21157);
nand U22210 (N_22210,N_21261,N_21704);
and U22211 (N_22211,N_21375,N_21382);
xor U22212 (N_22212,N_21740,N_21583);
nor U22213 (N_22213,N_21084,N_21594);
nor U22214 (N_22214,N_21938,N_21570);
or U22215 (N_22215,N_21208,N_21836);
nor U22216 (N_22216,N_21075,N_21123);
and U22217 (N_22217,N_21528,N_21787);
nand U22218 (N_22218,N_21315,N_21957);
nor U22219 (N_22219,N_21249,N_21352);
or U22220 (N_22220,N_21695,N_21071);
and U22221 (N_22221,N_21502,N_21333);
nor U22222 (N_22222,N_21063,N_21247);
nand U22223 (N_22223,N_21257,N_21673);
and U22224 (N_22224,N_21878,N_21343);
xor U22225 (N_22225,N_21974,N_21007);
and U22226 (N_22226,N_21130,N_21601);
nand U22227 (N_22227,N_21532,N_21140);
xor U22228 (N_22228,N_21275,N_21622);
nor U22229 (N_22229,N_21871,N_21989);
or U22230 (N_22230,N_21215,N_21843);
nor U22231 (N_22231,N_21024,N_21874);
and U22232 (N_22232,N_21334,N_21329);
nor U22233 (N_22233,N_21441,N_21131);
or U22234 (N_22234,N_21902,N_21819);
or U22235 (N_22235,N_21699,N_21485);
nor U22236 (N_22236,N_21498,N_21656);
nor U22237 (N_22237,N_21104,N_21776);
or U22238 (N_22238,N_21093,N_21775);
and U22239 (N_22239,N_21198,N_21784);
xnor U22240 (N_22240,N_21276,N_21429);
nor U22241 (N_22241,N_21475,N_21762);
nand U22242 (N_22242,N_21413,N_21612);
nor U22243 (N_22243,N_21817,N_21144);
nand U22244 (N_22244,N_21940,N_21501);
nand U22245 (N_22245,N_21565,N_21001);
xor U22246 (N_22246,N_21455,N_21492);
and U22247 (N_22247,N_21815,N_21164);
nor U22248 (N_22248,N_21428,N_21508);
nand U22249 (N_22249,N_21120,N_21129);
nand U22250 (N_22250,N_21092,N_21151);
nand U22251 (N_22251,N_21856,N_21361);
nand U22252 (N_22252,N_21737,N_21389);
or U22253 (N_22253,N_21731,N_21308);
nand U22254 (N_22254,N_21289,N_21348);
nor U22255 (N_22255,N_21056,N_21789);
or U22256 (N_22256,N_21790,N_21582);
xor U22257 (N_22257,N_21417,N_21530);
or U22258 (N_22258,N_21632,N_21158);
nor U22259 (N_22259,N_21892,N_21154);
nand U22260 (N_22260,N_21223,N_21014);
or U22261 (N_22261,N_21219,N_21430);
xnor U22262 (N_22262,N_21403,N_21669);
nand U22263 (N_22263,N_21377,N_21891);
xor U22264 (N_22264,N_21376,N_21497);
or U22265 (N_22265,N_21190,N_21270);
nor U22266 (N_22266,N_21196,N_21125);
nor U22267 (N_22267,N_21863,N_21657);
and U22268 (N_22268,N_21241,N_21709);
and U22269 (N_22269,N_21493,N_21145);
nand U22270 (N_22270,N_21338,N_21768);
nor U22271 (N_22271,N_21559,N_21310);
nand U22272 (N_22272,N_21756,N_21188);
nand U22273 (N_22273,N_21829,N_21613);
nor U22274 (N_22274,N_21936,N_21710);
nand U22275 (N_22275,N_21580,N_21050);
or U22276 (N_22276,N_21544,N_21774);
and U22277 (N_22277,N_21931,N_21945);
and U22278 (N_22278,N_21728,N_21879);
or U22279 (N_22279,N_21543,N_21653);
or U22280 (N_22280,N_21180,N_21547);
xor U22281 (N_22281,N_21479,N_21557);
and U22282 (N_22282,N_21631,N_21398);
nor U22283 (N_22283,N_21531,N_21160);
xnor U22284 (N_22284,N_21992,N_21720);
nor U22285 (N_22285,N_21825,N_21581);
xor U22286 (N_22286,N_21734,N_21554);
and U22287 (N_22287,N_21453,N_21489);
and U22288 (N_22288,N_21998,N_21930);
xnor U22289 (N_22289,N_21117,N_21142);
or U22290 (N_22290,N_21685,N_21496);
nand U22291 (N_22291,N_21115,N_21848);
nand U22292 (N_22292,N_21462,N_21970);
nor U22293 (N_22293,N_21694,N_21823);
or U22294 (N_22294,N_21647,N_21840);
nand U22295 (N_22295,N_21842,N_21859);
or U22296 (N_22296,N_21013,N_21194);
and U22297 (N_22297,N_21857,N_21681);
and U22298 (N_22298,N_21245,N_21184);
xor U22299 (N_22299,N_21354,N_21717);
nand U22300 (N_22300,N_21337,N_21365);
nand U22301 (N_22301,N_21255,N_21670);
nor U22302 (N_22302,N_21687,N_21359);
or U22303 (N_22303,N_21206,N_21321);
nor U22304 (N_22304,N_21751,N_21965);
or U22305 (N_22305,N_21667,N_21224);
nor U22306 (N_22306,N_21724,N_21634);
or U22307 (N_22307,N_21676,N_21039);
xor U22308 (N_22308,N_21103,N_21978);
and U22309 (N_22309,N_21946,N_21943);
xor U22310 (N_22310,N_21602,N_21060);
nand U22311 (N_22311,N_21553,N_21099);
and U22312 (N_22312,N_21341,N_21416);
or U22313 (N_22313,N_21069,N_21054);
xor U22314 (N_22314,N_21993,N_21434);
xor U22315 (N_22315,N_21648,N_21795);
nor U22316 (N_22316,N_21282,N_21966);
or U22317 (N_22317,N_21490,N_21418);
and U22318 (N_22318,N_21332,N_21064);
nand U22319 (N_22319,N_21606,N_21805);
nand U22320 (N_22320,N_21536,N_21391);
xor U22321 (N_22321,N_21168,N_21915);
nand U22322 (N_22322,N_21664,N_21314);
nor U22323 (N_22323,N_21869,N_21368);
xor U22324 (N_22324,N_21868,N_21546);
nor U22325 (N_22325,N_21445,N_21189);
nor U22326 (N_22326,N_21366,N_21969);
xnor U22327 (N_22327,N_21114,N_21921);
and U22328 (N_22328,N_21138,N_21052);
nand U22329 (N_22329,N_21349,N_21451);
xnor U22330 (N_22330,N_21828,N_21197);
and U22331 (N_22331,N_21861,N_21222);
nor U22332 (N_22332,N_21234,N_21169);
and U22333 (N_22333,N_21463,N_21016);
nand U22334 (N_22334,N_21405,N_21061);
and U22335 (N_22335,N_21963,N_21510);
nor U22336 (N_22336,N_21833,N_21225);
xor U22337 (N_22337,N_21295,N_21091);
xnor U22338 (N_22338,N_21262,N_21882);
nand U22339 (N_22339,N_21614,N_21268);
and U22340 (N_22340,N_21284,N_21080);
and U22341 (N_22341,N_21844,N_21203);
xnor U22342 (N_22342,N_21330,N_21564);
nand U22343 (N_22343,N_21094,N_21535);
or U22344 (N_22344,N_21772,N_21072);
or U22345 (N_22345,N_21107,N_21178);
nor U22346 (N_22346,N_21745,N_21662);
or U22347 (N_22347,N_21822,N_21577);
nand U22348 (N_22348,N_21723,N_21595);
nor U22349 (N_22349,N_21927,N_21058);
and U22350 (N_22350,N_21077,N_21193);
or U22351 (N_22351,N_21523,N_21779);
nor U22352 (N_22352,N_21297,N_21788);
nor U22353 (N_22353,N_21702,N_21446);
and U22354 (N_22354,N_21645,N_21202);
nand U22355 (N_22355,N_21873,N_21122);
xnor U22356 (N_22356,N_21611,N_21814);
or U22357 (N_22357,N_21272,N_21901);
nand U22358 (N_22358,N_21736,N_21469);
and U22359 (N_22359,N_21305,N_21031);
xnor U22360 (N_22360,N_21494,N_21119);
or U22361 (N_22361,N_21851,N_21307);
xnor U22362 (N_22362,N_21832,N_21813);
nand U22363 (N_22363,N_21294,N_21791);
nand U22364 (N_22364,N_21703,N_21585);
nand U22365 (N_22365,N_21541,N_21780);
xnor U22366 (N_22366,N_21616,N_21415);
xor U22367 (N_22367,N_21487,N_21511);
xor U22368 (N_22368,N_21108,N_21073);
and U22369 (N_22369,N_21513,N_21356);
nand U22370 (N_22370,N_21033,N_21715);
nor U22371 (N_22371,N_21527,N_21505);
nand U22372 (N_22372,N_21095,N_21841);
xnor U22373 (N_22373,N_21087,N_21409);
xnor U22374 (N_22374,N_21471,N_21311);
xor U22375 (N_22375,N_21719,N_21419);
nand U22376 (N_22376,N_21952,N_21217);
or U22377 (N_22377,N_21781,N_21951);
nor U22378 (N_22378,N_21542,N_21796);
nor U22379 (N_22379,N_21584,N_21909);
nor U22380 (N_22380,N_21928,N_21867);
nand U22381 (N_22381,N_21079,N_21067);
nor U22382 (N_22382,N_21732,N_21890);
nand U22383 (N_22383,N_21621,N_21285);
or U22384 (N_22384,N_21038,N_21153);
nand U22385 (N_22385,N_21579,N_21089);
nor U22386 (N_22386,N_21711,N_21753);
nand U22387 (N_22387,N_21568,N_21296);
or U22388 (N_22388,N_21112,N_21147);
xor U22389 (N_22389,N_21537,N_21773);
or U22390 (N_22390,N_21847,N_21586);
nand U22391 (N_22391,N_21948,N_21975);
xnor U22392 (N_22392,N_21040,N_21097);
nor U22393 (N_22393,N_21812,N_21444);
nor U22394 (N_22394,N_21991,N_21166);
and U22395 (N_22395,N_21739,N_21253);
or U22396 (N_22396,N_21534,N_21051);
nand U22397 (N_22397,N_21105,N_21472);
or U22398 (N_22398,N_21150,N_21967);
or U22399 (N_22399,N_21474,N_21905);
and U22400 (N_22400,N_21560,N_21816);
or U22401 (N_22401,N_21818,N_21414);
or U22402 (N_22402,N_21990,N_21355);
xor U22403 (N_22403,N_21335,N_21821);
or U22404 (N_22404,N_21517,N_21545);
xnor U22405 (N_22405,N_21226,N_21053);
and U22406 (N_22406,N_21432,N_21396);
or U22407 (N_22407,N_21649,N_21344);
xor U22408 (N_22408,N_21009,N_21897);
and U22409 (N_22409,N_21484,N_21934);
or U22410 (N_22410,N_21404,N_21894);
and U22411 (N_22411,N_21036,N_21949);
xnor U22412 (N_22412,N_21211,N_21605);
and U22413 (N_22413,N_21629,N_21402);
and U22414 (N_22414,N_21981,N_21525);
nor U22415 (N_22415,N_21465,N_21068);
nand U22416 (N_22416,N_21319,N_21733);
nand U22417 (N_22417,N_21916,N_21271);
nor U22418 (N_22418,N_21317,N_21491);
nand U22419 (N_22419,N_21227,N_21328);
and U22420 (N_22420,N_21803,N_21533);
xnor U22421 (N_22421,N_21232,N_21682);
nand U22422 (N_22422,N_21283,N_21835);
nand U22423 (N_22423,N_21179,N_21101);
and U22424 (N_22424,N_21228,N_21291);
xnor U22425 (N_22425,N_21747,N_21174);
or U22426 (N_22426,N_21340,N_21865);
xnor U22427 (N_22427,N_21637,N_21926);
and U22428 (N_22428,N_21028,N_21017);
nor U22429 (N_22429,N_21516,N_21288);
and U22430 (N_22430,N_21567,N_21364);
or U22431 (N_22431,N_21301,N_21005);
or U22432 (N_22432,N_21686,N_21700);
or U22433 (N_22433,N_21237,N_21454);
nor U22434 (N_22434,N_21886,N_21210);
xor U22435 (N_22435,N_21925,N_21155);
xnor U22436 (N_22436,N_21526,N_21911);
and U22437 (N_22437,N_21139,N_21524);
nor U22438 (N_22438,N_21336,N_21477);
or U22439 (N_22439,N_21235,N_21342);
nor U22440 (N_22440,N_21551,N_21721);
or U22441 (N_22441,N_21996,N_21691);
or U22442 (N_22442,N_21438,N_21437);
nor U22443 (N_22443,N_21744,N_21022);
or U22444 (N_22444,N_21908,N_21300);
nand U22445 (N_22445,N_21110,N_21167);
nand U22446 (N_22446,N_21246,N_21636);
and U22447 (N_22447,N_21127,N_21372);
and U22448 (N_22448,N_21864,N_21604);
and U22449 (N_22449,N_21708,N_21034);
xor U22450 (N_22450,N_21810,N_21875);
nand U22451 (N_22451,N_21713,N_21668);
nand U22452 (N_22452,N_21457,N_21248);
or U22453 (N_22453,N_21573,N_21556);
nand U22454 (N_22454,N_21769,N_21985);
nor U22455 (N_22455,N_21019,N_21442);
or U22456 (N_22456,N_21373,N_21260);
nor U22457 (N_22457,N_21118,N_21143);
nor U22458 (N_22458,N_21997,N_21885);
xor U22459 (N_22459,N_21309,N_21126);
or U22460 (N_22460,N_21683,N_21712);
and U22461 (N_22461,N_21593,N_21883);
and U22462 (N_22462,N_21630,N_21677);
or U22463 (N_22463,N_21020,N_21912);
and U22464 (N_22464,N_21023,N_21610);
xor U22465 (N_22465,N_21654,N_21666);
and U22466 (N_22466,N_21187,N_21571);
or U22467 (N_22467,N_21243,N_21887);
nor U22468 (N_22468,N_21642,N_21136);
nand U22469 (N_22469,N_21066,N_21671);
nor U22470 (N_22470,N_21495,N_21504);
nor U22471 (N_22471,N_21448,N_21156);
xor U22472 (N_22472,N_21692,N_21201);
nand U22473 (N_22473,N_21347,N_21360);
and U22474 (N_22474,N_21707,N_21346);
and U22475 (N_22475,N_21591,N_21236);
nor U22476 (N_22476,N_21323,N_21800);
xor U22477 (N_22477,N_21698,N_21421);
nor U22478 (N_22478,N_21575,N_21083);
nor U22479 (N_22479,N_21220,N_21010);
and U22480 (N_22480,N_21741,N_21218);
nor U22481 (N_22481,N_21440,N_21738);
nor U22482 (N_22482,N_21006,N_21076);
xor U22483 (N_22483,N_21846,N_21460);
xor U22484 (N_22484,N_21082,N_21363);
or U22485 (N_22485,N_21116,N_21302);
nand U22486 (N_22486,N_21552,N_21633);
or U22487 (N_22487,N_21767,N_21562);
or U22488 (N_22488,N_21357,N_21675);
nor U22489 (N_22489,N_21620,N_21183);
xnor U22490 (N_22490,N_21618,N_21956);
and U22491 (N_22491,N_21640,N_21678);
xor U22492 (N_22492,N_21999,N_21597);
nand U22493 (N_22493,N_21468,N_21499);
nand U22494 (N_22494,N_21088,N_21644);
nand U22495 (N_22495,N_21561,N_21893);
and U22496 (N_22496,N_21980,N_21055);
and U22497 (N_22497,N_21615,N_21628);
or U22498 (N_22498,N_21589,N_21750);
nand U22499 (N_22499,N_21486,N_21233);
nand U22500 (N_22500,N_21878,N_21681);
or U22501 (N_22501,N_21437,N_21826);
nand U22502 (N_22502,N_21239,N_21063);
xnor U22503 (N_22503,N_21832,N_21952);
xor U22504 (N_22504,N_21489,N_21233);
nor U22505 (N_22505,N_21002,N_21309);
and U22506 (N_22506,N_21245,N_21470);
nor U22507 (N_22507,N_21148,N_21843);
nor U22508 (N_22508,N_21277,N_21064);
nand U22509 (N_22509,N_21190,N_21698);
nand U22510 (N_22510,N_21009,N_21151);
xor U22511 (N_22511,N_21205,N_21654);
nor U22512 (N_22512,N_21675,N_21297);
or U22513 (N_22513,N_21262,N_21226);
nor U22514 (N_22514,N_21329,N_21041);
xnor U22515 (N_22515,N_21170,N_21562);
nand U22516 (N_22516,N_21760,N_21174);
or U22517 (N_22517,N_21277,N_21292);
xnor U22518 (N_22518,N_21075,N_21546);
xor U22519 (N_22519,N_21407,N_21990);
nand U22520 (N_22520,N_21283,N_21124);
nand U22521 (N_22521,N_21225,N_21157);
nor U22522 (N_22522,N_21325,N_21697);
or U22523 (N_22523,N_21362,N_21625);
or U22524 (N_22524,N_21150,N_21611);
nand U22525 (N_22525,N_21141,N_21427);
nand U22526 (N_22526,N_21443,N_21161);
nor U22527 (N_22527,N_21897,N_21127);
nand U22528 (N_22528,N_21191,N_21686);
xor U22529 (N_22529,N_21882,N_21451);
or U22530 (N_22530,N_21751,N_21979);
nor U22531 (N_22531,N_21087,N_21160);
nand U22532 (N_22532,N_21308,N_21567);
and U22533 (N_22533,N_21112,N_21295);
nand U22534 (N_22534,N_21304,N_21957);
nor U22535 (N_22535,N_21477,N_21228);
and U22536 (N_22536,N_21080,N_21176);
nand U22537 (N_22537,N_21398,N_21875);
nor U22538 (N_22538,N_21598,N_21871);
xor U22539 (N_22539,N_21574,N_21952);
nand U22540 (N_22540,N_21964,N_21624);
nor U22541 (N_22541,N_21921,N_21041);
xor U22542 (N_22542,N_21991,N_21737);
and U22543 (N_22543,N_21125,N_21103);
nand U22544 (N_22544,N_21388,N_21843);
or U22545 (N_22545,N_21055,N_21356);
nor U22546 (N_22546,N_21259,N_21361);
or U22547 (N_22547,N_21256,N_21471);
xor U22548 (N_22548,N_21237,N_21612);
nand U22549 (N_22549,N_21322,N_21209);
and U22550 (N_22550,N_21933,N_21742);
nand U22551 (N_22551,N_21773,N_21054);
nor U22552 (N_22552,N_21732,N_21600);
and U22553 (N_22553,N_21638,N_21540);
xor U22554 (N_22554,N_21119,N_21056);
xnor U22555 (N_22555,N_21131,N_21738);
nand U22556 (N_22556,N_21153,N_21290);
nor U22557 (N_22557,N_21289,N_21719);
and U22558 (N_22558,N_21230,N_21401);
nand U22559 (N_22559,N_21947,N_21221);
nand U22560 (N_22560,N_21811,N_21053);
nor U22561 (N_22561,N_21546,N_21464);
nand U22562 (N_22562,N_21322,N_21833);
and U22563 (N_22563,N_21924,N_21766);
nor U22564 (N_22564,N_21659,N_21258);
nand U22565 (N_22565,N_21568,N_21030);
nor U22566 (N_22566,N_21452,N_21550);
and U22567 (N_22567,N_21243,N_21961);
nand U22568 (N_22568,N_21410,N_21378);
and U22569 (N_22569,N_21727,N_21674);
or U22570 (N_22570,N_21348,N_21988);
or U22571 (N_22571,N_21885,N_21182);
or U22572 (N_22572,N_21067,N_21142);
nand U22573 (N_22573,N_21993,N_21170);
nand U22574 (N_22574,N_21905,N_21532);
nor U22575 (N_22575,N_21483,N_21304);
xor U22576 (N_22576,N_21954,N_21632);
nand U22577 (N_22577,N_21802,N_21474);
or U22578 (N_22578,N_21887,N_21640);
xnor U22579 (N_22579,N_21784,N_21699);
and U22580 (N_22580,N_21780,N_21924);
and U22581 (N_22581,N_21492,N_21313);
nand U22582 (N_22582,N_21882,N_21735);
and U22583 (N_22583,N_21474,N_21274);
nand U22584 (N_22584,N_21765,N_21454);
and U22585 (N_22585,N_21708,N_21450);
or U22586 (N_22586,N_21827,N_21264);
xor U22587 (N_22587,N_21503,N_21780);
xnor U22588 (N_22588,N_21414,N_21551);
nand U22589 (N_22589,N_21272,N_21328);
xnor U22590 (N_22590,N_21113,N_21260);
nor U22591 (N_22591,N_21400,N_21375);
xnor U22592 (N_22592,N_21656,N_21285);
nand U22593 (N_22593,N_21588,N_21480);
nor U22594 (N_22594,N_21757,N_21520);
or U22595 (N_22595,N_21663,N_21435);
and U22596 (N_22596,N_21853,N_21421);
and U22597 (N_22597,N_21215,N_21107);
and U22598 (N_22598,N_21098,N_21846);
and U22599 (N_22599,N_21301,N_21361);
nor U22600 (N_22600,N_21956,N_21914);
and U22601 (N_22601,N_21011,N_21467);
nor U22602 (N_22602,N_21163,N_21091);
xor U22603 (N_22603,N_21171,N_21078);
and U22604 (N_22604,N_21173,N_21305);
or U22605 (N_22605,N_21384,N_21339);
nand U22606 (N_22606,N_21286,N_21602);
and U22607 (N_22607,N_21369,N_21566);
and U22608 (N_22608,N_21361,N_21023);
and U22609 (N_22609,N_21231,N_21310);
xor U22610 (N_22610,N_21213,N_21399);
xor U22611 (N_22611,N_21045,N_21676);
xor U22612 (N_22612,N_21964,N_21122);
or U22613 (N_22613,N_21514,N_21193);
and U22614 (N_22614,N_21538,N_21773);
xor U22615 (N_22615,N_21035,N_21291);
and U22616 (N_22616,N_21409,N_21934);
and U22617 (N_22617,N_21574,N_21739);
nand U22618 (N_22618,N_21941,N_21294);
or U22619 (N_22619,N_21761,N_21979);
xnor U22620 (N_22620,N_21763,N_21168);
nor U22621 (N_22621,N_21595,N_21092);
xnor U22622 (N_22622,N_21976,N_21365);
nand U22623 (N_22623,N_21713,N_21940);
and U22624 (N_22624,N_21165,N_21958);
xor U22625 (N_22625,N_21692,N_21898);
and U22626 (N_22626,N_21842,N_21609);
nand U22627 (N_22627,N_21393,N_21333);
nand U22628 (N_22628,N_21422,N_21108);
or U22629 (N_22629,N_21260,N_21415);
xor U22630 (N_22630,N_21614,N_21549);
xnor U22631 (N_22631,N_21946,N_21654);
or U22632 (N_22632,N_21836,N_21504);
and U22633 (N_22633,N_21628,N_21855);
nand U22634 (N_22634,N_21902,N_21305);
and U22635 (N_22635,N_21357,N_21598);
and U22636 (N_22636,N_21656,N_21417);
and U22637 (N_22637,N_21273,N_21190);
nand U22638 (N_22638,N_21240,N_21770);
xor U22639 (N_22639,N_21538,N_21860);
nand U22640 (N_22640,N_21093,N_21606);
and U22641 (N_22641,N_21238,N_21272);
xor U22642 (N_22642,N_21237,N_21183);
and U22643 (N_22643,N_21720,N_21821);
and U22644 (N_22644,N_21767,N_21117);
and U22645 (N_22645,N_21034,N_21730);
nand U22646 (N_22646,N_21687,N_21276);
nor U22647 (N_22647,N_21722,N_21796);
nand U22648 (N_22648,N_21186,N_21394);
or U22649 (N_22649,N_21131,N_21027);
nand U22650 (N_22650,N_21279,N_21659);
and U22651 (N_22651,N_21805,N_21786);
nand U22652 (N_22652,N_21250,N_21292);
nor U22653 (N_22653,N_21530,N_21043);
or U22654 (N_22654,N_21849,N_21784);
or U22655 (N_22655,N_21001,N_21020);
and U22656 (N_22656,N_21699,N_21083);
or U22657 (N_22657,N_21718,N_21525);
and U22658 (N_22658,N_21772,N_21738);
or U22659 (N_22659,N_21732,N_21548);
or U22660 (N_22660,N_21114,N_21874);
nor U22661 (N_22661,N_21262,N_21951);
or U22662 (N_22662,N_21249,N_21050);
nand U22663 (N_22663,N_21402,N_21166);
nor U22664 (N_22664,N_21556,N_21078);
nor U22665 (N_22665,N_21053,N_21381);
xnor U22666 (N_22666,N_21326,N_21438);
and U22667 (N_22667,N_21681,N_21300);
nand U22668 (N_22668,N_21733,N_21430);
and U22669 (N_22669,N_21635,N_21851);
nor U22670 (N_22670,N_21333,N_21317);
xnor U22671 (N_22671,N_21430,N_21122);
xnor U22672 (N_22672,N_21529,N_21340);
or U22673 (N_22673,N_21952,N_21220);
and U22674 (N_22674,N_21129,N_21965);
xor U22675 (N_22675,N_21911,N_21278);
nor U22676 (N_22676,N_21620,N_21964);
xnor U22677 (N_22677,N_21293,N_21860);
or U22678 (N_22678,N_21469,N_21535);
nand U22679 (N_22679,N_21861,N_21903);
xnor U22680 (N_22680,N_21640,N_21114);
nor U22681 (N_22681,N_21478,N_21126);
xnor U22682 (N_22682,N_21714,N_21879);
nand U22683 (N_22683,N_21848,N_21605);
nand U22684 (N_22684,N_21449,N_21073);
nor U22685 (N_22685,N_21897,N_21539);
and U22686 (N_22686,N_21399,N_21013);
xor U22687 (N_22687,N_21437,N_21578);
xor U22688 (N_22688,N_21566,N_21319);
xor U22689 (N_22689,N_21154,N_21091);
and U22690 (N_22690,N_21923,N_21647);
and U22691 (N_22691,N_21299,N_21716);
or U22692 (N_22692,N_21682,N_21849);
nor U22693 (N_22693,N_21735,N_21342);
nand U22694 (N_22694,N_21650,N_21146);
nand U22695 (N_22695,N_21597,N_21784);
nand U22696 (N_22696,N_21503,N_21970);
xnor U22697 (N_22697,N_21375,N_21609);
xor U22698 (N_22698,N_21838,N_21508);
nor U22699 (N_22699,N_21916,N_21799);
or U22700 (N_22700,N_21731,N_21256);
or U22701 (N_22701,N_21603,N_21423);
xor U22702 (N_22702,N_21072,N_21817);
and U22703 (N_22703,N_21410,N_21343);
and U22704 (N_22704,N_21837,N_21085);
or U22705 (N_22705,N_21181,N_21411);
and U22706 (N_22706,N_21235,N_21021);
nor U22707 (N_22707,N_21068,N_21760);
nor U22708 (N_22708,N_21028,N_21013);
xnor U22709 (N_22709,N_21875,N_21400);
or U22710 (N_22710,N_21813,N_21278);
and U22711 (N_22711,N_21192,N_21988);
and U22712 (N_22712,N_21216,N_21441);
and U22713 (N_22713,N_21983,N_21728);
nand U22714 (N_22714,N_21951,N_21260);
nand U22715 (N_22715,N_21639,N_21665);
nor U22716 (N_22716,N_21193,N_21215);
nor U22717 (N_22717,N_21201,N_21478);
xnor U22718 (N_22718,N_21375,N_21015);
and U22719 (N_22719,N_21917,N_21507);
nor U22720 (N_22720,N_21558,N_21935);
or U22721 (N_22721,N_21989,N_21693);
nand U22722 (N_22722,N_21427,N_21657);
nor U22723 (N_22723,N_21484,N_21402);
or U22724 (N_22724,N_21348,N_21614);
and U22725 (N_22725,N_21282,N_21530);
or U22726 (N_22726,N_21243,N_21709);
or U22727 (N_22727,N_21300,N_21105);
and U22728 (N_22728,N_21408,N_21890);
and U22729 (N_22729,N_21475,N_21633);
or U22730 (N_22730,N_21773,N_21095);
and U22731 (N_22731,N_21989,N_21532);
nand U22732 (N_22732,N_21770,N_21877);
nand U22733 (N_22733,N_21510,N_21026);
and U22734 (N_22734,N_21582,N_21654);
nor U22735 (N_22735,N_21828,N_21107);
nor U22736 (N_22736,N_21705,N_21800);
and U22737 (N_22737,N_21778,N_21676);
xnor U22738 (N_22738,N_21997,N_21902);
or U22739 (N_22739,N_21117,N_21161);
and U22740 (N_22740,N_21918,N_21191);
or U22741 (N_22741,N_21540,N_21616);
xor U22742 (N_22742,N_21863,N_21913);
nor U22743 (N_22743,N_21802,N_21584);
and U22744 (N_22744,N_21371,N_21141);
or U22745 (N_22745,N_21447,N_21956);
nand U22746 (N_22746,N_21972,N_21431);
or U22747 (N_22747,N_21271,N_21821);
or U22748 (N_22748,N_21016,N_21640);
nor U22749 (N_22749,N_21755,N_21485);
nor U22750 (N_22750,N_21153,N_21771);
or U22751 (N_22751,N_21837,N_21759);
and U22752 (N_22752,N_21953,N_21494);
nor U22753 (N_22753,N_21578,N_21366);
nor U22754 (N_22754,N_21815,N_21655);
nand U22755 (N_22755,N_21619,N_21246);
and U22756 (N_22756,N_21515,N_21401);
or U22757 (N_22757,N_21302,N_21890);
or U22758 (N_22758,N_21998,N_21617);
and U22759 (N_22759,N_21695,N_21144);
nor U22760 (N_22760,N_21608,N_21286);
or U22761 (N_22761,N_21226,N_21299);
nor U22762 (N_22762,N_21612,N_21376);
nand U22763 (N_22763,N_21287,N_21672);
or U22764 (N_22764,N_21924,N_21840);
or U22765 (N_22765,N_21751,N_21898);
or U22766 (N_22766,N_21963,N_21461);
xnor U22767 (N_22767,N_21307,N_21063);
or U22768 (N_22768,N_21839,N_21728);
nor U22769 (N_22769,N_21568,N_21566);
nor U22770 (N_22770,N_21979,N_21285);
nand U22771 (N_22771,N_21666,N_21020);
nor U22772 (N_22772,N_21524,N_21642);
xor U22773 (N_22773,N_21770,N_21703);
or U22774 (N_22774,N_21660,N_21365);
xnor U22775 (N_22775,N_21733,N_21358);
and U22776 (N_22776,N_21494,N_21708);
nand U22777 (N_22777,N_21650,N_21161);
or U22778 (N_22778,N_21902,N_21906);
nor U22779 (N_22779,N_21260,N_21090);
or U22780 (N_22780,N_21138,N_21959);
xnor U22781 (N_22781,N_21386,N_21941);
xor U22782 (N_22782,N_21172,N_21181);
nor U22783 (N_22783,N_21125,N_21778);
nand U22784 (N_22784,N_21197,N_21092);
nand U22785 (N_22785,N_21982,N_21032);
or U22786 (N_22786,N_21951,N_21451);
or U22787 (N_22787,N_21456,N_21792);
and U22788 (N_22788,N_21090,N_21702);
nor U22789 (N_22789,N_21569,N_21978);
or U22790 (N_22790,N_21749,N_21721);
nand U22791 (N_22791,N_21041,N_21639);
and U22792 (N_22792,N_21708,N_21436);
nor U22793 (N_22793,N_21899,N_21315);
nor U22794 (N_22794,N_21562,N_21161);
nor U22795 (N_22795,N_21355,N_21422);
xor U22796 (N_22796,N_21385,N_21793);
or U22797 (N_22797,N_21073,N_21521);
xnor U22798 (N_22798,N_21709,N_21331);
and U22799 (N_22799,N_21548,N_21827);
or U22800 (N_22800,N_21961,N_21238);
nand U22801 (N_22801,N_21867,N_21936);
nor U22802 (N_22802,N_21830,N_21904);
or U22803 (N_22803,N_21610,N_21848);
xor U22804 (N_22804,N_21059,N_21540);
and U22805 (N_22805,N_21251,N_21643);
and U22806 (N_22806,N_21019,N_21729);
nand U22807 (N_22807,N_21886,N_21605);
and U22808 (N_22808,N_21165,N_21638);
or U22809 (N_22809,N_21697,N_21004);
or U22810 (N_22810,N_21336,N_21414);
and U22811 (N_22811,N_21466,N_21367);
xor U22812 (N_22812,N_21851,N_21768);
xnor U22813 (N_22813,N_21030,N_21132);
or U22814 (N_22814,N_21592,N_21193);
or U22815 (N_22815,N_21209,N_21132);
xnor U22816 (N_22816,N_21864,N_21427);
nand U22817 (N_22817,N_21127,N_21884);
and U22818 (N_22818,N_21356,N_21345);
nor U22819 (N_22819,N_21299,N_21522);
and U22820 (N_22820,N_21935,N_21096);
and U22821 (N_22821,N_21653,N_21913);
or U22822 (N_22822,N_21370,N_21028);
nand U22823 (N_22823,N_21983,N_21380);
nor U22824 (N_22824,N_21656,N_21721);
xor U22825 (N_22825,N_21061,N_21006);
nand U22826 (N_22826,N_21108,N_21715);
nand U22827 (N_22827,N_21218,N_21603);
or U22828 (N_22828,N_21266,N_21861);
and U22829 (N_22829,N_21177,N_21262);
and U22830 (N_22830,N_21989,N_21552);
xnor U22831 (N_22831,N_21467,N_21385);
nor U22832 (N_22832,N_21324,N_21920);
nor U22833 (N_22833,N_21461,N_21903);
nand U22834 (N_22834,N_21924,N_21171);
nand U22835 (N_22835,N_21655,N_21538);
or U22836 (N_22836,N_21730,N_21380);
nor U22837 (N_22837,N_21366,N_21249);
and U22838 (N_22838,N_21578,N_21860);
nor U22839 (N_22839,N_21594,N_21803);
and U22840 (N_22840,N_21889,N_21719);
or U22841 (N_22841,N_21426,N_21496);
xor U22842 (N_22842,N_21053,N_21050);
nand U22843 (N_22843,N_21251,N_21537);
and U22844 (N_22844,N_21836,N_21309);
nor U22845 (N_22845,N_21502,N_21835);
and U22846 (N_22846,N_21836,N_21982);
or U22847 (N_22847,N_21864,N_21984);
or U22848 (N_22848,N_21734,N_21472);
and U22849 (N_22849,N_21447,N_21966);
nor U22850 (N_22850,N_21833,N_21698);
or U22851 (N_22851,N_21298,N_21131);
xor U22852 (N_22852,N_21473,N_21983);
xnor U22853 (N_22853,N_21606,N_21862);
nand U22854 (N_22854,N_21586,N_21899);
or U22855 (N_22855,N_21077,N_21655);
and U22856 (N_22856,N_21179,N_21886);
nand U22857 (N_22857,N_21058,N_21845);
or U22858 (N_22858,N_21111,N_21388);
or U22859 (N_22859,N_21186,N_21666);
xnor U22860 (N_22860,N_21105,N_21674);
nor U22861 (N_22861,N_21986,N_21080);
nor U22862 (N_22862,N_21136,N_21397);
nor U22863 (N_22863,N_21464,N_21101);
nor U22864 (N_22864,N_21966,N_21408);
nand U22865 (N_22865,N_21047,N_21265);
and U22866 (N_22866,N_21533,N_21816);
and U22867 (N_22867,N_21627,N_21882);
xor U22868 (N_22868,N_21369,N_21338);
nor U22869 (N_22869,N_21693,N_21380);
xnor U22870 (N_22870,N_21507,N_21233);
or U22871 (N_22871,N_21130,N_21653);
xor U22872 (N_22872,N_21914,N_21288);
xnor U22873 (N_22873,N_21274,N_21263);
and U22874 (N_22874,N_21217,N_21420);
and U22875 (N_22875,N_21885,N_21705);
or U22876 (N_22876,N_21237,N_21880);
xnor U22877 (N_22877,N_21417,N_21589);
or U22878 (N_22878,N_21973,N_21829);
nor U22879 (N_22879,N_21386,N_21355);
xor U22880 (N_22880,N_21887,N_21742);
or U22881 (N_22881,N_21522,N_21122);
nor U22882 (N_22882,N_21261,N_21993);
and U22883 (N_22883,N_21584,N_21632);
or U22884 (N_22884,N_21510,N_21612);
nor U22885 (N_22885,N_21478,N_21826);
nor U22886 (N_22886,N_21658,N_21713);
and U22887 (N_22887,N_21923,N_21081);
nor U22888 (N_22888,N_21805,N_21209);
and U22889 (N_22889,N_21020,N_21194);
and U22890 (N_22890,N_21896,N_21795);
and U22891 (N_22891,N_21542,N_21175);
xor U22892 (N_22892,N_21888,N_21737);
or U22893 (N_22893,N_21944,N_21982);
and U22894 (N_22894,N_21240,N_21911);
and U22895 (N_22895,N_21240,N_21678);
xor U22896 (N_22896,N_21988,N_21609);
and U22897 (N_22897,N_21424,N_21432);
nor U22898 (N_22898,N_21243,N_21661);
nand U22899 (N_22899,N_21345,N_21458);
nand U22900 (N_22900,N_21533,N_21645);
xnor U22901 (N_22901,N_21382,N_21298);
and U22902 (N_22902,N_21151,N_21542);
xnor U22903 (N_22903,N_21636,N_21888);
nor U22904 (N_22904,N_21705,N_21934);
nor U22905 (N_22905,N_21654,N_21322);
xnor U22906 (N_22906,N_21357,N_21902);
nand U22907 (N_22907,N_21060,N_21878);
nor U22908 (N_22908,N_21454,N_21887);
xnor U22909 (N_22909,N_21736,N_21074);
or U22910 (N_22910,N_21309,N_21397);
and U22911 (N_22911,N_21779,N_21442);
nand U22912 (N_22912,N_21578,N_21423);
and U22913 (N_22913,N_21534,N_21497);
nor U22914 (N_22914,N_21941,N_21787);
nand U22915 (N_22915,N_21304,N_21528);
nor U22916 (N_22916,N_21041,N_21360);
xor U22917 (N_22917,N_21293,N_21143);
and U22918 (N_22918,N_21962,N_21754);
and U22919 (N_22919,N_21096,N_21028);
or U22920 (N_22920,N_21562,N_21583);
and U22921 (N_22921,N_21858,N_21633);
xor U22922 (N_22922,N_21577,N_21671);
and U22923 (N_22923,N_21018,N_21961);
and U22924 (N_22924,N_21012,N_21883);
nor U22925 (N_22925,N_21489,N_21801);
nor U22926 (N_22926,N_21069,N_21922);
nand U22927 (N_22927,N_21291,N_21310);
nor U22928 (N_22928,N_21325,N_21977);
nand U22929 (N_22929,N_21406,N_21504);
nor U22930 (N_22930,N_21637,N_21203);
xor U22931 (N_22931,N_21009,N_21460);
or U22932 (N_22932,N_21184,N_21599);
nand U22933 (N_22933,N_21155,N_21203);
or U22934 (N_22934,N_21991,N_21393);
nand U22935 (N_22935,N_21856,N_21876);
and U22936 (N_22936,N_21513,N_21227);
and U22937 (N_22937,N_21828,N_21098);
xnor U22938 (N_22938,N_21340,N_21693);
and U22939 (N_22939,N_21178,N_21240);
xnor U22940 (N_22940,N_21532,N_21855);
xnor U22941 (N_22941,N_21206,N_21114);
nor U22942 (N_22942,N_21088,N_21676);
nand U22943 (N_22943,N_21402,N_21790);
nor U22944 (N_22944,N_21347,N_21134);
xor U22945 (N_22945,N_21665,N_21575);
nor U22946 (N_22946,N_21727,N_21486);
nor U22947 (N_22947,N_21871,N_21402);
nor U22948 (N_22948,N_21665,N_21808);
and U22949 (N_22949,N_21417,N_21225);
xnor U22950 (N_22950,N_21269,N_21128);
or U22951 (N_22951,N_21656,N_21048);
nor U22952 (N_22952,N_21879,N_21353);
or U22953 (N_22953,N_21461,N_21322);
xnor U22954 (N_22954,N_21770,N_21796);
or U22955 (N_22955,N_21052,N_21151);
and U22956 (N_22956,N_21563,N_21095);
xor U22957 (N_22957,N_21531,N_21425);
nand U22958 (N_22958,N_21598,N_21257);
or U22959 (N_22959,N_21042,N_21027);
or U22960 (N_22960,N_21466,N_21952);
nor U22961 (N_22961,N_21029,N_21576);
or U22962 (N_22962,N_21993,N_21829);
nor U22963 (N_22963,N_21859,N_21093);
xor U22964 (N_22964,N_21224,N_21501);
nand U22965 (N_22965,N_21819,N_21552);
or U22966 (N_22966,N_21827,N_21636);
nand U22967 (N_22967,N_21965,N_21587);
nand U22968 (N_22968,N_21191,N_21469);
and U22969 (N_22969,N_21080,N_21085);
and U22970 (N_22970,N_21567,N_21762);
or U22971 (N_22971,N_21380,N_21665);
or U22972 (N_22972,N_21049,N_21379);
and U22973 (N_22973,N_21538,N_21244);
and U22974 (N_22974,N_21881,N_21406);
or U22975 (N_22975,N_21390,N_21601);
or U22976 (N_22976,N_21570,N_21356);
nor U22977 (N_22977,N_21865,N_21264);
or U22978 (N_22978,N_21000,N_21620);
nand U22979 (N_22979,N_21763,N_21871);
and U22980 (N_22980,N_21948,N_21432);
nand U22981 (N_22981,N_21398,N_21326);
nor U22982 (N_22982,N_21973,N_21581);
xnor U22983 (N_22983,N_21559,N_21397);
nand U22984 (N_22984,N_21807,N_21131);
and U22985 (N_22985,N_21794,N_21965);
nor U22986 (N_22986,N_21969,N_21037);
nor U22987 (N_22987,N_21483,N_21936);
and U22988 (N_22988,N_21762,N_21481);
nor U22989 (N_22989,N_21509,N_21751);
and U22990 (N_22990,N_21212,N_21202);
xnor U22991 (N_22991,N_21196,N_21186);
xor U22992 (N_22992,N_21715,N_21671);
and U22993 (N_22993,N_21382,N_21316);
or U22994 (N_22994,N_21608,N_21344);
or U22995 (N_22995,N_21110,N_21920);
and U22996 (N_22996,N_21859,N_21655);
nand U22997 (N_22997,N_21631,N_21143);
xor U22998 (N_22998,N_21180,N_21496);
nand U22999 (N_22999,N_21080,N_21261);
xor U23000 (N_23000,N_22244,N_22669);
nand U23001 (N_23001,N_22896,N_22114);
nor U23002 (N_23002,N_22163,N_22905);
xor U23003 (N_23003,N_22290,N_22561);
nand U23004 (N_23004,N_22463,N_22128);
nand U23005 (N_23005,N_22493,N_22357);
nor U23006 (N_23006,N_22386,N_22331);
xor U23007 (N_23007,N_22547,N_22122);
xor U23008 (N_23008,N_22292,N_22639);
or U23009 (N_23009,N_22974,N_22057);
nor U23010 (N_23010,N_22693,N_22278);
nor U23011 (N_23011,N_22123,N_22619);
xor U23012 (N_23012,N_22069,N_22954);
and U23013 (N_23013,N_22621,N_22439);
nand U23014 (N_23014,N_22470,N_22835);
xnor U23015 (N_23015,N_22277,N_22403);
nor U23016 (N_23016,N_22207,N_22537);
nor U23017 (N_23017,N_22409,N_22883);
or U23018 (N_23018,N_22016,N_22670);
xnor U23019 (N_23019,N_22127,N_22713);
or U23020 (N_23020,N_22592,N_22526);
and U23021 (N_23021,N_22906,N_22364);
nor U23022 (N_23022,N_22134,N_22600);
xnor U23023 (N_23023,N_22838,N_22220);
and U23024 (N_23024,N_22106,N_22732);
or U23025 (N_23025,N_22646,N_22901);
xnor U23026 (N_23026,N_22170,N_22869);
and U23027 (N_23027,N_22973,N_22860);
xnor U23028 (N_23028,N_22807,N_22475);
xnor U23029 (N_23029,N_22831,N_22532);
and U23030 (N_23030,N_22994,N_22897);
and U23031 (N_23031,N_22792,N_22744);
and U23032 (N_23032,N_22485,N_22446);
xnor U23033 (N_23033,N_22109,N_22243);
nor U23034 (N_23034,N_22614,N_22967);
nand U23035 (N_23035,N_22242,N_22467);
nor U23036 (N_23036,N_22022,N_22024);
xnor U23037 (N_23037,N_22484,N_22859);
nand U23038 (N_23038,N_22260,N_22136);
xnor U23039 (N_23039,N_22236,N_22714);
and U23040 (N_23040,N_22779,N_22202);
xnor U23041 (N_23041,N_22487,N_22165);
xnor U23042 (N_23042,N_22917,N_22519);
and U23043 (N_23043,N_22179,N_22815);
or U23044 (N_23044,N_22118,N_22448);
and U23045 (N_23045,N_22960,N_22011);
or U23046 (N_23046,N_22461,N_22706);
xnor U23047 (N_23047,N_22410,N_22098);
nor U23048 (N_23048,N_22015,N_22794);
nand U23049 (N_23049,N_22054,N_22237);
nand U23050 (N_23050,N_22301,N_22340);
and U23051 (N_23051,N_22483,N_22751);
and U23052 (N_23052,N_22727,N_22328);
xor U23053 (N_23053,N_22767,N_22125);
nand U23054 (N_23054,N_22650,N_22817);
nand U23055 (N_23055,N_22394,N_22846);
or U23056 (N_23056,N_22628,N_22658);
and U23057 (N_23057,N_22629,N_22685);
nand U23058 (N_23058,N_22848,N_22659);
and U23059 (N_23059,N_22987,N_22647);
or U23060 (N_23060,N_22262,N_22212);
nand U23061 (N_23061,N_22030,N_22186);
xor U23062 (N_23062,N_22655,N_22888);
nor U23063 (N_23063,N_22983,N_22351);
nand U23064 (N_23064,N_22197,N_22059);
nor U23065 (N_23065,N_22456,N_22551);
nor U23066 (N_23066,N_22944,N_22874);
xnor U23067 (N_23067,N_22607,N_22490);
nand U23068 (N_23068,N_22512,N_22899);
xor U23069 (N_23069,N_22821,N_22985);
and U23070 (N_23070,N_22230,N_22460);
xor U23071 (N_23071,N_22427,N_22316);
or U23072 (N_23072,N_22671,N_22667);
xor U23073 (N_23073,N_22133,N_22677);
nand U23074 (N_23074,N_22454,N_22653);
xor U23075 (N_23075,N_22847,N_22044);
xor U23076 (N_23076,N_22472,N_22080);
or U23077 (N_23077,N_22257,N_22157);
nor U23078 (N_23078,N_22405,N_22689);
or U23079 (N_23079,N_22238,N_22267);
nand U23080 (N_23080,N_22712,N_22595);
nor U23081 (N_23081,N_22217,N_22661);
or U23082 (N_23082,N_22963,N_22434);
nor U23083 (N_23083,N_22842,N_22618);
or U23084 (N_23084,N_22458,N_22012);
nor U23085 (N_23085,N_22844,N_22418);
nand U23086 (N_23086,N_22604,N_22552);
or U23087 (N_23087,N_22545,N_22746);
or U23088 (N_23088,N_22310,N_22766);
and U23089 (N_23089,N_22092,N_22222);
or U23090 (N_23090,N_22353,N_22910);
xor U23091 (N_23091,N_22715,N_22201);
xor U23092 (N_23092,N_22797,N_22895);
or U23093 (N_23093,N_22969,N_22249);
nor U23094 (N_23094,N_22749,N_22450);
or U23095 (N_23095,N_22793,N_22005);
xor U23096 (N_23096,N_22337,N_22473);
and U23097 (N_23097,N_22681,N_22912);
xnor U23098 (N_23098,N_22943,N_22162);
nor U23099 (N_23099,N_22980,N_22853);
nand U23100 (N_23100,N_22644,N_22977);
nor U23101 (N_23101,N_22900,N_22088);
nand U23102 (N_23102,N_22754,N_22185);
and U23103 (N_23103,N_22705,N_22199);
xnor U23104 (N_23104,N_22708,N_22465);
or U23105 (N_23105,N_22914,N_22579);
and U23106 (N_23106,N_22272,N_22510);
and U23107 (N_23107,N_22582,N_22726);
xor U23108 (N_23108,N_22503,N_22096);
nand U23109 (N_23109,N_22697,N_22298);
or U23110 (N_23110,N_22025,N_22297);
or U23111 (N_23111,N_22389,N_22840);
xnor U23112 (N_23112,N_22599,N_22145);
nor U23113 (N_23113,N_22589,N_22733);
and U23114 (N_23114,N_22919,N_22362);
or U23115 (N_23115,N_22894,N_22884);
or U23116 (N_23116,N_22887,N_22303);
and U23117 (N_23117,N_22314,N_22507);
nand U23118 (N_23118,N_22055,N_22701);
or U23119 (N_23119,N_22221,N_22986);
nor U23120 (N_23120,N_22245,N_22940);
and U23121 (N_23121,N_22391,N_22802);
or U23122 (N_23122,N_22023,N_22839);
and U23123 (N_23123,N_22956,N_22882);
xnor U23124 (N_23124,N_22769,N_22097);
xor U23125 (N_23125,N_22190,N_22375);
nor U23126 (N_23126,N_22094,N_22319);
or U23127 (N_23127,N_22181,N_22989);
xnor U23128 (N_23128,N_22227,N_22971);
nand U23129 (N_23129,N_22892,N_22739);
and U23130 (N_23130,N_22823,N_22610);
nand U23131 (N_23131,N_22730,N_22160);
xor U23132 (N_23132,N_22654,N_22570);
or U23133 (N_23133,N_22388,N_22327);
or U23134 (N_23134,N_22982,N_22194);
xor U23135 (N_23135,N_22111,N_22077);
and U23136 (N_23136,N_22294,N_22567);
or U23137 (N_23137,N_22379,N_22945);
xor U23138 (N_23138,N_22790,N_22332);
nand U23139 (N_23139,N_22756,N_22735);
or U23140 (N_23140,N_22393,N_22976);
nor U23141 (N_23141,N_22430,N_22010);
and U23142 (N_23142,N_22696,N_22398);
and U23143 (N_23143,N_22431,N_22368);
xor U23144 (N_23144,N_22466,N_22642);
nand U23145 (N_23145,N_22514,N_22281);
or U23146 (N_23146,N_22166,N_22075);
nor U23147 (N_23147,N_22304,N_22371);
and U23148 (N_23148,N_22288,N_22192);
xnor U23149 (N_23149,N_22593,N_22759);
xnor U23150 (N_23150,N_22033,N_22755);
and U23151 (N_23151,N_22486,N_22280);
nor U23152 (N_23152,N_22284,N_22648);
or U23153 (N_23153,N_22862,N_22521);
xor U23154 (N_23154,N_22326,N_22259);
nand U23155 (N_23155,N_22343,N_22949);
or U23156 (N_23156,N_22529,N_22341);
nand U23157 (N_23157,N_22694,N_22235);
and U23158 (N_23158,N_22908,N_22401);
and U23159 (N_23159,N_22468,N_22496);
or U23160 (N_23160,N_22921,N_22013);
nand U23161 (N_23161,N_22355,N_22711);
nand U23162 (N_23162,N_22999,N_22348);
nand U23163 (N_23163,N_22336,N_22066);
or U23164 (N_23164,N_22482,N_22680);
and U23165 (N_23165,N_22035,N_22443);
xnor U23166 (N_23166,N_22966,N_22876);
or U23167 (N_23167,N_22345,N_22953);
nor U23168 (N_23168,N_22885,N_22110);
nor U23169 (N_23169,N_22675,N_22904);
and U23170 (N_23170,N_22499,N_22923);
xnor U23171 (N_23171,N_22911,N_22494);
or U23172 (N_23172,N_22652,N_22232);
xor U23173 (N_23173,N_22951,N_22620);
nand U23174 (N_23174,N_22826,N_22682);
nor U23175 (N_23175,N_22084,N_22400);
nor U23176 (N_23176,N_22692,N_22959);
nand U23177 (N_23177,N_22038,N_22104);
or U23178 (N_23178,N_22891,N_22935);
and U23179 (N_23179,N_22662,N_22979);
and U23180 (N_23180,N_22928,N_22285);
and U23181 (N_23181,N_22083,N_22086);
and U23182 (N_23182,N_22700,N_22852);
nand U23183 (N_23183,N_22676,N_22073);
nor U23184 (N_23184,N_22287,N_22598);
nand U23185 (N_23185,N_22383,N_22783);
nand U23186 (N_23186,N_22760,N_22736);
or U23187 (N_23187,N_22991,N_22143);
xnor U23188 (N_23188,N_22441,N_22832);
nand U23189 (N_23189,N_22528,N_22218);
or U23190 (N_23190,N_22556,N_22695);
nor U23191 (N_23191,N_22321,N_22256);
or U23192 (N_23192,N_22742,N_22435);
xor U23193 (N_23193,N_22141,N_22812);
xnor U23194 (N_23194,N_22602,N_22672);
and U23195 (N_23195,N_22034,N_22861);
nand U23196 (N_23196,N_22215,N_22572);
and U23197 (N_23197,N_22274,N_22890);
nand U23198 (N_23198,N_22381,N_22455);
or U23199 (N_23199,N_22037,N_22497);
or U23200 (N_23200,N_22268,N_22698);
nor U23201 (N_23201,N_22481,N_22845);
nand U23202 (N_23202,N_22723,N_22729);
or U23203 (N_23203,N_22469,N_22703);
nand U23204 (N_23204,N_22995,N_22725);
or U23205 (N_23205,N_22007,N_22413);
nand U23206 (N_23206,N_22827,N_22524);
and U23207 (N_23207,N_22153,N_22990);
and U23208 (N_23208,N_22131,N_22169);
and U23209 (N_23209,N_22219,N_22154);
nor U23210 (N_23210,N_22254,N_22253);
and U23211 (N_23211,N_22178,N_22741);
and U23212 (N_23212,N_22523,N_22382);
and U23213 (N_23213,N_22422,N_22877);
or U23214 (N_23214,N_22651,N_22854);
nand U23215 (N_23215,N_22056,N_22031);
and U23216 (N_23216,N_22563,N_22590);
nand U23217 (N_23217,N_22116,N_22631);
nand U23218 (N_23218,N_22216,N_22509);
nor U23219 (N_23219,N_22189,N_22541);
and U23220 (N_23220,N_22863,N_22691);
and U23221 (N_23221,N_22932,N_22565);
xnor U23222 (N_23222,N_22006,N_22323);
and U23223 (N_23223,N_22615,N_22471);
or U23224 (N_23224,N_22603,N_22085);
and U23225 (N_23225,N_22550,N_22231);
xnor U23226 (N_23226,N_22063,N_22338);
nand U23227 (N_23227,N_22295,N_22402);
and U23228 (N_23228,N_22018,N_22941);
nand U23229 (N_23229,N_22071,N_22040);
nor U23230 (N_23230,N_22571,N_22089);
and U23231 (N_23231,N_22188,N_22922);
and U23232 (N_23232,N_22506,N_22819);
nor U23233 (N_23233,N_22805,N_22168);
xnor U23234 (N_23234,N_22775,N_22252);
nor U23235 (N_23235,N_22738,N_22058);
or U23236 (N_23236,N_22183,N_22993);
or U23237 (N_23237,N_22330,N_22029);
or U23238 (N_23238,N_22067,N_22717);
and U23239 (N_23239,N_22346,N_22569);
nor U23240 (N_23240,N_22907,N_22968);
nand U23241 (N_23241,N_22873,N_22743);
nand U23242 (N_23242,N_22074,N_22502);
and U23243 (N_23243,N_22009,N_22788);
nor U23244 (N_23244,N_22004,N_22442);
xor U23245 (N_23245,N_22665,N_22539);
nor U23246 (N_23246,N_22833,N_22830);
or U23247 (N_23247,N_22271,N_22702);
xor U23248 (N_23248,N_22273,N_22246);
nor U23249 (N_23249,N_22119,N_22961);
nand U23250 (N_23250,N_22684,N_22938);
nor U23251 (N_23251,N_22302,N_22308);
and U23252 (N_23252,N_22061,N_22361);
xnor U23253 (N_23253,N_22228,N_22344);
xnor U23254 (N_23254,N_22881,N_22462);
or U23255 (N_23255,N_22734,N_22180);
nand U23256 (N_23256,N_22645,N_22606);
and U23257 (N_23257,N_22198,N_22666);
and U23258 (N_23258,N_22660,N_22791);
nor U23259 (N_23259,N_22924,N_22079);
and U23260 (N_23260,N_22584,N_22200);
nand U23261 (N_23261,N_22206,N_22320);
nor U23262 (N_23262,N_22078,N_22070);
nor U23263 (N_23263,N_22930,N_22837);
or U23264 (N_23264,N_22453,N_22449);
and U23265 (N_23265,N_22474,N_22177);
or U23266 (N_23266,N_22047,N_22637);
nor U23267 (N_23267,N_22359,N_22421);
or U23268 (N_23268,N_22709,N_22477);
nor U23269 (N_23269,N_22605,N_22082);
xnor U23270 (N_23270,N_22927,N_22313);
or U23271 (N_23271,N_22390,N_22126);
xnor U23272 (N_23272,N_22039,N_22491);
nor U23273 (N_23273,N_22184,N_22611);
nand U23274 (N_23274,N_22886,N_22624);
nand U23275 (N_23275,N_22534,N_22356);
xor U23276 (N_23276,N_22289,N_22656);
and U23277 (N_23277,N_22064,N_22370);
nand U23278 (N_23278,N_22360,N_22223);
nand U23279 (N_23279,N_22801,N_22596);
or U23280 (N_23280,N_22609,N_22857);
nand U23281 (N_23281,N_22668,N_22002);
nor U23282 (N_23282,N_22003,N_22574);
xor U23283 (N_23283,N_22630,N_22091);
nand U23284 (N_23284,N_22750,N_22722);
xor U23285 (N_23285,N_22334,N_22772);
and U23286 (N_23286,N_22553,N_22478);
xor U23287 (N_23287,N_22374,N_22315);
nor U23288 (N_23288,N_22452,N_22001);
and U23289 (N_23289,N_22411,N_22377);
nand U23290 (N_23290,N_22120,N_22538);
xnor U23291 (N_23291,N_22311,N_22934);
nor U23292 (N_23292,N_22690,N_22947);
xnor U23293 (N_23293,N_22798,N_22404);
xor U23294 (N_23294,N_22972,N_22417);
xnor U23295 (N_23295,N_22804,N_22814);
nand U23296 (N_23296,N_22585,N_22283);
and U23297 (N_23297,N_22841,N_22781);
or U23298 (N_23298,N_22543,N_22740);
xor U23299 (N_23299,N_22581,N_22721);
and U23300 (N_23300,N_22597,N_22822);
and U23301 (N_23301,N_22988,N_22363);
xor U23302 (N_23302,N_22420,N_22042);
xor U23303 (N_23303,N_22027,N_22352);
nand U23304 (N_23304,N_22785,N_22195);
and U23305 (N_23305,N_22021,N_22796);
or U23306 (N_23306,N_22335,N_22350);
nor U23307 (N_23307,N_22366,N_22053);
and U23308 (N_23308,N_22121,N_22445);
nor U23309 (N_23309,N_22770,N_22043);
and U23310 (N_23310,N_22850,N_22488);
and U23311 (N_23311,N_22856,N_22636);
nand U23312 (N_23312,N_22210,N_22171);
nand U23313 (N_23313,N_22699,N_22554);
nand U23314 (N_23314,N_22041,N_22265);
xor U23315 (N_23315,N_22107,N_22834);
nor U23316 (N_23316,N_22204,N_22557);
xnor U23317 (N_23317,N_22981,N_22312);
and U23318 (N_23318,N_22673,N_22432);
xnor U23319 (N_23319,N_22925,N_22492);
nand U23320 (N_23320,N_22447,N_22763);
nor U23321 (N_23321,N_22076,N_22889);
and U23322 (N_23322,N_22373,N_22419);
and U23323 (N_23323,N_22719,N_22992);
xnor U23324 (N_23324,N_22777,N_22385);
nand U23325 (N_23325,N_22437,N_22436);
and U23326 (N_23326,N_22208,N_22898);
xor U23327 (N_23327,N_22933,N_22778);
nor U23328 (N_23328,N_22587,N_22068);
nand U23329 (N_23329,N_22247,N_22229);
nand U23330 (N_23330,N_22000,N_22975);
xor U23331 (N_23331,N_22872,N_22263);
and U23332 (N_23332,N_22558,N_22451);
and U23333 (N_23333,N_22014,N_22573);
or U23334 (N_23334,N_22588,N_22578);
nor U23335 (N_23335,N_22564,N_22372);
nor U23336 (N_23336,N_22132,N_22099);
or U23337 (N_23337,N_22984,N_22129);
nor U23338 (N_23338,N_22008,N_22929);
nand U23339 (N_23339,N_22544,N_22789);
nand U23340 (N_23340,N_22540,N_22962);
xnor U23341 (N_23341,N_22048,N_22151);
nor U23342 (N_23342,N_22635,N_22851);
xor U23343 (N_23343,N_22376,N_22396);
nor U23344 (N_23344,N_22867,N_22757);
nand U23345 (N_23345,N_22081,N_22317);
xnor U23346 (N_23346,N_22731,N_22423);
nor U23347 (N_23347,N_22358,N_22060);
xnor U23348 (N_23348,N_22322,N_22264);
xor U23349 (N_23349,N_22625,N_22580);
or U23350 (N_23350,N_22365,N_22875);
xnor U23351 (N_23351,N_22276,N_22286);
xnor U23352 (N_23352,N_22148,N_22918);
xor U23353 (N_23353,N_22810,N_22638);
or U23354 (N_23354,N_22296,N_22480);
and U23355 (N_23355,N_22771,N_22761);
nand U23356 (N_23356,N_22601,N_22633);
and U23357 (N_23357,N_22517,N_22150);
nand U23358 (N_23358,N_22809,N_22787);
or U23359 (N_23359,N_22130,N_22065);
or U23360 (N_23360,N_22843,N_22498);
or U23361 (N_23361,N_22258,N_22586);
or U23362 (N_23362,N_22028,N_22307);
nor U23363 (N_23363,N_22146,N_22535);
nand U23364 (N_23364,N_22026,N_22641);
xnor U23365 (N_23365,N_22270,N_22158);
and U23366 (N_23366,N_22138,N_22542);
nand U23367 (N_23367,N_22248,N_22868);
or U23368 (N_23368,N_22479,N_22623);
nor U23369 (N_23369,N_22046,N_22407);
or U23370 (N_23370,N_22627,N_22428);
nand U23371 (N_23371,N_22384,N_22515);
and U23372 (N_23372,N_22634,N_22864);
or U23373 (N_23373,N_22632,N_22855);
or U23374 (N_23374,N_22902,N_22415);
nor U23375 (N_23375,N_22926,N_22347);
nand U23376 (N_23376,N_22626,N_22191);
or U23377 (N_23377,N_22870,N_22576);
nand U23378 (N_23378,N_22032,N_22103);
xor U23379 (N_23379,N_22559,N_22704);
xnor U23380 (N_23380,N_22108,N_22978);
nand U23381 (N_23381,N_22594,N_22836);
nand U23382 (N_23382,N_22871,N_22664);
or U23383 (N_23383,N_22957,N_22858);
and U23384 (N_23384,N_22019,N_22829);
or U23385 (N_23385,N_22500,N_22806);
and U23386 (N_23386,N_22737,N_22017);
nor U23387 (N_23387,N_22768,N_22282);
xnor U23388 (N_23388,N_22747,N_22142);
or U23389 (N_23389,N_22795,N_22250);
or U23390 (N_23390,N_22459,N_22224);
nand U23391 (N_23391,N_22147,N_22367);
or U23392 (N_23392,N_22354,N_22920);
or U23393 (N_23393,N_22205,N_22765);
nor U23394 (N_23394,N_22786,N_22879);
nor U23395 (N_23395,N_22530,N_22511);
and U23396 (N_23396,N_22213,N_22780);
or U23397 (N_23397,N_22239,N_22279);
and U23398 (N_23398,N_22566,N_22516);
and U23399 (N_23399,N_22102,N_22764);
or U23400 (N_23400,N_22996,N_22758);
xnor U23401 (N_23401,N_22679,N_22489);
and U23402 (N_23402,N_22718,N_22965);
xor U23403 (N_23403,N_22115,N_22309);
and U23404 (N_23404,N_22800,N_22062);
nand U23405 (N_23405,N_22745,N_22051);
nor U23406 (N_23406,N_22903,N_22406);
and U23407 (N_23407,N_22050,N_22617);
xnor U23408 (N_23408,N_22657,N_22090);
and U23409 (N_23409,N_22997,N_22349);
nand U23410 (N_23410,N_22612,N_22525);
nor U23411 (N_23411,N_22339,N_22172);
or U23412 (N_23412,N_22329,N_22369);
xor U23413 (N_23413,N_22955,N_22608);
and U23414 (N_23414,N_22137,N_22531);
xnor U23415 (N_23415,N_22513,N_22378);
nor U23416 (N_23416,N_22380,N_22139);
xnor U23417 (N_23417,N_22225,N_22438);
and U23418 (N_23418,N_22266,N_22416);
xor U23419 (N_23419,N_22426,N_22164);
nand U23420 (N_23420,N_22408,N_22762);
nand U23421 (N_23421,N_22549,N_22240);
nand U23422 (N_23422,N_22187,N_22209);
or U23423 (N_23423,N_22562,N_22176);
nand U23424 (N_23424,N_22156,N_22520);
or U23425 (N_23425,N_22583,N_22135);
nor U23426 (N_23426,N_22942,N_22970);
nor U23427 (N_23427,N_22649,N_22049);
or U23428 (N_23428,N_22707,N_22144);
or U23429 (N_23429,N_22808,N_22117);
nand U23430 (N_23430,N_22211,N_22964);
xnor U23431 (N_23431,N_22952,N_22299);
nor U23432 (N_23432,N_22774,N_22203);
and U23433 (N_23433,N_22261,N_22752);
or U23434 (N_23434,N_22683,N_22577);
nor U23435 (N_23435,N_22939,N_22306);
and U23436 (N_23436,N_22936,N_22174);
nor U23437 (N_23437,N_22782,N_22728);
xor U23438 (N_23438,N_22533,N_22811);
and U23439 (N_23439,N_22916,N_22504);
nand U23440 (N_23440,N_22878,N_22546);
nand U23441 (N_23441,N_22214,N_22568);
nand U23442 (N_23442,N_22226,N_22865);
xnor U23443 (N_23443,N_22958,N_22342);
nor U23444 (N_23444,N_22036,N_22395);
nand U23445 (N_23445,N_22182,N_22175);
nand U23446 (N_23446,N_22687,N_22255);
nor U23447 (N_23447,N_22101,N_22816);
xnor U23448 (N_23448,N_22152,N_22622);
nor U23449 (N_23449,N_22444,N_22616);
nor U23450 (N_23450,N_22196,N_22536);
or U23451 (N_23451,N_22575,N_22518);
and U23452 (N_23452,N_22909,N_22849);
nor U23453 (N_23453,N_22663,N_22776);
xor U23454 (N_23454,N_22560,N_22155);
nor U23455 (N_23455,N_22020,N_22440);
nor U23456 (N_23456,N_22140,N_22159);
xnor U23457 (N_23457,N_22397,N_22464);
xor U23458 (N_23458,N_22052,N_22674);
nor U23459 (N_23459,N_22325,N_22799);
and U23460 (N_23460,N_22613,N_22476);
or U23461 (N_23461,N_22501,N_22784);
nand U23462 (N_23462,N_22946,N_22045);
and U23463 (N_23463,N_22591,N_22710);
or U23464 (N_23464,N_22112,N_22748);
or U23465 (N_23465,N_22087,N_22813);
xnor U23466 (N_23466,N_22998,N_22724);
nor U23467 (N_23467,N_22866,N_22716);
xor U23468 (N_23468,N_22173,N_22399);
or U23469 (N_23469,N_22234,N_22251);
or U23470 (N_23470,N_22291,N_22167);
nand U23471 (N_23471,N_22233,N_22548);
nor U23472 (N_23472,N_22429,N_22149);
or U23473 (N_23473,N_22318,N_22773);
nor U23474 (N_23474,N_22269,N_22161);
xnor U23475 (N_23475,N_22424,N_22275);
nor U23476 (N_23476,N_22495,N_22113);
or U23477 (N_23477,N_22324,N_22937);
xnor U23478 (N_23478,N_22640,N_22893);
nor U23479 (N_23479,N_22555,N_22124);
and U23480 (N_23480,N_22688,N_22948);
xor U23481 (N_23481,N_22508,N_22803);
and U23482 (N_23482,N_22824,N_22950);
nor U23483 (N_23483,N_22720,N_22425);
and U23484 (N_23484,N_22505,N_22880);
and U23485 (N_23485,N_22333,N_22825);
nor U23486 (N_23486,N_22093,N_22931);
nand U23487 (N_23487,N_22527,N_22392);
or U23488 (N_23488,N_22105,N_22293);
nand U23489 (N_23489,N_22305,N_22433);
or U23490 (N_23490,N_22300,N_22522);
and U23491 (N_23491,N_22072,N_22387);
or U23492 (N_23492,N_22095,N_22678);
xnor U23493 (N_23493,N_22818,N_22457);
xnor U23494 (N_23494,N_22686,N_22414);
xor U23495 (N_23495,N_22193,N_22915);
and U23496 (N_23496,N_22820,N_22913);
nor U23497 (N_23497,N_22753,N_22643);
and U23498 (N_23498,N_22241,N_22412);
and U23499 (N_23499,N_22100,N_22828);
and U23500 (N_23500,N_22797,N_22648);
nor U23501 (N_23501,N_22009,N_22593);
and U23502 (N_23502,N_22085,N_22571);
nand U23503 (N_23503,N_22954,N_22242);
and U23504 (N_23504,N_22000,N_22192);
nor U23505 (N_23505,N_22894,N_22037);
nor U23506 (N_23506,N_22200,N_22803);
nor U23507 (N_23507,N_22776,N_22190);
nand U23508 (N_23508,N_22153,N_22365);
xnor U23509 (N_23509,N_22355,N_22047);
nor U23510 (N_23510,N_22288,N_22256);
xnor U23511 (N_23511,N_22607,N_22454);
xnor U23512 (N_23512,N_22392,N_22300);
or U23513 (N_23513,N_22372,N_22063);
xor U23514 (N_23514,N_22460,N_22822);
nor U23515 (N_23515,N_22437,N_22443);
and U23516 (N_23516,N_22273,N_22221);
xor U23517 (N_23517,N_22377,N_22384);
nor U23518 (N_23518,N_22284,N_22139);
and U23519 (N_23519,N_22556,N_22950);
or U23520 (N_23520,N_22496,N_22162);
or U23521 (N_23521,N_22948,N_22325);
nand U23522 (N_23522,N_22656,N_22660);
nand U23523 (N_23523,N_22583,N_22551);
or U23524 (N_23524,N_22778,N_22163);
nor U23525 (N_23525,N_22514,N_22105);
and U23526 (N_23526,N_22876,N_22649);
nor U23527 (N_23527,N_22156,N_22185);
and U23528 (N_23528,N_22956,N_22931);
or U23529 (N_23529,N_22636,N_22021);
nor U23530 (N_23530,N_22743,N_22135);
and U23531 (N_23531,N_22148,N_22342);
nand U23532 (N_23532,N_22569,N_22486);
nor U23533 (N_23533,N_22414,N_22843);
and U23534 (N_23534,N_22113,N_22345);
xor U23535 (N_23535,N_22182,N_22790);
and U23536 (N_23536,N_22981,N_22679);
nor U23537 (N_23537,N_22121,N_22527);
nand U23538 (N_23538,N_22076,N_22551);
or U23539 (N_23539,N_22755,N_22538);
nor U23540 (N_23540,N_22494,N_22997);
nand U23541 (N_23541,N_22921,N_22706);
xor U23542 (N_23542,N_22104,N_22147);
nand U23543 (N_23543,N_22799,N_22693);
nand U23544 (N_23544,N_22219,N_22004);
and U23545 (N_23545,N_22801,N_22606);
nand U23546 (N_23546,N_22085,N_22771);
nand U23547 (N_23547,N_22742,N_22581);
or U23548 (N_23548,N_22569,N_22531);
and U23549 (N_23549,N_22129,N_22119);
nand U23550 (N_23550,N_22893,N_22189);
nand U23551 (N_23551,N_22382,N_22271);
nor U23552 (N_23552,N_22718,N_22040);
nand U23553 (N_23553,N_22855,N_22643);
or U23554 (N_23554,N_22280,N_22741);
and U23555 (N_23555,N_22991,N_22497);
nor U23556 (N_23556,N_22634,N_22782);
nand U23557 (N_23557,N_22717,N_22611);
xnor U23558 (N_23558,N_22583,N_22542);
nand U23559 (N_23559,N_22212,N_22258);
nand U23560 (N_23560,N_22095,N_22065);
and U23561 (N_23561,N_22683,N_22004);
nand U23562 (N_23562,N_22960,N_22617);
nand U23563 (N_23563,N_22385,N_22281);
nor U23564 (N_23564,N_22120,N_22128);
xor U23565 (N_23565,N_22535,N_22730);
nand U23566 (N_23566,N_22085,N_22718);
or U23567 (N_23567,N_22239,N_22717);
nor U23568 (N_23568,N_22997,N_22888);
nor U23569 (N_23569,N_22670,N_22227);
xnor U23570 (N_23570,N_22149,N_22877);
xor U23571 (N_23571,N_22787,N_22859);
nand U23572 (N_23572,N_22625,N_22107);
and U23573 (N_23573,N_22270,N_22282);
xnor U23574 (N_23574,N_22447,N_22370);
nor U23575 (N_23575,N_22602,N_22868);
nand U23576 (N_23576,N_22203,N_22242);
and U23577 (N_23577,N_22095,N_22081);
nor U23578 (N_23578,N_22603,N_22901);
nor U23579 (N_23579,N_22623,N_22786);
xor U23580 (N_23580,N_22073,N_22502);
nor U23581 (N_23581,N_22236,N_22060);
xnor U23582 (N_23582,N_22567,N_22431);
and U23583 (N_23583,N_22901,N_22415);
and U23584 (N_23584,N_22123,N_22509);
nor U23585 (N_23585,N_22991,N_22441);
nand U23586 (N_23586,N_22493,N_22096);
nor U23587 (N_23587,N_22099,N_22819);
nand U23588 (N_23588,N_22000,N_22864);
nand U23589 (N_23589,N_22946,N_22871);
nor U23590 (N_23590,N_22519,N_22616);
nor U23591 (N_23591,N_22638,N_22758);
nand U23592 (N_23592,N_22429,N_22971);
nor U23593 (N_23593,N_22998,N_22134);
xnor U23594 (N_23594,N_22166,N_22467);
xor U23595 (N_23595,N_22173,N_22493);
xor U23596 (N_23596,N_22894,N_22697);
or U23597 (N_23597,N_22653,N_22938);
and U23598 (N_23598,N_22478,N_22584);
nor U23599 (N_23599,N_22344,N_22247);
nor U23600 (N_23600,N_22044,N_22062);
or U23601 (N_23601,N_22917,N_22290);
and U23602 (N_23602,N_22294,N_22650);
nor U23603 (N_23603,N_22582,N_22666);
and U23604 (N_23604,N_22428,N_22382);
nand U23605 (N_23605,N_22581,N_22448);
nand U23606 (N_23606,N_22488,N_22407);
xor U23607 (N_23607,N_22488,N_22985);
nor U23608 (N_23608,N_22305,N_22203);
or U23609 (N_23609,N_22122,N_22633);
xor U23610 (N_23610,N_22702,N_22676);
nand U23611 (N_23611,N_22833,N_22598);
nor U23612 (N_23612,N_22653,N_22019);
or U23613 (N_23613,N_22386,N_22553);
or U23614 (N_23614,N_22700,N_22197);
or U23615 (N_23615,N_22518,N_22718);
or U23616 (N_23616,N_22714,N_22400);
nand U23617 (N_23617,N_22338,N_22617);
nor U23618 (N_23618,N_22615,N_22795);
and U23619 (N_23619,N_22333,N_22123);
and U23620 (N_23620,N_22584,N_22934);
nand U23621 (N_23621,N_22379,N_22373);
xnor U23622 (N_23622,N_22833,N_22954);
or U23623 (N_23623,N_22996,N_22702);
xnor U23624 (N_23624,N_22908,N_22110);
and U23625 (N_23625,N_22512,N_22959);
xnor U23626 (N_23626,N_22328,N_22909);
xor U23627 (N_23627,N_22869,N_22436);
nor U23628 (N_23628,N_22873,N_22044);
or U23629 (N_23629,N_22127,N_22646);
or U23630 (N_23630,N_22680,N_22810);
nor U23631 (N_23631,N_22288,N_22706);
or U23632 (N_23632,N_22164,N_22715);
nand U23633 (N_23633,N_22987,N_22583);
nand U23634 (N_23634,N_22963,N_22106);
xor U23635 (N_23635,N_22535,N_22376);
nand U23636 (N_23636,N_22328,N_22962);
or U23637 (N_23637,N_22645,N_22778);
or U23638 (N_23638,N_22992,N_22361);
nand U23639 (N_23639,N_22808,N_22439);
or U23640 (N_23640,N_22374,N_22412);
xnor U23641 (N_23641,N_22391,N_22037);
and U23642 (N_23642,N_22247,N_22757);
xnor U23643 (N_23643,N_22112,N_22608);
and U23644 (N_23644,N_22052,N_22299);
or U23645 (N_23645,N_22473,N_22173);
nand U23646 (N_23646,N_22113,N_22550);
and U23647 (N_23647,N_22158,N_22777);
and U23648 (N_23648,N_22859,N_22382);
or U23649 (N_23649,N_22695,N_22023);
nor U23650 (N_23650,N_22349,N_22182);
nand U23651 (N_23651,N_22617,N_22153);
or U23652 (N_23652,N_22612,N_22266);
and U23653 (N_23653,N_22321,N_22253);
nor U23654 (N_23654,N_22361,N_22339);
and U23655 (N_23655,N_22478,N_22447);
xor U23656 (N_23656,N_22606,N_22560);
or U23657 (N_23657,N_22330,N_22098);
and U23658 (N_23658,N_22153,N_22154);
or U23659 (N_23659,N_22241,N_22576);
xor U23660 (N_23660,N_22691,N_22631);
xnor U23661 (N_23661,N_22669,N_22045);
or U23662 (N_23662,N_22822,N_22572);
or U23663 (N_23663,N_22450,N_22612);
xnor U23664 (N_23664,N_22078,N_22092);
xor U23665 (N_23665,N_22352,N_22104);
xnor U23666 (N_23666,N_22125,N_22696);
nor U23667 (N_23667,N_22370,N_22177);
and U23668 (N_23668,N_22031,N_22589);
and U23669 (N_23669,N_22362,N_22134);
nor U23670 (N_23670,N_22585,N_22562);
xnor U23671 (N_23671,N_22781,N_22739);
and U23672 (N_23672,N_22017,N_22348);
xnor U23673 (N_23673,N_22847,N_22033);
and U23674 (N_23674,N_22112,N_22048);
xnor U23675 (N_23675,N_22995,N_22109);
xnor U23676 (N_23676,N_22402,N_22894);
xor U23677 (N_23677,N_22806,N_22645);
nand U23678 (N_23678,N_22401,N_22131);
xor U23679 (N_23679,N_22461,N_22661);
nand U23680 (N_23680,N_22833,N_22744);
and U23681 (N_23681,N_22297,N_22351);
nand U23682 (N_23682,N_22580,N_22460);
or U23683 (N_23683,N_22728,N_22127);
or U23684 (N_23684,N_22737,N_22210);
and U23685 (N_23685,N_22505,N_22895);
and U23686 (N_23686,N_22565,N_22878);
xor U23687 (N_23687,N_22232,N_22983);
nand U23688 (N_23688,N_22102,N_22847);
xnor U23689 (N_23689,N_22262,N_22340);
and U23690 (N_23690,N_22933,N_22733);
xnor U23691 (N_23691,N_22578,N_22623);
nand U23692 (N_23692,N_22574,N_22046);
and U23693 (N_23693,N_22389,N_22951);
nand U23694 (N_23694,N_22742,N_22019);
xor U23695 (N_23695,N_22318,N_22203);
nor U23696 (N_23696,N_22822,N_22516);
and U23697 (N_23697,N_22757,N_22903);
or U23698 (N_23698,N_22629,N_22251);
and U23699 (N_23699,N_22632,N_22545);
and U23700 (N_23700,N_22446,N_22936);
nor U23701 (N_23701,N_22624,N_22041);
nor U23702 (N_23702,N_22782,N_22683);
and U23703 (N_23703,N_22265,N_22748);
and U23704 (N_23704,N_22643,N_22261);
and U23705 (N_23705,N_22937,N_22075);
and U23706 (N_23706,N_22826,N_22709);
xor U23707 (N_23707,N_22118,N_22316);
nor U23708 (N_23708,N_22725,N_22432);
nand U23709 (N_23709,N_22583,N_22924);
nor U23710 (N_23710,N_22771,N_22653);
nor U23711 (N_23711,N_22758,N_22887);
nor U23712 (N_23712,N_22543,N_22354);
and U23713 (N_23713,N_22537,N_22194);
nand U23714 (N_23714,N_22659,N_22496);
xnor U23715 (N_23715,N_22405,N_22138);
and U23716 (N_23716,N_22244,N_22198);
nand U23717 (N_23717,N_22760,N_22699);
nand U23718 (N_23718,N_22490,N_22204);
nand U23719 (N_23719,N_22194,N_22504);
and U23720 (N_23720,N_22045,N_22303);
or U23721 (N_23721,N_22820,N_22484);
xor U23722 (N_23722,N_22540,N_22684);
or U23723 (N_23723,N_22796,N_22044);
nor U23724 (N_23724,N_22438,N_22953);
and U23725 (N_23725,N_22751,N_22802);
nor U23726 (N_23726,N_22276,N_22029);
xor U23727 (N_23727,N_22873,N_22852);
and U23728 (N_23728,N_22344,N_22070);
nand U23729 (N_23729,N_22979,N_22823);
and U23730 (N_23730,N_22209,N_22308);
nand U23731 (N_23731,N_22070,N_22924);
nor U23732 (N_23732,N_22984,N_22258);
nand U23733 (N_23733,N_22410,N_22933);
and U23734 (N_23734,N_22167,N_22348);
nor U23735 (N_23735,N_22013,N_22754);
or U23736 (N_23736,N_22617,N_22158);
nor U23737 (N_23737,N_22177,N_22864);
nor U23738 (N_23738,N_22645,N_22812);
xnor U23739 (N_23739,N_22741,N_22604);
nand U23740 (N_23740,N_22949,N_22019);
nand U23741 (N_23741,N_22616,N_22758);
nand U23742 (N_23742,N_22493,N_22327);
nor U23743 (N_23743,N_22542,N_22569);
nor U23744 (N_23744,N_22572,N_22155);
nor U23745 (N_23745,N_22183,N_22154);
and U23746 (N_23746,N_22674,N_22091);
nor U23747 (N_23747,N_22691,N_22383);
nor U23748 (N_23748,N_22464,N_22085);
xor U23749 (N_23749,N_22493,N_22484);
xor U23750 (N_23750,N_22654,N_22258);
nor U23751 (N_23751,N_22897,N_22651);
nor U23752 (N_23752,N_22338,N_22131);
nand U23753 (N_23753,N_22715,N_22779);
nand U23754 (N_23754,N_22914,N_22471);
and U23755 (N_23755,N_22022,N_22490);
and U23756 (N_23756,N_22730,N_22311);
or U23757 (N_23757,N_22512,N_22001);
nor U23758 (N_23758,N_22683,N_22064);
or U23759 (N_23759,N_22063,N_22174);
xnor U23760 (N_23760,N_22644,N_22252);
or U23761 (N_23761,N_22159,N_22424);
xor U23762 (N_23762,N_22755,N_22391);
or U23763 (N_23763,N_22956,N_22621);
xnor U23764 (N_23764,N_22270,N_22033);
nor U23765 (N_23765,N_22356,N_22475);
nor U23766 (N_23766,N_22645,N_22134);
and U23767 (N_23767,N_22405,N_22849);
or U23768 (N_23768,N_22627,N_22004);
nand U23769 (N_23769,N_22900,N_22943);
nor U23770 (N_23770,N_22949,N_22566);
nor U23771 (N_23771,N_22223,N_22529);
nand U23772 (N_23772,N_22089,N_22423);
nor U23773 (N_23773,N_22625,N_22079);
nand U23774 (N_23774,N_22694,N_22785);
and U23775 (N_23775,N_22905,N_22559);
or U23776 (N_23776,N_22350,N_22758);
xnor U23777 (N_23777,N_22474,N_22163);
xor U23778 (N_23778,N_22219,N_22987);
nand U23779 (N_23779,N_22872,N_22266);
nor U23780 (N_23780,N_22981,N_22592);
xor U23781 (N_23781,N_22542,N_22987);
nand U23782 (N_23782,N_22131,N_22729);
nor U23783 (N_23783,N_22143,N_22969);
or U23784 (N_23784,N_22285,N_22523);
xnor U23785 (N_23785,N_22055,N_22793);
nand U23786 (N_23786,N_22545,N_22836);
nand U23787 (N_23787,N_22031,N_22266);
nand U23788 (N_23788,N_22460,N_22581);
and U23789 (N_23789,N_22082,N_22372);
nor U23790 (N_23790,N_22609,N_22104);
nor U23791 (N_23791,N_22488,N_22154);
or U23792 (N_23792,N_22923,N_22676);
xnor U23793 (N_23793,N_22737,N_22361);
or U23794 (N_23794,N_22117,N_22426);
nand U23795 (N_23795,N_22691,N_22865);
xor U23796 (N_23796,N_22859,N_22145);
xnor U23797 (N_23797,N_22705,N_22985);
xnor U23798 (N_23798,N_22585,N_22985);
and U23799 (N_23799,N_22271,N_22095);
and U23800 (N_23800,N_22430,N_22474);
nor U23801 (N_23801,N_22211,N_22899);
and U23802 (N_23802,N_22313,N_22948);
nor U23803 (N_23803,N_22161,N_22107);
or U23804 (N_23804,N_22982,N_22038);
nor U23805 (N_23805,N_22266,N_22749);
or U23806 (N_23806,N_22534,N_22686);
or U23807 (N_23807,N_22246,N_22257);
or U23808 (N_23808,N_22783,N_22875);
and U23809 (N_23809,N_22243,N_22239);
or U23810 (N_23810,N_22400,N_22841);
or U23811 (N_23811,N_22248,N_22960);
or U23812 (N_23812,N_22234,N_22873);
nand U23813 (N_23813,N_22392,N_22635);
or U23814 (N_23814,N_22142,N_22022);
or U23815 (N_23815,N_22793,N_22946);
nand U23816 (N_23816,N_22071,N_22195);
or U23817 (N_23817,N_22226,N_22413);
nor U23818 (N_23818,N_22455,N_22705);
nor U23819 (N_23819,N_22587,N_22002);
and U23820 (N_23820,N_22398,N_22935);
and U23821 (N_23821,N_22141,N_22631);
nand U23822 (N_23822,N_22422,N_22518);
nand U23823 (N_23823,N_22482,N_22700);
nand U23824 (N_23824,N_22158,N_22699);
or U23825 (N_23825,N_22871,N_22134);
nand U23826 (N_23826,N_22538,N_22790);
xor U23827 (N_23827,N_22397,N_22683);
nor U23828 (N_23828,N_22719,N_22938);
or U23829 (N_23829,N_22242,N_22481);
nor U23830 (N_23830,N_22277,N_22404);
xnor U23831 (N_23831,N_22656,N_22858);
or U23832 (N_23832,N_22845,N_22196);
nand U23833 (N_23833,N_22321,N_22004);
xnor U23834 (N_23834,N_22330,N_22214);
or U23835 (N_23835,N_22431,N_22631);
and U23836 (N_23836,N_22224,N_22379);
xnor U23837 (N_23837,N_22086,N_22247);
xnor U23838 (N_23838,N_22770,N_22181);
or U23839 (N_23839,N_22840,N_22980);
nand U23840 (N_23840,N_22131,N_22756);
xor U23841 (N_23841,N_22564,N_22701);
and U23842 (N_23842,N_22109,N_22264);
xnor U23843 (N_23843,N_22335,N_22046);
or U23844 (N_23844,N_22684,N_22611);
nor U23845 (N_23845,N_22640,N_22913);
xor U23846 (N_23846,N_22093,N_22641);
or U23847 (N_23847,N_22040,N_22563);
nor U23848 (N_23848,N_22450,N_22896);
or U23849 (N_23849,N_22972,N_22936);
xnor U23850 (N_23850,N_22548,N_22674);
xnor U23851 (N_23851,N_22758,N_22850);
xor U23852 (N_23852,N_22747,N_22818);
and U23853 (N_23853,N_22554,N_22057);
xnor U23854 (N_23854,N_22984,N_22754);
nand U23855 (N_23855,N_22664,N_22578);
or U23856 (N_23856,N_22384,N_22791);
nand U23857 (N_23857,N_22638,N_22785);
nand U23858 (N_23858,N_22482,N_22260);
xnor U23859 (N_23859,N_22407,N_22914);
and U23860 (N_23860,N_22274,N_22188);
xnor U23861 (N_23861,N_22481,N_22580);
xnor U23862 (N_23862,N_22724,N_22230);
xor U23863 (N_23863,N_22766,N_22090);
nor U23864 (N_23864,N_22499,N_22715);
and U23865 (N_23865,N_22681,N_22537);
and U23866 (N_23866,N_22487,N_22488);
xnor U23867 (N_23867,N_22718,N_22908);
xor U23868 (N_23868,N_22645,N_22736);
nor U23869 (N_23869,N_22077,N_22793);
and U23870 (N_23870,N_22271,N_22622);
nand U23871 (N_23871,N_22071,N_22917);
and U23872 (N_23872,N_22746,N_22972);
nor U23873 (N_23873,N_22265,N_22836);
nor U23874 (N_23874,N_22700,N_22334);
nor U23875 (N_23875,N_22302,N_22088);
nand U23876 (N_23876,N_22704,N_22010);
or U23877 (N_23877,N_22208,N_22818);
nand U23878 (N_23878,N_22139,N_22492);
nor U23879 (N_23879,N_22159,N_22747);
nand U23880 (N_23880,N_22783,N_22739);
or U23881 (N_23881,N_22600,N_22556);
or U23882 (N_23882,N_22087,N_22280);
nand U23883 (N_23883,N_22577,N_22658);
nor U23884 (N_23884,N_22024,N_22857);
and U23885 (N_23885,N_22536,N_22165);
nand U23886 (N_23886,N_22854,N_22182);
nor U23887 (N_23887,N_22204,N_22797);
xnor U23888 (N_23888,N_22655,N_22996);
or U23889 (N_23889,N_22794,N_22080);
xnor U23890 (N_23890,N_22656,N_22678);
and U23891 (N_23891,N_22382,N_22420);
nand U23892 (N_23892,N_22507,N_22303);
and U23893 (N_23893,N_22454,N_22433);
xor U23894 (N_23894,N_22985,N_22953);
or U23895 (N_23895,N_22397,N_22803);
nand U23896 (N_23896,N_22967,N_22589);
xor U23897 (N_23897,N_22712,N_22186);
nand U23898 (N_23898,N_22102,N_22897);
nor U23899 (N_23899,N_22845,N_22460);
and U23900 (N_23900,N_22140,N_22209);
or U23901 (N_23901,N_22806,N_22844);
or U23902 (N_23902,N_22189,N_22579);
or U23903 (N_23903,N_22260,N_22021);
nand U23904 (N_23904,N_22393,N_22851);
nand U23905 (N_23905,N_22062,N_22461);
xnor U23906 (N_23906,N_22457,N_22831);
nand U23907 (N_23907,N_22373,N_22946);
nand U23908 (N_23908,N_22424,N_22735);
nand U23909 (N_23909,N_22368,N_22393);
nand U23910 (N_23910,N_22941,N_22099);
or U23911 (N_23911,N_22358,N_22997);
nor U23912 (N_23912,N_22843,N_22693);
and U23913 (N_23913,N_22031,N_22883);
nand U23914 (N_23914,N_22289,N_22201);
or U23915 (N_23915,N_22838,N_22966);
and U23916 (N_23916,N_22088,N_22969);
or U23917 (N_23917,N_22677,N_22356);
nand U23918 (N_23918,N_22374,N_22998);
or U23919 (N_23919,N_22957,N_22782);
nor U23920 (N_23920,N_22680,N_22578);
nand U23921 (N_23921,N_22835,N_22303);
and U23922 (N_23922,N_22002,N_22183);
xnor U23923 (N_23923,N_22358,N_22129);
or U23924 (N_23924,N_22630,N_22675);
nand U23925 (N_23925,N_22417,N_22671);
xor U23926 (N_23926,N_22501,N_22492);
and U23927 (N_23927,N_22691,N_22221);
nand U23928 (N_23928,N_22940,N_22154);
nor U23929 (N_23929,N_22047,N_22679);
and U23930 (N_23930,N_22322,N_22944);
and U23931 (N_23931,N_22916,N_22696);
or U23932 (N_23932,N_22453,N_22037);
or U23933 (N_23933,N_22690,N_22612);
and U23934 (N_23934,N_22455,N_22013);
nor U23935 (N_23935,N_22908,N_22713);
nor U23936 (N_23936,N_22703,N_22556);
nor U23937 (N_23937,N_22361,N_22689);
or U23938 (N_23938,N_22344,N_22369);
nor U23939 (N_23939,N_22517,N_22908);
nand U23940 (N_23940,N_22662,N_22390);
nor U23941 (N_23941,N_22966,N_22620);
nor U23942 (N_23942,N_22026,N_22378);
nand U23943 (N_23943,N_22390,N_22262);
or U23944 (N_23944,N_22362,N_22664);
and U23945 (N_23945,N_22536,N_22579);
nand U23946 (N_23946,N_22043,N_22712);
nand U23947 (N_23947,N_22041,N_22701);
nor U23948 (N_23948,N_22560,N_22800);
xor U23949 (N_23949,N_22969,N_22749);
and U23950 (N_23950,N_22925,N_22237);
or U23951 (N_23951,N_22510,N_22089);
nor U23952 (N_23952,N_22582,N_22900);
nand U23953 (N_23953,N_22408,N_22155);
xor U23954 (N_23954,N_22063,N_22855);
and U23955 (N_23955,N_22729,N_22510);
or U23956 (N_23956,N_22365,N_22163);
xor U23957 (N_23957,N_22752,N_22935);
nor U23958 (N_23958,N_22837,N_22904);
xnor U23959 (N_23959,N_22452,N_22584);
xnor U23960 (N_23960,N_22180,N_22730);
or U23961 (N_23961,N_22427,N_22839);
or U23962 (N_23962,N_22077,N_22850);
and U23963 (N_23963,N_22182,N_22083);
xor U23964 (N_23964,N_22965,N_22582);
nand U23965 (N_23965,N_22041,N_22136);
and U23966 (N_23966,N_22108,N_22830);
and U23967 (N_23967,N_22888,N_22415);
or U23968 (N_23968,N_22048,N_22633);
and U23969 (N_23969,N_22171,N_22706);
or U23970 (N_23970,N_22453,N_22367);
and U23971 (N_23971,N_22429,N_22703);
and U23972 (N_23972,N_22125,N_22839);
xnor U23973 (N_23973,N_22843,N_22842);
xnor U23974 (N_23974,N_22472,N_22210);
and U23975 (N_23975,N_22832,N_22840);
xor U23976 (N_23976,N_22743,N_22814);
and U23977 (N_23977,N_22740,N_22227);
or U23978 (N_23978,N_22490,N_22321);
or U23979 (N_23979,N_22999,N_22151);
nand U23980 (N_23980,N_22284,N_22510);
xor U23981 (N_23981,N_22701,N_22661);
nand U23982 (N_23982,N_22638,N_22705);
nor U23983 (N_23983,N_22503,N_22950);
or U23984 (N_23984,N_22555,N_22510);
or U23985 (N_23985,N_22060,N_22286);
xor U23986 (N_23986,N_22979,N_22014);
nand U23987 (N_23987,N_22196,N_22828);
nand U23988 (N_23988,N_22412,N_22564);
or U23989 (N_23989,N_22464,N_22175);
xnor U23990 (N_23990,N_22885,N_22482);
nand U23991 (N_23991,N_22257,N_22699);
nand U23992 (N_23992,N_22731,N_22180);
nand U23993 (N_23993,N_22630,N_22610);
xnor U23994 (N_23994,N_22776,N_22492);
nand U23995 (N_23995,N_22582,N_22675);
nand U23996 (N_23996,N_22620,N_22661);
nor U23997 (N_23997,N_22008,N_22487);
nand U23998 (N_23998,N_22770,N_22651);
xor U23999 (N_23999,N_22552,N_22701);
xnor U24000 (N_24000,N_23952,N_23039);
nor U24001 (N_24001,N_23909,N_23262);
or U24002 (N_24002,N_23484,N_23071);
and U24003 (N_24003,N_23654,N_23973);
or U24004 (N_24004,N_23562,N_23928);
or U24005 (N_24005,N_23549,N_23038);
xor U24006 (N_24006,N_23075,N_23347);
xor U24007 (N_24007,N_23255,N_23689);
nand U24008 (N_24008,N_23425,N_23923);
nor U24009 (N_24009,N_23503,N_23486);
nor U24010 (N_24010,N_23462,N_23559);
xor U24011 (N_24011,N_23374,N_23107);
xor U24012 (N_24012,N_23382,N_23676);
and U24013 (N_24013,N_23324,N_23800);
and U24014 (N_24014,N_23989,N_23623);
nor U24015 (N_24015,N_23550,N_23763);
or U24016 (N_24016,N_23210,N_23584);
xnor U24017 (N_24017,N_23352,N_23275);
xnor U24018 (N_24018,N_23509,N_23793);
and U24019 (N_24019,N_23116,N_23687);
nor U24020 (N_24020,N_23381,N_23703);
xor U24021 (N_24021,N_23734,N_23314);
and U24022 (N_24022,N_23596,N_23375);
nor U24023 (N_24023,N_23451,N_23536);
and U24024 (N_24024,N_23790,N_23480);
and U24025 (N_24025,N_23894,N_23294);
nand U24026 (N_24026,N_23638,N_23662);
nor U24027 (N_24027,N_23061,N_23343);
and U24028 (N_24028,N_23619,N_23735);
nand U24029 (N_24029,N_23185,N_23518);
or U24030 (N_24030,N_23749,N_23203);
nand U24031 (N_24031,N_23776,N_23620);
or U24032 (N_24032,N_23050,N_23191);
nand U24033 (N_24033,N_23753,N_23574);
nor U24034 (N_24034,N_23320,N_23283);
nand U24035 (N_24035,N_23254,N_23293);
nor U24036 (N_24036,N_23525,N_23821);
xnor U24037 (N_24037,N_23969,N_23552);
nor U24038 (N_24038,N_23477,N_23491);
and U24039 (N_24039,N_23169,N_23972);
xnor U24040 (N_24040,N_23471,N_23863);
or U24041 (N_24041,N_23630,N_23811);
or U24042 (N_24042,N_23545,N_23230);
or U24043 (N_24043,N_23267,N_23240);
xor U24044 (N_24044,N_23888,N_23505);
or U24045 (N_24045,N_23558,N_23166);
nor U24046 (N_24046,N_23031,N_23557);
xor U24047 (N_24047,N_23807,N_23367);
and U24048 (N_24048,N_23996,N_23951);
xor U24049 (N_24049,N_23015,N_23898);
and U24050 (N_24050,N_23042,N_23163);
or U24051 (N_24051,N_23111,N_23658);
or U24052 (N_24052,N_23601,N_23511);
or U24053 (N_24053,N_23692,N_23049);
nor U24054 (N_24054,N_23448,N_23987);
or U24055 (N_24055,N_23946,N_23351);
and U24056 (N_24056,N_23006,N_23300);
or U24057 (N_24057,N_23548,N_23943);
xnor U24058 (N_24058,N_23177,N_23616);
nand U24059 (N_24059,N_23740,N_23154);
or U24060 (N_24060,N_23791,N_23472);
nand U24061 (N_24061,N_23962,N_23804);
xnor U24062 (N_24062,N_23681,N_23919);
nand U24063 (N_24063,N_23520,N_23048);
nor U24064 (N_24064,N_23277,N_23865);
xor U24065 (N_24065,N_23290,N_23436);
nand U24066 (N_24066,N_23498,N_23745);
nand U24067 (N_24067,N_23473,N_23282);
xnor U24068 (N_24068,N_23529,N_23986);
nor U24069 (N_24069,N_23308,N_23705);
and U24070 (N_24070,N_23820,N_23795);
xor U24071 (N_24071,N_23074,N_23433);
nand U24072 (N_24072,N_23813,N_23312);
and U24073 (N_24073,N_23570,N_23147);
xor U24074 (N_24074,N_23418,N_23337);
nor U24075 (N_24075,N_23205,N_23591);
nand U24076 (N_24076,N_23104,N_23011);
xor U24077 (N_24077,N_23594,N_23141);
nor U24078 (N_24078,N_23396,N_23195);
xnor U24079 (N_24079,N_23652,N_23452);
nor U24080 (N_24080,N_23516,N_23773);
nor U24081 (N_24081,N_23435,N_23744);
nor U24082 (N_24082,N_23234,N_23657);
or U24083 (N_24083,N_23856,N_23767);
nor U24084 (N_24084,N_23138,N_23698);
or U24085 (N_24085,N_23463,N_23615);
nor U24086 (N_24086,N_23904,N_23880);
and U24087 (N_24087,N_23489,N_23707);
or U24088 (N_24088,N_23675,N_23515);
nor U24089 (N_24089,N_23642,N_23886);
nand U24090 (N_24090,N_23231,N_23899);
or U24091 (N_24091,N_23441,N_23128);
xnor U24092 (N_24092,N_23432,N_23572);
or U24093 (N_24093,N_23431,N_23326);
or U24094 (N_24094,N_23781,N_23988);
nor U24095 (N_24095,N_23582,N_23391);
nand U24096 (N_24096,N_23304,N_23901);
nor U24097 (N_24097,N_23787,N_23087);
nand U24098 (N_24098,N_23236,N_23702);
xor U24099 (N_24099,N_23526,N_23633);
nor U24100 (N_24100,N_23841,N_23174);
or U24101 (N_24101,N_23991,N_23933);
nor U24102 (N_24102,N_23335,N_23667);
and U24103 (N_24103,N_23510,N_23537);
or U24104 (N_24104,N_23941,N_23858);
and U24105 (N_24105,N_23051,N_23069);
xnor U24106 (N_24106,N_23656,N_23175);
and U24107 (N_24107,N_23819,N_23028);
and U24108 (N_24108,N_23045,N_23760);
nor U24109 (N_24109,N_23982,N_23672);
nand U24110 (N_24110,N_23133,N_23772);
nor U24111 (N_24111,N_23215,N_23338);
nand U24112 (N_24112,N_23523,N_23132);
or U24113 (N_24113,N_23189,N_23739);
xnor U24114 (N_24114,N_23782,N_23990);
nor U24115 (N_24115,N_23757,N_23243);
or U24116 (N_24116,N_23378,N_23409);
xnor U24117 (N_24117,N_23651,N_23030);
and U24118 (N_24118,N_23403,N_23640);
nor U24119 (N_24119,N_23578,N_23186);
nor U24120 (N_24120,N_23710,N_23871);
or U24121 (N_24121,N_23036,N_23876);
xnor U24122 (N_24122,N_23118,N_23994);
nand U24123 (N_24123,N_23096,N_23490);
or U24124 (N_24124,N_23910,N_23029);
or U24125 (N_24125,N_23634,N_23497);
nand U24126 (N_24126,N_23540,N_23291);
xnor U24127 (N_24127,N_23302,N_23386);
and U24128 (N_24128,N_23065,N_23199);
xor U24129 (N_24129,N_23274,N_23709);
or U24130 (N_24130,N_23999,N_23353);
or U24131 (N_24131,N_23602,N_23395);
or U24132 (N_24132,N_23164,N_23964);
xor U24133 (N_24133,N_23475,N_23853);
nand U24134 (N_24134,N_23697,N_23522);
xnor U24135 (N_24135,N_23421,N_23256);
and U24136 (N_24136,N_23513,N_23182);
nand U24137 (N_24137,N_23592,N_23053);
xnor U24138 (N_24138,N_23556,N_23336);
and U24139 (N_24139,N_23339,N_23464);
xnor U24140 (N_24140,N_23750,N_23514);
nor U24141 (N_24141,N_23612,N_23555);
xnor U24142 (N_24142,N_23142,N_23424);
and U24143 (N_24143,N_23001,N_23771);
and U24144 (N_24144,N_23057,N_23468);
or U24145 (N_24145,N_23945,N_23362);
xnor U24146 (N_24146,N_23092,N_23754);
and U24147 (N_24147,N_23450,N_23410);
and U24148 (N_24148,N_23541,N_23140);
and U24149 (N_24149,N_23077,N_23276);
or U24150 (N_24150,N_23350,N_23222);
or U24151 (N_24151,N_23492,N_23062);
nor U24152 (N_24152,N_23229,N_23701);
xnor U24153 (N_24153,N_23837,N_23444);
xor U24154 (N_24154,N_23249,N_23369);
nor U24155 (N_24155,N_23836,N_23816);
and U24156 (N_24156,N_23632,N_23020);
or U24157 (N_24157,N_23170,N_23825);
nand U24158 (N_24158,N_23948,N_23085);
and U24159 (N_24159,N_23748,N_23298);
or U24160 (N_24160,N_23217,N_23089);
nand U24161 (N_24161,N_23785,N_23358);
and U24162 (N_24162,N_23686,N_23938);
or U24163 (N_24163,N_23402,N_23542);
nand U24164 (N_24164,N_23332,N_23136);
xnor U24165 (N_24165,N_23830,N_23495);
nor U24166 (N_24166,N_23252,N_23932);
and U24167 (N_24167,N_23636,N_23700);
or U24168 (N_24168,N_23152,N_23090);
nand U24169 (N_24169,N_23883,N_23405);
or U24170 (N_24170,N_23034,N_23947);
or U24171 (N_24171,N_23198,N_23289);
xor U24172 (N_24172,N_23784,N_23942);
and U24173 (N_24173,N_23327,N_23388);
nand U24174 (N_24174,N_23280,N_23608);
nor U24175 (N_24175,N_23478,N_23607);
xor U24176 (N_24176,N_23007,N_23390);
or U24177 (N_24177,N_23538,N_23966);
and U24178 (N_24178,N_23233,N_23621);
nand U24179 (N_24179,N_23650,N_23512);
xor U24180 (N_24180,N_23611,N_23159);
xor U24181 (N_24181,N_23213,N_23708);
xnor U24182 (N_24182,N_23997,N_23370);
nand U24183 (N_24183,N_23653,N_23237);
xor U24184 (N_24184,N_23766,N_23023);
or U24185 (N_24185,N_23900,N_23924);
and U24186 (N_24186,N_23995,N_23397);
and U24187 (N_24187,N_23221,N_23119);
nand U24188 (N_24188,N_23927,N_23417);
nand U24189 (N_24189,N_23356,N_23931);
and U24190 (N_24190,N_23521,N_23984);
or U24191 (N_24191,N_23416,N_23377);
nor U24192 (N_24192,N_23171,N_23906);
or U24193 (N_24193,N_23714,N_23852);
nor U24194 (N_24194,N_23585,N_23588);
nand U24195 (N_24195,N_23590,N_23737);
nor U24196 (N_24196,N_23190,N_23114);
xnor U24197 (N_24197,N_23398,N_23798);
and U24198 (N_24198,N_23564,N_23976);
nand U24199 (N_24199,N_23551,N_23895);
xnor U24200 (N_24200,N_23258,N_23225);
xnor U24201 (N_24201,N_23902,N_23631);
or U24202 (N_24202,N_23004,N_23037);
nand U24203 (N_24203,N_23694,N_23861);
and U24204 (N_24204,N_23779,N_23364);
nor U24205 (N_24205,N_23010,N_23150);
nor U24206 (N_24206,N_23288,N_23840);
or U24207 (N_24207,N_23683,N_23359);
xnor U24208 (N_24208,N_23553,N_23148);
nand U24209 (N_24209,N_23859,N_23103);
nand U24210 (N_24210,N_23868,N_23789);
or U24211 (N_24211,N_23595,N_23106);
xor U24212 (N_24212,N_23257,N_23670);
nand U24213 (N_24213,N_23660,N_23829);
xor U24214 (N_24214,N_23875,N_23019);
xnor U24215 (N_24215,N_23183,N_23950);
or U24216 (N_24216,N_23794,N_23008);
nor U24217 (N_24217,N_23157,N_23822);
or U24218 (N_24218,N_23470,N_23309);
nand U24219 (N_24219,N_23907,N_23959);
or U24220 (N_24220,N_23812,N_23306);
xnor U24221 (N_24221,N_23372,N_23073);
nor U24222 (N_24222,N_23809,N_23622);
nand U24223 (N_24223,N_23122,N_23724);
nor U24224 (N_24224,N_23072,N_23671);
nor U24225 (N_24225,N_23730,N_23922);
and U24226 (N_24226,N_23896,N_23882);
nor U24227 (N_24227,N_23581,N_23586);
or U24228 (N_24228,N_23055,N_23466);
nand U24229 (N_24229,N_23801,N_23867);
nand U24230 (N_24230,N_23635,N_23979);
and U24231 (N_24231,N_23604,N_23218);
xor U24232 (N_24232,N_23488,N_23021);
and U24233 (N_24233,N_23415,N_23626);
and U24234 (N_24234,N_23135,N_23838);
and U24235 (N_24235,N_23501,N_23628);
or U24236 (N_24236,N_23404,N_23725);
xor U24237 (N_24237,N_23869,N_23862);
and U24238 (N_24238,N_23117,N_23400);
or U24239 (N_24239,N_23704,N_23691);
nand U24240 (N_24240,N_23531,N_23303);
nor U24241 (N_24241,N_23802,N_23000);
and U24242 (N_24242,N_23481,N_23956);
and U24243 (N_24243,N_23295,N_23877);
xnor U24244 (N_24244,N_23682,N_23134);
xnor U24245 (N_24245,N_23329,N_23696);
or U24246 (N_24246,N_23067,N_23736);
and U24247 (N_24247,N_23884,N_23647);
nand U24248 (N_24248,N_23720,N_23539);
nand U24249 (N_24249,N_23426,N_23831);
nor U24250 (N_24250,N_23476,N_23474);
and U24251 (N_24251,N_23914,N_23663);
or U24252 (N_24252,N_23086,N_23769);
nand U24253 (N_24253,N_23098,N_23017);
and U24254 (N_24254,N_23235,N_23674);
nor U24255 (N_24255,N_23496,N_23747);
or U24256 (N_24256,N_23155,N_23456);
nand U24257 (N_24257,N_23271,N_23685);
nor U24258 (N_24258,N_23301,N_23544);
nand U24259 (N_24259,N_23768,N_23153);
xnor U24260 (N_24260,N_23340,N_23315);
xor U24261 (N_24261,N_23115,N_23325);
and U24262 (N_24262,N_23399,N_23944);
or U24263 (N_24263,N_23746,N_23461);
or U24264 (N_24264,N_23669,N_23003);
or U24265 (N_24265,N_23597,N_23824);
nor U24266 (N_24266,N_23296,N_23219);
nor U24267 (N_24267,N_23331,N_23874);
nor U24268 (N_24268,N_23617,N_23835);
and U24269 (N_24269,N_23500,N_23130);
nor U24270 (N_24270,N_23160,N_23127);
and U24271 (N_24271,N_23251,N_23547);
or U24272 (N_24272,N_23908,N_23832);
or U24273 (N_24273,N_23527,N_23530);
and U24274 (N_24274,N_23729,N_23977);
and U24275 (N_24275,N_23953,N_23202);
or U24276 (N_24276,N_23911,N_23920);
and U24277 (N_24277,N_23376,N_23680);
and U24278 (N_24278,N_23726,N_23712);
and U24279 (N_24279,N_23070,N_23655);
and U24280 (N_24280,N_23286,N_23846);
xor U24281 (N_24281,N_23033,N_23365);
nand U24282 (N_24282,N_23892,N_23406);
xnor U24283 (N_24283,N_23806,N_23778);
nor U24284 (N_24284,N_23968,N_23125);
or U24285 (N_24285,N_23483,N_23212);
and U24286 (N_24286,N_23105,N_23643);
nand U24287 (N_24287,N_23796,N_23528);
or U24288 (N_24288,N_23571,N_23723);
nor U24289 (N_24289,N_23921,N_23613);
xor U24290 (N_24290,N_23756,N_23775);
or U24291 (N_24291,N_23245,N_23885);
nor U24292 (N_24292,N_23091,N_23046);
nor U24293 (N_24293,N_23854,N_23380);
or U24294 (N_24294,N_23196,N_23567);
nand U24295 (N_24295,N_23903,N_23279);
nand U24296 (N_24296,N_23583,N_23600);
xnor U24297 (N_24297,N_23810,N_23833);
xor U24298 (N_24298,N_23373,N_23214);
nand U24299 (N_24299,N_23009,N_23447);
nand U24300 (N_24300,N_23563,N_23847);
and U24301 (N_24301,N_23200,N_23392);
and U24302 (N_24302,N_23284,N_23459);
and U24303 (N_24303,N_23383,N_23318);
and U24304 (N_24304,N_23741,N_23316);
nand U24305 (N_24305,N_23223,N_23637);
and U24306 (N_24306,N_23285,N_23259);
or U24307 (N_24307,N_23094,N_23440);
nand U24308 (N_24308,N_23546,N_23063);
and U24309 (N_24309,N_23248,N_23269);
nand U24310 (N_24310,N_23580,N_23935);
or U24311 (N_24311,N_23129,N_23649);
and U24312 (N_24312,N_23879,N_23348);
nor U24313 (N_24313,N_23864,N_23797);
nor U24314 (N_24314,N_23679,N_23434);
or U24315 (N_24315,N_23961,N_23803);
xnor U24316 (N_24316,N_23139,N_23076);
xor U24317 (N_24317,N_23644,N_23305);
or U24318 (N_24318,N_23458,N_23207);
and U24319 (N_24319,N_23851,N_23016);
or U24320 (N_24320,N_23534,N_23176);
and U24321 (N_24321,N_23272,N_23341);
nand U24322 (N_24322,N_23241,N_23664);
nor U24323 (N_24323,N_23560,N_23764);
nor U24324 (N_24324,N_23442,N_23342);
or U24325 (N_24325,N_23079,N_23715);
nand U24326 (N_24326,N_23428,N_23731);
and U24327 (N_24327,N_23201,N_23957);
nor U24328 (N_24328,N_23661,N_23121);
xor U24329 (N_24329,N_23713,N_23026);
and U24330 (N_24330,N_23083,N_23519);
nand U24331 (N_24331,N_23101,N_23849);
nand U24332 (N_24332,N_23204,N_23208);
or U24333 (N_24333,N_23244,N_23307);
nand U24334 (N_24334,N_23706,N_23887);
nor U24335 (N_24335,N_23487,N_23445);
and U24336 (N_24336,N_23759,N_23273);
or U24337 (N_24337,N_23354,N_23743);
or U24338 (N_24338,N_23937,N_23261);
or U24339 (N_24339,N_23673,N_23823);
xor U24340 (N_24340,N_23872,N_23455);
and U24341 (N_24341,N_23845,N_23060);
or U24342 (N_24342,N_23247,N_23814);
and U24343 (N_24343,N_23504,N_23143);
and U24344 (N_24344,N_23268,N_23227);
nand U24345 (N_24345,N_23716,N_23641);
xor U24346 (N_24346,N_23024,N_23606);
or U24347 (N_24347,N_23093,N_23149);
xnor U24348 (N_24348,N_23639,N_23047);
nand U24349 (N_24349,N_23345,N_23842);
nor U24350 (N_24350,N_23913,N_23568);
and U24351 (N_24351,N_23454,N_23082);
nand U24352 (N_24352,N_23224,N_23178);
nor U24353 (N_24353,N_23081,N_23179);
and U24354 (N_24354,N_23690,N_23971);
nor U24355 (N_24355,N_23226,N_23014);
nor U24356 (N_24356,N_23394,N_23321);
or U24357 (N_24357,N_23493,N_23733);
nand U24358 (N_24358,N_23792,N_23893);
or U24359 (N_24359,N_23479,N_23099);
or U24360 (N_24360,N_23678,N_23565);
nor U24361 (N_24361,N_23366,N_23242);
nor U24362 (N_24362,N_23770,N_23438);
nand U24363 (N_24363,N_23985,N_23603);
and U24364 (N_24364,N_23981,N_23439);
nor U24365 (N_24365,N_23818,N_23870);
or U24366 (N_24366,N_23323,N_23333);
nand U24367 (N_24367,N_23629,N_23449);
and U24368 (N_24368,N_23156,N_23855);
nor U24369 (N_24369,N_23145,N_23808);
xor U24370 (N_24370,N_23843,N_23752);
nor U24371 (N_24371,N_23992,N_23317);
nand U24372 (N_24372,N_23022,N_23677);
nor U24373 (N_24373,N_23013,N_23533);
and U24374 (N_24374,N_23936,N_23209);
nor U24375 (N_24375,N_23192,N_23609);
and U24376 (N_24376,N_23384,N_23625);
nand U24377 (N_24377,N_23328,N_23446);
or U24378 (N_24378,N_23173,N_23905);
xnor U24379 (N_24379,N_23088,N_23577);
or U24380 (N_24380,N_23659,N_23827);
nor U24381 (N_24381,N_23206,N_23618);
xnor U24382 (N_24382,N_23151,N_23012);
or U24383 (N_24383,N_23299,N_23429);
xnor U24384 (N_24384,N_23355,N_23799);
or U24385 (N_24385,N_23889,N_23025);
nor U24386 (N_24386,N_23162,N_23524);
or U24387 (N_24387,N_23963,N_23181);
nor U24388 (N_24388,N_23881,N_23385);
and U24389 (N_24389,N_23357,N_23543);
nand U24390 (N_24390,N_23860,N_23379);
or U24391 (N_24391,N_23980,N_23780);
nor U24392 (N_24392,N_23124,N_23805);
or U24393 (N_24393,N_23507,N_23918);
nor U24394 (N_24394,N_23460,N_23246);
nand U24395 (N_24395,N_23742,N_23761);
nand U24396 (N_24396,N_23967,N_23535);
xor U24397 (N_24397,N_23915,N_23322);
nand U24398 (N_24398,N_23939,N_23593);
and U24399 (N_24399,N_23297,N_23457);
and U24400 (N_24400,N_23313,N_23826);
or U24401 (N_24401,N_23197,N_23068);
xor U24402 (N_24402,N_23878,N_23998);
nor U24403 (N_24403,N_23975,N_23018);
and U24404 (N_24404,N_23955,N_23232);
xor U24405 (N_24405,N_23420,N_23589);
nand U24406 (N_24406,N_23437,N_23281);
and U24407 (N_24407,N_23897,N_23755);
and U24408 (N_24408,N_23940,N_23123);
nand U24409 (N_24409,N_23187,N_23393);
or U24410 (N_24410,N_23949,N_23762);
and U24411 (N_24411,N_23738,N_23108);
and U24412 (N_24412,N_23857,N_23167);
and U24413 (N_24413,N_23408,N_23368);
nand U24414 (N_24414,N_23250,N_23110);
nor U24415 (N_24415,N_23080,N_23926);
and U24416 (N_24416,N_23239,N_23517);
nand U24417 (N_24417,N_23278,N_23684);
xnor U24418 (N_24418,N_23646,N_23165);
nor U24419 (N_24419,N_23718,N_23126);
xor U24420 (N_24420,N_23828,N_23566);
or U24421 (N_24421,N_23954,N_23993);
and U24422 (N_24422,N_23668,N_23506);
or U24423 (N_24423,N_23228,N_23413);
and U24424 (N_24424,N_23839,N_23005);
or U24425 (N_24425,N_23645,N_23777);
nor U24426 (N_24426,N_23587,N_23044);
nor U24427 (N_24427,N_23508,N_23066);
xor U24428 (N_24428,N_23978,N_23266);
nor U24429 (N_24429,N_23109,N_23168);
nand U24430 (N_24430,N_23172,N_23817);
and U24431 (N_24431,N_23220,N_23264);
nor U24432 (N_24432,N_23719,N_23158);
or U24433 (N_24433,N_23598,N_23387);
and U24434 (N_24434,N_23873,N_23054);
and U24435 (N_24435,N_23866,N_23211);
xor U24436 (N_24436,N_23443,N_23788);
nand U24437 (N_24437,N_23035,N_23319);
or U24438 (N_24438,N_23263,N_23575);
and U24439 (N_24439,N_23561,N_23002);
xor U24440 (N_24440,N_23310,N_23040);
or U24441 (N_24441,N_23965,N_23699);
xnor U24442 (N_24442,N_23064,N_23131);
nor U24443 (N_24443,N_23371,N_23688);
xnor U24444 (N_24444,N_23974,N_23848);
or U24445 (N_24445,N_23576,N_23648);
nor U24446 (N_24446,N_23502,N_23711);
nor U24447 (N_24447,N_23056,N_23722);
xnor U24448 (N_24448,N_23311,N_23027);
xor U24449 (N_24449,N_23614,N_23412);
or U24450 (N_24450,N_23260,N_23732);
nor U24451 (N_24451,N_23058,N_23180);
or U24452 (N_24452,N_23120,N_23467);
or U24453 (N_24453,N_23188,N_23624);
or U24454 (N_24454,N_23850,N_23097);
nor U24455 (N_24455,N_23579,N_23666);
nand U24456 (N_24456,N_23930,N_23569);
nand U24457 (N_24457,N_23929,N_23482);
or U24458 (N_24458,N_23721,N_23144);
nor U24459 (N_24459,N_23346,N_23960);
nor U24460 (N_24460,N_23728,N_23786);
nor U24461 (N_24461,N_23344,N_23934);
and U24462 (N_24462,N_23717,N_23727);
xor U24463 (N_24463,N_23925,N_23890);
nor U24464 (N_24464,N_23610,N_23407);
nand U24465 (N_24465,N_23958,N_23485);
xor U24466 (N_24466,N_23360,N_23161);
xor U24467 (N_24467,N_23422,N_23554);
nor U24468 (N_24468,N_23265,N_23453);
nand U24469 (N_24469,N_23084,N_23059);
xnor U24470 (N_24470,N_23627,N_23430);
nor U24471 (N_24471,N_23834,N_23253);
nand U24472 (N_24472,N_23216,N_23100);
and U24473 (N_24473,N_23917,N_23334);
and U24474 (N_24474,N_23815,N_23765);
nor U24475 (N_24475,N_23891,N_23599);
and U24476 (N_24476,N_23389,N_23783);
or U24477 (N_24477,N_23423,N_23270);
nand U24478 (N_24478,N_23043,N_23844);
nand U24479 (N_24479,N_23499,N_23494);
and U24480 (N_24480,N_23532,N_23665);
nand U24481 (N_24481,N_23363,N_23238);
or U24482 (N_24482,N_23465,N_23041);
and U24483 (N_24483,N_23695,N_23401);
nand U24484 (N_24484,N_23052,N_23427);
xor U24485 (N_24485,N_23970,N_23112);
nor U24486 (N_24486,N_23758,N_23102);
and U24487 (N_24487,N_23419,N_23146);
and U24488 (N_24488,N_23916,N_23912);
or U24489 (N_24489,N_23983,N_23194);
nand U24490 (N_24490,N_23193,N_23032);
and U24491 (N_24491,N_23469,N_23411);
nor U24492 (N_24492,N_23184,N_23573);
xor U24493 (N_24493,N_23292,N_23113);
and U24494 (N_24494,N_23774,N_23361);
nor U24495 (N_24495,N_23287,N_23751);
nor U24496 (N_24496,N_23693,N_23137);
nor U24497 (N_24497,N_23095,N_23349);
nor U24498 (N_24498,N_23414,N_23605);
and U24499 (N_24499,N_23330,N_23078);
nor U24500 (N_24500,N_23964,N_23829);
nand U24501 (N_24501,N_23338,N_23846);
and U24502 (N_24502,N_23384,N_23397);
nand U24503 (N_24503,N_23410,N_23497);
xor U24504 (N_24504,N_23467,N_23219);
nand U24505 (N_24505,N_23514,N_23337);
nor U24506 (N_24506,N_23219,N_23481);
nand U24507 (N_24507,N_23694,N_23543);
nor U24508 (N_24508,N_23205,N_23189);
and U24509 (N_24509,N_23857,N_23902);
nand U24510 (N_24510,N_23747,N_23467);
nor U24511 (N_24511,N_23663,N_23450);
and U24512 (N_24512,N_23804,N_23652);
xnor U24513 (N_24513,N_23236,N_23743);
and U24514 (N_24514,N_23228,N_23534);
nor U24515 (N_24515,N_23817,N_23717);
and U24516 (N_24516,N_23313,N_23507);
and U24517 (N_24517,N_23214,N_23220);
nor U24518 (N_24518,N_23680,N_23022);
nor U24519 (N_24519,N_23581,N_23755);
xor U24520 (N_24520,N_23865,N_23081);
nor U24521 (N_24521,N_23271,N_23896);
nor U24522 (N_24522,N_23276,N_23890);
nand U24523 (N_24523,N_23018,N_23103);
xnor U24524 (N_24524,N_23915,N_23057);
xor U24525 (N_24525,N_23615,N_23408);
xnor U24526 (N_24526,N_23675,N_23780);
nor U24527 (N_24527,N_23193,N_23412);
nor U24528 (N_24528,N_23946,N_23115);
nor U24529 (N_24529,N_23101,N_23937);
and U24530 (N_24530,N_23429,N_23316);
nor U24531 (N_24531,N_23721,N_23785);
xor U24532 (N_24532,N_23289,N_23255);
xnor U24533 (N_24533,N_23160,N_23761);
or U24534 (N_24534,N_23075,N_23858);
nor U24535 (N_24535,N_23927,N_23091);
nand U24536 (N_24536,N_23594,N_23063);
or U24537 (N_24537,N_23017,N_23549);
and U24538 (N_24538,N_23587,N_23797);
nand U24539 (N_24539,N_23735,N_23578);
xnor U24540 (N_24540,N_23868,N_23834);
and U24541 (N_24541,N_23876,N_23987);
or U24542 (N_24542,N_23407,N_23872);
or U24543 (N_24543,N_23470,N_23722);
xnor U24544 (N_24544,N_23659,N_23221);
nand U24545 (N_24545,N_23374,N_23042);
or U24546 (N_24546,N_23721,N_23371);
xor U24547 (N_24547,N_23214,N_23335);
and U24548 (N_24548,N_23566,N_23137);
and U24549 (N_24549,N_23324,N_23398);
nand U24550 (N_24550,N_23245,N_23402);
nand U24551 (N_24551,N_23084,N_23809);
and U24552 (N_24552,N_23271,N_23718);
xor U24553 (N_24553,N_23937,N_23104);
nor U24554 (N_24554,N_23677,N_23243);
or U24555 (N_24555,N_23588,N_23664);
nand U24556 (N_24556,N_23302,N_23496);
nand U24557 (N_24557,N_23488,N_23074);
nand U24558 (N_24558,N_23806,N_23047);
or U24559 (N_24559,N_23653,N_23606);
and U24560 (N_24560,N_23838,N_23853);
nor U24561 (N_24561,N_23477,N_23269);
xnor U24562 (N_24562,N_23118,N_23843);
and U24563 (N_24563,N_23872,N_23896);
xnor U24564 (N_24564,N_23118,N_23596);
nand U24565 (N_24565,N_23348,N_23150);
nor U24566 (N_24566,N_23622,N_23764);
and U24567 (N_24567,N_23012,N_23345);
nor U24568 (N_24568,N_23034,N_23368);
or U24569 (N_24569,N_23916,N_23522);
xor U24570 (N_24570,N_23224,N_23633);
xor U24571 (N_24571,N_23472,N_23559);
nand U24572 (N_24572,N_23194,N_23771);
xor U24573 (N_24573,N_23906,N_23363);
nand U24574 (N_24574,N_23029,N_23586);
nor U24575 (N_24575,N_23567,N_23460);
nor U24576 (N_24576,N_23575,N_23602);
nor U24577 (N_24577,N_23852,N_23906);
or U24578 (N_24578,N_23739,N_23812);
and U24579 (N_24579,N_23355,N_23495);
or U24580 (N_24580,N_23662,N_23392);
xor U24581 (N_24581,N_23944,N_23369);
and U24582 (N_24582,N_23068,N_23417);
or U24583 (N_24583,N_23430,N_23622);
nand U24584 (N_24584,N_23778,N_23688);
and U24585 (N_24585,N_23063,N_23670);
xor U24586 (N_24586,N_23666,N_23728);
or U24587 (N_24587,N_23522,N_23481);
xor U24588 (N_24588,N_23489,N_23164);
nor U24589 (N_24589,N_23321,N_23702);
nor U24590 (N_24590,N_23714,N_23737);
nor U24591 (N_24591,N_23816,N_23665);
or U24592 (N_24592,N_23638,N_23214);
nand U24593 (N_24593,N_23380,N_23771);
nor U24594 (N_24594,N_23079,N_23610);
nor U24595 (N_24595,N_23555,N_23984);
or U24596 (N_24596,N_23273,N_23368);
xor U24597 (N_24597,N_23711,N_23786);
and U24598 (N_24598,N_23678,N_23329);
and U24599 (N_24599,N_23612,N_23550);
or U24600 (N_24600,N_23620,N_23500);
or U24601 (N_24601,N_23053,N_23406);
or U24602 (N_24602,N_23309,N_23479);
or U24603 (N_24603,N_23856,N_23469);
and U24604 (N_24604,N_23709,N_23891);
xnor U24605 (N_24605,N_23250,N_23438);
nand U24606 (N_24606,N_23961,N_23818);
xnor U24607 (N_24607,N_23112,N_23170);
and U24608 (N_24608,N_23277,N_23987);
or U24609 (N_24609,N_23864,N_23647);
xor U24610 (N_24610,N_23026,N_23601);
xnor U24611 (N_24611,N_23044,N_23941);
or U24612 (N_24612,N_23389,N_23228);
xor U24613 (N_24613,N_23745,N_23816);
xnor U24614 (N_24614,N_23424,N_23474);
nand U24615 (N_24615,N_23650,N_23282);
nor U24616 (N_24616,N_23431,N_23168);
nand U24617 (N_24617,N_23263,N_23197);
xnor U24618 (N_24618,N_23686,N_23596);
or U24619 (N_24619,N_23393,N_23378);
nand U24620 (N_24620,N_23850,N_23846);
nand U24621 (N_24621,N_23274,N_23344);
or U24622 (N_24622,N_23021,N_23101);
nor U24623 (N_24623,N_23899,N_23691);
or U24624 (N_24624,N_23394,N_23486);
xnor U24625 (N_24625,N_23516,N_23711);
nand U24626 (N_24626,N_23487,N_23759);
nor U24627 (N_24627,N_23591,N_23179);
nand U24628 (N_24628,N_23026,N_23485);
or U24629 (N_24629,N_23916,N_23104);
nand U24630 (N_24630,N_23634,N_23674);
nor U24631 (N_24631,N_23248,N_23449);
or U24632 (N_24632,N_23644,N_23268);
nor U24633 (N_24633,N_23712,N_23233);
nand U24634 (N_24634,N_23674,N_23525);
nor U24635 (N_24635,N_23452,N_23850);
nor U24636 (N_24636,N_23909,N_23380);
xor U24637 (N_24637,N_23767,N_23227);
xnor U24638 (N_24638,N_23051,N_23952);
and U24639 (N_24639,N_23197,N_23296);
and U24640 (N_24640,N_23659,N_23153);
xnor U24641 (N_24641,N_23207,N_23975);
and U24642 (N_24642,N_23484,N_23115);
xnor U24643 (N_24643,N_23152,N_23089);
and U24644 (N_24644,N_23868,N_23505);
and U24645 (N_24645,N_23102,N_23333);
or U24646 (N_24646,N_23149,N_23195);
nor U24647 (N_24647,N_23516,N_23983);
and U24648 (N_24648,N_23600,N_23005);
and U24649 (N_24649,N_23514,N_23067);
nand U24650 (N_24650,N_23881,N_23936);
nor U24651 (N_24651,N_23827,N_23535);
and U24652 (N_24652,N_23321,N_23441);
nor U24653 (N_24653,N_23118,N_23923);
xnor U24654 (N_24654,N_23426,N_23479);
xnor U24655 (N_24655,N_23401,N_23559);
and U24656 (N_24656,N_23923,N_23022);
nand U24657 (N_24657,N_23434,N_23887);
xor U24658 (N_24658,N_23005,N_23853);
nand U24659 (N_24659,N_23048,N_23723);
and U24660 (N_24660,N_23397,N_23072);
or U24661 (N_24661,N_23385,N_23617);
and U24662 (N_24662,N_23892,N_23752);
xnor U24663 (N_24663,N_23879,N_23778);
xor U24664 (N_24664,N_23076,N_23587);
nand U24665 (N_24665,N_23095,N_23202);
or U24666 (N_24666,N_23633,N_23328);
and U24667 (N_24667,N_23470,N_23082);
xnor U24668 (N_24668,N_23658,N_23511);
xor U24669 (N_24669,N_23664,N_23962);
nand U24670 (N_24670,N_23178,N_23572);
nor U24671 (N_24671,N_23693,N_23007);
xnor U24672 (N_24672,N_23738,N_23342);
xor U24673 (N_24673,N_23605,N_23550);
nand U24674 (N_24674,N_23406,N_23142);
or U24675 (N_24675,N_23218,N_23877);
or U24676 (N_24676,N_23701,N_23561);
or U24677 (N_24677,N_23745,N_23490);
nand U24678 (N_24678,N_23868,N_23021);
and U24679 (N_24679,N_23881,N_23447);
and U24680 (N_24680,N_23283,N_23540);
or U24681 (N_24681,N_23440,N_23850);
nand U24682 (N_24682,N_23608,N_23173);
xnor U24683 (N_24683,N_23298,N_23098);
nand U24684 (N_24684,N_23433,N_23341);
xor U24685 (N_24685,N_23892,N_23946);
nor U24686 (N_24686,N_23398,N_23723);
or U24687 (N_24687,N_23047,N_23730);
xor U24688 (N_24688,N_23018,N_23243);
and U24689 (N_24689,N_23030,N_23513);
or U24690 (N_24690,N_23239,N_23792);
nor U24691 (N_24691,N_23757,N_23990);
nor U24692 (N_24692,N_23447,N_23292);
or U24693 (N_24693,N_23053,N_23631);
xor U24694 (N_24694,N_23071,N_23401);
xnor U24695 (N_24695,N_23865,N_23073);
xnor U24696 (N_24696,N_23429,N_23212);
nor U24697 (N_24697,N_23513,N_23663);
or U24698 (N_24698,N_23803,N_23584);
nand U24699 (N_24699,N_23094,N_23153);
xor U24700 (N_24700,N_23072,N_23949);
or U24701 (N_24701,N_23644,N_23190);
nand U24702 (N_24702,N_23221,N_23716);
nor U24703 (N_24703,N_23437,N_23682);
nor U24704 (N_24704,N_23374,N_23982);
and U24705 (N_24705,N_23603,N_23721);
or U24706 (N_24706,N_23210,N_23695);
or U24707 (N_24707,N_23800,N_23809);
or U24708 (N_24708,N_23973,N_23917);
nor U24709 (N_24709,N_23212,N_23249);
nor U24710 (N_24710,N_23243,N_23887);
or U24711 (N_24711,N_23438,N_23497);
nand U24712 (N_24712,N_23746,N_23789);
and U24713 (N_24713,N_23146,N_23954);
and U24714 (N_24714,N_23473,N_23358);
nor U24715 (N_24715,N_23797,N_23167);
xnor U24716 (N_24716,N_23335,N_23115);
xnor U24717 (N_24717,N_23117,N_23515);
and U24718 (N_24718,N_23371,N_23201);
or U24719 (N_24719,N_23395,N_23824);
and U24720 (N_24720,N_23021,N_23191);
xnor U24721 (N_24721,N_23963,N_23253);
nor U24722 (N_24722,N_23500,N_23290);
xor U24723 (N_24723,N_23788,N_23130);
or U24724 (N_24724,N_23065,N_23034);
xor U24725 (N_24725,N_23255,N_23608);
or U24726 (N_24726,N_23898,N_23823);
nor U24727 (N_24727,N_23759,N_23813);
or U24728 (N_24728,N_23594,N_23215);
nor U24729 (N_24729,N_23923,N_23901);
xnor U24730 (N_24730,N_23914,N_23529);
or U24731 (N_24731,N_23843,N_23225);
nand U24732 (N_24732,N_23237,N_23880);
or U24733 (N_24733,N_23102,N_23806);
or U24734 (N_24734,N_23971,N_23200);
nand U24735 (N_24735,N_23827,N_23390);
xnor U24736 (N_24736,N_23415,N_23528);
nor U24737 (N_24737,N_23369,N_23702);
and U24738 (N_24738,N_23299,N_23909);
nand U24739 (N_24739,N_23617,N_23774);
or U24740 (N_24740,N_23222,N_23518);
nor U24741 (N_24741,N_23419,N_23023);
nor U24742 (N_24742,N_23675,N_23129);
or U24743 (N_24743,N_23423,N_23132);
xnor U24744 (N_24744,N_23573,N_23010);
and U24745 (N_24745,N_23328,N_23580);
nor U24746 (N_24746,N_23218,N_23713);
nand U24747 (N_24747,N_23465,N_23567);
and U24748 (N_24748,N_23934,N_23748);
nor U24749 (N_24749,N_23399,N_23587);
nand U24750 (N_24750,N_23303,N_23336);
and U24751 (N_24751,N_23449,N_23746);
and U24752 (N_24752,N_23059,N_23238);
xnor U24753 (N_24753,N_23002,N_23803);
nor U24754 (N_24754,N_23385,N_23565);
xnor U24755 (N_24755,N_23161,N_23734);
nand U24756 (N_24756,N_23348,N_23543);
xnor U24757 (N_24757,N_23436,N_23558);
nand U24758 (N_24758,N_23826,N_23162);
xnor U24759 (N_24759,N_23859,N_23789);
xor U24760 (N_24760,N_23371,N_23650);
or U24761 (N_24761,N_23198,N_23274);
or U24762 (N_24762,N_23608,N_23213);
nand U24763 (N_24763,N_23579,N_23631);
and U24764 (N_24764,N_23969,N_23627);
and U24765 (N_24765,N_23440,N_23909);
and U24766 (N_24766,N_23484,N_23804);
nor U24767 (N_24767,N_23561,N_23774);
and U24768 (N_24768,N_23382,N_23070);
nand U24769 (N_24769,N_23276,N_23263);
and U24770 (N_24770,N_23885,N_23066);
nand U24771 (N_24771,N_23814,N_23176);
or U24772 (N_24772,N_23773,N_23843);
nand U24773 (N_24773,N_23548,N_23354);
and U24774 (N_24774,N_23724,N_23430);
nor U24775 (N_24775,N_23049,N_23519);
xor U24776 (N_24776,N_23696,N_23502);
nand U24777 (N_24777,N_23621,N_23572);
nand U24778 (N_24778,N_23481,N_23841);
nor U24779 (N_24779,N_23099,N_23379);
nor U24780 (N_24780,N_23255,N_23624);
nand U24781 (N_24781,N_23087,N_23465);
or U24782 (N_24782,N_23330,N_23382);
nor U24783 (N_24783,N_23784,N_23207);
nand U24784 (N_24784,N_23571,N_23700);
nor U24785 (N_24785,N_23661,N_23238);
nor U24786 (N_24786,N_23479,N_23534);
nor U24787 (N_24787,N_23043,N_23965);
nor U24788 (N_24788,N_23157,N_23733);
and U24789 (N_24789,N_23784,N_23022);
nand U24790 (N_24790,N_23927,N_23554);
and U24791 (N_24791,N_23282,N_23774);
nand U24792 (N_24792,N_23575,N_23153);
xnor U24793 (N_24793,N_23148,N_23563);
and U24794 (N_24794,N_23637,N_23188);
nor U24795 (N_24795,N_23654,N_23215);
nor U24796 (N_24796,N_23821,N_23533);
nor U24797 (N_24797,N_23112,N_23275);
xnor U24798 (N_24798,N_23589,N_23034);
xnor U24799 (N_24799,N_23375,N_23547);
xor U24800 (N_24800,N_23766,N_23021);
xnor U24801 (N_24801,N_23012,N_23271);
nand U24802 (N_24802,N_23135,N_23832);
nand U24803 (N_24803,N_23137,N_23871);
nand U24804 (N_24804,N_23138,N_23614);
nor U24805 (N_24805,N_23051,N_23953);
nand U24806 (N_24806,N_23389,N_23064);
and U24807 (N_24807,N_23019,N_23258);
or U24808 (N_24808,N_23010,N_23990);
nand U24809 (N_24809,N_23329,N_23009);
xnor U24810 (N_24810,N_23079,N_23073);
and U24811 (N_24811,N_23618,N_23015);
nor U24812 (N_24812,N_23874,N_23983);
nor U24813 (N_24813,N_23190,N_23068);
nand U24814 (N_24814,N_23235,N_23767);
and U24815 (N_24815,N_23609,N_23307);
nor U24816 (N_24816,N_23002,N_23765);
or U24817 (N_24817,N_23815,N_23683);
nor U24818 (N_24818,N_23749,N_23492);
and U24819 (N_24819,N_23919,N_23479);
nand U24820 (N_24820,N_23140,N_23240);
xor U24821 (N_24821,N_23279,N_23453);
nor U24822 (N_24822,N_23592,N_23465);
and U24823 (N_24823,N_23182,N_23996);
or U24824 (N_24824,N_23390,N_23473);
and U24825 (N_24825,N_23931,N_23678);
nand U24826 (N_24826,N_23101,N_23460);
nand U24827 (N_24827,N_23354,N_23442);
nand U24828 (N_24828,N_23494,N_23590);
nor U24829 (N_24829,N_23126,N_23472);
nand U24830 (N_24830,N_23479,N_23676);
or U24831 (N_24831,N_23073,N_23098);
nand U24832 (N_24832,N_23470,N_23266);
nand U24833 (N_24833,N_23892,N_23235);
and U24834 (N_24834,N_23261,N_23938);
nor U24835 (N_24835,N_23872,N_23270);
nand U24836 (N_24836,N_23074,N_23845);
and U24837 (N_24837,N_23200,N_23914);
or U24838 (N_24838,N_23305,N_23967);
or U24839 (N_24839,N_23135,N_23351);
or U24840 (N_24840,N_23728,N_23787);
nor U24841 (N_24841,N_23429,N_23954);
nor U24842 (N_24842,N_23648,N_23020);
or U24843 (N_24843,N_23823,N_23493);
nand U24844 (N_24844,N_23074,N_23965);
nor U24845 (N_24845,N_23241,N_23821);
nand U24846 (N_24846,N_23925,N_23458);
nor U24847 (N_24847,N_23898,N_23181);
or U24848 (N_24848,N_23487,N_23135);
xor U24849 (N_24849,N_23451,N_23575);
and U24850 (N_24850,N_23536,N_23214);
or U24851 (N_24851,N_23325,N_23763);
nand U24852 (N_24852,N_23858,N_23489);
and U24853 (N_24853,N_23102,N_23346);
nor U24854 (N_24854,N_23878,N_23917);
or U24855 (N_24855,N_23994,N_23249);
and U24856 (N_24856,N_23115,N_23423);
or U24857 (N_24857,N_23131,N_23336);
or U24858 (N_24858,N_23959,N_23124);
nor U24859 (N_24859,N_23757,N_23383);
nand U24860 (N_24860,N_23267,N_23998);
nand U24861 (N_24861,N_23397,N_23663);
nor U24862 (N_24862,N_23903,N_23095);
nand U24863 (N_24863,N_23864,N_23489);
nor U24864 (N_24864,N_23849,N_23311);
nand U24865 (N_24865,N_23757,N_23513);
nand U24866 (N_24866,N_23126,N_23188);
and U24867 (N_24867,N_23039,N_23131);
or U24868 (N_24868,N_23006,N_23690);
and U24869 (N_24869,N_23630,N_23626);
nor U24870 (N_24870,N_23561,N_23737);
nor U24871 (N_24871,N_23563,N_23855);
nand U24872 (N_24872,N_23324,N_23654);
xor U24873 (N_24873,N_23761,N_23888);
xor U24874 (N_24874,N_23261,N_23010);
and U24875 (N_24875,N_23048,N_23295);
nor U24876 (N_24876,N_23304,N_23224);
xnor U24877 (N_24877,N_23690,N_23261);
and U24878 (N_24878,N_23857,N_23493);
or U24879 (N_24879,N_23202,N_23638);
and U24880 (N_24880,N_23964,N_23266);
or U24881 (N_24881,N_23940,N_23767);
nor U24882 (N_24882,N_23814,N_23735);
or U24883 (N_24883,N_23052,N_23795);
xor U24884 (N_24884,N_23137,N_23339);
and U24885 (N_24885,N_23196,N_23105);
nor U24886 (N_24886,N_23712,N_23442);
nand U24887 (N_24887,N_23535,N_23035);
xor U24888 (N_24888,N_23666,N_23305);
nor U24889 (N_24889,N_23469,N_23107);
nor U24890 (N_24890,N_23821,N_23028);
xor U24891 (N_24891,N_23969,N_23916);
or U24892 (N_24892,N_23672,N_23019);
nand U24893 (N_24893,N_23929,N_23170);
xnor U24894 (N_24894,N_23902,N_23862);
nand U24895 (N_24895,N_23651,N_23560);
and U24896 (N_24896,N_23361,N_23093);
or U24897 (N_24897,N_23448,N_23251);
and U24898 (N_24898,N_23539,N_23908);
nor U24899 (N_24899,N_23204,N_23197);
nand U24900 (N_24900,N_23610,N_23508);
xnor U24901 (N_24901,N_23397,N_23045);
xnor U24902 (N_24902,N_23960,N_23503);
or U24903 (N_24903,N_23948,N_23181);
xor U24904 (N_24904,N_23002,N_23850);
xor U24905 (N_24905,N_23841,N_23364);
and U24906 (N_24906,N_23925,N_23133);
xor U24907 (N_24907,N_23562,N_23969);
or U24908 (N_24908,N_23790,N_23986);
or U24909 (N_24909,N_23613,N_23261);
nor U24910 (N_24910,N_23641,N_23358);
and U24911 (N_24911,N_23787,N_23296);
nand U24912 (N_24912,N_23198,N_23749);
nor U24913 (N_24913,N_23058,N_23170);
or U24914 (N_24914,N_23793,N_23763);
nor U24915 (N_24915,N_23236,N_23446);
xnor U24916 (N_24916,N_23754,N_23044);
xor U24917 (N_24917,N_23075,N_23712);
nand U24918 (N_24918,N_23189,N_23442);
nand U24919 (N_24919,N_23642,N_23321);
nand U24920 (N_24920,N_23524,N_23901);
xor U24921 (N_24921,N_23797,N_23364);
nand U24922 (N_24922,N_23806,N_23307);
and U24923 (N_24923,N_23983,N_23488);
nand U24924 (N_24924,N_23013,N_23261);
nand U24925 (N_24925,N_23225,N_23299);
nand U24926 (N_24926,N_23592,N_23819);
xor U24927 (N_24927,N_23827,N_23838);
nor U24928 (N_24928,N_23965,N_23830);
nand U24929 (N_24929,N_23016,N_23416);
or U24930 (N_24930,N_23245,N_23742);
and U24931 (N_24931,N_23902,N_23118);
or U24932 (N_24932,N_23377,N_23045);
or U24933 (N_24933,N_23765,N_23596);
nand U24934 (N_24934,N_23029,N_23136);
nand U24935 (N_24935,N_23186,N_23118);
and U24936 (N_24936,N_23575,N_23448);
xnor U24937 (N_24937,N_23493,N_23559);
and U24938 (N_24938,N_23813,N_23776);
and U24939 (N_24939,N_23786,N_23725);
or U24940 (N_24940,N_23976,N_23955);
and U24941 (N_24941,N_23472,N_23918);
xnor U24942 (N_24942,N_23297,N_23196);
or U24943 (N_24943,N_23865,N_23124);
or U24944 (N_24944,N_23637,N_23726);
nor U24945 (N_24945,N_23587,N_23740);
nand U24946 (N_24946,N_23963,N_23293);
or U24947 (N_24947,N_23724,N_23105);
xor U24948 (N_24948,N_23520,N_23079);
or U24949 (N_24949,N_23927,N_23889);
and U24950 (N_24950,N_23677,N_23478);
and U24951 (N_24951,N_23427,N_23639);
or U24952 (N_24952,N_23051,N_23400);
or U24953 (N_24953,N_23307,N_23728);
xnor U24954 (N_24954,N_23312,N_23279);
xor U24955 (N_24955,N_23706,N_23168);
xnor U24956 (N_24956,N_23851,N_23473);
or U24957 (N_24957,N_23825,N_23322);
or U24958 (N_24958,N_23766,N_23280);
and U24959 (N_24959,N_23641,N_23004);
nand U24960 (N_24960,N_23036,N_23030);
nor U24961 (N_24961,N_23278,N_23243);
and U24962 (N_24962,N_23601,N_23770);
nand U24963 (N_24963,N_23211,N_23048);
or U24964 (N_24964,N_23746,N_23870);
xnor U24965 (N_24965,N_23986,N_23148);
nor U24966 (N_24966,N_23136,N_23285);
and U24967 (N_24967,N_23431,N_23151);
nor U24968 (N_24968,N_23845,N_23234);
nor U24969 (N_24969,N_23919,N_23207);
or U24970 (N_24970,N_23970,N_23063);
nand U24971 (N_24971,N_23853,N_23978);
nor U24972 (N_24972,N_23252,N_23535);
xor U24973 (N_24973,N_23714,N_23564);
xnor U24974 (N_24974,N_23159,N_23772);
xor U24975 (N_24975,N_23068,N_23125);
xnor U24976 (N_24976,N_23305,N_23748);
nand U24977 (N_24977,N_23018,N_23802);
nor U24978 (N_24978,N_23361,N_23484);
xnor U24979 (N_24979,N_23600,N_23585);
or U24980 (N_24980,N_23320,N_23173);
nor U24981 (N_24981,N_23392,N_23177);
and U24982 (N_24982,N_23896,N_23410);
and U24983 (N_24983,N_23670,N_23590);
nor U24984 (N_24984,N_23984,N_23278);
xnor U24985 (N_24985,N_23957,N_23530);
xor U24986 (N_24986,N_23190,N_23895);
and U24987 (N_24987,N_23313,N_23123);
xor U24988 (N_24988,N_23370,N_23237);
and U24989 (N_24989,N_23269,N_23157);
xnor U24990 (N_24990,N_23517,N_23391);
nor U24991 (N_24991,N_23853,N_23867);
and U24992 (N_24992,N_23064,N_23459);
or U24993 (N_24993,N_23805,N_23560);
and U24994 (N_24994,N_23768,N_23879);
and U24995 (N_24995,N_23295,N_23667);
nand U24996 (N_24996,N_23537,N_23505);
nand U24997 (N_24997,N_23918,N_23977);
nor U24998 (N_24998,N_23767,N_23735);
nand U24999 (N_24999,N_23586,N_23322);
xnor U25000 (N_25000,N_24626,N_24613);
xnor U25001 (N_25001,N_24127,N_24726);
xnor U25002 (N_25002,N_24885,N_24916);
xor U25003 (N_25003,N_24826,N_24511);
nand U25004 (N_25004,N_24773,N_24807);
nand U25005 (N_25005,N_24015,N_24934);
nor U25006 (N_25006,N_24164,N_24049);
or U25007 (N_25007,N_24908,N_24258);
xor U25008 (N_25008,N_24308,N_24640);
or U25009 (N_25009,N_24556,N_24922);
xor U25010 (N_25010,N_24116,N_24946);
nand U25011 (N_25011,N_24064,N_24328);
nor U25012 (N_25012,N_24639,N_24973);
nand U25013 (N_25013,N_24827,N_24464);
or U25014 (N_25014,N_24789,N_24354);
nand U25015 (N_25015,N_24383,N_24525);
nand U25016 (N_25016,N_24332,N_24369);
and U25017 (N_25017,N_24970,N_24986);
and U25018 (N_25018,N_24954,N_24999);
nor U25019 (N_25019,N_24452,N_24251);
nor U25020 (N_25020,N_24204,N_24526);
nor U25021 (N_25021,N_24581,N_24804);
xor U25022 (N_25022,N_24947,N_24189);
nand U25023 (N_25023,N_24753,N_24521);
and U25024 (N_25024,N_24889,N_24886);
or U25025 (N_25025,N_24829,N_24077);
nor U25026 (N_25026,N_24645,N_24341);
and U25027 (N_25027,N_24048,N_24103);
xor U25028 (N_25028,N_24244,N_24429);
or U25029 (N_25029,N_24472,N_24470);
nor U25030 (N_25030,N_24536,N_24881);
nand U25031 (N_25031,N_24256,N_24478);
or U25032 (N_25032,N_24025,N_24122);
xnor U25033 (N_25033,N_24690,N_24373);
or U25034 (N_25034,N_24008,N_24051);
or U25035 (N_25035,N_24495,N_24945);
nor U25036 (N_25036,N_24683,N_24317);
or U25037 (N_25037,N_24824,N_24076);
xnor U25038 (N_25038,N_24158,N_24742);
nand U25039 (N_25039,N_24548,N_24567);
or U25040 (N_25040,N_24532,N_24877);
nand U25041 (N_25041,N_24516,N_24798);
nand U25042 (N_25042,N_24388,N_24345);
or U25043 (N_25043,N_24176,N_24738);
nor U25044 (N_25044,N_24502,N_24187);
or U25045 (N_25045,N_24871,N_24361);
and U25046 (N_25046,N_24230,N_24601);
or U25047 (N_25047,N_24146,N_24861);
nand U25048 (N_25048,N_24141,N_24591);
or U25049 (N_25049,N_24099,N_24374);
and U25050 (N_25050,N_24392,N_24352);
or U25051 (N_25051,N_24566,N_24208);
xor U25052 (N_25052,N_24370,N_24089);
nor U25053 (N_25053,N_24062,N_24961);
xnor U25054 (N_25054,N_24842,N_24437);
and U25055 (N_25055,N_24086,N_24597);
nor U25056 (N_25056,N_24702,N_24013);
or U25057 (N_25057,N_24156,N_24305);
and U25058 (N_25058,N_24896,N_24594);
nand U25059 (N_25059,N_24151,N_24041);
xnor U25060 (N_25060,N_24817,N_24764);
nor U25061 (N_25061,N_24215,N_24979);
and U25062 (N_25062,N_24682,N_24194);
nor U25063 (N_25063,N_24912,N_24781);
or U25064 (N_25064,N_24704,N_24299);
and U25065 (N_25065,N_24544,N_24273);
or U25066 (N_25066,N_24606,N_24972);
xnor U25067 (N_25067,N_24319,N_24366);
and U25068 (N_25068,N_24350,N_24130);
nand U25069 (N_25069,N_24096,N_24291);
xnor U25070 (N_25070,N_24925,N_24834);
nand U25071 (N_25071,N_24977,N_24859);
or U25072 (N_25072,N_24170,N_24811);
or U25073 (N_25073,N_24648,N_24178);
nand U25074 (N_25074,N_24175,N_24019);
or U25075 (N_25075,N_24862,N_24372);
nand U25076 (N_25076,N_24236,N_24882);
and U25077 (N_25077,N_24349,N_24381);
xnor U25078 (N_25078,N_24368,N_24783);
nor U25079 (N_25079,N_24253,N_24902);
or U25080 (N_25080,N_24277,N_24759);
xnor U25081 (N_25081,N_24568,N_24869);
xor U25082 (N_25082,N_24416,N_24237);
xnor U25083 (N_25083,N_24489,N_24184);
nand U25084 (N_25084,N_24782,N_24285);
nand U25085 (N_25085,N_24234,N_24444);
nand U25086 (N_25086,N_24557,N_24670);
and U25087 (N_25087,N_24754,N_24917);
nor U25088 (N_25088,N_24615,N_24734);
and U25089 (N_25089,N_24538,N_24728);
nand U25090 (N_25090,N_24075,N_24125);
nor U25091 (N_25091,N_24045,N_24772);
xnor U25092 (N_25092,N_24828,N_24306);
or U25093 (N_25093,N_24380,N_24745);
and U25094 (N_25094,N_24646,N_24152);
or U25095 (N_25095,N_24118,N_24643);
nor U25096 (N_25096,N_24649,N_24039);
and U25097 (N_25097,N_24985,N_24638);
or U25098 (N_25098,N_24029,N_24128);
or U25099 (N_25099,N_24873,N_24731);
or U25100 (N_25100,N_24456,N_24776);
nor U25101 (N_25101,N_24523,N_24002);
nor U25102 (N_25102,N_24609,N_24625);
or U25103 (N_25103,N_24515,N_24172);
xor U25104 (N_25104,N_24706,N_24496);
nor U25105 (N_25105,N_24522,N_24534);
and U25106 (N_25106,N_24485,N_24092);
xor U25107 (N_25107,N_24679,N_24962);
nand U25108 (N_25108,N_24936,N_24185);
and U25109 (N_25109,N_24992,N_24927);
nor U25110 (N_25110,N_24803,N_24990);
nor U25111 (N_25111,N_24790,N_24589);
or U25112 (N_25112,N_24115,N_24004);
xor U25113 (N_25113,N_24967,N_24020);
nand U25114 (N_25114,N_24499,N_24330);
and U25115 (N_25115,N_24677,N_24246);
nor U25116 (N_25116,N_24845,N_24909);
and U25117 (N_25117,N_24447,N_24364);
or U25118 (N_25118,N_24367,N_24688);
nor U25119 (N_25119,N_24242,N_24743);
nand U25120 (N_25120,N_24475,N_24147);
nand U25121 (N_25121,N_24011,N_24405);
xnor U25122 (N_25122,N_24695,N_24524);
and U25123 (N_25123,N_24428,N_24935);
xnor U25124 (N_25124,N_24174,N_24698);
nand U25125 (N_25125,N_24982,N_24576);
xor U25126 (N_25126,N_24740,N_24188);
nand U25127 (N_25127,N_24837,N_24124);
xor U25128 (N_25128,N_24056,N_24821);
xnor U25129 (N_25129,N_24852,N_24995);
nand U25130 (N_25130,N_24671,N_24540);
xor U25131 (N_25131,N_24232,N_24850);
xor U25132 (N_25132,N_24797,N_24655);
nand U25133 (N_25133,N_24211,N_24757);
or U25134 (N_25134,N_24887,N_24402);
nor U25135 (N_25135,N_24167,N_24436);
or U25136 (N_25136,N_24951,N_24697);
nor U25137 (N_25137,N_24500,N_24250);
nor U25138 (N_25138,N_24203,N_24888);
or U25139 (N_25139,N_24030,N_24966);
nand U25140 (N_25140,N_24446,N_24238);
nor U25141 (N_25141,N_24653,N_24458);
nand U25142 (N_25142,N_24055,N_24528);
nor U25143 (N_25143,N_24841,N_24315);
and U25144 (N_25144,N_24988,N_24053);
xor U25145 (N_25145,N_24413,N_24097);
nand U25146 (N_25146,N_24295,N_24200);
nor U25147 (N_25147,N_24565,N_24135);
nor U25148 (N_25148,N_24832,N_24825);
nand U25149 (N_25149,N_24036,N_24357);
or U25150 (N_25150,N_24598,N_24035);
nor U25151 (N_25151,N_24262,N_24353);
or U25152 (N_25152,N_24219,N_24260);
and U25153 (N_25153,N_24978,N_24080);
nand U25154 (N_25154,N_24586,N_24289);
and U25155 (N_25155,N_24445,N_24650);
xnor U25156 (N_25156,N_24914,N_24198);
and U25157 (N_25157,N_24145,N_24157);
or U25158 (N_25158,N_24223,N_24870);
and U25159 (N_25159,N_24968,N_24279);
and U25160 (N_25160,N_24162,N_24038);
nand U25161 (N_25161,N_24477,N_24104);
nor U25162 (N_25162,N_24297,N_24663);
or U25163 (N_25163,N_24755,N_24898);
nor U25164 (N_25164,N_24390,N_24919);
nor U25165 (N_25165,N_24513,N_24150);
nor U25166 (N_25166,N_24263,N_24471);
nor U25167 (N_25167,N_24788,N_24142);
nand U25168 (N_25168,N_24705,N_24415);
xor U25169 (N_25169,N_24137,N_24033);
and U25170 (N_25170,N_24535,N_24320);
xor U25171 (N_25171,N_24059,N_24708);
nor U25172 (N_25172,N_24133,N_24854);
nor U25173 (N_25173,N_24774,N_24490);
nor U25174 (N_25174,N_24042,N_24217);
nor U25175 (N_25175,N_24072,N_24703);
xnor U25176 (N_25176,N_24266,N_24376);
nand U25177 (N_25177,N_24681,N_24216);
or U25178 (N_25178,N_24239,N_24460);
nand U25179 (N_25179,N_24001,N_24732);
and U25180 (N_25180,N_24621,N_24220);
nand U25181 (N_25181,N_24274,N_24214);
nand U25182 (N_25182,N_24300,N_24819);
nand U25183 (N_25183,N_24699,N_24083);
and U25184 (N_25184,N_24387,N_24867);
nand U25185 (N_25185,N_24780,N_24406);
nor U25186 (N_25186,N_24541,N_24483);
and U25187 (N_25187,N_24894,N_24659);
or U25188 (N_25188,N_24459,N_24716);
or U25189 (N_25189,N_24231,N_24635);
xnor U25190 (N_25190,N_24857,N_24616);
nor U25191 (N_25191,N_24389,N_24424);
nand U25192 (N_25192,N_24915,N_24775);
nand U25193 (N_25193,N_24021,N_24675);
and U25194 (N_25194,N_24093,N_24517);
nand U25195 (N_25195,N_24180,N_24910);
nand U25196 (N_25196,N_24102,N_24044);
nand U25197 (N_25197,N_24201,N_24084);
nand U25198 (N_25198,N_24666,N_24562);
and U25199 (N_25199,N_24512,N_24469);
or U25200 (N_25200,N_24191,N_24747);
xor U25201 (N_25201,N_24131,N_24937);
nand U25202 (N_25202,N_24356,N_24667);
xor U25203 (N_25203,N_24377,N_24725);
xor U25204 (N_25204,N_24923,N_24421);
and U25205 (N_25205,N_24482,N_24132);
nand U25206 (N_25206,N_24006,N_24868);
nor U25207 (N_25207,N_24363,N_24052);
xnor U25208 (N_25208,N_24281,N_24550);
or U25209 (N_25209,N_24903,N_24644);
or U25210 (N_25210,N_24940,N_24094);
nand U25211 (N_25211,N_24139,N_24235);
nand U25212 (N_25212,N_24805,N_24358);
nand U25213 (N_25213,N_24518,N_24901);
and U25214 (N_25214,N_24778,N_24014);
nand U25215 (N_25215,N_24543,N_24040);
and U25216 (N_25216,N_24617,N_24467);
and U25217 (N_25217,N_24955,N_24920);
xnor U25218 (N_25218,N_24953,N_24272);
and U25219 (N_25219,N_24455,N_24883);
nand U25220 (N_25220,N_24864,N_24555);
xor U25221 (N_25221,N_24929,N_24282);
and U25222 (N_25222,N_24507,N_24023);
xnor U25223 (N_25223,N_24787,N_24610);
xnor U25224 (N_25224,N_24439,N_24312);
xnor U25225 (N_25225,N_24199,N_24719);
nor U25226 (N_25226,N_24549,N_24442);
or U25227 (N_25227,N_24339,N_24872);
nor U25228 (N_25228,N_24931,N_24193);
nor U25229 (N_25229,N_24971,N_24957);
xor U25230 (N_25230,N_24839,N_24993);
nand U25231 (N_25231,N_24007,N_24656);
nand U25232 (N_25232,N_24713,N_24949);
and U25233 (N_25233,N_24823,N_24100);
nor U25234 (N_25234,N_24722,N_24047);
xor U25235 (N_25235,N_24795,N_24275);
and U25236 (N_25236,N_24323,N_24637);
or U25237 (N_25237,N_24382,N_24874);
nor U25238 (N_25238,N_24183,N_24109);
xor U25239 (N_25239,N_24570,N_24451);
nand U25240 (N_25240,N_24710,N_24501);
nor U25241 (N_25241,N_24662,N_24848);
xnor U25242 (N_25242,N_24347,N_24425);
xor U25243 (N_25243,N_24433,N_24751);
xnor U25244 (N_25244,N_24321,N_24840);
nand U25245 (N_25245,N_24965,N_24816);
and U25246 (N_25246,N_24375,N_24326);
or U25247 (N_25247,N_24346,N_24689);
and U25248 (N_25248,N_24851,N_24588);
or U25249 (N_25249,N_24687,N_24561);
and U25250 (N_25250,N_24335,N_24709);
and U25251 (N_25251,N_24830,N_24652);
nand U25252 (N_25252,N_24192,N_24032);
xnor U25253 (N_25253,N_24454,N_24060);
and U25254 (N_25254,N_24197,N_24026);
nor U25255 (N_25255,N_24417,N_24660);
nor U25256 (N_25256,N_24765,N_24207);
nand U25257 (N_25257,N_24891,N_24494);
nand U25258 (N_25258,N_24784,N_24505);
nor U25259 (N_25259,N_24860,N_24975);
nor U25260 (N_25260,N_24212,N_24756);
nor U25261 (N_25261,N_24559,N_24057);
nand U25262 (N_25262,N_24546,N_24527);
nor U25263 (N_25263,N_24195,N_24835);
nand U25264 (N_25264,N_24680,N_24159);
xnor U25265 (N_25265,N_24067,N_24209);
or U25266 (N_25266,N_24969,N_24791);
xnor U25267 (N_25267,N_24712,N_24463);
nand U25268 (N_25268,N_24136,N_24717);
or U25269 (N_25269,N_24580,N_24202);
xor U25270 (N_25270,N_24658,N_24287);
or U25271 (N_25271,N_24989,N_24818);
and U25272 (N_25272,N_24426,N_24736);
nor U25273 (N_25273,N_24984,N_24331);
nand U25274 (N_25274,N_24061,N_24813);
and U25275 (N_25275,N_24431,N_24264);
and U25276 (N_25276,N_24276,N_24280);
xnor U25277 (N_25277,N_24430,N_24397);
nor U25278 (N_25278,N_24723,N_24572);
or U25279 (N_25279,N_24661,N_24620);
nor U25280 (N_25280,N_24179,N_24654);
or U25281 (N_25281,N_24700,N_24288);
or U25282 (N_25282,N_24213,N_24409);
or U25283 (N_25283,N_24342,N_24584);
nor U25284 (N_25284,N_24952,N_24027);
xor U25285 (N_25285,N_24991,N_24553);
xnor U25286 (N_25286,N_24907,N_24278);
or U25287 (N_25287,N_24696,N_24095);
xor U25288 (N_25288,N_24569,N_24892);
nor U25289 (N_25289,N_24578,N_24558);
xnor U25290 (N_25290,N_24800,N_24769);
nor U25291 (N_25291,N_24879,N_24403);
nand U25292 (N_25292,N_24066,N_24404);
xor U25293 (N_25293,N_24324,N_24880);
nand U25294 (N_25294,N_24296,N_24833);
or U25295 (N_25295,N_24693,N_24614);
nor U25296 (N_25296,N_24493,N_24504);
nand U25297 (N_25297,N_24810,N_24466);
or U25298 (N_25298,N_24632,N_24895);
and U25299 (N_25299,N_24733,N_24843);
and U25300 (N_25300,N_24893,N_24657);
xor U25301 (N_25301,N_24926,N_24865);
and U25302 (N_25302,N_24497,N_24412);
nand U25303 (N_25303,N_24301,N_24484);
xnor U25304 (N_25304,N_24334,N_24542);
nand U25305 (N_25305,N_24487,N_24016);
nor U25306 (N_25306,N_24932,N_24906);
nand U25307 (N_25307,N_24313,N_24360);
xnor U25308 (N_25308,N_24058,N_24590);
nor U25309 (N_25309,N_24206,N_24627);
or U25310 (N_25310,N_24913,N_24254);
or U25311 (N_25311,N_24017,N_24473);
and U25312 (N_25312,N_24960,N_24240);
and U25313 (N_25313,N_24794,N_24711);
xor U25314 (N_25314,N_24408,N_24351);
or U25315 (N_25315,N_24166,N_24612);
nand U25316 (N_25316,N_24010,N_24749);
and U25317 (N_25317,N_24340,N_24453);
nand U25318 (N_25318,N_24107,N_24292);
nor U25319 (N_25319,N_24079,N_24441);
xnor U25320 (N_25320,N_24123,N_24786);
and U25321 (N_25321,N_24009,N_24509);
xnor U25322 (N_25322,N_24293,N_24603);
xnor U25323 (N_25323,N_24267,N_24619);
nand U25324 (N_25324,N_24585,N_24227);
nor U25325 (N_25325,N_24629,N_24943);
or U25326 (N_25326,N_24685,N_24435);
and U25327 (N_25327,N_24846,N_24983);
and U25328 (N_25328,N_24365,N_24304);
xor U25329 (N_25329,N_24249,N_24081);
or U25330 (N_25330,N_24302,N_24149);
xor U25331 (N_25331,N_24651,N_24101);
xor U25332 (N_25332,N_24336,N_24085);
or U25333 (N_25333,N_24924,N_24046);
nor U25334 (N_25334,N_24574,N_24838);
or U25335 (N_25335,N_24420,N_24963);
or U25336 (N_25336,N_24715,N_24031);
or U25337 (N_25337,N_24457,N_24672);
nor U25338 (N_25338,N_24269,N_24318);
nand U25339 (N_25339,N_24801,N_24480);
or U25340 (N_25340,N_24537,N_24596);
or U25341 (N_25341,N_24050,N_24307);
nand U25342 (N_25342,N_24605,N_24218);
nor U25343 (N_25343,N_24153,N_24034);
nor U25344 (N_25344,N_24434,N_24043);
nand U25345 (N_25345,N_24228,N_24855);
nand U25346 (N_25346,N_24322,N_24465);
nor U25347 (N_25347,N_24673,N_24766);
nor U25348 (N_25348,N_24438,N_24996);
nand U25349 (N_25349,N_24890,N_24071);
xnor U25350 (N_25350,N_24310,N_24255);
and U25351 (N_25351,N_24763,N_24000);
nand U25352 (N_25352,N_24163,N_24796);
nor U25353 (N_25353,N_24779,N_24737);
nor U25354 (N_25354,N_24897,N_24468);
xnor U25355 (N_25355,N_24849,N_24106);
nand U25356 (N_25356,N_24386,N_24564);
nand U25357 (N_25357,N_24268,N_24866);
nand U25358 (N_25358,N_24899,N_24551);
or U25359 (N_25359,N_24165,N_24224);
xor U25360 (N_25360,N_24607,N_24694);
nand U25361 (N_25361,N_24221,N_24283);
xnor U25362 (N_25362,N_24314,N_24593);
or U25363 (N_25363,N_24822,N_24608);
xnor U25364 (N_25364,N_24563,N_24847);
and U25365 (N_25365,N_24508,N_24647);
nor U25366 (N_25366,N_24577,N_24812);
or U25367 (N_25367,N_24762,N_24210);
or U25368 (N_25368,N_24088,N_24476);
xor U25369 (N_25369,N_24126,N_24875);
or U25370 (N_25370,N_24618,N_24718);
or U25371 (N_25371,N_24091,N_24247);
xnor U25372 (N_25372,N_24583,N_24600);
xor U25373 (N_25373,N_24665,N_24474);
xnor U25374 (N_25374,N_24411,N_24245);
and U25375 (N_25375,N_24068,N_24371);
or U25376 (N_25376,N_24836,N_24750);
xor U25377 (N_25377,N_24082,N_24394);
xor U25378 (N_25378,N_24785,N_24820);
nand U25379 (N_25379,N_24063,N_24105);
nor U25380 (N_25380,N_24491,N_24410);
xor U25381 (N_25381,N_24806,N_24604);
and U25382 (N_25382,N_24950,N_24793);
or U25383 (N_25383,N_24630,N_24155);
or U25384 (N_25384,N_24707,N_24552);
or U25385 (N_25385,N_24018,N_24190);
nor U25386 (N_25386,N_24391,N_24933);
xor U25387 (N_25387,N_24037,N_24503);
xnor U25388 (N_25388,N_24090,N_24396);
and U25389 (N_25389,N_24461,N_24575);
nor U25390 (N_25390,N_24120,N_24259);
nor U25391 (N_25391,N_24746,N_24595);
nor U25392 (N_25392,N_24355,N_24941);
or U25393 (N_25393,N_24257,N_24222);
nor U25394 (N_25394,N_24814,N_24530);
xor U25395 (N_25395,N_24065,N_24173);
nand U25396 (N_25396,N_24691,N_24098);
and U25397 (N_25397,N_24311,N_24233);
or U25398 (N_25398,N_24271,N_24900);
nor U25399 (N_25399,N_24752,N_24448);
and U25400 (N_25400,N_24529,N_24486);
or U25401 (N_25401,N_24186,N_24270);
and U25402 (N_25402,N_24114,N_24348);
xnor U25403 (N_25403,N_24395,N_24768);
nand U25404 (N_25404,N_24144,N_24930);
xnor U25405 (N_25405,N_24261,N_24545);
nor U25406 (N_25406,N_24110,N_24714);
nand U25407 (N_25407,N_24054,N_24964);
nor U25408 (N_25408,N_24161,N_24831);
nand U25409 (N_25409,N_24692,N_24730);
nor U25410 (N_25410,N_24168,N_24171);
nand U25411 (N_25411,N_24294,N_24419);
nand U25412 (N_25412,N_24815,N_24359);
and U25413 (N_25413,N_24520,N_24265);
nor U25414 (N_25414,N_24676,N_24181);
nand U25415 (N_25415,N_24987,N_24863);
nand U25416 (N_25416,N_24622,N_24325);
xnor U25417 (N_25417,N_24884,N_24414);
xor U25418 (N_25418,N_24309,N_24005);
xor U25419 (N_25419,N_24422,N_24286);
or U25420 (N_25420,N_24587,N_24108);
nand U25421 (N_25421,N_24393,N_24143);
nand U25422 (N_25422,N_24160,N_24298);
and U25423 (N_25423,N_24229,N_24809);
nor U25424 (N_25424,N_24028,N_24720);
nand U25425 (N_25425,N_24560,N_24138);
and U25426 (N_25426,N_24876,N_24440);
or U25427 (N_25427,N_24479,N_24069);
or U25428 (N_25428,N_24904,N_24290);
nand U25429 (N_25429,N_24078,N_24344);
and U25430 (N_25430,N_24498,N_24533);
and U25431 (N_25431,N_24674,N_24087);
and U25432 (N_25432,N_24449,N_24959);
or U25433 (N_25433,N_24856,N_24928);
or U25434 (N_25434,N_24802,N_24631);
or U25435 (N_25435,N_24327,N_24140);
nor U25436 (N_25436,N_24177,N_24024);
or U25437 (N_25437,N_24853,N_24664);
and U25438 (N_25438,N_24129,N_24938);
nand U25439 (N_25439,N_24771,N_24303);
or U25440 (N_25440,N_24554,N_24400);
and U25441 (N_25441,N_24997,N_24686);
xor U25442 (N_25442,N_24378,N_24974);
nand U25443 (N_25443,N_24182,N_24510);
nor U25444 (N_25444,N_24748,N_24329);
or U25445 (N_25445,N_24226,N_24134);
nand U25446 (N_25446,N_24111,N_24844);
xor U25447 (N_25447,N_24248,N_24423);
xnor U25448 (N_25448,N_24582,N_24642);
nand U25449 (N_25449,N_24744,N_24942);
nand U25450 (N_25450,N_24994,N_24980);
xnor U25451 (N_25451,N_24944,N_24878);
or U25452 (N_25452,N_24760,N_24724);
or U25453 (N_25453,N_24003,N_24792);
and U25454 (N_25454,N_24611,N_24316);
and U25455 (N_25455,N_24998,N_24721);
nand U25456 (N_25456,N_24729,N_24514);
nor U25457 (N_25457,N_24571,N_24905);
or U25458 (N_25458,N_24385,N_24112);
and U25459 (N_25459,N_24252,N_24338);
nor U25460 (N_25460,N_24624,N_24243);
or U25461 (N_25461,N_24636,N_24384);
or U25462 (N_25462,N_24948,N_24633);
nand U25463 (N_25463,N_24573,N_24432);
xor U25464 (N_25464,N_24956,N_24154);
xor U25465 (N_25465,N_24592,N_24958);
nand U25466 (N_25466,N_24727,N_24858);
nand U25467 (N_25467,N_24808,N_24599);
xnor U25468 (N_25468,N_24735,N_24799);
or U25469 (N_25469,N_24399,N_24379);
nand U25470 (N_25470,N_24741,N_24333);
and U25471 (N_25471,N_24488,N_24121);
and U25472 (N_25472,N_24921,N_24668);
or U25473 (N_25473,N_24450,N_24918);
nor U25474 (N_25474,N_24401,N_24241);
nand U25475 (N_25475,N_24547,N_24169);
or U25476 (N_25476,N_24225,N_24074);
xor U25477 (N_25477,N_24531,N_24669);
nand U25478 (N_25478,N_24022,N_24602);
and U25479 (N_25479,N_24739,N_24070);
nand U25480 (N_25480,N_24427,N_24196);
and U25481 (N_25481,N_24579,N_24506);
nand U25482 (N_25482,N_24462,N_24701);
nand U25483 (N_25483,N_24343,N_24641);
and U25484 (N_25484,N_24981,N_24119);
xnor U25485 (N_25485,N_24634,N_24777);
nor U25486 (N_25486,N_24761,N_24117);
or U25487 (N_25487,N_24205,N_24623);
and U25488 (N_25488,N_24418,N_24443);
nand U25489 (N_25489,N_24519,N_24284);
xor U25490 (N_25490,N_24481,N_24148);
nor U25491 (N_25491,N_24398,N_24758);
or U25492 (N_25492,N_24073,N_24678);
nand U25493 (N_25493,N_24628,N_24911);
and U25494 (N_25494,N_24767,N_24976);
xnor U25495 (N_25495,N_24407,N_24684);
and U25496 (N_25496,N_24113,N_24492);
nand U25497 (N_25497,N_24939,N_24362);
xor U25498 (N_25498,N_24337,N_24012);
and U25499 (N_25499,N_24539,N_24770);
xor U25500 (N_25500,N_24316,N_24743);
nor U25501 (N_25501,N_24875,N_24085);
or U25502 (N_25502,N_24457,N_24731);
nand U25503 (N_25503,N_24837,N_24802);
nor U25504 (N_25504,N_24862,N_24380);
nand U25505 (N_25505,N_24978,N_24481);
or U25506 (N_25506,N_24084,N_24108);
and U25507 (N_25507,N_24461,N_24972);
xor U25508 (N_25508,N_24616,N_24289);
nor U25509 (N_25509,N_24473,N_24369);
nand U25510 (N_25510,N_24269,N_24311);
xnor U25511 (N_25511,N_24971,N_24367);
nand U25512 (N_25512,N_24350,N_24750);
nor U25513 (N_25513,N_24119,N_24989);
nand U25514 (N_25514,N_24815,N_24076);
and U25515 (N_25515,N_24168,N_24435);
xnor U25516 (N_25516,N_24236,N_24791);
nor U25517 (N_25517,N_24263,N_24833);
or U25518 (N_25518,N_24924,N_24739);
xnor U25519 (N_25519,N_24588,N_24089);
and U25520 (N_25520,N_24764,N_24246);
or U25521 (N_25521,N_24990,N_24519);
or U25522 (N_25522,N_24124,N_24033);
nor U25523 (N_25523,N_24159,N_24477);
and U25524 (N_25524,N_24503,N_24412);
or U25525 (N_25525,N_24616,N_24992);
nor U25526 (N_25526,N_24980,N_24706);
nand U25527 (N_25527,N_24023,N_24651);
or U25528 (N_25528,N_24317,N_24971);
and U25529 (N_25529,N_24349,N_24919);
xnor U25530 (N_25530,N_24378,N_24116);
nand U25531 (N_25531,N_24527,N_24946);
nand U25532 (N_25532,N_24722,N_24328);
nand U25533 (N_25533,N_24127,N_24142);
or U25534 (N_25534,N_24072,N_24510);
or U25535 (N_25535,N_24296,N_24232);
or U25536 (N_25536,N_24086,N_24071);
or U25537 (N_25537,N_24393,N_24608);
or U25538 (N_25538,N_24325,N_24609);
nand U25539 (N_25539,N_24392,N_24534);
xor U25540 (N_25540,N_24020,N_24330);
nor U25541 (N_25541,N_24713,N_24749);
or U25542 (N_25542,N_24257,N_24986);
or U25543 (N_25543,N_24552,N_24087);
and U25544 (N_25544,N_24145,N_24794);
nor U25545 (N_25545,N_24228,N_24146);
or U25546 (N_25546,N_24408,N_24221);
xor U25547 (N_25547,N_24048,N_24864);
xnor U25548 (N_25548,N_24041,N_24999);
or U25549 (N_25549,N_24388,N_24487);
and U25550 (N_25550,N_24100,N_24828);
nand U25551 (N_25551,N_24248,N_24615);
nand U25552 (N_25552,N_24479,N_24844);
nand U25553 (N_25553,N_24208,N_24712);
or U25554 (N_25554,N_24380,N_24051);
xor U25555 (N_25555,N_24003,N_24854);
xor U25556 (N_25556,N_24827,N_24076);
nand U25557 (N_25557,N_24363,N_24981);
and U25558 (N_25558,N_24049,N_24574);
xor U25559 (N_25559,N_24297,N_24379);
xnor U25560 (N_25560,N_24993,N_24960);
or U25561 (N_25561,N_24370,N_24834);
nand U25562 (N_25562,N_24666,N_24259);
nor U25563 (N_25563,N_24589,N_24503);
nor U25564 (N_25564,N_24059,N_24776);
nor U25565 (N_25565,N_24144,N_24950);
and U25566 (N_25566,N_24552,N_24916);
nor U25567 (N_25567,N_24736,N_24860);
and U25568 (N_25568,N_24817,N_24105);
and U25569 (N_25569,N_24289,N_24563);
and U25570 (N_25570,N_24828,N_24708);
or U25571 (N_25571,N_24870,N_24368);
and U25572 (N_25572,N_24215,N_24185);
and U25573 (N_25573,N_24064,N_24432);
nand U25574 (N_25574,N_24864,N_24521);
xor U25575 (N_25575,N_24072,N_24131);
or U25576 (N_25576,N_24570,N_24162);
nor U25577 (N_25577,N_24919,N_24810);
nand U25578 (N_25578,N_24342,N_24590);
xor U25579 (N_25579,N_24446,N_24687);
nand U25580 (N_25580,N_24601,N_24528);
and U25581 (N_25581,N_24135,N_24727);
and U25582 (N_25582,N_24486,N_24891);
xnor U25583 (N_25583,N_24567,N_24794);
and U25584 (N_25584,N_24598,N_24419);
nor U25585 (N_25585,N_24589,N_24633);
and U25586 (N_25586,N_24318,N_24367);
xnor U25587 (N_25587,N_24324,N_24635);
or U25588 (N_25588,N_24919,N_24259);
or U25589 (N_25589,N_24502,N_24021);
nor U25590 (N_25590,N_24554,N_24500);
or U25591 (N_25591,N_24510,N_24068);
or U25592 (N_25592,N_24233,N_24256);
nor U25593 (N_25593,N_24658,N_24274);
xor U25594 (N_25594,N_24817,N_24074);
nor U25595 (N_25595,N_24878,N_24979);
xnor U25596 (N_25596,N_24728,N_24714);
nand U25597 (N_25597,N_24899,N_24546);
nor U25598 (N_25598,N_24189,N_24359);
nor U25599 (N_25599,N_24228,N_24825);
xor U25600 (N_25600,N_24129,N_24318);
xor U25601 (N_25601,N_24623,N_24621);
nor U25602 (N_25602,N_24226,N_24155);
nor U25603 (N_25603,N_24336,N_24981);
nand U25604 (N_25604,N_24672,N_24981);
nand U25605 (N_25605,N_24393,N_24737);
or U25606 (N_25606,N_24803,N_24507);
nor U25607 (N_25607,N_24512,N_24268);
xor U25608 (N_25608,N_24324,N_24101);
nand U25609 (N_25609,N_24645,N_24614);
xor U25610 (N_25610,N_24020,N_24271);
xor U25611 (N_25611,N_24369,N_24786);
xnor U25612 (N_25612,N_24731,N_24390);
xnor U25613 (N_25613,N_24455,N_24182);
and U25614 (N_25614,N_24481,N_24222);
nor U25615 (N_25615,N_24289,N_24363);
and U25616 (N_25616,N_24700,N_24350);
xnor U25617 (N_25617,N_24999,N_24517);
and U25618 (N_25618,N_24163,N_24756);
or U25619 (N_25619,N_24431,N_24666);
nor U25620 (N_25620,N_24312,N_24761);
nand U25621 (N_25621,N_24593,N_24275);
xor U25622 (N_25622,N_24260,N_24096);
and U25623 (N_25623,N_24247,N_24732);
xnor U25624 (N_25624,N_24566,N_24588);
nor U25625 (N_25625,N_24858,N_24893);
nand U25626 (N_25626,N_24873,N_24889);
xor U25627 (N_25627,N_24515,N_24595);
and U25628 (N_25628,N_24907,N_24043);
nand U25629 (N_25629,N_24020,N_24403);
or U25630 (N_25630,N_24888,N_24220);
and U25631 (N_25631,N_24239,N_24079);
nand U25632 (N_25632,N_24135,N_24961);
nand U25633 (N_25633,N_24832,N_24065);
nor U25634 (N_25634,N_24766,N_24044);
nand U25635 (N_25635,N_24074,N_24687);
nor U25636 (N_25636,N_24709,N_24216);
nor U25637 (N_25637,N_24720,N_24510);
nor U25638 (N_25638,N_24956,N_24874);
nand U25639 (N_25639,N_24124,N_24376);
xnor U25640 (N_25640,N_24549,N_24302);
xnor U25641 (N_25641,N_24398,N_24266);
and U25642 (N_25642,N_24249,N_24284);
and U25643 (N_25643,N_24484,N_24508);
nand U25644 (N_25644,N_24954,N_24903);
nor U25645 (N_25645,N_24365,N_24757);
nor U25646 (N_25646,N_24179,N_24450);
xnor U25647 (N_25647,N_24477,N_24185);
or U25648 (N_25648,N_24055,N_24174);
nor U25649 (N_25649,N_24578,N_24168);
or U25650 (N_25650,N_24316,N_24575);
nor U25651 (N_25651,N_24969,N_24970);
xnor U25652 (N_25652,N_24614,N_24375);
and U25653 (N_25653,N_24413,N_24354);
nor U25654 (N_25654,N_24893,N_24484);
nand U25655 (N_25655,N_24867,N_24002);
and U25656 (N_25656,N_24795,N_24023);
or U25657 (N_25657,N_24516,N_24643);
xor U25658 (N_25658,N_24978,N_24093);
nand U25659 (N_25659,N_24098,N_24925);
nand U25660 (N_25660,N_24210,N_24370);
nor U25661 (N_25661,N_24814,N_24915);
and U25662 (N_25662,N_24221,N_24603);
xnor U25663 (N_25663,N_24557,N_24481);
or U25664 (N_25664,N_24345,N_24682);
and U25665 (N_25665,N_24716,N_24129);
nor U25666 (N_25666,N_24788,N_24610);
nor U25667 (N_25667,N_24034,N_24400);
nor U25668 (N_25668,N_24881,N_24415);
nand U25669 (N_25669,N_24479,N_24024);
nor U25670 (N_25670,N_24222,N_24948);
nand U25671 (N_25671,N_24593,N_24400);
xor U25672 (N_25672,N_24680,N_24876);
and U25673 (N_25673,N_24349,N_24154);
xnor U25674 (N_25674,N_24029,N_24075);
or U25675 (N_25675,N_24038,N_24558);
or U25676 (N_25676,N_24717,N_24116);
nor U25677 (N_25677,N_24569,N_24010);
or U25678 (N_25678,N_24980,N_24549);
nand U25679 (N_25679,N_24502,N_24766);
or U25680 (N_25680,N_24605,N_24244);
or U25681 (N_25681,N_24815,N_24910);
and U25682 (N_25682,N_24208,N_24013);
nor U25683 (N_25683,N_24433,N_24130);
and U25684 (N_25684,N_24423,N_24722);
and U25685 (N_25685,N_24051,N_24498);
xnor U25686 (N_25686,N_24276,N_24095);
and U25687 (N_25687,N_24441,N_24479);
or U25688 (N_25688,N_24825,N_24868);
or U25689 (N_25689,N_24604,N_24935);
nor U25690 (N_25690,N_24160,N_24266);
nor U25691 (N_25691,N_24953,N_24300);
nand U25692 (N_25692,N_24310,N_24894);
or U25693 (N_25693,N_24863,N_24318);
or U25694 (N_25694,N_24065,N_24726);
nor U25695 (N_25695,N_24158,N_24586);
or U25696 (N_25696,N_24615,N_24744);
nor U25697 (N_25697,N_24834,N_24714);
and U25698 (N_25698,N_24727,N_24910);
nand U25699 (N_25699,N_24583,N_24781);
or U25700 (N_25700,N_24801,N_24343);
nand U25701 (N_25701,N_24223,N_24431);
xnor U25702 (N_25702,N_24528,N_24199);
xor U25703 (N_25703,N_24066,N_24910);
nand U25704 (N_25704,N_24203,N_24270);
nor U25705 (N_25705,N_24524,N_24907);
nand U25706 (N_25706,N_24448,N_24604);
nand U25707 (N_25707,N_24337,N_24827);
or U25708 (N_25708,N_24673,N_24972);
or U25709 (N_25709,N_24529,N_24880);
or U25710 (N_25710,N_24425,N_24740);
and U25711 (N_25711,N_24461,N_24513);
xnor U25712 (N_25712,N_24892,N_24368);
nor U25713 (N_25713,N_24927,N_24538);
xnor U25714 (N_25714,N_24172,N_24737);
nand U25715 (N_25715,N_24632,N_24433);
nor U25716 (N_25716,N_24741,N_24296);
or U25717 (N_25717,N_24973,N_24195);
or U25718 (N_25718,N_24109,N_24731);
nor U25719 (N_25719,N_24507,N_24581);
and U25720 (N_25720,N_24629,N_24296);
or U25721 (N_25721,N_24821,N_24265);
nor U25722 (N_25722,N_24957,N_24270);
xor U25723 (N_25723,N_24173,N_24813);
xnor U25724 (N_25724,N_24108,N_24295);
xor U25725 (N_25725,N_24096,N_24565);
or U25726 (N_25726,N_24626,N_24761);
and U25727 (N_25727,N_24168,N_24025);
or U25728 (N_25728,N_24357,N_24608);
and U25729 (N_25729,N_24830,N_24159);
xor U25730 (N_25730,N_24028,N_24102);
or U25731 (N_25731,N_24638,N_24780);
nand U25732 (N_25732,N_24021,N_24738);
xnor U25733 (N_25733,N_24164,N_24619);
or U25734 (N_25734,N_24441,N_24618);
or U25735 (N_25735,N_24936,N_24087);
or U25736 (N_25736,N_24552,N_24743);
or U25737 (N_25737,N_24455,N_24910);
or U25738 (N_25738,N_24777,N_24544);
or U25739 (N_25739,N_24583,N_24713);
nor U25740 (N_25740,N_24443,N_24310);
nor U25741 (N_25741,N_24200,N_24375);
or U25742 (N_25742,N_24092,N_24706);
and U25743 (N_25743,N_24906,N_24558);
xor U25744 (N_25744,N_24868,N_24300);
or U25745 (N_25745,N_24184,N_24947);
nand U25746 (N_25746,N_24314,N_24037);
and U25747 (N_25747,N_24935,N_24109);
nand U25748 (N_25748,N_24185,N_24254);
or U25749 (N_25749,N_24829,N_24657);
xnor U25750 (N_25750,N_24704,N_24020);
or U25751 (N_25751,N_24764,N_24714);
or U25752 (N_25752,N_24846,N_24017);
xnor U25753 (N_25753,N_24060,N_24703);
xor U25754 (N_25754,N_24248,N_24874);
or U25755 (N_25755,N_24329,N_24500);
nor U25756 (N_25756,N_24642,N_24041);
or U25757 (N_25757,N_24903,N_24684);
nand U25758 (N_25758,N_24951,N_24201);
or U25759 (N_25759,N_24031,N_24174);
nor U25760 (N_25760,N_24553,N_24095);
xor U25761 (N_25761,N_24669,N_24732);
or U25762 (N_25762,N_24810,N_24507);
xor U25763 (N_25763,N_24599,N_24368);
nand U25764 (N_25764,N_24560,N_24858);
nand U25765 (N_25765,N_24203,N_24478);
and U25766 (N_25766,N_24896,N_24049);
nor U25767 (N_25767,N_24383,N_24796);
and U25768 (N_25768,N_24538,N_24887);
xnor U25769 (N_25769,N_24893,N_24975);
or U25770 (N_25770,N_24198,N_24969);
nor U25771 (N_25771,N_24284,N_24388);
nor U25772 (N_25772,N_24478,N_24570);
and U25773 (N_25773,N_24608,N_24931);
or U25774 (N_25774,N_24417,N_24706);
nand U25775 (N_25775,N_24272,N_24273);
or U25776 (N_25776,N_24268,N_24655);
or U25777 (N_25777,N_24971,N_24587);
nor U25778 (N_25778,N_24578,N_24624);
nand U25779 (N_25779,N_24461,N_24609);
nor U25780 (N_25780,N_24548,N_24069);
xnor U25781 (N_25781,N_24705,N_24224);
or U25782 (N_25782,N_24793,N_24445);
or U25783 (N_25783,N_24249,N_24220);
nor U25784 (N_25784,N_24827,N_24971);
nand U25785 (N_25785,N_24144,N_24370);
nor U25786 (N_25786,N_24629,N_24377);
or U25787 (N_25787,N_24351,N_24125);
nand U25788 (N_25788,N_24936,N_24843);
and U25789 (N_25789,N_24296,N_24160);
or U25790 (N_25790,N_24232,N_24954);
nand U25791 (N_25791,N_24347,N_24814);
nor U25792 (N_25792,N_24952,N_24360);
xor U25793 (N_25793,N_24758,N_24771);
nand U25794 (N_25794,N_24188,N_24364);
or U25795 (N_25795,N_24502,N_24780);
or U25796 (N_25796,N_24023,N_24726);
nand U25797 (N_25797,N_24246,N_24215);
nor U25798 (N_25798,N_24455,N_24459);
and U25799 (N_25799,N_24774,N_24426);
xnor U25800 (N_25800,N_24424,N_24915);
xor U25801 (N_25801,N_24659,N_24568);
nor U25802 (N_25802,N_24688,N_24499);
nor U25803 (N_25803,N_24618,N_24975);
nor U25804 (N_25804,N_24401,N_24582);
or U25805 (N_25805,N_24214,N_24778);
nor U25806 (N_25806,N_24790,N_24884);
nand U25807 (N_25807,N_24675,N_24567);
nand U25808 (N_25808,N_24622,N_24701);
or U25809 (N_25809,N_24537,N_24065);
and U25810 (N_25810,N_24240,N_24926);
nor U25811 (N_25811,N_24150,N_24422);
nor U25812 (N_25812,N_24464,N_24506);
nand U25813 (N_25813,N_24896,N_24841);
nor U25814 (N_25814,N_24493,N_24582);
nand U25815 (N_25815,N_24916,N_24017);
or U25816 (N_25816,N_24108,N_24323);
or U25817 (N_25817,N_24048,N_24881);
or U25818 (N_25818,N_24396,N_24410);
nor U25819 (N_25819,N_24641,N_24446);
or U25820 (N_25820,N_24966,N_24557);
or U25821 (N_25821,N_24743,N_24831);
nor U25822 (N_25822,N_24445,N_24752);
xnor U25823 (N_25823,N_24934,N_24699);
xnor U25824 (N_25824,N_24472,N_24904);
nand U25825 (N_25825,N_24698,N_24761);
nand U25826 (N_25826,N_24456,N_24468);
and U25827 (N_25827,N_24890,N_24443);
nand U25828 (N_25828,N_24896,N_24345);
or U25829 (N_25829,N_24158,N_24041);
and U25830 (N_25830,N_24077,N_24801);
nor U25831 (N_25831,N_24712,N_24402);
nor U25832 (N_25832,N_24373,N_24483);
nand U25833 (N_25833,N_24660,N_24745);
nand U25834 (N_25834,N_24284,N_24320);
and U25835 (N_25835,N_24202,N_24651);
xor U25836 (N_25836,N_24757,N_24128);
xnor U25837 (N_25837,N_24286,N_24239);
xnor U25838 (N_25838,N_24293,N_24939);
and U25839 (N_25839,N_24991,N_24116);
or U25840 (N_25840,N_24561,N_24580);
and U25841 (N_25841,N_24204,N_24853);
and U25842 (N_25842,N_24957,N_24902);
nor U25843 (N_25843,N_24239,N_24266);
nor U25844 (N_25844,N_24672,N_24191);
nand U25845 (N_25845,N_24460,N_24491);
or U25846 (N_25846,N_24041,N_24630);
and U25847 (N_25847,N_24801,N_24187);
and U25848 (N_25848,N_24093,N_24323);
or U25849 (N_25849,N_24672,N_24554);
and U25850 (N_25850,N_24041,N_24496);
nor U25851 (N_25851,N_24380,N_24085);
nand U25852 (N_25852,N_24754,N_24633);
nor U25853 (N_25853,N_24060,N_24447);
xor U25854 (N_25854,N_24192,N_24095);
or U25855 (N_25855,N_24306,N_24639);
xnor U25856 (N_25856,N_24164,N_24304);
nor U25857 (N_25857,N_24299,N_24890);
or U25858 (N_25858,N_24903,N_24346);
nor U25859 (N_25859,N_24090,N_24156);
nor U25860 (N_25860,N_24455,N_24418);
xor U25861 (N_25861,N_24873,N_24297);
nand U25862 (N_25862,N_24855,N_24281);
xnor U25863 (N_25863,N_24041,N_24649);
or U25864 (N_25864,N_24407,N_24076);
or U25865 (N_25865,N_24175,N_24526);
nand U25866 (N_25866,N_24853,N_24458);
nand U25867 (N_25867,N_24749,N_24970);
or U25868 (N_25868,N_24882,N_24837);
and U25869 (N_25869,N_24003,N_24564);
xnor U25870 (N_25870,N_24657,N_24899);
xnor U25871 (N_25871,N_24893,N_24510);
and U25872 (N_25872,N_24809,N_24941);
xnor U25873 (N_25873,N_24608,N_24070);
xnor U25874 (N_25874,N_24799,N_24928);
xnor U25875 (N_25875,N_24884,N_24419);
xnor U25876 (N_25876,N_24975,N_24647);
xor U25877 (N_25877,N_24864,N_24277);
xnor U25878 (N_25878,N_24593,N_24934);
or U25879 (N_25879,N_24937,N_24653);
nand U25880 (N_25880,N_24486,N_24128);
nor U25881 (N_25881,N_24465,N_24468);
and U25882 (N_25882,N_24538,N_24693);
nand U25883 (N_25883,N_24534,N_24712);
nand U25884 (N_25884,N_24245,N_24629);
xnor U25885 (N_25885,N_24518,N_24301);
and U25886 (N_25886,N_24139,N_24504);
or U25887 (N_25887,N_24549,N_24186);
nor U25888 (N_25888,N_24616,N_24891);
nand U25889 (N_25889,N_24508,N_24310);
or U25890 (N_25890,N_24314,N_24898);
nand U25891 (N_25891,N_24123,N_24490);
and U25892 (N_25892,N_24907,N_24638);
xnor U25893 (N_25893,N_24709,N_24060);
or U25894 (N_25894,N_24876,N_24926);
nor U25895 (N_25895,N_24861,N_24811);
nand U25896 (N_25896,N_24552,N_24583);
and U25897 (N_25897,N_24932,N_24595);
or U25898 (N_25898,N_24231,N_24573);
and U25899 (N_25899,N_24117,N_24665);
or U25900 (N_25900,N_24461,N_24203);
and U25901 (N_25901,N_24081,N_24220);
nand U25902 (N_25902,N_24497,N_24356);
nand U25903 (N_25903,N_24783,N_24248);
xnor U25904 (N_25904,N_24260,N_24131);
and U25905 (N_25905,N_24904,N_24690);
nor U25906 (N_25906,N_24989,N_24894);
or U25907 (N_25907,N_24387,N_24832);
xnor U25908 (N_25908,N_24390,N_24425);
nand U25909 (N_25909,N_24046,N_24277);
xor U25910 (N_25910,N_24330,N_24690);
nand U25911 (N_25911,N_24881,N_24914);
or U25912 (N_25912,N_24628,N_24295);
and U25913 (N_25913,N_24484,N_24660);
and U25914 (N_25914,N_24243,N_24503);
nand U25915 (N_25915,N_24655,N_24774);
xor U25916 (N_25916,N_24954,N_24543);
and U25917 (N_25917,N_24174,N_24365);
nand U25918 (N_25918,N_24001,N_24908);
and U25919 (N_25919,N_24425,N_24849);
and U25920 (N_25920,N_24654,N_24555);
nor U25921 (N_25921,N_24081,N_24022);
or U25922 (N_25922,N_24578,N_24752);
xnor U25923 (N_25923,N_24884,N_24668);
xnor U25924 (N_25924,N_24814,N_24694);
or U25925 (N_25925,N_24775,N_24045);
xor U25926 (N_25926,N_24587,N_24139);
nor U25927 (N_25927,N_24232,N_24882);
xor U25928 (N_25928,N_24458,N_24697);
or U25929 (N_25929,N_24759,N_24551);
nor U25930 (N_25930,N_24650,N_24882);
or U25931 (N_25931,N_24804,N_24128);
and U25932 (N_25932,N_24453,N_24653);
xor U25933 (N_25933,N_24006,N_24136);
or U25934 (N_25934,N_24550,N_24461);
nand U25935 (N_25935,N_24188,N_24893);
and U25936 (N_25936,N_24734,N_24808);
and U25937 (N_25937,N_24184,N_24250);
and U25938 (N_25938,N_24523,N_24943);
or U25939 (N_25939,N_24258,N_24220);
and U25940 (N_25940,N_24541,N_24146);
or U25941 (N_25941,N_24009,N_24608);
or U25942 (N_25942,N_24285,N_24392);
or U25943 (N_25943,N_24408,N_24002);
and U25944 (N_25944,N_24730,N_24131);
and U25945 (N_25945,N_24677,N_24530);
and U25946 (N_25946,N_24945,N_24282);
nand U25947 (N_25947,N_24281,N_24560);
nand U25948 (N_25948,N_24622,N_24682);
nand U25949 (N_25949,N_24073,N_24139);
and U25950 (N_25950,N_24081,N_24387);
nor U25951 (N_25951,N_24139,N_24653);
nor U25952 (N_25952,N_24559,N_24047);
or U25953 (N_25953,N_24408,N_24054);
nor U25954 (N_25954,N_24879,N_24937);
nor U25955 (N_25955,N_24206,N_24178);
xor U25956 (N_25956,N_24157,N_24765);
nor U25957 (N_25957,N_24682,N_24077);
nor U25958 (N_25958,N_24480,N_24488);
or U25959 (N_25959,N_24818,N_24387);
and U25960 (N_25960,N_24229,N_24730);
or U25961 (N_25961,N_24927,N_24210);
nand U25962 (N_25962,N_24140,N_24627);
or U25963 (N_25963,N_24848,N_24879);
nand U25964 (N_25964,N_24563,N_24759);
and U25965 (N_25965,N_24142,N_24730);
and U25966 (N_25966,N_24797,N_24328);
or U25967 (N_25967,N_24027,N_24761);
and U25968 (N_25968,N_24127,N_24346);
nand U25969 (N_25969,N_24070,N_24869);
nor U25970 (N_25970,N_24980,N_24100);
or U25971 (N_25971,N_24819,N_24953);
xnor U25972 (N_25972,N_24417,N_24219);
and U25973 (N_25973,N_24453,N_24412);
xnor U25974 (N_25974,N_24562,N_24053);
xnor U25975 (N_25975,N_24875,N_24391);
or U25976 (N_25976,N_24209,N_24618);
and U25977 (N_25977,N_24653,N_24384);
and U25978 (N_25978,N_24566,N_24459);
nor U25979 (N_25979,N_24168,N_24043);
nand U25980 (N_25980,N_24654,N_24897);
xor U25981 (N_25981,N_24943,N_24231);
nor U25982 (N_25982,N_24597,N_24013);
nand U25983 (N_25983,N_24684,N_24766);
or U25984 (N_25984,N_24956,N_24123);
nor U25985 (N_25985,N_24903,N_24027);
or U25986 (N_25986,N_24391,N_24056);
and U25987 (N_25987,N_24653,N_24017);
nand U25988 (N_25988,N_24399,N_24387);
xnor U25989 (N_25989,N_24054,N_24683);
and U25990 (N_25990,N_24753,N_24416);
nand U25991 (N_25991,N_24735,N_24163);
xnor U25992 (N_25992,N_24342,N_24318);
or U25993 (N_25993,N_24728,N_24676);
xor U25994 (N_25994,N_24795,N_24906);
and U25995 (N_25995,N_24196,N_24203);
nand U25996 (N_25996,N_24189,N_24867);
nand U25997 (N_25997,N_24711,N_24176);
nor U25998 (N_25998,N_24875,N_24400);
nand U25999 (N_25999,N_24987,N_24828);
and U26000 (N_26000,N_25060,N_25525);
or U26001 (N_26001,N_25608,N_25615);
or U26002 (N_26002,N_25999,N_25952);
nor U26003 (N_26003,N_25225,N_25792);
or U26004 (N_26004,N_25658,N_25724);
nand U26005 (N_26005,N_25635,N_25119);
nand U26006 (N_26006,N_25392,N_25028);
xor U26007 (N_26007,N_25887,N_25921);
nand U26008 (N_26008,N_25316,N_25086);
nand U26009 (N_26009,N_25955,N_25477);
nand U26010 (N_26010,N_25871,N_25984);
xnor U26011 (N_26011,N_25321,N_25052);
nand U26012 (N_26012,N_25920,N_25003);
nand U26013 (N_26013,N_25718,N_25339);
xor U26014 (N_26014,N_25074,N_25352);
or U26015 (N_26015,N_25323,N_25319);
or U26016 (N_26016,N_25487,N_25864);
xnor U26017 (N_26017,N_25888,N_25757);
and U26018 (N_26018,N_25544,N_25341);
nor U26019 (N_26019,N_25970,N_25595);
or U26020 (N_26020,N_25551,N_25896);
and U26021 (N_26021,N_25479,N_25496);
xor U26022 (N_26022,N_25059,N_25428);
nor U26023 (N_26023,N_25278,N_25530);
nor U26024 (N_26024,N_25072,N_25235);
or U26025 (N_26025,N_25604,N_25163);
and U26026 (N_26026,N_25665,N_25553);
or U26027 (N_26027,N_25241,N_25651);
and U26028 (N_26028,N_25112,N_25866);
nor U26029 (N_26029,N_25532,N_25975);
nor U26030 (N_26030,N_25464,N_25337);
nor U26031 (N_26031,N_25550,N_25066);
nor U26032 (N_26032,N_25628,N_25476);
and U26033 (N_26033,N_25123,N_25274);
and U26034 (N_26034,N_25297,N_25960);
or U26035 (N_26035,N_25092,N_25312);
xor U26036 (N_26036,N_25560,N_25997);
or U26037 (N_26037,N_25648,N_25296);
and U26038 (N_26038,N_25490,N_25200);
nand U26039 (N_26039,N_25106,N_25307);
nor U26040 (N_26040,N_25799,N_25463);
and U26041 (N_26041,N_25501,N_25515);
and U26042 (N_26042,N_25317,N_25047);
xor U26043 (N_26043,N_25558,N_25855);
or U26044 (N_26044,N_25144,N_25354);
and U26045 (N_26045,N_25134,N_25742);
xor U26046 (N_26046,N_25861,N_25147);
or U26047 (N_26047,N_25713,N_25209);
nand U26048 (N_26048,N_25985,N_25589);
and U26049 (N_26049,N_25821,N_25454);
nand U26050 (N_26050,N_25671,N_25136);
or U26051 (N_26051,N_25865,N_25332);
xnor U26052 (N_26052,N_25900,N_25809);
and U26053 (N_26053,N_25655,N_25313);
or U26054 (N_26054,N_25329,N_25844);
nor U26055 (N_26055,N_25221,N_25305);
and U26056 (N_26056,N_25402,N_25890);
and U26057 (N_26057,N_25933,N_25183);
nor U26058 (N_26058,N_25504,N_25155);
xnor U26059 (N_26059,N_25989,N_25764);
nor U26060 (N_26060,N_25666,N_25617);
nor U26061 (N_26061,N_25364,N_25951);
nand U26062 (N_26062,N_25702,N_25720);
or U26063 (N_26063,N_25692,N_25990);
xor U26064 (N_26064,N_25877,N_25876);
nor U26065 (N_26065,N_25233,N_25991);
nand U26066 (N_26066,N_25872,N_25438);
and U26067 (N_26067,N_25475,N_25009);
xnor U26068 (N_26068,N_25973,N_25620);
nor U26069 (N_26069,N_25038,N_25171);
xnor U26070 (N_26070,N_25954,N_25996);
nor U26071 (N_26071,N_25609,N_25833);
or U26072 (N_26072,N_25491,N_25740);
nor U26073 (N_26073,N_25754,N_25619);
or U26074 (N_26074,N_25145,N_25253);
nand U26075 (N_26075,N_25415,N_25834);
nor U26076 (N_26076,N_25424,N_25068);
xnor U26077 (N_26077,N_25566,N_25979);
nand U26078 (N_26078,N_25265,N_25654);
or U26079 (N_26079,N_25852,N_25987);
nand U26080 (N_26080,N_25923,N_25892);
nor U26081 (N_26081,N_25478,N_25242);
nor U26082 (N_26082,N_25427,N_25036);
and U26083 (N_26083,N_25238,N_25937);
nand U26084 (N_26084,N_25875,N_25391);
nand U26085 (N_26085,N_25810,N_25444);
or U26086 (N_26086,N_25250,N_25484);
nand U26087 (N_26087,N_25800,N_25469);
nand U26088 (N_26088,N_25218,N_25915);
nor U26089 (N_26089,N_25432,N_25486);
or U26090 (N_26090,N_25456,N_25010);
nand U26091 (N_26091,N_25054,N_25593);
and U26092 (N_26092,N_25320,N_25738);
nand U26093 (N_26093,N_25000,N_25878);
nand U26094 (N_26094,N_25026,N_25545);
nand U26095 (N_26095,N_25939,N_25465);
nor U26096 (N_26096,N_25762,N_25466);
or U26097 (N_26097,N_25897,N_25363);
nor U26098 (N_26098,N_25790,N_25981);
nor U26099 (N_26099,N_25664,N_25945);
xor U26100 (N_26100,N_25188,N_25881);
nor U26101 (N_26101,N_25166,N_25239);
or U26102 (N_26102,N_25446,N_25344);
nand U26103 (N_26103,N_25678,N_25133);
nor U26104 (N_26104,N_25350,N_25378);
nand U26105 (N_26105,N_25690,N_25271);
and U26106 (N_26106,N_25728,N_25423);
nand U26107 (N_26107,N_25373,N_25934);
nand U26108 (N_26108,N_25051,N_25509);
xor U26109 (N_26109,N_25583,N_25027);
or U26110 (N_26110,N_25158,N_25828);
or U26111 (N_26111,N_25717,N_25013);
xor U26112 (N_26112,N_25244,N_25909);
and U26113 (N_26113,N_25121,N_25267);
and U26114 (N_26114,N_25669,N_25675);
or U26115 (N_26115,N_25845,N_25683);
nor U26116 (N_26116,N_25361,N_25856);
nor U26117 (N_26117,N_25642,N_25063);
or U26118 (N_26118,N_25266,N_25025);
and U26119 (N_26119,N_25611,N_25110);
or U26120 (N_26120,N_25747,N_25069);
and U26121 (N_26121,N_25331,N_25785);
nor U26122 (N_26122,N_25524,N_25204);
nor U26123 (N_26123,N_25021,N_25260);
xor U26124 (N_26124,N_25150,N_25622);
nand U26125 (N_26125,N_25906,N_25837);
nor U26126 (N_26126,N_25259,N_25410);
and U26127 (N_26127,N_25198,N_25342);
or U26128 (N_26128,N_25294,N_25540);
and U26129 (N_26129,N_25967,N_25169);
or U26130 (N_26130,N_25002,N_25753);
nor U26131 (N_26131,N_25722,N_25959);
xnor U26132 (N_26132,N_25823,N_25217);
and U26133 (N_26133,N_25776,N_25505);
nand U26134 (N_26134,N_25159,N_25101);
nor U26135 (N_26135,N_25767,N_25399);
and U26136 (N_26136,N_25448,N_25458);
xor U26137 (N_26137,N_25914,N_25625);
or U26138 (N_26138,N_25298,N_25349);
or U26139 (N_26139,N_25383,N_25246);
xor U26140 (N_26140,N_25730,N_25761);
nor U26141 (N_26141,N_25450,N_25228);
or U26142 (N_26142,N_25019,N_25936);
or U26143 (N_26143,N_25766,N_25699);
or U26144 (N_26144,N_25404,N_25289);
nor U26145 (N_26145,N_25388,N_25237);
xor U26146 (N_26146,N_25079,N_25340);
or U26147 (N_26147,N_25483,N_25122);
nor U26148 (N_26148,N_25971,N_25174);
nor U26149 (N_26149,N_25902,N_25506);
and U26150 (N_26150,N_25771,N_25706);
xor U26151 (N_26151,N_25760,N_25192);
or U26152 (N_26152,N_25024,N_25394);
and U26153 (N_26153,N_25795,N_25310);
nor U26154 (N_26154,N_25564,N_25202);
nand U26155 (N_26155,N_25829,N_25974);
nand U26156 (N_26156,N_25911,N_25338);
nand U26157 (N_26157,N_25847,N_25127);
nand U26158 (N_26158,N_25721,N_25451);
nand U26159 (N_26159,N_25813,N_25115);
nor U26160 (N_26160,N_25434,N_25597);
xor U26161 (N_26161,N_25326,N_25536);
or U26162 (N_26162,N_25226,N_25108);
and U26163 (N_26163,N_25559,N_25268);
xnor U26164 (N_26164,N_25455,N_25901);
xor U26165 (N_26165,N_25033,N_25537);
or U26166 (N_26166,N_25325,N_25711);
nor U26167 (N_26167,N_25978,N_25435);
nor U26168 (N_26168,N_25579,N_25899);
nor U26169 (N_26169,N_25563,N_25815);
nor U26170 (N_26170,N_25705,N_25156);
and U26171 (N_26171,N_25502,N_25405);
nand U26172 (N_26172,N_25610,N_25020);
nor U26173 (N_26173,N_25263,N_25085);
or U26174 (N_26174,N_25205,N_25324);
nand U26175 (N_26175,N_25646,N_25976);
or U26176 (N_26176,N_25222,N_25637);
or U26177 (N_26177,N_25613,N_25950);
nand U26178 (N_26178,N_25573,N_25472);
or U26179 (N_26179,N_25408,N_25067);
or U26180 (N_26180,N_25947,N_25614);
nor U26181 (N_26181,N_25531,N_25445);
or U26182 (N_26182,N_25499,N_25512);
xnor U26183 (N_26183,N_25634,N_25431);
or U26184 (N_26184,N_25756,N_25172);
and U26185 (N_26185,N_25302,N_25794);
nor U26186 (N_26186,N_25346,N_25406);
nand U26187 (N_26187,N_25356,N_25503);
nor U26188 (N_26188,N_25520,N_25014);
xnor U26189 (N_26189,N_25516,N_25149);
nor U26190 (N_26190,N_25796,N_25759);
xnor U26191 (N_26191,N_25591,N_25416);
xor U26192 (N_26192,N_25439,N_25644);
xor U26193 (N_26193,N_25390,N_25585);
nand U26194 (N_26194,N_25175,N_25311);
nand U26195 (N_26195,N_25953,N_25588);
nor U26196 (N_26196,N_25592,N_25443);
nor U26197 (N_26197,N_25185,N_25701);
nand U26198 (N_26198,N_25091,N_25836);
and U26199 (N_26199,N_25519,N_25220);
or U26200 (N_26200,N_25090,N_25186);
or U26201 (N_26201,N_25913,N_25521);
nand U26202 (N_26202,N_25858,N_25929);
nor U26203 (N_26203,N_25602,N_25807);
nor U26204 (N_26204,N_25963,N_25641);
nand U26205 (N_26205,N_25938,N_25420);
xnor U26206 (N_26206,N_25005,N_25926);
nor U26207 (N_26207,N_25284,N_25194);
nand U26208 (N_26208,N_25574,N_25181);
nand U26209 (N_26209,N_25376,N_25853);
or U26210 (N_26210,N_25212,N_25269);
or U26211 (N_26211,N_25580,N_25142);
nor U26212 (N_26212,N_25076,N_25078);
and U26213 (N_26213,N_25965,N_25179);
or U26214 (N_26214,N_25726,N_25854);
and U26215 (N_26215,N_25830,N_25749);
or U26216 (N_26216,N_25869,N_25173);
nand U26217 (N_26217,N_25282,N_25417);
nand U26218 (N_26218,N_25995,N_25680);
xor U26219 (N_26219,N_25916,N_25895);
nor U26220 (N_26220,N_25710,N_25201);
nand U26221 (N_26221,N_25791,N_25359);
nand U26222 (N_26222,N_25782,N_25165);
nand U26223 (N_26223,N_25116,N_25022);
nor U26224 (N_26224,N_25734,N_25017);
nand U26225 (N_26225,N_25983,N_25467);
and U26226 (N_26226,N_25577,N_25774);
and U26227 (N_26227,N_25224,N_25482);
xor U26228 (N_26228,N_25733,N_25429);
nor U26229 (N_26229,N_25012,N_25040);
xor U26230 (N_26230,N_25743,N_25393);
nand U26231 (N_26231,N_25397,N_25041);
nand U26232 (N_26232,N_25696,N_25309);
nor U26233 (N_26233,N_25961,N_25632);
and U26234 (N_26234,N_25640,N_25154);
xor U26235 (N_26235,N_25351,N_25409);
or U26236 (N_26236,N_25568,N_25780);
nand U26237 (N_26237,N_25746,N_25880);
and U26238 (N_26238,N_25407,N_25518);
and U26239 (N_26239,N_25709,N_25177);
nor U26240 (N_26240,N_25453,N_25264);
xor U26241 (N_26241,N_25249,N_25691);
xnor U26242 (N_26242,N_25770,N_25223);
nor U26243 (N_26243,N_25668,N_25629);
nand U26244 (N_26244,N_25578,N_25258);
xnor U26245 (N_26245,N_25657,N_25576);
and U26246 (N_26246,N_25290,N_25081);
or U26247 (N_26247,N_25280,N_25497);
xor U26248 (N_26248,N_25411,N_25300);
xor U26249 (N_26249,N_25414,N_25131);
nor U26250 (N_26250,N_25433,N_25527);
xor U26251 (N_26251,N_25748,N_25046);
or U26252 (N_26252,N_25386,N_25943);
nor U26253 (N_26253,N_25215,N_25379);
xor U26254 (N_26254,N_25584,N_25304);
or U26255 (N_26255,N_25511,N_25184);
or U26256 (N_26256,N_25306,N_25167);
xor U26257 (N_26257,N_25686,N_25492);
nor U26258 (N_26258,N_25885,N_25120);
xor U26259 (N_26259,N_25928,N_25917);
nor U26260 (N_26260,N_25286,N_25562);
nor U26261 (N_26261,N_25396,N_25883);
or U26262 (N_26262,N_25840,N_25548);
nand U26263 (N_26263,N_25698,N_25931);
nand U26264 (N_26264,N_25045,N_25832);
nand U26265 (N_26265,N_25526,N_25556);
nand U26266 (N_26266,N_25822,N_25168);
nand U26267 (N_26267,N_25073,N_25732);
or U26268 (N_26268,N_25114,N_25755);
nand U26269 (N_26269,N_25727,N_25839);
nand U26270 (N_26270,N_25797,N_25571);
xnor U26271 (N_26271,N_25130,N_25627);
nand U26272 (N_26272,N_25542,N_25102);
or U26273 (N_26273,N_25164,N_25247);
or U26274 (N_26274,N_25964,N_25712);
and U26275 (N_26275,N_25170,N_25656);
or U26276 (N_26276,N_25368,N_25485);
nor U26277 (N_26277,N_25500,N_25674);
nand U26278 (N_26278,N_25663,N_25030);
xor U26279 (N_26279,N_25176,N_25365);
nand U26280 (N_26280,N_25057,N_25196);
nand U26281 (N_26281,N_25043,N_25327);
xnor U26282 (N_26282,N_25137,N_25787);
xnor U26283 (N_26283,N_25489,N_25135);
nor U26284 (N_26284,N_25422,N_25208);
xnor U26285 (N_26285,N_25703,N_25334);
nand U26286 (N_26286,N_25898,N_25605);
and U26287 (N_26287,N_25626,N_25940);
xor U26288 (N_26288,N_25752,N_25513);
or U26289 (N_26289,N_25843,N_25214);
nand U26290 (N_26290,N_25372,N_25357);
nand U26291 (N_26291,N_25660,N_25251);
and U26292 (N_26292,N_25004,N_25918);
or U26293 (N_26293,N_25105,N_25704);
nor U26294 (N_26294,N_25825,N_25650);
or U26295 (N_26295,N_25211,N_25495);
nand U26296 (N_26296,N_25946,N_25670);
or U26297 (N_26297,N_25412,N_25460);
and U26298 (N_26298,N_25874,N_25886);
or U26299 (N_26299,N_25784,N_25581);
nand U26300 (N_26300,N_25193,N_25459);
or U26301 (N_26301,N_25835,N_25925);
and U26302 (N_26302,N_25380,N_25493);
or U26303 (N_26303,N_25023,N_25889);
and U26304 (N_26304,N_25143,N_25707);
nor U26305 (N_26305,N_25860,N_25178);
xor U26306 (N_26306,N_25769,N_25811);
and U26307 (N_26307,N_25227,N_25859);
xnor U26308 (N_26308,N_25494,N_25461);
or U26309 (N_26309,N_25481,N_25977);
nand U26310 (N_26310,N_25343,N_25160);
nand U26311 (N_26311,N_25744,N_25993);
or U26312 (N_26312,N_25647,N_25189);
xor U26313 (N_26313,N_25814,N_25262);
xor U26314 (N_26314,N_25912,N_25695);
or U26315 (N_26315,N_25089,N_25803);
xor U26316 (N_26316,N_25180,N_25944);
and U26317 (N_26317,N_25930,N_25863);
or U26318 (N_26318,N_25042,N_25058);
and U26319 (N_26319,N_25333,N_25561);
or U26320 (N_26320,N_25206,N_25956);
nor U26321 (N_26321,N_25624,N_25100);
or U26322 (N_26322,N_25598,N_25232);
nor U26323 (N_26323,N_25781,N_25008);
nand U26324 (N_26324,N_25966,N_25449);
xor U26325 (N_26325,N_25590,N_25295);
xor U26326 (N_26326,N_25255,N_25011);
nand U26327 (N_26327,N_25162,N_25270);
and U26328 (N_26328,N_25685,N_25768);
xnor U26329 (N_26329,N_25681,N_25739);
and U26330 (N_26330,N_25355,N_25216);
nor U26331 (N_26331,N_25533,N_25549);
nand U26332 (N_26332,N_25037,N_25015);
nor U26333 (N_26333,N_25082,N_25219);
or U26334 (N_26334,N_25245,N_25382);
or U26335 (N_26335,N_25161,N_25430);
or U26336 (N_26336,N_25437,N_25841);
xor U26337 (N_26337,N_25032,N_25293);
nor U26338 (N_26338,N_25735,N_25994);
or U26339 (N_26339,N_25229,N_25285);
nand U26340 (N_26340,N_25345,N_25824);
nand U26341 (N_26341,N_25389,N_25367);
nor U26342 (N_26342,N_25689,N_25031);
xor U26343 (N_26343,N_25126,N_25603);
nor U26344 (N_26344,N_25498,N_25371);
and U26345 (N_26345,N_25777,N_25765);
or U26346 (N_26346,N_25779,N_25827);
xor U26347 (N_26347,N_25029,N_25109);
nand U26348 (N_26348,N_25441,N_25099);
and U26349 (N_26349,N_25398,N_25948);
or U26350 (N_26350,N_25488,N_25426);
nand U26351 (N_26351,N_25335,N_25256);
and U26352 (N_26352,N_25056,N_25210);
and U26353 (N_26353,N_25972,N_25107);
and U26354 (N_26354,N_25132,N_25567);
nand U26355 (N_26355,N_25236,N_25187);
nor U26356 (N_26356,N_25862,N_25763);
nor U26357 (N_26357,N_25207,N_25927);
nor U26358 (N_26358,N_25276,N_25694);
or U26359 (N_26359,N_25653,N_25893);
or U26360 (N_26360,N_25384,N_25330);
or U26361 (N_26361,N_25808,N_25922);
and U26362 (N_26362,N_25894,N_25191);
or U26363 (N_26363,N_25572,N_25879);
nor U26364 (N_26364,N_25070,N_25118);
xnor U26365 (N_26365,N_25700,N_25804);
or U26366 (N_26366,N_25789,N_25962);
nand U26367 (N_26367,N_25360,N_25715);
xor U26368 (N_26368,N_25254,N_25197);
nor U26369 (N_26369,N_25607,N_25601);
nor U26370 (N_26370,N_25374,N_25786);
or U26371 (N_26371,N_25273,N_25992);
nor U26372 (N_26372,N_25838,N_25908);
nor U26373 (N_26373,N_25462,N_25805);
nor U26374 (N_26374,N_25366,N_25693);
or U26375 (N_26375,N_25633,N_25231);
xor U26376 (N_26376,N_25287,N_25958);
or U26377 (N_26377,N_25528,N_25016);
nand U26378 (N_26378,N_25793,N_25138);
xor U26379 (N_26379,N_25942,N_25292);
nand U26380 (N_26380,N_25075,N_25140);
nor U26381 (N_26381,N_25124,N_25514);
or U26382 (N_26382,N_25870,N_25157);
nor U26383 (N_26383,N_25190,N_25905);
nand U26384 (N_26384,N_25554,N_25148);
or U26385 (N_26385,N_25095,N_25988);
or U26386 (N_26386,N_25385,N_25903);
or U26387 (N_26387,N_25842,N_25778);
and U26388 (N_26388,N_25358,N_25517);
and U26389 (N_26389,N_25006,N_25606);
nor U26390 (N_26390,N_25322,N_25257);
nor U26391 (N_26391,N_25638,N_25203);
nand U26392 (N_26392,N_25672,N_25275);
or U26393 (N_26393,N_25812,N_25652);
or U26394 (N_26394,N_25725,N_25096);
nand U26395 (N_26395,N_25400,N_25375);
and U26396 (N_26396,N_25369,N_25111);
or U26397 (N_26397,N_25403,N_25139);
or U26398 (N_26398,N_25104,N_25649);
or U26399 (N_26399,N_25783,N_25473);
nand U26400 (N_26400,N_25442,N_25141);
nand U26401 (N_26401,N_25729,N_25555);
or U26402 (N_26402,N_25071,N_25570);
and U26403 (N_26403,N_25199,N_25234);
nand U26404 (N_26404,N_25684,N_25088);
or U26405 (N_26405,N_25094,N_25596);
xor U26406 (N_26406,N_25818,N_25957);
or U26407 (N_26407,N_25529,N_25968);
xor U26408 (N_26408,N_25986,N_25582);
xor U26409 (N_26409,N_25117,N_25687);
and U26410 (N_26410,N_25087,N_25736);
or U26411 (N_26411,N_25884,N_25594);
nand U26412 (N_26412,N_25065,N_25418);
xnor U26413 (N_26413,N_25639,N_25819);
or U26414 (N_26414,N_25851,N_25673);
and U26415 (N_26415,N_25452,N_25053);
xor U26416 (N_26416,N_25806,N_25659);
xnor U26417 (N_26417,N_25662,N_25301);
nor U26418 (N_26418,N_25569,N_25826);
nor U26419 (N_26419,N_25077,N_25539);
or U26420 (N_26420,N_25924,N_25919);
or U26421 (N_26421,N_25623,N_25314);
nor U26422 (N_26422,N_25534,N_25281);
and U26423 (N_26423,N_25816,N_25631);
xnor U26424 (N_26424,N_25413,N_25001);
xnor U26425 (N_26425,N_25867,N_25708);
or U26426 (N_26426,N_25440,N_25616);
and U26427 (N_26427,N_25347,N_25480);
nor U26428 (N_26428,N_25758,N_25291);
and U26429 (N_26429,N_25688,N_25612);
and U26430 (N_26430,N_25788,N_25745);
nand U26431 (N_26431,N_25436,N_25272);
and U26432 (N_26432,N_25050,N_25677);
nor U26433 (N_26433,N_25510,N_25381);
nand U26434 (N_26434,N_25716,N_25507);
nor U26435 (N_26435,N_25261,N_25538);
nand U26436 (N_26436,N_25575,N_25007);
or U26437 (N_26437,N_25714,N_25868);
nor U26438 (N_26438,N_25128,N_25831);
nor U26439 (N_26439,N_25565,N_25543);
nor U26440 (N_26440,N_25820,N_25103);
nand U26441 (N_26441,N_25857,N_25801);
and U26442 (N_26442,N_25775,N_25315);
nor U26443 (N_26443,N_25904,N_25750);
and U26444 (N_26444,N_25048,N_25798);
xnor U26445 (N_26445,N_25283,N_25395);
nand U26446 (N_26446,N_25679,N_25098);
or U26447 (N_26447,N_25719,N_25998);
or U26448 (N_26448,N_25370,N_25636);
xor U26449 (N_26449,N_25277,N_25055);
xnor U26450 (N_26450,N_25093,N_25299);
or U26451 (N_26451,N_25034,N_25535);
nor U26452 (N_26452,N_25982,N_25949);
and U26453 (N_26453,N_25308,N_25471);
and U26454 (N_26454,N_25248,N_25547);
or U26455 (N_26455,N_25802,N_25113);
nor U26456 (N_26456,N_25252,N_25129);
nor U26457 (N_26457,N_25362,N_25062);
nor U26458 (N_26458,N_25523,N_25682);
nor U26459 (N_26459,N_25049,N_25064);
nor U26460 (N_26460,N_25522,N_25097);
xnor U26461 (N_26461,N_25980,N_25891);
xnor U26462 (N_26462,N_25546,N_25941);
nand U26463 (N_26463,N_25773,N_25600);
or U26464 (N_26464,N_25661,N_25772);
or U26465 (N_26465,N_25039,N_25182);
nand U26466 (N_26466,N_25468,N_25318);
xor U26467 (N_26467,N_25586,N_25969);
nor U26468 (N_26468,N_25035,N_25401);
xor U26469 (N_26469,N_25645,N_25723);
xor U26470 (N_26470,N_25932,N_25817);
nor U26471 (N_26471,N_25353,N_25618);
nand U26472 (N_26472,N_25676,N_25080);
or U26473 (N_26473,N_25470,N_25328);
xor U26474 (N_26474,N_25213,N_25146);
xor U26475 (N_26475,N_25377,N_25474);
xor U26476 (N_26476,N_25731,N_25387);
xnor U26477 (N_26477,N_25425,N_25552);
nand U26478 (N_26478,N_25421,N_25419);
nand U26479 (N_26479,N_25152,N_25240);
xnor U26480 (N_26480,N_25348,N_25195);
and U26481 (N_26481,N_25667,N_25083);
and U26482 (N_26482,N_25910,N_25279);
or U26483 (N_26483,N_25630,N_25741);
xor U26484 (N_26484,N_25873,N_25850);
or U26485 (N_26485,N_25751,N_25907);
or U26486 (N_26486,N_25541,N_25848);
nor U26487 (N_26487,N_25846,N_25336);
xor U26488 (N_26488,N_25508,N_25303);
or U26489 (N_26489,N_25288,N_25737);
xnor U26490 (N_26490,N_25061,N_25882);
nand U26491 (N_26491,N_25044,N_25084);
xor U26492 (N_26492,N_25557,N_25153);
nand U26493 (N_26493,N_25230,N_25457);
nand U26494 (N_26494,N_25849,N_25599);
and U26495 (N_26495,N_25621,N_25125);
xnor U26496 (N_26496,N_25697,N_25447);
nor U26497 (N_26497,N_25935,N_25643);
nand U26498 (N_26498,N_25151,N_25243);
nand U26499 (N_26499,N_25587,N_25018);
xor U26500 (N_26500,N_25824,N_25328);
xor U26501 (N_26501,N_25339,N_25097);
nand U26502 (N_26502,N_25235,N_25076);
and U26503 (N_26503,N_25968,N_25704);
and U26504 (N_26504,N_25363,N_25400);
or U26505 (N_26505,N_25237,N_25571);
nor U26506 (N_26506,N_25294,N_25962);
nor U26507 (N_26507,N_25119,N_25574);
nor U26508 (N_26508,N_25394,N_25671);
nor U26509 (N_26509,N_25378,N_25647);
or U26510 (N_26510,N_25997,N_25802);
nor U26511 (N_26511,N_25600,N_25531);
or U26512 (N_26512,N_25362,N_25998);
and U26513 (N_26513,N_25826,N_25196);
or U26514 (N_26514,N_25522,N_25929);
nor U26515 (N_26515,N_25156,N_25101);
or U26516 (N_26516,N_25925,N_25898);
nand U26517 (N_26517,N_25721,N_25529);
or U26518 (N_26518,N_25891,N_25787);
or U26519 (N_26519,N_25772,N_25482);
or U26520 (N_26520,N_25853,N_25136);
nand U26521 (N_26521,N_25629,N_25418);
nor U26522 (N_26522,N_25781,N_25777);
or U26523 (N_26523,N_25008,N_25278);
nor U26524 (N_26524,N_25872,N_25489);
nand U26525 (N_26525,N_25646,N_25027);
nand U26526 (N_26526,N_25267,N_25924);
nand U26527 (N_26527,N_25552,N_25189);
and U26528 (N_26528,N_25583,N_25741);
nand U26529 (N_26529,N_25302,N_25595);
or U26530 (N_26530,N_25043,N_25695);
and U26531 (N_26531,N_25677,N_25071);
and U26532 (N_26532,N_25570,N_25930);
or U26533 (N_26533,N_25646,N_25767);
nor U26534 (N_26534,N_25602,N_25434);
xnor U26535 (N_26535,N_25624,N_25348);
nand U26536 (N_26536,N_25124,N_25698);
nor U26537 (N_26537,N_25758,N_25729);
and U26538 (N_26538,N_25393,N_25588);
nand U26539 (N_26539,N_25753,N_25413);
xor U26540 (N_26540,N_25522,N_25895);
or U26541 (N_26541,N_25342,N_25321);
xor U26542 (N_26542,N_25200,N_25102);
and U26543 (N_26543,N_25283,N_25435);
and U26544 (N_26544,N_25437,N_25770);
xor U26545 (N_26545,N_25906,N_25863);
or U26546 (N_26546,N_25787,N_25032);
nor U26547 (N_26547,N_25640,N_25867);
nand U26548 (N_26548,N_25442,N_25832);
or U26549 (N_26549,N_25003,N_25821);
nor U26550 (N_26550,N_25443,N_25303);
nor U26551 (N_26551,N_25144,N_25969);
or U26552 (N_26552,N_25786,N_25655);
xnor U26553 (N_26553,N_25078,N_25871);
or U26554 (N_26554,N_25505,N_25257);
xor U26555 (N_26555,N_25145,N_25084);
or U26556 (N_26556,N_25556,N_25580);
nand U26557 (N_26557,N_25889,N_25965);
nor U26558 (N_26558,N_25019,N_25657);
or U26559 (N_26559,N_25077,N_25047);
xnor U26560 (N_26560,N_25544,N_25319);
xor U26561 (N_26561,N_25444,N_25003);
or U26562 (N_26562,N_25040,N_25561);
nor U26563 (N_26563,N_25958,N_25994);
nand U26564 (N_26564,N_25287,N_25851);
or U26565 (N_26565,N_25375,N_25783);
xor U26566 (N_26566,N_25540,N_25738);
or U26567 (N_26567,N_25726,N_25580);
nand U26568 (N_26568,N_25500,N_25768);
or U26569 (N_26569,N_25939,N_25467);
nand U26570 (N_26570,N_25667,N_25336);
nand U26571 (N_26571,N_25180,N_25943);
and U26572 (N_26572,N_25651,N_25017);
nand U26573 (N_26573,N_25516,N_25735);
xnor U26574 (N_26574,N_25650,N_25455);
nor U26575 (N_26575,N_25229,N_25539);
or U26576 (N_26576,N_25413,N_25889);
and U26577 (N_26577,N_25700,N_25989);
or U26578 (N_26578,N_25042,N_25913);
xnor U26579 (N_26579,N_25940,N_25314);
xor U26580 (N_26580,N_25692,N_25721);
nor U26581 (N_26581,N_25541,N_25190);
nor U26582 (N_26582,N_25594,N_25488);
nor U26583 (N_26583,N_25333,N_25448);
and U26584 (N_26584,N_25328,N_25118);
nand U26585 (N_26585,N_25991,N_25887);
nand U26586 (N_26586,N_25029,N_25980);
xnor U26587 (N_26587,N_25414,N_25693);
or U26588 (N_26588,N_25022,N_25095);
xnor U26589 (N_26589,N_25791,N_25100);
nand U26590 (N_26590,N_25405,N_25698);
nand U26591 (N_26591,N_25227,N_25189);
or U26592 (N_26592,N_25551,N_25248);
nand U26593 (N_26593,N_25196,N_25915);
nand U26594 (N_26594,N_25842,N_25421);
and U26595 (N_26595,N_25105,N_25266);
or U26596 (N_26596,N_25369,N_25632);
nand U26597 (N_26597,N_25232,N_25825);
xor U26598 (N_26598,N_25519,N_25912);
xnor U26599 (N_26599,N_25015,N_25910);
nand U26600 (N_26600,N_25715,N_25154);
nand U26601 (N_26601,N_25266,N_25628);
or U26602 (N_26602,N_25420,N_25281);
nand U26603 (N_26603,N_25212,N_25168);
nand U26604 (N_26604,N_25947,N_25783);
nor U26605 (N_26605,N_25479,N_25958);
nand U26606 (N_26606,N_25822,N_25092);
and U26607 (N_26607,N_25873,N_25105);
nand U26608 (N_26608,N_25181,N_25394);
or U26609 (N_26609,N_25291,N_25319);
nor U26610 (N_26610,N_25586,N_25495);
xnor U26611 (N_26611,N_25544,N_25439);
or U26612 (N_26612,N_25653,N_25457);
nor U26613 (N_26613,N_25674,N_25506);
and U26614 (N_26614,N_25303,N_25522);
and U26615 (N_26615,N_25284,N_25676);
or U26616 (N_26616,N_25385,N_25150);
or U26617 (N_26617,N_25347,N_25774);
and U26618 (N_26618,N_25359,N_25199);
and U26619 (N_26619,N_25917,N_25252);
and U26620 (N_26620,N_25146,N_25725);
xor U26621 (N_26621,N_25473,N_25121);
nand U26622 (N_26622,N_25865,N_25624);
nor U26623 (N_26623,N_25498,N_25459);
or U26624 (N_26624,N_25619,N_25067);
or U26625 (N_26625,N_25227,N_25758);
or U26626 (N_26626,N_25743,N_25185);
nor U26627 (N_26627,N_25858,N_25513);
and U26628 (N_26628,N_25294,N_25848);
xor U26629 (N_26629,N_25036,N_25639);
nand U26630 (N_26630,N_25846,N_25765);
and U26631 (N_26631,N_25450,N_25430);
or U26632 (N_26632,N_25426,N_25101);
and U26633 (N_26633,N_25812,N_25444);
nand U26634 (N_26634,N_25274,N_25140);
or U26635 (N_26635,N_25208,N_25165);
xor U26636 (N_26636,N_25684,N_25937);
or U26637 (N_26637,N_25673,N_25855);
nand U26638 (N_26638,N_25681,N_25853);
and U26639 (N_26639,N_25073,N_25383);
or U26640 (N_26640,N_25873,N_25484);
nor U26641 (N_26641,N_25754,N_25168);
nor U26642 (N_26642,N_25008,N_25512);
nand U26643 (N_26643,N_25816,N_25428);
nor U26644 (N_26644,N_25852,N_25014);
xor U26645 (N_26645,N_25633,N_25749);
and U26646 (N_26646,N_25486,N_25066);
or U26647 (N_26647,N_25944,N_25442);
or U26648 (N_26648,N_25246,N_25650);
xnor U26649 (N_26649,N_25864,N_25182);
xnor U26650 (N_26650,N_25971,N_25162);
and U26651 (N_26651,N_25579,N_25907);
or U26652 (N_26652,N_25598,N_25253);
nand U26653 (N_26653,N_25811,N_25923);
nor U26654 (N_26654,N_25589,N_25267);
xor U26655 (N_26655,N_25891,N_25185);
nor U26656 (N_26656,N_25663,N_25659);
xnor U26657 (N_26657,N_25390,N_25711);
xnor U26658 (N_26658,N_25405,N_25513);
nor U26659 (N_26659,N_25995,N_25508);
nor U26660 (N_26660,N_25201,N_25669);
and U26661 (N_26661,N_25930,N_25046);
or U26662 (N_26662,N_25074,N_25975);
nand U26663 (N_26663,N_25857,N_25358);
and U26664 (N_26664,N_25813,N_25870);
nand U26665 (N_26665,N_25886,N_25100);
nor U26666 (N_26666,N_25429,N_25613);
and U26667 (N_26667,N_25608,N_25574);
or U26668 (N_26668,N_25490,N_25839);
nor U26669 (N_26669,N_25756,N_25664);
nand U26670 (N_26670,N_25224,N_25884);
or U26671 (N_26671,N_25560,N_25943);
or U26672 (N_26672,N_25105,N_25887);
or U26673 (N_26673,N_25418,N_25241);
nor U26674 (N_26674,N_25847,N_25387);
nand U26675 (N_26675,N_25487,N_25617);
or U26676 (N_26676,N_25860,N_25639);
or U26677 (N_26677,N_25939,N_25940);
or U26678 (N_26678,N_25383,N_25530);
or U26679 (N_26679,N_25193,N_25079);
nor U26680 (N_26680,N_25023,N_25706);
nand U26681 (N_26681,N_25396,N_25924);
and U26682 (N_26682,N_25145,N_25081);
xor U26683 (N_26683,N_25021,N_25172);
and U26684 (N_26684,N_25188,N_25623);
nand U26685 (N_26685,N_25341,N_25641);
and U26686 (N_26686,N_25449,N_25367);
nor U26687 (N_26687,N_25006,N_25918);
or U26688 (N_26688,N_25682,N_25973);
nand U26689 (N_26689,N_25733,N_25291);
and U26690 (N_26690,N_25850,N_25514);
and U26691 (N_26691,N_25968,N_25370);
and U26692 (N_26692,N_25129,N_25965);
xor U26693 (N_26693,N_25306,N_25583);
and U26694 (N_26694,N_25553,N_25518);
nand U26695 (N_26695,N_25404,N_25218);
nand U26696 (N_26696,N_25035,N_25629);
and U26697 (N_26697,N_25610,N_25974);
nand U26698 (N_26698,N_25829,N_25509);
nor U26699 (N_26699,N_25572,N_25856);
or U26700 (N_26700,N_25724,N_25321);
nand U26701 (N_26701,N_25270,N_25733);
and U26702 (N_26702,N_25650,N_25190);
and U26703 (N_26703,N_25317,N_25080);
xor U26704 (N_26704,N_25399,N_25205);
and U26705 (N_26705,N_25074,N_25120);
or U26706 (N_26706,N_25164,N_25701);
or U26707 (N_26707,N_25705,N_25358);
nand U26708 (N_26708,N_25561,N_25054);
or U26709 (N_26709,N_25806,N_25614);
or U26710 (N_26710,N_25660,N_25404);
or U26711 (N_26711,N_25585,N_25527);
xnor U26712 (N_26712,N_25511,N_25046);
nand U26713 (N_26713,N_25962,N_25151);
xnor U26714 (N_26714,N_25988,N_25322);
xor U26715 (N_26715,N_25504,N_25282);
or U26716 (N_26716,N_25378,N_25980);
and U26717 (N_26717,N_25726,N_25544);
nor U26718 (N_26718,N_25278,N_25204);
nor U26719 (N_26719,N_25016,N_25398);
nor U26720 (N_26720,N_25632,N_25956);
nand U26721 (N_26721,N_25802,N_25722);
nand U26722 (N_26722,N_25416,N_25715);
nand U26723 (N_26723,N_25966,N_25442);
nand U26724 (N_26724,N_25909,N_25894);
xor U26725 (N_26725,N_25444,N_25599);
nor U26726 (N_26726,N_25430,N_25635);
xor U26727 (N_26727,N_25641,N_25660);
nor U26728 (N_26728,N_25307,N_25789);
xnor U26729 (N_26729,N_25609,N_25685);
nand U26730 (N_26730,N_25382,N_25814);
nor U26731 (N_26731,N_25359,N_25215);
xnor U26732 (N_26732,N_25856,N_25803);
nor U26733 (N_26733,N_25654,N_25233);
or U26734 (N_26734,N_25058,N_25772);
xor U26735 (N_26735,N_25536,N_25053);
nand U26736 (N_26736,N_25472,N_25395);
and U26737 (N_26737,N_25121,N_25919);
and U26738 (N_26738,N_25189,N_25480);
xnor U26739 (N_26739,N_25526,N_25519);
nand U26740 (N_26740,N_25184,N_25898);
and U26741 (N_26741,N_25956,N_25512);
nand U26742 (N_26742,N_25312,N_25512);
and U26743 (N_26743,N_25071,N_25543);
nand U26744 (N_26744,N_25570,N_25827);
nand U26745 (N_26745,N_25406,N_25936);
nor U26746 (N_26746,N_25762,N_25249);
xor U26747 (N_26747,N_25548,N_25124);
and U26748 (N_26748,N_25909,N_25905);
and U26749 (N_26749,N_25282,N_25137);
xnor U26750 (N_26750,N_25465,N_25579);
or U26751 (N_26751,N_25355,N_25188);
and U26752 (N_26752,N_25012,N_25197);
or U26753 (N_26753,N_25386,N_25913);
nand U26754 (N_26754,N_25189,N_25271);
nor U26755 (N_26755,N_25274,N_25999);
nor U26756 (N_26756,N_25006,N_25936);
and U26757 (N_26757,N_25112,N_25483);
xnor U26758 (N_26758,N_25681,N_25430);
or U26759 (N_26759,N_25693,N_25656);
or U26760 (N_26760,N_25912,N_25626);
nand U26761 (N_26761,N_25389,N_25905);
and U26762 (N_26762,N_25493,N_25663);
and U26763 (N_26763,N_25751,N_25147);
nor U26764 (N_26764,N_25074,N_25055);
or U26765 (N_26765,N_25112,N_25011);
nand U26766 (N_26766,N_25789,N_25205);
xor U26767 (N_26767,N_25061,N_25634);
nor U26768 (N_26768,N_25286,N_25046);
nand U26769 (N_26769,N_25436,N_25449);
nor U26770 (N_26770,N_25720,N_25673);
or U26771 (N_26771,N_25790,N_25798);
nor U26772 (N_26772,N_25726,N_25063);
nand U26773 (N_26773,N_25345,N_25095);
nor U26774 (N_26774,N_25576,N_25364);
or U26775 (N_26775,N_25036,N_25941);
nor U26776 (N_26776,N_25327,N_25623);
nor U26777 (N_26777,N_25838,N_25468);
nor U26778 (N_26778,N_25891,N_25616);
xor U26779 (N_26779,N_25147,N_25034);
xor U26780 (N_26780,N_25631,N_25082);
nand U26781 (N_26781,N_25738,N_25537);
nor U26782 (N_26782,N_25613,N_25829);
or U26783 (N_26783,N_25011,N_25387);
nand U26784 (N_26784,N_25390,N_25956);
nor U26785 (N_26785,N_25086,N_25134);
nor U26786 (N_26786,N_25853,N_25689);
nand U26787 (N_26787,N_25800,N_25539);
or U26788 (N_26788,N_25337,N_25364);
nand U26789 (N_26789,N_25857,N_25729);
nor U26790 (N_26790,N_25244,N_25700);
or U26791 (N_26791,N_25453,N_25466);
nor U26792 (N_26792,N_25796,N_25349);
nand U26793 (N_26793,N_25744,N_25959);
nand U26794 (N_26794,N_25368,N_25026);
xnor U26795 (N_26795,N_25506,N_25887);
or U26796 (N_26796,N_25056,N_25398);
xor U26797 (N_26797,N_25392,N_25358);
xnor U26798 (N_26798,N_25041,N_25827);
nand U26799 (N_26799,N_25501,N_25587);
nand U26800 (N_26800,N_25001,N_25855);
nor U26801 (N_26801,N_25623,N_25573);
and U26802 (N_26802,N_25011,N_25699);
and U26803 (N_26803,N_25075,N_25415);
xnor U26804 (N_26804,N_25043,N_25213);
xnor U26805 (N_26805,N_25064,N_25939);
and U26806 (N_26806,N_25235,N_25383);
or U26807 (N_26807,N_25205,N_25748);
and U26808 (N_26808,N_25734,N_25919);
xor U26809 (N_26809,N_25166,N_25777);
xnor U26810 (N_26810,N_25878,N_25846);
or U26811 (N_26811,N_25096,N_25508);
and U26812 (N_26812,N_25551,N_25449);
or U26813 (N_26813,N_25590,N_25767);
or U26814 (N_26814,N_25134,N_25492);
nor U26815 (N_26815,N_25740,N_25321);
and U26816 (N_26816,N_25569,N_25191);
and U26817 (N_26817,N_25449,N_25321);
or U26818 (N_26818,N_25867,N_25921);
xor U26819 (N_26819,N_25354,N_25458);
and U26820 (N_26820,N_25189,N_25358);
and U26821 (N_26821,N_25361,N_25532);
or U26822 (N_26822,N_25803,N_25866);
xor U26823 (N_26823,N_25206,N_25017);
nor U26824 (N_26824,N_25405,N_25221);
xnor U26825 (N_26825,N_25125,N_25791);
nor U26826 (N_26826,N_25774,N_25861);
xnor U26827 (N_26827,N_25725,N_25399);
or U26828 (N_26828,N_25731,N_25943);
or U26829 (N_26829,N_25576,N_25451);
and U26830 (N_26830,N_25809,N_25163);
and U26831 (N_26831,N_25918,N_25516);
nand U26832 (N_26832,N_25875,N_25649);
nand U26833 (N_26833,N_25175,N_25995);
or U26834 (N_26834,N_25946,N_25673);
or U26835 (N_26835,N_25984,N_25826);
and U26836 (N_26836,N_25382,N_25088);
xor U26837 (N_26837,N_25805,N_25083);
and U26838 (N_26838,N_25439,N_25017);
and U26839 (N_26839,N_25504,N_25358);
nor U26840 (N_26840,N_25029,N_25825);
nand U26841 (N_26841,N_25116,N_25701);
and U26842 (N_26842,N_25035,N_25459);
and U26843 (N_26843,N_25242,N_25067);
and U26844 (N_26844,N_25375,N_25931);
or U26845 (N_26845,N_25772,N_25459);
nand U26846 (N_26846,N_25746,N_25382);
and U26847 (N_26847,N_25917,N_25299);
or U26848 (N_26848,N_25481,N_25546);
and U26849 (N_26849,N_25893,N_25149);
and U26850 (N_26850,N_25815,N_25235);
or U26851 (N_26851,N_25665,N_25452);
xnor U26852 (N_26852,N_25986,N_25025);
and U26853 (N_26853,N_25767,N_25668);
and U26854 (N_26854,N_25861,N_25571);
nor U26855 (N_26855,N_25391,N_25658);
xnor U26856 (N_26856,N_25403,N_25315);
nor U26857 (N_26857,N_25635,N_25349);
xor U26858 (N_26858,N_25540,N_25918);
nor U26859 (N_26859,N_25869,N_25672);
or U26860 (N_26860,N_25790,N_25480);
xor U26861 (N_26861,N_25919,N_25134);
or U26862 (N_26862,N_25434,N_25059);
nand U26863 (N_26863,N_25391,N_25051);
nor U26864 (N_26864,N_25233,N_25492);
nand U26865 (N_26865,N_25551,N_25767);
nor U26866 (N_26866,N_25126,N_25549);
xor U26867 (N_26867,N_25998,N_25755);
or U26868 (N_26868,N_25416,N_25744);
or U26869 (N_26869,N_25795,N_25827);
nor U26870 (N_26870,N_25863,N_25097);
or U26871 (N_26871,N_25392,N_25373);
nor U26872 (N_26872,N_25218,N_25758);
nor U26873 (N_26873,N_25702,N_25385);
nor U26874 (N_26874,N_25245,N_25408);
nor U26875 (N_26875,N_25490,N_25472);
xnor U26876 (N_26876,N_25119,N_25117);
or U26877 (N_26877,N_25369,N_25682);
and U26878 (N_26878,N_25502,N_25687);
and U26879 (N_26879,N_25757,N_25967);
xnor U26880 (N_26880,N_25003,N_25186);
nor U26881 (N_26881,N_25962,N_25589);
and U26882 (N_26882,N_25976,N_25550);
or U26883 (N_26883,N_25131,N_25477);
and U26884 (N_26884,N_25373,N_25947);
xnor U26885 (N_26885,N_25779,N_25280);
or U26886 (N_26886,N_25685,N_25514);
nand U26887 (N_26887,N_25041,N_25233);
or U26888 (N_26888,N_25215,N_25723);
nand U26889 (N_26889,N_25122,N_25356);
or U26890 (N_26890,N_25725,N_25083);
xor U26891 (N_26891,N_25286,N_25469);
or U26892 (N_26892,N_25852,N_25303);
nand U26893 (N_26893,N_25332,N_25499);
or U26894 (N_26894,N_25102,N_25787);
nand U26895 (N_26895,N_25361,N_25714);
xor U26896 (N_26896,N_25711,N_25589);
nor U26897 (N_26897,N_25203,N_25801);
nor U26898 (N_26898,N_25340,N_25104);
or U26899 (N_26899,N_25358,N_25641);
or U26900 (N_26900,N_25047,N_25897);
nand U26901 (N_26901,N_25472,N_25328);
and U26902 (N_26902,N_25258,N_25988);
xor U26903 (N_26903,N_25315,N_25615);
nand U26904 (N_26904,N_25851,N_25083);
and U26905 (N_26905,N_25561,N_25269);
xnor U26906 (N_26906,N_25738,N_25994);
nor U26907 (N_26907,N_25110,N_25586);
nand U26908 (N_26908,N_25189,N_25028);
and U26909 (N_26909,N_25478,N_25237);
xnor U26910 (N_26910,N_25911,N_25557);
xnor U26911 (N_26911,N_25393,N_25071);
nand U26912 (N_26912,N_25363,N_25795);
xnor U26913 (N_26913,N_25284,N_25539);
nand U26914 (N_26914,N_25169,N_25399);
xor U26915 (N_26915,N_25839,N_25313);
nor U26916 (N_26916,N_25397,N_25191);
nor U26917 (N_26917,N_25153,N_25882);
nor U26918 (N_26918,N_25679,N_25074);
or U26919 (N_26919,N_25933,N_25399);
xnor U26920 (N_26920,N_25116,N_25989);
or U26921 (N_26921,N_25266,N_25443);
or U26922 (N_26922,N_25989,N_25799);
nand U26923 (N_26923,N_25490,N_25427);
nand U26924 (N_26924,N_25085,N_25001);
nor U26925 (N_26925,N_25849,N_25797);
and U26926 (N_26926,N_25092,N_25082);
xnor U26927 (N_26927,N_25855,N_25579);
nor U26928 (N_26928,N_25199,N_25655);
xnor U26929 (N_26929,N_25385,N_25681);
nor U26930 (N_26930,N_25818,N_25361);
or U26931 (N_26931,N_25964,N_25257);
nor U26932 (N_26932,N_25763,N_25133);
and U26933 (N_26933,N_25540,N_25705);
and U26934 (N_26934,N_25576,N_25455);
xnor U26935 (N_26935,N_25639,N_25592);
nand U26936 (N_26936,N_25883,N_25143);
and U26937 (N_26937,N_25407,N_25790);
and U26938 (N_26938,N_25460,N_25933);
or U26939 (N_26939,N_25089,N_25854);
xor U26940 (N_26940,N_25083,N_25736);
nand U26941 (N_26941,N_25690,N_25038);
nor U26942 (N_26942,N_25804,N_25336);
or U26943 (N_26943,N_25712,N_25899);
or U26944 (N_26944,N_25700,N_25634);
and U26945 (N_26945,N_25096,N_25573);
nor U26946 (N_26946,N_25128,N_25730);
or U26947 (N_26947,N_25032,N_25087);
xnor U26948 (N_26948,N_25530,N_25879);
xor U26949 (N_26949,N_25851,N_25784);
or U26950 (N_26950,N_25443,N_25044);
nand U26951 (N_26951,N_25294,N_25089);
and U26952 (N_26952,N_25886,N_25077);
or U26953 (N_26953,N_25094,N_25470);
nor U26954 (N_26954,N_25708,N_25168);
nand U26955 (N_26955,N_25293,N_25706);
or U26956 (N_26956,N_25081,N_25197);
nand U26957 (N_26957,N_25056,N_25264);
nand U26958 (N_26958,N_25623,N_25934);
or U26959 (N_26959,N_25425,N_25280);
nor U26960 (N_26960,N_25591,N_25555);
or U26961 (N_26961,N_25252,N_25705);
xor U26962 (N_26962,N_25633,N_25115);
and U26963 (N_26963,N_25786,N_25621);
nand U26964 (N_26964,N_25540,N_25211);
nand U26965 (N_26965,N_25134,N_25907);
or U26966 (N_26966,N_25299,N_25664);
xnor U26967 (N_26967,N_25945,N_25210);
xor U26968 (N_26968,N_25710,N_25923);
or U26969 (N_26969,N_25631,N_25801);
xor U26970 (N_26970,N_25031,N_25238);
or U26971 (N_26971,N_25372,N_25375);
nand U26972 (N_26972,N_25035,N_25660);
and U26973 (N_26973,N_25197,N_25340);
and U26974 (N_26974,N_25589,N_25618);
xnor U26975 (N_26975,N_25605,N_25646);
or U26976 (N_26976,N_25945,N_25254);
nor U26977 (N_26977,N_25990,N_25303);
nand U26978 (N_26978,N_25800,N_25039);
nand U26979 (N_26979,N_25291,N_25781);
nand U26980 (N_26980,N_25031,N_25767);
nand U26981 (N_26981,N_25960,N_25545);
xnor U26982 (N_26982,N_25358,N_25589);
nand U26983 (N_26983,N_25052,N_25918);
nand U26984 (N_26984,N_25088,N_25463);
and U26985 (N_26985,N_25301,N_25960);
xor U26986 (N_26986,N_25272,N_25842);
or U26987 (N_26987,N_25289,N_25789);
nor U26988 (N_26988,N_25771,N_25207);
and U26989 (N_26989,N_25457,N_25080);
nand U26990 (N_26990,N_25514,N_25823);
nor U26991 (N_26991,N_25247,N_25092);
xor U26992 (N_26992,N_25338,N_25676);
or U26993 (N_26993,N_25016,N_25879);
and U26994 (N_26994,N_25970,N_25360);
or U26995 (N_26995,N_25858,N_25612);
nand U26996 (N_26996,N_25237,N_25397);
nand U26997 (N_26997,N_25748,N_25350);
or U26998 (N_26998,N_25741,N_25237);
and U26999 (N_26999,N_25973,N_25351);
nor U27000 (N_27000,N_26267,N_26630);
xor U27001 (N_27001,N_26305,N_26432);
xnor U27002 (N_27002,N_26521,N_26936);
xor U27003 (N_27003,N_26357,N_26196);
nor U27004 (N_27004,N_26029,N_26700);
nand U27005 (N_27005,N_26637,N_26145);
xor U27006 (N_27006,N_26580,N_26031);
xor U27007 (N_27007,N_26655,N_26034);
nor U27008 (N_27008,N_26293,N_26923);
and U27009 (N_27009,N_26578,N_26807);
nor U27010 (N_27010,N_26524,N_26394);
or U27011 (N_27011,N_26307,N_26174);
xnor U27012 (N_27012,N_26334,N_26484);
xor U27013 (N_27013,N_26072,N_26037);
nand U27014 (N_27014,N_26232,N_26438);
nand U27015 (N_27015,N_26532,N_26822);
nand U27016 (N_27016,N_26440,N_26392);
and U27017 (N_27017,N_26560,N_26974);
xnor U27018 (N_27018,N_26418,N_26523);
and U27019 (N_27019,N_26618,N_26097);
or U27020 (N_27020,N_26405,N_26938);
nand U27021 (N_27021,N_26791,N_26793);
or U27022 (N_27022,N_26841,N_26537);
nor U27023 (N_27023,N_26350,N_26644);
and U27024 (N_27024,N_26699,N_26614);
and U27025 (N_27025,N_26991,N_26879);
nand U27026 (N_27026,N_26850,N_26483);
or U27027 (N_27027,N_26076,N_26608);
nor U27028 (N_27028,N_26672,N_26148);
or U27029 (N_27029,N_26409,N_26878);
xnor U27030 (N_27030,N_26475,N_26961);
or U27031 (N_27031,N_26772,N_26570);
nand U27032 (N_27032,N_26368,N_26309);
and U27033 (N_27033,N_26340,N_26834);
nand U27034 (N_27034,N_26083,N_26898);
and U27035 (N_27035,N_26248,N_26194);
and U27036 (N_27036,N_26000,N_26740);
and U27037 (N_27037,N_26458,N_26369);
and U27038 (N_27038,N_26456,N_26652);
nor U27039 (N_27039,N_26538,N_26103);
or U27040 (N_27040,N_26735,N_26866);
nor U27041 (N_27041,N_26245,N_26055);
xnor U27042 (N_27042,N_26513,N_26059);
xnor U27043 (N_27043,N_26378,N_26612);
nand U27044 (N_27044,N_26292,N_26184);
and U27045 (N_27045,N_26052,N_26909);
and U27046 (N_27046,N_26211,N_26095);
nor U27047 (N_27047,N_26945,N_26497);
and U27048 (N_27048,N_26121,N_26529);
and U27049 (N_27049,N_26075,N_26188);
and U27050 (N_27050,N_26605,N_26453);
xnor U27051 (N_27051,N_26476,N_26415);
nand U27052 (N_27052,N_26178,N_26287);
nor U27053 (N_27053,N_26279,N_26362);
nor U27054 (N_27054,N_26092,N_26761);
xnor U27055 (N_27055,N_26470,N_26645);
and U27056 (N_27056,N_26077,N_26270);
and U27057 (N_27057,N_26955,N_26534);
xor U27058 (N_27058,N_26498,N_26046);
and U27059 (N_27059,N_26199,N_26204);
nor U27060 (N_27060,N_26238,N_26601);
or U27061 (N_27061,N_26796,N_26568);
nor U27062 (N_27062,N_26976,N_26054);
xor U27063 (N_27063,N_26284,N_26774);
nor U27064 (N_27064,N_26242,N_26814);
nand U27065 (N_27065,N_26901,N_26480);
or U27066 (N_27066,N_26230,N_26698);
nor U27067 (N_27067,N_26330,N_26710);
xnor U27068 (N_27068,N_26314,N_26024);
xor U27069 (N_27069,N_26831,N_26530);
xnor U27070 (N_27070,N_26094,N_26897);
nor U27071 (N_27071,N_26039,N_26706);
nor U27072 (N_27072,N_26787,N_26869);
xor U27073 (N_27073,N_26439,N_26249);
nor U27074 (N_27074,N_26262,N_26682);
nand U27075 (N_27075,N_26195,N_26861);
or U27076 (N_27076,N_26753,N_26506);
xor U27077 (N_27077,N_26124,N_26499);
nand U27078 (N_27078,N_26659,N_26624);
or U27079 (N_27079,N_26582,N_26694);
nor U27080 (N_27080,N_26801,N_26301);
xnor U27081 (N_27081,N_26719,N_26143);
nand U27082 (N_27082,N_26149,N_26776);
xnor U27083 (N_27083,N_26466,N_26220);
and U27084 (N_27084,N_26020,N_26080);
and U27085 (N_27085,N_26893,N_26079);
or U27086 (N_27086,N_26353,N_26692);
nand U27087 (N_27087,N_26808,N_26565);
xor U27088 (N_27088,N_26584,N_26541);
and U27089 (N_27089,N_26328,N_26531);
nor U27090 (N_27090,N_26452,N_26864);
nand U27091 (N_27091,N_26918,N_26952);
xnor U27092 (N_27092,N_26583,N_26345);
or U27093 (N_27093,N_26297,N_26332);
or U27094 (N_27094,N_26826,N_26844);
nand U27095 (N_27095,N_26109,N_26561);
and U27096 (N_27096,N_26081,N_26727);
nand U27097 (N_27097,N_26004,N_26957);
xor U27098 (N_27098,N_26329,N_26997);
nand U27099 (N_27099,N_26900,N_26283);
nor U27100 (N_27100,N_26315,N_26090);
or U27101 (N_27101,N_26554,N_26701);
and U27102 (N_27102,N_26001,N_26402);
or U27103 (N_27103,N_26794,N_26854);
and U27104 (N_27104,N_26414,N_26713);
and U27105 (N_27105,N_26060,N_26091);
nor U27106 (N_27106,N_26073,N_26413);
nor U27107 (N_27107,N_26326,N_26216);
and U27108 (N_27108,N_26300,N_26349);
xnor U27109 (N_27109,N_26503,N_26653);
or U27110 (N_27110,N_26087,N_26880);
xnor U27111 (N_27111,N_26858,N_26697);
and U27112 (N_27112,N_26009,N_26832);
and U27113 (N_27113,N_26425,N_26535);
and U27114 (N_27114,N_26755,N_26299);
or U27115 (N_27115,N_26022,N_26112);
and U27116 (N_27116,N_26189,N_26745);
nand U27117 (N_27117,N_26343,N_26288);
xnor U27118 (N_27118,N_26750,N_26639);
and U27119 (N_27119,N_26904,N_26254);
nand U27120 (N_27120,N_26712,N_26346);
xor U27121 (N_27121,N_26258,N_26014);
xor U27122 (N_27122,N_26200,N_26275);
and U27123 (N_27123,N_26295,N_26224);
and U27124 (N_27124,N_26686,N_26434);
or U27125 (N_27125,N_26208,N_26114);
or U27126 (N_27126,N_26627,N_26044);
nor U27127 (N_27127,N_26606,N_26367);
xnor U27128 (N_27128,N_26871,N_26975);
nand U27129 (N_27129,N_26210,N_26212);
xor U27130 (N_27130,N_26252,N_26572);
nor U27131 (N_27131,N_26983,N_26151);
nand U27132 (N_27132,N_26795,N_26587);
or U27133 (N_27133,N_26322,N_26320);
xor U27134 (N_27134,N_26430,N_26967);
nand U27135 (N_27135,N_26388,N_26839);
and U27136 (N_27136,N_26058,N_26882);
nand U27137 (N_27137,N_26276,N_26168);
nand U27138 (N_27138,N_26336,N_26985);
xnor U27139 (N_27139,N_26744,N_26240);
nor U27140 (N_27140,N_26585,N_26549);
nand U27141 (N_27141,N_26335,N_26280);
nor U27142 (N_27142,N_26355,N_26131);
nor U27143 (N_27143,N_26954,N_26061);
nand U27144 (N_27144,N_26469,N_26633);
or U27145 (N_27145,N_26036,N_26045);
nand U27146 (N_27146,N_26323,N_26217);
or U27147 (N_27147,N_26333,N_26960);
and U27148 (N_27148,N_26908,N_26681);
xnor U27149 (N_27149,N_26944,N_26389);
nor U27150 (N_27150,N_26198,N_26948);
nor U27151 (N_27151,N_26514,N_26100);
or U27152 (N_27152,N_26781,N_26972);
or U27153 (N_27153,N_26290,N_26312);
nor U27154 (N_27154,N_26096,N_26166);
nand U27155 (N_27155,N_26445,N_26939);
or U27156 (N_27156,N_26576,N_26684);
and U27157 (N_27157,N_26610,N_26730);
or U27158 (N_27158,N_26851,N_26819);
nor U27159 (N_27159,N_26116,N_26631);
or U27160 (N_27160,N_26107,N_26797);
or U27161 (N_27161,N_26958,N_26071);
or U27162 (N_27162,N_26435,N_26613);
and U27163 (N_27163,N_26640,N_26370);
nor U27164 (N_27164,N_26015,N_26696);
or U27165 (N_27165,N_26042,N_26830);
or U27166 (N_27166,N_26722,N_26743);
or U27167 (N_27167,N_26751,N_26454);
nand U27168 (N_27168,N_26959,N_26737);
xor U27169 (N_27169,N_26708,N_26899);
and U27170 (N_27170,N_26995,N_26520);
xor U27171 (N_27171,N_26665,N_26347);
or U27172 (N_27172,N_26442,N_26175);
nor U27173 (N_27173,N_26494,N_26308);
and U27174 (N_27174,N_26542,N_26725);
nand U27175 (N_27175,N_26790,N_26703);
or U27176 (N_27176,N_26956,N_26410);
and U27177 (N_27177,N_26126,N_26051);
nand U27178 (N_27178,N_26233,N_26845);
or U27179 (N_27179,N_26950,N_26688);
xor U27180 (N_27180,N_26050,N_26236);
and U27181 (N_27181,N_26374,N_26888);
nand U27182 (N_27182,N_26611,N_26543);
nor U27183 (N_27183,N_26342,N_26732);
or U27184 (N_27184,N_26815,N_26496);
nand U27185 (N_27185,N_26176,N_26734);
nand U27186 (N_27186,N_26657,N_26012);
and U27187 (N_27187,N_26666,N_26433);
xor U27188 (N_27188,N_26085,N_26816);
xor U27189 (N_27189,N_26250,N_26495);
nand U27190 (N_27190,N_26462,N_26979);
or U27191 (N_27191,N_26931,N_26467);
and U27192 (N_27192,N_26827,N_26406);
or U27193 (N_27193,N_26846,N_26241);
xnor U27194 (N_27194,N_26182,N_26843);
and U27195 (N_27195,N_26172,N_26662);
nand U27196 (N_27196,N_26978,N_26677);
nand U27197 (N_27197,N_26987,N_26487);
nor U27198 (N_27198,N_26482,N_26977);
or U27199 (N_27199,N_26912,N_26747);
nand U27200 (N_27200,N_26853,N_26920);
xnor U27201 (N_27201,N_26273,N_26206);
and U27202 (N_27202,N_26449,N_26226);
and U27203 (N_27203,N_26567,N_26999);
nand U27204 (N_27204,N_26768,N_26461);
nand U27205 (N_27205,N_26748,N_26836);
nand U27206 (N_27206,N_26375,N_26835);
or U27207 (N_27207,N_26491,N_26229);
or U27208 (N_27208,N_26949,N_26400);
or U27209 (N_27209,N_26234,N_26988);
xnor U27210 (N_27210,N_26393,N_26180);
and U27211 (N_27211,N_26030,N_26792);
xor U27212 (N_27212,N_26604,N_26770);
or U27213 (N_27213,N_26274,N_26887);
and U27214 (N_27214,N_26237,N_26401);
or U27215 (N_27215,N_26186,N_26398);
xor U27216 (N_27216,N_26886,N_26255);
nand U27217 (N_27217,N_26619,N_26767);
or U27218 (N_27218,N_26152,N_26005);
and U27219 (N_27219,N_26313,N_26946);
xor U27220 (N_27220,N_26916,N_26579);
nor U27221 (N_27221,N_26327,N_26870);
xor U27222 (N_27222,N_26381,N_26099);
or U27223 (N_27223,N_26577,N_26215);
and U27224 (N_27224,N_26306,N_26629);
xnor U27225 (N_27225,N_26765,N_26132);
xor U27226 (N_27226,N_26875,N_26154);
nand U27227 (N_27227,N_26522,N_26364);
nand U27228 (N_27228,N_26218,N_26857);
nand U27229 (N_27229,N_26125,N_26019);
and U27230 (N_27230,N_26086,N_26294);
nand U27231 (N_27231,N_26661,N_26980);
xor U27232 (N_27232,N_26557,N_26160);
nand U27233 (N_27233,N_26511,N_26408);
xor U27234 (N_27234,N_26041,N_26926);
and U27235 (N_27235,N_26028,N_26225);
nand U27236 (N_27236,N_26481,N_26894);
or U27237 (N_27237,N_26507,N_26164);
or U27238 (N_27238,N_26011,N_26066);
or U27239 (N_27239,N_26360,N_26108);
xnor U27240 (N_27240,N_26338,N_26444);
or U27241 (N_27241,N_26563,N_26070);
or U27242 (N_27242,N_26986,N_26764);
and U27243 (N_27243,N_26399,N_26352);
nand U27244 (N_27244,N_26914,N_26032);
and U27245 (N_27245,N_26865,N_26508);
nand U27246 (N_27246,N_26915,N_26463);
and U27247 (N_27247,N_26104,N_26113);
xor U27248 (N_27248,N_26187,N_26040);
and U27249 (N_27249,N_26785,N_26302);
nand U27250 (N_27250,N_26473,N_26318);
or U27251 (N_27251,N_26896,N_26754);
xor U27252 (N_27252,N_26924,N_26246);
nand U27253 (N_27253,N_26884,N_26358);
and U27254 (N_27254,N_26155,N_26356);
xnor U27255 (N_27255,N_26033,N_26634);
nand U27256 (N_27256,N_26500,N_26192);
nor U27257 (N_27257,N_26384,N_26996);
or U27258 (N_27258,N_26856,N_26726);
nand U27259 (N_27259,N_26859,N_26123);
xnor U27260 (N_27260,N_26840,N_26376);
and U27261 (N_27261,N_26990,N_26065);
nand U27262 (N_27262,N_26063,N_26266);
nand U27263 (N_27263,N_26197,N_26025);
nand U27264 (N_27264,N_26942,N_26902);
xnor U27265 (N_27265,N_26622,N_26419);
or U27266 (N_27266,N_26680,N_26027);
and U27267 (N_27267,N_26729,N_26150);
xor U27268 (N_27268,N_26739,N_26472);
nor U27269 (N_27269,N_26371,N_26253);
xor U27270 (N_27270,N_26526,N_26239);
xnor U27271 (N_27271,N_26365,N_26800);
nor U27272 (N_27272,N_26695,N_26867);
or U27273 (N_27273,N_26407,N_26319);
nand U27274 (N_27274,N_26423,N_26304);
and U27275 (N_27275,N_26922,N_26474);
and U27276 (N_27276,N_26047,N_26115);
nand U27277 (N_27277,N_26023,N_26420);
nor U27278 (N_27278,N_26510,N_26251);
and U27279 (N_27279,N_26105,N_26581);
or U27280 (N_27280,N_26903,N_26465);
nand U27281 (N_27281,N_26286,N_26679);
nor U27282 (N_27282,N_26228,N_26013);
nand U27283 (N_27283,N_26264,N_26282);
and U27284 (N_27284,N_26518,N_26683);
or U27285 (N_27285,N_26501,N_26436);
or U27286 (N_27286,N_26147,N_26517);
nand U27287 (N_27287,N_26933,N_26678);
nor U27288 (N_27288,N_26404,N_26782);
nor U27289 (N_27289,N_26426,N_26907);
or U27290 (N_27290,N_26962,N_26354);
or U27291 (N_27291,N_26341,N_26642);
nand U27292 (N_27292,N_26177,N_26925);
nor U27293 (N_27293,N_26895,N_26162);
and U27294 (N_27294,N_26704,N_26139);
or U27295 (N_27295,N_26707,N_26167);
nand U27296 (N_27296,N_26303,N_26209);
nand U27297 (N_27297,N_26431,N_26421);
xor U27298 (N_27298,N_26675,N_26820);
nand U27299 (N_27299,N_26589,N_26257);
and U27300 (N_27300,N_26635,N_26868);
nand U27301 (N_27301,N_26658,N_26648);
xnor U27302 (N_27302,N_26890,N_26008);
nand U27303 (N_27303,N_26599,N_26311);
nand U27304 (N_27304,N_26715,N_26968);
nor U27305 (N_27305,N_26057,N_26982);
nand U27306 (N_27306,N_26069,N_26053);
nor U27307 (N_27307,N_26366,N_26883);
and U27308 (N_27308,N_26847,N_26855);
nand U27309 (N_27309,N_26396,N_26447);
nor U27310 (N_27310,N_26163,N_26161);
xor U27311 (N_27311,N_26746,N_26574);
nand U27312 (N_27312,N_26459,N_26383);
or U27313 (N_27313,N_26016,N_26395);
nand U27314 (N_27314,N_26120,N_26263);
or U27315 (N_27315,N_26324,N_26935);
or U27316 (N_27316,N_26766,N_26272);
or U27317 (N_27317,N_26590,N_26930);
or U27318 (N_27318,N_26762,N_26636);
nor U27319 (N_27319,N_26504,N_26718);
or U27320 (N_27320,N_26992,N_26667);
or U27321 (N_27321,N_26736,N_26351);
or U27322 (N_27322,N_26673,N_26664);
nand U27323 (N_27323,N_26268,N_26603);
and U27324 (N_27324,N_26779,N_26823);
or U27325 (N_27325,N_26359,N_26687);
nand U27326 (N_27326,N_26643,N_26488);
xor U27327 (N_27327,N_26848,N_26716);
nor U27328 (N_27328,N_26026,N_26321);
nand U27329 (N_27329,N_26752,N_26674);
xor U27330 (N_27330,N_26153,N_26628);
nand U27331 (N_27331,N_26783,N_26377);
xor U27332 (N_27332,N_26721,N_26539);
nand U27333 (N_27333,N_26490,N_26049);
and U27334 (N_27334,N_26965,N_26102);
nand U27335 (N_27335,N_26331,N_26221);
nand U27336 (N_27336,N_26759,N_26201);
nor U27337 (N_27337,N_26205,N_26141);
and U27338 (N_27338,N_26758,N_26993);
or U27339 (N_27339,N_26852,N_26600);
nor U27340 (N_27340,N_26111,N_26428);
or U27341 (N_27341,N_26806,N_26285);
nor U27342 (N_27342,N_26862,N_26344);
xnor U27343 (N_27343,N_26575,N_26422);
and U27344 (N_27344,N_26705,N_26810);
or U27345 (N_27345,N_26670,N_26390);
or U27346 (N_27346,N_26382,N_26068);
nor U27347 (N_27347,N_26728,N_26825);
nand U27348 (N_27348,N_26158,N_26966);
and U27349 (N_27349,N_26243,N_26720);
and U27350 (N_27350,N_26760,N_26873);
and U27351 (N_27351,N_26559,N_26512);
or U27352 (N_27352,N_26742,N_26119);
or U27353 (N_27353,N_26138,N_26615);
nor U27354 (N_27354,N_26919,N_26464);
xor U27355 (N_27355,N_26555,N_26235);
xnor U27356 (N_27356,N_26062,N_26802);
nor U27357 (N_27357,N_26289,N_26676);
nand U27358 (N_27358,N_26872,N_26165);
xnor U27359 (N_27359,N_26485,N_26159);
nand U27360 (N_27360,N_26460,N_26714);
nand U27361 (N_27361,N_26117,N_26892);
nor U27362 (N_27362,N_26078,N_26553);
nor U27363 (N_27363,N_26573,N_26717);
nand U27364 (N_27364,N_26593,N_26821);
nand U27365 (N_27365,N_26056,N_26828);
xor U27366 (N_27366,N_26777,N_26649);
and U27367 (N_27367,N_26185,N_26773);
nand U27368 (N_27368,N_26527,N_26778);
or U27369 (N_27369,N_26809,N_26741);
and U27370 (N_27370,N_26617,N_26571);
or U27371 (N_27371,N_26876,N_26118);
or U27372 (N_27372,N_26064,N_26550);
nor U27373 (N_27373,N_26891,N_26877);
and U27374 (N_27374,N_26951,N_26799);
nor U27375 (N_27375,N_26265,N_26397);
and U27376 (N_27376,N_26609,N_26906);
nor U27377 (N_27377,N_26446,N_26455);
and U27378 (N_27378,N_26492,N_26231);
or U27379 (N_27379,N_26525,N_26937);
and U27380 (N_27380,N_26805,N_26595);
xnor U27381 (N_27381,N_26971,N_26271);
and U27382 (N_27382,N_26690,N_26849);
xnor U27383 (N_27383,N_26203,N_26157);
and U27384 (N_27384,N_26784,N_26566);
nor U27385 (N_27385,N_26838,N_26973);
nor U27386 (N_27386,N_26339,N_26219);
nor U27387 (N_27387,N_26602,N_26963);
xnor U27388 (N_27388,N_26417,N_26786);
nand U27389 (N_27389,N_26010,N_26913);
and U27390 (N_27390,N_26372,N_26989);
nand U27391 (N_27391,N_26552,N_26947);
nand U27392 (N_27392,N_26547,N_26917);
nand U27393 (N_27393,N_26656,N_26693);
and U27394 (N_27394,N_26711,N_26214);
and U27395 (N_27395,N_26471,N_26556);
and U27396 (N_27396,N_26911,N_26486);
nor U27397 (N_27397,N_26098,N_26144);
and U27398 (N_27398,N_26457,N_26142);
nand U27399 (N_27399,N_26756,N_26509);
and U27400 (N_27400,N_26544,N_26190);
xor U27401 (N_27401,N_26594,N_26591);
and U27402 (N_27402,N_26860,N_26934);
or U27403 (N_27403,N_26932,N_26540);
nand U27404 (N_27404,N_26626,N_26493);
xnor U27405 (N_27405,N_26137,N_26478);
nand U27406 (N_27406,N_26207,N_26837);
xor U27407 (N_27407,N_26450,N_26881);
nor U27408 (N_27408,N_26516,N_26607);
or U27409 (N_27409,N_26548,N_26502);
or U27410 (N_27410,N_26183,N_26437);
nand U27411 (N_27411,N_26889,N_26179);
nor U27412 (N_27412,N_26003,N_26261);
nand U27413 (N_27413,N_26632,N_26489);
nand U27414 (N_27414,N_26416,N_26448);
or U27415 (N_27415,N_26998,N_26135);
and U27416 (N_27416,N_26002,N_26278);
nand U27417 (N_27417,N_26256,N_26733);
or U27418 (N_27418,N_26337,N_26325);
nor U27419 (N_27419,N_26647,N_26110);
or U27420 (N_27420,N_26620,N_26101);
nor U27421 (N_27421,N_26874,N_26953);
or U27422 (N_27422,N_26021,N_26702);
nor U27423 (N_27423,N_26411,N_26477);
xnor U27424 (N_27424,N_26363,N_26441);
nand U27425 (N_27425,N_26043,N_26621);
nor U27426 (N_27426,N_26597,N_26391);
xnor U27427 (N_27427,N_26586,N_26412);
and U27428 (N_27428,N_26663,N_26505);
or U27429 (N_27429,N_26074,N_26775);
and U27430 (N_27430,N_26387,N_26905);
and U27431 (N_27431,N_26093,N_26385);
and U27432 (N_27432,N_26863,N_26173);
xnor U27433 (N_27433,N_26723,N_26451);
nor U27434 (N_27434,N_26193,N_26269);
and U27435 (N_27435,N_26928,N_26646);
nand U27436 (N_27436,N_26929,N_26106);
nand U27437 (N_27437,N_26921,N_26519);
nand U27438 (N_27438,N_26943,N_26833);
nand U27439 (N_27439,N_26569,N_26803);
and U27440 (N_27440,N_26038,N_26545);
or U27441 (N_27441,N_26592,N_26386);
nand U27442 (N_27442,N_26804,N_26088);
nor U27443 (N_27443,N_26048,N_26317);
and U27444 (N_27444,N_26244,N_26169);
and U27445 (N_27445,N_26616,N_26479);
xor U27446 (N_27446,N_26780,N_26927);
xor U27447 (N_27447,N_26136,N_26316);
nor U27448 (N_27448,N_26361,N_26650);
nor U27449 (N_27449,N_26006,N_26994);
or U27450 (N_27450,N_26171,N_26981);
xnor U27451 (N_27451,N_26533,N_26724);
or U27452 (N_27452,N_26140,N_26130);
and U27453 (N_27453,N_26007,N_26625);
nor U27454 (N_27454,N_26379,N_26082);
xor U27455 (N_27455,N_26018,N_26281);
nand U27456 (N_27456,N_26651,N_26310);
xor U27457 (N_27457,N_26984,N_26146);
nand U27458 (N_27458,N_26181,N_26035);
nor U27459 (N_27459,N_26223,N_26660);
nand U27460 (N_27460,N_26222,N_26156);
nor U27461 (N_27461,N_26769,N_26528);
xor U27462 (N_27462,N_26813,N_26403);
nor U27463 (N_27463,N_26668,N_26424);
nand U27464 (N_27464,N_26551,N_26964);
xnor U27465 (N_27465,N_26443,N_26170);
nand U27466 (N_27466,N_26817,N_26691);
or U27467 (N_27467,N_26129,N_26468);
nand U27468 (N_27468,N_26685,N_26824);
nor U27469 (N_27469,N_26128,N_26564);
nand U27470 (N_27470,N_26812,N_26067);
and U27471 (N_27471,N_26134,N_26298);
nand U27472 (N_27472,N_26277,N_26731);
nor U27473 (N_27473,N_26191,N_26738);
or U27474 (N_27474,N_26709,N_26940);
xor U27475 (N_27475,N_26789,N_26122);
or U27476 (N_27476,N_26127,N_26885);
nand U27477 (N_27477,N_26515,N_26757);
xor U27478 (N_27478,N_26818,N_26588);
and U27479 (N_27479,N_26348,N_26829);
nand U27480 (N_27480,N_26133,N_26910);
or U27481 (N_27481,N_26291,N_26641);
and U27482 (N_27482,N_26596,N_26260);
xnor U27483 (N_27483,N_26798,N_26671);
nand U27484 (N_27484,N_26623,N_26562);
nand U27485 (N_27485,N_26380,N_26558);
nand U27486 (N_27486,N_26969,N_26763);
or U27487 (N_27487,N_26689,N_26373);
xor U27488 (N_27488,N_26788,N_26202);
nor U27489 (N_27489,N_26811,N_26941);
nand U27490 (N_27490,N_26427,N_26017);
xor U27491 (N_27491,N_26247,N_26084);
and U27492 (N_27492,N_26598,N_26429);
nand U27493 (N_27493,N_26771,N_26749);
or U27494 (N_27494,N_26970,N_26546);
nand U27495 (N_27495,N_26638,N_26669);
or U27496 (N_27496,N_26089,N_26296);
and U27497 (N_27497,N_26213,N_26227);
and U27498 (N_27498,N_26259,N_26536);
nor U27499 (N_27499,N_26842,N_26654);
or U27500 (N_27500,N_26059,N_26822);
and U27501 (N_27501,N_26852,N_26571);
nand U27502 (N_27502,N_26851,N_26089);
nor U27503 (N_27503,N_26419,N_26258);
or U27504 (N_27504,N_26752,N_26430);
or U27505 (N_27505,N_26450,N_26222);
xor U27506 (N_27506,N_26387,N_26239);
xnor U27507 (N_27507,N_26054,N_26956);
and U27508 (N_27508,N_26136,N_26275);
or U27509 (N_27509,N_26845,N_26443);
nand U27510 (N_27510,N_26691,N_26322);
nor U27511 (N_27511,N_26284,N_26868);
nand U27512 (N_27512,N_26257,N_26937);
and U27513 (N_27513,N_26681,N_26742);
or U27514 (N_27514,N_26053,N_26978);
nand U27515 (N_27515,N_26925,N_26567);
nand U27516 (N_27516,N_26289,N_26635);
or U27517 (N_27517,N_26265,N_26610);
nor U27518 (N_27518,N_26135,N_26727);
nor U27519 (N_27519,N_26226,N_26420);
and U27520 (N_27520,N_26763,N_26582);
nor U27521 (N_27521,N_26616,N_26245);
nand U27522 (N_27522,N_26403,N_26274);
or U27523 (N_27523,N_26560,N_26420);
nand U27524 (N_27524,N_26442,N_26313);
nand U27525 (N_27525,N_26721,N_26480);
and U27526 (N_27526,N_26703,N_26289);
xor U27527 (N_27527,N_26127,N_26433);
nor U27528 (N_27528,N_26399,N_26114);
or U27529 (N_27529,N_26080,N_26857);
and U27530 (N_27530,N_26643,N_26493);
xnor U27531 (N_27531,N_26422,N_26547);
nand U27532 (N_27532,N_26054,N_26485);
or U27533 (N_27533,N_26579,N_26862);
and U27534 (N_27534,N_26659,N_26440);
or U27535 (N_27535,N_26239,N_26786);
xnor U27536 (N_27536,N_26811,N_26592);
or U27537 (N_27537,N_26452,N_26487);
nand U27538 (N_27538,N_26562,N_26760);
nor U27539 (N_27539,N_26798,N_26992);
nand U27540 (N_27540,N_26511,N_26947);
nor U27541 (N_27541,N_26551,N_26136);
nand U27542 (N_27542,N_26030,N_26274);
and U27543 (N_27543,N_26386,N_26863);
nand U27544 (N_27544,N_26126,N_26498);
or U27545 (N_27545,N_26033,N_26344);
and U27546 (N_27546,N_26190,N_26629);
nand U27547 (N_27547,N_26260,N_26558);
or U27548 (N_27548,N_26997,N_26745);
nand U27549 (N_27549,N_26132,N_26290);
nor U27550 (N_27550,N_26061,N_26100);
nor U27551 (N_27551,N_26036,N_26586);
nor U27552 (N_27552,N_26483,N_26816);
nor U27553 (N_27553,N_26194,N_26455);
nand U27554 (N_27554,N_26544,N_26001);
or U27555 (N_27555,N_26855,N_26297);
xor U27556 (N_27556,N_26923,N_26549);
xor U27557 (N_27557,N_26844,N_26939);
nand U27558 (N_27558,N_26204,N_26485);
and U27559 (N_27559,N_26859,N_26710);
nor U27560 (N_27560,N_26007,N_26768);
and U27561 (N_27561,N_26280,N_26664);
and U27562 (N_27562,N_26266,N_26840);
or U27563 (N_27563,N_26521,N_26645);
and U27564 (N_27564,N_26940,N_26639);
nand U27565 (N_27565,N_26673,N_26761);
and U27566 (N_27566,N_26852,N_26836);
and U27567 (N_27567,N_26599,N_26526);
nor U27568 (N_27568,N_26547,N_26003);
nor U27569 (N_27569,N_26161,N_26841);
nor U27570 (N_27570,N_26278,N_26822);
xor U27571 (N_27571,N_26141,N_26157);
or U27572 (N_27572,N_26727,N_26773);
nand U27573 (N_27573,N_26282,N_26951);
or U27574 (N_27574,N_26552,N_26263);
nor U27575 (N_27575,N_26131,N_26861);
nand U27576 (N_27576,N_26472,N_26692);
xnor U27577 (N_27577,N_26506,N_26636);
xor U27578 (N_27578,N_26174,N_26634);
xnor U27579 (N_27579,N_26696,N_26224);
and U27580 (N_27580,N_26286,N_26248);
and U27581 (N_27581,N_26774,N_26589);
nand U27582 (N_27582,N_26263,N_26727);
nand U27583 (N_27583,N_26275,N_26644);
nand U27584 (N_27584,N_26589,N_26445);
nor U27585 (N_27585,N_26144,N_26419);
or U27586 (N_27586,N_26587,N_26988);
xnor U27587 (N_27587,N_26783,N_26677);
nand U27588 (N_27588,N_26941,N_26778);
or U27589 (N_27589,N_26455,N_26916);
nand U27590 (N_27590,N_26186,N_26482);
and U27591 (N_27591,N_26592,N_26548);
nor U27592 (N_27592,N_26552,N_26825);
or U27593 (N_27593,N_26544,N_26239);
and U27594 (N_27594,N_26464,N_26402);
nand U27595 (N_27595,N_26450,N_26021);
nor U27596 (N_27596,N_26163,N_26721);
or U27597 (N_27597,N_26740,N_26622);
and U27598 (N_27598,N_26498,N_26010);
or U27599 (N_27599,N_26091,N_26046);
nor U27600 (N_27600,N_26886,N_26374);
or U27601 (N_27601,N_26880,N_26303);
or U27602 (N_27602,N_26149,N_26569);
nor U27603 (N_27603,N_26405,N_26698);
nor U27604 (N_27604,N_26302,N_26512);
and U27605 (N_27605,N_26047,N_26167);
or U27606 (N_27606,N_26681,N_26202);
nor U27607 (N_27607,N_26894,N_26599);
nor U27608 (N_27608,N_26888,N_26174);
or U27609 (N_27609,N_26525,N_26829);
nand U27610 (N_27610,N_26122,N_26806);
nand U27611 (N_27611,N_26408,N_26454);
xor U27612 (N_27612,N_26302,N_26905);
or U27613 (N_27613,N_26234,N_26700);
and U27614 (N_27614,N_26047,N_26518);
nand U27615 (N_27615,N_26212,N_26341);
xnor U27616 (N_27616,N_26297,N_26635);
nand U27617 (N_27617,N_26690,N_26036);
nor U27618 (N_27618,N_26013,N_26299);
or U27619 (N_27619,N_26550,N_26375);
nor U27620 (N_27620,N_26330,N_26385);
and U27621 (N_27621,N_26217,N_26815);
or U27622 (N_27622,N_26773,N_26292);
and U27623 (N_27623,N_26259,N_26730);
nor U27624 (N_27624,N_26859,N_26582);
or U27625 (N_27625,N_26994,N_26737);
and U27626 (N_27626,N_26128,N_26911);
nand U27627 (N_27627,N_26855,N_26903);
and U27628 (N_27628,N_26117,N_26692);
and U27629 (N_27629,N_26463,N_26166);
xnor U27630 (N_27630,N_26509,N_26045);
and U27631 (N_27631,N_26243,N_26618);
nor U27632 (N_27632,N_26503,N_26479);
xnor U27633 (N_27633,N_26229,N_26635);
nand U27634 (N_27634,N_26629,N_26426);
and U27635 (N_27635,N_26245,N_26464);
xor U27636 (N_27636,N_26855,N_26342);
nor U27637 (N_27637,N_26373,N_26862);
or U27638 (N_27638,N_26899,N_26990);
nor U27639 (N_27639,N_26224,N_26317);
nand U27640 (N_27640,N_26699,N_26903);
xnor U27641 (N_27641,N_26026,N_26711);
and U27642 (N_27642,N_26521,N_26418);
and U27643 (N_27643,N_26370,N_26538);
xor U27644 (N_27644,N_26282,N_26758);
nor U27645 (N_27645,N_26266,N_26860);
or U27646 (N_27646,N_26955,N_26543);
or U27647 (N_27647,N_26629,N_26054);
nor U27648 (N_27648,N_26511,N_26736);
nand U27649 (N_27649,N_26119,N_26468);
nand U27650 (N_27650,N_26940,N_26271);
xnor U27651 (N_27651,N_26675,N_26718);
xor U27652 (N_27652,N_26339,N_26568);
xnor U27653 (N_27653,N_26983,N_26265);
and U27654 (N_27654,N_26336,N_26331);
or U27655 (N_27655,N_26465,N_26104);
nor U27656 (N_27656,N_26482,N_26014);
or U27657 (N_27657,N_26087,N_26105);
nor U27658 (N_27658,N_26108,N_26082);
xor U27659 (N_27659,N_26287,N_26227);
or U27660 (N_27660,N_26749,N_26428);
and U27661 (N_27661,N_26607,N_26871);
nand U27662 (N_27662,N_26181,N_26768);
or U27663 (N_27663,N_26693,N_26883);
and U27664 (N_27664,N_26996,N_26000);
and U27665 (N_27665,N_26636,N_26927);
nor U27666 (N_27666,N_26628,N_26112);
and U27667 (N_27667,N_26974,N_26064);
and U27668 (N_27668,N_26403,N_26769);
or U27669 (N_27669,N_26455,N_26521);
or U27670 (N_27670,N_26221,N_26363);
or U27671 (N_27671,N_26788,N_26368);
xor U27672 (N_27672,N_26012,N_26263);
and U27673 (N_27673,N_26694,N_26576);
or U27674 (N_27674,N_26185,N_26911);
and U27675 (N_27675,N_26406,N_26127);
or U27676 (N_27676,N_26683,N_26417);
and U27677 (N_27677,N_26689,N_26739);
and U27678 (N_27678,N_26209,N_26449);
nor U27679 (N_27679,N_26639,N_26848);
and U27680 (N_27680,N_26250,N_26802);
and U27681 (N_27681,N_26623,N_26038);
and U27682 (N_27682,N_26788,N_26491);
and U27683 (N_27683,N_26778,N_26960);
nand U27684 (N_27684,N_26174,N_26331);
and U27685 (N_27685,N_26829,N_26544);
nor U27686 (N_27686,N_26685,N_26028);
nand U27687 (N_27687,N_26573,N_26460);
or U27688 (N_27688,N_26413,N_26733);
and U27689 (N_27689,N_26783,N_26780);
or U27690 (N_27690,N_26369,N_26478);
and U27691 (N_27691,N_26781,N_26195);
or U27692 (N_27692,N_26244,N_26482);
nor U27693 (N_27693,N_26231,N_26350);
or U27694 (N_27694,N_26150,N_26234);
nand U27695 (N_27695,N_26385,N_26271);
nand U27696 (N_27696,N_26681,N_26602);
nor U27697 (N_27697,N_26348,N_26572);
or U27698 (N_27698,N_26717,N_26221);
and U27699 (N_27699,N_26154,N_26153);
nand U27700 (N_27700,N_26509,N_26230);
or U27701 (N_27701,N_26868,N_26398);
xnor U27702 (N_27702,N_26360,N_26953);
xor U27703 (N_27703,N_26297,N_26583);
nand U27704 (N_27704,N_26912,N_26299);
and U27705 (N_27705,N_26746,N_26826);
xnor U27706 (N_27706,N_26195,N_26048);
nor U27707 (N_27707,N_26384,N_26103);
nand U27708 (N_27708,N_26243,N_26166);
and U27709 (N_27709,N_26314,N_26101);
xor U27710 (N_27710,N_26145,N_26505);
nor U27711 (N_27711,N_26134,N_26297);
and U27712 (N_27712,N_26841,N_26281);
or U27713 (N_27713,N_26991,N_26472);
and U27714 (N_27714,N_26263,N_26966);
nor U27715 (N_27715,N_26483,N_26995);
nand U27716 (N_27716,N_26476,N_26044);
xnor U27717 (N_27717,N_26554,N_26086);
nor U27718 (N_27718,N_26992,N_26491);
nand U27719 (N_27719,N_26134,N_26252);
or U27720 (N_27720,N_26870,N_26322);
and U27721 (N_27721,N_26664,N_26250);
and U27722 (N_27722,N_26007,N_26172);
nor U27723 (N_27723,N_26475,N_26027);
and U27724 (N_27724,N_26288,N_26415);
or U27725 (N_27725,N_26442,N_26674);
and U27726 (N_27726,N_26400,N_26723);
nor U27727 (N_27727,N_26564,N_26654);
or U27728 (N_27728,N_26143,N_26489);
and U27729 (N_27729,N_26036,N_26105);
xor U27730 (N_27730,N_26096,N_26810);
xnor U27731 (N_27731,N_26509,N_26331);
nor U27732 (N_27732,N_26308,N_26574);
and U27733 (N_27733,N_26571,N_26077);
nand U27734 (N_27734,N_26866,N_26569);
nor U27735 (N_27735,N_26478,N_26442);
nand U27736 (N_27736,N_26460,N_26626);
xor U27737 (N_27737,N_26661,N_26935);
nor U27738 (N_27738,N_26567,N_26742);
nand U27739 (N_27739,N_26176,N_26872);
and U27740 (N_27740,N_26297,N_26149);
nor U27741 (N_27741,N_26160,N_26991);
xor U27742 (N_27742,N_26697,N_26881);
xnor U27743 (N_27743,N_26683,N_26835);
and U27744 (N_27744,N_26116,N_26645);
nor U27745 (N_27745,N_26251,N_26515);
and U27746 (N_27746,N_26463,N_26608);
nor U27747 (N_27747,N_26682,N_26261);
or U27748 (N_27748,N_26142,N_26095);
and U27749 (N_27749,N_26600,N_26737);
xnor U27750 (N_27750,N_26864,N_26993);
or U27751 (N_27751,N_26140,N_26611);
xor U27752 (N_27752,N_26083,N_26643);
and U27753 (N_27753,N_26334,N_26335);
and U27754 (N_27754,N_26159,N_26400);
nor U27755 (N_27755,N_26968,N_26582);
nor U27756 (N_27756,N_26873,N_26590);
xor U27757 (N_27757,N_26992,N_26539);
and U27758 (N_27758,N_26307,N_26992);
nand U27759 (N_27759,N_26181,N_26860);
or U27760 (N_27760,N_26471,N_26504);
xnor U27761 (N_27761,N_26263,N_26155);
or U27762 (N_27762,N_26436,N_26424);
nor U27763 (N_27763,N_26218,N_26685);
and U27764 (N_27764,N_26227,N_26489);
and U27765 (N_27765,N_26418,N_26590);
nand U27766 (N_27766,N_26172,N_26500);
nand U27767 (N_27767,N_26452,N_26581);
and U27768 (N_27768,N_26084,N_26879);
nand U27769 (N_27769,N_26195,N_26455);
and U27770 (N_27770,N_26707,N_26008);
and U27771 (N_27771,N_26883,N_26586);
or U27772 (N_27772,N_26464,N_26818);
nand U27773 (N_27773,N_26375,N_26398);
nand U27774 (N_27774,N_26707,N_26324);
and U27775 (N_27775,N_26663,N_26430);
xnor U27776 (N_27776,N_26116,N_26848);
nor U27777 (N_27777,N_26032,N_26232);
nand U27778 (N_27778,N_26115,N_26031);
or U27779 (N_27779,N_26943,N_26175);
nor U27780 (N_27780,N_26591,N_26053);
nand U27781 (N_27781,N_26682,N_26451);
or U27782 (N_27782,N_26204,N_26704);
or U27783 (N_27783,N_26724,N_26302);
and U27784 (N_27784,N_26357,N_26193);
nand U27785 (N_27785,N_26302,N_26130);
nand U27786 (N_27786,N_26753,N_26071);
xnor U27787 (N_27787,N_26588,N_26959);
nand U27788 (N_27788,N_26221,N_26423);
nand U27789 (N_27789,N_26123,N_26534);
nand U27790 (N_27790,N_26461,N_26487);
nand U27791 (N_27791,N_26348,N_26601);
or U27792 (N_27792,N_26762,N_26850);
xor U27793 (N_27793,N_26956,N_26236);
or U27794 (N_27794,N_26477,N_26250);
or U27795 (N_27795,N_26725,N_26069);
nand U27796 (N_27796,N_26330,N_26595);
nor U27797 (N_27797,N_26163,N_26556);
nor U27798 (N_27798,N_26286,N_26700);
xnor U27799 (N_27799,N_26780,N_26919);
or U27800 (N_27800,N_26155,N_26917);
nand U27801 (N_27801,N_26456,N_26540);
and U27802 (N_27802,N_26462,N_26334);
or U27803 (N_27803,N_26941,N_26246);
xnor U27804 (N_27804,N_26010,N_26352);
or U27805 (N_27805,N_26999,N_26086);
or U27806 (N_27806,N_26352,N_26547);
or U27807 (N_27807,N_26201,N_26121);
xor U27808 (N_27808,N_26496,N_26160);
xor U27809 (N_27809,N_26927,N_26917);
or U27810 (N_27810,N_26518,N_26037);
xor U27811 (N_27811,N_26979,N_26008);
and U27812 (N_27812,N_26693,N_26502);
or U27813 (N_27813,N_26897,N_26363);
xnor U27814 (N_27814,N_26424,N_26473);
or U27815 (N_27815,N_26061,N_26858);
or U27816 (N_27816,N_26637,N_26322);
nand U27817 (N_27817,N_26858,N_26415);
nor U27818 (N_27818,N_26252,N_26292);
nand U27819 (N_27819,N_26933,N_26462);
nor U27820 (N_27820,N_26911,N_26699);
and U27821 (N_27821,N_26213,N_26570);
and U27822 (N_27822,N_26659,N_26613);
and U27823 (N_27823,N_26442,N_26344);
or U27824 (N_27824,N_26066,N_26588);
xor U27825 (N_27825,N_26198,N_26575);
xor U27826 (N_27826,N_26800,N_26450);
or U27827 (N_27827,N_26945,N_26489);
or U27828 (N_27828,N_26747,N_26400);
xnor U27829 (N_27829,N_26562,N_26723);
nand U27830 (N_27830,N_26585,N_26026);
or U27831 (N_27831,N_26316,N_26697);
or U27832 (N_27832,N_26551,N_26113);
xor U27833 (N_27833,N_26985,N_26590);
or U27834 (N_27834,N_26144,N_26327);
xnor U27835 (N_27835,N_26960,N_26368);
and U27836 (N_27836,N_26264,N_26849);
nand U27837 (N_27837,N_26483,N_26819);
or U27838 (N_27838,N_26342,N_26335);
nor U27839 (N_27839,N_26091,N_26810);
nand U27840 (N_27840,N_26742,N_26936);
or U27841 (N_27841,N_26333,N_26059);
xnor U27842 (N_27842,N_26094,N_26169);
xor U27843 (N_27843,N_26292,N_26213);
xnor U27844 (N_27844,N_26610,N_26208);
nand U27845 (N_27845,N_26088,N_26523);
nand U27846 (N_27846,N_26644,N_26097);
or U27847 (N_27847,N_26590,N_26509);
and U27848 (N_27848,N_26580,N_26962);
and U27849 (N_27849,N_26562,N_26707);
nor U27850 (N_27850,N_26090,N_26274);
and U27851 (N_27851,N_26888,N_26785);
nor U27852 (N_27852,N_26778,N_26340);
xnor U27853 (N_27853,N_26531,N_26876);
nor U27854 (N_27854,N_26618,N_26293);
and U27855 (N_27855,N_26272,N_26054);
nand U27856 (N_27856,N_26254,N_26924);
or U27857 (N_27857,N_26931,N_26230);
or U27858 (N_27858,N_26118,N_26827);
nand U27859 (N_27859,N_26994,N_26686);
xnor U27860 (N_27860,N_26189,N_26568);
nand U27861 (N_27861,N_26224,N_26563);
xnor U27862 (N_27862,N_26581,N_26410);
xnor U27863 (N_27863,N_26836,N_26848);
nor U27864 (N_27864,N_26131,N_26296);
nand U27865 (N_27865,N_26580,N_26305);
or U27866 (N_27866,N_26075,N_26470);
nand U27867 (N_27867,N_26830,N_26564);
nand U27868 (N_27868,N_26024,N_26301);
nand U27869 (N_27869,N_26797,N_26536);
and U27870 (N_27870,N_26888,N_26821);
nor U27871 (N_27871,N_26768,N_26583);
or U27872 (N_27872,N_26497,N_26803);
nand U27873 (N_27873,N_26165,N_26044);
nand U27874 (N_27874,N_26854,N_26245);
and U27875 (N_27875,N_26782,N_26792);
xor U27876 (N_27876,N_26760,N_26468);
and U27877 (N_27877,N_26483,N_26609);
and U27878 (N_27878,N_26865,N_26126);
or U27879 (N_27879,N_26506,N_26944);
xnor U27880 (N_27880,N_26262,N_26330);
and U27881 (N_27881,N_26445,N_26506);
nand U27882 (N_27882,N_26047,N_26242);
or U27883 (N_27883,N_26944,N_26957);
nor U27884 (N_27884,N_26380,N_26553);
or U27885 (N_27885,N_26339,N_26125);
and U27886 (N_27886,N_26568,N_26464);
and U27887 (N_27887,N_26588,N_26261);
nor U27888 (N_27888,N_26817,N_26908);
and U27889 (N_27889,N_26227,N_26628);
xor U27890 (N_27890,N_26368,N_26926);
nor U27891 (N_27891,N_26244,N_26503);
and U27892 (N_27892,N_26224,N_26314);
or U27893 (N_27893,N_26318,N_26156);
or U27894 (N_27894,N_26489,N_26218);
xor U27895 (N_27895,N_26432,N_26775);
or U27896 (N_27896,N_26009,N_26073);
nor U27897 (N_27897,N_26568,N_26601);
and U27898 (N_27898,N_26182,N_26005);
nor U27899 (N_27899,N_26438,N_26419);
xor U27900 (N_27900,N_26594,N_26133);
and U27901 (N_27901,N_26348,N_26206);
xnor U27902 (N_27902,N_26844,N_26722);
nand U27903 (N_27903,N_26451,N_26356);
and U27904 (N_27904,N_26624,N_26509);
or U27905 (N_27905,N_26387,N_26245);
nand U27906 (N_27906,N_26261,N_26892);
nor U27907 (N_27907,N_26426,N_26446);
xnor U27908 (N_27908,N_26529,N_26665);
xnor U27909 (N_27909,N_26756,N_26246);
xor U27910 (N_27910,N_26023,N_26063);
nand U27911 (N_27911,N_26958,N_26542);
and U27912 (N_27912,N_26952,N_26865);
xnor U27913 (N_27913,N_26826,N_26612);
xnor U27914 (N_27914,N_26284,N_26341);
and U27915 (N_27915,N_26178,N_26032);
or U27916 (N_27916,N_26719,N_26219);
xor U27917 (N_27917,N_26070,N_26848);
nor U27918 (N_27918,N_26179,N_26182);
xnor U27919 (N_27919,N_26955,N_26307);
and U27920 (N_27920,N_26829,N_26009);
nand U27921 (N_27921,N_26414,N_26408);
or U27922 (N_27922,N_26041,N_26652);
and U27923 (N_27923,N_26704,N_26479);
and U27924 (N_27924,N_26711,N_26579);
nand U27925 (N_27925,N_26845,N_26070);
xnor U27926 (N_27926,N_26196,N_26166);
or U27927 (N_27927,N_26693,N_26200);
nor U27928 (N_27928,N_26887,N_26123);
nor U27929 (N_27929,N_26058,N_26144);
xnor U27930 (N_27930,N_26157,N_26791);
nor U27931 (N_27931,N_26538,N_26479);
or U27932 (N_27932,N_26378,N_26802);
xor U27933 (N_27933,N_26194,N_26405);
nand U27934 (N_27934,N_26046,N_26300);
or U27935 (N_27935,N_26931,N_26660);
nand U27936 (N_27936,N_26482,N_26266);
or U27937 (N_27937,N_26005,N_26255);
or U27938 (N_27938,N_26307,N_26322);
or U27939 (N_27939,N_26687,N_26474);
and U27940 (N_27940,N_26351,N_26559);
nand U27941 (N_27941,N_26035,N_26762);
nand U27942 (N_27942,N_26839,N_26859);
nor U27943 (N_27943,N_26111,N_26284);
and U27944 (N_27944,N_26954,N_26399);
nor U27945 (N_27945,N_26931,N_26149);
and U27946 (N_27946,N_26634,N_26539);
nor U27947 (N_27947,N_26897,N_26004);
nand U27948 (N_27948,N_26834,N_26386);
and U27949 (N_27949,N_26528,N_26013);
and U27950 (N_27950,N_26882,N_26303);
and U27951 (N_27951,N_26501,N_26839);
and U27952 (N_27952,N_26827,N_26080);
nand U27953 (N_27953,N_26247,N_26014);
nor U27954 (N_27954,N_26838,N_26713);
xor U27955 (N_27955,N_26668,N_26978);
and U27956 (N_27956,N_26423,N_26283);
nand U27957 (N_27957,N_26305,N_26618);
nor U27958 (N_27958,N_26182,N_26453);
and U27959 (N_27959,N_26535,N_26266);
nand U27960 (N_27960,N_26307,N_26348);
xor U27961 (N_27961,N_26571,N_26175);
or U27962 (N_27962,N_26110,N_26336);
xor U27963 (N_27963,N_26850,N_26593);
and U27964 (N_27964,N_26044,N_26569);
nor U27965 (N_27965,N_26463,N_26354);
nor U27966 (N_27966,N_26606,N_26487);
nor U27967 (N_27967,N_26392,N_26153);
xor U27968 (N_27968,N_26249,N_26379);
xor U27969 (N_27969,N_26045,N_26661);
nand U27970 (N_27970,N_26121,N_26433);
nor U27971 (N_27971,N_26147,N_26340);
or U27972 (N_27972,N_26943,N_26381);
and U27973 (N_27973,N_26670,N_26740);
and U27974 (N_27974,N_26172,N_26713);
and U27975 (N_27975,N_26745,N_26635);
and U27976 (N_27976,N_26267,N_26490);
nand U27977 (N_27977,N_26748,N_26404);
and U27978 (N_27978,N_26741,N_26762);
or U27979 (N_27979,N_26600,N_26224);
and U27980 (N_27980,N_26202,N_26204);
xnor U27981 (N_27981,N_26277,N_26161);
or U27982 (N_27982,N_26957,N_26553);
and U27983 (N_27983,N_26216,N_26798);
nor U27984 (N_27984,N_26549,N_26613);
xnor U27985 (N_27985,N_26136,N_26736);
nor U27986 (N_27986,N_26460,N_26692);
nand U27987 (N_27987,N_26599,N_26883);
nor U27988 (N_27988,N_26083,N_26041);
or U27989 (N_27989,N_26435,N_26587);
and U27990 (N_27990,N_26894,N_26002);
nor U27991 (N_27991,N_26567,N_26012);
nor U27992 (N_27992,N_26775,N_26844);
nand U27993 (N_27993,N_26992,N_26966);
nand U27994 (N_27994,N_26456,N_26575);
or U27995 (N_27995,N_26971,N_26525);
nor U27996 (N_27996,N_26285,N_26562);
or U27997 (N_27997,N_26840,N_26962);
nand U27998 (N_27998,N_26485,N_26851);
nand U27999 (N_27999,N_26635,N_26428);
and U28000 (N_28000,N_27151,N_27037);
or U28001 (N_28001,N_27223,N_27296);
xor U28002 (N_28002,N_27504,N_27174);
and U28003 (N_28003,N_27340,N_27819);
nor U28004 (N_28004,N_27890,N_27372);
nand U28005 (N_28005,N_27994,N_27526);
nand U28006 (N_28006,N_27239,N_27142);
nor U28007 (N_28007,N_27782,N_27592);
nand U28008 (N_28008,N_27569,N_27393);
nand U28009 (N_28009,N_27662,N_27789);
or U28010 (N_28010,N_27052,N_27824);
nand U28011 (N_28011,N_27800,N_27289);
nand U28012 (N_28012,N_27314,N_27651);
xor U28013 (N_28013,N_27904,N_27531);
xor U28014 (N_28014,N_27941,N_27780);
nand U28015 (N_28015,N_27452,N_27901);
and U28016 (N_28016,N_27467,N_27205);
nand U28017 (N_28017,N_27398,N_27292);
nand U28018 (N_28018,N_27230,N_27363);
nand U28019 (N_28019,N_27401,N_27466);
or U28020 (N_28020,N_27803,N_27365);
or U28021 (N_28021,N_27951,N_27758);
and U28022 (N_28022,N_27720,N_27505);
xnor U28023 (N_28023,N_27529,N_27284);
and U28024 (N_28024,N_27606,N_27442);
nor U28025 (N_28025,N_27580,N_27138);
or U28026 (N_28026,N_27278,N_27282);
nor U28027 (N_28027,N_27381,N_27222);
and U28028 (N_28028,N_27648,N_27764);
nand U28029 (N_28029,N_27128,N_27243);
or U28030 (N_28030,N_27013,N_27250);
or U28031 (N_28031,N_27029,N_27836);
nand U28032 (N_28032,N_27736,N_27880);
or U28033 (N_28033,N_27136,N_27208);
or U28034 (N_28034,N_27711,N_27067);
xnor U28035 (N_28035,N_27016,N_27443);
nor U28036 (N_28036,N_27772,N_27021);
nor U28037 (N_28037,N_27301,N_27437);
and U28038 (N_28038,N_27154,N_27558);
or U28039 (N_28039,N_27487,N_27462);
xor U28040 (N_28040,N_27137,N_27435);
nand U28041 (N_28041,N_27910,N_27473);
and U28042 (N_28042,N_27086,N_27105);
nor U28043 (N_28043,N_27429,N_27081);
or U28044 (N_28044,N_27089,N_27455);
and U28045 (N_28045,N_27659,N_27533);
xnor U28046 (N_28046,N_27317,N_27325);
or U28047 (N_28047,N_27678,N_27369);
or U28048 (N_28048,N_27109,N_27760);
xor U28049 (N_28049,N_27516,N_27981);
xnor U28050 (N_28050,N_27980,N_27170);
xnor U28051 (N_28051,N_27943,N_27729);
or U28052 (N_28052,N_27033,N_27256);
xor U28053 (N_28053,N_27589,N_27091);
nand U28054 (N_28054,N_27587,N_27274);
xnor U28055 (N_28055,N_27578,N_27049);
and U28056 (N_28056,N_27936,N_27433);
xor U28057 (N_28057,N_27629,N_27975);
or U28058 (N_28058,N_27619,N_27304);
xor U28059 (N_28059,N_27641,N_27309);
nor U28060 (N_28060,N_27116,N_27148);
xnor U28061 (N_28061,N_27852,N_27560);
nand U28062 (N_28062,N_27618,N_27972);
and U28063 (N_28063,N_27127,N_27934);
nand U28064 (N_28064,N_27906,N_27734);
nor U28065 (N_28065,N_27679,N_27242);
nor U28066 (N_28066,N_27746,N_27547);
nor U28067 (N_28067,N_27545,N_27155);
xnor U28068 (N_28068,N_27152,N_27140);
xor U28069 (N_28069,N_27982,N_27347);
nor U28070 (N_28070,N_27887,N_27312);
and U28071 (N_28071,N_27791,N_27761);
and U28072 (N_28072,N_27179,N_27123);
and U28073 (N_28073,N_27874,N_27319);
or U28074 (N_28074,N_27058,N_27804);
and U28075 (N_28075,N_27601,N_27733);
xnor U28076 (N_28076,N_27438,N_27693);
xnor U28077 (N_28077,N_27330,N_27846);
nand U28078 (N_28078,N_27502,N_27444);
xnor U28079 (N_28079,N_27726,N_27360);
xor U28080 (N_28080,N_27054,N_27549);
xor U28081 (N_28081,N_27479,N_27719);
nor U28082 (N_28082,N_27106,N_27638);
nor U28083 (N_28083,N_27451,N_27815);
nand U28084 (N_28084,N_27645,N_27305);
xor U28085 (N_28085,N_27912,N_27881);
or U28086 (N_28086,N_27446,N_27318);
xor U28087 (N_28087,N_27627,N_27642);
or U28088 (N_28088,N_27749,N_27727);
nand U28089 (N_28089,N_27050,N_27680);
xnor U28090 (N_28090,N_27053,N_27192);
xor U28091 (N_28091,N_27066,N_27022);
nor U28092 (N_28092,N_27861,N_27636);
or U28093 (N_28093,N_27828,N_27079);
or U28094 (N_28094,N_27345,N_27808);
or U28095 (N_28095,N_27386,N_27624);
xor U28096 (N_28096,N_27577,N_27182);
or U28097 (N_28097,N_27489,N_27919);
and U28098 (N_28098,N_27474,N_27658);
or U28099 (N_28099,N_27983,N_27088);
and U28100 (N_28100,N_27354,N_27788);
nor U28101 (N_28101,N_27425,N_27896);
nand U28102 (N_28102,N_27617,N_27084);
nand U28103 (N_28103,N_27457,N_27279);
and U28104 (N_28104,N_27867,N_27739);
or U28105 (N_28105,N_27161,N_27078);
nor U28106 (N_28106,N_27838,N_27376);
xor U28107 (N_28107,N_27774,N_27754);
nor U28108 (N_28108,N_27518,N_27285);
nor U28109 (N_28109,N_27604,N_27979);
xor U28110 (N_28110,N_27732,N_27610);
or U28111 (N_28111,N_27190,N_27100);
nand U28112 (N_28112,N_27857,N_27463);
nand U28113 (N_28113,N_27620,N_27383);
and U28114 (N_28114,N_27108,N_27964);
and U28115 (N_28115,N_27897,N_27969);
or U28116 (N_28116,N_27527,N_27935);
or U28117 (N_28117,N_27870,N_27656);
nor U28118 (N_28118,N_27755,N_27267);
nand U28119 (N_28119,N_27675,N_27952);
nor U28120 (N_28120,N_27894,N_27763);
xor U28121 (N_28121,N_27023,N_27776);
nor U28122 (N_28122,N_27769,N_27453);
nor U28123 (N_28123,N_27832,N_27588);
and U28124 (N_28124,N_27717,N_27903);
nor U28125 (N_28125,N_27117,N_27930);
nand U28126 (N_28126,N_27441,N_27528);
xor U28127 (N_28127,N_27503,N_27522);
nor U28128 (N_28128,N_27051,N_27406);
xor U28129 (N_28129,N_27408,N_27364);
nor U28130 (N_28130,N_27160,N_27667);
nor U28131 (N_28131,N_27166,N_27963);
nand U28132 (N_28132,N_27775,N_27946);
xnor U28133 (N_28133,N_27576,N_27722);
xnor U28134 (N_28134,N_27837,N_27269);
nor U28135 (N_28135,N_27008,N_27327);
and U28136 (N_28136,N_27939,N_27960);
and U28137 (N_28137,N_27783,N_27920);
nor U28138 (N_28138,N_27011,N_27272);
or U28139 (N_28139,N_27508,N_27598);
or U28140 (N_28140,N_27640,N_27876);
or U28141 (N_28141,N_27388,N_27218);
or U28142 (N_28142,N_27770,N_27114);
xnor U28143 (N_28143,N_27805,N_27225);
or U28144 (N_28144,N_27333,N_27993);
and U28145 (N_28145,N_27958,N_27193);
and U28146 (N_28146,N_27111,N_27907);
xor U28147 (N_28147,N_27976,N_27131);
xor U28148 (N_28148,N_27368,N_27322);
nand U28149 (N_28149,N_27034,N_27180);
nand U28150 (N_28150,N_27313,N_27194);
nand U28151 (N_28151,N_27584,N_27581);
or U28152 (N_28152,N_27570,N_27197);
and U28153 (N_28153,N_27967,N_27071);
xor U28154 (N_28154,N_27921,N_27677);
nor U28155 (N_28155,N_27602,N_27083);
and U28156 (N_28156,N_27821,N_27559);
and U28157 (N_28157,N_27759,N_27799);
xor U28158 (N_28158,N_27063,N_27530);
or U28159 (N_28159,N_27048,N_27352);
and U28160 (N_28160,N_27227,N_27315);
nor U28161 (N_28161,N_27382,N_27355);
xor U28162 (N_28162,N_27399,N_27010);
nand U28163 (N_28163,N_27026,N_27794);
xnor U28164 (N_28164,N_27186,N_27346);
xnor U28165 (N_28165,N_27260,N_27966);
or U28166 (N_28166,N_27064,N_27405);
nand U28167 (N_28167,N_27700,N_27188);
or U28168 (N_28168,N_27778,N_27573);
nand U28169 (N_28169,N_27816,N_27582);
xnor U28170 (N_28170,N_27998,N_27988);
and U28171 (N_28171,N_27370,N_27215);
nand U28172 (N_28172,N_27686,N_27075);
or U28173 (N_28173,N_27594,N_27682);
nor U28174 (N_28174,N_27657,N_27695);
nor U28175 (N_28175,N_27195,N_27377);
nand U28176 (N_28176,N_27575,N_27858);
xnor U28177 (N_28177,N_27019,N_27884);
nor U28178 (N_28178,N_27351,N_27786);
xnor U28179 (N_28179,N_27449,N_27600);
nand U28180 (N_28180,N_27691,N_27673);
and U28181 (N_28181,N_27603,N_27495);
nand U28182 (N_28182,N_27970,N_27550);
and U28183 (N_28183,N_27835,N_27481);
xnor U28184 (N_28184,N_27099,N_27141);
nand U28185 (N_28185,N_27430,N_27404);
nand U28186 (N_28186,N_27510,N_27925);
nor U28187 (N_28187,N_27756,N_27150);
and U28188 (N_28188,N_27506,N_27189);
nand U28189 (N_28189,N_27751,N_27073);
or U28190 (N_28190,N_27830,N_27744);
and U28191 (N_28191,N_27834,N_27057);
or U28192 (N_28192,N_27059,N_27613);
xor U28193 (N_28193,N_27146,N_27974);
and U28194 (N_28194,N_27548,N_27986);
nand U28195 (N_28195,N_27110,N_27041);
and U28196 (N_28196,N_27889,N_27633);
xnor U28197 (N_28197,N_27556,N_27992);
or U28198 (N_28198,N_27701,N_27519);
nor U28199 (N_28199,N_27712,N_27124);
nor U28200 (N_28200,N_27025,N_27220);
or U28201 (N_28201,N_27038,N_27028);
nor U28202 (N_28202,N_27813,N_27321);
xor U28203 (N_28203,N_27164,N_27915);
and U28204 (N_28204,N_27149,N_27997);
nand U28205 (N_28205,N_27737,N_27644);
or U28206 (N_28206,N_27514,N_27294);
nand U28207 (N_28207,N_27718,N_27568);
and U28208 (N_28208,N_27047,N_27157);
nor U28209 (N_28209,N_27216,N_27913);
or U28210 (N_28210,N_27199,N_27286);
nor U28211 (N_28211,N_27407,N_27681);
or U28212 (N_28212,N_27706,N_27426);
xnor U28213 (N_28213,N_27178,N_27924);
or U28214 (N_28214,N_27748,N_27103);
or U28215 (N_28215,N_27043,N_27233);
nor U28216 (N_28216,N_27517,N_27647);
xnor U28217 (N_28217,N_27203,N_27854);
and U28218 (N_28218,N_27957,N_27561);
nor U28219 (N_28219,N_27412,N_27863);
nor U28220 (N_28220,N_27507,N_27524);
xor U28221 (N_28221,N_27480,N_27829);
or U28222 (N_28222,N_27596,N_27090);
and U28223 (N_28223,N_27002,N_27012);
nor U28224 (N_28224,N_27181,N_27177);
or U28225 (N_28225,N_27878,N_27820);
or U28226 (N_28226,N_27932,N_27862);
nor U28227 (N_28227,N_27623,N_27985);
and U28228 (N_28228,N_27306,N_27490);
xnor U28229 (N_28229,N_27886,N_27302);
xnor U28230 (N_28230,N_27696,N_27564);
nor U28231 (N_28231,N_27280,N_27424);
or U28232 (N_28232,N_27167,N_27344);
xor U28233 (N_28233,N_27221,N_27822);
or U28234 (N_28234,N_27316,N_27501);
nand U28235 (N_28235,N_27687,N_27663);
and U28236 (N_28236,N_27851,N_27534);
nor U28237 (N_28237,N_27055,N_27204);
or U28238 (N_28238,N_27491,N_27175);
or U28239 (N_28239,N_27420,N_27207);
and U28240 (N_28240,N_27937,N_27692);
xor U28241 (N_28241,N_27511,N_27035);
xor U28242 (N_28242,N_27273,N_27427);
nor U28243 (N_28243,N_27373,N_27290);
nand U28244 (N_28244,N_27085,N_27353);
nand U28245 (N_28245,N_27908,N_27923);
nor U28246 (N_28246,N_27162,N_27554);
nor U28247 (N_28247,N_27823,N_27866);
or U28248 (N_28248,N_27042,N_27902);
and U28249 (N_28249,N_27076,N_27421);
or U28250 (N_28250,N_27145,N_27459);
nor U28251 (N_28251,N_27056,N_27978);
or U28252 (N_28252,N_27888,N_27999);
and U28253 (N_28253,N_27850,N_27477);
xor U28254 (N_28254,N_27210,N_27120);
or U28255 (N_28255,N_27212,N_27133);
nor U28256 (N_28256,N_27062,N_27525);
nor U28257 (N_28257,N_27509,N_27539);
and U28258 (N_28258,N_27872,N_27257);
or U28259 (N_28259,N_27074,N_27349);
xor U28260 (N_28260,N_27483,N_27882);
nand U28261 (N_28261,N_27476,N_27411);
or U28262 (N_28262,N_27032,N_27336);
and U28263 (N_28263,N_27332,N_27024);
nand U28264 (N_28264,N_27521,N_27699);
or U28265 (N_28265,N_27563,N_27655);
or U28266 (N_28266,N_27731,N_27445);
and U28267 (N_28267,N_27262,N_27567);
or U28268 (N_28268,N_27342,N_27634);
nand U28269 (N_28269,N_27428,N_27362);
xor U28270 (N_28270,N_27367,N_27311);
nor U28271 (N_28271,N_27263,N_27551);
xor U28272 (N_28272,N_27498,N_27209);
xor U28273 (N_28273,N_27949,N_27609);
nand U28274 (N_28274,N_27101,N_27542);
nor U28275 (N_28275,N_27231,N_27134);
xor U28276 (N_28276,N_27954,N_27017);
or U28277 (N_28277,N_27436,N_27320);
xnor U28278 (N_28278,N_27771,N_27684);
and U28279 (N_28279,N_27806,N_27144);
nand U28280 (N_28280,N_27987,N_27891);
xor U28281 (N_28281,N_27069,N_27948);
nand U28282 (N_28282,N_27129,N_27465);
or U28283 (N_28283,N_27859,N_27802);
and U28284 (N_28284,N_27541,N_27817);
nor U28285 (N_28285,N_27475,N_27747);
and U28286 (N_28286,N_27942,N_27478);
xnor U28287 (N_28287,N_27757,N_27909);
xnor U28288 (N_28288,N_27893,N_27497);
or U28289 (N_28289,N_27000,N_27738);
nor U28290 (N_28290,N_27093,N_27403);
nand U28291 (N_28291,N_27014,N_27703);
nor U28292 (N_28292,N_27845,N_27259);
or U28293 (N_28293,N_27841,N_27121);
nand U28294 (N_28294,N_27869,N_27672);
nand U28295 (N_28295,N_27329,N_27400);
and U28296 (N_28296,N_27217,N_27653);
xnor U28297 (N_28297,N_27579,N_27612);
or U28298 (N_28298,N_27730,N_27380);
nor U28299 (N_28299,N_27523,N_27750);
or U28300 (N_28300,N_27065,N_27200);
nor U28301 (N_28301,N_27702,N_27326);
nand U28302 (N_28302,N_27631,N_27665);
xnor U28303 (N_28303,N_27855,N_27875);
and U28304 (N_28304,N_27807,N_27499);
and U28305 (N_28305,N_27307,N_27118);
and U28306 (N_28306,N_27918,N_27469);
xor U28307 (N_28307,N_27268,N_27825);
nand U28308 (N_28308,N_27068,N_27798);
nor U28309 (N_28309,N_27229,N_27356);
xor U28310 (N_28310,N_27418,N_27275);
and U28311 (N_28311,N_27784,N_27070);
nor U28312 (N_28312,N_27096,N_27709);
or U28313 (N_28313,N_27486,N_27255);
and U28314 (N_28314,N_27040,N_27899);
nand U28315 (N_28315,N_27454,N_27295);
or U28316 (N_28316,N_27661,N_27077);
xnor U28317 (N_28317,N_27104,N_27379);
nor U28318 (N_28318,N_27385,N_27300);
nand U28319 (N_28319,N_27842,N_27461);
xor U28320 (N_28320,N_27928,N_27871);
or U28321 (N_28321,N_27753,N_27698);
and U28322 (N_28322,N_27632,N_27538);
nor U28323 (N_28323,N_27323,N_27605);
nor U28324 (N_28324,N_27812,N_27310);
nor U28325 (N_28325,N_27130,N_27492);
nor U28326 (N_28326,N_27950,N_27676);
nand U28327 (N_28327,N_27006,N_27163);
and U28328 (N_28328,N_27060,N_27236);
nor U28329 (N_28329,N_27625,N_27697);
or U28330 (N_28330,N_27585,N_27098);
xor U28331 (N_28331,N_27650,N_27586);
and U28332 (N_28332,N_27571,N_27253);
xor U28333 (N_28333,N_27394,N_27219);
or U28334 (N_28334,N_27015,N_27044);
nor U28335 (N_28335,N_27402,N_27643);
nor U28336 (N_28336,N_27061,N_27991);
or U28337 (N_28337,N_27552,N_27628);
xnor U28338 (N_28338,N_27343,N_27843);
or U28339 (N_28339,N_27003,N_27752);
nand U28340 (N_28340,N_27777,N_27328);
and U28341 (N_28341,N_27536,N_27818);
or U28342 (N_28342,N_27287,N_27254);
or U28343 (N_28343,N_27968,N_27206);
or U28344 (N_28344,N_27947,N_27557);
xor U28345 (N_28345,N_27005,N_27113);
nor U28346 (N_28346,N_27112,N_27690);
nor U28347 (N_28347,N_27555,N_27595);
or U28348 (N_28348,N_27728,N_27288);
and U28349 (N_28349,N_27308,N_27324);
or U28350 (N_28350,N_27856,N_27971);
xor U28351 (N_28351,N_27688,N_27244);
xnor U28352 (N_28352,N_27202,N_27668);
nand U28353 (N_28353,N_27270,N_27371);
nand U28354 (N_28354,N_27996,N_27847);
nor U28355 (N_28355,N_27892,N_27809);
xor U28356 (N_28356,N_27168,N_27674);
and U28357 (N_28357,N_27714,N_27097);
or U28358 (N_28358,N_27652,N_27940);
nand U28359 (N_28359,N_27072,N_27922);
or U28360 (N_28360,N_27434,N_27198);
nand U28361 (N_28361,N_27962,N_27416);
nor U28362 (N_28362,N_27046,N_27515);
nand U28363 (N_28363,N_27384,N_27027);
and U28364 (N_28364,N_27868,N_27249);
xnor U28365 (N_28365,N_27214,N_27773);
nand U28366 (N_28366,N_27251,N_27839);
nand U28367 (N_28367,N_27339,N_27335);
nand U28368 (N_28368,N_27795,N_27258);
and U28369 (N_28369,N_27271,N_27574);
nand U28370 (N_28370,N_27281,N_27460);
nand U28371 (N_28371,N_27735,N_27397);
or U28372 (N_28372,N_27766,N_27018);
xor U28373 (N_28373,N_27448,N_27224);
nand U28374 (N_28374,N_27107,N_27826);
xor U28375 (N_28375,N_27338,N_27183);
xor U28376 (N_28376,N_27172,N_27860);
and U28377 (N_28377,N_27297,N_27520);
nand U28378 (N_28378,N_27187,N_27470);
xnor U28379 (N_28379,N_27785,N_27590);
xnor U28380 (N_28380,N_27374,N_27392);
nor U28381 (N_28381,N_27810,N_27740);
or U28382 (N_28382,N_27710,N_27790);
nor U28383 (N_28383,N_27762,N_27685);
or U28384 (N_28384,N_27119,N_27264);
and U28385 (N_28385,N_27546,N_27705);
xor U28386 (N_28386,N_27626,N_27543);
xor U28387 (N_28387,N_27196,N_27493);
or U28388 (N_28388,N_27669,N_27646);
xor U28389 (N_28389,N_27366,N_27911);
nand U28390 (N_28390,N_27248,N_27599);
xor U28391 (N_28391,N_27126,N_27485);
and U28392 (N_28392,N_27989,N_27361);
or U28393 (N_28393,N_27622,N_27234);
and U28394 (N_28394,N_27955,N_27232);
nor U28395 (N_28395,N_27844,N_27811);
xor U28396 (N_28396,N_27413,N_27637);
nor U28397 (N_28397,N_27608,N_27092);
or U28398 (N_28398,N_27905,N_27494);
or U28399 (N_28399,N_27607,N_27931);
xor U28400 (N_28400,N_27898,N_27431);
or U28401 (N_28401,N_27848,N_27419);
nor U28402 (N_28402,N_27916,N_27593);
and U28403 (N_28403,N_27357,N_27303);
nand U28404 (N_28404,N_27337,N_27139);
nand U28405 (N_28405,N_27191,N_27537);
nand U28406 (N_28406,N_27885,N_27562);
xor U28407 (N_28407,N_27375,N_27879);
and U28408 (N_28408,N_27864,N_27990);
and U28409 (N_28409,N_27649,N_27156);
nand U28410 (N_28410,N_27953,N_27378);
nor U28411 (N_28411,N_27395,N_27414);
nand U28412 (N_28412,N_27410,N_27660);
nor U28413 (N_28413,N_27933,N_27045);
nor U28414 (N_28414,N_27779,N_27241);
and U28415 (N_28415,N_27616,N_27787);
xnor U28416 (N_28416,N_27927,N_27961);
nand U28417 (N_28417,N_27350,N_27597);
or U28418 (N_28418,N_27277,N_27283);
or U28419 (N_28419,N_27873,N_27132);
and U28420 (N_28420,N_27237,N_27840);
and U28421 (N_28421,N_27184,N_27147);
nand U28422 (N_28422,N_27211,N_27488);
or U28423 (N_28423,N_27849,N_27039);
and U28424 (N_28424,N_27664,N_27228);
nor U28425 (N_28425,N_27235,N_27796);
and U28426 (N_28426,N_27725,N_27417);
nor U28427 (N_28427,N_27389,N_27814);
nand U28428 (N_28428,N_27995,N_27447);
or U28429 (N_28429,N_27635,N_27439);
or U28430 (N_28430,N_27895,N_27298);
xor U28431 (N_28431,N_27007,N_27591);
nor U28432 (N_28432,N_27713,N_27291);
nor U28433 (N_28433,N_27456,N_27768);
nor U28434 (N_28434,N_27716,N_27391);
xor U28435 (N_28435,N_27415,N_27082);
nand U28436 (N_28436,N_27036,N_27793);
nand U28437 (N_28437,N_27334,N_27422);
and U28438 (N_28438,N_27240,N_27938);
or U28439 (N_28439,N_27471,N_27977);
or U28440 (N_28440,N_27261,N_27171);
nor U28441 (N_28441,N_27831,N_27293);
nand U28442 (N_28442,N_27185,N_27201);
and U28443 (N_28443,N_27169,N_27423);
xnor U28444 (N_28444,N_27331,N_27031);
nor U28445 (N_28445,N_27801,N_27276);
or U28446 (N_28446,N_27572,N_27009);
xnor U28447 (N_28447,N_27238,N_27125);
and U28448 (N_28448,N_27513,N_27566);
xor U28449 (N_28449,N_27135,N_27450);
xnor U28450 (N_28450,N_27745,N_27689);
xnor U28451 (N_28451,N_27917,N_27512);
or U28452 (N_28452,N_27944,N_27540);
and U28453 (N_28453,N_27080,N_27914);
xor U28454 (N_28454,N_27707,N_27496);
nor U28455 (N_28455,N_27468,N_27544);
xor U28456 (N_28456,N_27724,N_27926);
nor U28457 (N_28457,N_27670,N_27159);
and U28458 (N_28458,N_27797,N_27553);
and U28459 (N_28459,N_27409,N_27615);
xor U28460 (N_28460,N_27165,N_27900);
or U28461 (N_28461,N_27247,N_27266);
nor U28462 (N_28462,N_27348,N_27095);
xor U28463 (N_28463,N_27611,N_27341);
or U28464 (N_28464,N_27458,N_27583);
or U28465 (N_28465,N_27153,N_27956);
xor U28466 (N_28466,N_27765,N_27500);
nor U28467 (N_28467,N_27715,N_27158);
nand U28468 (N_28468,N_27621,N_27143);
nand U28469 (N_28469,N_27020,N_27959);
nor U28470 (N_28470,N_27767,N_27265);
nor U28471 (N_28471,N_27877,N_27472);
or U28472 (N_28472,N_27464,N_27929);
xnor U28473 (N_28473,N_27087,N_27654);
nor U28474 (N_28474,N_27226,N_27094);
nor U28475 (N_28475,N_27173,N_27865);
nand U28476 (N_28476,N_27245,N_27299);
or U28477 (N_28477,N_27827,N_27359);
nor U28478 (N_28478,N_27945,N_27535);
nand U28479 (N_28479,N_27630,N_27639);
nor U28480 (N_28480,N_27246,N_27390);
and U28481 (N_28481,N_27792,N_27742);
nor U28482 (N_28482,N_27484,N_27666);
and U28483 (N_28483,N_27853,N_27358);
and U28484 (N_28484,N_27973,N_27102);
or U28485 (N_28485,N_27440,N_27741);
and U28486 (N_28486,N_27708,N_27001);
or U28487 (N_28487,N_27532,N_27176);
or U28488 (N_28488,N_27213,N_27781);
xor U28489 (N_28489,N_27030,N_27671);
nor U28490 (N_28490,N_27252,N_27004);
xnor U28491 (N_28491,N_27432,N_27387);
nor U28492 (N_28492,N_27883,N_27723);
xnor U28493 (N_28493,N_27694,N_27115);
or U28494 (N_28494,N_27683,N_27614);
or U28495 (N_28495,N_27721,N_27984);
or U28496 (N_28496,N_27743,N_27482);
or U28497 (N_28497,N_27704,N_27396);
xor U28498 (N_28498,N_27122,N_27833);
or U28499 (N_28499,N_27965,N_27565);
or U28500 (N_28500,N_27388,N_27508);
and U28501 (N_28501,N_27301,N_27621);
or U28502 (N_28502,N_27274,N_27014);
or U28503 (N_28503,N_27306,N_27254);
nor U28504 (N_28504,N_27169,N_27047);
nor U28505 (N_28505,N_27750,N_27386);
and U28506 (N_28506,N_27679,N_27299);
xnor U28507 (N_28507,N_27175,N_27350);
and U28508 (N_28508,N_27552,N_27612);
nand U28509 (N_28509,N_27912,N_27805);
xor U28510 (N_28510,N_27951,N_27539);
and U28511 (N_28511,N_27236,N_27888);
xor U28512 (N_28512,N_27153,N_27352);
xnor U28513 (N_28513,N_27509,N_27357);
or U28514 (N_28514,N_27113,N_27401);
and U28515 (N_28515,N_27549,N_27974);
xnor U28516 (N_28516,N_27350,N_27725);
nand U28517 (N_28517,N_27923,N_27975);
nor U28518 (N_28518,N_27173,N_27267);
nor U28519 (N_28519,N_27491,N_27568);
nand U28520 (N_28520,N_27097,N_27533);
or U28521 (N_28521,N_27428,N_27509);
nor U28522 (N_28522,N_27915,N_27566);
nor U28523 (N_28523,N_27950,N_27440);
nor U28524 (N_28524,N_27733,N_27985);
or U28525 (N_28525,N_27975,N_27254);
and U28526 (N_28526,N_27516,N_27939);
nand U28527 (N_28527,N_27173,N_27593);
or U28528 (N_28528,N_27258,N_27657);
and U28529 (N_28529,N_27463,N_27802);
or U28530 (N_28530,N_27627,N_27982);
nor U28531 (N_28531,N_27309,N_27496);
and U28532 (N_28532,N_27930,N_27454);
and U28533 (N_28533,N_27106,N_27034);
xor U28534 (N_28534,N_27235,N_27458);
nor U28535 (N_28535,N_27759,N_27468);
or U28536 (N_28536,N_27083,N_27518);
and U28537 (N_28537,N_27164,N_27282);
or U28538 (N_28538,N_27360,N_27172);
and U28539 (N_28539,N_27576,N_27633);
nand U28540 (N_28540,N_27739,N_27855);
and U28541 (N_28541,N_27311,N_27530);
nand U28542 (N_28542,N_27800,N_27428);
nor U28543 (N_28543,N_27313,N_27163);
nand U28544 (N_28544,N_27801,N_27158);
or U28545 (N_28545,N_27192,N_27448);
nor U28546 (N_28546,N_27152,N_27993);
and U28547 (N_28547,N_27594,N_27553);
nand U28548 (N_28548,N_27666,N_27834);
or U28549 (N_28549,N_27694,N_27570);
nand U28550 (N_28550,N_27940,N_27970);
xor U28551 (N_28551,N_27405,N_27641);
xnor U28552 (N_28552,N_27861,N_27974);
or U28553 (N_28553,N_27217,N_27453);
xnor U28554 (N_28554,N_27683,N_27898);
xor U28555 (N_28555,N_27451,N_27979);
or U28556 (N_28556,N_27506,N_27358);
and U28557 (N_28557,N_27469,N_27211);
or U28558 (N_28558,N_27904,N_27826);
or U28559 (N_28559,N_27956,N_27075);
nand U28560 (N_28560,N_27115,N_27428);
or U28561 (N_28561,N_27274,N_27462);
and U28562 (N_28562,N_27594,N_27873);
and U28563 (N_28563,N_27519,N_27805);
xor U28564 (N_28564,N_27595,N_27429);
nor U28565 (N_28565,N_27335,N_27804);
nand U28566 (N_28566,N_27446,N_27925);
or U28567 (N_28567,N_27989,N_27725);
or U28568 (N_28568,N_27132,N_27701);
and U28569 (N_28569,N_27805,N_27625);
nor U28570 (N_28570,N_27993,N_27896);
nand U28571 (N_28571,N_27879,N_27476);
nand U28572 (N_28572,N_27649,N_27981);
and U28573 (N_28573,N_27840,N_27841);
nand U28574 (N_28574,N_27065,N_27439);
or U28575 (N_28575,N_27636,N_27396);
nor U28576 (N_28576,N_27076,N_27942);
nand U28577 (N_28577,N_27747,N_27952);
or U28578 (N_28578,N_27149,N_27365);
xor U28579 (N_28579,N_27293,N_27645);
xor U28580 (N_28580,N_27225,N_27197);
or U28581 (N_28581,N_27773,N_27911);
nor U28582 (N_28582,N_27114,N_27805);
xnor U28583 (N_28583,N_27222,N_27095);
nor U28584 (N_28584,N_27268,N_27700);
or U28585 (N_28585,N_27681,N_27388);
nand U28586 (N_28586,N_27562,N_27538);
or U28587 (N_28587,N_27762,N_27894);
or U28588 (N_28588,N_27909,N_27792);
nor U28589 (N_28589,N_27936,N_27413);
nand U28590 (N_28590,N_27413,N_27521);
and U28591 (N_28591,N_27253,N_27003);
and U28592 (N_28592,N_27361,N_27211);
and U28593 (N_28593,N_27803,N_27640);
and U28594 (N_28594,N_27579,N_27099);
xor U28595 (N_28595,N_27328,N_27043);
or U28596 (N_28596,N_27210,N_27189);
nor U28597 (N_28597,N_27057,N_27662);
nor U28598 (N_28598,N_27440,N_27617);
or U28599 (N_28599,N_27838,N_27080);
xor U28600 (N_28600,N_27536,N_27568);
nand U28601 (N_28601,N_27615,N_27204);
xor U28602 (N_28602,N_27607,N_27412);
and U28603 (N_28603,N_27355,N_27131);
nor U28604 (N_28604,N_27899,N_27302);
nand U28605 (N_28605,N_27383,N_27626);
nand U28606 (N_28606,N_27682,N_27070);
nor U28607 (N_28607,N_27901,N_27489);
or U28608 (N_28608,N_27539,N_27156);
and U28609 (N_28609,N_27396,N_27763);
or U28610 (N_28610,N_27133,N_27773);
and U28611 (N_28611,N_27267,N_27923);
nor U28612 (N_28612,N_27451,N_27443);
xor U28613 (N_28613,N_27966,N_27616);
nor U28614 (N_28614,N_27315,N_27100);
nor U28615 (N_28615,N_27272,N_27384);
xnor U28616 (N_28616,N_27380,N_27874);
and U28617 (N_28617,N_27428,N_27149);
or U28618 (N_28618,N_27863,N_27734);
or U28619 (N_28619,N_27341,N_27825);
nor U28620 (N_28620,N_27972,N_27210);
xor U28621 (N_28621,N_27780,N_27445);
nor U28622 (N_28622,N_27288,N_27658);
nand U28623 (N_28623,N_27988,N_27337);
or U28624 (N_28624,N_27358,N_27906);
xor U28625 (N_28625,N_27538,N_27120);
or U28626 (N_28626,N_27067,N_27827);
nor U28627 (N_28627,N_27344,N_27005);
nor U28628 (N_28628,N_27161,N_27273);
nor U28629 (N_28629,N_27874,N_27355);
or U28630 (N_28630,N_27704,N_27465);
nand U28631 (N_28631,N_27297,N_27364);
nor U28632 (N_28632,N_27931,N_27989);
xnor U28633 (N_28633,N_27851,N_27483);
nor U28634 (N_28634,N_27854,N_27911);
and U28635 (N_28635,N_27692,N_27610);
or U28636 (N_28636,N_27040,N_27107);
xor U28637 (N_28637,N_27759,N_27712);
or U28638 (N_28638,N_27573,N_27706);
or U28639 (N_28639,N_27353,N_27196);
xor U28640 (N_28640,N_27026,N_27362);
xor U28641 (N_28641,N_27349,N_27292);
or U28642 (N_28642,N_27622,N_27834);
nor U28643 (N_28643,N_27936,N_27641);
nand U28644 (N_28644,N_27757,N_27254);
nor U28645 (N_28645,N_27050,N_27870);
xor U28646 (N_28646,N_27676,N_27922);
nand U28647 (N_28647,N_27369,N_27956);
and U28648 (N_28648,N_27683,N_27158);
nand U28649 (N_28649,N_27192,N_27535);
nor U28650 (N_28650,N_27615,N_27317);
nand U28651 (N_28651,N_27408,N_27197);
nand U28652 (N_28652,N_27877,N_27823);
nor U28653 (N_28653,N_27783,N_27940);
xor U28654 (N_28654,N_27038,N_27566);
nand U28655 (N_28655,N_27144,N_27304);
xor U28656 (N_28656,N_27954,N_27253);
nor U28657 (N_28657,N_27136,N_27129);
xor U28658 (N_28658,N_27954,N_27329);
nand U28659 (N_28659,N_27402,N_27489);
xor U28660 (N_28660,N_27569,N_27787);
nor U28661 (N_28661,N_27228,N_27762);
or U28662 (N_28662,N_27929,N_27499);
nor U28663 (N_28663,N_27501,N_27249);
or U28664 (N_28664,N_27746,N_27715);
xnor U28665 (N_28665,N_27426,N_27021);
xor U28666 (N_28666,N_27038,N_27374);
nand U28667 (N_28667,N_27097,N_27860);
nor U28668 (N_28668,N_27591,N_27020);
or U28669 (N_28669,N_27291,N_27398);
or U28670 (N_28670,N_27837,N_27461);
nor U28671 (N_28671,N_27450,N_27256);
and U28672 (N_28672,N_27737,N_27776);
or U28673 (N_28673,N_27721,N_27440);
nor U28674 (N_28674,N_27860,N_27210);
or U28675 (N_28675,N_27935,N_27096);
xnor U28676 (N_28676,N_27366,N_27808);
xor U28677 (N_28677,N_27205,N_27372);
xnor U28678 (N_28678,N_27370,N_27577);
nor U28679 (N_28679,N_27404,N_27638);
nand U28680 (N_28680,N_27740,N_27216);
xnor U28681 (N_28681,N_27655,N_27325);
nand U28682 (N_28682,N_27497,N_27730);
or U28683 (N_28683,N_27292,N_27875);
nand U28684 (N_28684,N_27604,N_27349);
or U28685 (N_28685,N_27412,N_27202);
xor U28686 (N_28686,N_27867,N_27381);
nor U28687 (N_28687,N_27657,N_27779);
xnor U28688 (N_28688,N_27540,N_27547);
and U28689 (N_28689,N_27798,N_27037);
nor U28690 (N_28690,N_27748,N_27148);
nand U28691 (N_28691,N_27937,N_27326);
nor U28692 (N_28692,N_27364,N_27586);
or U28693 (N_28693,N_27883,N_27478);
xnor U28694 (N_28694,N_27879,N_27419);
nor U28695 (N_28695,N_27209,N_27360);
xor U28696 (N_28696,N_27321,N_27614);
or U28697 (N_28697,N_27986,N_27518);
xor U28698 (N_28698,N_27809,N_27729);
xor U28699 (N_28699,N_27461,N_27343);
nand U28700 (N_28700,N_27252,N_27459);
or U28701 (N_28701,N_27377,N_27436);
nor U28702 (N_28702,N_27211,N_27683);
nor U28703 (N_28703,N_27732,N_27944);
nand U28704 (N_28704,N_27257,N_27347);
nor U28705 (N_28705,N_27264,N_27241);
nand U28706 (N_28706,N_27362,N_27331);
or U28707 (N_28707,N_27991,N_27455);
nor U28708 (N_28708,N_27449,N_27989);
nor U28709 (N_28709,N_27009,N_27083);
or U28710 (N_28710,N_27721,N_27604);
and U28711 (N_28711,N_27908,N_27477);
xnor U28712 (N_28712,N_27108,N_27089);
nor U28713 (N_28713,N_27200,N_27554);
xor U28714 (N_28714,N_27265,N_27463);
xor U28715 (N_28715,N_27410,N_27163);
nor U28716 (N_28716,N_27624,N_27983);
nor U28717 (N_28717,N_27704,N_27670);
nand U28718 (N_28718,N_27737,N_27078);
nor U28719 (N_28719,N_27249,N_27207);
or U28720 (N_28720,N_27167,N_27142);
xor U28721 (N_28721,N_27077,N_27321);
xor U28722 (N_28722,N_27176,N_27265);
and U28723 (N_28723,N_27299,N_27437);
nor U28724 (N_28724,N_27930,N_27177);
or U28725 (N_28725,N_27134,N_27287);
or U28726 (N_28726,N_27062,N_27808);
or U28727 (N_28727,N_27250,N_27129);
xor U28728 (N_28728,N_27803,N_27919);
and U28729 (N_28729,N_27257,N_27555);
and U28730 (N_28730,N_27746,N_27107);
xor U28731 (N_28731,N_27525,N_27153);
and U28732 (N_28732,N_27869,N_27521);
or U28733 (N_28733,N_27640,N_27009);
and U28734 (N_28734,N_27363,N_27310);
nor U28735 (N_28735,N_27168,N_27265);
or U28736 (N_28736,N_27735,N_27301);
and U28737 (N_28737,N_27063,N_27269);
and U28738 (N_28738,N_27960,N_27950);
nand U28739 (N_28739,N_27569,N_27699);
nor U28740 (N_28740,N_27143,N_27994);
nand U28741 (N_28741,N_27572,N_27674);
xor U28742 (N_28742,N_27584,N_27962);
nand U28743 (N_28743,N_27990,N_27200);
xnor U28744 (N_28744,N_27664,N_27005);
or U28745 (N_28745,N_27393,N_27866);
and U28746 (N_28746,N_27002,N_27297);
xnor U28747 (N_28747,N_27652,N_27350);
and U28748 (N_28748,N_27477,N_27020);
nor U28749 (N_28749,N_27907,N_27501);
or U28750 (N_28750,N_27193,N_27949);
nor U28751 (N_28751,N_27901,N_27725);
nand U28752 (N_28752,N_27665,N_27733);
and U28753 (N_28753,N_27174,N_27806);
and U28754 (N_28754,N_27469,N_27758);
and U28755 (N_28755,N_27840,N_27813);
nand U28756 (N_28756,N_27777,N_27500);
and U28757 (N_28757,N_27389,N_27580);
or U28758 (N_28758,N_27727,N_27282);
or U28759 (N_28759,N_27087,N_27265);
nand U28760 (N_28760,N_27495,N_27482);
nor U28761 (N_28761,N_27407,N_27024);
and U28762 (N_28762,N_27114,N_27389);
or U28763 (N_28763,N_27197,N_27114);
xnor U28764 (N_28764,N_27339,N_27629);
nand U28765 (N_28765,N_27761,N_27899);
or U28766 (N_28766,N_27744,N_27869);
xor U28767 (N_28767,N_27443,N_27225);
nor U28768 (N_28768,N_27725,N_27895);
or U28769 (N_28769,N_27596,N_27024);
nor U28770 (N_28770,N_27774,N_27729);
or U28771 (N_28771,N_27057,N_27375);
nand U28772 (N_28772,N_27562,N_27393);
and U28773 (N_28773,N_27794,N_27741);
and U28774 (N_28774,N_27674,N_27979);
or U28775 (N_28775,N_27475,N_27870);
nand U28776 (N_28776,N_27010,N_27387);
xnor U28777 (N_28777,N_27715,N_27312);
and U28778 (N_28778,N_27538,N_27122);
nand U28779 (N_28779,N_27380,N_27519);
nand U28780 (N_28780,N_27832,N_27161);
nor U28781 (N_28781,N_27964,N_27680);
and U28782 (N_28782,N_27597,N_27158);
nand U28783 (N_28783,N_27674,N_27983);
xor U28784 (N_28784,N_27974,N_27294);
nand U28785 (N_28785,N_27291,N_27053);
nand U28786 (N_28786,N_27920,N_27119);
nand U28787 (N_28787,N_27788,N_27450);
or U28788 (N_28788,N_27642,N_27391);
or U28789 (N_28789,N_27294,N_27078);
nor U28790 (N_28790,N_27914,N_27364);
nor U28791 (N_28791,N_27430,N_27695);
xor U28792 (N_28792,N_27327,N_27096);
and U28793 (N_28793,N_27971,N_27726);
and U28794 (N_28794,N_27101,N_27525);
nand U28795 (N_28795,N_27621,N_27282);
xor U28796 (N_28796,N_27577,N_27994);
or U28797 (N_28797,N_27585,N_27798);
nand U28798 (N_28798,N_27729,N_27520);
xor U28799 (N_28799,N_27998,N_27294);
or U28800 (N_28800,N_27173,N_27806);
nor U28801 (N_28801,N_27378,N_27251);
or U28802 (N_28802,N_27499,N_27471);
nand U28803 (N_28803,N_27490,N_27249);
or U28804 (N_28804,N_27603,N_27418);
nor U28805 (N_28805,N_27038,N_27886);
nand U28806 (N_28806,N_27050,N_27556);
nand U28807 (N_28807,N_27979,N_27849);
or U28808 (N_28808,N_27158,N_27621);
nor U28809 (N_28809,N_27584,N_27748);
or U28810 (N_28810,N_27566,N_27972);
nand U28811 (N_28811,N_27964,N_27167);
nand U28812 (N_28812,N_27047,N_27516);
and U28813 (N_28813,N_27902,N_27893);
or U28814 (N_28814,N_27735,N_27373);
and U28815 (N_28815,N_27075,N_27558);
nand U28816 (N_28816,N_27560,N_27714);
xnor U28817 (N_28817,N_27684,N_27400);
and U28818 (N_28818,N_27279,N_27476);
xnor U28819 (N_28819,N_27991,N_27783);
or U28820 (N_28820,N_27168,N_27964);
or U28821 (N_28821,N_27809,N_27206);
xor U28822 (N_28822,N_27810,N_27675);
or U28823 (N_28823,N_27691,N_27022);
nor U28824 (N_28824,N_27359,N_27397);
or U28825 (N_28825,N_27885,N_27320);
nand U28826 (N_28826,N_27476,N_27761);
xor U28827 (N_28827,N_27510,N_27173);
or U28828 (N_28828,N_27944,N_27135);
nand U28829 (N_28829,N_27122,N_27368);
nand U28830 (N_28830,N_27419,N_27195);
nand U28831 (N_28831,N_27540,N_27009);
nor U28832 (N_28832,N_27904,N_27995);
xor U28833 (N_28833,N_27012,N_27058);
xnor U28834 (N_28834,N_27774,N_27545);
xnor U28835 (N_28835,N_27873,N_27531);
and U28836 (N_28836,N_27897,N_27112);
and U28837 (N_28837,N_27495,N_27925);
nor U28838 (N_28838,N_27290,N_27308);
and U28839 (N_28839,N_27763,N_27070);
and U28840 (N_28840,N_27343,N_27955);
nand U28841 (N_28841,N_27909,N_27979);
nand U28842 (N_28842,N_27955,N_27739);
and U28843 (N_28843,N_27780,N_27823);
and U28844 (N_28844,N_27375,N_27551);
and U28845 (N_28845,N_27558,N_27083);
and U28846 (N_28846,N_27663,N_27623);
nor U28847 (N_28847,N_27264,N_27080);
or U28848 (N_28848,N_27107,N_27450);
nand U28849 (N_28849,N_27180,N_27453);
or U28850 (N_28850,N_27473,N_27917);
xnor U28851 (N_28851,N_27865,N_27785);
nor U28852 (N_28852,N_27476,N_27510);
and U28853 (N_28853,N_27415,N_27976);
and U28854 (N_28854,N_27174,N_27725);
nand U28855 (N_28855,N_27752,N_27926);
or U28856 (N_28856,N_27063,N_27900);
nand U28857 (N_28857,N_27042,N_27193);
or U28858 (N_28858,N_27830,N_27132);
or U28859 (N_28859,N_27667,N_27236);
xor U28860 (N_28860,N_27128,N_27122);
or U28861 (N_28861,N_27937,N_27539);
or U28862 (N_28862,N_27669,N_27499);
xor U28863 (N_28863,N_27357,N_27067);
and U28864 (N_28864,N_27100,N_27714);
nor U28865 (N_28865,N_27784,N_27007);
xor U28866 (N_28866,N_27450,N_27488);
or U28867 (N_28867,N_27000,N_27988);
nand U28868 (N_28868,N_27975,N_27047);
nor U28869 (N_28869,N_27316,N_27649);
and U28870 (N_28870,N_27842,N_27336);
nand U28871 (N_28871,N_27714,N_27567);
xnor U28872 (N_28872,N_27522,N_27121);
nor U28873 (N_28873,N_27371,N_27029);
and U28874 (N_28874,N_27028,N_27941);
nor U28875 (N_28875,N_27071,N_27442);
nand U28876 (N_28876,N_27051,N_27180);
nor U28877 (N_28877,N_27487,N_27800);
xor U28878 (N_28878,N_27132,N_27280);
or U28879 (N_28879,N_27455,N_27684);
xor U28880 (N_28880,N_27695,N_27476);
and U28881 (N_28881,N_27965,N_27863);
or U28882 (N_28882,N_27935,N_27590);
xor U28883 (N_28883,N_27874,N_27029);
nor U28884 (N_28884,N_27527,N_27601);
or U28885 (N_28885,N_27432,N_27323);
xor U28886 (N_28886,N_27990,N_27208);
or U28887 (N_28887,N_27849,N_27168);
nand U28888 (N_28888,N_27600,N_27837);
nand U28889 (N_28889,N_27865,N_27211);
xor U28890 (N_28890,N_27832,N_27887);
and U28891 (N_28891,N_27371,N_27684);
nor U28892 (N_28892,N_27657,N_27749);
nor U28893 (N_28893,N_27762,N_27276);
nand U28894 (N_28894,N_27718,N_27319);
xor U28895 (N_28895,N_27714,N_27828);
and U28896 (N_28896,N_27288,N_27838);
or U28897 (N_28897,N_27475,N_27857);
or U28898 (N_28898,N_27735,N_27425);
or U28899 (N_28899,N_27112,N_27865);
nand U28900 (N_28900,N_27065,N_27127);
xor U28901 (N_28901,N_27978,N_27981);
and U28902 (N_28902,N_27312,N_27943);
and U28903 (N_28903,N_27821,N_27885);
xor U28904 (N_28904,N_27979,N_27415);
nand U28905 (N_28905,N_27700,N_27383);
nor U28906 (N_28906,N_27804,N_27141);
nor U28907 (N_28907,N_27237,N_27471);
xnor U28908 (N_28908,N_27138,N_27802);
nand U28909 (N_28909,N_27403,N_27356);
or U28910 (N_28910,N_27285,N_27835);
xnor U28911 (N_28911,N_27629,N_27882);
nand U28912 (N_28912,N_27011,N_27956);
and U28913 (N_28913,N_27779,N_27873);
nand U28914 (N_28914,N_27703,N_27420);
xor U28915 (N_28915,N_27390,N_27946);
nand U28916 (N_28916,N_27642,N_27230);
nand U28917 (N_28917,N_27221,N_27011);
or U28918 (N_28918,N_27413,N_27350);
nor U28919 (N_28919,N_27389,N_27142);
or U28920 (N_28920,N_27724,N_27409);
nand U28921 (N_28921,N_27376,N_27985);
nor U28922 (N_28922,N_27627,N_27481);
xnor U28923 (N_28923,N_27055,N_27249);
or U28924 (N_28924,N_27660,N_27596);
nor U28925 (N_28925,N_27062,N_27477);
nor U28926 (N_28926,N_27607,N_27115);
nor U28927 (N_28927,N_27634,N_27419);
nand U28928 (N_28928,N_27794,N_27413);
or U28929 (N_28929,N_27625,N_27750);
nor U28930 (N_28930,N_27639,N_27279);
nand U28931 (N_28931,N_27113,N_27884);
or U28932 (N_28932,N_27529,N_27991);
and U28933 (N_28933,N_27634,N_27533);
nor U28934 (N_28934,N_27647,N_27701);
xor U28935 (N_28935,N_27217,N_27353);
nand U28936 (N_28936,N_27759,N_27679);
nand U28937 (N_28937,N_27588,N_27105);
and U28938 (N_28938,N_27515,N_27382);
nand U28939 (N_28939,N_27963,N_27874);
or U28940 (N_28940,N_27122,N_27100);
xnor U28941 (N_28941,N_27915,N_27253);
or U28942 (N_28942,N_27389,N_27406);
xnor U28943 (N_28943,N_27661,N_27025);
or U28944 (N_28944,N_27190,N_27966);
xor U28945 (N_28945,N_27428,N_27407);
nor U28946 (N_28946,N_27236,N_27755);
xnor U28947 (N_28947,N_27560,N_27407);
or U28948 (N_28948,N_27571,N_27119);
nand U28949 (N_28949,N_27827,N_27200);
xor U28950 (N_28950,N_27657,N_27304);
and U28951 (N_28951,N_27335,N_27860);
or U28952 (N_28952,N_27378,N_27700);
and U28953 (N_28953,N_27089,N_27884);
xor U28954 (N_28954,N_27741,N_27639);
nor U28955 (N_28955,N_27873,N_27825);
xnor U28956 (N_28956,N_27078,N_27081);
xor U28957 (N_28957,N_27011,N_27608);
xor U28958 (N_28958,N_27494,N_27733);
or U28959 (N_28959,N_27804,N_27930);
and U28960 (N_28960,N_27921,N_27990);
and U28961 (N_28961,N_27970,N_27962);
nor U28962 (N_28962,N_27894,N_27253);
xor U28963 (N_28963,N_27929,N_27222);
and U28964 (N_28964,N_27530,N_27565);
or U28965 (N_28965,N_27745,N_27027);
nand U28966 (N_28966,N_27228,N_27060);
and U28967 (N_28967,N_27518,N_27558);
and U28968 (N_28968,N_27032,N_27769);
xor U28969 (N_28969,N_27860,N_27556);
nor U28970 (N_28970,N_27987,N_27484);
or U28971 (N_28971,N_27870,N_27166);
and U28972 (N_28972,N_27744,N_27764);
and U28973 (N_28973,N_27969,N_27906);
or U28974 (N_28974,N_27893,N_27095);
and U28975 (N_28975,N_27637,N_27550);
nor U28976 (N_28976,N_27457,N_27791);
xor U28977 (N_28977,N_27338,N_27827);
and U28978 (N_28978,N_27438,N_27690);
nor U28979 (N_28979,N_27142,N_27081);
nor U28980 (N_28980,N_27679,N_27486);
nand U28981 (N_28981,N_27071,N_27532);
xor U28982 (N_28982,N_27099,N_27885);
xnor U28983 (N_28983,N_27007,N_27929);
nor U28984 (N_28984,N_27675,N_27608);
and U28985 (N_28985,N_27173,N_27386);
or U28986 (N_28986,N_27849,N_27938);
or U28987 (N_28987,N_27881,N_27914);
nor U28988 (N_28988,N_27501,N_27334);
nand U28989 (N_28989,N_27219,N_27095);
nor U28990 (N_28990,N_27455,N_27906);
xor U28991 (N_28991,N_27486,N_27268);
and U28992 (N_28992,N_27341,N_27216);
nand U28993 (N_28993,N_27958,N_27671);
or U28994 (N_28994,N_27796,N_27080);
nor U28995 (N_28995,N_27243,N_27253);
nand U28996 (N_28996,N_27581,N_27492);
and U28997 (N_28997,N_27380,N_27812);
nor U28998 (N_28998,N_27995,N_27059);
or U28999 (N_28999,N_27010,N_27548);
nor U29000 (N_29000,N_28406,N_28057);
xor U29001 (N_29001,N_28125,N_28313);
or U29002 (N_29002,N_28303,N_28873);
xor U29003 (N_29003,N_28823,N_28563);
xor U29004 (N_29004,N_28705,N_28960);
nor U29005 (N_29005,N_28207,N_28425);
and U29006 (N_29006,N_28424,N_28200);
nand U29007 (N_29007,N_28131,N_28037);
nor U29008 (N_29008,N_28801,N_28712);
xor U29009 (N_29009,N_28306,N_28470);
nand U29010 (N_29010,N_28983,N_28187);
nand U29011 (N_29011,N_28922,N_28546);
nand U29012 (N_29012,N_28522,N_28161);
nor U29013 (N_29013,N_28496,N_28595);
xor U29014 (N_29014,N_28608,N_28897);
nand U29015 (N_29015,N_28638,N_28391);
xnor U29016 (N_29016,N_28921,N_28173);
xor U29017 (N_29017,N_28211,N_28484);
xor U29018 (N_29018,N_28039,N_28888);
or U29019 (N_29019,N_28596,N_28442);
and U29020 (N_29020,N_28277,N_28414);
nand U29021 (N_29021,N_28066,N_28042);
or U29022 (N_29022,N_28491,N_28507);
xor U29023 (N_29023,N_28091,N_28052);
xnor U29024 (N_29024,N_28453,N_28808);
xor U29025 (N_29025,N_28217,N_28165);
and U29026 (N_29026,N_28630,N_28196);
nand U29027 (N_29027,N_28986,N_28845);
nor U29028 (N_29028,N_28375,N_28138);
and U29029 (N_29029,N_28872,N_28376);
nand U29030 (N_29030,N_28299,N_28417);
and U29031 (N_29031,N_28623,N_28833);
xor U29032 (N_29032,N_28243,N_28092);
nand U29033 (N_29033,N_28169,N_28981);
or U29034 (N_29034,N_28641,N_28392);
xor U29035 (N_29035,N_28731,N_28818);
or U29036 (N_29036,N_28298,N_28756);
xnor U29037 (N_29037,N_28836,N_28191);
nor U29038 (N_29038,N_28755,N_28167);
nor U29039 (N_29039,N_28025,N_28995);
nand U29040 (N_29040,N_28743,N_28610);
nor U29041 (N_29041,N_28830,N_28010);
xnor U29042 (N_29042,N_28552,N_28397);
and U29043 (N_29043,N_28401,N_28603);
xor U29044 (N_29044,N_28718,N_28395);
nor U29045 (N_29045,N_28604,N_28297);
nor U29046 (N_29046,N_28624,N_28103);
xor U29047 (N_29047,N_28148,N_28617);
xor U29048 (N_29048,N_28933,N_28330);
nor U29049 (N_29049,N_28855,N_28308);
nand U29050 (N_29050,N_28223,N_28478);
xnor U29051 (N_29051,N_28096,N_28162);
or U29052 (N_29052,N_28707,N_28904);
nand U29053 (N_29053,N_28652,N_28744);
and U29054 (N_29054,N_28027,N_28422);
nor U29055 (N_29055,N_28253,N_28141);
nor U29056 (N_29056,N_28254,N_28727);
nand U29057 (N_29057,N_28771,N_28321);
or U29058 (N_29058,N_28068,N_28002);
or U29059 (N_29059,N_28047,N_28016);
xnor U29060 (N_29060,N_28111,N_28980);
and U29061 (N_29061,N_28784,N_28877);
nand U29062 (N_29062,N_28806,N_28432);
or U29063 (N_29063,N_28046,N_28653);
xor U29064 (N_29064,N_28445,N_28267);
nand U29065 (N_29065,N_28816,N_28402);
xor U29066 (N_29066,N_28700,N_28945);
nand U29067 (N_29067,N_28155,N_28074);
nand U29068 (N_29068,N_28225,N_28991);
xor U29069 (N_29069,N_28544,N_28998);
xor U29070 (N_29070,N_28221,N_28740);
nand U29071 (N_29071,N_28671,N_28136);
nand U29072 (N_29072,N_28972,N_28334);
and U29073 (N_29073,N_28849,N_28714);
and U29074 (N_29074,N_28631,N_28661);
xor U29075 (N_29075,N_28423,N_28782);
and U29076 (N_29076,N_28748,N_28182);
or U29077 (N_29077,N_28017,N_28408);
and U29078 (N_29078,N_28149,N_28073);
or U29079 (N_29079,N_28911,N_28702);
nand U29080 (N_29080,N_28664,N_28372);
nand U29081 (N_29081,N_28870,N_28699);
nand U29082 (N_29082,N_28411,N_28809);
nand U29083 (N_29083,N_28795,N_28434);
or U29084 (N_29084,N_28576,N_28193);
xor U29085 (N_29085,N_28270,N_28464);
or U29086 (N_29086,N_28691,N_28900);
nand U29087 (N_29087,N_28914,N_28446);
xnor U29088 (N_29088,N_28222,N_28050);
and U29089 (N_29089,N_28110,N_28421);
nand U29090 (N_29090,N_28764,N_28465);
nand U29091 (N_29091,N_28515,N_28942);
nand U29092 (N_29092,N_28481,N_28118);
and U29093 (N_29093,N_28435,N_28257);
nor U29094 (N_29094,N_28909,N_28988);
nand U29095 (N_29095,N_28218,N_28710);
or U29096 (N_29096,N_28301,N_28529);
xnor U29097 (N_29097,N_28399,N_28085);
and U29098 (N_29098,N_28082,N_28412);
nor U29099 (N_29099,N_28394,N_28834);
or U29100 (N_29100,N_28679,N_28452);
nand U29101 (N_29101,N_28647,N_28662);
xnor U29102 (N_29102,N_28612,N_28997);
or U29103 (N_29103,N_28670,N_28498);
and U29104 (N_29104,N_28785,N_28711);
xnor U29105 (N_29105,N_28355,N_28677);
nor U29106 (N_29106,N_28393,N_28541);
nor U29107 (N_29107,N_28437,N_28163);
or U29108 (N_29108,N_28772,N_28956);
and U29109 (N_29109,N_28658,N_28593);
and U29110 (N_29110,N_28143,N_28494);
and U29111 (N_29111,N_28121,N_28789);
and U29112 (N_29112,N_28788,N_28485);
nand U29113 (N_29113,N_28466,N_28890);
nor U29114 (N_29114,N_28179,N_28255);
and U29115 (N_29115,N_28787,N_28007);
nand U29116 (N_29116,N_28918,N_28463);
or U29117 (N_29117,N_28347,N_28560);
and U29118 (N_29118,N_28689,N_28053);
nor U29119 (N_29119,N_28248,N_28850);
nor U29120 (N_29120,N_28455,N_28095);
nand U29121 (N_29121,N_28305,N_28116);
and U29122 (N_29122,N_28729,N_28793);
nand U29123 (N_29123,N_28746,N_28886);
or U29124 (N_29124,N_28356,N_28229);
nand U29125 (N_29125,N_28086,N_28587);
nor U29126 (N_29126,N_28528,N_28087);
xor U29127 (N_29127,N_28759,N_28589);
nand U29128 (N_29128,N_28965,N_28390);
nand U29129 (N_29129,N_28773,N_28917);
xnor U29130 (N_29130,N_28339,N_28758);
or U29131 (N_29131,N_28451,N_28135);
nor U29132 (N_29132,N_28471,N_28343);
and U29133 (N_29133,N_28561,N_28475);
nand U29134 (N_29134,N_28547,N_28480);
and U29135 (N_29135,N_28246,N_28693);
nor U29136 (N_29136,N_28558,N_28774);
xnor U29137 (N_29137,N_28197,N_28287);
or U29138 (N_29138,N_28366,N_28540);
nand U29139 (N_29139,N_28613,N_28205);
nand U29140 (N_29140,N_28504,N_28106);
and U29141 (N_29141,N_28724,N_28537);
xor U29142 (N_29142,N_28079,N_28611);
nor U29143 (N_29143,N_28049,N_28098);
xnor U29144 (N_29144,N_28635,N_28646);
xor U29145 (N_29145,N_28667,N_28265);
nor U29146 (N_29146,N_28012,N_28151);
nand U29147 (N_29147,N_28358,N_28654);
nor U29148 (N_29148,N_28987,N_28876);
xnor U29149 (N_29149,N_28508,N_28717);
nand U29150 (N_29150,N_28014,N_28230);
or U29151 (N_29151,N_28967,N_28913);
nand U29152 (N_29152,N_28949,N_28420);
nor U29153 (N_29153,N_28860,N_28260);
xor U29154 (N_29154,N_28499,N_28129);
and U29155 (N_29155,N_28869,N_28716);
or U29156 (N_29156,N_28770,N_28235);
xor U29157 (N_29157,N_28353,N_28227);
nand U29158 (N_29158,N_28682,N_28698);
and U29159 (N_29159,N_28418,N_28269);
xor U29160 (N_29160,N_28362,N_28814);
nor U29161 (N_29161,N_28524,N_28794);
xnor U29162 (N_29162,N_28977,N_28473);
nor U29163 (N_29163,N_28078,N_28331);
or U29164 (N_29164,N_28032,N_28684);
or U29165 (N_29165,N_28573,N_28634);
or U29166 (N_29166,N_28800,N_28365);
xor U29167 (N_29167,N_28309,N_28985);
and U29168 (N_29168,N_28999,N_28805);
nand U29169 (N_29169,N_28273,N_28447);
or U29170 (N_29170,N_28351,N_28288);
or U29171 (N_29171,N_28174,N_28368);
nand U29172 (N_29172,N_28268,N_28974);
or U29173 (N_29173,N_28363,N_28655);
xor U29174 (N_29174,N_28064,N_28577);
xor U29175 (N_29175,N_28796,N_28732);
xor U29176 (N_29176,N_28500,N_28206);
nor U29177 (N_29177,N_28530,N_28233);
nand U29178 (N_29178,N_28361,N_28370);
nand U29179 (N_29179,N_28345,N_28673);
nor U29180 (N_29180,N_28036,N_28152);
and U29181 (N_29181,N_28307,N_28685);
nand U29182 (N_29182,N_28113,N_28591);
or U29183 (N_29183,N_28648,N_28090);
or U29184 (N_29184,N_28578,N_28950);
or U29185 (N_29185,N_28492,N_28571);
and U29186 (N_29186,N_28033,N_28626);
or U29187 (N_29187,N_28030,N_28185);
and U29188 (N_29188,N_28512,N_28158);
nand U29189 (N_29189,N_28847,N_28164);
xnor U29190 (N_29190,N_28760,N_28848);
and U29191 (N_29191,N_28493,N_28409);
nor U29192 (N_29192,N_28168,N_28134);
and U29193 (N_29193,N_28943,N_28990);
nor U29194 (N_29194,N_28826,N_28386);
nand U29195 (N_29195,N_28346,N_28019);
nor U29196 (N_29196,N_28973,N_28031);
and U29197 (N_29197,N_28448,N_28958);
nand U29198 (N_29198,N_28340,N_28342);
nor U29199 (N_29199,N_28660,N_28767);
nor U29200 (N_29200,N_28857,N_28328);
nor U29201 (N_29201,N_28176,N_28837);
or U29202 (N_29202,N_28310,N_28088);
and U29203 (N_29203,N_28559,N_28632);
nor U29204 (N_29204,N_28278,N_28602);
nor U29205 (N_29205,N_28289,N_28831);
xor U29206 (N_29206,N_28879,N_28929);
nor U29207 (N_29207,N_28752,N_28215);
nor U29208 (N_29208,N_28332,N_28865);
nor U29209 (N_29209,N_28349,N_28966);
and U29210 (N_29210,N_28853,N_28201);
nand U29211 (N_29211,N_28864,N_28659);
or U29212 (N_29212,N_28359,N_28526);
and U29213 (N_29213,N_28780,N_28245);
nand U29214 (N_29214,N_28214,N_28145);
nand U29215 (N_29215,N_28107,N_28083);
nor U29216 (N_29216,N_28315,N_28244);
nor U29217 (N_29217,N_28543,N_28458);
and U29218 (N_29218,N_28615,N_28912);
nor U29219 (N_29219,N_28625,N_28542);
nor U29220 (N_29220,N_28013,N_28264);
nor U29221 (N_29221,N_28825,N_28114);
or U29222 (N_29222,N_28557,N_28124);
xnor U29223 (N_29223,N_28776,N_28675);
or U29224 (N_29224,N_28819,N_28266);
xnor U29225 (N_29225,N_28940,N_28804);
nor U29226 (N_29226,N_28583,N_28018);
nor U29227 (N_29227,N_28622,N_28548);
nor U29228 (N_29228,N_28198,N_28687);
and U29229 (N_29229,N_28069,N_28450);
nor U29230 (N_29230,N_28599,N_28004);
nand U29231 (N_29231,N_28226,N_28766);
xor U29232 (N_29232,N_28271,N_28666);
and U29233 (N_29233,N_28859,N_28275);
nand U29234 (N_29234,N_28621,N_28497);
nor U29235 (N_29235,N_28517,N_28505);
nor U29236 (N_29236,N_28735,N_28854);
nor U29237 (N_29237,N_28065,N_28817);
and U29238 (N_29238,N_28798,N_28482);
or U29239 (N_29239,N_28021,N_28204);
nor U29240 (N_29240,N_28590,N_28120);
or U29241 (N_29241,N_28020,N_28416);
and U29242 (N_29242,N_28938,N_28649);
or U29243 (N_29243,N_28713,N_28915);
nor U29244 (N_29244,N_28678,N_28778);
or U29245 (N_29245,N_28968,N_28150);
and U29246 (N_29246,N_28656,N_28436);
nand U29247 (N_29247,N_28348,N_28931);
and U29248 (N_29248,N_28585,N_28302);
nand U29249 (N_29249,N_28979,N_28026);
xnor U29250 (N_29250,N_28947,N_28754);
xnor U29251 (N_29251,N_28644,N_28285);
xnor U29252 (N_29252,N_28570,N_28381);
nand U29253 (N_29253,N_28304,N_28574);
and U29254 (N_29254,N_28170,N_28373);
nand U29255 (N_29255,N_28063,N_28133);
xor U29256 (N_29256,N_28868,N_28993);
nand U29257 (N_29257,N_28367,N_28650);
or U29258 (N_29258,N_28609,N_28629);
and U29259 (N_29259,N_28927,N_28829);
nand U29260 (N_29260,N_28194,N_28534);
or U29261 (N_29261,N_28300,N_28751);
or U29262 (N_29262,N_28156,N_28028);
xnor U29263 (N_29263,N_28140,N_28415);
nand U29264 (N_29264,N_28694,N_28186);
and U29265 (N_29265,N_28329,N_28384);
xnor U29266 (N_29266,N_28123,N_28127);
nor U29267 (N_29267,N_28856,N_28213);
xor U29268 (N_29268,N_28620,N_28430);
nor U29269 (N_29269,N_28606,N_28538);
or U29270 (N_29270,N_28044,N_28554);
xor U29271 (N_29271,N_28935,N_28601);
nand U29272 (N_29272,N_28252,N_28188);
xnor U29273 (N_29273,N_28290,N_28405);
or U29274 (N_29274,N_28954,N_28696);
nor U29275 (N_29275,N_28352,N_28022);
nor U29276 (N_29276,N_28531,N_28396);
and U29277 (N_29277,N_28584,N_28525);
nor U29278 (N_29278,N_28093,N_28467);
and U29279 (N_29279,N_28462,N_28688);
nor U29280 (N_29280,N_28040,N_28511);
nand U29281 (N_29281,N_28906,N_28075);
and U29282 (N_29282,N_28479,N_28487);
or U29283 (N_29283,N_28941,N_28011);
and U29284 (N_29284,N_28109,N_28383);
and U29285 (N_29285,N_28104,N_28535);
nand U29286 (N_29286,N_28468,N_28726);
xor U29287 (N_29287,N_28739,N_28317);
xor U29288 (N_29288,N_28338,N_28736);
xnor U29289 (N_29289,N_28628,N_28282);
or U29290 (N_29290,N_28490,N_28923);
or U29291 (N_29291,N_28592,N_28378);
xnor U29292 (N_29292,N_28477,N_28055);
nand U29293 (N_29293,N_28884,N_28841);
nand U29294 (N_29294,N_28210,N_28518);
and U29295 (N_29295,N_28240,N_28750);
nor U29296 (N_29296,N_28586,N_28874);
nand U29297 (N_29297,N_28902,N_28828);
or U29298 (N_29298,N_28761,N_28296);
nand U29299 (N_29299,N_28946,N_28749);
nand U29300 (N_29300,N_28089,N_28719);
or U29301 (N_29301,N_28720,N_28242);
xor U29302 (N_29302,N_28827,N_28216);
nand U29303 (N_29303,N_28371,N_28157);
or U29304 (N_29304,N_28431,N_28976);
or U29305 (N_29305,N_28400,N_28812);
nor U29306 (N_29306,N_28539,N_28891);
nor U29307 (N_29307,N_28322,N_28842);
and U29308 (N_29308,N_28180,N_28427);
or U29309 (N_29309,N_28051,N_28926);
xor U29310 (N_29310,N_28564,N_28283);
or U29311 (N_29311,N_28443,N_28100);
nand U29312 (N_29312,N_28821,N_28549);
nand U29313 (N_29313,N_28737,N_28896);
or U29314 (N_29314,N_28777,N_28994);
and U29315 (N_29315,N_28438,N_28035);
nor U29316 (N_29316,N_28212,N_28117);
nand U29317 (N_29317,N_28597,N_28080);
nor U29318 (N_29318,N_28311,N_28676);
xor U29319 (N_29319,N_28247,N_28144);
xor U29320 (N_29320,N_28324,N_28234);
nand U29321 (N_29321,N_28516,N_28130);
nor U29322 (N_29322,N_28503,N_28318);
and U29323 (N_29323,N_28284,N_28489);
and U29324 (N_29324,N_28272,N_28762);
xnor U29325 (N_29325,N_28892,N_28159);
nor U29326 (N_29326,N_28952,N_28721);
or U29327 (N_29327,N_28404,N_28619);
nand U29328 (N_29328,N_28429,N_28996);
nor U29329 (N_29329,N_28236,N_28637);
xnor U29330 (N_29330,N_28005,N_28108);
xor U29331 (N_29331,N_28824,N_28202);
nor U29332 (N_29332,N_28851,N_28439);
nand U29333 (N_29333,N_28276,N_28895);
nor U29334 (N_29334,N_28969,N_28887);
nand U29335 (N_29335,N_28779,N_28871);
nor U29336 (N_29336,N_28875,N_28286);
nor U29337 (N_29337,N_28344,N_28822);
and U29338 (N_29338,N_28757,N_28792);
xor U29339 (N_29339,N_28483,N_28861);
nand U29340 (N_29340,N_28775,N_28060);
and U29341 (N_29341,N_28459,N_28734);
or U29342 (N_29342,N_28295,N_28097);
xor U29343 (N_29343,N_28094,N_28146);
nand U29344 (N_29344,N_28820,N_28250);
and U29345 (N_29345,N_28815,N_28070);
or U29346 (N_29346,N_28697,N_28665);
and U29347 (N_29347,N_28034,N_28072);
nand U29348 (N_29348,N_28279,N_28708);
nand U29349 (N_29349,N_28605,N_28893);
and U29350 (N_29350,N_28259,N_28398);
nand U29351 (N_29351,N_28325,N_28651);
nor U29352 (N_29352,N_28843,N_28454);
nor U29353 (N_29353,N_28354,N_28799);
nand U29354 (N_29354,N_28992,N_28840);
xor U29355 (N_29355,N_28600,N_28192);
or U29356 (N_29356,N_28076,N_28939);
or U29357 (N_29357,N_28701,N_28115);
xnor U29358 (N_29358,N_28102,N_28963);
nor U29359 (N_29359,N_28880,N_28261);
nor U29360 (N_29360,N_28101,N_28388);
nor U29361 (N_29361,N_28633,N_28208);
nand U29362 (N_29362,N_28126,N_28738);
and U29363 (N_29363,N_28572,N_28533);
and U29364 (N_29364,N_28341,N_28907);
and U29365 (N_29365,N_28009,N_28955);
xor U29366 (N_29366,N_28061,N_28449);
and U29367 (N_29367,N_28195,N_28166);
and U29368 (N_29368,N_28071,N_28407);
and U29369 (N_29369,N_28209,N_28642);
nand U29370 (N_29370,N_28582,N_28723);
nor U29371 (N_29371,N_28580,N_28054);
and U29372 (N_29372,N_28566,N_28501);
nor U29373 (N_29373,N_28728,N_28618);
nor U29374 (N_29374,N_28228,N_28357);
xnor U29375 (N_29375,N_28374,N_28084);
xor U29376 (N_29376,N_28350,N_28335);
and U29377 (N_29377,N_28280,N_28137);
nand U29378 (N_29378,N_28327,N_28048);
and U29379 (N_29379,N_28813,N_28172);
and U29380 (N_29380,N_28569,N_28742);
nand U29381 (N_29381,N_28506,N_28041);
or U29382 (N_29382,N_28457,N_28781);
nor U29383 (N_29383,N_28669,N_28132);
and U29384 (N_29384,N_28262,N_28364);
or U29385 (N_29385,N_28128,N_28835);
nor U29386 (N_29386,N_28686,N_28695);
or U29387 (N_29387,N_28360,N_28765);
xnor U29388 (N_29388,N_28680,N_28241);
and U29389 (N_29389,N_28936,N_28062);
or U29390 (N_29390,N_28614,N_28232);
nor U29391 (N_29391,N_28369,N_28183);
nor U29392 (N_29392,N_28502,N_28419);
and U29393 (N_29393,N_28745,N_28249);
nor U29394 (N_29394,N_28811,N_28038);
nor U29395 (N_29395,N_28753,N_28099);
nor U29396 (N_29396,N_28389,N_28783);
xor U29397 (N_29397,N_28903,N_28703);
xor U29398 (N_29398,N_28444,N_28510);
xor U29399 (N_29399,N_28948,N_28486);
nand U29400 (N_29400,N_28239,N_28640);
and U29401 (N_29401,N_28153,N_28989);
and U29402 (N_29402,N_28177,N_28844);
xnor U29403 (N_29403,N_28220,N_28672);
nor U29404 (N_29404,N_28867,N_28930);
xor U29405 (N_29405,N_28058,N_28883);
xor U29406 (N_29406,N_28476,N_28521);
or U29407 (N_29407,N_28567,N_28953);
and U29408 (N_29408,N_28725,N_28692);
xnor U29409 (N_29409,N_28281,N_28919);
xnor U29410 (N_29410,N_28937,N_28668);
nand U29411 (N_29411,N_28741,N_28456);
or U29412 (N_29412,N_28568,N_28863);
and U29413 (N_29413,N_28527,N_28681);
xnor U29414 (N_29414,N_28003,N_28790);
or U29415 (N_29415,N_28433,N_28551);
nor U29416 (N_29416,N_28565,N_28077);
nor U29417 (N_29417,N_28460,N_28190);
or U29418 (N_29418,N_28056,N_28112);
nand U29419 (N_29419,N_28024,N_28553);
and U29420 (N_29420,N_28594,N_28978);
nor U29421 (N_29421,N_28067,N_28333);
xnor U29422 (N_29422,N_28984,N_28730);
nor U29423 (N_29423,N_28905,N_28519);
or U29424 (N_29424,N_28959,N_28488);
nand U29425 (N_29425,N_28410,N_28722);
nand U29426 (N_29426,N_28474,N_28294);
or U29427 (N_29427,N_28555,N_28881);
or U29428 (N_29428,N_28536,N_28171);
and U29429 (N_29429,N_28957,N_28832);
nor U29430 (N_29430,N_28181,N_28690);
or U29431 (N_29431,N_28175,N_28337);
xor U29432 (N_29432,N_28920,N_28461);
and U29433 (N_29433,N_28178,N_28291);
or U29434 (N_29434,N_28683,N_28323);
nand U29435 (N_29435,N_28643,N_28320);
xnor U29436 (N_29436,N_28961,N_28231);
nor U29437 (N_29437,N_28203,N_28899);
xor U29438 (N_29438,N_28440,N_28663);
or U29439 (N_29439,N_28403,N_28224);
nand U29440 (N_29440,N_28747,N_28575);
and U29441 (N_29441,N_28426,N_28803);
or U29442 (N_29442,N_28184,N_28982);
xnor U29443 (N_29443,N_28377,N_28607);
xnor U29444 (N_29444,N_28858,N_28975);
xor U29445 (N_29445,N_28081,N_28791);
nand U29446 (N_29446,N_28043,N_28562);
xor U29447 (N_29447,N_28704,N_28263);
nand U29448 (N_29448,N_28878,N_28105);
xnor U29449 (N_29449,N_28674,N_28316);
and U29450 (N_29450,N_28319,N_28910);
and U29451 (N_29451,N_28616,N_28015);
or U29452 (N_29452,N_28059,N_28520);
xnor U29453 (N_29453,N_28219,N_28706);
nor U29454 (N_29454,N_28885,N_28513);
xor U29455 (N_29455,N_28379,N_28581);
nor U29456 (N_29456,N_28908,N_28258);
nor U29457 (N_29457,N_28898,N_28951);
xor U29458 (N_29458,N_28769,N_28495);
nor U29459 (N_29459,N_28532,N_28029);
or U29460 (N_29460,N_28639,N_28944);
nor U29461 (N_29461,N_28802,N_28292);
nor U29462 (N_29462,N_28925,N_28514);
and U29463 (N_29463,N_28550,N_28000);
or U29464 (N_29464,N_28924,N_28971);
nand U29465 (N_29465,N_28901,N_28810);
xnor U29466 (N_29466,N_28509,N_28006);
nor U29467 (N_29467,N_28962,N_28932);
nand U29468 (N_29468,N_28147,N_28916);
xor U29469 (N_29469,N_28715,N_28807);
xor U29470 (N_29470,N_28797,N_28636);
nand U29471 (N_29471,N_28657,N_28314);
nand U29472 (N_29472,N_28469,N_28598);
and U29473 (N_29473,N_28627,N_28023);
nand U29474 (N_29474,N_28545,N_28312);
nor U29475 (N_29475,N_28385,N_28472);
nand U29476 (N_29476,N_28238,N_28189);
nor U29477 (N_29477,N_28326,N_28882);
xor U29478 (N_29478,N_28336,N_28142);
nor U29479 (N_29479,N_28139,N_28768);
nor U29480 (N_29480,N_28251,N_28428);
or U29481 (N_29481,N_28122,N_28523);
nand U29482 (N_29482,N_28846,N_28934);
nand U29483 (N_29483,N_28862,N_28645);
or U29484 (N_29484,N_28588,N_28763);
nor U29485 (N_29485,N_28008,N_28838);
and U29486 (N_29486,N_28387,N_28256);
or U29487 (N_29487,N_28928,N_28786);
and U29488 (N_29488,N_28380,N_28866);
or U29489 (N_29489,N_28045,N_28894);
or U29490 (N_29490,N_28274,N_28413);
and U29491 (N_29491,N_28852,N_28293);
nand U29492 (N_29492,N_28001,N_28839);
nor U29493 (N_29493,N_28964,N_28382);
and U29494 (N_29494,N_28199,N_28733);
or U29495 (N_29495,N_28889,N_28154);
xnor U29496 (N_29496,N_28709,N_28237);
nand U29497 (N_29497,N_28160,N_28579);
nand U29498 (N_29498,N_28441,N_28970);
or U29499 (N_29499,N_28119,N_28556);
nor U29500 (N_29500,N_28448,N_28766);
xnor U29501 (N_29501,N_28668,N_28174);
and U29502 (N_29502,N_28187,N_28021);
xnor U29503 (N_29503,N_28299,N_28618);
nand U29504 (N_29504,N_28035,N_28810);
xor U29505 (N_29505,N_28042,N_28972);
and U29506 (N_29506,N_28208,N_28163);
and U29507 (N_29507,N_28343,N_28125);
nor U29508 (N_29508,N_28555,N_28788);
nor U29509 (N_29509,N_28629,N_28645);
xnor U29510 (N_29510,N_28868,N_28194);
and U29511 (N_29511,N_28331,N_28200);
nand U29512 (N_29512,N_28305,N_28185);
xor U29513 (N_29513,N_28288,N_28776);
xor U29514 (N_29514,N_28501,N_28806);
or U29515 (N_29515,N_28966,N_28023);
or U29516 (N_29516,N_28339,N_28178);
and U29517 (N_29517,N_28977,N_28382);
xnor U29518 (N_29518,N_28111,N_28501);
nor U29519 (N_29519,N_28712,N_28211);
or U29520 (N_29520,N_28477,N_28937);
and U29521 (N_29521,N_28151,N_28545);
nor U29522 (N_29522,N_28378,N_28905);
and U29523 (N_29523,N_28547,N_28018);
nand U29524 (N_29524,N_28477,N_28387);
and U29525 (N_29525,N_28529,N_28878);
nand U29526 (N_29526,N_28411,N_28368);
or U29527 (N_29527,N_28558,N_28598);
xor U29528 (N_29528,N_28134,N_28343);
nor U29529 (N_29529,N_28757,N_28627);
nand U29530 (N_29530,N_28188,N_28793);
and U29531 (N_29531,N_28796,N_28902);
nor U29532 (N_29532,N_28851,N_28639);
or U29533 (N_29533,N_28968,N_28751);
and U29534 (N_29534,N_28286,N_28970);
nor U29535 (N_29535,N_28099,N_28644);
or U29536 (N_29536,N_28173,N_28113);
xor U29537 (N_29537,N_28208,N_28852);
or U29538 (N_29538,N_28406,N_28074);
and U29539 (N_29539,N_28237,N_28674);
and U29540 (N_29540,N_28138,N_28880);
nor U29541 (N_29541,N_28138,N_28295);
and U29542 (N_29542,N_28054,N_28118);
and U29543 (N_29543,N_28329,N_28182);
nand U29544 (N_29544,N_28272,N_28402);
nor U29545 (N_29545,N_28780,N_28611);
nand U29546 (N_29546,N_28578,N_28876);
or U29547 (N_29547,N_28745,N_28401);
xor U29548 (N_29548,N_28326,N_28848);
nand U29549 (N_29549,N_28432,N_28976);
nor U29550 (N_29550,N_28017,N_28500);
nor U29551 (N_29551,N_28630,N_28346);
nand U29552 (N_29552,N_28828,N_28884);
nand U29553 (N_29553,N_28003,N_28387);
and U29554 (N_29554,N_28196,N_28473);
xor U29555 (N_29555,N_28806,N_28206);
and U29556 (N_29556,N_28611,N_28213);
nand U29557 (N_29557,N_28898,N_28080);
or U29558 (N_29558,N_28648,N_28888);
and U29559 (N_29559,N_28460,N_28077);
xnor U29560 (N_29560,N_28366,N_28719);
nand U29561 (N_29561,N_28356,N_28075);
nor U29562 (N_29562,N_28808,N_28730);
xnor U29563 (N_29563,N_28000,N_28914);
nor U29564 (N_29564,N_28838,N_28942);
and U29565 (N_29565,N_28615,N_28128);
and U29566 (N_29566,N_28687,N_28287);
xor U29567 (N_29567,N_28948,N_28272);
or U29568 (N_29568,N_28202,N_28497);
xnor U29569 (N_29569,N_28940,N_28933);
and U29570 (N_29570,N_28615,N_28400);
or U29571 (N_29571,N_28049,N_28213);
or U29572 (N_29572,N_28534,N_28461);
nand U29573 (N_29573,N_28832,N_28439);
nand U29574 (N_29574,N_28944,N_28259);
nor U29575 (N_29575,N_28819,N_28749);
nand U29576 (N_29576,N_28580,N_28266);
xnor U29577 (N_29577,N_28739,N_28253);
nand U29578 (N_29578,N_28511,N_28572);
nor U29579 (N_29579,N_28954,N_28834);
or U29580 (N_29580,N_28845,N_28247);
xnor U29581 (N_29581,N_28142,N_28282);
xnor U29582 (N_29582,N_28562,N_28811);
nand U29583 (N_29583,N_28273,N_28551);
nand U29584 (N_29584,N_28078,N_28830);
nor U29585 (N_29585,N_28253,N_28913);
or U29586 (N_29586,N_28815,N_28936);
xor U29587 (N_29587,N_28890,N_28066);
nand U29588 (N_29588,N_28726,N_28883);
or U29589 (N_29589,N_28215,N_28926);
or U29590 (N_29590,N_28953,N_28614);
and U29591 (N_29591,N_28708,N_28331);
nor U29592 (N_29592,N_28154,N_28749);
and U29593 (N_29593,N_28129,N_28613);
xor U29594 (N_29594,N_28048,N_28835);
and U29595 (N_29595,N_28855,N_28742);
nand U29596 (N_29596,N_28342,N_28315);
nor U29597 (N_29597,N_28833,N_28314);
nand U29598 (N_29598,N_28858,N_28451);
xor U29599 (N_29599,N_28013,N_28135);
or U29600 (N_29600,N_28594,N_28200);
or U29601 (N_29601,N_28779,N_28824);
nor U29602 (N_29602,N_28176,N_28371);
nor U29603 (N_29603,N_28179,N_28764);
nand U29604 (N_29604,N_28917,N_28315);
nand U29605 (N_29605,N_28285,N_28635);
or U29606 (N_29606,N_28478,N_28636);
nand U29607 (N_29607,N_28413,N_28285);
xor U29608 (N_29608,N_28596,N_28429);
and U29609 (N_29609,N_28434,N_28526);
and U29610 (N_29610,N_28331,N_28608);
xor U29611 (N_29611,N_28526,N_28680);
xnor U29612 (N_29612,N_28560,N_28209);
nand U29613 (N_29613,N_28324,N_28008);
and U29614 (N_29614,N_28020,N_28904);
or U29615 (N_29615,N_28064,N_28467);
or U29616 (N_29616,N_28404,N_28193);
nand U29617 (N_29617,N_28739,N_28676);
xnor U29618 (N_29618,N_28765,N_28679);
nor U29619 (N_29619,N_28032,N_28127);
xnor U29620 (N_29620,N_28194,N_28296);
xor U29621 (N_29621,N_28869,N_28312);
nand U29622 (N_29622,N_28638,N_28777);
xor U29623 (N_29623,N_28196,N_28339);
xor U29624 (N_29624,N_28045,N_28381);
nand U29625 (N_29625,N_28228,N_28258);
nor U29626 (N_29626,N_28951,N_28335);
and U29627 (N_29627,N_28412,N_28100);
nor U29628 (N_29628,N_28279,N_28937);
nor U29629 (N_29629,N_28338,N_28291);
xnor U29630 (N_29630,N_28639,N_28398);
or U29631 (N_29631,N_28792,N_28204);
nand U29632 (N_29632,N_28333,N_28990);
or U29633 (N_29633,N_28567,N_28397);
xnor U29634 (N_29634,N_28067,N_28034);
and U29635 (N_29635,N_28817,N_28337);
nor U29636 (N_29636,N_28638,N_28987);
xor U29637 (N_29637,N_28145,N_28852);
nor U29638 (N_29638,N_28938,N_28643);
nor U29639 (N_29639,N_28877,N_28837);
and U29640 (N_29640,N_28610,N_28307);
nand U29641 (N_29641,N_28858,N_28389);
xor U29642 (N_29642,N_28881,N_28675);
and U29643 (N_29643,N_28616,N_28174);
or U29644 (N_29644,N_28638,N_28282);
and U29645 (N_29645,N_28896,N_28099);
and U29646 (N_29646,N_28042,N_28523);
and U29647 (N_29647,N_28485,N_28653);
xor U29648 (N_29648,N_28452,N_28082);
or U29649 (N_29649,N_28501,N_28897);
or U29650 (N_29650,N_28542,N_28154);
and U29651 (N_29651,N_28574,N_28861);
xnor U29652 (N_29652,N_28458,N_28792);
or U29653 (N_29653,N_28380,N_28412);
and U29654 (N_29654,N_28555,N_28469);
and U29655 (N_29655,N_28563,N_28255);
nor U29656 (N_29656,N_28162,N_28631);
xor U29657 (N_29657,N_28517,N_28602);
or U29658 (N_29658,N_28116,N_28119);
xnor U29659 (N_29659,N_28169,N_28126);
and U29660 (N_29660,N_28606,N_28689);
or U29661 (N_29661,N_28017,N_28617);
xnor U29662 (N_29662,N_28044,N_28568);
nand U29663 (N_29663,N_28761,N_28981);
xnor U29664 (N_29664,N_28827,N_28067);
nor U29665 (N_29665,N_28748,N_28185);
xor U29666 (N_29666,N_28318,N_28429);
or U29667 (N_29667,N_28415,N_28677);
nor U29668 (N_29668,N_28205,N_28176);
xnor U29669 (N_29669,N_28448,N_28618);
and U29670 (N_29670,N_28759,N_28739);
xnor U29671 (N_29671,N_28385,N_28749);
nand U29672 (N_29672,N_28454,N_28211);
nand U29673 (N_29673,N_28128,N_28131);
nor U29674 (N_29674,N_28326,N_28625);
xnor U29675 (N_29675,N_28834,N_28115);
or U29676 (N_29676,N_28057,N_28973);
or U29677 (N_29677,N_28269,N_28836);
and U29678 (N_29678,N_28950,N_28972);
nor U29679 (N_29679,N_28902,N_28473);
xor U29680 (N_29680,N_28989,N_28373);
nor U29681 (N_29681,N_28859,N_28337);
and U29682 (N_29682,N_28029,N_28254);
nor U29683 (N_29683,N_28274,N_28155);
or U29684 (N_29684,N_28735,N_28920);
and U29685 (N_29685,N_28314,N_28720);
and U29686 (N_29686,N_28575,N_28015);
xor U29687 (N_29687,N_28365,N_28515);
xnor U29688 (N_29688,N_28227,N_28015);
xnor U29689 (N_29689,N_28331,N_28260);
nor U29690 (N_29690,N_28376,N_28944);
or U29691 (N_29691,N_28077,N_28266);
and U29692 (N_29692,N_28760,N_28212);
nor U29693 (N_29693,N_28767,N_28005);
and U29694 (N_29694,N_28079,N_28912);
nor U29695 (N_29695,N_28533,N_28853);
or U29696 (N_29696,N_28601,N_28246);
or U29697 (N_29697,N_28242,N_28127);
or U29698 (N_29698,N_28993,N_28625);
nand U29699 (N_29699,N_28585,N_28209);
xor U29700 (N_29700,N_28401,N_28064);
xnor U29701 (N_29701,N_28204,N_28209);
xnor U29702 (N_29702,N_28946,N_28150);
xnor U29703 (N_29703,N_28608,N_28449);
nand U29704 (N_29704,N_28144,N_28886);
or U29705 (N_29705,N_28434,N_28145);
or U29706 (N_29706,N_28845,N_28144);
xor U29707 (N_29707,N_28957,N_28082);
nor U29708 (N_29708,N_28762,N_28425);
and U29709 (N_29709,N_28706,N_28393);
or U29710 (N_29710,N_28577,N_28928);
and U29711 (N_29711,N_28682,N_28441);
and U29712 (N_29712,N_28864,N_28204);
or U29713 (N_29713,N_28907,N_28653);
nor U29714 (N_29714,N_28292,N_28655);
nor U29715 (N_29715,N_28666,N_28481);
and U29716 (N_29716,N_28275,N_28100);
nand U29717 (N_29717,N_28697,N_28888);
nand U29718 (N_29718,N_28260,N_28196);
xor U29719 (N_29719,N_28046,N_28770);
nand U29720 (N_29720,N_28518,N_28552);
or U29721 (N_29721,N_28345,N_28661);
and U29722 (N_29722,N_28240,N_28833);
xor U29723 (N_29723,N_28684,N_28224);
xnor U29724 (N_29724,N_28378,N_28081);
and U29725 (N_29725,N_28373,N_28121);
nand U29726 (N_29726,N_28985,N_28338);
nand U29727 (N_29727,N_28511,N_28148);
nor U29728 (N_29728,N_28562,N_28127);
xnor U29729 (N_29729,N_28170,N_28838);
and U29730 (N_29730,N_28669,N_28605);
nor U29731 (N_29731,N_28150,N_28516);
nand U29732 (N_29732,N_28767,N_28965);
or U29733 (N_29733,N_28058,N_28596);
nor U29734 (N_29734,N_28580,N_28761);
nor U29735 (N_29735,N_28287,N_28474);
nand U29736 (N_29736,N_28592,N_28761);
or U29737 (N_29737,N_28286,N_28613);
nand U29738 (N_29738,N_28226,N_28495);
xnor U29739 (N_29739,N_28423,N_28273);
or U29740 (N_29740,N_28672,N_28408);
xnor U29741 (N_29741,N_28044,N_28111);
or U29742 (N_29742,N_28060,N_28520);
nor U29743 (N_29743,N_28717,N_28534);
nand U29744 (N_29744,N_28109,N_28290);
nor U29745 (N_29745,N_28190,N_28142);
nor U29746 (N_29746,N_28609,N_28340);
or U29747 (N_29747,N_28439,N_28914);
and U29748 (N_29748,N_28717,N_28912);
nand U29749 (N_29749,N_28614,N_28196);
or U29750 (N_29750,N_28724,N_28388);
and U29751 (N_29751,N_28227,N_28702);
xnor U29752 (N_29752,N_28709,N_28190);
or U29753 (N_29753,N_28965,N_28201);
nand U29754 (N_29754,N_28975,N_28877);
and U29755 (N_29755,N_28326,N_28853);
xnor U29756 (N_29756,N_28030,N_28022);
nand U29757 (N_29757,N_28249,N_28317);
xor U29758 (N_29758,N_28904,N_28329);
xnor U29759 (N_29759,N_28600,N_28911);
and U29760 (N_29760,N_28575,N_28436);
nand U29761 (N_29761,N_28971,N_28992);
and U29762 (N_29762,N_28778,N_28691);
or U29763 (N_29763,N_28836,N_28421);
nor U29764 (N_29764,N_28247,N_28479);
xnor U29765 (N_29765,N_28638,N_28677);
xor U29766 (N_29766,N_28246,N_28426);
and U29767 (N_29767,N_28837,N_28654);
xnor U29768 (N_29768,N_28334,N_28427);
xor U29769 (N_29769,N_28007,N_28857);
or U29770 (N_29770,N_28653,N_28657);
and U29771 (N_29771,N_28999,N_28670);
or U29772 (N_29772,N_28065,N_28788);
nand U29773 (N_29773,N_28933,N_28904);
nand U29774 (N_29774,N_28202,N_28915);
xor U29775 (N_29775,N_28568,N_28163);
nor U29776 (N_29776,N_28790,N_28231);
and U29777 (N_29777,N_28651,N_28874);
nand U29778 (N_29778,N_28628,N_28213);
nand U29779 (N_29779,N_28672,N_28625);
and U29780 (N_29780,N_28860,N_28225);
nor U29781 (N_29781,N_28019,N_28349);
nor U29782 (N_29782,N_28637,N_28113);
and U29783 (N_29783,N_28135,N_28448);
nor U29784 (N_29784,N_28262,N_28500);
and U29785 (N_29785,N_28409,N_28426);
and U29786 (N_29786,N_28848,N_28822);
or U29787 (N_29787,N_28641,N_28151);
or U29788 (N_29788,N_28151,N_28181);
nor U29789 (N_29789,N_28987,N_28325);
and U29790 (N_29790,N_28598,N_28100);
and U29791 (N_29791,N_28374,N_28631);
nor U29792 (N_29792,N_28274,N_28546);
nor U29793 (N_29793,N_28311,N_28191);
xor U29794 (N_29794,N_28498,N_28798);
xor U29795 (N_29795,N_28686,N_28415);
or U29796 (N_29796,N_28571,N_28895);
and U29797 (N_29797,N_28439,N_28078);
nand U29798 (N_29798,N_28831,N_28629);
and U29799 (N_29799,N_28606,N_28566);
xnor U29800 (N_29800,N_28353,N_28388);
and U29801 (N_29801,N_28142,N_28502);
nor U29802 (N_29802,N_28758,N_28646);
xnor U29803 (N_29803,N_28628,N_28515);
xnor U29804 (N_29804,N_28311,N_28129);
xor U29805 (N_29805,N_28194,N_28843);
xnor U29806 (N_29806,N_28433,N_28084);
xor U29807 (N_29807,N_28255,N_28913);
xor U29808 (N_29808,N_28902,N_28885);
or U29809 (N_29809,N_28165,N_28019);
nand U29810 (N_29810,N_28888,N_28060);
nand U29811 (N_29811,N_28852,N_28529);
nand U29812 (N_29812,N_28252,N_28957);
and U29813 (N_29813,N_28278,N_28869);
nand U29814 (N_29814,N_28355,N_28005);
and U29815 (N_29815,N_28808,N_28872);
nor U29816 (N_29816,N_28975,N_28404);
or U29817 (N_29817,N_28953,N_28906);
nand U29818 (N_29818,N_28506,N_28826);
and U29819 (N_29819,N_28943,N_28186);
or U29820 (N_29820,N_28999,N_28119);
or U29821 (N_29821,N_28526,N_28820);
nand U29822 (N_29822,N_28145,N_28265);
nor U29823 (N_29823,N_28161,N_28856);
xnor U29824 (N_29824,N_28901,N_28958);
and U29825 (N_29825,N_28459,N_28237);
xor U29826 (N_29826,N_28696,N_28515);
xor U29827 (N_29827,N_28932,N_28426);
nand U29828 (N_29828,N_28161,N_28325);
nand U29829 (N_29829,N_28314,N_28060);
or U29830 (N_29830,N_28003,N_28621);
and U29831 (N_29831,N_28014,N_28579);
xor U29832 (N_29832,N_28364,N_28674);
nand U29833 (N_29833,N_28113,N_28199);
xnor U29834 (N_29834,N_28785,N_28805);
or U29835 (N_29835,N_28130,N_28909);
or U29836 (N_29836,N_28682,N_28713);
nor U29837 (N_29837,N_28124,N_28105);
nor U29838 (N_29838,N_28898,N_28429);
nor U29839 (N_29839,N_28859,N_28452);
nand U29840 (N_29840,N_28420,N_28208);
nand U29841 (N_29841,N_28651,N_28520);
nand U29842 (N_29842,N_28427,N_28020);
nand U29843 (N_29843,N_28000,N_28800);
and U29844 (N_29844,N_28234,N_28618);
or U29845 (N_29845,N_28331,N_28102);
nor U29846 (N_29846,N_28382,N_28457);
nor U29847 (N_29847,N_28439,N_28674);
or U29848 (N_29848,N_28663,N_28165);
or U29849 (N_29849,N_28034,N_28798);
or U29850 (N_29850,N_28842,N_28073);
xnor U29851 (N_29851,N_28288,N_28215);
nand U29852 (N_29852,N_28934,N_28633);
or U29853 (N_29853,N_28510,N_28473);
and U29854 (N_29854,N_28150,N_28325);
nor U29855 (N_29855,N_28115,N_28438);
xor U29856 (N_29856,N_28385,N_28712);
xor U29857 (N_29857,N_28642,N_28610);
nand U29858 (N_29858,N_28907,N_28329);
nor U29859 (N_29859,N_28766,N_28480);
xor U29860 (N_29860,N_28295,N_28568);
nand U29861 (N_29861,N_28441,N_28156);
nor U29862 (N_29862,N_28017,N_28495);
nor U29863 (N_29863,N_28924,N_28041);
xor U29864 (N_29864,N_28265,N_28548);
and U29865 (N_29865,N_28041,N_28989);
and U29866 (N_29866,N_28452,N_28089);
nand U29867 (N_29867,N_28299,N_28414);
nor U29868 (N_29868,N_28362,N_28636);
and U29869 (N_29869,N_28296,N_28067);
xnor U29870 (N_29870,N_28995,N_28074);
nor U29871 (N_29871,N_28912,N_28610);
nor U29872 (N_29872,N_28738,N_28015);
xor U29873 (N_29873,N_28068,N_28213);
or U29874 (N_29874,N_28746,N_28161);
xor U29875 (N_29875,N_28930,N_28048);
xor U29876 (N_29876,N_28944,N_28453);
nor U29877 (N_29877,N_28424,N_28355);
or U29878 (N_29878,N_28437,N_28927);
xor U29879 (N_29879,N_28170,N_28930);
or U29880 (N_29880,N_28498,N_28195);
xor U29881 (N_29881,N_28734,N_28307);
xor U29882 (N_29882,N_28371,N_28727);
nor U29883 (N_29883,N_28278,N_28501);
and U29884 (N_29884,N_28139,N_28958);
nor U29885 (N_29885,N_28863,N_28784);
nand U29886 (N_29886,N_28831,N_28358);
nand U29887 (N_29887,N_28592,N_28040);
and U29888 (N_29888,N_28041,N_28527);
nand U29889 (N_29889,N_28400,N_28937);
or U29890 (N_29890,N_28481,N_28075);
or U29891 (N_29891,N_28866,N_28062);
nor U29892 (N_29892,N_28883,N_28494);
nor U29893 (N_29893,N_28214,N_28462);
or U29894 (N_29894,N_28696,N_28924);
xor U29895 (N_29895,N_28845,N_28079);
nor U29896 (N_29896,N_28158,N_28209);
nand U29897 (N_29897,N_28466,N_28090);
nor U29898 (N_29898,N_28791,N_28645);
nor U29899 (N_29899,N_28545,N_28621);
nor U29900 (N_29900,N_28329,N_28203);
or U29901 (N_29901,N_28592,N_28984);
nor U29902 (N_29902,N_28941,N_28602);
nand U29903 (N_29903,N_28879,N_28384);
and U29904 (N_29904,N_28557,N_28695);
nor U29905 (N_29905,N_28189,N_28842);
xor U29906 (N_29906,N_28079,N_28052);
xor U29907 (N_29907,N_28892,N_28470);
nand U29908 (N_29908,N_28310,N_28251);
nand U29909 (N_29909,N_28158,N_28948);
or U29910 (N_29910,N_28929,N_28994);
nand U29911 (N_29911,N_28840,N_28000);
and U29912 (N_29912,N_28484,N_28116);
and U29913 (N_29913,N_28912,N_28580);
or U29914 (N_29914,N_28524,N_28473);
nor U29915 (N_29915,N_28423,N_28165);
nand U29916 (N_29916,N_28122,N_28575);
or U29917 (N_29917,N_28563,N_28655);
and U29918 (N_29918,N_28128,N_28428);
nor U29919 (N_29919,N_28501,N_28738);
xor U29920 (N_29920,N_28333,N_28496);
and U29921 (N_29921,N_28540,N_28430);
and U29922 (N_29922,N_28387,N_28604);
xnor U29923 (N_29923,N_28440,N_28775);
or U29924 (N_29924,N_28190,N_28001);
xor U29925 (N_29925,N_28444,N_28491);
and U29926 (N_29926,N_28020,N_28103);
and U29927 (N_29927,N_28845,N_28778);
nand U29928 (N_29928,N_28653,N_28102);
xor U29929 (N_29929,N_28257,N_28720);
xor U29930 (N_29930,N_28301,N_28099);
nand U29931 (N_29931,N_28727,N_28305);
xnor U29932 (N_29932,N_28960,N_28524);
and U29933 (N_29933,N_28595,N_28361);
nor U29934 (N_29934,N_28085,N_28577);
xor U29935 (N_29935,N_28904,N_28274);
nand U29936 (N_29936,N_28544,N_28970);
xnor U29937 (N_29937,N_28069,N_28433);
xor U29938 (N_29938,N_28417,N_28895);
or U29939 (N_29939,N_28253,N_28262);
xnor U29940 (N_29940,N_28665,N_28860);
and U29941 (N_29941,N_28996,N_28711);
nand U29942 (N_29942,N_28951,N_28185);
nand U29943 (N_29943,N_28939,N_28003);
xnor U29944 (N_29944,N_28648,N_28698);
and U29945 (N_29945,N_28705,N_28889);
or U29946 (N_29946,N_28828,N_28236);
xor U29947 (N_29947,N_28871,N_28455);
nand U29948 (N_29948,N_28481,N_28039);
nand U29949 (N_29949,N_28543,N_28183);
nor U29950 (N_29950,N_28981,N_28724);
xnor U29951 (N_29951,N_28743,N_28788);
and U29952 (N_29952,N_28743,N_28760);
or U29953 (N_29953,N_28737,N_28125);
nor U29954 (N_29954,N_28976,N_28157);
nor U29955 (N_29955,N_28570,N_28188);
and U29956 (N_29956,N_28666,N_28097);
nand U29957 (N_29957,N_28643,N_28248);
or U29958 (N_29958,N_28624,N_28510);
and U29959 (N_29959,N_28825,N_28563);
nor U29960 (N_29960,N_28809,N_28229);
xnor U29961 (N_29961,N_28959,N_28883);
nor U29962 (N_29962,N_28187,N_28794);
xor U29963 (N_29963,N_28917,N_28782);
nand U29964 (N_29964,N_28460,N_28158);
xnor U29965 (N_29965,N_28771,N_28261);
nand U29966 (N_29966,N_28954,N_28894);
or U29967 (N_29967,N_28465,N_28217);
and U29968 (N_29968,N_28212,N_28944);
xor U29969 (N_29969,N_28569,N_28914);
or U29970 (N_29970,N_28150,N_28681);
and U29971 (N_29971,N_28890,N_28364);
or U29972 (N_29972,N_28586,N_28392);
nand U29973 (N_29973,N_28809,N_28100);
xnor U29974 (N_29974,N_28459,N_28472);
nor U29975 (N_29975,N_28235,N_28523);
and U29976 (N_29976,N_28362,N_28732);
nand U29977 (N_29977,N_28495,N_28253);
and U29978 (N_29978,N_28060,N_28948);
nand U29979 (N_29979,N_28677,N_28437);
or U29980 (N_29980,N_28096,N_28899);
nor U29981 (N_29981,N_28466,N_28722);
and U29982 (N_29982,N_28125,N_28623);
nand U29983 (N_29983,N_28050,N_28034);
and U29984 (N_29984,N_28597,N_28392);
or U29985 (N_29985,N_28933,N_28993);
and U29986 (N_29986,N_28927,N_28234);
xor U29987 (N_29987,N_28255,N_28831);
xor U29988 (N_29988,N_28073,N_28345);
xor U29989 (N_29989,N_28489,N_28714);
nand U29990 (N_29990,N_28846,N_28792);
xor U29991 (N_29991,N_28957,N_28821);
nor U29992 (N_29992,N_28505,N_28052);
xor U29993 (N_29993,N_28779,N_28240);
nand U29994 (N_29994,N_28832,N_28417);
or U29995 (N_29995,N_28485,N_28869);
xnor U29996 (N_29996,N_28636,N_28329);
xnor U29997 (N_29997,N_28099,N_28100);
xnor U29998 (N_29998,N_28338,N_28022);
or U29999 (N_29999,N_28937,N_28543);
or U30000 (N_30000,N_29562,N_29694);
nor U30001 (N_30001,N_29351,N_29388);
nand U30002 (N_30002,N_29407,N_29802);
nor U30003 (N_30003,N_29534,N_29746);
or U30004 (N_30004,N_29137,N_29197);
nor U30005 (N_30005,N_29069,N_29902);
xor U30006 (N_30006,N_29289,N_29028);
and U30007 (N_30007,N_29195,N_29477);
or U30008 (N_30008,N_29501,N_29699);
and U30009 (N_30009,N_29352,N_29659);
xnor U30010 (N_30010,N_29359,N_29913);
nand U30011 (N_30011,N_29241,N_29267);
nor U30012 (N_30012,N_29758,N_29506);
nor U30013 (N_30013,N_29532,N_29492);
and U30014 (N_30014,N_29148,N_29441);
and U30015 (N_30015,N_29608,N_29291);
xnor U30016 (N_30016,N_29507,N_29414);
nand U30017 (N_30017,N_29191,N_29718);
and U30018 (N_30018,N_29033,N_29225);
and U30019 (N_30019,N_29838,N_29223);
or U30020 (N_30020,N_29049,N_29382);
xnor U30021 (N_30021,N_29229,N_29383);
and U30022 (N_30022,N_29164,N_29323);
nand U30023 (N_30023,N_29811,N_29543);
xor U30024 (N_30024,N_29607,N_29252);
nand U30025 (N_30025,N_29023,N_29194);
nor U30026 (N_30026,N_29186,N_29064);
or U30027 (N_30027,N_29832,N_29431);
nor U30028 (N_30028,N_29960,N_29258);
or U30029 (N_30029,N_29588,N_29944);
xor U30030 (N_30030,N_29379,N_29867);
nand U30031 (N_30031,N_29039,N_29785);
xor U30032 (N_30032,N_29560,N_29862);
nand U30033 (N_30033,N_29423,N_29417);
or U30034 (N_30034,N_29858,N_29278);
nor U30035 (N_30035,N_29146,N_29226);
xnor U30036 (N_30036,N_29422,N_29539);
and U30037 (N_30037,N_29956,N_29232);
nand U30038 (N_30038,N_29974,N_29181);
nand U30039 (N_30039,N_29579,N_29502);
or U30040 (N_30040,N_29962,N_29798);
nor U30041 (N_30041,N_29985,N_29932);
or U30042 (N_30042,N_29580,N_29171);
nor U30043 (N_30043,N_29903,N_29337);
xor U30044 (N_30044,N_29312,N_29533);
and U30045 (N_30045,N_29888,N_29854);
and U30046 (N_30046,N_29037,N_29819);
nand U30047 (N_30047,N_29822,N_29676);
xor U30048 (N_30048,N_29602,N_29056);
xnor U30049 (N_30049,N_29322,N_29150);
nor U30050 (N_30050,N_29106,N_29524);
nand U30051 (N_30051,N_29619,N_29459);
xor U30052 (N_30052,N_29749,N_29405);
xnor U30053 (N_30053,N_29935,N_29839);
or U30054 (N_30054,N_29736,N_29724);
and U30055 (N_30055,N_29347,N_29270);
and U30056 (N_30056,N_29683,N_29961);
xnor U30057 (N_30057,N_29329,N_29376);
nor U30058 (N_30058,N_29889,N_29713);
nand U30059 (N_30059,N_29666,N_29178);
xor U30060 (N_30060,N_29308,N_29877);
xor U30061 (N_30061,N_29470,N_29964);
and U30062 (N_30062,N_29705,N_29034);
nor U30063 (N_30063,N_29016,N_29269);
and U30064 (N_30064,N_29615,N_29440);
or U30065 (N_30065,N_29170,N_29429);
xor U30066 (N_30066,N_29552,N_29314);
or U30067 (N_30067,N_29192,N_29404);
and U30068 (N_30068,N_29018,N_29793);
nand U30069 (N_30069,N_29138,N_29499);
nor U30070 (N_30070,N_29936,N_29795);
nand U30071 (N_30071,N_29378,N_29456);
xnor U30072 (N_30072,N_29331,N_29045);
nand U30073 (N_30073,N_29915,N_29344);
nor U30074 (N_30074,N_29693,N_29397);
nor U30075 (N_30075,N_29717,N_29887);
and U30076 (N_30076,N_29824,N_29630);
nor U30077 (N_30077,N_29024,N_29471);
xor U30078 (N_30078,N_29756,N_29846);
or U30079 (N_30079,N_29450,N_29516);
or U30080 (N_30080,N_29334,N_29131);
or U30081 (N_30081,N_29398,N_29276);
and U30082 (N_30082,N_29409,N_29430);
nor U30083 (N_30083,N_29255,N_29317);
xor U30084 (N_30084,N_29467,N_29361);
nor U30085 (N_30085,N_29975,N_29777);
and U30086 (N_30086,N_29074,N_29006);
nand U30087 (N_30087,N_29592,N_29446);
nor U30088 (N_30088,N_29239,N_29906);
nor U30089 (N_30089,N_29771,N_29894);
and U30090 (N_30090,N_29628,N_29301);
and U30091 (N_30091,N_29432,N_29940);
xnor U30092 (N_30092,N_29814,N_29859);
or U30093 (N_30093,N_29380,N_29061);
and U30094 (N_30094,N_29973,N_29554);
or U30095 (N_30095,N_29408,N_29399);
nand U30096 (N_30096,N_29556,N_29685);
or U30097 (N_30097,N_29110,N_29221);
nor U30098 (N_30098,N_29385,N_29618);
nand U30099 (N_30099,N_29062,N_29410);
or U30100 (N_30100,N_29078,N_29265);
nor U30101 (N_30101,N_29236,N_29969);
nor U30102 (N_30102,N_29548,N_29230);
or U30103 (N_30103,N_29466,N_29884);
and U30104 (N_30104,N_29157,N_29369);
xnor U30105 (N_30105,N_29797,N_29967);
or U30106 (N_30106,N_29848,N_29711);
and U30107 (N_30107,N_29594,N_29886);
nor U30108 (N_30108,N_29104,N_29261);
or U30109 (N_30109,N_29368,N_29480);
nand U30110 (N_30110,N_29327,N_29752);
nand U30111 (N_30111,N_29463,N_29719);
xor U30112 (N_30112,N_29143,N_29631);
nand U30113 (N_30113,N_29183,N_29864);
nand U30114 (N_30114,N_29773,N_29803);
nand U30115 (N_30115,N_29710,N_29203);
xnor U30116 (N_30116,N_29122,N_29675);
and U30117 (N_30117,N_29306,N_29402);
and U30118 (N_30118,N_29916,N_29545);
or U30119 (N_30119,N_29836,N_29790);
nand U30120 (N_30120,N_29395,N_29165);
nand U30121 (N_30121,N_29792,N_29521);
nand U30122 (N_30122,N_29680,N_29815);
nor U30123 (N_30123,N_29870,N_29907);
nor U30124 (N_30124,N_29294,N_29500);
nor U30125 (N_30125,N_29387,N_29584);
nand U30126 (N_30126,N_29831,N_29332);
nor U30127 (N_30127,N_29875,N_29233);
nand U30128 (N_30128,N_29072,N_29005);
or U30129 (N_30129,N_29564,N_29338);
xor U30130 (N_30130,N_29610,N_29652);
xor U30131 (N_30131,N_29498,N_29511);
and U30132 (N_30132,N_29707,N_29517);
nand U30133 (N_30133,N_29527,N_29739);
nor U30134 (N_30134,N_29412,N_29144);
xnor U30135 (N_30135,N_29198,N_29257);
xnor U30136 (N_30136,N_29966,N_29504);
xnor U30137 (N_30137,N_29476,N_29159);
xor U30138 (N_30138,N_29085,N_29857);
nand U30139 (N_30139,N_29460,N_29433);
and U30140 (N_30140,N_29212,N_29162);
xnor U30141 (N_30141,N_29179,N_29883);
or U30142 (N_30142,N_29125,N_29780);
nand U30143 (N_30143,N_29420,N_29097);
nand U30144 (N_30144,N_29860,N_29763);
and U30145 (N_30145,N_29978,N_29977);
or U30146 (N_30146,N_29931,N_29003);
nand U30147 (N_30147,N_29950,N_29597);
nor U30148 (N_30148,N_29565,N_29211);
nor U30149 (N_30149,N_29572,N_29546);
or U30150 (N_30150,N_29885,N_29434);
xor U30151 (N_30151,N_29172,N_29288);
and U30152 (N_30152,N_29114,N_29734);
xnor U30153 (N_30153,N_29362,N_29720);
nor U30154 (N_30154,N_29520,N_29928);
nor U30155 (N_30155,N_29444,N_29447);
xor U30156 (N_30156,N_29919,N_29304);
nand U30157 (N_30157,N_29817,N_29508);
nor U30158 (N_30158,N_29356,N_29243);
or U30159 (N_30159,N_29394,N_29140);
xor U30160 (N_30160,N_29868,N_29712);
or U30161 (N_30161,N_29000,N_29567);
nor U30162 (N_30162,N_29954,N_29569);
xor U30163 (N_30163,N_29677,N_29462);
or U30164 (N_30164,N_29904,N_29672);
or U30165 (N_30165,N_29601,N_29593);
and U30166 (N_30166,N_29249,N_29073);
nand U30167 (N_30167,N_29353,N_29644);
nor U30168 (N_30168,N_29514,N_29899);
xnor U30169 (N_30169,N_29551,N_29706);
nor U30170 (N_30170,N_29829,N_29156);
and U30171 (N_30171,N_29363,N_29390);
xor U30172 (N_30172,N_29939,N_29094);
nand U30173 (N_30173,N_29487,N_29266);
xnor U30174 (N_30174,N_29737,N_29367);
and U30175 (N_30175,N_29059,N_29806);
and U30176 (N_30176,N_29897,N_29934);
nor U30177 (N_30177,N_29090,N_29174);
nand U30178 (N_30178,N_29577,N_29244);
xnor U30179 (N_30179,N_29365,N_29808);
nand U30180 (N_30180,N_29688,N_29188);
and U30181 (N_30181,N_29151,N_29264);
nand U30182 (N_30182,N_29823,N_29512);
and U30183 (N_30183,N_29496,N_29438);
xor U30184 (N_30184,N_29624,N_29871);
and U30185 (N_30185,N_29340,N_29224);
nor U30186 (N_30186,N_29687,N_29099);
nor U30187 (N_30187,N_29484,N_29299);
nor U30188 (N_30188,N_29645,N_29637);
xor U30189 (N_30189,N_29210,N_29494);
xnor U30190 (N_30190,N_29972,N_29290);
nand U30191 (N_30191,N_29287,N_29284);
nor U30192 (N_30192,N_29566,N_29686);
nor U30193 (N_30193,N_29425,N_29008);
nand U30194 (N_30194,N_29598,N_29155);
and U30195 (N_30195,N_29336,N_29891);
and U30196 (N_30196,N_29482,N_29286);
xor U30197 (N_30197,N_29735,N_29012);
xnor U30198 (N_30198,N_29472,N_29640);
or U30199 (N_30199,N_29704,N_29297);
xnor U30200 (N_30200,N_29120,N_29537);
and U30201 (N_30201,N_29757,N_29483);
nand U30202 (N_30202,N_29994,N_29816);
or U30203 (N_30203,N_29949,N_29561);
and U30204 (N_30204,N_29358,N_29614);
nand U30205 (N_30205,N_29318,N_29851);
xor U30206 (N_30206,N_29055,N_29127);
or U30207 (N_30207,N_29855,N_29673);
nand U30208 (N_30208,N_29182,N_29493);
nor U30209 (N_30209,N_29136,N_29922);
nor U30210 (N_30210,N_29419,N_29648);
or U30211 (N_30211,N_29540,N_29963);
and U30212 (N_30212,N_29957,N_29842);
xnor U30213 (N_30213,N_29087,N_29166);
nor U30214 (N_30214,N_29600,N_29001);
nor U30215 (N_30215,N_29464,N_29307);
or U30216 (N_30216,N_29530,N_29636);
and U30217 (N_30217,N_29830,N_29701);
or U30218 (N_30218,N_29599,N_29914);
nand U30219 (N_30219,N_29998,N_29669);
nand U30220 (N_30220,N_29054,N_29947);
nand U30221 (N_30221,N_29945,N_29519);
nand U30222 (N_30222,N_29247,N_29568);
nor U30223 (N_30223,N_29050,N_29981);
nand U30224 (N_30224,N_29925,N_29702);
xnor U30225 (N_30225,N_29733,N_29818);
nor U30226 (N_30226,N_29727,N_29285);
or U30227 (N_30227,N_29215,N_29523);
xor U30228 (N_30228,N_29726,N_29918);
and U30229 (N_30229,N_29077,N_29202);
xnor U30230 (N_30230,N_29133,N_29794);
nand U30231 (N_30231,N_29346,N_29730);
or U30232 (N_30232,N_29841,N_29373);
nor U30233 (N_30233,N_29542,N_29279);
nand U30234 (N_30234,N_29696,N_29253);
xnor U30235 (N_30235,N_29242,N_29199);
or U30236 (N_30236,N_29176,N_29684);
nor U30237 (N_30237,N_29789,N_29315);
nor U30238 (N_30238,N_29582,N_29139);
or U30239 (N_30239,N_29910,N_29457);
nor U30240 (N_30240,N_29117,N_29043);
xnor U30241 (N_30241,N_29449,N_29873);
nor U30242 (N_30242,N_29112,N_29142);
or U30243 (N_30243,N_29465,N_29098);
xnor U30244 (N_30244,N_29679,N_29213);
and U30245 (N_30245,N_29262,N_29128);
nand U30246 (N_30246,N_29990,N_29435);
and U30247 (N_30247,N_29651,N_29744);
nor U30248 (N_30248,N_29053,N_29088);
and U30249 (N_30249,N_29850,N_29130);
nand U30250 (N_30250,N_29153,N_29451);
nand U30251 (N_30251,N_29065,N_29901);
and U30252 (N_30252,N_29513,N_29031);
xnor U30253 (N_30253,N_29107,N_29427);
xnor U30254 (N_30254,N_29671,N_29013);
or U30255 (N_30255,N_29011,N_29703);
and U30256 (N_30256,N_29075,N_29189);
nor U30257 (N_30257,N_29999,N_29807);
or U30258 (N_30258,N_29782,N_29812);
nor U30259 (N_30259,N_29313,N_29436);
nor U30260 (N_30260,N_29827,N_29118);
and U30261 (N_30261,N_29204,N_29102);
and U30262 (N_30262,N_29987,N_29613);
or U30263 (N_30263,N_29218,N_29282);
nor U30264 (N_30264,N_29759,N_29788);
nand U30265 (N_30265,N_29946,N_29277);
xnor U30266 (N_30266,N_29765,N_29660);
nand U30267 (N_30267,N_29691,N_29019);
or U30268 (N_30268,N_29762,N_29665);
nor U30269 (N_30269,N_29141,N_29917);
nor U30270 (N_30270,N_29207,N_29926);
nor U30271 (N_30271,N_29856,N_29081);
or U30272 (N_30272,N_29661,N_29145);
nor U30273 (N_30273,N_29428,N_29343);
or U30274 (N_30274,N_29052,N_29058);
xnor U30275 (N_30275,N_29168,N_29769);
or U30276 (N_30276,N_29035,N_29784);
nand U30277 (N_30277,N_29820,N_29559);
or U30278 (N_30278,N_29214,N_29324);
or U30279 (N_30279,N_29022,N_29587);
xnor U30280 (N_30280,N_29689,N_29124);
nor U30281 (N_30281,N_29032,N_29080);
nand U30282 (N_30282,N_29263,N_29796);
and U30283 (N_30283,N_29834,N_29905);
nor U30284 (N_30284,N_29046,N_29132);
xnor U30285 (N_30285,N_29386,N_29027);
nand U30286 (N_30286,N_29030,N_29595);
nor U30287 (N_30287,N_29938,N_29256);
and U30288 (N_30288,N_29360,N_29246);
xnor U30289 (N_30289,N_29861,N_29729);
and U30290 (N_30290,N_29007,N_29259);
and U30291 (N_30291,N_29840,N_29623);
and U30292 (N_30292,N_29646,N_29892);
or U30293 (N_30293,N_29632,N_29328);
nor U30294 (N_30294,N_29716,N_29103);
nand U30295 (N_30295,N_29021,N_29206);
or U30296 (N_30296,N_29180,N_29201);
nand U30297 (N_30297,N_29714,N_29955);
xor U30298 (N_30298,N_29590,N_29424);
nor U30299 (N_30299,N_29874,N_29863);
nand U30300 (N_30300,N_29774,N_29400);
nand U30301 (N_30301,N_29895,N_29952);
xnor U30302 (N_30302,N_29538,N_29237);
and U30303 (N_30303,N_29478,N_29578);
nand U30304 (N_30304,N_29510,N_29020);
nor U30305 (N_30305,N_29108,N_29093);
and U30306 (N_30306,N_29657,N_29654);
and U30307 (N_30307,N_29017,N_29800);
nand U30308 (N_30308,N_29647,N_29416);
nor U30309 (N_30309,N_29929,N_29339);
nor U30310 (N_30310,N_29461,N_29219);
or U30311 (N_30311,N_29292,N_29042);
nand U30312 (N_30312,N_29603,N_29709);
xor U30313 (N_30313,N_29234,N_29574);
or U30314 (N_30314,N_29573,N_29240);
xor U30315 (N_30315,N_29555,N_29341);
nor U30316 (N_30316,N_29943,N_29750);
or U30317 (N_30317,N_29531,N_29937);
or U30318 (N_30318,N_29779,N_29448);
nor U30319 (N_30319,N_29682,N_29876);
or U30320 (N_30320,N_29082,N_29616);
or U30321 (N_30321,N_29222,N_29366);
nand U30322 (N_30322,N_29541,N_29649);
nor U30323 (N_30323,N_29326,N_29123);
nor U30324 (N_30324,N_29515,N_29029);
and U30325 (N_30325,N_29325,N_29342);
and U30326 (N_30326,N_29528,N_29813);
nand U30327 (N_30327,N_29664,N_29695);
nor U30328 (N_30328,N_29604,N_29828);
xor U30329 (N_30329,N_29298,N_29674);
nor U30330 (N_30330,N_29272,N_29333);
xor U30331 (N_30331,N_29173,N_29129);
and U30332 (N_30332,N_29479,N_29621);
or U30333 (N_30333,N_29575,N_29804);
and U30334 (N_30334,N_29731,N_29633);
nor U30335 (N_30335,N_29335,N_29658);
nand U30336 (N_30336,N_29303,N_29505);
and U30337 (N_30337,N_29583,N_29473);
and U30338 (N_30338,N_29389,N_29992);
or U30339 (N_30339,N_29100,N_29205);
nand U30340 (N_30340,N_29475,N_29909);
and U30341 (N_30341,N_29025,N_29890);
nand U30342 (N_30342,N_29445,N_29767);
and U30343 (N_30343,N_29634,N_29134);
or U30344 (N_30344,N_29160,N_29079);
or U30345 (N_30345,N_29866,N_29743);
and U30346 (N_30346,N_29921,N_29535);
nand U30347 (N_30347,N_29766,N_29667);
and U30348 (N_30348,N_29778,N_29349);
or U30349 (N_30349,N_29522,N_29437);
or U30350 (N_30350,N_29837,N_29606);
and U30351 (N_30351,N_29948,N_29576);
nor U30352 (N_30352,N_29439,N_29670);
nor U30353 (N_30353,N_29260,N_29912);
nor U30354 (N_30354,N_29489,N_29852);
and U30355 (N_30355,N_29930,N_29791);
nand U30356 (N_30356,N_29865,N_29070);
and U30357 (N_30357,N_29549,N_29725);
nand U30358 (N_30358,N_29849,N_29115);
nor U30359 (N_30359,N_29585,N_29642);
nor U30360 (N_30360,N_29663,N_29959);
xor U30361 (N_30361,N_29989,N_29655);
and U30362 (N_30362,N_29067,N_29968);
and U30363 (N_30363,N_29825,N_29495);
nand U30364 (N_30364,N_29392,N_29776);
and U30365 (N_30365,N_29754,N_29638);
or U30366 (N_30366,N_29163,N_29063);
nand U30367 (N_30367,N_29760,N_29089);
nor U30368 (N_30368,N_29620,N_29497);
or U30369 (N_30369,N_29452,N_29896);
xor U30370 (N_30370,N_29413,N_29997);
and U30371 (N_30371,N_29415,N_29311);
nor U30372 (N_30372,N_29271,N_29982);
and U30373 (N_30373,N_29933,N_29217);
and U30374 (N_30374,N_29309,N_29544);
nand U30375 (N_30375,N_29845,N_29996);
nand U30376 (N_30376,N_29485,N_29971);
and U30377 (N_30377,N_29988,N_29668);
and U30378 (N_30378,N_29200,N_29442);
nor U30379 (N_30379,N_29723,N_29557);
xnor U30380 (N_30380,N_29503,N_29563);
nand U30381 (N_30381,N_29167,N_29844);
nand U30382 (N_30382,N_29348,N_29426);
or U30383 (N_30383,N_29721,N_29458);
and U30384 (N_30384,N_29391,N_29364);
nand U30385 (N_30385,N_29740,N_29152);
and U30386 (N_30386,N_29810,N_29208);
nor U30387 (N_30387,N_29051,N_29722);
nor U30388 (N_30388,N_29612,N_29293);
or U30389 (N_30389,N_29320,N_29553);
or U30390 (N_30390,N_29095,N_29036);
or U30391 (N_30391,N_29228,N_29635);
nand U30392 (N_30392,N_29396,N_29154);
and U30393 (N_30393,N_29040,N_29443);
nor U30394 (N_30394,N_29923,N_29653);
xnor U30395 (N_30395,N_29591,N_29371);
or U30396 (N_30396,N_29741,N_29372);
nor U30397 (N_30397,N_29662,N_29609);
nand U30398 (N_30398,N_29084,N_29627);
or U30399 (N_30399,N_29274,N_29786);
xor U30400 (N_30400,N_29126,N_29295);
and U30401 (N_30401,N_29980,N_29009);
nand U30402 (N_30402,N_29302,N_29586);
nand U30403 (N_30403,N_29418,N_29281);
and U30404 (N_30404,N_29015,N_29403);
nor U30405 (N_30405,N_29105,N_29715);
xor U30406 (N_30406,N_29625,N_29014);
or U30407 (N_30407,N_29526,N_29924);
xnor U30408 (N_30408,N_29490,N_29374);
or U30409 (N_30409,N_29571,N_29421);
nor U30410 (N_30410,N_29393,N_29066);
xor U30411 (N_30411,N_29781,N_29927);
xor U30412 (N_30412,N_29193,N_29622);
nor U30413 (N_30413,N_29958,N_29345);
nor U30414 (N_30414,N_29872,N_29469);
nor U30415 (N_30415,N_29908,N_29384);
or U30416 (N_30416,N_29488,N_29639);
or U30417 (N_30417,N_29184,N_29708);
and U30418 (N_30418,N_29690,N_29250);
xnor U30419 (N_30419,N_29251,N_29091);
nor U30420 (N_30420,N_29231,N_29805);
and U30421 (N_30421,N_29216,N_29799);
nand U30422 (N_30422,N_29570,N_29847);
nand U30423 (N_30423,N_29377,N_29355);
nor U30424 (N_30424,N_29026,N_29190);
xor U30425 (N_30425,N_29698,N_29509);
and U30426 (N_30426,N_29310,N_29581);
nor U30427 (N_30427,N_29738,N_29004);
or U30428 (N_30428,N_29518,N_29275);
and U30429 (N_30429,N_29911,N_29953);
and U30430 (N_30430,N_29745,N_29135);
nand U30431 (N_30431,N_29083,N_29678);
and U30432 (N_30432,N_29468,N_29991);
nand U30433 (N_30433,N_29254,N_29057);
xnor U30434 (N_30434,N_29942,N_29161);
xor U30435 (N_30435,N_29984,N_29536);
and U30436 (N_30436,N_29898,N_29406);
nor U30437 (N_30437,N_29280,N_29605);
nand U30438 (N_30438,N_29048,N_29986);
nand U30439 (N_30439,N_29761,N_29770);
xor U30440 (N_30440,N_29965,N_29976);
nand U30441 (N_30441,N_29900,N_29196);
nor U30442 (N_30442,N_29881,N_29656);
and U30443 (N_30443,N_29060,N_29177);
nand U30444 (N_30444,N_29751,N_29641);
nand U30445 (N_30445,N_29768,N_29357);
or U30446 (N_30446,N_29076,N_29092);
nand U30447 (N_30447,N_29038,N_29728);
and U30448 (N_30448,N_29316,N_29116);
nor U30449 (N_30449,N_29010,N_29697);
or U30450 (N_30450,N_29617,N_29983);
xor U30451 (N_30451,N_29121,N_29227);
or U30452 (N_30452,N_29330,N_29764);
nand U30453 (N_30453,N_29300,N_29611);
xnor U30454 (N_30454,N_29629,N_29273);
and U30455 (N_30455,N_29558,N_29732);
or U30456 (N_30456,N_29550,N_29835);
and U30457 (N_30457,N_29350,N_29086);
nand U30458 (N_30458,N_29354,N_29755);
xnor U30459 (N_30459,N_29993,N_29941);
nand U30460 (N_30460,N_29772,N_29596);
or U30461 (N_30461,N_29650,N_29375);
and U30462 (N_30462,N_29296,N_29692);
and U30463 (N_30463,N_29821,N_29893);
nand U30464 (N_30464,N_29748,N_29455);
and U30465 (N_30465,N_29589,N_29370);
or U30466 (N_30466,N_29319,N_29843);
or U30467 (N_30467,N_29175,N_29169);
xor U30468 (N_30468,N_29185,N_29486);
nor U30469 (N_30469,N_29970,N_29809);
and U30470 (N_30470,N_29833,N_29381);
and U30471 (N_30471,N_29096,N_29305);
nor U30472 (N_30472,N_29979,N_29547);
nor U30473 (N_30473,N_29041,N_29109);
and U30474 (N_30474,N_29700,N_29113);
or U30475 (N_30475,N_29826,N_29783);
nand U30476 (N_30476,N_29787,N_29742);
nor U30477 (N_30477,N_29491,N_29853);
and U30478 (N_30478,N_29220,N_29283);
nor U30479 (N_30479,N_29878,N_29454);
nor U30480 (N_30480,N_29147,N_29995);
nor U30481 (N_30481,N_29071,N_29401);
and U30482 (N_30482,N_29111,N_29775);
and U30483 (N_30483,N_29474,N_29453);
and U30484 (N_30484,N_29068,N_29747);
nand U30485 (N_30485,N_29245,N_29481);
nor U30486 (N_30486,N_29951,N_29411);
or U30487 (N_30487,N_29187,N_29753);
xnor U30488 (N_30488,N_29119,N_29002);
and U30489 (N_30489,N_29880,N_29529);
and U30490 (N_30490,N_29643,N_29158);
xor U30491 (N_30491,N_29920,N_29801);
nand U30492 (N_30492,N_29681,N_29268);
nand U30493 (N_30493,N_29879,N_29321);
xnor U30494 (N_30494,N_29238,N_29047);
nand U30495 (N_30495,N_29882,N_29525);
xnor U30496 (N_30496,N_29209,N_29248);
nand U30497 (N_30497,N_29235,N_29044);
nand U30498 (N_30498,N_29101,N_29869);
nand U30499 (N_30499,N_29149,N_29626);
nor U30500 (N_30500,N_29179,N_29311);
and U30501 (N_30501,N_29864,N_29356);
nand U30502 (N_30502,N_29929,N_29208);
or U30503 (N_30503,N_29707,N_29067);
nor U30504 (N_30504,N_29080,N_29340);
xor U30505 (N_30505,N_29605,N_29340);
nor U30506 (N_30506,N_29052,N_29136);
or U30507 (N_30507,N_29328,N_29246);
nor U30508 (N_30508,N_29580,N_29977);
nor U30509 (N_30509,N_29354,N_29709);
and U30510 (N_30510,N_29043,N_29230);
xor U30511 (N_30511,N_29294,N_29767);
nand U30512 (N_30512,N_29114,N_29468);
nor U30513 (N_30513,N_29520,N_29647);
nand U30514 (N_30514,N_29667,N_29305);
xor U30515 (N_30515,N_29824,N_29864);
xnor U30516 (N_30516,N_29998,N_29074);
xor U30517 (N_30517,N_29262,N_29340);
or U30518 (N_30518,N_29586,N_29413);
nor U30519 (N_30519,N_29508,N_29045);
nand U30520 (N_30520,N_29797,N_29609);
or U30521 (N_30521,N_29978,N_29627);
xor U30522 (N_30522,N_29477,N_29598);
nand U30523 (N_30523,N_29924,N_29850);
nor U30524 (N_30524,N_29698,N_29180);
or U30525 (N_30525,N_29845,N_29241);
nand U30526 (N_30526,N_29233,N_29811);
xnor U30527 (N_30527,N_29691,N_29238);
nand U30528 (N_30528,N_29062,N_29046);
nand U30529 (N_30529,N_29276,N_29184);
nor U30530 (N_30530,N_29411,N_29682);
or U30531 (N_30531,N_29576,N_29179);
nand U30532 (N_30532,N_29898,N_29016);
nor U30533 (N_30533,N_29881,N_29122);
nor U30534 (N_30534,N_29156,N_29193);
nand U30535 (N_30535,N_29004,N_29111);
nor U30536 (N_30536,N_29959,N_29415);
xnor U30537 (N_30537,N_29009,N_29080);
and U30538 (N_30538,N_29592,N_29005);
xor U30539 (N_30539,N_29388,N_29496);
and U30540 (N_30540,N_29478,N_29239);
or U30541 (N_30541,N_29360,N_29100);
and U30542 (N_30542,N_29184,N_29254);
and U30543 (N_30543,N_29144,N_29633);
nand U30544 (N_30544,N_29120,N_29119);
and U30545 (N_30545,N_29226,N_29290);
nand U30546 (N_30546,N_29292,N_29655);
nor U30547 (N_30547,N_29946,N_29935);
or U30548 (N_30548,N_29237,N_29272);
or U30549 (N_30549,N_29925,N_29529);
and U30550 (N_30550,N_29008,N_29035);
xnor U30551 (N_30551,N_29623,N_29998);
and U30552 (N_30552,N_29016,N_29271);
nand U30553 (N_30553,N_29776,N_29397);
or U30554 (N_30554,N_29543,N_29460);
and U30555 (N_30555,N_29537,N_29037);
and U30556 (N_30556,N_29306,N_29149);
nor U30557 (N_30557,N_29625,N_29277);
nand U30558 (N_30558,N_29932,N_29566);
nand U30559 (N_30559,N_29681,N_29756);
or U30560 (N_30560,N_29054,N_29079);
and U30561 (N_30561,N_29810,N_29612);
or U30562 (N_30562,N_29697,N_29624);
or U30563 (N_30563,N_29657,N_29237);
xnor U30564 (N_30564,N_29173,N_29786);
or U30565 (N_30565,N_29330,N_29862);
and U30566 (N_30566,N_29960,N_29340);
xor U30567 (N_30567,N_29260,N_29784);
xor U30568 (N_30568,N_29732,N_29981);
nand U30569 (N_30569,N_29197,N_29997);
or U30570 (N_30570,N_29704,N_29423);
or U30571 (N_30571,N_29671,N_29679);
nor U30572 (N_30572,N_29862,N_29195);
xor U30573 (N_30573,N_29832,N_29383);
xnor U30574 (N_30574,N_29587,N_29028);
nor U30575 (N_30575,N_29373,N_29526);
nor U30576 (N_30576,N_29431,N_29446);
nand U30577 (N_30577,N_29675,N_29845);
or U30578 (N_30578,N_29022,N_29720);
or U30579 (N_30579,N_29839,N_29569);
nor U30580 (N_30580,N_29577,N_29347);
xnor U30581 (N_30581,N_29776,N_29327);
nor U30582 (N_30582,N_29324,N_29180);
nor U30583 (N_30583,N_29190,N_29767);
or U30584 (N_30584,N_29372,N_29966);
or U30585 (N_30585,N_29292,N_29174);
nor U30586 (N_30586,N_29311,N_29107);
nand U30587 (N_30587,N_29479,N_29008);
or U30588 (N_30588,N_29493,N_29396);
nor U30589 (N_30589,N_29246,N_29942);
or U30590 (N_30590,N_29520,N_29724);
nor U30591 (N_30591,N_29759,N_29821);
nor U30592 (N_30592,N_29477,N_29282);
xnor U30593 (N_30593,N_29240,N_29116);
nor U30594 (N_30594,N_29434,N_29930);
or U30595 (N_30595,N_29264,N_29738);
nor U30596 (N_30596,N_29794,N_29007);
nand U30597 (N_30597,N_29287,N_29113);
nor U30598 (N_30598,N_29186,N_29080);
and U30599 (N_30599,N_29032,N_29838);
nor U30600 (N_30600,N_29126,N_29768);
xnor U30601 (N_30601,N_29205,N_29996);
xnor U30602 (N_30602,N_29543,N_29727);
nand U30603 (N_30603,N_29721,N_29662);
nand U30604 (N_30604,N_29732,N_29352);
nand U30605 (N_30605,N_29042,N_29618);
nor U30606 (N_30606,N_29738,N_29586);
or U30607 (N_30607,N_29291,N_29744);
nand U30608 (N_30608,N_29223,N_29039);
xor U30609 (N_30609,N_29374,N_29551);
or U30610 (N_30610,N_29334,N_29358);
and U30611 (N_30611,N_29013,N_29479);
or U30612 (N_30612,N_29858,N_29180);
and U30613 (N_30613,N_29595,N_29223);
xnor U30614 (N_30614,N_29175,N_29624);
nor U30615 (N_30615,N_29273,N_29150);
nor U30616 (N_30616,N_29905,N_29375);
nor U30617 (N_30617,N_29727,N_29100);
and U30618 (N_30618,N_29385,N_29536);
xnor U30619 (N_30619,N_29421,N_29511);
nor U30620 (N_30620,N_29783,N_29386);
nor U30621 (N_30621,N_29792,N_29785);
or U30622 (N_30622,N_29959,N_29932);
nand U30623 (N_30623,N_29649,N_29291);
xnor U30624 (N_30624,N_29567,N_29992);
xnor U30625 (N_30625,N_29311,N_29229);
xor U30626 (N_30626,N_29287,N_29957);
and U30627 (N_30627,N_29999,N_29260);
nor U30628 (N_30628,N_29972,N_29181);
xnor U30629 (N_30629,N_29499,N_29769);
or U30630 (N_30630,N_29442,N_29910);
nand U30631 (N_30631,N_29221,N_29283);
nor U30632 (N_30632,N_29167,N_29939);
and U30633 (N_30633,N_29580,N_29652);
nor U30634 (N_30634,N_29741,N_29710);
or U30635 (N_30635,N_29629,N_29556);
or U30636 (N_30636,N_29680,N_29348);
xor U30637 (N_30637,N_29681,N_29912);
xnor U30638 (N_30638,N_29050,N_29124);
nor U30639 (N_30639,N_29297,N_29151);
nor U30640 (N_30640,N_29230,N_29799);
or U30641 (N_30641,N_29637,N_29105);
and U30642 (N_30642,N_29517,N_29639);
nand U30643 (N_30643,N_29571,N_29070);
xnor U30644 (N_30644,N_29684,N_29711);
and U30645 (N_30645,N_29390,N_29728);
nor U30646 (N_30646,N_29676,N_29351);
nand U30647 (N_30647,N_29463,N_29306);
nor U30648 (N_30648,N_29093,N_29106);
nand U30649 (N_30649,N_29152,N_29072);
xor U30650 (N_30650,N_29006,N_29930);
xor U30651 (N_30651,N_29746,N_29852);
nand U30652 (N_30652,N_29760,N_29104);
xor U30653 (N_30653,N_29198,N_29734);
or U30654 (N_30654,N_29463,N_29027);
xor U30655 (N_30655,N_29248,N_29726);
and U30656 (N_30656,N_29545,N_29979);
nor U30657 (N_30657,N_29438,N_29392);
or U30658 (N_30658,N_29227,N_29744);
and U30659 (N_30659,N_29857,N_29005);
xor U30660 (N_30660,N_29501,N_29225);
nand U30661 (N_30661,N_29222,N_29008);
or U30662 (N_30662,N_29223,N_29704);
xnor U30663 (N_30663,N_29657,N_29443);
nand U30664 (N_30664,N_29691,N_29854);
nand U30665 (N_30665,N_29207,N_29773);
and U30666 (N_30666,N_29664,N_29470);
and U30667 (N_30667,N_29672,N_29776);
nor U30668 (N_30668,N_29681,N_29495);
nand U30669 (N_30669,N_29692,N_29469);
xor U30670 (N_30670,N_29863,N_29292);
nand U30671 (N_30671,N_29554,N_29791);
xor U30672 (N_30672,N_29418,N_29848);
nor U30673 (N_30673,N_29198,N_29286);
xnor U30674 (N_30674,N_29020,N_29477);
nor U30675 (N_30675,N_29884,N_29732);
xor U30676 (N_30676,N_29981,N_29590);
nor U30677 (N_30677,N_29001,N_29020);
and U30678 (N_30678,N_29039,N_29177);
xor U30679 (N_30679,N_29562,N_29420);
and U30680 (N_30680,N_29513,N_29221);
nor U30681 (N_30681,N_29284,N_29355);
nor U30682 (N_30682,N_29662,N_29885);
nand U30683 (N_30683,N_29549,N_29919);
nand U30684 (N_30684,N_29542,N_29086);
or U30685 (N_30685,N_29212,N_29620);
xor U30686 (N_30686,N_29725,N_29399);
and U30687 (N_30687,N_29854,N_29923);
xnor U30688 (N_30688,N_29764,N_29401);
xnor U30689 (N_30689,N_29563,N_29746);
nand U30690 (N_30690,N_29286,N_29804);
and U30691 (N_30691,N_29454,N_29537);
and U30692 (N_30692,N_29771,N_29258);
nor U30693 (N_30693,N_29919,N_29186);
nand U30694 (N_30694,N_29509,N_29941);
xnor U30695 (N_30695,N_29228,N_29775);
nand U30696 (N_30696,N_29503,N_29659);
nand U30697 (N_30697,N_29118,N_29246);
xor U30698 (N_30698,N_29050,N_29811);
or U30699 (N_30699,N_29912,N_29208);
and U30700 (N_30700,N_29418,N_29884);
nor U30701 (N_30701,N_29667,N_29521);
and U30702 (N_30702,N_29549,N_29956);
xnor U30703 (N_30703,N_29079,N_29788);
or U30704 (N_30704,N_29324,N_29220);
nand U30705 (N_30705,N_29359,N_29574);
nand U30706 (N_30706,N_29564,N_29225);
nor U30707 (N_30707,N_29447,N_29007);
and U30708 (N_30708,N_29578,N_29741);
xor U30709 (N_30709,N_29163,N_29211);
xor U30710 (N_30710,N_29387,N_29943);
and U30711 (N_30711,N_29078,N_29108);
xnor U30712 (N_30712,N_29261,N_29941);
and U30713 (N_30713,N_29695,N_29250);
nand U30714 (N_30714,N_29783,N_29389);
xnor U30715 (N_30715,N_29514,N_29926);
nor U30716 (N_30716,N_29356,N_29086);
xor U30717 (N_30717,N_29760,N_29225);
nand U30718 (N_30718,N_29887,N_29755);
or U30719 (N_30719,N_29536,N_29277);
nor U30720 (N_30720,N_29868,N_29904);
nor U30721 (N_30721,N_29521,N_29465);
or U30722 (N_30722,N_29574,N_29057);
and U30723 (N_30723,N_29079,N_29777);
nor U30724 (N_30724,N_29655,N_29928);
nor U30725 (N_30725,N_29658,N_29042);
nor U30726 (N_30726,N_29158,N_29238);
and U30727 (N_30727,N_29547,N_29978);
nor U30728 (N_30728,N_29242,N_29195);
nand U30729 (N_30729,N_29594,N_29996);
nor U30730 (N_30730,N_29211,N_29779);
nand U30731 (N_30731,N_29089,N_29735);
and U30732 (N_30732,N_29015,N_29720);
xor U30733 (N_30733,N_29918,N_29078);
nand U30734 (N_30734,N_29440,N_29327);
nor U30735 (N_30735,N_29310,N_29748);
and U30736 (N_30736,N_29521,N_29793);
xnor U30737 (N_30737,N_29036,N_29649);
xor U30738 (N_30738,N_29329,N_29937);
nand U30739 (N_30739,N_29585,N_29837);
or U30740 (N_30740,N_29805,N_29017);
nor U30741 (N_30741,N_29102,N_29537);
nor U30742 (N_30742,N_29031,N_29989);
and U30743 (N_30743,N_29183,N_29218);
or U30744 (N_30744,N_29491,N_29495);
or U30745 (N_30745,N_29204,N_29303);
nand U30746 (N_30746,N_29494,N_29561);
or U30747 (N_30747,N_29545,N_29567);
nand U30748 (N_30748,N_29588,N_29860);
xor U30749 (N_30749,N_29871,N_29898);
or U30750 (N_30750,N_29121,N_29070);
and U30751 (N_30751,N_29771,N_29188);
and U30752 (N_30752,N_29864,N_29465);
nand U30753 (N_30753,N_29416,N_29855);
or U30754 (N_30754,N_29466,N_29477);
nor U30755 (N_30755,N_29668,N_29674);
nand U30756 (N_30756,N_29528,N_29124);
xnor U30757 (N_30757,N_29548,N_29703);
xnor U30758 (N_30758,N_29172,N_29024);
or U30759 (N_30759,N_29093,N_29985);
or U30760 (N_30760,N_29883,N_29063);
nand U30761 (N_30761,N_29305,N_29209);
xor U30762 (N_30762,N_29547,N_29329);
nand U30763 (N_30763,N_29548,N_29571);
nor U30764 (N_30764,N_29508,N_29052);
nor U30765 (N_30765,N_29957,N_29807);
and U30766 (N_30766,N_29010,N_29128);
and U30767 (N_30767,N_29244,N_29448);
xnor U30768 (N_30768,N_29630,N_29063);
nand U30769 (N_30769,N_29743,N_29868);
and U30770 (N_30770,N_29473,N_29940);
nor U30771 (N_30771,N_29640,N_29101);
nand U30772 (N_30772,N_29767,N_29512);
and U30773 (N_30773,N_29781,N_29879);
and U30774 (N_30774,N_29649,N_29683);
nand U30775 (N_30775,N_29753,N_29943);
or U30776 (N_30776,N_29248,N_29961);
and U30777 (N_30777,N_29907,N_29082);
or U30778 (N_30778,N_29248,N_29426);
nand U30779 (N_30779,N_29988,N_29933);
or U30780 (N_30780,N_29311,N_29769);
and U30781 (N_30781,N_29411,N_29352);
or U30782 (N_30782,N_29865,N_29048);
nor U30783 (N_30783,N_29316,N_29622);
xor U30784 (N_30784,N_29988,N_29119);
and U30785 (N_30785,N_29307,N_29207);
nor U30786 (N_30786,N_29265,N_29922);
nand U30787 (N_30787,N_29895,N_29431);
xor U30788 (N_30788,N_29761,N_29197);
or U30789 (N_30789,N_29505,N_29518);
or U30790 (N_30790,N_29517,N_29207);
and U30791 (N_30791,N_29388,N_29715);
nor U30792 (N_30792,N_29240,N_29514);
or U30793 (N_30793,N_29459,N_29307);
nor U30794 (N_30794,N_29301,N_29163);
and U30795 (N_30795,N_29659,N_29943);
nor U30796 (N_30796,N_29829,N_29637);
nand U30797 (N_30797,N_29356,N_29007);
or U30798 (N_30798,N_29612,N_29461);
or U30799 (N_30799,N_29969,N_29651);
nand U30800 (N_30800,N_29479,N_29857);
or U30801 (N_30801,N_29943,N_29217);
nor U30802 (N_30802,N_29892,N_29842);
nor U30803 (N_30803,N_29627,N_29439);
xor U30804 (N_30804,N_29987,N_29786);
and U30805 (N_30805,N_29979,N_29396);
nor U30806 (N_30806,N_29273,N_29604);
nor U30807 (N_30807,N_29056,N_29505);
nand U30808 (N_30808,N_29127,N_29534);
and U30809 (N_30809,N_29093,N_29993);
xnor U30810 (N_30810,N_29648,N_29099);
nand U30811 (N_30811,N_29362,N_29606);
xnor U30812 (N_30812,N_29616,N_29940);
or U30813 (N_30813,N_29910,N_29797);
nor U30814 (N_30814,N_29484,N_29951);
and U30815 (N_30815,N_29163,N_29828);
xor U30816 (N_30816,N_29955,N_29086);
xnor U30817 (N_30817,N_29588,N_29348);
nand U30818 (N_30818,N_29305,N_29499);
xnor U30819 (N_30819,N_29398,N_29155);
and U30820 (N_30820,N_29397,N_29329);
xor U30821 (N_30821,N_29099,N_29255);
nand U30822 (N_30822,N_29481,N_29836);
nor U30823 (N_30823,N_29424,N_29835);
nor U30824 (N_30824,N_29772,N_29696);
nor U30825 (N_30825,N_29167,N_29207);
xor U30826 (N_30826,N_29732,N_29515);
and U30827 (N_30827,N_29649,N_29932);
or U30828 (N_30828,N_29381,N_29459);
and U30829 (N_30829,N_29694,N_29459);
xnor U30830 (N_30830,N_29159,N_29402);
nor U30831 (N_30831,N_29784,N_29379);
nor U30832 (N_30832,N_29998,N_29515);
nor U30833 (N_30833,N_29781,N_29615);
nor U30834 (N_30834,N_29036,N_29895);
nor U30835 (N_30835,N_29514,N_29667);
and U30836 (N_30836,N_29314,N_29403);
or U30837 (N_30837,N_29344,N_29484);
or U30838 (N_30838,N_29469,N_29814);
xnor U30839 (N_30839,N_29183,N_29579);
and U30840 (N_30840,N_29776,N_29199);
nor U30841 (N_30841,N_29348,N_29415);
xnor U30842 (N_30842,N_29216,N_29466);
or U30843 (N_30843,N_29124,N_29393);
nand U30844 (N_30844,N_29236,N_29488);
nand U30845 (N_30845,N_29412,N_29125);
xor U30846 (N_30846,N_29959,N_29917);
and U30847 (N_30847,N_29589,N_29630);
and U30848 (N_30848,N_29854,N_29563);
xor U30849 (N_30849,N_29408,N_29441);
or U30850 (N_30850,N_29518,N_29492);
or U30851 (N_30851,N_29586,N_29669);
nor U30852 (N_30852,N_29983,N_29568);
xnor U30853 (N_30853,N_29107,N_29648);
and U30854 (N_30854,N_29791,N_29049);
xor U30855 (N_30855,N_29213,N_29765);
or U30856 (N_30856,N_29191,N_29374);
and U30857 (N_30857,N_29924,N_29546);
and U30858 (N_30858,N_29811,N_29114);
nand U30859 (N_30859,N_29677,N_29927);
nor U30860 (N_30860,N_29782,N_29847);
nand U30861 (N_30861,N_29226,N_29038);
nor U30862 (N_30862,N_29945,N_29203);
nor U30863 (N_30863,N_29125,N_29761);
xor U30864 (N_30864,N_29000,N_29379);
or U30865 (N_30865,N_29571,N_29193);
nand U30866 (N_30866,N_29550,N_29859);
and U30867 (N_30867,N_29137,N_29998);
xor U30868 (N_30868,N_29664,N_29810);
nor U30869 (N_30869,N_29796,N_29440);
and U30870 (N_30870,N_29178,N_29660);
nand U30871 (N_30871,N_29759,N_29436);
nand U30872 (N_30872,N_29712,N_29690);
and U30873 (N_30873,N_29636,N_29109);
or U30874 (N_30874,N_29243,N_29058);
nor U30875 (N_30875,N_29828,N_29807);
and U30876 (N_30876,N_29374,N_29787);
and U30877 (N_30877,N_29066,N_29222);
nand U30878 (N_30878,N_29194,N_29995);
xnor U30879 (N_30879,N_29719,N_29649);
nor U30880 (N_30880,N_29579,N_29967);
and U30881 (N_30881,N_29352,N_29275);
xnor U30882 (N_30882,N_29834,N_29692);
xnor U30883 (N_30883,N_29949,N_29126);
xor U30884 (N_30884,N_29186,N_29035);
nand U30885 (N_30885,N_29905,N_29389);
or U30886 (N_30886,N_29900,N_29510);
or U30887 (N_30887,N_29216,N_29606);
or U30888 (N_30888,N_29498,N_29460);
and U30889 (N_30889,N_29654,N_29971);
and U30890 (N_30890,N_29228,N_29086);
or U30891 (N_30891,N_29386,N_29200);
xor U30892 (N_30892,N_29293,N_29605);
nor U30893 (N_30893,N_29509,N_29795);
nor U30894 (N_30894,N_29705,N_29873);
and U30895 (N_30895,N_29527,N_29721);
or U30896 (N_30896,N_29850,N_29938);
xor U30897 (N_30897,N_29793,N_29370);
nor U30898 (N_30898,N_29819,N_29838);
or U30899 (N_30899,N_29385,N_29596);
and U30900 (N_30900,N_29796,N_29280);
and U30901 (N_30901,N_29618,N_29019);
or U30902 (N_30902,N_29316,N_29256);
and U30903 (N_30903,N_29635,N_29053);
and U30904 (N_30904,N_29834,N_29609);
and U30905 (N_30905,N_29343,N_29100);
or U30906 (N_30906,N_29920,N_29580);
and U30907 (N_30907,N_29286,N_29363);
or U30908 (N_30908,N_29741,N_29034);
or U30909 (N_30909,N_29910,N_29060);
and U30910 (N_30910,N_29483,N_29023);
nand U30911 (N_30911,N_29342,N_29219);
and U30912 (N_30912,N_29993,N_29126);
nand U30913 (N_30913,N_29291,N_29391);
nor U30914 (N_30914,N_29029,N_29273);
nor U30915 (N_30915,N_29285,N_29411);
nor U30916 (N_30916,N_29389,N_29523);
and U30917 (N_30917,N_29941,N_29838);
xnor U30918 (N_30918,N_29400,N_29224);
nor U30919 (N_30919,N_29461,N_29610);
nor U30920 (N_30920,N_29169,N_29296);
nor U30921 (N_30921,N_29683,N_29441);
nor U30922 (N_30922,N_29665,N_29070);
and U30923 (N_30923,N_29904,N_29676);
nor U30924 (N_30924,N_29875,N_29336);
nand U30925 (N_30925,N_29006,N_29953);
nand U30926 (N_30926,N_29204,N_29772);
nor U30927 (N_30927,N_29030,N_29991);
or U30928 (N_30928,N_29221,N_29415);
xnor U30929 (N_30929,N_29000,N_29480);
nand U30930 (N_30930,N_29393,N_29360);
and U30931 (N_30931,N_29376,N_29454);
or U30932 (N_30932,N_29723,N_29262);
and U30933 (N_30933,N_29761,N_29099);
and U30934 (N_30934,N_29621,N_29172);
nand U30935 (N_30935,N_29522,N_29872);
or U30936 (N_30936,N_29999,N_29980);
xnor U30937 (N_30937,N_29165,N_29921);
nor U30938 (N_30938,N_29050,N_29194);
nor U30939 (N_30939,N_29604,N_29219);
nor U30940 (N_30940,N_29863,N_29484);
and U30941 (N_30941,N_29910,N_29111);
or U30942 (N_30942,N_29983,N_29902);
xor U30943 (N_30943,N_29540,N_29327);
xnor U30944 (N_30944,N_29276,N_29268);
and U30945 (N_30945,N_29295,N_29720);
nand U30946 (N_30946,N_29537,N_29383);
or U30947 (N_30947,N_29222,N_29727);
nand U30948 (N_30948,N_29458,N_29468);
xnor U30949 (N_30949,N_29951,N_29241);
nand U30950 (N_30950,N_29593,N_29936);
or U30951 (N_30951,N_29431,N_29307);
xnor U30952 (N_30952,N_29964,N_29882);
xor U30953 (N_30953,N_29606,N_29011);
nor U30954 (N_30954,N_29338,N_29429);
or U30955 (N_30955,N_29326,N_29412);
nor U30956 (N_30956,N_29648,N_29100);
or U30957 (N_30957,N_29870,N_29168);
nor U30958 (N_30958,N_29492,N_29983);
or U30959 (N_30959,N_29353,N_29825);
xor U30960 (N_30960,N_29262,N_29695);
nor U30961 (N_30961,N_29399,N_29940);
nand U30962 (N_30962,N_29050,N_29886);
nand U30963 (N_30963,N_29732,N_29115);
nand U30964 (N_30964,N_29327,N_29850);
nand U30965 (N_30965,N_29121,N_29572);
and U30966 (N_30966,N_29460,N_29043);
nor U30967 (N_30967,N_29287,N_29426);
nor U30968 (N_30968,N_29722,N_29697);
nand U30969 (N_30969,N_29039,N_29299);
or U30970 (N_30970,N_29972,N_29827);
nand U30971 (N_30971,N_29829,N_29489);
or U30972 (N_30972,N_29916,N_29612);
and U30973 (N_30973,N_29351,N_29300);
nand U30974 (N_30974,N_29738,N_29948);
xnor U30975 (N_30975,N_29345,N_29904);
and U30976 (N_30976,N_29770,N_29165);
and U30977 (N_30977,N_29509,N_29719);
nor U30978 (N_30978,N_29890,N_29960);
nor U30979 (N_30979,N_29818,N_29588);
nand U30980 (N_30980,N_29774,N_29118);
nand U30981 (N_30981,N_29979,N_29755);
xor U30982 (N_30982,N_29880,N_29221);
xor U30983 (N_30983,N_29847,N_29322);
nand U30984 (N_30984,N_29946,N_29770);
nand U30985 (N_30985,N_29367,N_29491);
xnor U30986 (N_30986,N_29993,N_29695);
nor U30987 (N_30987,N_29385,N_29451);
xnor U30988 (N_30988,N_29736,N_29505);
or U30989 (N_30989,N_29066,N_29832);
nor U30990 (N_30990,N_29687,N_29164);
nand U30991 (N_30991,N_29987,N_29337);
nand U30992 (N_30992,N_29467,N_29739);
and U30993 (N_30993,N_29962,N_29295);
nor U30994 (N_30994,N_29096,N_29412);
or U30995 (N_30995,N_29152,N_29630);
nor U30996 (N_30996,N_29741,N_29210);
nand U30997 (N_30997,N_29187,N_29099);
or U30998 (N_30998,N_29647,N_29383);
and U30999 (N_30999,N_29209,N_29452);
and U31000 (N_31000,N_30440,N_30523);
nand U31001 (N_31001,N_30683,N_30166);
nand U31002 (N_31002,N_30762,N_30056);
nand U31003 (N_31003,N_30303,N_30107);
or U31004 (N_31004,N_30252,N_30322);
nand U31005 (N_31005,N_30837,N_30239);
xor U31006 (N_31006,N_30779,N_30456);
and U31007 (N_31007,N_30896,N_30789);
and U31008 (N_31008,N_30085,N_30805);
and U31009 (N_31009,N_30241,N_30876);
or U31010 (N_31010,N_30644,N_30582);
nor U31011 (N_31011,N_30945,N_30980);
and U31012 (N_31012,N_30257,N_30767);
and U31013 (N_31013,N_30591,N_30246);
and U31014 (N_31014,N_30677,N_30502);
and U31015 (N_31015,N_30367,N_30357);
nand U31016 (N_31016,N_30231,N_30399);
nand U31017 (N_31017,N_30288,N_30610);
and U31018 (N_31018,N_30658,N_30974);
and U31019 (N_31019,N_30254,N_30422);
xor U31020 (N_31020,N_30300,N_30569);
nor U31021 (N_31021,N_30574,N_30401);
and U31022 (N_31022,N_30988,N_30943);
or U31023 (N_31023,N_30018,N_30940);
or U31024 (N_31024,N_30327,N_30337);
and U31025 (N_31025,N_30784,N_30102);
nor U31026 (N_31026,N_30335,N_30522);
and U31027 (N_31027,N_30823,N_30245);
xor U31028 (N_31028,N_30792,N_30728);
nand U31029 (N_31029,N_30135,N_30383);
and U31030 (N_31030,N_30167,N_30978);
or U31031 (N_31031,N_30060,N_30958);
and U31032 (N_31032,N_30841,N_30140);
xnor U31033 (N_31033,N_30911,N_30725);
or U31034 (N_31034,N_30509,N_30982);
nand U31035 (N_31035,N_30206,N_30799);
xnor U31036 (N_31036,N_30520,N_30479);
nor U31037 (N_31037,N_30312,N_30680);
xnor U31038 (N_31038,N_30602,N_30636);
nand U31039 (N_31039,N_30626,N_30439);
xnor U31040 (N_31040,N_30096,N_30143);
xor U31041 (N_31041,N_30656,N_30998);
nand U31042 (N_31042,N_30123,N_30459);
nand U31043 (N_31043,N_30153,N_30547);
xor U31044 (N_31044,N_30764,N_30358);
or U31045 (N_31045,N_30209,N_30187);
xnor U31046 (N_31046,N_30718,N_30601);
nor U31047 (N_31047,N_30179,N_30645);
and U31048 (N_31048,N_30593,N_30804);
and U31049 (N_31049,N_30320,N_30647);
or U31050 (N_31050,N_30203,N_30304);
and U31051 (N_31051,N_30605,N_30164);
xor U31052 (N_31052,N_30470,N_30724);
nor U31053 (N_31053,N_30268,N_30546);
xnor U31054 (N_31054,N_30460,N_30863);
and U31055 (N_31055,N_30033,N_30753);
nand U31056 (N_31056,N_30256,N_30771);
nand U31057 (N_31057,N_30833,N_30247);
and U31058 (N_31058,N_30759,N_30008);
nor U31059 (N_31059,N_30934,N_30519);
nor U31060 (N_31060,N_30735,N_30169);
and U31061 (N_31061,N_30156,N_30510);
xnor U31062 (N_31062,N_30035,N_30009);
or U31063 (N_31063,N_30219,N_30892);
xnor U31064 (N_31064,N_30275,N_30390);
xor U31065 (N_31065,N_30448,N_30310);
xnor U31066 (N_31066,N_30617,N_30961);
xor U31067 (N_31067,N_30816,N_30525);
nor U31068 (N_31068,N_30483,N_30027);
nor U31069 (N_31069,N_30270,N_30369);
nand U31070 (N_31070,N_30919,N_30318);
or U31071 (N_31071,N_30738,N_30671);
and U31072 (N_31072,N_30936,N_30603);
or U31073 (N_31073,N_30824,N_30580);
or U31074 (N_31074,N_30098,N_30737);
or U31075 (N_31075,N_30877,N_30365);
and U31076 (N_31076,N_30248,N_30400);
nand U31077 (N_31077,N_30886,N_30114);
nor U31078 (N_31078,N_30971,N_30229);
nand U31079 (N_31079,N_30014,N_30561);
xor U31080 (N_31080,N_30531,N_30711);
or U31081 (N_31081,N_30797,N_30528);
nor U31082 (N_31082,N_30878,N_30050);
xnor U31083 (N_31083,N_30585,N_30362);
nand U31084 (N_31084,N_30484,N_30859);
nand U31085 (N_31085,N_30161,N_30492);
xor U31086 (N_31086,N_30409,N_30534);
xnor U31087 (N_31087,N_30118,N_30223);
nand U31088 (N_31088,N_30986,N_30893);
and U31089 (N_31089,N_30101,N_30111);
nor U31090 (N_31090,N_30627,N_30091);
nor U31091 (N_31091,N_30088,N_30914);
nor U31092 (N_31092,N_30827,N_30127);
nand U31093 (N_31093,N_30653,N_30652);
xor U31094 (N_31094,N_30935,N_30095);
nor U31095 (N_31095,N_30145,N_30214);
or U31096 (N_31096,N_30800,N_30541);
and U31097 (N_31097,N_30146,N_30190);
nor U31098 (N_31098,N_30630,N_30477);
xnor U31099 (N_31099,N_30366,N_30493);
and U31100 (N_31100,N_30432,N_30716);
xor U31101 (N_31101,N_30259,N_30427);
and U31102 (N_31102,N_30845,N_30193);
xor U31103 (N_31103,N_30103,N_30951);
nand U31104 (N_31104,N_30150,N_30504);
and U31105 (N_31105,N_30371,N_30685);
and U31106 (N_31106,N_30973,N_30556);
nor U31107 (N_31107,N_30545,N_30213);
xor U31108 (N_31108,N_30537,N_30070);
or U31109 (N_31109,N_30813,N_30202);
nand U31110 (N_31110,N_30115,N_30794);
nor U31111 (N_31111,N_30138,N_30864);
and U31112 (N_31112,N_30195,N_30281);
or U31113 (N_31113,N_30368,N_30861);
nor U31114 (N_31114,N_30862,N_30632);
nand U31115 (N_31115,N_30544,N_30681);
or U31116 (N_31116,N_30831,N_30210);
xnor U31117 (N_31117,N_30567,N_30807);
nor U31118 (N_31118,N_30575,N_30468);
xor U31119 (N_31119,N_30727,N_30324);
or U31120 (N_31120,N_30490,N_30404);
and U31121 (N_31121,N_30676,N_30385);
or U31122 (N_31122,N_30419,N_30461);
nand U31123 (N_31123,N_30899,N_30836);
and U31124 (N_31124,N_30551,N_30624);
and U31125 (N_31125,N_30990,N_30392);
nor U31126 (N_31126,N_30158,N_30446);
or U31127 (N_31127,N_30377,N_30352);
nor U31128 (N_31128,N_30301,N_30177);
nand U31129 (N_31129,N_30080,N_30218);
nand U31130 (N_31130,N_30879,N_30772);
nand U31131 (N_31131,N_30809,N_30758);
xor U31132 (N_31132,N_30444,N_30710);
xor U31133 (N_31133,N_30696,N_30273);
or U31134 (N_31134,N_30686,N_30276);
nand U31135 (N_31135,N_30277,N_30678);
nor U31136 (N_31136,N_30489,N_30554);
or U31137 (N_31137,N_30756,N_30396);
xor U31138 (N_31138,N_30408,N_30898);
nand U31139 (N_31139,N_30242,N_30511);
or U31140 (N_31140,N_30433,N_30840);
or U31141 (N_31141,N_30105,N_30126);
nor U31142 (N_31142,N_30702,N_30949);
and U31143 (N_31143,N_30704,N_30306);
and U31144 (N_31144,N_30506,N_30733);
or U31145 (N_31145,N_30010,N_30669);
nand U31146 (N_31146,N_30852,N_30835);
and U31147 (N_31147,N_30969,N_30082);
or U31148 (N_31148,N_30550,N_30089);
or U31149 (N_31149,N_30142,N_30494);
nor U31150 (N_31150,N_30130,N_30113);
xor U31151 (N_31151,N_30598,N_30995);
and U31152 (N_31152,N_30395,N_30053);
or U31153 (N_31153,N_30761,N_30321);
nand U31154 (N_31154,N_30013,N_30372);
and U31155 (N_31155,N_30250,N_30673);
nor U31156 (N_31156,N_30355,N_30810);
or U31157 (N_31157,N_30781,N_30224);
nand U31158 (N_31158,N_30110,N_30768);
nand U31159 (N_31159,N_30315,N_30564);
and U31160 (N_31160,N_30578,N_30415);
nor U31161 (N_31161,N_30867,N_30019);
or U31162 (N_31162,N_30116,N_30482);
and U31163 (N_31163,N_30613,N_30665);
and U31164 (N_31164,N_30348,N_30611);
nor U31165 (N_31165,N_30924,N_30264);
or U31166 (N_31166,N_30894,N_30297);
and U31167 (N_31167,N_30104,N_30720);
or U31168 (N_31168,N_30350,N_30151);
xor U31169 (N_31169,N_30087,N_30866);
and U31170 (N_31170,N_30317,N_30684);
xor U31171 (N_31171,N_30072,N_30251);
nand U31172 (N_31172,N_30455,N_30125);
or U31173 (N_31173,N_30488,N_30289);
nor U31174 (N_31174,N_30044,N_30594);
or U31175 (N_31175,N_30891,N_30438);
xor U31176 (N_31176,N_30382,N_30705);
nand U31177 (N_31177,N_30638,N_30485);
nand U31178 (N_31178,N_30787,N_30829);
nor U31179 (N_31179,N_30948,N_30347);
xor U31180 (N_31180,N_30486,N_30856);
nand U31181 (N_31181,N_30571,N_30992);
xnor U31182 (N_31182,N_30426,N_30664);
and U31183 (N_31183,N_30715,N_30425);
and U31184 (N_31184,N_30985,N_30222);
and U31185 (N_31185,N_30930,N_30933);
nor U31186 (N_31186,N_30041,N_30015);
or U31187 (N_31187,N_30962,N_30849);
and U31188 (N_31188,N_30148,N_30240);
or U31189 (N_31189,N_30843,N_30283);
nor U31190 (N_31190,N_30436,N_30929);
or U31191 (N_31191,N_30428,N_30631);
and U31192 (N_31192,N_30063,N_30064);
xor U31193 (N_31193,N_30901,N_30539);
nor U31194 (N_31194,N_30858,N_30212);
and U31195 (N_31195,N_30650,N_30712);
xnor U31196 (N_31196,N_30073,N_30555);
and U31197 (N_31197,N_30803,N_30540);
nor U31198 (N_31198,N_30783,N_30029);
or U31199 (N_31199,N_30905,N_30048);
or U31200 (N_31200,N_30947,N_30183);
or U31201 (N_31201,N_30773,N_30120);
and U31202 (N_31202,N_30134,N_30532);
nand U31203 (N_31203,N_30196,N_30174);
xnor U31204 (N_31204,N_30162,N_30917);
and U31205 (N_31205,N_30131,N_30584);
nor U31206 (N_31206,N_30868,N_30625);
and U31207 (N_31207,N_30937,N_30228);
nand U31208 (N_31208,N_30999,N_30388);
and U31209 (N_31209,N_30966,N_30291);
nor U31210 (N_31210,N_30959,N_30765);
xnor U31211 (N_31211,N_30463,N_30791);
nor U31212 (N_31212,N_30552,N_30386);
nor U31213 (N_31213,N_30307,N_30269);
xnor U31214 (N_31214,N_30021,N_30648);
or U31215 (N_31215,N_30394,N_30354);
nor U31216 (N_31216,N_30994,N_30046);
nor U31217 (N_31217,N_30749,N_30192);
nor U31218 (N_31218,N_30478,N_30236);
nor U31219 (N_31219,N_30530,N_30067);
xor U31220 (N_31220,N_30227,N_30298);
nand U31221 (N_31221,N_30071,N_30047);
nand U31222 (N_31222,N_30215,N_30380);
nand U31223 (N_31223,N_30039,N_30576);
and U31224 (N_31224,N_30226,N_30154);
nor U31225 (N_31225,N_30562,N_30639);
nand U31226 (N_31226,N_30526,N_30378);
nor U31227 (N_31227,N_30560,N_30643);
xor U31228 (N_31228,N_30972,N_30147);
or U31229 (N_31229,N_30946,N_30186);
xnor U31230 (N_31230,N_30991,N_30069);
xnor U31231 (N_31231,N_30821,N_30445);
nor U31232 (N_31232,N_30882,N_30722);
nor U31233 (N_31233,N_30234,N_30370);
nand U31234 (N_31234,N_30729,N_30667);
xor U31235 (N_31235,N_30697,N_30828);
nor U31236 (N_31236,N_30129,N_30418);
xor U31237 (N_31237,N_30331,N_30583);
and U31238 (N_31238,N_30491,N_30723);
or U31239 (N_31239,N_30932,N_30458);
and U31240 (N_31240,N_30052,N_30373);
nor U31241 (N_31241,N_30323,N_30391);
nand U31242 (N_31242,N_30182,N_30201);
nor U31243 (N_31243,N_30589,N_30927);
and U31244 (N_31244,N_30338,N_30498);
nor U31245 (N_31245,N_30597,N_30587);
nand U31246 (N_31246,N_30022,N_30709);
nand U31247 (N_31247,N_30614,N_30920);
xor U31248 (N_31248,N_30881,N_30319);
or U31249 (N_31249,N_30847,N_30062);
and U31250 (N_31250,N_30001,N_30913);
or U31251 (N_31251,N_30983,N_30640);
xnor U31252 (N_31252,N_30000,N_30457);
xnor U31253 (N_31253,N_30031,N_30449);
nor U31254 (N_31254,N_30529,N_30916);
nand U31255 (N_31255,N_30160,N_30925);
nand U31256 (N_31256,N_30065,N_30078);
nand U31257 (N_31257,N_30199,N_30180);
and U31258 (N_31258,N_30476,N_30634);
or U31259 (N_31259,N_30176,N_30608);
nand U31260 (N_31260,N_30698,N_30284);
nor U31261 (N_31261,N_30443,N_30020);
nor U31262 (N_31262,N_30453,N_30083);
nor U31263 (N_31263,N_30612,N_30204);
nand U31264 (N_31264,N_30410,N_30462);
nor U31265 (N_31265,N_30207,N_30641);
or U31266 (N_31266,N_30513,N_30258);
xnor U31267 (N_31267,N_30588,N_30785);
nor U31268 (N_31268,N_30379,N_30984);
xnor U31269 (N_31269,N_30353,N_30345);
or U31270 (N_31270,N_30777,N_30235);
or U31271 (N_31271,N_30880,N_30155);
nand U31272 (N_31272,N_30407,N_30790);
xor U31273 (N_31273,N_30061,N_30726);
and U31274 (N_31274,N_30708,N_30049);
xnor U31275 (N_31275,N_30171,N_30865);
xor U31276 (N_31276,N_30117,N_30743);
xnor U31277 (N_31277,N_30747,N_30189);
or U31278 (N_31278,N_30466,N_30744);
xnor U31279 (N_31279,N_30007,N_30757);
nand U31280 (N_31280,N_30136,N_30993);
nand U31281 (N_31281,N_30542,N_30329);
and U31282 (N_31282,N_30233,N_30055);
nor U31283 (N_31283,N_30121,N_30441);
nor U31284 (N_31284,N_30848,N_30548);
nor U31285 (N_31285,N_30360,N_30745);
nand U31286 (N_31286,N_30817,N_30170);
nand U31287 (N_31287,N_30870,N_30682);
nor U31288 (N_31288,N_30157,N_30280);
nor U31289 (N_31289,N_30507,N_30294);
or U31290 (N_31290,N_30912,N_30850);
or U31291 (N_31291,N_30695,N_30017);
or U31292 (N_31292,N_30883,N_30406);
or U31293 (N_31293,N_30006,N_30282);
xnor U31294 (N_31294,N_30620,N_30420);
xnor U31295 (N_31295,N_30622,N_30076);
or U31296 (N_31296,N_30475,N_30344);
and U31297 (N_31297,N_30243,N_30346);
nand U31298 (N_31298,N_30826,N_30742);
or U31299 (N_31299,N_30713,N_30944);
nor U31300 (N_31300,N_30030,N_30132);
and U31301 (N_31301,N_30606,N_30795);
xnor U31302 (N_31302,N_30706,N_30802);
nand U31303 (N_31303,N_30793,N_30314);
or U31304 (N_31304,N_30516,N_30987);
or U31305 (N_31305,N_30108,N_30465);
or U31306 (N_31306,N_30398,N_30558);
nand U31307 (N_31307,N_30707,N_30825);
nor U31308 (N_31308,N_30568,N_30043);
xnor U31309 (N_31309,N_30628,N_30265);
nand U31310 (N_31310,N_30232,N_30262);
nand U31311 (N_31311,N_30471,N_30042);
nor U31312 (N_31312,N_30796,N_30496);
xnor U31313 (N_31313,N_30435,N_30660);
and U31314 (N_31314,N_30953,N_30128);
or U31315 (N_31315,N_30618,N_30662);
nand U31316 (N_31316,N_30834,N_30389);
or U31317 (N_31317,N_30846,N_30600);
nor U31318 (N_31318,N_30616,N_30092);
nand U31319 (N_31319,N_30910,N_30375);
nand U31320 (N_31320,N_30191,N_30577);
and U31321 (N_31321,N_30026,N_30703);
xor U31322 (N_31322,N_30693,N_30290);
nor U31323 (N_31323,N_30874,N_30093);
and U31324 (N_31324,N_30424,N_30887);
xor U31325 (N_31325,N_30997,N_30557);
nand U31326 (N_31326,N_30194,N_30975);
or U31327 (N_31327,N_30249,N_30688);
nand U31328 (N_31328,N_30687,N_30633);
xnor U31329 (N_31329,N_30099,N_30906);
and U31330 (N_31330,N_30518,N_30374);
xnor U31331 (N_31331,N_30672,N_30607);
nand U31332 (N_31332,N_30302,N_30165);
nand U31333 (N_31333,N_30152,N_30253);
xor U31334 (N_31334,N_30524,N_30292);
and U31335 (N_31335,N_30909,N_30731);
or U31336 (N_31336,N_30037,N_30381);
nor U31337 (N_31337,N_30330,N_30918);
or U31338 (N_31338,N_30168,N_30596);
nor U31339 (N_31339,N_30989,N_30950);
and U31340 (N_31340,N_30261,N_30885);
or U31341 (N_31341,N_30734,N_30003);
xnor U31342 (N_31342,N_30328,N_30811);
or U31343 (N_31343,N_30889,N_30512);
nand U31344 (N_31344,N_30563,N_30413);
and U31345 (N_31345,N_30349,N_30717);
and U31346 (N_31346,N_30780,N_30818);
nor U31347 (N_31347,N_30079,N_30939);
or U31348 (N_31348,N_30635,N_30938);
or U31349 (N_31349,N_30351,N_30172);
nor U31350 (N_31350,N_30205,N_30527);
and U31351 (N_31351,N_30336,N_30699);
xnor U31352 (N_31352,N_30333,N_30670);
nor U31353 (N_31353,N_30860,N_30957);
or U31354 (N_31354,N_30244,N_30119);
nand U31355 (N_31355,N_30573,N_30842);
and U31356 (N_31356,N_30739,N_30272);
or U31357 (N_31357,N_30267,N_30163);
nor U31358 (N_31358,N_30801,N_30430);
xnor U31359 (N_31359,N_30295,N_30472);
or U31360 (N_31360,N_30313,N_30719);
nor U31361 (N_31361,N_30904,N_30536);
and U31362 (N_31362,N_30769,N_30996);
nor U31363 (N_31363,N_30815,N_30871);
nor U31364 (N_31364,N_30450,N_30387);
nand U31365 (N_31365,N_30402,N_30500);
nor U31366 (N_31366,N_30403,N_30051);
and U31367 (N_31367,N_30657,N_30299);
or U31368 (N_31368,N_30122,N_30356);
nand U31369 (N_31369,N_30872,N_30004);
xor U31370 (N_31370,N_30890,N_30808);
xnor U31371 (N_31371,N_30970,N_30642);
xor U31372 (N_31372,N_30309,N_30260);
xnor U31373 (N_31373,N_30188,N_30084);
nor U31374 (N_31374,N_30361,N_30581);
nand U31375 (N_31375,N_30454,N_30287);
or U31376 (N_31376,N_30760,N_30873);
nor U31377 (N_31377,N_30895,N_30661);
xnor U31378 (N_31378,N_30763,N_30505);
nand U31379 (N_31379,N_30363,N_30820);
and U31380 (N_31380,N_30431,N_30057);
xor U31381 (N_31381,N_30595,N_30200);
nor U31382 (N_31382,N_30417,N_30032);
or U31383 (N_31383,N_30181,N_30884);
nand U31384 (N_31384,N_30217,N_30746);
xor U31385 (N_31385,N_30045,N_30888);
nor U31386 (N_31386,N_30654,N_30497);
nand U31387 (N_31387,N_30124,N_30159);
nand U31388 (N_31388,N_30334,N_30853);
xor U31389 (N_31389,N_30691,N_30646);
nand U31390 (N_31390,N_30806,N_30832);
xor U31391 (N_31391,N_30754,N_30133);
or U31392 (N_31392,N_30736,N_30752);
and U31393 (N_31393,N_30308,N_30649);
nand U31394 (N_31394,N_30305,N_30036);
nand U31395 (N_31395,N_30086,N_30968);
and U31396 (N_31396,N_30926,N_30238);
xnor U31397 (N_31397,N_30106,N_30679);
nor U31398 (N_31398,N_30579,N_30819);
or U31399 (N_31399,N_30464,N_30501);
or U31400 (N_31400,N_30663,N_30514);
nand U31401 (N_31401,N_30732,N_30225);
xor U31402 (N_31402,N_30416,N_30921);
or U31403 (N_31403,N_30776,N_30012);
nand U31404 (N_31404,N_30941,N_30255);
nand U31405 (N_31405,N_30112,N_30090);
or U31406 (N_31406,N_30293,N_30963);
or U31407 (N_31407,N_30565,N_30059);
nand U31408 (N_31408,N_30751,N_30414);
or U31409 (N_31409,N_30359,N_30766);
nand U31410 (N_31410,N_30689,N_30508);
or U31411 (N_31411,N_30740,N_30499);
or U31412 (N_31412,N_30339,N_30830);
nor U31413 (N_31413,N_30094,N_30467);
or U31414 (N_31414,N_30674,N_30474);
xnor U31415 (N_31415,N_30332,N_30198);
xor U31416 (N_31416,N_30981,N_30572);
nand U31417 (N_31417,N_30692,N_30405);
or U31418 (N_31418,N_30619,N_30411);
or U31419 (N_31419,N_30495,N_30964);
or U31420 (N_31420,N_30447,N_30659);
nand U31421 (N_31421,N_30184,N_30237);
and U31422 (N_31422,N_30016,N_30025);
nor U31423 (N_31423,N_30109,N_30034);
xnor U31424 (N_31424,N_30434,N_30137);
xor U31425 (N_31425,N_30178,N_30005);
xnor U31426 (N_31426,N_30521,N_30325);
xor U31427 (N_31427,N_30623,N_30755);
and U31428 (N_31428,N_30002,N_30469);
and U31429 (N_31429,N_30637,N_30741);
xor U31430 (N_31430,N_30721,N_30028);
nand U31431 (N_31431,N_30977,N_30139);
nand U31432 (N_31432,N_30965,N_30480);
or U31433 (N_31433,N_30778,N_30221);
nand U31434 (N_31434,N_30144,N_30376);
nand U31435 (N_31435,N_30857,N_30604);
nand U31436 (N_31436,N_30175,N_30839);
or U31437 (N_31437,N_30296,N_30694);
nand U31438 (N_31438,N_30915,N_30979);
xnor U31439 (N_31439,N_30266,N_30040);
or U31440 (N_31440,N_30285,N_30535);
nand U31441 (N_31441,N_30928,N_30629);
nor U31442 (N_31442,N_30149,N_30216);
nor U31443 (N_31443,N_30533,N_30286);
nor U31444 (N_31444,N_30515,N_30609);
and U31445 (N_31445,N_30077,N_30271);
nand U31446 (N_31446,N_30931,N_30024);
nand U31447 (N_31447,N_30701,N_30263);
nand U31448 (N_31448,N_30897,N_30316);
nand U31449 (N_31449,N_30675,N_30437);
and U31450 (N_31450,N_30423,N_30621);
nor U31451 (N_31451,N_30473,N_30342);
and U31452 (N_31452,N_30855,N_30812);
nor U31453 (N_31453,N_30774,N_30908);
or U31454 (N_31454,N_30566,N_30503);
xnor U31455 (N_31455,N_30690,N_30788);
nor U31456 (N_31456,N_30786,N_30900);
nand U31457 (N_31457,N_30869,N_30770);
xnor U31458 (N_31458,N_30851,N_30775);
or U31459 (N_31459,N_30730,N_30902);
xor U31460 (N_31460,N_30100,N_30066);
and U31461 (N_31461,N_30844,N_30421);
nand U31462 (N_31462,N_30054,N_30451);
and U31463 (N_31463,N_30279,N_30955);
xnor U31464 (N_31464,N_30553,N_30549);
nor U31465 (N_31465,N_30750,N_30274);
or U31466 (N_31466,N_30487,N_30666);
and U31467 (N_31467,N_30097,N_30942);
nand U31468 (N_31468,N_30854,N_30038);
nor U31469 (N_31469,N_30278,N_30173);
xor U31470 (N_31470,N_30798,N_30141);
xor U31471 (N_31471,N_30954,N_30875);
xor U31472 (N_31472,N_30592,N_30429);
xor U31473 (N_31473,N_30923,N_30960);
xor U31474 (N_31474,N_30058,N_30903);
nor U31475 (N_31475,N_30075,N_30822);
nor U31476 (N_31476,N_30341,N_30068);
or U31477 (N_31477,N_30700,N_30586);
and U31478 (N_31478,N_30023,N_30081);
nand U31479 (N_31479,N_30074,N_30838);
or U31480 (N_31480,N_30326,N_30590);
xnor U31481 (N_31481,N_30907,N_30517);
and U31482 (N_31482,N_30340,N_30384);
nor U31483 (N_31483,N_30668,N_30922);
xor U31484 (N_31484,N_30651,N_30599);
and U31485 (N_31485,N_30543,N_30814);
and U31486 (N_31486,N_30343,N_30976);
nand U31487 (N_31487,N_30397,N_30364);
and U31488 (N_31488,N_30538,N_30442);
nor U31489 (N_31489,N_30655,N_30452);
nand U31490 (N_31490,N_30211,N_30952);
xnor U31491 (N_31491,N_30748,N_30197);
and U31492 (N_31492,N_30393,N_30956);
and U31493 (N_31493,N_30185,N_30559);
or U31494 (N_31494,N_30481,N_30230);
or U31495 (N_31495,N_30208,N_30220);
or U31496 (N_31496,N_30782,N_30967);
xor U31497 (N_31497,N_30615,N_30311);
nand U31498 (N_31498,N_30570,N_30714);
nand U31499 (N_31499,N_30011,N_30412);
nand U31500 (N_31500,N_30980,N_30507);
xor U31501 (N_31501,N_30321,N_30736);
and U31502 (N_31502,N_30085,N_30272);
and U31503 (N_31503,N_30264,N_30774);
and U31504 (N_31504,N_30598,N_30753);
and U31505 (N_31505,N_30946,N_30144);
and U31506 (N_31506,N_30380,N_30242);
or U31507 (N_31507,N_30019,N_30902);
nor U31508 (N_31508,N_30190,N_30661);
nand U31509 (N_31509,N_30989,N_30273);
and U31510 (N_31510,N_30746,N_30390);
xnor U31511 (N_31511,N_30828,N_30243);
and U31512 (N_31512,N_30121,N_30893);
nor U31513 (N_31513,N_30167,N_30747);
and U31514 (N_31514,N_30807,N_30801);
xor U31515 (N_31515,N_30740,N_30779);
or U31516 (N_31516,N_30410,N_30799);
xor U31517 (N_31517,N_30208,N_30792);
or U31518 (N_31518,N_30674,N_30654);
xor U31519 (N_31519,N_30906,N_30439);
or U31520 (N_31520,N_30923,N_30587);
nand U31521 (N_31521,N_30066,N_30039);
and U31522 (N_31522,N_30307,N_30633);
nand U31523 (N_31523,N_30002,N_30907);
nand U31524 (N_31524,N_30021,N_30328);
and U31525 (N_31525,N_30304,N_30385);
and U31526 (N_31526,N_30849,N_30635);
xnor U31527 (N_31527,N_30922,N_30795);
or U31528 (N_31528,N_30978,N_30553);
nor U31529 (N_31529,N_30553,N_30213);
nand U31530 (N_31530,N_30129,N_30913);
nor U31531 (N_31531,N_30987,N_30346);
xnor U31532 (N_31532,N_30584,N_30286);
nor U31533 (N_31533,N_30774,N_30789);
nor U31534 (N_31534,N_30719,N_30070);
or U31535 (N_31535,N_30707,N_30276);
xnor U31536 (N_31536,N_30804,N_30589);
or U31537 (N_31537,N_30201,N_30532);
nor U31538 (N_31538,N_30725,N_30225);
and U31539 (N_31539,N_30958,N_30986);
or U31540 (N_31540,N_30654,N_30026);
xor U31541 (N_31541,N_30768,N_30547);
or U31542 (N_31542,N_30597,N_30367);
nand U31543 (N_31543,N_30351,N_30905);
or U31544 (N_31544,N_30258,N_30704);
xnor U31545 (N_31545,N_30941,N_30741);
nand U31546 (N_31546,N_30264,N_30008);
nor U31547 (N_31547,N_30745,N_30577);
nand U31548 (N_31548,N_30291,N_30246);
nor U31549 (N_31549,N_30678,N_30970);
or U31550 (N_31550,N_30306,N_30429);
nand U31551 (N_31551,N_30621,N_30561);
nand U31552 (N_31552,N_30919,N_30422);
and U31553 (N_31553,N_30665,N_30864);
nand U31554 (N_31554,N_30367,N_30829);
and U31555 (N_31555,N_30042,N_30079);
and U31556 (N_31556,N_30856,N_30489);
xor U31557 (N_31557,N_30652,N_30044);
and U31558 (N_31558,N_30264,N_30030);
and U31559 (N_31559,N_30703,N_30323);
or U31560 (N_31560,N_30033,N_30330);
and U31561 (N_31561,N_30593,N_30518);
xor U31562 (N_31562,N_30329,N_30142);
nand U31563 (N_31563,N_30002,N_30607);
nand U31564 (N_31564,N_30569,N_30370);
nand U31565 (N_31565,N_30901,N_30009);
nand U31566 (N_31566,N_30287,N_30198);
or U31567 (N_31567,N_30188,N_30584);
nor U31568 (N_31568,N_30115,N_30245);
nand U31569 (N_31569,N_30697,N_30701);
or U31570 (N_31570,N_30898,N_30956);
nor U31571 (N_31571,N_30569,N_30782);
and U31572 (N_31572,N_30109,N_30651);
nor U31573 (N_31573,N_30274,N_30962);
nor U31574 (N_31574,N_30949,N_30059);
xor U31575 (N_31575,N_30966,N_30550);
xor U31576 (N_31576,N_30172,N_30032);
xor U31577 (N_31577,N_30175,N_30164);
nand U31578 (N_31578,N_30310,N_30954);
xor U31579 (N_31579,N_30552,N_30641);
xor U31580 (N_31580,N_30293,N_30678);
xor U31581 (N_31581,N_30462,N_30445);
and U31582 (N_31582,N_30028,N_30021);
nor U31583 (N_31583,N_30698,N_30720);
and U31584 (N_31584,N_30425,N_30507);
and U31585 (N_31585,N_30550,N_30944);
or U31586 (N_31586,N_30728,N_30558);
or U31587 (N_31587,N_30148,N_30052);
nand U31588 (N_31588,N_30663,N_30533);
nand U31589 (N_31589,N_30734,N_30531);
xor U31590 (N_31590,N_30116,N_30496);
xnor U31591 (N_31591,N_30319,N_30426);
nor U31592 (N_31592,N_30332,N_30408);
xnor U31593 (N_31593,N_30065,N_30540);
and U31594 (N_31594,N_30072,N_30215);
nor U31595 (N_31595,N_30934,N_30888);
or U31596 (N_31596,N_30657,N_30222);
and U31597 (N_31597,N_30904,N_30887);
and U31598 (N_31598,N_30245,N_30424);
xnor U31599 (N_31599,N_30543,N_30681);
nand U31600 (N_31600,N_30836,N_30012);
nor U31601 (N_31601,N_30650,N_30795);
or U31602 (N_31602,N_30667,N_30316);
xor U31603 (N_31603,N_30970,N_30715);
nor U31604 (N_31604,N_30693,N_30582);
or U31605 (N_31605,N_30373,N_30613);
or U31606 (N_31606,N_30830,N_30677);
nand U31607 (N_31607,N_30639,N_30775);
nand U31608 (N_31608,N_30329,N_30786);
xor U31609 (N_31609,N_30095,N_30658);
nand U31610 (N_31610,N_30412,N_30410);
and U31611 (N_31611,N_30340,N_30747);
xnor U31612 (N_31612,N_30772,N_30985);
and U31613 (N_31613,N_30186,N_30292);
nor U31614 (N_31614,N_30392,N_30089);
nor U31615 (N_31615,N_30304,N_30989);
nand U31616 (N_31616,N_30953,N_30616);
nand U31617 (N_31617,N_30602,N_30755);
nand U31618 (N_31618,N_30126,N_30399);
nor U31619 (N_31619,N_30032,N_30986);
xnor U31620 (N_31620,N_30879,N_30952);
or U31621 (N_31621,N_30162,N_30572);
and U31622 (N_31622,N_30658,N_30174);
and U31623 (N_31623,N_30939,N_30931);
nor U31624 (N_31624,N_30416,N_30561);
xor U31625 (N_31625,N_30008,N_30035);
and U31626 (N_31626,N_30533,N_30372);
xor U31627 (N_31627,N_30542,N_30867);
nor U31628 (N_31628,N_30871,N_30217);
xnor U31629 (N_31629,N_30770,N_30651);
nand U31630 (N_31630,N_30979,N_30884);
nand U31631 (N_31631,N_30159,N_30400);
xnor U31632 (N_31632,N_30177,N_30665);
or U31633 (N_31633,N_30964,N_30327);
or U31634 (N_31634,N_30810,N_30205);
xor U31635 (N_31635,N_30469,N_30461);
nor U31636 (N_31636,N_30449,N_30398);
xor U31637 (N_31637,N_30139,N_30108);
and U31638 (N_31638,N_30045,N_30163);
nor U31639 (N_31639,N_30630,N_30859);
or U31640 (N_31640,N_30787,N_30666);
nor U31641 (N_31641,N_30033,N_30078);
and U31642 (N_31642,N_30019,N_30749);
nand U31643 (N_31643,N_30693,N_30116);
or U31644 (N_31644,N_30106,N_30535);
or U31645 (N_31645,N_30660,N_30304);
nand U31646 (N_31646,N_30043,N_30164);
nand U31647 (N_31647,N_30032,N_30583);
and U31648 (N_31648,N_30395,N_30906);
xor U31649 (N_31649,N_30994,N_30109);
nor U31650 (N_31650,N_30735,N_30153);
xor U31651 (N_31651,N_30574,N_30279);
nor U31652 (N_31652,N_30732,N_30207);
nor U31653 (N_31653,N_30544,N_30584);
nand U31654 (N_31654,N_30340,N_30434);
nand U31655 (N_31655,N_30998,N_30001);
nor U31656 (N_31656,N_30736,N_30989);
nand U31657 (N_31657,N_30013,N_30394);
nor U31658 (N_31658,N_30521,N_30425);
xor U31659 (N_31659,N_30260,N_30975);
nand U31660 (N_31660,N_30676,N_30411);
nand U31661 (N_31661,N_30279,N_30845);
and U31662 (N_31662,N_30590,N_30963);
xor U31663 (N_31663,N_30418,N_30532);
or U31664 (N_31664,N_30838,N_30642);
nand U31665 (N_31665,N_30656,N_30573);
nor U31666 (N_31666,N_30013,N_30450);
xnor U31667 (N_31667,N_30373,N_30020);
nand U31668 (N_31668,N_30079,N_30468);
xnor U31669 (N_31669,N_30533,N_30267);
and U31670 (N_31670,N_30869,N_30836);
xnor U31671 (N_31671,N_30923,N_30975);
nor U31672 (N_31672,N_30995,N_30162);
and U31673 (N_31673,N_30705,N_30513);
nand U31674 (N_31674,N_30863,N_30634);
nand U31675 (N_31675,N_30278,N_30491);
nand U31676 (N_31676,N_30936,N_30924);
or U31677 (N_31677,N_30093,N_30616);
nand U31678 (N_31678,N_30249,N_30363);
nor U31679 (N_31679,N_30305,N_30798);
nand U31680 (N_31680,N_30001,N_30950);
or U31681 (N_31681,N_30593,N_30412);
or U31682 (N_31682,N_30683,N_30554);
nor U31683 (N_31683,N_30900,N_30529);
nand U31684 (N_31684,N_30368,N_30724);
or U31685 (N_31685,N_30294,N_30571);
or U31686 (N_31686,N_30610,N_30514);
nor U31687 (N_31687,N_30855,N_30577);
nand U31688 (N_31688,N_30006,N_30301);
and U31689 (N_31689,N_30070,N_30488);
xor U31690 (N_31690,N_30291,N_30334);
or U31691 (N_31691,N_30357,N_30902);
nor U31692 (N_31692,N_30630,N_30608);
nor U31693 (N_31693,N_30022,N_30071);
or U31694 (N_31694,N_30914,N_30013);
and U31695 (N_31695,N_30925,N_30909);
and U31696 (N_31696,N_30195,N_30076);
nand U31697 (N_31697,N_30760,N_30318);
xor U31698 (N_31698,N_30152,N_30061);
and U31699 (N_31699,N_30830,N_30223);
or U31700 (N_31700,N_30425,N_30404);
and U31701 (N_31701,N_30463,N_30438);
xor U31702 (N_31702,N_30696,N_30307);
and U31703 (N_31703,N_30674,N_30242);
nor U31704 (N_31704,N_30019,N_30576);
xnor U31705 (N_31705,N_30105,N_30138);
nand U31706 (N_31706,N_30206,N_30741);
xor U31707 (N_31707,N_30625,N_30524);
xor U31708 (N_31708,N_30194,N_30263);
nand U31709 (N_31709,N_30641,N_30984);
nor U31710 (N_31710,N_30869,N_30642);
nor U31711 (N_31711,N_30326,N_30017);
xor U31712 (N_31712,N_30780,N_30316);
and U31713 (N_31713,N_30838,N_30883);
xnor U31714 (N_31714,N_30436,N_30501);
nor U31715 (N_31715,N_30621,N_30349);
or U31716 (N_31716,N_30306,N_30761);
xnor U31717 (N_31717,N_30349,N_30627);
or U31718 (N_31718,N_30114,N_30544);
and U31719 (N_31719,N_30618,N_30058);
xor U31720 (N_31720,N_30509,N_30460);
xnor U31721 (N_31721,N_30085,N_30217);
and U31722 (N_31722,N_30892,N_30820);
and U31723 (N_31723,N_30491,N_30149);
and U31724 (N_31724,N_30003,N_30621);
or U31725 (N_31725,N_30598,N_30954);
nand U31726 (N_31726,N_30840,N_30610);
and U31727 (N_31727,N_30727,N_30787);
nor U31728 (N_31728,N_30196,N_30390);
nand U31729 (N_31729,N_30698,N_30670);
nand U31730 (N_31730,N_30159,N_30736);
nand U31731 (N_31731,N_30167,N_30153);
nand U31732 (N_31732,N_30821,N_30949);
or U31733 (N_31733,N_30611,N_30563);
nand U31734 (N_31734,N_30031,N_30979);
or U31735 (N_31735,N_30413,N_30833);
xor U31736 (N_31736,N_30333,N_30567);
nor U31737 (N_31737,N_30765,N_30718);
nand U31738 (N_31738,N_30777,N_30257);
nand U31739 (N_31739,N_30442,N_30842);
xnor U31740 (N_31740,N_30331,N_30174);
or U31741 (N_31741,N_30634,N_30910);
xnor U31742 (N_31742,N_30560,N_30207);
nor U31743 (N_31743,N_30715,N_30624);
xor U31744 (N_31744,N_30611,N_30540);
xnor U31745 (N_31745,N_30590,N_30731);
xor U31746 (N_31746,N_30566,N_30327);
nand U31747 (N_31747,N_30940,N_30881);
nand U31748 (N_31748,N_30572,N_30647);
xnor U31749 (N_31749,N_30756,N_30296);
nand U31750 (N_31750,N_30290,N_30962);
and U31751 (N_31751,N_30709,N_30162);
nand U31752 (N_31752,N_30465,N_30385);
and U31753 (N_31753,N_30587,N_30454);
and U31754 (N_31754,N_30646,N_30310);
and U31755 (N_31755,N_30433,N_30444);
nand U31756 (N_31756,N_30829,N_30439);
or U31757 (N_31757,N_30125,N_30475);
xnor U31758 (N_31758,N_30659,N_30137);
nor U31759 (N_31759,N_30743,N_30929);
or U31760 (N_31760,N_30314,N_30063);
xor U31761 (N_31761,N_30293,N_30740);
xnor U31762 (N_31762,N_30645,N_30258);
xnor U31763 (N_31763,N_30341,N_30199);
nand U31764 (N_31764,N_30667,N_30798);
nand U31765 (N_31765,N_30730,N_30337);
and U31766 (N_31766,N_30892,N_30187);
nand U31767 (N_31767,N_30206,N_30993);
nand U31768 (N_31768,N_30806,N_30676);
or U31769 (N_31769,N_30925,N_30930);
nand U31770 (N_31770,N_30199,N_30750);
nand U31771 (N_31771,N_30796,N_30024);
xnor U31772 (N_31772,N_30410,N_30276);
nor U31773 (N_31773,N_30220,N_30553);
nor U31774 (N_31774,N_30606,N_30675);
xnor U31775 (N_31775,N_30840,N_30290);
xnor U31776 (N_31776,N_30392,N_30496);
and U31777 (N_31777,N_30191,N_30720);
or U31778 (N_31778,N_30018,N_30401);
xnor U31779 (N_31779,N_30066,N_30359);
and U31780 (N_31780,N_30938,N_30994);
nand U31781 (N_31781,N_30293,N_30311);
nor U31782 (N_31782,N_30296,N_30272);
and U31783 (N_31783,N_30946,N_30010);
xor U31784 (N_31784,N_30267,N_30532);
nor U31785 (N_31785,N_30963,N_30161);
nor U31786 (N_31786,N_30465,N_30980);
or U31787 (N_31787,N_30374,N_30183);
nor U31788 (N_31788,N_30864,N_30627);
nand U31789 (N_31789,N_30633,N_30819);
xor U31790 (N_31790,N_30436,N_30927);
xor U31791 (N_31791,N_30810,N_30586);
and U31792 (N_31792,N_30417,N_30607);
and U31793 (N_31793,N_30535,N_30745);
nand U31794 (N_31794,N_30806,N_30052);
or U31795 (N_31795,N_30854,N_30776);
xnor U31796 (N_31796,N_30608,N_30254);
and U31797 (N_31797,N_30793,N_30653);
nand U31798 (N_31798,N_30268,N_30785);
and U31799 (N_31799,N_30298,N_30278);
or U31800 (N_31800,N_30938,N_30110);
and U31801 (N_31801,N_30984,N_30025);
nand U31802 (N_31802,N_30118,N_30665);
and U31803 (N_31803,N_30233,N_30039);
and U31804 (N_31804,N_30995,N_30838);
or U31805 (N_31805,N_30166,N_30978);
and U31806 (N_31806,N_30744,N_30903);
nor U31807 (N_31807,N_30823,N_30195);
nand U31808 (N_31808,N_30028,N_30298);
or U31809 (N_31809,N_30389,N_30736);
nand U31810 (N_31810,N_30064,N_30872);
nor U31811 (N_31811,N_30460,N_30995);
or U31812 (N_31812,N_30464,N_30353);
nand U31813 (N_31813,N_30917,N_30223);
or U31814 (N_31814,N_30691,N_30569);
nor U31815 (N_31815,N_30073,N_30296);
or U31816 (N_31816,N_30057,N_30012);
xnor U31817 (N_31817,N_30291,N_30102);
or U31818 (N_31818,N_30580,N_30050);
and U31819 (N_31819,N_30500,N_30933);
xor U31820 (N_31820,N_30401,N_30362);
nor U31821 (N_31821,N_30404,N_30211);
xnor U31822 (N_31822,N_30117,N_30094);
nand U31823 (N_31823,N_30099,N_30688);
and U31824 (N_31824,N_30691,N_30171);
or U31825 (N_31825,N_30240,N_30082);
or U31826 (N_31826,N_30369,N_30218);
or U31827 (N_31827,N_30560,N_30113);
or U31828 (N_31828,N_30315,N_30311);
nor U31829 (N_31829,N_30372,N_30398);
and U31830 (N_31830,N_30518,N_30971);
and U31831 (N_31831,N_30193,N_30392);
xnor U31832 (N_31832,N_30849,N_30576);
xnor U31833 (N_31833,N_30646,N_30687);
nand U31834 (N_31834,N_30842,N_30574);
nand U31835 (N_31835,N_30229,N_30374);
and U31836 (N_31836,N_30716,N_30558);
nand U31837 (N_31837,N_30683,N_30558);
and U31838 (N_31838,N_30584,N_30792);
nor U31839 (N_31839,N_30972,N_30663);
and U31840 (N_31840,N_30561,N_30234);
nor U31841 (N_31841,N_30389,N_30861);
or U31842 (N_31842,N_30512,N_30590);
nor U31843 (N_31843,N_30088,N_30789);
and U31844 (N_31844,N_30760,N_30509);
nor U31845 (N_31845,N_30686,N_30262);
nand U31846 (N_31846,N_30407,N_30204);
and U31847 (N_31847,N_30138,N_30678);
nor U31848 (N_31848,N_30921,N_30881);
and U31849 (N_31849,N_30253,N_30192);
nor U31850 (N_31850,N_30477,N_30995);
and U31851 (N_31851,N_30385,N_30759);
or U31852 (N_31852,N_30133,N_30597);
or U31853 (N_31853,N_30954,N_30411);
nor U31854 (N_31854,N_30745,N_30036);
nor U31855 (N_31855,N_30549,N_30261);
nor U31856 (N_31856,N_30722,N_30256);
nand U31857 (N_31857,N_30965,N_30422);
xor U31858 (N_31858,N_30005,N_30272);
nand U31859 (N_31859,N_30004,N_30603);
nor U31860 (N_31860,N_30378,N_30499);
nand U31861 (N_31861,N_30546,N_30792);
nor U31862 (N_31862,N_30069,N_30075);
or U31863 (N_31863,N_30167,N_30724);
nor U31864 (N_31864,N_30398,N_30386);
xor U31865 (N_31865,N_30951,N_30112);
nor U31866 (N_31866,N_30443,N_30255);
nor U31867 (N_31867,N_30720,N_30842);
xnor U31868 (N_31868,N_30161,N_30919);
and U31869 (N_31869,N_30169,N_30512);
xor U31870 (N_31870,N_30354,N_30115);
and U31871 (N_31871,N_30087,N_30228);
or U31872 (N_31872,N_30603,N_30450);
nand U31873 (N_31873,N_30777,N_30064);
nand U31874 (N_31874,N_30784,N_30030);
nand U31875 (N_31875,N_30680,N_30286);
or U31876 (N_31876,N_30450,N_30191);
or U31877 (N_31877,N_30192,N_30564);
xor U31878 (N_31878,N_30216,N_30053);
nand U31879 (N_31879,N_30375,N_30026);
or U31880 (N_31880,N_30351,N_30900);
nor U31881 (N_31881,N_30228,N_30893);
xor U31882 (N_31882,N_30809,N_30191);
nor U31883 (N_31883,N_30828,N_30271);
and U31884 (N_31884,N_30197,N_30788);
or U31885 (N_31885,N_30639,N_30300);
xor U31886 (N_31886,N_30707,N_30941);
and U31887 (N_31887,N_30702,N_30575);
or U31888 (N_31888,N_30188,N_30788);
or U31889 (N_31889,N_30030,N_30289);
nor U31890 (N_31890,N_30904,N_30647);
and U31891 (N_31891,N_30485,N_30605);
and U31892 (N_31892,N_30396,N_30460);
nor U31893 (N_31893,N_30324,N_30338);
and U31894 (N_31894,N_30568,N_30048);
or U31895 (N_31895,N_30139,N_30519);
nand U31896 (N_31896,N_30924,N_30062);
nand U31897 (N_31897,N_30610,N_30301);
nor U31898 (N_31898,N_30543,N_30615);
xnor U31899 (N_31899,N_30797,N_30491);
nor U31900 (N_31900,N_30469,N_30096);
xor U31901 (N_31901,N_30212,N_30549);
xnor U31902 (N_31902,N_30913,N_30706);
xnor U31903 (N_31903,N_30536,N_30712);
xor U31904 (N_31904,N_30320,N_30289);
or U31905 (N_31905,N_30562,N_30893);
nand U31906 (N_31906,N_30670,N_30370);
nor U31907 (N_31907,N_30720,N_30790);
nand U31908 (N_31908,N_30873,N_30546);
and U31909 (N_31909,N_30513,N_30918);
xnor U31910 (N_31910,N_30142,N_30881);
or U31911 (N_31911,N_30535,N_30002);
or U31912 (N_31912,N_30920,N_30254);
or U31913 (N_31913,N_30448,N_30302);
or U31914 (N_31914,N_30724,N_30758);
nor U31915 (N_31915,N_30247,N_30989);
or U31916 (N_31916,N_30976,N_30376);
xor U31917 (N_31917,N_30547,N_30910);
nor U31918 (N_31918,N_30312,N_30945);
nor U31919 (N_31919,N_30553,N_30367);
nand U31920 (N_31920,N_30478,N_30042);
or U31921 (N_31921,N_30725,N_30737);
xnor U31922 (N_31922,N_30268,N_30060);
nor U31923 (N_31923,N_30735,N_30537);
nor U31924 (N_31924,N_30648,N_30057);
nor U31925 (N_31925,N_30665,N_30647);
or U31926 (N_31926,N_30572,N_30225);
xor U31927 (N_31927,N_30254,N_30069);
nand U31928 (N_31928,N_30993,N_30681);
and U31929 (N_31929,N_30270,N_30857);
or U31930 (N_31930,N_30846,N_30450);
nor U31931 (N_31931,N_30645,N_30104);
xor U31932 (N_31932,N_30229,N_30561);
or U31933 (N_31933,N_30032,N_30131);
or U31934 (N_31934,N_30582,N_30086);
xor U31935 (N_31935,N_30694,N_30369);
nor U31936 (N_31936,N_30204,N_30125);
nor U31937 (N_31937,N_30114,N_30126);
nor U31938 (N_31938,N_30725,N_30960);
or U31939 (N_31939,N_30443,N_30196);
nor U31940 (N_31940,N_30012,N_30659);
xnor U31941 (N_31941,N_30001,N_30548);
and U31942 (N_31942,N_30366,N_30249);
xor U31943 (N_31943,N_30114,N_30976);
xor U31944 (N_31944,N_30060,N_30309);
and U31945 (N_31945,N_30883,N_30616);
nor U31946 (N_31946,N_30302,N_30402);
and U31947 (N_31947,N_30563,N_30873);
or U31948 (N_31948,N_30513,N_30437);
nor U31949 (N_31949,N_30702,N_30699);
or U31950 (N_31950,N_30779,N_30836);
or U31951 (N_31951,N_30992,N_30490);
or U31952 (N_31952,N_30574,N_30147);
and U31953 (N_31953,N_30161,N_30632);
nor U31954 (N_31954,N_30356,N_30285);
and U31955 (N_31955,N_30428,N_30812);
nor U31956 (N_31956,N_30120,N_30754);
and U31957 (N_31957,N_30855,N_30516);
nor U31958 (N_31958,N_30282,N_30242);
xor U31959 (N_31959,N_30284,N_30522);
xor U31960 (N_31960,N_30729,N_30053);
nand U31961 (N_31961,N_30294,N_30651);
and U31962 (N_31962,N_30923,N_30260);
and U31963 (N_31963,N_30965,N_30452);
or U31964 (N_31964,N_30563,N_30647);
nor U31965 (N_31965,N_30374,N_30601);
or U31966 (N_31966,N_30544,N_30496);
nand U31967 (N_31967,N_30889,N_30249);
and U31968 (N_31968,N_30212,N_30408);
or U31969 (N_31969,N_30268,N_30965);
and U31970 (N_31970,N_30698,N_30237);
or U31971 (N_31971,N_30289,N_30284);
xor U31972 (N_31972,N_30183,N_30568);
nand U31973 (N_31973,N_30109,N_30169);
nor U31974 (N_31974,N_30893,N_30503);
or U31975 (N_31975,N_30692,N_30004);
nor U31976 (N_31976,N_30179,N_30136);
or U31977 (N_31977,N_30445,N_30016);
nand U31978 (N_31978,N_30849,N_30593);
or U31979 (N_31979,N_30087,N_30837);
xnor U31980 (N_31980,N_30146,N_30865);
xnor U31981 (N_31981,N_30205,N_30404);
xor U31982 (N_31982,N_30785,N_30729);
nor U31983 (N_31983,N_30571,N_30145);
or U31984 (N_31984,N_30383,N_30750);
xor U31985 (N_31985,N_30591,N_30985);
or U31986 (N_31986,N_30025,N_30640);
and U31987 (N_31987,N_30808,N_30103);
or U31988 (N_31988,N_30661,N_30033);
and U31989 (N_31989,N_30947,N_30244);
or U31990 (N_31990,N_30515,N_30875);
xor U31991 (N_31991,N_30872,N_30631);
nand U31992 (N_31992,N_30892,N_30214);
xnor U31993 (N_31993,N_30996,N_30581);
xor U31994 (N_31994,N_30826,N_30647);
and U31995 (N_31995,N_30586,N_30666);
xor U31996 (N_31996,N_30007,N_30315);
nand U31997 (N_31997,N_30055,N_30813);
and U31998 (N_31998,N_30636,N_30164);
and U31999 (N_31999,N_30120,N_30879);
nor U32000 (N_32000,N_31241,N_31236);
xor U32001 (N_32001,N_31436,N_31254);
or U32002 (N_32002,N_31712,N_31710);
xor U32003 (N_32003,N_31224,N_31217);
xor U32004 (N_32004,N_31315,N_31935);
xor U32005 (N_32005,N_31419,N_31119);
or U32006 (N_32006,N_31028,N_31588);
and U32007 (N_32007,N_31742,N_31370);
nand U32008 (N_32008,N_31335,N_31507);
and U32009 (N_32009,N_31936,N_31675);
nand U32010 (N_32010,N_31100,N_31910);
nor U32011 (N_32011,N_31685,N_31841);
xnor U32012 (N_32012,N_31558,N_31459);
nor U32013 (N_32013,N_31299,N_31662);
and U32014 (N_32014,N_31041,N_31914);
nor U32015 (N_32015,N_31819,N_31622);
xnor U32016 (N_32016,N_31255,N_31748);
nand U32017 (N_32017,N_31294,N_31767);
and U32018 (N_32018,N_31930,N_31725);
nor U32019 (N_32019,N_31623,N_31238);
and U32020 (N_32020,N_31406,N_31133);
nand U32021 (N_32021,N_31547,N_31153);
xor U32022 (N_32022,N_31503,N_31145);
nand U32023 (N_32023,N_31293,N_31468);
and U32024 (N_32024,N_31773,N_31491);
nand U32025 (N_32025,N_31209,N_31783);
or U32026 (N_32026,N_31178,N_31303);
nor U32027 (N_32027,N_31235,N_31135);
xor U32028 (N_32028,N_31518,N_31475);
or U32029 (N_32029,N_31489,N_31581);
nand U32030 (N_32030,N_31388,N_31892);
or U32031 (N_32031,N_31340,N_31015);
and U32032 (N_32032,N_31760,N_31152);
nand U32033 (N_32033,N_31321,N_31789);
and U32034 (N_32034,N_31988,N_31213);
or U32035 (N_32035,N_31441,N_31927);
nand U32036 (N_32036,N_31312,N_31182);
nor U32037 (N_32037,N_31113,N_31267);
xor U32038 (N_32038,N_31449,N_31647);
nor U32039 (N_32039,N_31517,N_31967);
xor U32040 (N_32040,N_31323,N_31928);
and U32041 (N_32041,N_31476,N_31649);
nand U32042 (N_32042,N_31895,N_31657);
or U32043 (N_32043,N_31477,N_31852);
or U32044 (N_32044,N_31328,N_31885);
and U32045 (N_32045,N_31242,N_31557);
nand U32046 (N_32046,N_31362,N_31204);
or U32047 (N_32047,N_31250,N_31755);
and U32048 (N_32048,N_31521,N_31946);
and U32049 (N_32049,N_31126,N_31976);
xnor U32050 (N_32050,N_31114,N_31600);
xor U32051 (N_32051,N_31369,N_31799);
nor U32052 (N_32052,N_31616,N_31906);
and U32053 (N_32053,N_31563,N_31635);
xnor U32054 (N_32054,N_31107,N_31764);
xor U32055 (N_32055,N_31684,N_31593);
nor U32056 (N_32056,N_31103,N_31645);
nand U32057 (N_32057,N_31448,N_31637);
nor U32058 (N_32058,N_31161,N_31019);
nand U32059 (N_32059,N_31543,N_31598);
and U32060 (N_32060,N_31067,N_31035);
or U32061 (N_32061,N_31822,N_31246);
or U32062 (N_32062,N_31160,N_31724);
nand U32063 (N_32063,N_31354,N_31347);
and U32064 (N_32064,N_31751,N_31458);
nor U32065 (N_32065,N_31351,N_31384);
and U32066 (N_32066,N_31147,N_31956);
nor U32067 (N_32067,N_31648,N_31229);
nand U32068 (N_32068,N_31486,N_31579);
xor U32069 (N_32069,N_31508,N_31814);
nand U32070 (N_32070,N_31654,N_31118);
and U32071 (N_32071,N_31903,N_31284);
or U32072 (N_32072,N_31410,N_31442);
or U32073 (N_32073,N_31296,N_31257);
nand U32074 (N_32074,N_31243,N_31465);
nor U32075 (N_32075,N_31047,N_31539);
xor U32076 (N_32076,N_31317,N_31225);
and U32077 (N_32077,N_31496,N_31787);
xnor U32078 (N_32078,N_31151,N_31377);
nand U32079 (N_32079,N_31332,N_31427);
and U32080 (N_32080,N_31553,N_31909);
nor U32081 (N_32081,N_31298,N_31269);
or U32082 (N_32082,N_31173,N_31105);
nor U32083 (N_32083,N_31717,N_31215);
or U32084 (N_32084,N_31848,N_31096);
xnor U32085 (N_32085,N_31037,N_31313);
and U32086 (N_32086,N_31044,N_31308);
xnor U32087 (N_32087,N_31820,N_31580);
nand U32088 (N_32088,N_31502,N_31682);
and U32089 (N_32089,N_31847,N_31853);
or U32090 (N_32090,N_31971,N_31206);
or U32091 (N_32091,N_31450,N_31703);
nand U32092 (N_32092,N_31858,N_31075);
nand U32093 (N_32093,N_31098,N_31271);
xor U32094 (N_32094,N_31346,N_31387);
nand U32095 (N_32095,N_31955,N_31097);
xnor U32096 (N_32096,N_31739,N_31089);
nand U32097 (N_32097,N_31584,N_31365);
and U32098 (N_32098,N_31921,N_31112);
nand U32099 (N_32099,N_31690,N_31643);
nor U32100 (N_32100,N_31537,N_31569);
and U32101 (N_32101,N_31551,N_31827);
nor U32102 (N_32102,N_31883,N_31433);
nand U32103 (N_32103,N_31493,N_31179);
or U32104 (N_32104,N_31626,N_31741);
and U32105 (N_32105,N_31793,N_31149);
or U32106 (N_32106,N_31248,N_31472);
or U32107 (N_32107,N_31252,N_31779);
nor U32108 (N_32108,N_31355,N_31263);
and U32109 (N_32109,N_31307,N_31786);
xnor U32110 (N_32110,N_31667,N_31878);
and U32111 (N_32111,N_31265,N_31951);
and U32112 (N_32112,N_31838,N_31804);
nand U32113 (N_32113,N_31031,N_31210);
or U32114 (N_32114,N_31691,N_31713);
and U32115 (N_32115,N_31368,N_31898);
or U32116 (N_32116,N_31631,N_31360);
or U32117 (N_32117,N_31302,N_31201);
xnor U32118 (N_32118,N_31064,N_31027);
nor U32119 (N_32119,N_31524,N_31777);
nand U32120 (N_32120,N_31234,N_31745);
or U32121 (N_32121,N_31942,N_31208);
nand U32122 (N_32122,N_31081,N_31871);
nor U32123 (N_32123,N_31451,N_31619);
nand U32124 (N_32124,N_31632,N_31156);
nor U32125 (N_32125,N_31911,N_31708);
nand U32126 (N_32126,N_31919,N_31576);
nor U32127 (N_32127,N_31912,N_31385);
xnor U32128 (N_32128,N_31146,N_31494);
and U32129 (N_32129,N_31072,N_31945);
or U32130 (N_32130,N_31087,N_31615);
xor U32131 (N_32131,N_31875,N_31050);
and U32132 (N_32132,N_31851,N_31661);
nand U32133 (N_32133,N_31900,N_31595);
nor U32134 (N_32134,N_31653,N_31348);
nor U32135 (N_32135,N_31761,N_31404);
nor U32136 (N_32136,N_31401,N_31994);
and U32137 (N_32137,N_31000,N_31642);
or U32138 (N_32138,N_31197,N_31108);
and U32139 (N_32139,N_31589,N_31556);
nand U32140 (N_32140,N_31809,N_31093);
nor U32141 (N_32141,N_31915,N_31253);
xor U32142 (N_32142,N_31621,N_31057);
or U32143 (N_32143,N_31357,N_31538);
nand U32144 (N_32144,N_31830,N_31240);
xnor U32145 (N_32145,N_31414,N_31350);
and U32146 (N_32146,N_31867,N_31002);
or U32147 (N_32147,N_31017,N_31609);
or U32148 (N_32148,N_31053,N_31762);
nor U32149 (N_32149,N_31484,N_31567);
and U32150 (N_32150,N_31702,N_31523);
and U32151 (N_32151,N_31715,N_31397);
nor U32152 (N_32152,N_31226,N_31172);
nand U32153 (N_32153,N_31689,N_31099);
nand U32154 (N_32154,N_31826,N_31954);
nand U32155 (N_32155,N_31602,N_31984);
nor U32156 (N_32156,N_31409,N_31203);
and U32157 (N_32157,N_31310,N_31925);
xor U32158 (N_32158,N_31260,N_31636);
or U32159 (N_32159,N_31601,N_31222);
xor U32160 (N_32160,N_31991,N_31627);
xor U32161 (N_32161,N_31012,N_31613);
xnor U32162 (N_32162,N_31599,N_31926);
and U32163 (N_32163,N_31447,N_31824);
nor U32164 (N_32164,N_31273,N_31375);
or U32165 (N_32165,N_31190,N_31233);
or U32166 (N_32166,N_31688,N_31757);
and U32167 (N_32167,N_31681,N_31902);
xnor U32168 (N_32168,N_31586,N_31756);
or U32169 (N_32169,N_31083,N_31987);
nand U32170 (N_32170,N_31931,N_31535);
or U32171 (N_32171,N_31192,N_31032);
or U32172 (N_32172,N_31174,N_31102);
or U32173 (N_32173,N_31191,N_31356);
xnor U32174 (N_32174,N_31542,N_31262);
nor U32175 (N_32175,N_31221,N_31776);
nand U32176 (N_32176,N_31300,N_31337);
xnor U32177 (N_32177,N_31792,N_31747);
xor U32178 (N_32178,N_31358,N_31698);
or U32179 (N_32179,N_31443,N_31051);
and U32180 (N_32180,N_31887,N_31620);
and U32181 (N_32181,N_31614,N_31658);
nand U32182 (N_32182,N_31177,N_31500);
or U32183 (N_32183,N_31295,N_31343);
nor U32184 (N_32184,N_31574,N_31975);
nand U32185 (N_32185,N_31664,N_31407);
or U32186 (N_32186,N_31752,N_31923);
and U32187 (N_32187,N_31120,N_31292);
and U32188 (N_32188,N_31430,N_31495);
xnor U32189 (N_32189,N_31216,N_31726);
and U32190 (N_32190,N_31391,N_31680);
and U32191 (N_32191,N_31142,N_31837);
xor U32192 (N_32192,N_31398,N_31711);
xor U32193 (N_32193,N_31462,N_31929);
and U32194 (N_32194,N_31048,N_31036);
nor U32195 (N_32195,N_31924,N_31979);
and U32196 (N_32196,N_31533,N_31882);
and U32197 (N_32197,N_31150,N_31772);
and U32198 (N_32198,N_31554,N_31270);
or U32199 (N_32199,N_31256,N_31080);
nor U32200 (N_32200,N_31808,N_31810);
nor U32201 (N_32201,N_31677,N_31816);
nand U32202 (N_32202,N_31129,N_31237);
or U32203 (N_32203,N_31536,N_31952);
or U32204 (N_32204,N_31501,N_31605);
nor U32205 (N_32205,N_31003,N_31873);
and U32206 (N_32206,N_31437,N_31577);
nor U32207 (N_32207,N_31422,N_31386);
and U32208 (N_32208,N_31683,N_31498);
and U32209 (N_32209,N_31587,N_31066);
nand U32210 (N_32210,N_31941,N_31947);
or U32211 (N_32211,N_31176,N_31288);
nor U32212 (N_32212,N_31978,N_31272);
nand U32213 (N_32213,N_31797,N_31042);
nand U32214 (N_32214,N_31718,N_31162);
nor U32215 (N_32215,N_31261,N_31652);
nand U32216 (N_32216,N_31069,N_31466);
or U32217 (N_32217,N_31548,N_31877);
nand U32218 (N_32218,N_31095,N_31429);
xor U32219 (N_32219,N_31399,N_31479);
or U32220 (N_32220,N_31734,N_31559);
and U32221 (N_32221,N_31467,N_31607);
and U32222 (N_32222,N_31106,N_31231);
nor U32223 (N_32223,N_31396,N_31336);
nor U32224 (N_32224,N_31771,N_31525);
nor U32225 (N_32225,N_31737,N_31639);
or U32226 (N_32226,N_31074,N_31738);
nor U32227 (N_32227,N_31169,N_31371);
nand U32228 (N_32228,N_31101,N_31259);
xnor U32229 (N_32229,N_31730,N_31800);
nor U32230 (N_32230,N_31727,N_31412);
nand U32231 (N_32231,N_31117,N_31416);
or U32232 (N_32232,N_31531,N_31520);
nand U32233 (N_32233,N_31469,N_31076);
xor U32234 (N_32234,N_31965,N_31038);
nor U32235 (N_32235,N_31832,N_31431);
or U32236 (N_32236,N_31891,N_31045);
xnor U32237 (N_32237,N_31749,N_31140);
xor U32238 (N_32238,N_31194,N_31818);
or U32239 (N_32239,N_31624,N_31562);
and U32240 (N_32240,N_31471,N_31361);
or U32241 (N_32241,N_31839,N_31608);
or U32242 (N_32242,N_31457,N_31700);
or U32243 (N_32243,N_31957,N_31784);
and U32244 (N_32244,N_31944,N_31940);
nand U32245 (N_32245,N_31446,N_31813);
nand U32246 (N_32246,N_31707,N_31993);
nand U32247 (N_32247,N_31187,N_31011);
nand U32248 (N_32248,N_31803,N_31181);
xor U32249 (N_32249,N_31731,N_31905);
or U32250 (N_32250,N_31281,N_31372);
nand U32251 (N_32251,N_31546,N_31342);
or U32252 (N_32252,N_31175,N_31382);
and U32253 (N_32253,N_31844,N_31277);
xor U32254 (N_32254,N_31716,N_31408);
xnor U32255 (N_32255,N_31025,N_31750);
nand U32256 (N_32256,N_31363,N_31625);
or U32257 (N_32257,N_31040,N_31485);
nand U32258 (N_32258,N_31068,N_31515);
and U32259 (N_32259,N_31132,N_31630);
nor U32260 (N_32260,N_31165,N_31781);
nand U32261 (N_32261,N_31456,N_31163);
xnor U32262 (N_32262,N_31864,N_31510);
nor U32263 (N_32263,N_31001,N_31141);
xor U32264 (N_32264,N_31913,N_31973);
xnor U32265 (N_32265,N_31950,N_31374);
and U32266 (N_32266,N_31088,N_31529);
or U32267 (N_32267,N_31247,N_31733);
or U32268 (N_32268,N_31695,N_31744);
nand U32269 (N_32269,N_31540,N_31344);
nor U32270 (N_32270,N_31629,N_31960);
nor U32271 (N_32271,N_31030,N_31334);
nor U32272 (N_32272,N_31815,N_31918);
nor U32273 (N_32273,N_31782,N_31005);
or U32274 (N_32274,N_31908,N_31568);
xor U32275 (N_32275,N_31056,N_31861);
nor U32276 (N_32276,N_31981,N_31555);
or U32277 (N_32277,N_31154,N_31167);
nand U32278 (N_32278,N_31802,N_31244);
nand U32279 (N_32279,N_31010,N_31856);
xor U32280 (N_32280,N_31701,N_31729);
nand U32281 (N_32281,N_31881,N_31478);
nor U32282 (N_32282,N_31322,N_31159);
or U32283 (N_32283,N_31704,N_31660);
and U32284 (N_32284,N_31998,N_31301);
nand U32285 (N_32285,N_31470,N_31732);
xor U32286 (N_32286,N_31862,N_31638);
xnor U32287 (N_32287,N_31673,N_31612);
and U32288 (N_32288,N_31541,N_31420);
and U32289 (N_32289,N_31582,N_31668);
nor U32290 (N_32290,N_31144,N_31591);
nor U32291 (N_32291,N_31227,N_31021);
or U32292 (N_32292,N_31986,N_31434);
and U32293 (N_32293,N_31880,N_31046);
xor U32294 (N_32294,N_31890,N_31610);
xnor U32295 (N_32295,N_31290,N_31659);
or U32296 (N_32296,N_31872,N_31364);
and U32297 (N_32297,N_31214,N_31383);
nor U32298 (N_32298,N_31759,N_31884);
nand U32299 (N_32299,N_31780,N_31833);
nand U32300 (N_32300,N_31999,N_31969);
xnor U32301 (N_32301,N_31709,N_31943);
xor U32302 (N_32302,N_31868,N_31338);
or U32303 (N_32303,N_31527,N_31306);
nor U32304 (N_32304,N_31352,N_31611);
or U32305 (N_32305,N_31575,N_31220);
and U32306 (N_32306,N_31073,N_31394);
nand U32307 (N_32307,N_31488,N_31171);
or U32308 (N_32308,N_31544,N_31128);
nand U32309 (N_32309,N_31345,N_31696);
xnor U32310 (N_32310,N_31378,N_31843);
and U32311 (N_32311,N_31679,N_31874);
and U32312 (N_32312,N_31245,N_31722);
and U32313 (N_32313,N_31060,N_31440);
xor U32314 (N_32314,N_31740,N_31428);
or U32315 (N_32315,N_31617,N_31086);
nor U32316 (N_32316,N_31164,N_31723);
and U32317 (N_32317,N_31148,N_31481);
nor U32318 (N_32318,N_31655,N_31699);
nor U32319 (N_32319,N_31676,N_31207);
xor U32320 (N_32320,N_31033,N_31970);
or U32321 (N_32321,N_31678,N_31445);
and U32322 (N_32322,N_31949,N_31550);
and U32323 (N_32323,N_31403,N_31644);
xor U32324 (N_32324,N_31180,N_31850);
and U32325 (N_32325,N_31845,N_31893);
and U32326 (N_32326,N_31886,N_31061);
xnor U32327 (N_32327,N_31251,N_31721);
nor U32328 (N_32328,N_31219,N_31687);
nor U32329 (N_32329,N_31425,N_31139);
xor U32330 (N_32330,N_31094,N_31506);
xor U32331 (N_32331,N_31656,N_31013);
nand U32332 (N_32332,N_31314,N_31438);
and U32333 (N_32333,N_31560,N_31669);
xor U32334 (N_32334,N_31821,N_31009);
xor U32335 (N_32335,N_31865,N_31239);
xnor U32336 (N_32336,N_31572,N_31665);
nor U32337 (N_32337,N_31166,N_31590);
xor U32338 (N_32338,N_31327,N_31855);
xor U32339 (N_32339,N_31463,N_31058);
or U32340 (N_32340,N_31258,N_31202);
and U32341 (N_32341,N_31170,N_31798);
or U32342 (N_32342,N_31024,N_31788);
nor U32343 (N_32343,N_31565,N_31116);
xnor U32344 (N_32344,N_31423,N_31325);
and U32345 (N_32345,N_31817,N_31519);
xnor U32346 (N_32346,N_31829,N_31333);
and U32347 (N_32347,N_31534,N_31395);
nand U32348 (N_32348,N_31136,N_31860);
and U32349 (N_32349,N_31505,N_31266);
and U32350 (N_32350,N_31052,N_31794);
nor U32351 (N_32351,N_31131,N_31007);
nor U32352 (N_32352,N_31522,N_31079);
nand U32353 (N_32353,N_31483,N_31938);
and U32354 (N_32354,N_31359,N_31415);
or U32355 (N_32355,N_31907,N_31373);
or U32356 (N_32356,N_31487,N_31380);
xnor U32357 (N_32357,N_31719,N_31592);
nand U32358 (N_32358,N_31863,N_31492);
or U32359 (N_32359,N_31426,N_31670);
xor U32360 (N_32360,N_31029,N_31720);
xor U32361 (N_32361,N_31922,N_31846);
and U32362 (N_32362,N_31071,N_31806);
or U32363 (N_32363,N_31996,N_31917);
nor U32364 (N_32364,N_31020,N_31916);
nor U32365 (N_32365,N_31249,N_31432);
or U32366 (N_32366,N_31795,N_31444);
xnor U32367 (N_32367,N_31694,N_31276);
or U32368 (N_32368,N_31990,N_31801);
nor U32369 (N_32369,N_31513,N_31995);
and U32370 (N_32370,N_31157,N_31278);
and U32371 (N_32371,N_31183,N_31530);
xor U32372 (N_32372,N_31212,N_31275);
nor U32373 (N_32373,N_31974,N_31758);
xor U32374 (N_32374,N_31305,N_31583);
xnor U32375 (N_32375,N_31511,N_31353);
nor U32376 (N_32376,N_31418,N_31796);
nor U32377 (N_32377,N_31084,N_31980);
xor U32378 (N_32378,N_31211,N_31200);
and U32379 (N_32379,N_31115,N_31320);
nor U32380 (N_32380,N_31640,N_31666);
and U32381 (N_32381,N_31596,N_31143);
nor U32382 (N_32382,N_31859,N_31034);
nor U32383 (N_32383,N_31082,N_31769);
or U32384 (N_32384,N_31514,N_31566);
or U32385 (N_32385,N_31285,N_31381);
nand U32386 (N_32386,N_31366,N_31393);
or U32387 (N_32387,N_31823,N_31497);
xor U32388 (N_32388,N_31920,N_31022);
nand U32389 (N_32389,N_31904,N_31754);
and U32390 (N_32390,N_31571,N_31532);
nand U32391 (N_32391,N_31791,N_31641);
xnor U32392 (N_32392,N_31196,N_31585);
and U32393 (N_32393,N_31078,N_31706);
nand U32394 (N_32394,N_31043,N_31090);
or U32395 (N_32395,N_31953,N_31059);
or U32396 (N_32396,N_31834,N_31774);
and U32397 (N_32397,N_31512,N_31528);
or U32398 (N_32398,N_31339,N_31123);
xor U32399 (N_32399,N_31070,N_31134);
and U32400 (N_32400,N_31693,N_31894);
and U32401 (N_32401,N_31121,N_31473);
xor U32402 (N_32402,N_31650,N_31932);
nand U32403 (N_32403,N_31122,N_31026);
or U32404 (N_32404,N_31634,N_31606);
nand U32405 (N_32405,N_31876,N_31937);
or U32406 (N_32406,N_31453,N_31091);
xnor U32407 (N_32407,N_31092,N_31870);
nor U32408 (N_32408,N_31016,N_31006);
or U32409 (N_32409,N_31109,N_31085);
nor U32410 (N_32410,N_31223,N_31111);
nand U32411 (N_32411,N_31018,N_31198);
nor U32412 (N_32412,N_31618,N_31933);
xor U32413 (N_32413,N_31454,N_31633);
or U32414 (N_32414,N_31104,N_31743);
nand U32415 (N_32415,N_31379,N_31959);
nor U32416 (N_32416,N_31274,N_31297);
and U32417 (N_32417,N_31948,N_31735);
xor U32418 (N_32418,N_31768,N_31869);
xnor U32419 (N_32419,N_31474,N_31480);
or U32420 (N_32420,N_31286,N_31746);
and U32421 (N_32421,N_31705,N_31836);
nor U32422 (N_32422,N_31509,N_31455);
nand U32423 (N_32423,N_31594,N_31966);
nor U32424 (N_32424,N_31977,N_31766);
and U32425 (N_32425,N_31205,N_31840);
or U32426 (N_32426,N_31697,N_31763);
xnor U32427 (N_32427,N_31324,N_31831);
nand U32428 (N_32428,N_31304,N_31228);
and U32429 (N_32429,N_31127,N_31264);
nor U32430 (N_32430,N_31311,N_31055);
nor U32431 (N_32431,N_31331,N_31125);
or U32432 (N_32432,N_31597,N_31997);
xor U32433 (N_32433,N_31663,N_31482);
nand U32434 (N_32434,N_31155,N_31189);
nor U32435 (N_32435,N_31138,N_31842);
xnor U32436 (N_32436,N_31545,N_31291);
nor U32437 (N_32437,N_31674,N_31158);
xor U32438 (N_32438,N_31417,N_31199);
nand U32439 (N_32439,N_31460,N_31400);
and U32440 (N_32440,N_31790,N_31828);
nor U32441 (N_32441,N_31854,N_31014);
xor U32442 (N_32442,N_31232,N_31807);
and U32443 (N_32443,N_31958,N_31464);
and U32444 (N_32444,N_31962,N_31062);
xnor U32445 (N_32445,N_31785,N_31686);
xnor U32446 (N_32446,N_31023,N_31499);
xor U32447 (N_32447,N_31490,N_31218);
or U32448 (N_32448,N_31516,N_31972);
xor U32449 (N_32449,N_31318,N_31889);
xnor U32450 (N_32450,N_31753,N_31603);
nor U32451 (N_32451,N_31054,N_31065);
and U32452 (N_32452,N_31341,N_31063);
or U32453 (N_32453,N_31435,N_31736);
nand U32454 (N_32454,N_31287,N_31628);
and U32455 (N_32455,N_31390,N_31982);
or U32456 (N_32456,N_31901,N_31039);
or U32457 (N_32457,N_31309,N_31985);
and U32458 (N_32458,N_31413,N_31367);
nand U32459 (N_32459,N_31421,N_31411);
or U32460 (N_32460,N_31825,N_31268);
nor U32461 (N_32461,N_31184,N_31230);
or U32462 (N_32462,N_31578,N_31714);
xnor U32463 (N_32463,N_31195,N_31004);
and U32464 (N_32464,N_31646,N_31124);
xnor U32465 (N_32465,N_31552,N_31775);
nor U32466 (N_32466,N_31983,N_31692);
xnor U32467 (N_32467,N_31137,N_31186);
or U32468 (N_32468,N_31963,N_31168);
and U32469 (N_32469,N_31879,N_31961);
xor U32470 (N_32470,N_31193,N_31805);
and U32471 (N_32471,N_31282,N_31049);
and U32472 (N_32472,N_31326,N_31778);
or U32473 (N_32473,N_31405,N_31329);
or U32474 (N_32474,N_31564,N_31188);
xnor U32475 (N_32475,N_31283,N_31077);
and U32476 (N_32476,N_31316,N_31439);
and U32477 (N_32477,N_31008,N_31934);
nor U32478 (N_32478,N_31604,N_31899);
xnor U32479 (N_32479,N_31835,N_31319);
xor U32480 (N_32480,N_31349,N_31992);
or U32481 (N_32481,N_31765,N_31728);
and U32482 (N_32482,N_31968,N_31812);
or U32483 (N_32483,N_31811,N_31573);
and U32484 (N_32484,N_31461,N_31964);
nand U32485 (N_32485,N_31452,N_31989);
xor U32486 (N_32486,N_31939,N_31130);
xor U32487 (N_32487,N_31849,N_31330);
and U32488 (N_32488,N_31896,N_31570);
nand U32489 (N_32489,N_31897,N_31279);
nor U32490 (N_32490,N_31389,N_31402);
xnor U32491 (N_32491,N_31504,N_31857);
or U32492 (N_32492,N_31392,N_31280);
and U32493 (N_32493,N_31866,N_31561);
nor U32494 (N_32494,N_31424,N_31888);
and U32495 (N_32495,N_31526,N_31651);
and U32496 (N_32496,N_31289,N_31110);
or U32497 (N_32497,N_31770,N_31376);
and U32498 (N_32498,N_31549,N_31671);
or U32499 (N_32499,N_31672,N_31185);
and U32500 (N_32500,N_31015,N_31105);
nor U32501 (N_32501,N_31261,N_31847);
and U32502 (N_32502,N_31577,N_31598);
nand U32503 (N_32503,N_31763,N_31810);
nor U32504 (N_32504,N_31802,N_31047);
xnor U32505 (N_32505,N_31553,N_31493);
nand U32506 (N_32506,N_31539,N_31098);
nor U32507 (N_32507,N_31544,N_31751);
nor U32508 (N_32508,N_31719,N_31578);
nand U32509 (N_32509,N_31634,N_31618);
xor U32510 (N_32510,N_31997,N_31628);
or U32511 (N_32511,N_31479,N_31627);
nand U32512 (N_32512,N_31074,N_31865);
nor U32513 (N_32513,N_31083,N_31401);
nand U32514 (N_32514,N_31472,N_31036);
nand U32515 (N_32515,N_31960,N_31713);
xor U32516 (N_32516,N_31438,N_31738);
nor U32517 (N_32517,N_31270,N_31294);
and U32518 (N_32518,N_31689,N_31302);
and U32519 (N_32519,N_31040,N_31532);
xor U32520 (N_32520,N_31528,N_31926);
nor U32521 (N_32521,N_31632,N_31691);
nand U32522 (N_32522,N_31620,N_31385);
or U32523 (N_32523,N_31757,N_31616);
nor U32524 (N_32524,N_31719,N_31133);
nor U32525 (N_32525,N_31157,N_31136);
xnor U32526 (N_32526,N_31544,N_31203);
nor U32527 (N_32527,N_31972,N_31234);
xnor U32528 (N_32528,N_31993,N_31525);
nand U32529 (N_32529,N_31975,N_31120);
or U32530 (N_32530,N_31192,N_31556);
and U32531 (N_32531,N_31780,N_31082);
nand U32532 (N_32532,N_31896,N_31215);
and U32533 (N_32533,N_31159,N_31968);
nand U32534 (N_32534,N_31850,N_31156);
nor U32535 (N_32535,N_31565,N_31273);
and U32536 (N_32536,N_31500,N_31579);
xnor U32537 (N_32537,N_31117,N_31729);
nand U32538 (N_32538,N_31139,N_31782);
or U32539 (N_32539,N_31805,N_31106);
nor U32540 (N_32540,N_31298,N_31562);
nand U32541 (N_32541,N_31845,N_31936);
or U32542 (N_32542,N_31003,N_31119);
nor U32543 (N_32543,N_31356,N_31277);
nor U32544 (N_32544,N_31993,N_31671);
and U32545 (N_32545,N_31985,N_31786);
nor U32546 (N_32546,N_31388,N_31567);
and U32547 (N_32547,N_31434,N_31236);
or U32548 (N_32548,N_31773,N_31394);
nand U32549 (N_32549,N_31737,N_31408);
nand U32550 (N_32550,N_31605,N_31907);
nand U32551 (N_32551,N_31026,N_31437);
or U32552 (N_32552,N_31686,N_31732);
xnor U32553 (N_32553,N_31829,N_31819);
nand U32554 (N_32554,N_31944,N_31101);
nor U32555 (N_32555,N_31881,N_31585);
xnor U32556 (N_32556,N_31661,N_31519);
or U32557 (N_32557,N_31279,N_31558);
nor U32558 (N_32558,N_31539,N_31091);
or U32559 (N_32559,N_31500,N_31513);
or U32560 (N_32560,N_31806,N_31669);
and U32561 (N_32561,N_31585,N_31995);
nand U32562 (N_32562,N_31169,N_31221);
xnor U32563 (N_32563,N_31613,N_31652);
nand U32564 (N_32564,N_31664,N_31879);
or U32565 (N_32565,N_31274,N_31863);
xnor U32566 (N_32566,N_31708,N_31553);
xor U32567 (N_32567,N_31872,N_31021);
or U32568 (N_32568,N_31568,N_31144);
nand U32569 (N_32569,N_31892,N_31158);
or U32570 (N_32570,N_31933,N_31240);
xnor U32571 (N_32571,N_31188,N_31209);
nor U32572 (N_32572,N_31494,N_31859);
xor U32573 (N_32573,N_31455,N_31838);
nand U32574 (N_32574,N_31920,N_31218);
nand U32575 (N_32575,N_31586,N_31456);
or U32576 (N_32576,N_31607,N_31640);
or U32577 (N_32577,N_31993,N_31849);
xnor U32578 (N_32578,N_31441,N_31933);
or U32579 (N_32579,N_31886,N_31105);
nand U32580 (N_32580,N_31324,N_31564);
nor U32581 (N_32581,N_31558,N_31990);
nor U32582 (N_32582,N_31434,N_31332);
nand U32583 (N_32583,N_31138,N_31239);
nand U32584 (N_32584,N_31912,N_31347);
xor U32585 (N_32585,N_31340,N_31394);
or U32586 (N_32586,N_31366,N_31612);
or U32587 (N_32587,N_31109,N_31195);
and U32588 (N_32588,N_31594,N_31717);
xor U32589 (N_32589,N_31518,N_31525);
xor U32590 (N_32590,N_31504,N_31772);
nand U32591 (N_32591,N_31102,N_31256);
or U32592 (N_32592,N_31730,N_31180);
or U32593 (N_32593,N_31838,N_31444);
or U32594 (N_32594,N_31573,N_31138);
xnor U32595 (N_32595,N_31717,N_31535);
nand U32596 (N_32596,N_31175,N_31542);
and U32597 (N_32597,N_31027,N_31525);
or U32598 (N_32598,N_31200,N_31022);
and U32599 (N_32599,N_31198,N_31309);
or U32600 (N_32600,N_31517,N_31364);
or U32601 (N_32601,N_31378,N_31181);
or U32602 (N_32602,N_31737,N_31420);
nor U32603 (N_32603,N_31255,N_31214);
and U32604 (N_32604,N_31191,N_31710);
or U32605 (N_32605,N_31047,N_31677);
or U32606 (N_32606,N_31985,N_31714);
xnor U32607 (N_32607,N_31072,N_31297);
and U32608 (N_32608,N_31359,N_31776);
nand U32609 (N_32609,N_31702,N_31580);
nand U32610 (N_32610,N_31992,N_31383);
nand U32611 (N_32611,N_31621,N_31009);
xor U32612 (N_32612,N_31653,N_31454);
and U32613 (N_32613,N_31253,N_31295);
or U32614 (N_32614,N_31572,N_31855);
and U32615 (N_32615,N_31607,N_31845);
nand U32616 (N_32616,N_31070,N_31580);
or U32617 (N_32617,N_31342,N_31021);
and U32618 (N_32618,N_31223,N_31106);
or U32619 (N_32619,N_31423,N_31631);
and U32620 (N_32620,N_31180,N_31382);
and U32621 (N_32621,N_31405,N_31073);
nor U32622 (N_32622,N_31608,N_31812);
nor U32623 (N_32623,N_31488,N_31889);
xnor U32624 (N_32624,N_31385,N_31276);
or U32625 (N_32625,N_31939,N_31448);
nand U32626 (N_32626,N_31447,N_31109);
and U32627 (N_32627,N_31121,N_31068);
nand U32628 (N_32628,N_31722,N_31517);
xnor U32629 (N_32629,N_31843,N_31272);
and U32630 (N_32630,N_31075,N_31340);
xor U32631 (N_32631,N_31293,N_31959);
and U32632 (N_32632,N_31005,N_31755);
nand U32633 (N_32633,N_31015,N_31363);
nor U32634 (N_32634,N_31412,N_31841);
xnor U32635 (N_32635,N_31994,N_31303);
nand U32636 (N_32636,N_31575,N_31477);
xnor U32637 (N_32637,N_31586,N_31241);
nand U32638 (N_32638,N_31727,N_31231);
or U32639 (N_32639,N_31364,N_31024);
xnor U32640 (N_32640,N_31201,N_31480);
or U32641 (N_32641,N_31362,N_31461);
xnor U32642 (N_32642,N_31355,N_31285);
nor U32643 (N_32643,N_31235,N_31237);
nor U32644 (N_32644,N_31141,N_31158);
xor U32645 (N_32645,N_31686,N_31198);
and U32646 (N_32646,N_31757,N_31956);
or U32647 (N_32647,N_31583,N_31414);
xor U32648 (N_32648,N_31046,N_31718);
and U32649 (N_32649,N_31591,N_31825);
nor U32650 (N_32650,N_31362,N_31249);
nand U32651 (N_32651,N_31540,N_31628);
nand U32652 (N_32652,N_31428,N_31796);
xor U32653 (N_32653,N_31580,N_31337);
and U32654 (N_32654,N_31378,N_31529);
and U32655 (N_32655,N_31921,N_31039);
nand U32656 (N_32656,N_31623,N_31020);
xnor U32657 (N_32657,N_31128,N_31434);
nand U32658 (N_32658,N_31593,N_31505);
and U32659 (N_32659,N_31321,N_31995);
nand U32660 (N_32660,N_31610,N_31742);
nand U32661 (N_32661,N_31222,N_31437);
nand U32662 (N_32662,N_31648,N_31841);
nand U32663 (N_32663,N_31205,N_31725);
or U32664 (N_32664,N_31646,N_31957);
nor U32665 (N_32665,N_31636,N_31665);
nor U32666 (N_32666,N_31210,N_31457);
nor U32667 (N_32667,N_31017,N_31587);
nand U32668 (N_32668,N_31430,N_31259);
nand U32669 (N_32669,N_31971,N_31359);
or U32670 (N_32670,N_31470,N_31799);
and U32671 (N_32671,N_31806,N_31486);
nor U32672 (N_32672,N_31726,N_31384);
and U32673 (N_32673,N_31921,N_31326);
nor U32674 (N_32674,N_31057,N_31377);
nand U32675 (N_32675,N_31060,N_31762);
nand U32676 (N_32676,N_31830,N_31652);
and U32677 (N_32677,N_31112,N_31822);
nand U32678 (N_32678,N_31455,N_31751);
or U32679 (N_32679,N_31136,N_31594);
nor U32680 (N_32680,N_31371,N_31525);
nand U32681 (N_32681,N_31061,N_31781);
nor U32682 (N_32682,N_31325,N_31115);
nand U32683 (N_32683,N_31888,N_31646);
and U32684 (N_32684,N_31240,N_31859);
or U32685 (N_32685,N_31292,N_31327);
xnor U32686 (N_32686,N_31138,N_31897);
nor U32687 (N_32687,N_31502,N_31116);
or U32688 (N_32688,N_31797,N_31290);
xor U32689 (N_32689,N_31305,N_31155);
or U32690 (N_32690,N_31761,N_31736);
nor U32691 (N_32691,N_31116,N_31820);
and U32692 (N_32692,N_31197,N_31154);
or U32693 (N_32693,N_31728,N_31794);
xnor U32694 (N_32694,N_31846,N_31251);
or U32695 (N_32695,N_31368,N_31692);
nand U32696 (N_32696,N_31378,N_31749);
or U32697 (N_32697,N_31096,N_31582);
nand U32698 (N_32698,N_31106,N_31005);
xor U32699 (N_32699,N_31522,N_31912);
and U32700 (N_32700,N_31123,N_31976);
nor U32701 (N_32701,N_31168,N_31578);
nor U32702 (N_32702,N_31200,N_31705);
xnor U32703 (N_32703,N_31642,N_31737);
xor U32704 (N_32704,N_31184,N_31535);
and U32705 (N_32705,N_31012,N_31078);
xnor U32706 (N_32706,N_31806,N_31513);
or U32707 (N_32707,N_31365,N_31201);
or U32708 (N_32708,N_31713,N_31814);
nor U32709 (N_32709,N_31836,N_31999);
nor U32710 (N_32710,N_31222,N_31640);
xnor U32711 (N_32711,N_31556,N_31749);
xor U32712 (N_32712,N_31757,N_31827);
and U32713 (N_32713,N_31452,N_31146);
nand U32714 (N_32714,N_31039,N_31629);
or U32715 (N_32715,N_31214,N_31922);
or U32716 (N_32716,N_31690,N_31736);
nand U32717 (N_32717,N_31870,N_31996);
or U32718 (N_32718,N_31522,N_31610);
and U32719 (N_32719,N_31928,N_31400);
xnor U32720 (N_32720,N_31474,N_31332);
nor U32721 (N_32721,N_31036,N_31105);
nor U32722 (N_32722,N_31430,N_31432);
xnor U32723 (N_32723,N_31067,N_31454);
or U32724 (N_32724,N_31299,N_31050);
and U32725 (N_32725,N_31789,N_31146);
or U32726 (N_32726,N_31009,N_31877);
and U32727 (N_32727,N_31455,N_31854);
or U32728 (N_32728,N_31814,N_31909);
or U32729 (N_32729,N_31555,N_31329);
and U32730 (N_32730,N_31486,N_31978);
or U32731 (N_32731,N_31723,N_31843);
xnor U32732 (N_32732,N_31623,N_31932);
or U32733 (N_32733,N_31424,N_31388);
nor U32734 (N_32734,N_31064,N_31455);
nand U32735 (N_32735,N_31122,N_31865);
nand U32736 (N_32736,N_31415,N_31338);
nand U32737 (N_32737,N_31448,N_31482);
or U32738 (N_32738,N_31609,N_31368);
or U32739 (N_32739,N_31334,N_31860);
nand U32740 (N_32740,N_31055,N_31435);
nand U32741 (N_32741,N_31196,N_31944);
nor U32742 (N_32742,N_31259,N_31894);
or U32743 (N_32743,N_31475,N_31016);
nor U32744 (N_32744,N_31301,N_31677);
and U32745 (N_32745,N_31713,N_31673);
or U32746 (N_32746,N_31857,N_31704);
or U32747 (N_32747,N_31327,N_31386);
nor U32748 (N_32748,N_31748,N_31187);
nor U32749 (N_32749,N_31674,N_31833);
and U32750 (N_32750,N_31974,N_31515);
nor U32751 (N_32751,N_31174,N_31760);
xnor U32752 (N_32752,N_31591,N_31745);
or U32753 (N_32753,N_31015,N_31539);
nand U32754 (N_32754,N_31491,N_31995);
xnor U32755 (N_32755,N_31209,N_31625);
and U32756 (N_32756,N_31574,N_31244);
xor U32757 (N_32757,N_31215,N_31156);
or U32758 (N_32758,N_31500,N_31053);
xor U32759 (N_32759,N_31625,N_31487);
or U32760 (N_32760,N_31162,N_31180);
nor U32761 (N_32761,N_31381,N_31992);
xor U32762 (N_32762,N_31471,N_31692);
nor U32763 (N_32763,N_31798,N_31342);
nand U32764 (N_32764,N_31312,N_31710);
or U32765 (N_32765,N_31997,N_31972);
nor U32766 (N_32766,N_31535,N_31864);
nand U32767 (N_32767,N_31572,N_31453);
nand U32768 (N_32768,N_31768,N_31128);
and U32769 (N_32769,N_31057,N_31101);
and U32770 (N_32770,N_31284,N_31588);
nand U32771 (N_32771,N_31207,N_31686);
and U32772 (N_32772,N_31143,N_31912);
and U32773 (N_32773,N_31103,N_31974);
and U32774 (N_32774,N_31987,N_31258);
xnor U32775 (N_32775,N_31694,N_31803);
nor U32776 (N_32776,N_31176,N_31143);
xor U32777 (N_32777,N_31872,N_31768);
nor U32778 (N_32778,N_31204,N_31167);
and U32779 (N_32779,N_31536,N_31357);
nor U32780 (N_32780,N_31145,N_31669);
nand U32781 (N_32781,N_31207,N_31809);
nand U32782 (N_32782,N_31591,N_31421);
nand U32783 (N_32783,N_31699,N_31546);
xor U32784 (N_32784,N_31495,N_31730);
xnor U32785 (N_32785,N_31920,N_31159);
nor U32786 (N_32786,N_31049,N_31038);
nand U32787 (N_32787,N_31970,N_31610);
xor U32788 (N_32788,N_31239,N_31602);
nor U32789 (N_32789,N_31384,N_31342);
and U32790 (N_32790,N_31170,N_31913);
nand U32791 (N_32791,N_31871,N_31029);
xor U32792 (N_32792,N_31092,N_31839);
or U32793 (N_32793,N_31319,N_31189);
xnor U32794 (N_32794,N_31789,N_31865);
or U32795 (N_32795,N_31676,N_31744);
nand U32796 (N_32796,N_31418,N_31094);
xnor U32797 (N_32797,N_31625,N_31899);
nor U32798 (N_32798,N_31251,N_31028);
and U32799 (N_32799,N_31499,N_31102);
xnor U32800 (N_32800,N_31941,N_31714);
xor U32801 (N_32801,N_31135,N_31304);
xnor U32802 (N_32802,N_31431,N_31656);
xor U32803 (N_32803,N_31606,N_31984);
or U32804 (N_32804,N_31643,N_31433);
and U32805 (N_32805,N_31466,N_31242);
nand U32806 (N_32806,N_31847,N_31308);
and U32807 (N_32807,N_31957,N_31210);
nor U32808 (N_32808,N_31337,N_31190);
nor U32809 (N_32809,N_31490,N_31205);
and U32810 (N_32810,N_31776,N_31136);
or U32811 (N_32811,N_31463,N_31461);
or U32812 (N_32812,N_31578,N_31744);
or U32813 (N_32813,N_31894,N_31252);
or U32814 (N_32814,N_31000,N_31211);
or U32815 (N_32815,N_31295,N_31989);
nor U32816 (N_32816,N_31056,N_31376);
xor U32817 (N_32817,N_31152,N_31780);
or U32818 (N_32818,N_31269,N_31288);
xor U32819 (N_32819,N_31866,N_31377);
and U32820 (N_32820,N_31408,N_31495);
nor U32821 (N_32821,N_31556,N_31429);
nor U32822 (N_32822,N_31812,N_31486);
xnor U32823 (N_32823,N_31723,N_31555);
nand U32824 (N_32824,N_31709,N_31380);
nor U32825 (N_32825,N_31682,N_31147);
and U32826 (N_32826,N_31358,N_31853);
xnor U32827 (N_32827,N_31729,N_31603);
xor U32828 (N_32828,N_31375,N_31712);
and U32829 (N_32829,N_31953,N_31036);
nor U32830 (N_32830,N_31679,N_31759);
nor U32831 (N_32831,N_31483,N_31606);
and U32832 (N_32832,N_31885,N_31132);
nor U32833 (N_32833,N_31481,N_31628);
nor U32834 (N_32834,N_31234,N_31308);
xnor U32835 (N_32835,N_31240,N_31522);
nor U32836 (N_32836,N_31593,N_31809);
nand U32837 (N_32837,N_31672,N_31966);
or U32838 (N_32838,N_31956,N_31628);
or U32839 (N_32839,N_31711,N_31886);
nand U32840 (N_32840,N_31047,N_31282);
nand U32841 (N_32841,N_31383,N_31429);
and U32842 (N_32842,N_31732,N_31593);
nor U32843 (N_32843,N_31842,N_31472);
nor U32844 (N_32844,N_31132,N_31932);
nor U32845 (N_32845,N_31127,N_31239);
or U32846 (N_32846,N_31546,N_31121);
xnor U32847 (N_32847,N_31998,N_31849);
nor U32848 (N_32848,N_31782,N_31286);
nor U32849 (N_32849,N_31984,N_31110);
nor U32850 (N_32850,N_31383,N_31036);
nand U32851 (N_32851,N_31701,N_31971);
and U32852 (N_32852,N_31967,N_31847);
or U32853 (N_32853,N_31376,N_31134);
and U32854 (N_32854,N_31067,N_31493);
and U32855 (N_32855,N_31206,N_31552);
or U32856 (N_32856,N_31229,N_31458);
or U32857 (N_32857,N_31953,N_31917);
or U32858 (N_32858,N_31638,N_31787);
or U32859 (N_32859,N_31585,N_31556);
nand U32860 (N_32860,N_31603,N_31559);
nand U32861 (N_32861,N_31373,N_31400);
or U32862 (N_32862,N_31716,N_31573);
nand U32863 (N_32863,N_31411,N_31789);
nand U32864 (N_32864,N_31093,N_31668);
nor U32865 (N_32865,N_31173,N_31070);
and U32866 (N_32866,N_31095,N_31453);
and U32867 (N_32867,N_31365,N_31140);
nor U32868 (N_32868,N_31177,N_31397);
xor U32869 (N_32869,N_31112,N_31607);
nor U32870 (N_32870,N_31447,N_31538);
and U32871 (N_32871,N_31577,N_31538);
xnor U32872 (N_32872,N_31303,N_31862);
nand U32873 (N_32873,N_31417,N_31732);
nand U32874 (N_32874,N_31375,N_31810);
xnor U32875 (N_32875,N_31152,N_31513);
and U32876 (N_32876,N_31109,N_31057);
xor U32877 (N_32877,N_31948,N_31344);
or U32878 (N_32878,N_31302,N_31135);
and U32879 (N_32879,N_31340,N_31993);
xor U32880 (N_32880,N_31208,N_31240);
nor U32881 (N_32881,N_31210,N_31415);
xnor U32882 (N_32882,N_31987,N_31921);
nor U32883 (N_32883,N_31535,N_31964);
nand U32884 (N_32884,N_31645,N_31900);
xor U32885 (N_32885,N_31548,N_31576);
and U32886 (N_32886,N_31447,N_31194);
nand U32887 (N_32887,N_31280,N_31361);
and U32888 (N_32888,N_31034,N_31747);
xnor U32889 (N_32889,N_31219,N_31232);
or U32890 (N_32890,N_31601,N_31139);
nor U32891 (N_32891,N_31770,N_31553);
xor U32892 (N_32892,N_31895,N_31291);
and U32893 (N_32893,N_31485,N_31851);
or U32894 (N_32894,N_31459,N_31423);
or U32895 (N_32895,N_31650,N_31986);
and U32896 (N_32896,N_31292,N_31049);
and U32897 (N_32897,N_31959,N_31137);
nand U32898 (N_32898,N_31054,N_31089);
xor U32899 (N_32899,N_31948,N_31159);
and U32900 (N_32900,N_31333,N_31596);
xnor U32901 (N_32901,N_31643,N_31731);
nand U32902 (N_32902,N_31795,N_31616);
nor U32903 (N_32903,N_31458,N_31326);
xor U32904 (N_32904,N_31263,N_31062);
nor U32905 (N_32905,N_31091,N_31102);
nor U32906 (N_32906,N_31863,N_31100);
and U32907 (N_32907,N_31013,N_31882);
xor U32908 (N_32908,N_31530,N_31506);
or U32909 (N_32909,N_31695,N_31921);
or U32910 (N_32910,N_31818,N_31556);
and U32911 (N_32911,N_31066,N_31366);
or U32912 (N_32912,N_31773,N_31641);
nand U32913 (N_32913,N_31795,N_31258);
xnor U32914 (N_32914,N_31287,N_31311);
xnor U32915 (N_32915,N_31849,N_31940);
nor U32916 (N_32916,N_31869,N_31690);
nand U32917 (N_32917,N_31746,N_31967);
nor U32918 (N_32918,N_31978,N_31208);
and U32919 (N_32919,N_31202,N_31701);
nor U32920 (N_32920,N_31875,N_31055);
nor U32921 (N_32921,N_31418,N_31251);
or U32922 (N_32922,N_31977,N_31187);
nor U32923 (N_32923,N_31426,N_31769);
nand U32924 (N_32924,N_31465,N_31410);
or U32925 (N_32925,N_31766,N_31285);
or U32926 (N_32926,N_31673,N_31848);
or U32927 (N_32927,N_31813,N_31615);
nor U32928 (N_32928,N_31714,N_31733);
nand U32929 (N_32929,N_31748,N_31614);
nand U32930 (N_32930,N_31931,N_31086);
nor U32931 (N_32931,N_31073,N_31481);
xnor U32932 (N_32932,N_31247,N_31060);
nor U32933 (N_32933,N_31599,N_31789);
nor U32934 (N_32934,N_31574,N_31426);
or U32935 (N_32935,N_31150,N_31517);
xor U32936 (N_32936,N_31794,N_31795);
nor U32937 (N_32937,N_31560,N_31202);
or U32938 (N_32938,N_31258,N_31966);
or U32939 (N_32939,N_31593,N_31839);
or U32940 (N_32940,N_31552,N_31276);
and U32941 (N_32941,N_31778,N_31595);
xor U32942 (N_32942,N_31085,N_31196);
nor U32943 (N_32943,N_31872,N_31617);
nand U32944 (N_32944,N_31238,N_31952);
and U32945 (N_32945,N_31764,N_31997);
or U32946 (N_32946,N_31549,N_31061);
nor U32947 (N_32947,N_31419,N_31465);
nor U32948 (N_32948,N_31292,N_31607);
xnor U32949 (N_32949,N_31764,N_31377);
or U32950 (N_32950,N_31397,N_31303);
xor U32951 (N_32951,N_31594,N_31304);
and U32952 (N_32952,N_31900,N_31094);
nand U32953 (N_32953,N_31589,N_31801);
and U32954 (N_32954,N_31168,N_31685);
nand U32955 (N_32955,N_31114,N_31040);
and U32956 (N_32956,N_31624,N_31271);
xor U32957 (N_32957,N_31970,N_31574);
nand U32958 (N_32958,N_31925,N_31476);
nand U32959 (N_32959,N_31895,N_31165);
nor U32960 (N_32960,N_31884,N_31922);
and U32961 (N_32961,N_31703,N_31420);
nand U32962 (N_32962,N_31866,N_31107);
nand U32963 (N_32963,N_31411,N_31375);
nand U32964 (N_32964,N_31375,N_31899);
xor U32965 (N_32965,N_31435,N_31550);
nand U32966 (N_32966,N_31554,N_31078);
nor U32967 (N_32967,N_31454,N_31613);
nand U32968 (N_32968,N_31505,N_31644);
or U32969 (N_32969,N_31227,N_31348);
and U32970 (N_32970,N_31162,N_31338);
nor U32971 (N_32971,N_31262,N_31441);
or U32972 (N_32972,N_31513,N_31548);
nor U32973 (N_32973,N_31321,N_31387);
or U32974 (N_32974,N_31857,N_31545);
and U32975 (N_32975,N_31019,N_31497);
nor U32976 (N_32976,N_31769,N_31692);
or U32977 (N_32977,N_31808,N_31988);
nor U32978 (N_32978,N_31773,N_31823);
xnor U32979 (N_32979,N_31710,N_31892);
or U32980 (N_32980,N_31339,N_31761);
nor U32981 (N_32981,N_31673,N_31631);
or U32982 (N_32982,N_31020,N_31734);
nor U32983 (N_32983,N_31771,N_31524);
xnor U32984 (N_32984,N_31186,N_31479);
or U32985 (N_32985,N_31081,N_31955);
nor U32986 (N_32986,N_31100,N_31987);
and U32987 (N_32987,N_31534,N_31934);
nor U32988 (N_32988,N_31014,N_31049);
and U32989 (N_32989,N_31780,N_31143);
or U32990 (N_32990,N_31790,N_31966);
nand U32991 (N_32991,N_31346,N_31928);
nand U32992 (N_32992,N_31848,N_31155);
and U32993 (N_32993,N_31092,N_31360);
or U32994 (N_32994,N_31102,N_31308);
or U32995 (N_32995,N_31390,N_31577);
and U32996 (N_32996,N_31629,N_31941);
or U32997 (N_32997,N_31878,N_31066);
xor U32998 (N_32998,N_31418,N_31002);
xor U32999 (N_32999,N_31421,N_31704);
or U33000 (N_33000,N_32682,N_32257);
nor U33001 (N_33001,N_32600,N_32037);
xnor U33002 (N_33002,N_32282,N_32482);
or U33003 (N_33003,N_32982,N_32613);
nand U33004 (N_33004,N_32462,N_32896);
nor U33005 (N_33005,N_32805,N_32430);
or U33006 (N_33006,N_32380,N_32798);
xor U33007 (N_33007,N_32581,N_32622);
xor U33008 (N_33008,N_32845,N_32969);
and U33009 (N_33009,N_32855,N_32728);
xor U33010 (N_33010,N_32510,N_32789);
nor U33011 (N_33011,N_32822,N_32379);
xor U33012 (N_33012,N_32154,N_32685);
xor U33013 (N_33013,N_32064,N_32126);
nand U33014 (N_33014,N_32409,N_32275);
nor U33015 (N_33015,N_32347,N_32865);
and U33016 (N_33016,N_32874,N_32922);
nor U33017 (N_33017,N_32860,N_32988);
nand U33018 (N_33018,N_32694,N_32315);
nand U33019 (N_33019,N_32444,N_32422);
nor U33020 (N_33020,N_32359,N_32455);
or U33021 (N_33021,N_32343,N_32313);
or U33022 (N_33022,N_32308,N_32425);
nand U33023 (N_33023,N_32353,N_32757);
and U33024 (N_33024,N_32345,N_32421);
xor U33025 (N_33025,N_32958,N_32610);
or U33026 (N_33026,N_32442,N_32990);
or U33027 (N_33027,N_32594,N_32941);
xor U33028 (N_33028,N_32734,N_32013);
nor U33029 (N_33029,N_32429,N_32036);
nor U33030 (N_33030,N_32180,N_32292);
xor U33031 (N_33031,N_32243,N_32493);
or U33032 (N_33032,N_32206,N_32119);
xor U33033 (N_33033,N_32265,N_32711);
xnor U33034 (N_33034,N_32813,N_32652);
and U33035 (N_33035,N_32057,N_32793);
xnor U33036 (N_33036,N_32673,N_32733);
and U33037 (N_33037,N_32800,N_32151);
or U33038 (N_33038,N_32513,N_32745);
xnor U33039 (N_33039,N_32964,N_32207);
and U33040 (N_33040,N_32973,N_32818);
or U33041 (N_33041,N_32386,N_32007);
nand U33042 (N_33042,N_32410,N_32008);
xnor U33043 (N_33043,N_32894,N_32092);
xor U33044 (N_33044,N_32428,N_32318);
and U33045 (N_33045,N_32411,N_32754);
or U33046 (N_33046,N_32231,N_32103);
and U33047 (N_33047,N_32340,N_32851);
and U33048 (N_33048,N_32893,N_32784);
nand U33049 (N_33049,N_32344,N_32885);
xnor U33050 (N_33050,N_32210,N_32978);
or U33051 (N_33051,N_32397,N_32545);
and U33052 (N_33052,N_32110,N_32461);
xnor U33053 (N_33053,N_32290,N_32396);
xnor U33054 (N_33054,N_32662,N_32432);
or U33055 (N_33055,N_32497,N_32371);
or U33056 (N_33056,N_32656,N_32624);
nand U33057 (N_33057,N_32633,N_32938);
or U33058 (N_33058,N_32394,N_32378);
nand U33059 (N_33059,N_32216,N_32528);
nor U33060 (N_33060,N_32141,N_32358);
xnor U33061 (N_33061,N_32055,N_32459);
xnor U33062 (N_33062,N_32752,N_32582);
nor U33063 (N_33063,N_32628,N_32066);
nor U33064 (N_33064,N_32399,N_32102);
nor U33065 (N_33065,N_32959,N_32834);
nand U33066 (N_33066,N_32569,N_32059);
nand U33067 (N_33067,N_32242,N_32289);
or U33068 (N_33068,N_32160,N_32142);
and U33069 (N_33069,N_32693,N_32599);
nand U33070 (N_33070,N_32952,N_32564);
nand U33071 (N_33071,N_32079,N_32786);
and U33072 (N_33072,N_32568,N_32288);
nor U33073 (N_33073,N_32269,N_32226);
nand U33074 (N_33074,N_32134,N_32362);
nand U33075 (N_33075,N_32520,N_32718);
or U33076 (N_33076,N_32476,N_32846);
xor U33077 (N_33077,N_32947,N_32112);
and U33078 (N_33078,N_32256,N_32299);
or U33079 (N_33079,N_32273,N_32368);
nor U33080 (N_33080,N_32720,N_32355);
nor U33081 (N_33081,N_32283,N_32566);
and U33082 (N_33082,N_32487,N_32584);
and U33083 (N_33083,N_32829,N_32635);
nor U33084 (N_33084,N_32611,N_32413);
and U33085 (N_33085,N_32872,N_32172);
or U33086 (N_33086,N_32350,N_32850);
nand U33087 (N_33087,N_32255,N_32637);
xnor U33088 (N_33088,N_32148,N_32418);
or U33089 (N_33089,N_32161,N_32506);
xor U33090 (N_33090,N_32909,N_32911);
and U33091 (N_33091,N_32515,N_32705);
nand U33092 (N_33092,N_32987,N_32348);
nor U33093 (N_33093,N_32446,N_32687);
and U33094 (N_33094,N_32565,N_32262);
or U33095 (N_33095,N_32251,N_32310);
xor U33096 (N_33096,N_32441,N_32073);
nand U33097 (N_33097,N_32069,N_32304);
and U33098 (N_33098,N_32127,N_32541);
xor U33099 (N_33099,N_32556,N_32090);
nand U33100 (N_33100,N_32732,N_32025);
nand U33101 (N_33101,N_32848,N_32701);
xor U33102 (N_33102,N_32181,N_32484);
or U33103 (N_33103,N_32391,N_32116);
xor U33104 (N_33104,N_32641,N_32495);
and U33105 (N_33105,N_32676,N_32217);
and U33106 (N_33106,N_32063,N_32955);
or U33107 (N_33107,N_32691,N_32963);
or U33108 (N_33108,N_32144,N_32370);
xnor U33109 (N_33109,N_32198,N_32212);
xor U33110 (N_33110,N_32724,N_32551);
or U33111 (N_33111,N_32264,N_32174);
nor U33112 (N_33112,N_32284,N_32535);
and U33113 (N_33113,N_32744,N_32143);
nand U33114 (N_33114,N_32714,N_32605);
nor U33115 (N_33115,N_32097,N_32763);
nand U33116 (N_33116,N_32638,N_32260);
xnor U33117 (N_33117,N_32113,N_32925);
xnor U33118 (N_33118,N_32547,N_32145);
and U33119 (N_33119,N_32155,N_32906);
or U33120 (N_33120,N_32042,N_32327);
and U33121 (N_33121,N_32808,N_32287);
and U33122 (N_33122,N_32470,N_32883);
nand U33123 (N_33123,N_32305,N_32105);
or U33124 (N_33124,N_32590,N_32050);
and U33125 (N_33125,N_32919,N_32831);
xor U33126 (N_33126,N_32956,N_32523);
or U33127 (N_33127,N_32940,N_32494);
and U33128 (N_33128,N_32248,N_32787);
and U33129 (N_33129,N_32489,N_32930);
nand U33130 (N_33130,N_32467,N_32749);
and U33131 (N_33131,N_32222,N_32406);
and U33132 (N_33132,N_32514,N_32086);
and U33133 (N_33133,N_32190,N_32375);
and U33134 (N_33134,N_32076,N_32196);
nor U33135 (N_33135,N_32768,N_32980);
nor U33136 (N_33136,N_32835,N_32507);
xnor U33137 (N_33137,N_32946,N_32435);
and U33138 (N_33138,N_32202,N_32286);
and U33139 (N_33139,N_32096,N_32616);
and U33140 (N_33140,N_32658,N_32739);
xor U33141 (N_33141,N_32115,N_32508);
nor U33142 (N_33142,N_32456,N_32093);
nor U33143 (N_33143,N_32049,N_32901);
nand U33144 (N_33144,N_32867,N_32424);
or U33145 (N_33145,N_32204,N_32402);
xor U33146 (N_33146,N_32769,N_32843);
nor U33147 (N_33147,N_32607,N_32542);
nor U33148 (N_33148,N_32663,N_32957);
or U33149 (N_33149,N_32838,N_32225);
or U33150 (N_33150,N_32385,N_32316);
nor U33151 (N_33151,N_32774,N_32821);
and U33152 (N_33152,N_32166,N_32747);
nor U33153 (N_33153,N_32229,N_32077);
or U33154 (N_33154,N_32029,N_32966);
nand U33155 (N_33155,N_32197,N_32892);
nor U33156 (N_33156,N_32950,N_32218);
xnor U33157 (N_33157,N_32490,N_32211);
nand U33158 (N_33158,N_32132,N_32052);
nand U33159 (N_33159,N_32992,N_32870);
or U33160 (N_33160,N_32912,N_32072);
and U33161 (N_33161,N_32554,N_32647);
or U33162 (N_33162,N_32239,N_32876);
xor U33163 (N_33163,N_32176,N_32241);
nor U33164 (N_33164,N_32031,N_32719);
nor U33165 (N_33165,N_32071,N_32777);
nor U33166 (N_33166,N_32708,N_32018);
or U33167 (N_33167,N_32233,N_32440);
and U33168 (N_33168,N_32125,N_32017);
nand U33169 (N_33169,N_32644,N_32136);
nand U33170 (N_33170,N_32479,N_32108);
nor U33171 (N_33171,N_32918,N_32496);
and U33172 (N_33172,N_32035,N_32875);
or U33173 (N_33173,N_32447,N_32192);
nor U33174 (N_33174,N_32175,N_32758);
xor U33175 (N_33175,N_32346,N_32903);
nand U33176 (N_33176,N_32157,N_32780);
nor U33177 (N_33177,N_32329,N_32153);
or U33178 (N_33178,N_32033,N_32139);
or U33179 (N_33179,N_32001,N_32801);
xnor U33180 (N_33180,N_32942,N_32555);
and U33181 (N_33181,N_32034,N_32664);
xor U33182 (N_33182,N_32756,N_32924);
xor U33183 (N_33183,N_32184,N_32640);
nor U33184 (N_33184,N_32254,N_32453);
nand U33185 (N_33185,N_32856,N_32056);
nor U33186 (N_33186,N_32936,N_32655);
xor U33187 (N_33187,N_32471,N_32372);
or U33188 (N_33188,N_32404,N_32140);
nor U33189 (N_33189,N_32913,N_32138);
and U33190 (N_33190,N_32983,N_32237);
xor U33191 (N_33191,N_32677,N_32303);
xor U33192 (N_33192,N_32560,N_32107);
or U33193 (N_33193,N_32989,N_32081);
nor U33194 (N_33194,N_32578,N_32833);
nand U33195 (N_33195,N_32252,N_32729);
or U33196 (N_33196,N_32999,N_32962);
or U33197 (N_33197,N_32579,N_32311);
or U33198 (N_33198,N_32213,N_32381);
or U33199 (N_33199,N_32512,N_32377);
and U33200 (N_33200,N_32690,N_32232);
nand U33201 (N_33201,N_32058,N_32791);
and U33202 (N_33202,N_32109,N_32890);
xnor U33203 (N_33203,N_32878,N_32889);
nor U33204 (N_33204,N_32934,N_32443);
nor U33205 (N_33205,N_32954,N_32880);
xor U33206 (N_33206,N_32117,N_32811);
nand U33207 (N_33207,N_32130,N_32356);
nor U33208 (N_33208,N_32367,N_32620);
xnor U33209 (N_33209,N_32186,N_32731);
nor U33210 (N_33210,N_32187,N_32928);
nand U33211 (N_33211,N_32464,N_32162);
or U33212 (N_33212,N_32245,N_32511);
xor U33213 (N_33213,N_32227,N_32672);
and U33214 (N_33214,N_32643,N_32006);
xnor U33215 (N_33215,N_32975,N_32539);
or U33216 (N_33216,N_32032,N_32009);
nor U33217 (N_33217,N_32738,N_32853);
xor U33218 (N_33218,N_32695,N_32585);
nor U33219 (N_33219,N_32707,N_32692);
nand U33220 (N_33220,N_32871,N_32965);
and U33221 (N_33221,N_32603,N_32448);
nand U33222 (N_33222,N_32261,N_32150);
nor U33223 (N_33223,N_32604,N_32984);
and U33224 (N_33224,N_32653,N_32706);
xor U33225 (N_33225,N_32067,N_32790);
and U33226 (N_33226,N_32334,N_32247);
or U33227 (N_33227,N_32812,N_32840);
nor U33228 (N_33228,N_32679,N_32098);
and U33229 (N_33229,N_32466,N_32700);
nand U33230 (N_33230,N_32949,N_32062);
xnor U33231 (N_33231,N_32991,N_32078);
and U33232 (N_33232,N_32179,N_32866);
nor U33233 (N_33233,N_32028,N_32328);
nor U33234 (N_33234,N_32163,N_32408);
xor U33235 (N_33235,N_32503,N_32048);
and U33236 (N_33236,N_32935,N_32819);
or U33237 (N_33237,N_32039,N_32760);
xnor U33238 (N_33238,N_32669,N_32689);
and U33239 (N_33239,N_32219,N_32713);
nor U33240 (N_33240,N_32319,N_32550);
nand U33241 (N_33241,N_32854,N_32671);
nand U33242 (N_33242,N_32426,N_32061);
or U33243 (N_33243,N_32549,N_32349);
or U33244 (N_33244,N_32236,N_32023);
nand U33245 (N_33245,N_32366,N_32333);
nand U33246 (N_33246,N_32369,N_32297);
or U33247 (N_33247,N_32960,N_32414);
and U33248 (N_33248,N_32400,N_32178);
nor U33249 (N_33249,N_32277,N_32193);
nor U33250 (N_33250,N_32214,N_32053);
and U33251 (N_33251,N_32398,N_32363);
nand U33252 (N_33252,N_32352,N_32735);
and U33253 (N_33253,N_32660,N_32882);
xor U33254 (N_33254,N_32606,N_32267);
nor U33255 (N_33255,N_32068,N_32223);
and U33256 (N_33256,N_32392,N_32419);
nand U33257 (N_33257,N_32612,N_32101);
nor U33258 (N_33258,N_32194,N_32026);
and U33259 (N_33259,N_32910,N_32712);
xnor U33260 (N_33260,N_32920,N_32552);
nand U33261 (N_33261,N_32976,N_32953);
and U33262 (N_33262,N_32085,N_32173);
or U33263 (N_33263,N_32575,N_32710);
nand U33264 (N_33264,N_32703,N_32626);
and U33265 (N_33265,N_32244,N_32208);
or U33266 (N_33266,N_32040,N_32771);
or U33267 (N_33267,N_32776,N_32985);
or U33268 (N_33268,N_32567,N_32937);
xor U33269 (N_33269,N_32841,N_32317);
nor U33270 (N_33270,N_32384,N_32617);
xor U33271 (N_33271,N_32452,N_32010);
or U33272 (N_33272,N_32128,N_32259);
and U33273 (N_33273,N_32773,N_32080);
nand U33274 (N_33274,N_32839,N_32051);
nor U33275 (N_33275,N_32230,N_32727);
or U33276 (N_33276,N_32544,N_32164);
xor U33277 (N_33277,N_32075,N_32133);
or U33278 (N_33278,N_32796,N_32281);
xnor U33279 (N_33279,N_32927,N_32608);
or U33280 (N_33280,N_32827,N_32401);
nand U33281 (N_33281,N_32804,N_32932);
nor U33282 (N_33282,N_32249,N_32521);
xor U33283 (N_33283,N_32580,N_32016);
or U33284 (N_33284,N_32864,N_32877);
and U33285 (N_33285,N_32169,N_32011);
and U33286 (N_33286,N_32388,N_32122);
nand U33287 (N_33287,N_32412,N_32041);
nand U33288 (N_33288,N_32881,N_32382);
xor U33289 (N_33289,N_32486,N_32004);
and U33290 (N_33290,N_32809,N_32478);
nor U33291 (N_33291,N_32824,N_32698);
and U33292 (N_33292,N_32374,N_32686);
xor U33293 (N_33293,N_32666,N_32759);
and U33294 (N_33294,N_32792,N_32751);
nand U33295 (N_33295,N_32038,N_32814);
nand U33296 (N_33296,N_32383,N_32997);
and U33297 (N_33297,N_32129,N_32054);
and U33298 (N_33298,N_32439,N_32330);
or U33299 (N_33299,N_32895,N_32200);
xor U33300 (N_33300,N_32312,N_32046);
or U33301 (N_33301,N_32639,N_32929);
and U33302 (N_33302,N_32525,N_32968);
xor U33303 (N_33303,N_32996,N_32088);
or U33304 (N_33304,N_32502,N_32403);
nor U33305 (N_33305,N_32314,N_32797);
nand U33306 (N_33306,N_32634,N_32407);
or U33307 (N_33307,N_32923,N_32291);
xor U33308 (N_33308,N_32124,N_32778);
nand U33309 (N_33309,N_32454,N_32994);
or U33310 (N_33310,N_32271,N_32817);
or U33311 (N_33311,N_32755,N_32389);
xor U33312 (N_33312,N_32948,N_32189);
or U33313 (N_33313,N_32279,N_32012);
and U33314 (N_33314,N_32268,N_32087);
xnor U33315 (N_33315,N_32301,N_32543);
xor U33316 (N_33316,N_32065,N_32737);
or U33317 (N_33317,N_32469,N_32837);
or U33318 (N_33318,N_32688,N_32320);
nor U33319 (N_33319,N_32898,N_32782);
nor U33320 (N_33320,N_32869,N_32240);
and U33321 (N_33321,N_32203,N_32030);
xor U33322 (N_33322,N_32699,N_32131);
nor U33323 (N_33323,N_32972,N_32785);
xor U33324 (N_33324,N_32250,N_32331);
nand U33325 (N_33325,N_32977,N_32858);
xnor U33326 (N_33326,N_32721,N_32530);
or U33327 (N_33327,N_32532,N_32593);
or U33328 (N_33328,N_32645,N_32517);
or U33329 (N_33329,N_32943,N_32651);
xor U33330 (N_33330,N_32583,N_32373);
or U33331 (N_33331,N_32609,N_32298);
and U33332 (N_33332,N_32205,N_32632);
nor U33333 (N_33333,N_32862,N_32003);
nand U33334 (N_33334,N_32123,N_32137);
nor U33335 (N_33335,N_32118,N_32019);
and U33336 (N_33336,N_32423,N_32657);
and U33337 (N_33337,N_32518,N_32696);
nand U33338 (N_33338,N_32188,N_32182);
nand U33339 (N_33339,N_32341,N_32816);
xor U33340 (N_33340,N_32601,N_32614);
or U33341 (N_33341,N_32723,N_32234);
nand U33342 (N_33342,N_32746,N_32631);
nor U33343 (N_33343,N_32149,N_32799);
nand U33344 (N_33344,N_32722,N_32084);
nand U33345 (N_33345,N_32027,N_32615);
nand U33346 (N_33346,N_32764,N_32522);
or U33347 (N_33347,N_32762,N_32309);
xor U33348 (N_33348,N_32165,N_32665);
nand U33349 (N_33349,N_32921,N_32852);
and U33350 (N_33350,N_32627,N_32725);
nor U33351 (N_33351,N_32621,N_32907);
or U33352 (N_33352,N_32884,N_32433);
nor U33353 (N_33353,N_32238,N_32646);
nand U33354 (N_33354,N_32888,N_32899);
nand U33355 (N_33355,N_32998,N_32158);
and U33356 (N_33356,N_32917,N_32020);
and U33357 (N_33357,N_32823,N_32415);
nor U33358 (N_33358,N_32451,N_32772);
xnor U33359 (N_33359,N_32357,N_32697);
and U33360 (N_33360,N_32104,N_32152);
or U33361 (N_33361,N_32887,N_32460);
nor U33362 (N_33362,N_32505,N_32595);
nor U33363 (N_33363,N_32168,N_32263);
and U33364 (N_33364,N_32726,N_32648);
nand U33365 (N_33365,N_32553,N_32806);
xor U33366 (N_33366,N_32434,N_32156);
or U33367 (N_33367,N_32570,N_32499);
nand U33368 (N_33368,N_32572,N_32736);
and U33369 (N_33369,N_32832,N_32465);
nand U33370 (N_33370,N_32364,N_32536);
nor U33371 (N_33371,N_32574,N_32859);
nand U33372 (N_33372,N_32043,N_32483);
or U33373 (N_33373,N_32857,N_32945);
or U33374 (N_33374,N_32961,N_32970);
nor U33375 (N_33375,N_32540,N_32005);
xor U33376 (N_33376,N_32681,N_32095);
and U33377 (N_33377,N_32235,N_32220);
nand U33378 (N_33378,N_32592,N_32060);
nand U33379 (N_33379,N_32390,N_32674);
xor U33380 (N_33380,N_32967,N_32675);
or U33381 (N_33381,N_32395,N_32477);
nand U33382 (N_33382,N_32070,N_32844);
or U33383 (N_33383,N_32559,N_32803);
and U33384 (N_33384,N_32596,N_32636);
or U33385 (N_33385,N_32417,N_32879);
or U33386 (N_33386,N_32278,N_32562);
nand U33387 (N_33387,N_32981,N_32002);
nand U33388 (N_33388,N_32828,N_32500);
nand U33389 (N_33389,N_32336,N_32258);
nor U33390 (N_33390,N_32836,N_32307);
nor U33391 (N_33391,N_32337,N_32668);
nand U33392 (N_33392,N_32683,N_32571);
xnor U33393 (N_33393,N_32767,N_32931);
or U33394 (N_33394,N_32427,N_32481);
nand U33395 (N_33395,N_32276,N_32170);
and U33396 (N_33396,N_32416,N_32509);
and U33397 (N_33397,N_32886,N_32159);
and U33398 (N_33398,N_32365,N_32015);
nor U33399 (N_33399,N_32993,N_32463);
nor U33400 (N_33400,N_32715,N_32387);
or U33401 (N_33401,N_32587,N_32891);
xnor U33402 (N_33402,N_32802,N_32360);
and U33403 (N_33403,N_32740,N_32472);
nor U33404 (N_33404,N_32121,N_32529);
and U33405 (N_33405,N_32215,N_32351);
xnor U33406 (N_33406,N_32504,N_32781);
xor U33407 (N_33407,N_32630,N_32557);
or U33408 (N_33408,N_32815,N_32642);
nand U33409 (N_33409,N_32944,N_32022);
and U33410 (N_33410,N_32742,N_32111);
or U33411 (N_33411,N_32100,N_32338);
xor U33412 (N_33412,N_32342,N_32702);
xnor U33413 (N_33413,N_32332,N_32974);
xnor U33414 (N_33414,N_32900,N_32868);
nor U33415 (N_33415,N_32563,N_32704);
xor U33416 (N_33416,N_32684,N_32516);
nor U33417 (N_33417,N_32221,N_32753);
or U33418 (N_33418,N_32519,N_32473);
or U33419 (N_33419,N_32717,N_32826);
and U33420 (N_33420,N_32306,N_32339);
nand U33421 (N_33421,N_32524,N_32475);
nor U33422 (N_33422,N_32591,N_32573);
or U33423 (N_33423,N_32625,N_32488);
or U33424 (N_33424,N_32485,N_32926);
nand U33425 (N_33425,N_32654,N_32376);
or U33426 (N_33426,N_32106,N_32830);
or U33427 (N_33427,N_32939,N_32171);
and U33428 (N_33428,N_32014,N_32561);
nor U33429 (N_33429,N_32548,N_32750);
nand U33430 (N_33430,N_32933,N_32266);
xor U33431 (N_33431,N_32094,N_32847);
nand U33432 (N_33432,N_32436,N_32321);
and U33433 (N_33433,N_32457,N_32272);
nor U33434 (N_33434,N_32576,N_32670);
and U33435 (N_33435,N_32849,N_32228);
or U33436 (N_33436,N_32597,N_32825);
and U33437 (N_33437,N_32649,N_32361);
and U33438 (N_33438,N_32979,N_32667);
nor U33439 (N_33439,N_32449,N_32294);
and U33440 (N_33440,N_32393,N_32765);
and U33441 (N_33441,N_32185,N_32322);
nand U33442 (N_33442,N_32420,N_32445);
and U33443 (N_33443,N_32325,N_32326);
or U33444 (N_33444,N_32114,N_32951);
xnor U33445 (N_33445,N_32783,N_32915);
and U33446 (N_33446,N_32533,N_32099);
or U33447 (N_33447,N_32024,N_32354);
nor U33448 (N_33448,N_32650,N_32191);
nor U33449 (N_33449,N_32761,N_32302);
nand U33450 (N_33450,N_32709,N_32904);
nand U33451 (N_33451,N_32468,N_32916);
nor U33452 (N_33452,N_32270,N_32253);
and U33453 (N_33453,N_32146,N_32498);
and U33454 (N_33454,N_32295,N_32558);
nor U33455 (N_33455,N_32450,N_32074);
xor U33456 (N_33456,N_32293,N_32986);
or U33457 (N_33457,N_32474,N_32788);
and U33458 (N_33458,N_32195,N_32795);
nor U33459 (N_33459,N_32598,N_32716);
nand U33460 (N_33460,N_32661,N_32438);
or U33461 (N_33461,N_32300,N_32209);
nand U33462 (N_33462,N_32602,N_32280);
nor U33463 (N_33463,N_32618,N_32770);
and U33464 (N_33464,N_32183,N_32246);
or U33465 (N_33465,N_32873,N_32995);
and U33466 (N_33466,N_32659,N_32861);
nand U33467 (N_33467,N_32678,N_32147);
nand U33468 (N_33468,N_32531,N_32274);
nor U33469 (N_33469,N_32082,N_32296);
xor U33470 (N_33470,N_32526,N_32807);
or U33471 (N_33471,N_32577,N_32748);
nor U33472 (N_33472,N_32091,N_32914);
xor U33473 (N_33473,N_32680,N_32021);
or U33474 (N_33474,N_32766,N_32089);
xor U33475 (N_33475,N_32629,N_32820);
and U33476 (N_33476,N_32405,N_32323);
nor U33477 (N_33477,N_32501,N_32458);
or U33478 (N_33478,N_32897,N_32971);
nor U33479 (N_33479,N_32083,N_32905);
xor U33480 (N_33480,N_32044,N_32537);
nor U33481 (N_33481,N_32902,N_32730);
nor U33482 (N_33482,N_32619,N_32588);
nor U33483 (N_33483,N_32779,N_32167);
and U33484 (N_33484,N_32045,N_32335);
nor U33485 (N_33485,N_32480,N_32538);
or U33486 (N_33486,N_32492,N_32491);
nand U33487 (N_33487,N_32743,N_32842);
nor U33488 (N_33488,N_32047,N_32177);
and U33489 (N_33489,N_32586,N_32810);
xor U33490 (N_33490,N_32135,N_32285);
or U33491 (N_33491,N_32863,N_32623);
nand U33492 (N_33492,N_32201,N_32120);
xor U33493 (N_33493,N_32199,N_32527);
nor U33494 (N_33494,N_32775,N_32534);
nor U33495 (N_33495,N_32908,N_32437);
and U33496 (N_33496,N_32546,N_32794);
and U33497 (N_33497,N_32431,N_32224);
nor U33498 (N_33498,N_32741,N_32324);
and U33499 (N_33499,N_32000,N_32589);
and U33500 (N_33500,N_32837,N_32334);
or U33501 (N_33501,N_32444,N_32869);
or U33502 (N_33502,N_32109,N_32805);
nand U33503 (N_33503,N_32096,N_32215);
nor U33504 (N_33504,N_32615,N_32443);
or U33505 (N_33505,N_32818,N_32102);
nand U33506 (N_33506,N_32816,N_32945);
nand U33507 (N_33507,N_32717,N_32355);
nor U33508 (N_33508,N_32546,N_32000);
nand U33509 (N_33509,N_32470,N_32162);
or U33510 (N_33510,N_32229,N_32924);
nand U33511 (N_33511,N_32958,N_32588);
xor U33512 (N_33512,N_32646,N_32728);
and U33513 (N_33513,N_32516,N_32360);
nor U33514 (N_33514,N_32724,N_32700);
and U33515 (N_33515,N_32105,N_32736);
nand U33516 (N_33516,N_32722,N_32716);
or U33517 (N_33517,N_32204,N_32431);
nor U33518 (N_33518,N_32893,N_32227);
and U33519 (N_33519,N_32953,N_32130);
or U33520 (N_33520,N_32123,N_32415);
or U33521 (N_33521,N_32317,N_32327);
xor U33522 (N_33522,N_32438,N_32235);
and U33523 (N_33523,N_32944,N_32205);
and U33524 (N_33524,N_32476,N_32776);
nor U33525 (N_33525,N_32115,N_32426);
nor U33526 (N_33526,N_32378,N_32050);
nand U33527 (N_33527,N_32885,N_32216);
xnor U33528 (N_33528,N_32025,N_32296);
xnor U33529 (N_33529,N_32659,N_32826);
and U33530 (N_33530,N_32649,N_32247);
or U33531 (N_33531,N_32441,N_32255);
nor U33532 (N_33532,N_32542,N_32637);
or U33533 (N_33533,N_32370,N_32656);
and U33534 (N_33534,N_32405,N_32436);
and U33535 (N_33535,N_32022,N_32772);
nand U33536 (N_33536,N_32344,N_32338);
nand U33537 (N_33537,N_32351,N_32766);
and U33538 (N_33538,N_32571,N_32789);
xnor U33539 (N_33539,N_32561,N_32027);
nand U33540 (N_33540,N_32138,N_32141);
nand U33541 (N_33541,N_32575,N_32741);
nor U33542 (N_33542,N_32427,N_32746);
and U33543 (N_33543,N_32698,N_32523);
nor U33544 (N_33544,N_32824,N_32101);
nor U33545 (N_33545,N_32352,N_32923);
nand U33546 (N_33546,N_32538,N_32805);
and U33547 (N_33547,N_32345,N_32199);
nor U33548 (N_33548,N_32644,N_32678);
nor U33549 (N_33549,N_32920,N_32290);
nand U33550 (N_33550,N_32514,N_32461);
xor U33551 (N_33551,N_32439,N_32153);
xor U33552 (N_33552,N_32239,N_32461);
nor U33553 (N_33553,N_32874,N_32539);
nor U33554 (N_33554,N_32967,N_32884);
nor U33555 (N_33555,N_32274,N_32169);
and U33556 (N_33556,N_32165,N_32326);
xnor U33557 (N_33557,N_32676,N_32515);
nor U33558 (N_33558,N_32700,N_32167);
nor U33559 (N_33559,N_32095,N_32980);
or U33560 (N_33560,N_32264,N_32397);
nor U33561 (N_33561,N_32245,N_32483);
nand U33562 (N_33562,N_32133,N_32875);
xnor U33563 (N_33563,N_32901,N_32606);
or U33564 (N_33564,N_32421,N_32721);
nand U33565 (N_33565,N_32712,N_32969);
or U33566 (N_33566,N_32242,N_32974);
nor U33567 (N_33567,N_32593,N_32175);
and U33568 (N_33568,N_32501,N_32957);
or U33569 (N_33569,N_32882,N_32536);
xor U33570 (N_33570,N_32404,N_32466);
and U33571 (N_33571,N_32345,N_32363);
or U33572 (N_33572,N_32428,N_32137);
and U33573 (N_33573,N_32318,N_32713);
and U33574 (N_33574,N_32487,N_32143);
and U33575 (N_33575,N_32242,N_32311);
xor U33576 (N_33576,N_32735,N_32215);
nor U33577 (N_33577,N_32894,N_32807);
nand U33578 (N_33578,N_32852,N_32672);
nand U33579 (N_33579,N_32953,N_32385);
or U33580 (N_33580,N_32500,N_32258);
nor U33581 (N_33581,N_32046,N_32181);
nor U33582 (N_33582,N_32090,N_32972);
or U33583 (N_33583,N_32919,N_32064);
xnor U33584 (N_33584,N_32250,N_32998);
or U33585 (N_33585,N_32222,N_32288);
xnor U33586 (N_33586,N_32548,N_32978);
nand U33587 (N_33587,N_32908,N_32594);
and U33588 (N_33588,N_32589,N_32540);
nand U33589 (N_33589,N_32182,N_32014);
nand U33590 (N_33590,N_32484,N_32359);
and U33591 (N_33591,N_32321,N_32377);
or U33592 (N_33592,N_32964,N_32466);
xnor U33593 (N_33593,N_32818,N_32999);
nor U33594 (N_33594,N_32605,N_32463);
nor U33595 (N_33595,N_32733,N_32392);
and U33596 (N_33596,N_32907,N_32023);
nand U33597 (N_33597,N_32857,N_32095);
nor U33598 (N_33598,N_32858,N_32603);
xnor U33599 (N_33599,N_32603,N_32203);
or U33600 (N_33600,N_32296,N_32875);
and U33601 (N_33601,N_32655,N_32876);
or U33602 (N_33602,N_32281,N_32896);
or U33603 (N_33603,N_32171,N_32554);
nor U33604 (N_33604,N_32666,N_32610);
and U33605 (N_33605,N_32336,N_32862);
nor U33606 (N_33606,N_32169,N_32045);
and U33607 (N_33607,N_32871,N_32096);
nand U33608 (N_33608,N_32360,N_32163);
xor U33609 (N_33609,N_32365,N_32690);
or U33610 (N_33610,N_32991,N_32172);
xnor U33611 (N_33611,N_32593,N_32983);
xor U33612 (N_33612,N_32519,N_32477);
and U33613 (N_33613,N_32066,N_32197);
and U33614 (N_33614,N_32026,N_32157);
or U33615 (N_33615,N_32385,N_32029);
or U33616 (N_33616,N_32189,N_32590);
xnor U33617 (N_33617,N_32179,N_32564);
or U33618 (N_33618,N_32482,N_32985);
and U33619 (N_33619,N_32865,N_32956);
and U33620 (N_33620,N_32562,N_32875);
and U33621 (N_33621,N_32408,N_32762);
and U33622 (N_33622,N_32088,N_32728);
nor U33623 (N_33623,N_32482,N_32481);
and U33624 (N_33624,N_32754,N_32867);
xnor U33625 (N_33625,N_32934,N_32736);
nor U33626 (N_33626,N_32684,N_32500);
nor U33627 (N_33627,N_32725,N_32826);
nor U33628 (N_33628,N_32228,N_32757);
or U33629 (N_33629,N_32909,N_32957);
and U33630 (N_33630,N_32870,N_32054);
or U33631 (N_33631,N_32128,N_32069);
xnor U33632 (N_33632,N_32278,N_32777);
xnor U33633 (N_33633,N_32397,N_32827);
or U33634 (N_33634,N_32862,N_32547);
nand U33635 (N_33635,N_32624,N_32698);
nand U33636 (N_33636,N_32442,N_32828);
or U33637 (N_33637,N_32829,N_32636);
nand U33638 (N_33638,N_32925,N_32678);
nand U33639 (N_33639,N_32780,N_32815);
xor U33640 (N_33640,N_32496,N_32930);
nand U33641 (N_33641,N_32870,N_32012);
or U33642 (N_33642,N_32058,N_32393);
nor U33643 (N_33643,N_32951,N_32574);
nand U33644 (N_33644,N_32584,N_32505);
nand U33645 (N_33645,N_32869,N_32604);
nand U33646 (N_33646,N_32356,N_32921);
or U33647 (N_33647,N_32757,N_32531);
or U33648 (N_33648,N_32765,N_32015);
and U33649 (N_33649,N_32012,N_32444);
xor U33650 (N_33650,N_32094,N_32630);
xor U33651 (N_33651,N_32837,N_32780);
or U33652 (N_33652,N_32082,N_32298);
or U33653 (N_33653,N_32879,N_32370);
or U33654 (N_33654,N_32836,N_32405);
xnor U33655 (N_33655,N_32248,N_32763);
and U33656 (N_33656,N_32640,N_32584);
and U33657 (N_33657,N_32120,N_32887);
nand U33658 (N_33658,N_32059,N_32701);
nor U33659 (N_33659,N_32395,N_32915);
nor U33660 (N_33660,N_32937,N_32882);
xor U33661 (N_33661,N_32156,N_32900);
or U33662 (N_33662,N_32079,N_32272);
or U33663 (N_33663,N_32489,N_32783);
nor U33664 (N_33664,N_32883,N_32983);
or U33665 (N_33665,N_32440,N_32155);
nor U33666 (N_33666,N_32163,N_32337);
and U33667 (N_33667,N_32839,N_32064);
nor U33668 (N_33668,N_32079,N_32442);
nand U33669 (N_33669,N_32526,N_32110);
or U33670 (N_33670,N_32270,N_32463);
nand U33671 (N_33671,N_32930,N_32611);
nand U33672 (N_33672,N_32412,N_32189);
and U33673 (N_33673,N_32634,N_32800);
and U33674 (N_33674,N_32110,N_32040);
or U33675 (N_33675,N_32778,N_32077);
and U33676 (N_33676,N_32104,N_32370);
nor U33677 (N_33677,N_32244,N_32826);
xnor U33678 (N_33678,N_32212,N_32021);
nor U33679 (N_33679,N_32485,N_32131);
or U33680 (N_33680,N_32645,N_32815);
xor U33681 (N_33681,N_32705,N_32124);
or U33682 (N_33682,N_32007,N_32991);
nor U33683 (N_33683,N_32040,N_32231);
nand U33684 (N_33684,N_32550,N_32463);
nor U33685 (N_33685,N_32124,N_32297);
or U33686 (N_33686,N_32362,N_32790);
or U33687 (N_33687,N_32566,N_32915);
or U33688 (N_33688,N_32737,N_32524);
and U33689 (N_33689,N_32024,N_32590);
and U33690 (N_33690,N_32177,N_32083);
and U33691 (N_33691,N_32473,N_32626);
xnor U33692 (N_33692,N_32961,N_32333);
nor U33693 (N_33693,N_32319,N_32875);
nand U33694 (N_33694,N_32190,N_32839);
xor U33695 (N_33695,N_32491,N_32078);
and U33696 (N_33696,N_32438,N_32957);
xor U33697 (N_33697,N_32923,N_32615);
and U33698 (N_33698,N_32484,N_32402);
nand U33699 (N_33699,N_32017,N_32893);
nor U33700 (N_33700,N_32668,N_32354);
nand U33701 (N_33701,N_32099,N_32791);
nand U33702 (N_33702,N_32490,N_32630);
nand U33703 (N_33703,N_32936,N_32020);
nor U33704 (N_33704,N_32641,N_32609);
or U33705 (N_33705,N_32297,N_32055);
and U33706 (N_33706,N_32891,N_32798);
or U33707 (N_33707,N_32524,N_32464);
xnor U33708 (N_33708,N_32484,N_32033);
nand U33709 (N_33709,N_32616,N_32026);
xnor U33710 (N_33710,N_32762,N_32931);
and U33711 (N_33711,N_32746,N_32389);
or U33712 (N_33712,N_32315,N_32884);
nor U33713 (N_33713,N_32819,N_32056);
nand U33714 (N_33714,N_32933,N_32048);
xor U33715 (N_33715,N_32368,N_32901);
xnor U33716 (N_33716,N_32791,N_32821);
nor U33717 (N_33717,N_32537,N_32555);
or U33718 (N_33718,N_32635,N_32733);
and U33719 (N_33719,N_32031,N_32726);
nor U33720 (N_33720,N_32763,N_32384);
and U33721 (N_33721,N_32898,N_32428);
and U33722 (N_33722,N_32136,N_32701);
and U33723 (N_33723,N_32743,N_32890);
or U33724 (N_33724,N_32115,N_32648);
nor U33725 (N_33725,N_32520,N_32508);
nand U33726 (N_33726,N_32224,N_32158);
nor U33727 (N_33727,N_32271,N_32048);
xnor U33728 (N_33728,N_32341,N_32896);
nand U33729 (N_33729,N_32176,N_32000);
xor U33730 (N_33730,N_32485,N_32496);
nand U33731 (N_33731,N_32850,N_32479);
or U33732 (N_33732,N_32388,N_32473);
nand U33733 (N_33733,N_32777,N_32691);
and U33734 (N_33734,N_32718,N_32949);
nor U33735 (N_33735,N_32489,N_32385);
xor U33736 (N_33736,N_32420,N_32628);
or U33737 (N_33737,N_32685,N_32292);
nor U33738 (N_33738,N_32242,N_32923);
or U33739 (N_33739,N_32667,N_32052);
and U33740 (N_33740,N_32278,N_32756);
nor U33741 (N_33741,N_32926,N_32082);
and U33742 (N_33742,N_32568,N_32038);
nand U33743 (N_33743,N_32653,N_32942);
nor U33744 (N_33744,N_32961,N_32683);
nor U33745 (N_33745,N_32352,N_32777);
or U33746 (N_33746,N_32716,N_32713);
or U33747 (N_33747,N_32983,N_32714);
and U33748 (N_33748,N_32432,N_32612);
or U33749 (N_33749,N_32550,N_32509);
nor U33750 (N_33750,N_32793,N_32357);
and U33751 (N_33751,N_32270,N_32310);
xor U33752 (N_33752,N_32938,N_32693);
nand U33753 (N_33753,N_32083,N_32706);
or U33754 (N_33754,N_32717,N_32997);
nand U33755 (N_33755,N_32920,N_32190);
or U33756 (N_33756,N_32889,N_32936);
or U33757 (N_33757,N_32287,N_32768);
nor U33758 (N_33758,N_32923,N_32883);
nand U33759 (N_33759,N_32860,N_32931);
xnor U33760 (N_33760,N_32581,N_32314);
or U33761 (N_33761,N_32486,N_32160);
nor U33762 (N_33762,N_32779,N_32761);
nor U33763 (N_33763,N_32182,N_32866);
nand U33764 (N_33764,N_32476,N_32681);
xnor U33765 (N_33765,N_32907,N_32260);
nand U33766 (N_33766,N_32324,N_32344);
xnor U33767 (N_33767,N_32292,N_32198);
xnor U33768 (N_33768,N_32763,N_32762);
and U33769 (N_33769,N_32176,N_32162);
and U33770 (N_33770,N_32484,N_32793);
and U33771 (N_33771,N_32498,N_32025);
xnor U33772 (N_33772,N_32337,N_32916);
and U33773 (N_33773,N_32295,N_32206);
or U33774 (N_33774,N_32610,N_32461);
nor U33775 (N_33775,N_32501,N_32174);
and U33776 (N_33776,N_32727,N_32688);
xor U33777 (N_33777,N_32933,N_32024);
nor U33778 (N_33778,N_32628,N_32368);
nor U33779 (N_33779,N_32885,N_32230);
and U33780 (N_33780,N_32035,N_32075);
nand U33781 (N_33781,N_32753,N_32805);
or U33782 (N_33782,N_32502,N_32060);
nor U33783 (N_33783,N_32084,N_32391);
nand U33784 (N_33784,N_32807,N_32302);
nor U33785 (N_33785,N_32722,N_32535);
nor U33786 (N_33786,N_32545,N_32381);
nand U33787 (N_33787,N_32060,N_32803);
nand U33788 (N_33788,N_32362,N_32754);
or U33789 (N_33789,N_32833,N_32480);
and U33790 (N_33790,N_32695,N_32201);
or U33791 (N_33791,N_32200,N_32321);
xnor U33792 (N_33792,N_32537,N_32666);
or U33793 (N_33793,N_32578,N_32301);
and U33794 (N_33794,N_32888,N_32911);
xor U33795 (N_33795,N_32007,N_32984);
nand U33796 (N_33796,N_32774,N_32854);
nor U33797 (N_33797,N_32988,N_32604);
nor U33798 (N_33798,N_32405,N_32221);
nand U33799 (N_33799,N_32318,N_32630);
nand U33800 (N_33800,N_32971,N_32099);
nand U33801 (N_33801,N_32553,N_32586);
xnor U33802 (N_33802,N_32005,N_32114);
nor U33803 (N_33803,N_32069,N_32971);
nor U33804 (N_33804,N_32408,N_32367);
xnor U33805 (N_33805,N_32018,N_32738);
xor U33806 (N_33806,N_32148,N_32149);
nand U33807 (N_33807,N_32079,N_32467);
nor U33808 (N_33808,N_32149,N_32397);
or U33809 (N_33809,N_32424,N_32042);
nor U33810 (N_33810,N_32233,N_32087);
or U33811 (N_33811,N_32071,N_32237);
nand U33812 (N_33812,N_32338,N_32475);
xor U33813 (N_33813,N_32389,N_32704);
or U33814 (N_33814,N_32297,N_32895);
and U33815 (N_33815,N_32235,N_32496);
or U33816 (N_33816,N_32147,N_32226);
or U33817 (N_33817,N_32125,N_32926);
nand U33818 (N_33818,N_32623,N_32061);
nor U33819 (N_33819,N_32736,N_32568);
nor U33820 (N_33820,N_32827,N_32909);
nor U33821 (N_33821,N_32980,N_32300);
nand U33822 (N_33822,N_32981,N_32293);
nand U33823 (N_33823,N_32350,N_32180);
and U33824 (N_33824,N_32550,N_32238);
nor U33825 (N_33825,N_32579,N_32246);
nand U33826 (N_33826,N_32483,N_32448);
xor U33827 (N_33827,N_32993,N_32009);
nand U33828 (N_33828,N_32127,N_32535);
xor U33829 (N_33829,N_32131,N_32653);
xor U33830 (N_33830,N_32745,N_32804);
nor U33831 (N_33831,N_32696,N_32714);
xnor U33832 (N_33832,N_32365,N_32735);
nor U33833 (N_33833,N_32936,N_32024);
xnor U33834 (N_33834,N_32711,N_32838);
or U33835 (N_33835,N_32022,N_32302);
or U33836 (N_33836,N_32203,N_32647);
xnor U33837 (N_33837,N_32782,N_32257);
xnor U33838 (N_33838,N_32467,N_32741);
nor U33839 (N_33839,N_32761,N_32723);
or U33840 (N_33840,N_32874,N_32926);
nand U33841 (N_33841,N_32470,N_32307);
nand U33842 (N_33842,N_32564,N_32483);
or U33843 (N_33843,N_32756,N_32569);
and U33844 (N_33844,N_32364,N_32604);
nand U33845 (N_33845,N_32492,N_32129);
nand U33846 (N_33846,N_32595,N_32314);
xnor U33847 (N_33847,N_32869,N_32809);
xor U33848 (N_33848,N_32936,N_32960);
xnor U33849 (N_33849,N_32419,N_32443);
nand U33850 (N_33850,N_32484,N_32001);
nand U33851 (N_33851,N_32390,N_32153);
xor U33852 (N_33852,N_32731,N_32202);
or U33853 (N_33853,N_32387,N_32983);
nor U33854 (N_33854,N_32753,N_32164);
xor U33855 (N_33855,N_32551,N_32746);
nand U33856 (N_33856,N_32168,N_32936);
xor U33857 (N_33857,N_32383,N_32808);
nor U33858 (N_33858,N_32335,N_32621);
and U33859 (N_33859,N_32383,N_32089);
nor U33860 (N_33860,N_32730,N_32845);
xnor U33861 (N_33861,N_32341,N_32659);
xnor U33862 (N_33862,N_32369,N_32566);
nor U33863 (N_33863,N_32098,N_32052);
nor U33864 (N_33864,N_32581,N_32529);
xnor U33865 (N_33865,N_32915,N_32943);
nor U33866 (N_33866,N_32904,N_32958);
nor U33867 (N_33867,N_32353,N_32539);
nand U33868 (N_33868,N_32185,N_32759);
or U33869 (N_33869,N_32888,N_32392);
and U33870 (N_33870,N_32488,N_32241);
nand U33871 (N_33871,N_32002,N_32669);
nand U33872 (N_33872,N_32954,N_32995);
and U33873 (N_33873,N_32257,N_32683);
nand U33874 (N_33874,N_32913,N_32476);
nand U33875 (N_33875,N_32135,N_32638);
nor U33876 (N_33876,N_32538,N_32791);
nand U33877 (N_33877,N_32062,N_32765);
nand U33878 (N_33878,N_32299,N_32597);
xor U33879 (N_33879,N_32985,N_32586);
nand U33880 (N_33880,N_32807,N_32939);
and U33881 (N_33881,N_32389,N_32904);
nor U33882 (N_33882,N_32323,N_32383);
nor U33883 (N_33883,N_32133,N_32565);
nand U33884 (N_33884,N_32717,N_32204);
nand U33885 (N_33885,N_32561,N_32698);
nor U33886 (N_33886,N_32287,N_32208);
nand U33887 (N_33887,N_32597,N_32701);
or U33888 (N_33888,N_32108,N_32730);
or U33889 (N_33889,N_32410,N_32104);
or U33890 (N_33890,N_32949,N_32257);
or U33891 (N_33891,N_32276,N_32396);
or U33892 (N_33892,N_32974,N_32777);
and U33893 (N_33893,N_32366,N_32022);
or U33894 (N_33894,N_32805,N_32149);
nand U33895 (N_33895,N_32721,N_32031);
nand U33896 (N_33896,N_32164,N_32713);
nor U33897 (N_33897,N_32592,N_32593);
nand U33898 (N_33898,N_32176,N_32535);
nand U33899 (N_33899,N_32082,N_32025);
and U33900 (N_33900,N_32219,N_32149);
nand U33901 (N_33901,N_32543,N_32168);
nand U33902 (N_33902,N_32088,N_32256);
nor U33903 (N_33903,N_32461,N_32839);
xnor U33904 (N_33904,N_32402,N_32598);
or U33905 (N_33905,N_32920,N_32132);
nor U33906 (N_33906,N_32442,N_32599);
nand U33907 (N_33907,N_32148,N_32729);
xor U33908 (N_33908,N_32381,N_32380);
nor U33909 (N_33909,N_32068,N_32783);
nor U33910 (N_33910,N_32161,N_32536);
nand U33911 (N_33911,N_32069,N_32757);
nand U33912 (N_33912,N_32124,N_32728);
or U33913 (N_33913,N_32831,N_32313);
and U33914 (N_33914,N_32757,N_32263);
and U33915 (N_33915,N_32373,N_32191);
or U33916 (N_33916,N_32312,N_32060);
or U33917 (N_33917,N_32098,N_32416);
nor U33918 (N_33918,N_32875,N_32660);
nor U33919 (N_33919,N_32514,N_32296);
nand U33920 (N_33920,N_32167,N_32413);
or U33921 (N_33921,N_32141,N_32709);
xor U33922 (N_33922,N_32460,N_32426);
and U33923 (N_33923,N_32515,N_32103);
nand U33924 (N_33924,N_32131,N_32868);
nor U33925 (N_33925,N_32475,N_32278);
xor U33926 (N_33926,N_32239,N_32573);
nor U33927 (N_33927,N_32017,N_32782);
or U33928 (N_33928,N_32074,N_32174);
nand U33929 (N_33929,N_32546,N_32139);
nor U33930 (N_33930,N_32354,N_32311);
or U33931 (N_33931,N_32899,N_32699);
nor U33932 (N_33932,N_32052,N_32454);
nand U33933 (N_33933,N_32493,N_32223);
or U33934 (N_33934,N_32274,N_32693);
xor U33935 (N_33935,N_32080,N_32116);
or U33936 (N_33936,N_32546,N_32103);
and U33937 (N_33937,N_32134,N_32775);
or U33938 (N_33938,N_32138,N_32071);
nand U33939 (N_33939,N_32096,N_32884);
nand U33940 (N_33940,N_32131,N_32711);
nor U33941 (N_33941,N_32548,N_32345);
nor U33942 (N_33942,N_32474,N_32088);
nor U33943 (N_33943,N_32737,N_32061);
nor U33944 (N_33944,N_32836,N_32406);
and U33945 (N_33945,N_32665,N_32249);
and U33946 (N_33946,N_32139,N_32611);
or U33947 (N_33947,N_32072,N_32821);
and U33948 (N_33948,N_32708,N_32627);
xnor U33949 (N_33949,N_32575,N_32554);
nand U33950 (N_33950,N_32173,N_32474);
and U33951 (N_33951,N_32277,N_32584);
or U33952 (N_33952,N_32069,N_32193);
xor U33953 (N_33953,N_32823,N_32954);
xor U33954 (N_33954,N_32617,N_32257);
nand U33955 (N_33955,N_32570,N_32491);
and U33956 (N_33956,N_32913,N_32958);
nand U33957 (N_33957,N_32239,N_32870);
nand U33958 (N_33958,N_32244,N_32963);
xor U33959 (N_33959,N_32800,N_32610);
and U33960 (N_33960,N_32267,N_32384);
nand U33961 (N_33961,N_32026,N_32130);
or U33962 (N_33962,N_32494,N_32704);
xor U33963 (N_33963,N_32539,N_32444);
nor U33964 (N_33964,N_32525,N_32239);
and U33965 (N_33965,N_32396,N_32350);
nand U33966 (N_33966,N_32882,N_32274);
nor U33967 (N_33967,N_32158,N_32567);
xnor U33968 (N_33968,N_32944,N_32755);
xnor U33969 (N_33969,N_32527,N_32814);
or U33970 (N_33970,N_32832,N_32943);
nand U33971 (N_33971,N_32917,N_32976);
xor U33972 (N_33972,N_32243,N_32868);
and U33973 (N_33973,N_32679,N_32393);
nor U33974 (N_33974,N_32052,N_32368);
or U33975 (N_33975,N_32461,N_32730);
nand U33976 (N_33976,N_32943,N_32590);
nand U33977 (N_33977,N_32327,N_32681);
and U33978 (N_33978,N_32115,N_32968);
nor U33979 (N_33979,N_32004,N_32359);
nor U33980 (N_33980,N_32398,N_32502);
nor U33981 (N_33981,N_32632,N_32053);
nand U33982 (N_33982,N_32335,N_32927);
and U33983 (N_33983,N_32184,N_32407);
or U33984 (N_33984,N_32607,N_32538);
or U33985 (N_33985,N_32368,N_32575);
and U33986 (N_33986,N_32826,N_32027);
nor U33987 (N_33987,N_32949,N_32799);
xor U33988 (N_33988,N_32390,N_32624);
xor U33989 (N_33989,N_32142,N_32217);
and U33990 (N_33990,N_32566,N_32762);
and U33991 (N_33991,N_32746,N_32925);
and U33992 (N_33992,N_32998,N_32119);
and U33993 (N_33993,N_32058,N_32707);
or U33994 (N_33994,N_32503,N_32656);
nand U33995 (N_33995,N_32469,N_32447);
nand U33996 (N_33996,N_32712,N_32063);
nor U33997 (N_33997,N_32574,N_32276);
and U33998 (N_33998,N_32098,N_32809);
xnor U33999 (N_33999,N_32711,N_32065);
nand U34000 (N_34000,N_33391,N_33093);
nand U34001 (N_34001,N_33244,N_33084);
nor U34002 (N_34002,N_33740,N_33025);
or U34003 (N_34003,N_33905,N_33778);
xnor U34004 (N_34004,N_33017,N_33976);
nand U34005 (N_34005,N_33207,N_33801);
nand U34006 (N_34006,N_33247,N_33262);
nand U34007 (N_34007,N_33121,N_33339);
xor U34008 (N_34008,N_33486,N_33419);
nor U34009 (N_34009,N_33162,N_33399);
xnor U34010 (N_34010,N_33811,N_33837);
or U34011 (N_34011,N_33474,N_33846);
or U34012 (N_34012,N_33444,N_33424);
and U34013 (N_34013,N_33351,N_33713);
or U34014 (N_34014,N_33089,N_33189);
nor U34015 (N_34015,N_33428,N_33029);
or U34016 (N_34016,N_33632,N_33874);
or U34017 (N_34017,N_33180,N_33500);
and U34018 (N_34018,N_33229,N_33015);
nand U34019 (N_34019,N_33758,N_33276);
nand U34020 (N_34020,N_33807,N_33042);
and U34021 (N_34021,N_33831,N_33800);
nor U34022 (N_34022,N_33509,N_33969);
or U34023 (N_34023,N_33642,N_33943);
or U34024 (N_34024,N_33558,N_33160);
or U34025 (N_34025,N_33527,N_33796);
and U34026 (N_34026,N_33265,N_33252);
nand U34027 (N_34027,N_33933,N_33885);
nor U34028 (N_34028,N_33454,N_33353);
and U34029 (N_34029,N_33103,N_33693);
or U34030 (N_34030,N_33838,N_33478);
xnor U34031 (N_34031,N_33350,N_33201);
xnor U34032 (N_34032,N_33716,N_33623);
nand U34033 (N_34033,N_33111,N_33222);
xor U34034 (N_34034,N_33223,N_33074);
xnor U34035 (N_34035,N_33116,N_33571);
or U34036 (N_34036,N_33856,N_33185);
and U34037 (N_34037,N_33128,N_33033);
xor U34038 (N_34038,N_33470,N_33132);
and U34039 (N_34039,N_33021,N_33375);
or U34040 (N_34040,N_33164,N_33117);
or U34041 (N_34041,N_33062,N_33555);
xnor U34042 (N_34042,N_33827,N_33651);
or U34043 (N_34043,N_33151,N_33621);
xor U34044 (N_34044,N_33041,N_33863);
or U34045 (N_34045,N_33982,N_33175);
nand U34046 (N_34046,N_33987,N_33589);
nor U34047 (N_34047,N_33767,N_33759);
xor U34048 (N_34048,N_33371,N_33163);
nor U34049 (N_34049,N_33464,N_33274);
and U34050 (N_34050,N_33110,N_33628);
nor U34051 (N_34051,N_33820,N_33453);
nand U34052 (N_34052,N_33303,N_33152);
or U34053 (N_34053,N_33726,N_33815);
nand U34054 (N_34054,N_33902,N_33887);
nand U34055 (N_34055,N_33279,N_33656);
xnor U34056 (N_34056,N_33173,N_33669);
nand U34057 (N_34057,N_33101,N_33365);
nand U34058 (N_34058,N_33433,N_33508);
and U34059 (N_34059,N_33733,N_33840);
nand U34060 (N_34060,N_33954,N_33872);
xor U34061 (N_34061,N_33217,N_33280);
or U34062 (N_34062,N_33978,N_33221);
nand U34063 (N_34063,N_33919,N_33067);
and U34064 (N_34064,N_33552,N_33005);
nand U34065 (N_34065,N_33209,N_33810);
and U34066 (N_34066,N_33225,N_33034);
and U34067 (N_34067,N_33519,N_33564);
or U34068 (N_34068,N_33142,N_33940);
nor U34069 (N_34069,N_33497,N_33580);
nand U34070 (N_34070,N_33451,N_33398);
nand U34071 (N_34071,N_33756,N_33772);
nor U34072 (N_34072,N_33836,N_33662);
nor U34073 (N_34073,N_33842,N_33996);
xnor U34074 (N_34074,N_33925,N_33789);
nand U34075 (N_34075,N_33737,N_33141);
or U34076 (N_34076,N_33296,N_33866);
or U34077 (N_34077,N_33561,N_33544);
and U34078 (N_34078,N_33430,N_33039);
or U34079 (N_34079,N_33283,N_33408);
xor U34080 (N_34080,N_33931,N_33830);
xor U34081 (N_34081,N_33968,N_33898);
and U34082 (N_34082,N_33546,N_33425);
nand U34083 (N_34083,N_33153,N_33698);
nor U34084 (N_34084,N_33166,N_33984);
nor U34085 (N_34085,N_33794,N_33333);
nor U34086 (N_34086,N_33625,N_33683);
xor U34087 (N_34087,N_33602,N_33514);
xnor U34088 (N_34088,N_33786,N_33790);
and U34089 (N_34089,N_33219,N_33300);
and U34090 (N_34090,N_33921,N_33890);
nand U34091 (N_34091,N_33374,N_33633);
nand U34092 (N_34092,N_33870,N_33728);
or U34093 (N_34093,N_33597,N_33009);
and U34094 (N_34094,N_33727,N_33073);
nand U34095 (N_34095,N_33245,N_33417);
xnor U34096 (N_34096,N_33441,N_33748);
nand U34097 (N_34097,N_33057,N_33672);
nand U34098 (N_34098,N_33338,N_33520);
or U34099 (N_34099,N_33904,N_33650);
nand U34100 (N_34100,N_33377,N_33473);
xnor U34101 (N_34101,N_33992,N_33566);
nor U34102 (N_34102,N_33403,N_33595);
xor U34103 (N_34103,N_33719,N_33886);
and U34104 (N_34104,N_33498,N_33354);
xor U34105 (N_34105,N_33055,N_33660);
nor U34106 (N_34106,N_33190,N_33257);
and U34107 (N_34107,N_33240,N_33658);
and U34108 (N_34108,N_33368,N_33634);
or U34109 (N_34109,N_33238,N_33367);
nor U34110 (N_34110,N_33620,N_33802);
nor U34111 (N_34111,N_33445,N_33576);
nand U34112 (N_34112,N_33619,N_33959);
nand U34113 (N_34113,N_33237,N_33636);
or U34114 (N_34114,N_33246,N_33673);
or U34115 (N_34115,N_33379,N_33331);
and U34116 (N_34116,N_33069,N_33168);
xor U34117 (N_34117,N_33948,N_33679);
nand U34118 (N_34118,N_33051,N_33819);
nand U34119 (N_34119,N_33458,N_33661);
and U34120 (N_34120,N_33394,N_33410);
and U34121 (N_34121,N_33926,N_33888);
nand U34122 (N_34122,N_33554,N_33980);
xor U34123 (N_34123,N_33951,N_33289);
nor U34124 (N_34124,N_33917,N_33321);
and U34125 (N_34125,N_33710,N_33050);
nor U34126 (N_34126,N_33202,N_33267);
and U34127 (N_34127,N_33239,N_33193);
or U34128 (N_34128,N_33220,N_33360);
or U34129 (N_34129,N_33357,N_33736);
nor U34130 (N_34130,N_33007,N_33730);
and U34131 (N_34131,N_33533,N_33569);
or U34132 (N_34132,N_33174,N_33944);
or U34133 (N_34133,N_33749,N_33287);
nand U34134 (N_34134,N_33884,N_33956);
xor U34135 (N_34135,N_33385,N_33143);
and U34136 (N_34136,N_33440,N_33938);
and U34137 (N_34137,N_33609,N_33182);
and U34138 (N_34138,N_33139,N_33889);
xnor U34139 (N_34139,N_33114,N_33415);
and U34140 (N_34140,N_33517,N_33288);
or U34141 (N_34141,N_33857,N_33102);
or U34142 (N_34142,N_33460,N_33924);
and U34143 (N_34143,N_33064,N_33438);
and U34144 (N_34144,N_33822,N_33032);
nand U34145 (N_34145,N_33195,N_33284);
xnor U34146 (N_34146,N_33665,N_33475);
nor U34147 (N_34147,N_33977,N_33323);
nor U34148 (N_34148,N_33918,N_33541);
xor U34149 (N_34149,N_33655,N_33027);
xor U34150 (N_34150,N_33178,N_33505);
nand U34151 (N_34151,N_33910,N_33694);
nand U34152 (N_34152,N_33332,N_33040);
or U34153 (N_34153,N_33056,N_33302);
nand U34154 (N_34154,N_33706,N_33528);
nor U34155 (N_34155,N_33226,N_33090);
nor U34156 (N_34156,N_33002,N_33799);
nor U34157 (N_34157,N_33426,N_33795);
nand U34158 (N_34158,N_33078,N_33753);
or U34159 (N_34159,N_33663,N_33932);
xor U34160 (N_34160,N_33316,N_33746);
xor U34161 (N_34161,N_33738,N_33306);
or U34162 (N_34162,N_33409,N_33031);
xor U34163 (N_34163,N_33477,N_33218);
xor U34164 (N_34164,N_33468,N_33515);
or U34165 (N_34165,N_33411,N_33404);
and U34166 (N_34166,N_33818,N_33605);
nand U34167 (N_34167,N_33309,N_33355);
and U34168 (N_34168,N_33305,N_33432);
xnor U34169 (N_34169,N_33135,N_33522);
xnor U34170 (N_34170,N_33825,N_33471);
or U34171 (N_34171,N_33494,N_33823);
and U34172 (N_34172,N_33947,N_33086);
and U34173 (N_34173,N_33942,N_33161);
nor U34174 (N_34174,N_33205,N_33782);
xnor U34175 (N_34175,N_33503,N_33028);
nand U34176 (N_34176,N_33264,N_33567);
or U34177 (N_34177,N_33638,N_33784);
nor U34178 (N_34178,N_33158,N_33608);
and U34179 (N_34179,N_33995,N_33349);
or U34180 (N_34180,N_33647,N_33115);
nor U34181 (N_34181,N_33335,N_33523);
nand U34182 (N_34182,N_33418,N_33540);
and U34183 (N_34183,N_33845,N_33294);
or U34184 (N_34184,N_33681,N_33715);
xnor U34185 (N_34185,N_33461,N_33450);
and U34186 (N_34186,N_33493,N_33388);
xnor U34187 (N_34187,N_33053,N_33573);
and U34188 (N_34188,N_33973,N_33868);
and U34189 (N_34189,N_33312,N_33295);
xor U34190 (N_34190,N_33853,N_33008);
and U34191 (N_34191,N_33490,N_33369);
nor U34192 (N_34192,N_33297,N_33072);
and U34193 (N_34193,N_33626,N_33939);
nand U34194 (N_34194,N_33991,N_33666);
nor U34195 (N_34195,N_33499,N_33582);
nand U34196 (N_34196,N_33641,N_33136);
xor U34197 (N_34197,N_33048,N_33556);
nor U34198 (N_34198,N_33196,N_33104);
xor U34199 (N_34199,N_33186,N_33495);
xor U34200 (N_34200,N_33725,N_33993);
nor U34201 (N_34201,N_33149,N_33382);
nand U34202 (N_34202,N_33763,N_33286);
and U34203 (N_34203,N_33322,N_33742);
or U34204 (N_34204,N_33496,N_33512);
nor U34205 (N_34205,N_33058,N_33913);
nand U34206 (N_34206,N_33466,N_33233);
nand U34207 (N_34207,N_33106,N_33584);
and U34208 (N_34208,N_33705,N_33272);
or U34209 (N_34209,N_33832,N_33934);
and U34210 (N_34210,N_33513,N_33397);
and U34211 (N_34211,N_33950,N_33762);
or U34212 (N_34212,N_33961,N_33347);
xor U34213 (N_34213,N_33212,N_33170);
or U34214 (N_34214,N_33861,N_33797);
and U34215 (N_34215,N_33405,N_33018);
or U34216 (N_34216,N_33817,N_33529);
and U34217 (N_34217,N_33277,N_33120);
or U34218 (N_34218,N_33336,N_33364);
xnor U34219 (N_34219,N_33834,N_33109);
and U34220 (N_34220,N_33974,N_33581);
nor U34221 (N_34221,N_33760,N_33975);
xnor U34222 (N_34222,N_33045,N_33629);
and U34223 (N_34223,N_33506,N_33376);
nor U34224 (N_34224,N_33776,N_33310);
and U34225 (N_34225,N_33957,N_33894);
xor U34226 (N_34226,N_33721,N_33682);
nand U34227 (N_34227,N_33821,N_33138);
nor U34228 (N_34228,N_33273,N_33215);
nor U34229 (N_34229,N_33436,N_33431);
nor U34230 (N_34230,N_33092,N_33646);
nor U34231 (N_34231,N_33537,N_33446);
nand U34232 (N_34232,N_33775,N_33687);
nor U34233 (N_34233,N_33159,N_33026);
nor U34234 (N_34234,N_33600,N_33402);
xnor U34235 (N_34235,N_33922,N_33019);
xor U34236 (N_34236,N_33812,N_33228);
nor U34237 (N_34237,N_33912,N_33911);
nor U34238 (N_34238,N_33697,N_33722);
xnor U34239 (N_34239,N_33971,N_33813);
nand U34240 (N_34240,N_33988,N_33044);
and U34241 (N_34241,N_33507,N_33862);
xor U34242 (N_34242,N_33770,N_33952);
nor U34243 (N_34243,N_33096,N_33439);
nand U34244 (N_34244,N_33614,N_33340);
xnor U34245 (N_34245,N_33598,N_33603);
xnor U34246 (N_34246,N_33230,N_33144);
and U34247 (N_34247,N_33407,N_33744);
or U34248 (N_34248,N_33345,N_33551);
or U34249 (N_34249,N_33105,N_33792);
nand U34250 (N_34250,N_33459,N_33396);
and U34251 (N_34251,N_33487,N_33895);
and U34252 (N_34252,N_33334,N_33085);
nand U34253 (N_34253,N_33291,N_33437);
nor U34254 (N_34254,N_33480,N_33516);
or U34255 (N_34255,N_33997,N_33774);
nor U34256 (N_34256,N_33081,N_33545);
xor U34257 (N_34257,N_33535,N_33615);
nor U34258 (N_34258,N_33877,N_33181);
xor U34259 (N_34259,N_33465,N_33577);
nand U34260 (N_34260,N_33717,N_33313);
xnor U34261 (N_34261,N_33701,N_33985);
and U34262 (N_34262,N_33501,N_33275);
nand U34263 (N_34263,N_33937,N_33955);
nand U34264 (N_34264,N_33667,N_33400);
and U34265 (N_34265,N_33876,N_33630);
or U34266 (N_34266,N_33518,N_33456);
and U34267 (N_34267,N_33611,N_33060);
or U34268 (N_34268,N_33263,N_33652);
xor U34269 (N_34269,N_33688,N_33356);
or U34270 (N_34270,N_33278,N_33617);
or U34271 (N_34271,N_33211,N_33986);
or U34272 (N_34272,N_33392,N_33147);
or U34273 (N_34273,N_33406,N_33686);
nor U34274 (N_34274,N_33401,N_33542);
nand U34275 (N_34275,N_33864,N_33140);
and U34276 (N_34276,N_33435,N_33935);
or U34277 (N_34277,N_33256,N_33750);
nor U34278 (N_34278,N_33447,N_33998);
xnor U34279 (N_34279,N_33122,N_33780);
nor U34280 (N_34280,N_33900,N_33261);
nand U34281 (N_34281,N_33668,N_33718);
or U34282 (N_34282,N_33378,N_33003);
xnor U34283 (N_34283,N_33735,N_33803);
nand U34284 (N_34284,N_33983,N_33671);
xor U34285 (N_34285,N_33188,N_33916);
and U34286 (N_34286,N_33119,N_33224);
or U34287 (N_34287,N_33416,N_33964);
xnor U34288 (N_34288,N_33013,N_33659);
nand U34289 (N_34289,N_33893,N_33269);
and U34290 (N_34290,N_33216,N_33878);
nand U34291 (N_34291,N_33414,N_33094);
nor U34292 (N_34292,N_33568,N_33268);
nor U34293 (N_34293,N_33348,N_33704);
nand U34294 (N_34294,N_33150,N_33685);
xor U34295 (N_34295,N_33071,N_33384);
xnor U34296 (N_34296,N_33881,N_33342);
nand U34297 (N_34297,N_33765,N_33046);
and U34298 (N_34298,N_33783,N_33363);
nor U34299 (N_34299,N_33729,N_33994);
or U34300 (N_34300,N_33443,N_33696);
nor U34301 (N_34301,N_33301,N_33107);
or U34302 (N_34302,N_33241,N_33747);
nor U34303 (N_34303,N_33361,N_33112);
or U34304 (N_34304,N_33066,N_33882);
and U34305 (N_34305,N_33847,N_33324);
or U34306 (N_34306,N_33359,N_33731);
and U34307 (N_34307,N_33526,N_33587);
or U34308 (N_34308,N_33087,N_33824);
and U34309 (N_34309,N_33012,N_33966);
nor U34310 (N_34310,N_33052,N_33664);
nand U34311 (N_34311,N_33036,N_33172);
or U34312 (N_34312,N_33165,N_33091);
or U34313 (N_34313,N_33734,N_33231);
xnor U34314 (N_34314,N_33849,N_33146);
xnor U34315 (N_34315,N_33328,N_33908);
nor U34316 (N_34316,N_33043,N_33548);
or U34317 (N_34317,N_33370,N_33627);
nand U34318 (N_34318,N_33179,N_33176);
or U34319 (N_34319,N_33023,N_33773);
nor U34320 (N_34320,N_33809,N_33213);
nand U34321 (N_34321,N_33206,N_33798);
nand U34322 (N_34322,N_33896,N_33909);
xnor U34323 (N_34323,N_33214,N_33826);
or U34324 (N_34324,N_33038,N_33427);
nor U34325 (N_34325,N_33907,N_33711);
nand U34326 (N_34326,N_33703,N_33253);
and U34327 (N_34327,N_33255,N_33967);
nand U34328 (N_34328,N_33549,N_33271);
nor U34329 (N_34329,N_33972,N_33199);
or U34330 (N_34330,N_33793,N_33344);
xor U34331 (N_34331,N_33386,N_33352);
or U34332 (N_34332,N_33787,N_33557);
and U34333 (N_34333,N_33184,N_33065);
or U34334 (N_34334,N_33599,N_33155);
or U34335 (N_34335,N_33327,N_33648);
and U34336 (N_34336,N_33844,N_33852);
or U34337 (N_34337,N_33137,N_33393);
nand U34338 (N_34338,N_33788,N_33806);
or U34339 (N_34339,N_33565,N_33127);
and U34340 (N_34340,N_33187,N_33607);
nand U34341 (N_34341,N_33011,N_33004);
nor U34342 (N_34342,N_33854,N_33936);
nor U34343 (N_34343,N_33691,N_33200);
and U34344 (N_34344,N_33743,N_33191);
nor U34345 (N_34345,N_33307,N_33962);
nor U34346 (N_34346,N_33892,N_33828);
or U34347 (N_34347,N_33290,N_33479);
or U34348 (N_34348,N_33583,N_33999);
and U34349 (N_34349,N_33875,N_33308);
nor U34350 (N_34350,N_33123,N_33644);
nor U34351 (N_34351,N_33572,N_33035);
nand U34352 (N_34352,N_33129,N_33330);
and U34353 (N_34353,N_33260,N_33304);
nor U34354 (N_34354,N_33755,N_33315);
nand U34355 (N_34355,N_33649,N_33871);
or U34356 (N_34356,N_33325,N_33539);
xor U34357 (N_34357,N_33848,N_33547);
nor U34358 (N_34358,N_33596,N_33457);
or U34359 (N_34359,N_33318,N_33741);
or U34360 (N_34360,N_33204,N_33841);
xnor U34361 (N_34361,N_33677,N_33593);
xor U34362 (N_34362,N_33346,N_33250);
nor U34363 (N_34363,N_33531,N_33097);
nor U34364 (N_34364,N_33413,N_33720);
nor U34365 (N_34365,N_33622,N_33192);
and U34366 (N_34366,N_33030,N_33242);
or U34367 (N_34367,N_33618,N_33859);
xor U34368 (N_34368,N_33771,N_33707);
and U34369 (N_34369,N_33024,N_33804);
nor U34370 (N_34370,N_33285,N_33873);
xnor U34371 (N_34371,N_33167,N_33754);
and U34372 (N_34372,N_33502,N_33157);
and U34373 (N_34373,N_33680,N_33927);
or U34374 (N_34374,N_33578,N_33319);
nand U34375 (N_34375,N_33326,N_33076);
nor U34376 (N_34376,N_33083,N_33850);
xnor U34377 (N_34377,N_33521,N_33098);
xnor U34378 (N_34378,N_33366,N_33752);
xor U34379 (N_34379,N_33171,N_33766);
and U34380 (N_34380,N_33169,N_33113);
or U34381 (N_34381,N_33234,N_33075);
nand U34382 (N_34382,N_33266,N_33805);
and U34383 (N_34383,N_33684,N_33610);
nand U34384 (N_34384,N_33254,N_33989);
or U34385 (N_34385,N_33640,N_33745);
nand U34386 (N_34386,N_33851,N_33880);
nand U34387 (N_34387,N_33695,N_33867);
or U34388 (N_34388,N_33063,N_33455);
xor U34389 (N_34389,N_33442,N_33777);
and U34390 (N_34390,N_33329,N_33906);
xnor U34391 (N_34391,N_33133,N_33243);
xor U34392 (N_34392,N_33963,N_33020);
nand U34393 (N_34393,N_33631,N_33899);
xnor U34394 (N_34394,N_33082,N_33420);
and U34395 (N_34395,N_33709,N_33785);
nand U34396 (N_34396,N_33808,N_33606);
nand U34397 (N_34397,N_33390,N_33643);
nand U34398 (N_34398,N_33362,N_33080);
nand U34399 (N_34399,N_33903,N_33270);
and U34400 (N_34400,N_33865,N_33492);
nand U34401 (N_34401,N_33714,N_33412);
xor U34402 (N_34402,N_33676,N_33941);
or U34403 (N_34403,N_33463,N_33945);
and U34404 (N_34404,N_33299,N_33781);
nor U34405 (N_34405,N_33482,N_33022);
xor U34406 (N_34406,N_33281,N_33645);
nor U34407 (N_34407,N_33177,N_33635);
or U34408 (N_34408,N_33381,N_33469);
or U34409 (N_34409,N_33485,N_33699);
or U34410 (N_34410,N_33203,N_33049);
xnor U34411 (N_34411,N_33897,N_33570);
xnor U34412 (N_34412,N_33946,N_33616);
nand U34413 (N_34413,N_33833,N_33197);
and U34414 (N_34414,N_33915,N_33990);
nand U34415 (N_34415,N_33488,N_33768);
and U34416 (N_34416,N_33511,N_33712);
nand U34417 (N_34417,N_33575,N_33449);
nor U34418 (N_34418,N_33525,N_33373);
nor U34419 (N_34419,N_33380,N_33708);
or U34420 (N_34420,N_33550,N_33586);
xor U34421 (N_34421,N_33452,N_33125);
or U34422 (N_34422,N_33757,N_33613);
xnor U34423 (N_34423,N_33657,N_33981);
nand U34424 (N_34424,N_33588,N_33965);
or U34425 (N_34425,N_33769,N_33227);
or U34426 (N_34426,N_33481,N_33108);
nor U34427 (N_34427,N_33949,N_33524);
nor U34428 (N_34428,N_33637,N_33429);
nor U34429 (N_34429,N_33958,N_33210);
and U34430 (N_34430,N_33732,N_33510);
nand U34431 (N_34431,N_33879,N_33145);
nor U34432 (N_34432,N_33387,N_33723);
nand U34433 (N_34433,N_33536,N_33010);
nor U34434 (N_34434,N_33670,N_33448);
nand U34435 (N_34435,N_33421,N_33592);
and U34436 (N_34436,N_33100,N_33118);
or U34437 (N_34437,N_33530,N_33692);
and U34438 (N_34438,N_33014,N_33232);
nand U34439 (N_34439,N_33534,N_33001);
nor U34440 (N_34440,N_33320,N_33483);
and U34441 (N_34441,N_33248,N_33395);
xnor U34442 (N_34442,N_33604,N_33675);
xnor U34443 (N_34443,N_33624,N_33532);
nand U34444 (N_34444,N_33960,N_33317);
xor U34445 (N_34445,N_33282,N_33472);
nor U34446 (N_34446,N_33061,N_33489);
or U34447 (N_34447,N_33389,N_33088);
nor U34448 (N_34448,N_33126,N_33923);
or U34449 (N_34449,N_33292,N_33343);
nand U34450 (N_34450,N_33654,N_33538);
xor U34451 (N_34451,N_33891,N_33678);
xnor U34452 (N_34452,N_33724,N_33970);
and U34453 (N_34453,N_33979,N_33124);
nor U34454 (N_34454,N_33869,N_33612);
or U34455 (N_34455,N_33068,N_33751);
nor U34456 (N_34456,N_33079,N_33835);
and U34457 (N_34457,N_33858,N_33953);
or U34458 (N_34458,N_33814,N_33690);
xnor U34459 (N_34459,N_33816,N_33249);
xnor U34460 (N_34460,N_33462,N_33594);
or U34461 (N_34461,N_33341,N_33562);
nand U34462 (N_34462,N_33761,N_33883);
xor U34463 (N_34463,N_33251,N_33423);
xnor U34464 (N_34464,N_33198,N_33259);
nor U34465 (N_34465,N_33574,N_33000);
and U34466 (N_34466,N_33553,N_33579);
and U34467 (N_34467,N_33131,N_33006);
and U34468 (N_34468,N_33689,N_33476);
nand U34469 (N_34469,N_33070,N_33543);
and U34470 (N_34470,N_33148,N_33860);
or U34471 (N_34471,N_33258,N_33099);
nand U34472 (N_34472,N_33559,N_33674);
nand U34473 (N_34473,N_33337,N_33059);
or U34474 (N_34474,N_33314,N_33134);
and U34475 (N_34475,N_33779,N_33194);
or U34476 (N_34476,N_33702,N_33653);
nand U34477 (N_34477,N_33920,N_33016);
nor U34478 (N_34478,N_33095,N_33372);
or U34479 (N_34479,N_33601,N_33563);
nand U34480 (N_34480,N_33739,N_33130);
xnor U34481 (N_34481,N_33358,N_33839);
or U34482 (N_34482,N_33235,N_33422);
or U34483 (N_34483,N_33764,N_33208);
xor U34484 (N_34484,N_33700,N_33484);
xor U34485 (N_34485,N_33293,N_33467);
nor U34486 (N_34486,N_33491,N_33560);
nor U34487 (N_34487,N_33591,N_33585);
or U34488 (N_34488,N_33914,N_33383);
or U34489 (N_34489,N_33077,N_33928);
or U34490 (N_34490,N_33791,N_33154);
or U34491 (N_34491,N_33639,N_33590);
nand U34492 (N_34492,N_33298,N_33434);
nand U34493 (N_34493,N_33929,N_33829);
nand U34494 (N_34494,N_33843,N_33054);
or U34495 (N_34495,N_33236,N_33037);
or U34496 (N_34496,N_33901,N_33047);
nor U34497 (N_34497,N_33311,N_33930);
xor U34498 (N_34498,N_33855,N_33156);
and U34499 (N_34499,N_33183,N_33504);
nand U34500 (N_34500,N_33608,N_33859);
xnor U34501 (N_34501,N_33112,N_33134);
nor U34502 (N_34502,N_33474,N_33306);
xor U34503 (N_34503,N_33390,N_33101);
nor U34504 (N_34504,N_33819,N_33802);
or U34505 (N_34505,N_33325,N_33796);
nand U34506 (N_34506,N_33945,N_33853);
xnor U34507 (N_34507,N_33084,N_33654);
xnor U34508 (N_34508,N_33282,N_33158);
nor U34509 (N_34509,N_33975,N_33321);
nand U34510 (N_34510,N_33279,N_33039);
nor U34511 (N_34511,N_33365,N_33219);
xor U34512 (N_34512,N_33175,N_33803);
or U34513 (N_34513,N_33251,N_33398);
nand U34514 (N_34514,N_33319,N_33240);
nand U34515 (N_34515,N_33807,N_33744);
nor U34516 (N_34516,N_33047,N_33977);
nand U34517 (N_34517,N_33608,N_33095);
nor U34518 (N_34518,N_33705,N_33309);
xnor U34519 (N_34519,N_33502,N_33356);
and U34520 (N_34520,N_33893,N_33088);
xnor U34521 (N_34521,N_33090,N_33549);
xnor U34522 (N_34522,N_33119,N_33282);
and U34523 (N_34523,N_33744,N_33797);
xor U34524 (N_34524,N_33626,N_33349);
xnor U34525 (N_34525,N_33438,N_33911);
xnor U34526 (N_34526,N_33972,N_33660);
nand U34527 (N_34527,N_33635,N_33842);
xor U34528 (N_34528,N_33835,N_33390);
xor U34529 (N_34529,N_33252,N_33083);
xnor U34530 (N_34530,N_33539,N_33349);
nand U34531 (N_34531,N_33124,N_33849);
nor U34532 (N_34532,N_33496,N_33078);
and U34533 (N_34533,N_33366,N_33111);
or U34534 (N_34534,N_33311,N_33604);
or U34535 (N_34535,N_33096,N_33226);
nor U34536 (N_34536,N_33685,N_33700);
and U34537 (N_34537,N_33515,N_33610);
nand U34538 (N_34538,N_33109,N_33986);
and U34539 (N_34539,N_33870,N_33934);
and U34540 (N_34540,N_33725,N_33268);
and U34541 (N_34541,N_33882,N_33281);
and U34542 (N_34542,N_33091,N_33737);
xnor U34543 (N_34543,N_33411,N_33986);
and U34544 (N_34544,N_33290,N_33084);
nand U34545 (N_34545,N_33990,N_33892);
xnor U34546 (N_34546,N_33289,N_33088);
and U34547 (N_34547,N_33388,N_33132);
nor U34548 (N_34548,N_33143,N_33021);
xnor U34549 (N_34549,N_33464,N_33382);
and U34550 (N_34550,N_33743,N_33412);
xor U34551 (N_34551,N_33163,N_33160);
nor U34552 (N_34552,N_33677,N_33503);
and U34553 (N_34553,N_33831,N_33945);
xnor U34554 (N_34554,N_33330,N_33063);
nor U34555 (N_34555,N_33843,N_33763);
and U34556 (N_34556,N_33259,N_33447);
nor U34557 (N_34557,N_33891,N_33938);
xnor U34558 (N_34558,N_33814,N_33874);
nand U34559 (N_34559,N_33786,N_33096);
xor U34560 (N_34560,N_33743,N_33749);
and U34561 (N_34561,N_33684,N_33536);
and U34562 (N_34562,N_33999,N_33326);
or U34563 (N_34563,N_33130,N_33890);
nand U34564 (N_34564,N_33694,N_33240);
and U34565 (N_34565,N_33831,N_33703);
nor U34566 (N_34566,N_33062,N_33619);
xnor U34567 (N_34567,N_33065,N_33463);
or U34568 (N_34568,N_33225,N_33957);
nand U34569 (N_34569,N_33890,N_33494);
xnor U34570 (N_34570,N_33560,N_33106);
xor U34571 (N_34571,N_33700,N_33593);
nand U34572 (N_34572,N_33215,N_33473);
or U34573 (N_34573,N_33453,N_33660);
nor U34574 (N_34574,N_33311,N_33082);
xnor U34575 (N_34575,N_33184,N_33648);
or U34576 (N_34576,N_33878,N_33914);
xnor U34577 (N_34577,N_33709,N_33320);
nand U34578 (N_34578,N_33377,N_33968);
nor U34579 (N_34579,N_33161,N_33447);
or U34580 (N_34580,N_33417,N_33351);
and U34581 (N_34581,N_33199,N_33413);
nand U34582 (N_34582,N_33528,N_33879);
xor U34583 (N_34583,N_33520,N_33029);
nand U34584 (N_34584,N_33991,N_33088);
nor U34585 (N_34585,N_33004,N_33733);
or U34586 (N_34586,N_33418,N_33662);
nand U34587 (N_34587,N_33848,N_33271);
nand U34588 (N_34588,N_33706,N_33476);
xor U34589 (N_34589,N_33353,N_33679);
and U34590 (N_34590,N_33042,N_33713);
and U34591 (N_34591,N_33824,N_33140);
nand U34592 (N_34592,N_33807,N_33326);
and U34593 (N_34593,N_33566,N_33623);
nor U34594 (N_34594,N_33353,N_33789);
and U34595 (N_34595,N_33897,N_33437);
and U34596 (N_34596,N_33366,N_33495);
nor U34597 (N_34597,N_33059,N_33792);
or U34598 (N_34598,N_33989,N_33456);
nand U34599 (N_34599,N_33847,N_33996);
nor U34600 (N_34600,N_33133,N_33417);
xnor U34601 (N_34601,N_33526,N_33474);
and U34602 (N_34602,N_33126,N_33749);
nand U34603 (N_34603,N_33879,N_33920);
nor U34604 (N_34604,N_33757,N_33426);
nor U34605 (N_34605,N_33340,N_33116);
nand U34606 (N_34606,N_33114,N_33384);
nand U34607 (N_34607,N_33866,N_33633);
or U34608 (N_34608,N_33400,N_33618);
nand U34609 (N_34609,N_33776,N_33685);
or U34610 (N_34610,N_33826,N_33980);
nand U34611 (N_34611,N_33885,N_33931);
and U34612 (N_34612,N_33991,N_33227);
nand U34613 (N_34613,N_33375,N_33573);
xor U34614 (N_34614,N_33781,N_33608);
nand U34615 (N_34615,N_33699,N_33797);
or U34616 (N_34616,N_33518,N_33234);
nor U34617 (N_34617,N_33209,N_33084);
nand U34618 (N_34618,N_33775,N_33304);
nor U34619 (N_34619,N_33310,N_33631);
and U34620 (N_34620,N_33249,N_33010);
and U34621 (N_34621,N_33326,N_33134);
nor U34622 (N_34622,N_33729,N_33012);
nand U34623 (N_34623,N_33937,N_33705);
nand U34624 (N_34624,N_33615,N_33165);
nand U34625 (N_34625,N_33803,N_33685);
and U34626 (N_34626,N_33814,N_33917);
nor U34627 (N_34627,N_33543,N_33423);
and U34628 (N_34628,N_33350,N_33275);
nor U34629 (N_34629,N_33189,N_33172);
nor U34630 (N_34630,N_33545,N_33741);
nor U34631 (N_34631,N_33384,N_33711);
nand U34632 (N_34632,N_33482,N_33081);
nor U34633 (N_34633,N_33797,N_33333);
nor U34634 (N_34634,N_33927,N_33693);
xor U34635 (N_34635,N_33674,N_33726);
or U34636 (N_34636,N_33837,N_33796);
xor U34637 (N_34637,N_33401,N_33623);
and U34638 (N_34638,N_33062,N_33262);
or U34639 (N_34639,N_33546,N_33861);
and U34640 (N_34640,N_33733,N_33097);
nand U34641 (N_34641,N_33117,N_33597);
or U34642 (N_34642,N_33151,N_33892);
or U34643 (N_34643,N_33104,N_33738);
and U34644 (N_34644,N_33100,N_33243);
and U34645 (N_34645,N_33687,N_33265);
and U34646 (N_34646,N_33286,N_33291);
or U34647 (N_34647,N_33283,N_33069);
nand U34648 (N_34648,N_33265,N_33904);
and U34649 (N_34649,N_33421,N_33042);
and U34650 (N_34650,N_33518,N_33306);
xnor U34651 (N_34651,N_33537,N_33449);
nor U34652 (N_34652,N_33993,N_33891);
and U34653 (N_34653,N_33151,N_33258);
nand U34654 (N_34654,N_33593,N_33327);
xor U34655 (N_34655,N_33328,N_33852);
xor U34656 (N_34656,N_33808,N_33051);
or U34657 (N_34657,N_33392,N_33998);
nor U34658 (N_34658,N_33483,N_33275);
and U34659 (N_34659,N_33749,N_33805);
and U34660 (N_34660,N_33026,N_33532);
nand U34661 (N_34661,N_33552,N_33058);
nor U34662 (N_34662,N_33969,N_33508);
xnor U34663 (N_34663,N_33373,N_33530);
and U34664 (N_34664,N_33957,N_33884);
nand U34665 (N_34665,N_33143,N_33389);
and U34666 (N_34666,N_33834,N_33120);
nor U34667 (N_34667,N_33157,N_33761);
and U34668 (N_34668,N_33977,N_33252);
nand U34669 (N_34669,N_33089,N_33256);
or U34670 (N_34670,N_33266,N_33759);
nand U34671 (N_34671,N_33484,N_33735);
nand U34672 (N_34672,N_33940,N_33299);
or U34673 (N_34673,N_33038,N_33562);
xnor U34674 (N_34674,N_33739,N_33000);
nor U34675 (N_34675,N_33648,N_33209);
and U34676 (N_34676,N_33814,N_33435);
or U34677 (N_34677,N_33522,N_33165);
nor U34678 (N_34678,N_33148,N_33433);
or U34679 (N_34679,N_33551,N_33936);
nor U34680 (N_34680,N_33196,N_33054);
and U34681 (N_34681,N_33793,N_33909);
nand U34682 (N_34682,N_33983,N_33722);
and U34683 (N_34683,N_33747,N_33598);
or U34684 (N_34684,N_33551,N_33154);
nand U34685 (N_34685,N_33113,N_33787);
and U34686 (N_34686,N_33395,N_33439);
and U34687 (N_34687,N_33869,N_33562);
and U34688 (N_34688,N_33308,N_33517);
and U34689 (N_34689,N_33538,N_33208);
and U34690 (N_34690,N_33226,N_33189);
and U34691 (N_34691,N_33213,N_33454);
or U34692 (N_34692,N_33173,N_33085);
nand U34693 (N_34693,N_33326,N_33933);
nand U34694 (N_34694,N_33923,N_33818);
xor U34695 (N_34695,N_33271,N_33721);
xor U34696 (N_34696,N_33766,N_33307);
nand U34697 (N_34697,N_33062,N_33171);
xnor U34698 (N_34698,N_33382,N_33970);
nor U34699 (N_34699,N_33378,N_33285);
or U34700 (N_34700,N_33052,N_33525);
nor U34701 (N_34701,N_33901,N_33672);
and U34702 (N_34702,N_33361,N_33040);
and U34703 (N_34703,N_33595,N_33408);
nand U34704 (N_34704,N_33988,N_33188);
xnor U34705 (N_34705,N_33929,N_33767);
nor U34706 (N_34706,N_33581,N_33856);
or U34707 (N_34707,N_33502,N_33908);
nand U34708 (N_34708,N_33113,N_33259);
nor U34709 (N_34709,N_33295,N_33946);
xnor U34710 (N_34710,N_33383,N_33879);
and U34711 (N_34711,N_33191,N_33325);
or U34712 (N_34712,N_33520,N_33618);
xnor U34713 (N_34713,N_33379,N_33069);
xor U34714 (N_34714,N_33478,N_33610);
or U34715 (N_34715,N_33729,N_33687);
xor U34716 (N_34716,N_33070,N_33443);
xor U34717 (N_34717,N_33719,N_33515);
xor U34718 (N_34718,N_33621,N_33522);
nand U34719 (N_34719,N_33739,N_33400);
xor U34720 (N_34720,N_33940,N_33564);
or U34721 (N_34721,N_33421,N_33099);
nor U34722 (N_34722,N_33750,N_33726);
nor U34723 (N_34723,N_33060,N_33722);
nand U34724 (N_34724,N_33919,N_33695);
nor U34725 (N_34725,N_33114,N_33434);
xor U34726 (N_34726,N_33647,N_33852);
xor U34727 (N_34727,N_33574,N_33381);
and U34728 (N_34728,N_33730,N_33387);
or U34729 (N_34729,N_33228,N_33715);
xor U34730 (N_34730,N_33035,N_33886);
or U34731 (N_34731,N_33995,N_33913);
nand U34732 (N_34732,N_33209,N_33902);
and U34733 (N_34733,N_33618,N_33037);
nand U34734 (N_34734,N_33856,N_33181);
nand U34735 (N_34735,N_33672,N_33791);
and U34736 (N_34736,N_33335,N_33191);
nor U34737 (N_34737,N_33065,N_33745);
or U34738 (N_34738,N_33103,N_33515);
nand U34739 (N_34739,N_33105,N_33900);
or U34740 (N_34740,N_33993,N_33784);
xor U34741 (N_34741,N_33864,N_33306);
xor U34742 (N_34742,N_33333,N_33459);
or U34743 (N_34743,N_33721,N_33486);
xor U34744 (N_34744,N_33343,N_33256);
xor U34745 (N_34745,N_33387,N_33538);
or U34746 (N_34746,N_33339,N_33272);
xor U34747 (N_34747,N_33223,N_33534);
nor U34748 (N_34748,N_33245,N_33552);
and U34749 (N_34749,N_33077,N_33459);
or U34750 (N_34750,N_33645,N_33863);
nand U34751 (N_34751,N_33880,N_33537);
nand U34752 (N_34752,N_33506,N_33824);
nand U34753 (N_34753,N_33138,N_33990);
and U34754 (N_34754,N_33265,N_33913);
xnor U34755 (N_34755,N_33678,N_33607);
xnor U34756 (N_34756,N_33097,N_33786);
nor U34757 (N_34757,N_33083,N_33156);
nand U34758 (N_34758,N_33758,N_33491);
xor U34759 (N_34759,N_33789,N_33990);
and U34760 (N_34760,N_33641,N_33702);
xnor U34761 (N_34761,N_33581,N_33645);
nor U34762 (N_34762,N_33981,N_33744);
or U34763 (N_34763,N_33109,N_33279);
xor U34764 (N_34764,N_33145,N_33249);
xnor U34765 (N_34765,N_33372,N_33505);
nand U34766 (N_34766,N_33131,N_33604);
nor U34767 (N_34767,N_33106,N_33145);
nor U34768 (N_34768,N_33867,N_33383);
xnor U34769 (N_34769,N_33832,N_33628);
nand U34770 (N_34770,N_33619,N_33796);
xor U34771 (N_34771,N_33323,N_33820);
nor U34772 (N_34772,N_33657,N_33214);
xnor U34773 (N_34773,N_33861,N_33483);
xnor U34774 (N_34774,N_33779,N_33053);
nor U34775 (N_34775,N_33019,N_33618);
or U34776 (N_34776,N_33882,N_33279);
or U34777 (N_34777,N_33607,N_33245);
xor U34778 (N_34778,N_33582,N_33672);
nand U34779 (N_34779,N_33488,N_33126);
and U34780 (N_34780,N_33412,N_33374);
and U34781 (N_34781,N_33727,N_33366);
and U34782 (N_34782,N_33644,N_33759);
nor U34783 (N_34783,N_33430,N_33316);
nand U34784 (N_34784,N_33479,N_33378);
or U34785 (N_34785,N_33658,N_33324);
nand U34786 (N_34786,N_33095,N_33911);
and U34787 (N_34787,N_33575,N_33034);
nand U34788 (N_34788,N_33157,N_33160);
xor U34789 (N_34789,N_33338,N_33221);
xnor U34790 (N_34790,N_33441,N_33885);
nand U34791 (N_34791,N_33661,N_33505);
or U34792 (N_34792,N_33142,N_33850);
or U34793 (N_34793,N_33323,N_33552);
and U34794 (N_34794,N_33962,N_33994);
nor U34795 (N_34795,N_33164,N_33378);
or U34796 (N_34796,N_33477,N_33457);
nor U34797 (N_34797,N_33170,N_33148);
nand U34798 (N_34798,N_33855,N_33814);
or U34799 (N_34799,N_33792,N_33351);
nand U34800 (N_34800,N_33964,N_33290);
or U34801 (N_34801,N_33813,N_33704);
and U34802 (N_34802,N_33462,N_33934);
and U34803 (N_34803,N_33248,N_33757);
nand U34804 (N_34804,N_33437,N_33551);
and U34805 (N_34805,N_33711,N_33235);
and U34806 (N_34806,N_33681,N_33564);
nand U34807 (N_34807,N_33469,N_33920);
nand U34808 (N_34808,N_33453,N_33518);
nor U34809 (N_34809,N_33233,N_33732);
xnor U34810 (N_34810,N_33917,N_33647);
nand U34811 (N_34811,N_33967,N_33266);
or U34812 (N_34812,N_33469,N_33768);
or U34813 (N_34813,N_33075,N_33068);
or U34814 (N_34814,N_33624,N_33440);
or U34815 (N_34815,N_33666,N_33048);
xnor U34816 (N_34816,N_33092,N_33340);
and U34817 (N_34817,N_33218,N_33213);
nand U34818 (N_34818,N_33247,N_33088);
nand U34819 (N_34819,N_33173,N_33226);
nand U34820 (N_34820,N_33474,N_33377);
and U34821 (N_34821,N_33916,N_33088);
nor U34822 (N_34822,N_33044,N_33740);
nor U34823 (N_34823,N_33088,N_33212);
or U34824 (N_34824,N_33987,N_33486);
or U34825 (N_34825,N_33199,N_33352);
nor U34826 (N_34826,N_33008,N_33467);
and U34827 (N_34827,N_33459,N_33738);
xnor U34828 (N_34828,N_33438,N_33218);
or U34829 (N_34829,N_33944,N_33033);
xnor U34830 (N_34830,N_33286,N_33391);
and U34831 (N_34831,N_33180,N_33375);
or U34832 (N_34832,N_33703,N_33545);
or U34833 (N_34833,N_33546,N_33521);
or U34834 (N_34834,N_33762,N_33073);
nor U34835 (N_34835,N_33521,N_33124);
nand U34836 (N_34836,N_33996,N_33567);
xnor U34837 (N_34837,N_33742,N_33236);
nand U34838 (N_34838,N_33716,N_33538);
and U34839 (N_34839,N_33207,N_33782);
nor U34840 (N_34840,N_33579,N_33742);
nand U34841 (N_34841,N_33040,N_33467);
nor U34842 (N_34842,N_33055,N_33900);
or U34843 (N_34843,N_33219,N_33777);
xor U34844 (N_34844,N_33095,N_33301);
xnor U34845 (N_34845,N_33619,N_33325);
and U34846 (N_34846,N_33962,N_33366);
or U34847 (N_34847,N_33113,N_33409);
or U34848 (N_34848,N_33478,N_33550);
and U34849 (N_34849,N_33982,N_33510);
nand U34850 (N_34850,N_33411,N_33560);
and U34851 (N_34851,N_33849,N_33074);
nor U34852 (N_34852,N_33722,N_33253);
or U34853 (N_34853,N_33672,N_33490);
and U34854 (N_34854,N_33336,N_33109);
nand U34855 (N_34855,N_33377,N_33655);
nand U34856 (N_34856,N_33017,N_33984);
nand U34857 (N_34857,N_33006,N_33969);
and U34858 (N_34858,N_33006,N_33279);
nand U34859 (N_34859,N_33947,N_33225);
nor U34860 (N_34860,N_33669,N_33550);
xor U34861 (N_34861,N_33641,N_33074);
nor U34862 (N_34862,N_33148,N_33239);
or U34863 (N_34863,N_33428,N_33862);
nor U34864 (N_34864,N_33398,N_33766);
nand U34865 (N_34865,N_33423,N_33997);
nor U34866 (N_34866,N_33762,N_33685);
xnor U34867 (N_34867,N_33669,N_33259);
nor U34868 (N_34868,N_33349,N_33680);
and U34869 (N_34869,N_33364,N_33775);
xor U34870 (N_34870,N_33197,N_33216);
and U34871 (N_34871,N_33004,N_33488);
xor U34872 (N_34872,N_33151,N_33389);
and U34873 (N_34873,N_33554,N_33255);
xor U34874 (N_34874,N_33223,N_33656);
and U34875 (N_34875,N_33702,N_33087);
or U34876 (N_34876,N_33313,N_33012);
xnor U34877 (N_34877,N_33691,N_33288);
and U34878 (N_34878,N_33823,N_33096);
nand U34879 (N_34879,N_33359,N_33289);
nand U34880 (N_34880,N_33955,N_33068);
nand U34881 (N_34881,N_33527,N_33831);
or U34882 (N_34882,N_33746,N_33991);
nand U34883 (N_34883,N_33672,N_33688);
nand U34884 (N_34884,N_33851,N_33463);
and U34885 (N_34885,N_33284,N_33803);
and U34886 (N_34886,N_33634,N_33225);
or U34887 (N_34887,N_33720,N_33236);
nand U34888 (N_34888,N_33729,N_33188);
nor U34889 (N_34889,N_33163,N_33857);
nand U34890 (N_34890,N_33789,N_33863);
and U34891 (N_34891,N_33842,N_33769);
nor U34892 (N_34892,N_33003,N_33215);
xnor U34893 (N_34893,N_33826,N_33512);
or U34894 (N_34894,N_33771,N_33818);
and U34895 (N_34895,N_33596,N_33384);
nor U34896 (N_34896,N_33327,N_33330);
or U34897 (N_34897,N_33287,N_33782);
nor U34898 (N_34898,N_33095,N_33912);
nand U34899 (N_34899,N_33153,N_33437);
nand U34900 (N_34900,N_33404,N_33175);
or U34901 (N_34901,N_33201,N_33178);
nor U34902 (N_34902,N_33398,N_33465);
xnor U34903 (N_34903,N_33055,N_33764);
nor U34904 (N_34904,N_33447,N_33745);
and U34905 (N_34905,N_33676,N_33179);
and U34906 (N_34906,N_33552,N_33010);
nor U34907 (N_34907,N_33682,N_33344);
or U34908 (N_34908,N_33920,N_33407);
or U34909 (N_34909,N_33356,N_33122);
or U34910 (N_34910,N_33227,N_33680);
and U34911 (N_34911,N_33177,N_33861);
xor U34912 (N_34912,N_33404,N_33636);
nand U34913 (N_34913,N_33447,N_33373);
and U34914 (N_34914,N_33563,N_33676);
nor U34915 (N_34915,N_33957,N_33341);
xor U34916 (N_34916,N_33487,N_33746);
or U34917 (N_34917,N_33392,N_33619);
or U34918 (N_34918,N_33307,N_33314);
and U34919 (N_34919,N_33024,N_33666);
and U34920 (N_34920,N_33265,N_33600);
nor U34921 (N_34921,N_33504,N_33844);
or U34922 (N_34922,N_33157,N_33999);
xor U34923 (N_34923,N_33780,N_33096);
nand U34924 (N_34924,N_33455,N_33591);
or U34925 (N_34925,N_33385,N_33412);
or U34926 (N_34926,N_33402,N_33057);
xor U34927 (N_34927,N_33948,N_33239);
nand U34928 (N_34928,N_33259,N_33825);
and U34929 (N_34929,N_33720,N_33274);
nand U34930 (N_34930,N_33030,N_33288);
xnor U34931 (N_34931,N_33291,N_33822);
or U34932 (N_34932,N_33554,N_33166);
xnor U34933 (N_34933,N_33233,N_33604);
nand U34934 (N_34934,N_33320,N_33045);
and U34935 (N_34935,N_33089,N_33001);
or U34936 (N_34936,N_33990,N_33452);
nor U34937 (N_34937,N_33734,N_33350);
nand U34938 (N_34938,N_33030,N_33668);
or U34939 (N_34939,N_33170,N_33090);
nand U34940 (N_34940,N_33635,N_33096);
and U34941 (N_34941,N_33373,N_33888);
xor U34942 (N_34942,N_33335,N_33947);
nand U34943 (N_34943,N_33668,N_33361);
nor U34944 (N_34944,N_33689,N_33446);
nor U34945 (N_34945,N_33769,N_33608);
xor U34946 (N_34946,N_33193,N_33693);
nand U34947 (N_34947,N_33568,N_33882);
xnor U34948 (N_34948,N_33836,N_33917);
and U34949 (N_34949,N_33807,N_33932);
nand U34950 (N_34950,N_33319,N_33432);
nor U34951 (N_34951,N_33076,N_33643);
nand U34952 (N_34952,N_33814,N_33207);
xnor U34953 (N_34953,N_33688,N_33608);
nand U34954 (N_34954,N_33541,N_33345);
nand U34955 (N_34955,N_33180,N_33721);
and U34956 (N_34956,N_33805,N_33599);
nor U34957 (N_34957,N_33925,N_33420);
nor U34958 (N_34958,N_33409,N_33120);
nor U34959 (N_34959,N_33212,N_33577);
or U34960 (N_34960,N_33708,N_33159);
and U34961 (N_34961,N_33749,N_33379);
nand U34962 (N_34962,N_33518,N_33674);
nand U34963 (N_34963,N_33656,N_33933);
nand U34964 (N_34964,N_33049,N_33439);
nor U34965 (N_34965,N_33130,N_33935);
nand U34966 (N_34966,N_33259,N_33322);
nor U34967 (N_34967,N_33860,N_33588);
and U34968 (N_34968,N_33848,N_33684);
xnor U34969 (N_34969,N_33403,N_33285);
xnor U34970 (N_34970,N_33439,N_33886);
xor U34971 (N_34971,N_33819,N_33921);
and U34972 (N_34972,N_33419,N_33422);
nor U34973 (N_34973,N_33394,N_33913);
or U34974 (N_34974,N_33265,N_33819);
or U34975 (N_34975,N_33344,N_33007);
nor U34976 (N_34976,N_33163,N_33545);
nand U34977 (N_34977,N_33979,N_33242);
and U34978 (N_34978,N_33906,N_33175);
nor U34979 (N_34979,N_33074,N_33229);
or U34980 (N_34980,N_33287,N_33205);
nor U34981 (N_34981,N_33287,N_33711);
nor U34982 (N_34982,N_33902,N_33115);
or U34983 (N_34983,N_33179,N_33823);
or U34984 (N_34984,N_33665,N_33852);
or U34985 (N_34985,N_33066,N_33459);
or U34986 (N_34986,N_33529,N_33396);
or U34987 (N_34987,N_33236,N_33521);
and U34988 (N_34988,N_33710,N_33588);
nand U34989 (N_34989,N_33751,N_33458);
or U34990 (N_34990,N_33763,N_33250);
nand U34991 (N_34991,N_33023,N_33556);
nor U34992 (N_34992,N_33284,N_33766);
and U34993 (N_34993,N_33590,N_33694);
nor U34994 (N_34994,N_33290,N_33799);
and U34995 (N_34995,N_33002,N_33191);
and U34996 (N_34996,N_33330,N_33280);
nor U34997 (N_34997,N_33528,N_33414);
or U34998 (N_34998,N_33984,N_33382);
xor U34999 (N_34999,N_33290,N_33762);
or U35000 (N_35000,N_34940,N_34144);
and U35001 (N_35001,N_34229,N_34002);
or U35002 (N_35002,N_34559,N_34181);
xnor U35003 (N_35003,N_34998,N_34233);
nand U35004 (N_35004,N_34049,N_34072);
and U35005 (N_35005,N_34914,N_34352);
nor U35006 (N_35006,N_34869,N_34619);
xor U35007 (N_35007,N_34259,N_34032);
xnor U35008 (N_35008,N_34408,N_34857);
and U35009 (N_35009,N_34560,N_34839);
and U35010 (N_35010,N_34491,N_34167);
xnor U35011 (N_35011,N_34249,N_34178);
nor U35012 (N_35012,N_34396,N_34689);
nor U35013 (N_35013,N_34083,N_34936);
and U35014 (N_35014,N_34846,N_34084);
and U35015 (N_35015,N_34412,N_34247);
or U35016 (N_35016,N_34526,N_34082);
or U35017 (N_35017,N_34294,N_34046);
and U35018 (N_35018,N_34146,N_34785);
nand U35019 (N_35019,N_34653,N_34777);
nor U35020 (N_35020,N_34636,N_34720);
nor U35021 (N_35021,N_34217,N_34342);
nor U35022 (N_35022,N_34005,N_34363);
xor U35023 (N_35023,N_34867,N_34456);
nand U35024 (N_35024,N_34351,N_34537);
and U35025 (N_35025,N_34614,N_34199);
or U35026 (N_35026,N_34933,N_34077);
nand U35027 (N_35027,N_34708,N_34542);
and U35028 (N_35028,N_34573,N_34316);
xor U35029 (N_35029,N_34011,N_34528);
nor U35030 (N_35030,N_34039,N_34382);
nor U35031 (N_35031,N_34643,N_34944);
and U35032 (N_35032,N_34424,N_34935);
or U35033 (N_35033,N_34320,N_34808);
and U35034 (N_35034,N_34538,N_34333);
nor U35035 (N_35035,N_34618,N_34563);
or U35036 (N_35036,N_34079,N_34306);
nor U35037 (N_35037,N_34864,N_34865);
and U35038 (N_35038,N_34147,N_34702);
and U35039 (N_35039,N_34277,N_34120);
or U35040 (N_35040,N_34763,N_34773);
or U35041 (N_35041,N_34851,N_34089);
or U35042 (N_35042,N_34654,N_34647);
or U35043 (N_35043,N_34623,N_34286);
nor U35044 (N_35044,N_34327,N_34965);
or U35045 (N_35045,N_34218,N_34238);
and U35046 (N_35046,N_34176,N_34004);
or U35047 (N_35047,N_34122,N_34261);
nand U35048 (N_35048,N_34161,N_34367);
nor U35049 (N_35049,N_34956,N_34904);
and U35050 (N_35050,N_34473,N_34972);
xor U35051 (N_35051,N_34855,N_34250);
nand U35052 (N_35052,N_34493,N_34097);
and U35053 (N_35053,N_34264,N_34335);
nand U35054 (N_35054,N_34530,N_34600);
nand U35055 (N_35055,N_34822,N_34738);
nor U35056 (N_35056,N_34877,N_34686);
nor U35057 (N_35057,N_34805,N_34765);
or U35058 (N_35058,N_34453,N_34583);
nor U35059 (N_35059,N_34760,N_34649);
xor U35060 (N_35060,N_34449,N_34389);
and U35061 (N_35061,N_34801,N_34878);
and U35062 (N_35062,N_34260,N_34546);
nand U35063 (N_35063,N_34321,N_34958);
xor U35064 (N_35064,N_34251,N_34479);
or U35065 (N_35065,N_34613,N_34932);
or U35066 (N_35066,N_34786,N_34273);
nor U35067 (N_35067,N_34244,N_34793);
and U35068 (N_35068,N_34691,N_34658);
or U35069 (N_35069,N_34927,N_34910);
xor U35070 (N_35070,N_34215,N_34754);
nor U35071 (N_35071,N_34432,N_34138);
nor U35072 (N_35072,N_34481,N_34888);
nand U35073 (N_35073,N_34924,N_34863);
nand U35074 (N_35074,N_34985,N_34565);
xor U35075 (N_35075,N_34687,N_34459);
nor U35076 (N_35076,N_34336,N_34207);
and U35077 (N_35077,N_34024,N_34885);
or U35078 (N_35078,N_34744,N_34671);
or U35079 (N_35079,N_34219,N_34392);
nand U35080 (N_35080,N_34081,N_34285);
nand U35081 (N_35081,N_34640,N_34446);
nor U35082 (N_35082,N_34920,N_34506);
and U35083 (N_35083,N_34007,N_34676);
or U35084 (N_35084,N_34873,N_34798);
nor U35085 (N_35085,N_34715,N_34678);
and U35086 (N_35086,N_34823,N_34299);
and U35087 (N_35087,N_34444,N_34633);
and U35088 (N_35088,N_34159,N_34609);
xor U35089 (N_35089,N_34736,N_34922);
nor U35090 (N_35090,N_34369,N_34796);
nand U35091 (N_35091,N_34111,N_34488);
xor U35092 (N_35092,N_34997,N_34588);
nor U35093 (N_35093,N_34045,N_34853);
or U35094 (N_35094,N_34228,N_34467);
and U35095 (N_35095,N_34917,N_34787);
and U35096 (N_35096,N_34463,N_34641);
xor U35097 (N_35097,N_34733,N_34766);
xor U35098 (N_35098,N_34764,N_34364);
nor U35099 (N_35099,N_34982,N_34790);
or U35100 (N_35100,N_34312,N_34026);
or U35101 (N_35101,N_34248,N_34431);
and U35102 (N_35102,N_34890,N_34582);
nor U35103 (N_35103,N_34554,N_34757);
nor U35104 (N_35104,N_34393,N_34443);
nand U35105 (N_35105,N_34242,N_34208);
xnor U35106 (N_35106,N_34806,N_34398);
and U35107 (N_35107,N_34862,N_34202);
xnor U35108 (N_35108,N_34502,N_34307);
xnor U35109 (N_35109,N_34988,N_34127);
nor U35110 (N_35110,N_34115,N_34001);
nand U35111 (N_35111,N_34939,N_34612);
nor U35112 (N_35112,N_34664,N_34071);
nor U35113 (N_35113,N_34732,N_34267);
and U35114 (N_35114,N_34572,N_34717);
xnor U35115 (N_35115,N_34707,N_34519);
xor U35116 (N_35116,N_34418,N_34714);
nor U35117 (N_35117,N_34523,N_34774);
xor U35118 (N_35118,N_34838,N_34213);
nor U35119 (N_35119,N_34941,N_34751);
and U35120 (N_35120,N_34227,N_34015);
nor U35121 (N_35121,N_34813,N_34953);
nor U35122 (N_35122,N_34378,N_34597);
nand U35123 (N_35123,N_34254,N_34324);
or U35124 (N_35124,N_34980,N_34870);
xnor U35125 (N_35125,N_34628,N_34986);
nor U35126 (N_35126,N_34427,N_34454);
nor U35127 (N_35127,N_34126,N_34395);
nor U35128 (N_35128,N_34517,N_34828);
and U35129 (N_35129,N_34076,N_34946);
and U35130 (N_35130,N_34522,N_34420);
or U35131 (N_35131,N_34718,N_34200);
or U35132 (N_35132,N_34727,N_34646);
nor U35133 (N_35133,N_34346,N_34644);
and U35134 (N_35134,N_34778,N_34203);
or U35135 (N_35135,N_34938,N_34314);
xnor U35136 (N_35136,N_34648,N_34610);
and U35137 (N_35137,N_34365,N_34655);
and U35138 (N_35138,N_34487,N_34353);
and U35139 (N_35139,N_34101,N_34128);
nor U35140 (N_35140,N_34087,N_34376);
nand U35141 (N_35141,N_34317,N_34848);
xor U35142 (N_35142,N_34734,N_34153);
and U35143 (N_35143,N_34674,N_34627);
nor U35144 (N_35144,N_34402,N_34595);
and U35145 (N_35145,N_34281,N_34679);
nor U35146 (N_35146,N_34657,N_34818);
nor U35147 (N_35147,N_34992,N_34241);
nand U35148 (N_35148,N_34670,N_34761);
nor U35149 (N_35149,N_34345,N_34704);
nand U35150 (N_35150,N_34113,N_34182);
xor U35151 (N_35151,N_34970,N_34685);
xor U35152 (N_35152,N_34021,N_34053);
nor U35153 (N_35153,N_34952,N_34239);
xnor U35154 (N_35154,N_34322,N_34293);
and U35155 (N_35155,N_34268,N_34103);
or U35156 (N_35156,N_34589,N_34692);
nand U35157 (N_35157,N_34812,N_34780);
nand U35158 (N_35158,N_34520,N_34503);
or U35159 (N_35159,N_34169,N_34642);
nand U35160 (N_35160,N_34879,N_34561);
xor U35161 (N_35161,N_34586,N_34634);
xor U35162 (N_35162,N_34132,N_34043);
and U35163 (N_35163,N_34031,N_34544);
xnor U35164 (N_35164,N_34051,N_34577);
or U35165 (N_35165,N_34852,N_34820);
nor U35166 (N_35166,N_34065,N_34223);
xnor U35167 (N_35167,N_34849,N_34912);
nor U35168 (N_35168,N_34310,N_34606);
or U35169 (N_35169,N_34137,N_34656);
xnor U35170 (N_35170,N_34745,N_34383);
nand U35171 (N_35171,N_34133,N_34694);
nor U35172 (N_35172,N_34050,N_34090);
nor U35173 (N_35173,N_34070,N_34105);
or U35174 (N_35174,N_34550,N_34964);
or U35175 (N_35175,N_34458,N_34168);
nand U35176 (N_35176,N_34188,N_34357);
nand U35177 (N_35177,N_34447,N_34541);
nor U35178 (N_35178,N_34698,N_34252);
xnor U35179 (N_35179,N_34638,N_34226);
xnor U35180 (N_35180,N_34684,N_34832);
xor U35181 (N_35181,N_34926,N_34729);
nor U35182 (N_35182,N_34255,N_34621);
nand U35183 (N_35183,N_34696,N_34602);
nand U35184 (N_35184,N_34305,N_34834);
nor U35185 (N_35185,N_34950,N_34377);
nor U35186 (N_35186,N_34154,N_34018);
nor U35187 (N_35187,N_34478,N_34349);
xor U35188 (N_35188,N_34150,N_34999);
and U35189 (N_35189,N_34419,N_34866);
or U35190 (N_35190,N_34934,N_34104);
or U35191 (N_35191,N_34022,N_34123);
and U35192 (N_35192,N_34788,N_34211);
and U35193 (N_35193,N_34880,N_34074);
and U35194 (N_35194,N_34085,N_34854);
nand U35195 (N_35195,N_34220,N_34030);
or U35196 (N_35196,N_34850,N_34124);
xor U35197 (N_35197,N_34500,N_34996);
or U35198 (N_35198,N_34406,N_34152);
xor U35199 (N_35199,N_34884,N_34682);
nand U35200 (N_35200,N_34501,N_34978);
xnor U35201 (N_35201,N_34983,N_34824);
nor U35202 (N_35202,N_34624,N_34792);
nand U35203 (N_35203,N_34882,N_34945);
nand U35204 (N_35204,N_34348,N_34416);
nand U35205 (N_35205,N_34375,N_34433);
xor U35206 (N_35206,N_34163,N_34555);
nand U35207 (N_35207,N_34338,N_34274);
nand U35208 (N_35208,N_34987,N_34186);
nand U35209 (N_35209,N_34632,N_34693);
nand U35210 (N_35210,N_34789,N_34170);
and U35211 (N_35211,N_34652,N_34499);
or U35212 (N_35212,N_34579,N_34210);
xor U35213 (N_35213,N_34302,N_34270);
nor U35214 (N_35214,N_34843,N_34323);
xnor U35215 (N_35215,N_34174,N_34460);
xnor U35216 (N_35216,N_34037,N_34486);
and U35217 (N_35217,N_34075,N_34112);
nor U35218 (N_35218,N_34771,N_34325);
and U35219 (N_35219,N_34189,N_34906);
nor U35220 (N_35220,N_34810,N_34334);
xnor U35221 (N_35221,N_34562,N_34054);
nor U35222 (N_35222,N_34058,N_34234);
or U35223 (N_35223,N_34620,N_34009);
and U35224 (N_35224,N_34036,N_34651);
nor U35225 (N_35225,N_34359,N_34581);
or U35226 (N_35226,N_34521,N_34728);
or U35227 (N_35227,N_34216,N_34557);
nand U35228 (N_35228,N_34288,N_34355);
and U35229 (N_35229,N_34148,N_34574);
nand U35230 (N_35230,N_34826,N_34536);
xnor U35231 (N_35231,N_34504,N_34006);
or U35232 (N_35232,N_34979,N_34162);
or U35233 (N_35233,N_34552,N_34272);
nor U35234 (N_35234,N_34308,N_34430);
and U35235 (N_35235,N_34096,N_34875);
xnor U35236 (N_35236,N_34731,N_34911);
xnor U35237 (N_35237,N_34008,N_34571);
and U35238 (N_35238,N_34937,N_34175);
and U35239 (N_35239,N_34508,N_34918);
nand U35240 (N_35240,N_34598,N_34010);
nor U35241 (N_35241,N_34516,N_34889);
nand U35242 (N_35242,N_34116,N_34165);
nor U35243 (N_35243,N_34991,N_34014);
or U35244 (N_35244,N_34587,N_34399);
or U35245 (N_35245,N_34844,N_34253);
xnor U35246 (N_35246,N_34100,N_34591);
xnor U35247 (N_35247,N_34360,N_34019);
xor U35248 (N_35248,N_34237,N_34845);
xnor U35249 (N_35249,N_34568,N_34388);
nand U35250 (N_35250,N_34118,N_34971);
and U35251 (N_35251,N_34056,N_34151);
xnor U35252 (N_35252,N_34358,N_34131);
nand U35253 (N_35253,N_34746,N_34993);
or U35254 (N_35254,N_34140,N_34361);
xor U35255 (N_35255,N_34027,N_34578);
nor U35256 (N_35256,N_34240,N_34584);
and U35257 (N_35257,N_34477,N_34129);
and U35258 (N_35258,N_34301,N_34821);
nand U35259 (N_35259,N_34404,N_34114);
and U35260 (N_35260,N_34830,N_34759);
nor U35261 (N_35261,N_34222,N_34603);
nand U35262 (N_35262,N_34794,N_34437);
nor U35263 (N_35263,N_34068,N_34608);
nor U35264 (N_35264,N_34062,N_34825);
nand U35265 (N_35265,N_34723,N_34527);
nor U35266 (N_35266,N_34016,N_34775);
or U35267 (N_35267,N_34748,N_34829);
nand U35268 (N_35268,N_34663,N_34896);
nor U35269 (N_35269,N_34407,N_34130);
and U35270 (N_35270,N_34119,N_34566);
nand U35271 (N_35271,N_34902,N_34883);
and U35272 (N_35272,N_34059,N_34145);
and U35273 (N_35273,N_34086,N_34332);
or U35274 (N_35274,N_34758,N_34108);
or U35275 (N_35275,N_34680,N_34413);
or U35276 (N_35276,N_34340,N_34534);
and U35277 (N_35277,N_34576,N_34747);
and U35278 (N_35278,N_34683,N_34204);
nand U35279 (N_35279,N_34331,N_34468);
nand U35280 (N_35280,N_34035,N_34384);
or U35281 (N_35281,N_34549,N_34650);
and U35282 (N_35282,N_34512,N_34923);
xor U35283 (N_35283,N_34954,N_34209);
or U35284 (N_35284,N_34817,N_34374);
nor U35285 (N_35285,N_34354,N_34498);
xor U35286 (N_35286,N_34814,N_34959);
and U35287 (N_35287,N_34662,N_34328);
or U35288 (N_35288,N_34990,N_34107);
nor U35289 (N_35289,N_34042,N_34706);
and U35290 (N_35290,N_34110,N_34300);
nand U35291 (N_35291,N_34452,N_34919);
or U35292 (N_35292,N_34703,N_34585);
xor U35293 (N_35293,N_34379,N_34318);
nor U35294 (N_35294,N_34756,N_34370);
nand U35295 (N_35295,N_34858,N_34256);
or U35296 (N_35296,N_34930,N_34496);
or U35297 (N_35297,N_34900,N_34411);
and U35298 (N_35298,N_34405,N_34386);
xnor U35299 (N_35299,N_34553,N_34055);
xnor U35300 (N_35300,N_34450,N_34038);
xnor U35301 (N_35301,N_34672,N_34387);
or U35302 (N_35302,N_34422,N_34121);
or U35303 (N_35303,N_34057,N_34073);
or U35304 (N_35304,N_34529,N_34770);
nand U35305 (N_35305,N_34596,N_34856);
xor U35306 (N_35306,N_34462,N_34371);
xor U35307 (N_35307,N_34063,N_34976);
nand U35308 (N_35308,N_34356,N_34507);
nor U35309 (N_35309,N_34088,N_34184);
nand U35310 (N_35310,N_34136,N_34795);
and U35311 (N_35311,N_34831,N_34630);
and U35312 (N_35312,N_34943,N_34475);
nand U35313 (N_35313,N_34868,N_34847);
and U35314 (N_35314,N_34668,N_34802);
nand U35315 (N_35315,N_34390,N_34994);
nor U35316 (N_35316,N_34872,N_34721);
and U35317 (N_35317,N_34401,N_34330);
or U35318 (N_35318,N_34909,N_34871);
nand U35319 (N_35319,N_34515,N_34017);
nand U35320 (N_35320,N_34969,N_34547);
nor U35321 (N_35321,N_34466,N_34190);
xnor U35322 (N_35322,N_34044,N_34901);
nand U35323 (N_35323,N_34837,N_34842);
nor U35324 (N_35324,N_34403,N_34490);
nor U35325 (N_35325,N_34962,N_34435);
and U35326 (N_35326,N_34908,N_34776);
and U35327 (N_35327,N_34807,N_34155);
nor U35328 (N_35328,N_34545,N_34380);
nor U35329 (N_35329,N_34567,N_34166);
and U35330 (N_35330,N_34569,N_34604);
xor U35331 (N_35331,N_34631,N_34091);
and U35332 (N_35332,N_34417,N_34726);
nor U35333 (N_35333,N_34492,N_34895);
or U35334 (N_35334,N_34309,N_34513);
nor U35335 (N_35335,N_34981,N_34881);
nor U35336 (N_35336,N_34713,N_34841);
and U35337 (N_35337,N_34665,N_34752);
nor U35338 (N_35338,N_34783,N_34931);
nor U35339 (N_35339,N_34280,N_34276);
or U35340 (N_35340,N_34673,N_34394);
nor U35341 (N_35341,N_34003,N_34894);
nor U35342 (N_35342,N_34341,N_34048);
or U35343 (N_35343,N_34258,N_34968);
nor U35344 (N_35344,N_34742,N_34960);
and U35345 (N_35345,N_34198,N_34347);
nand U35346 (N_35346,N_34712,N_34494);
nor U35347 (N_35347,N_34179,N_34064);
nand U35348 (N_35348,N_34929,N_34212);
nor U35349 (N_35349,N_34149,N_34196);
xor U35350 (N_35350,N_34551,N_34339);
and U35351 (N_35351,N_34262,N_34282);
xor U35352 (N_35352,N_34661,N_34350);
and U35353 (N_35353,N_34245,N_34474);
and U35354 (N_35354,N_34548,N_34495);
nor U35355 (N_35355,N_34961,N_34509);
xor U35356 (N_35356,N_34675,N_34230);
or U35357 (N_35357,N_34372,N_34289);
nor U35358 (N_35358,N_34069,N_34139);
or U35359 (N_35359,N_34607,N_34750);
or U35360 (N_35360,N_34947,N_34539);
nor U35361 (N_35361,N_34669,N_34797);
nand U35362 (N_35362,N_34429,N_34690);
nand U35363 (N_35363,N_34278,N_34060);
and U35364 (N_35364,N_34206,N_34362);
nor U35365 (N_35365,N_34514,N_34290);
and U35366 (N_35366,N_34013,N_34265);
xnor U35367 (N_35367,N_34622,N_34428);
nand U35368 (N_35368,N_34232,N_34617);
or U35369 (N_35369,N_34898,N_34033);
or U35370 (N_35370,N_34052,N_34094);
or U35371 (N_35371,N_34291,N_34225);
xnor U35372 (N_35372,N_34439,N_34667);
or U35373 (N_35373,N_34423,N_34158);
nor U35374 (N_35374,N_34205,N_34887);
or U35375 (N_35375,N_34611,N_34172);
nor U35376 (N_35376,N_34592,N_34815);
nand U35377 (N_35377,N_34243,N_34385);
xor U35378 (N_35378,N_34836,N_34730);
or U35379 (N_35379,N_34457,N_34414);
xor U35380 (N_35380,N_34191,N_34735);
xor U35381 (N_35381,N_34098,N_34221);
nand U35382 (N_35382,N_34283,N_34791);
xnor U35383 (N_35383,N_34533,N_34719);
or U35384 (N_35384,N_34187,N_34893);
xor U35385 (N_35385,N_34214,N_34762);
nor U35386 (N_35386,N_34185,N_34955);
and U35387 (N_35387,N_34483,N_34319);
nand U35388 (N_35388,N_34066,N_34311);
and U35389 (N_35389,N_34505,N_34381);
or U35390 (N_35390,N_34425,N_34025);
or U35391 (N_35391,N_34753,N_34171);
nand U35392 (N_35392,N_34368,N_34194);
and U35393 (N_35393,N_34164,N_34743);
nor U35394 (N_35394,N_34688,N_34942);
xnor U35395 (N_35395,N_34489,N_34575);
nand U35396 (N_35396,N_34445,N_34897);
xor U35397 (N_35397,N_34835,N_34740);
nor U35398 (N_35398,N_34768,N_34804);
xnor U35399 (N_35399,N_34767,N_34482);
or U35400 (N_35400,N_34779,N_34034);
xnor U35401 (N_35401,N_34967,N_34741);
or U35402 (N_35402,N_34716,N_34681);
xnor U35403 (N_35403,N_34092,N_34329);
xor U35404 (N_35404,N_34470,N_34023);
xnor U35405 (N_35405,N_34296,N_34705);
and U35406 (N_35406,N_34615,N_34304);
nor U35407 (N_35407,N_34629,N_34284);
xnor U35408 (N_35408,N_34840,N_34995);
or U35409 (N_35409,N_34224,N_34485);
or U35410 (N_35410,N_34710,N_34183);
or U35411 (N_35411,N_34029,N_34916);
or U35412 (N_35412,N_34800,N_34974);
and U35413 (N_35413,N_34160,N_34781);
nor U35414 (N_35414,N_34366,N_34269);
nor U35415 (N_35415,N_34195,N_34677);
or U35416 (N_35416,N_34749,N_34287);
nor U35417 (N_35417,N_34000,N_34373);
or U35418 (N_35418,N_34464,N_34886);
or U35419 (N_35419,N_34695,N_34484);
and U35420 (N_35420,N_34639,N_34951);
xor U35421 (N_35421,N_34297,N_34441);
xor U35422 (N_35422,N_34666,N_34518);
or U35423 (N_35423,N_34963,N_34616);
nand U35424 (N_35424,N_34438,N_34859);
or U35425 (N_35425,N_34469,N_34625);
and U35426 (N_35426,N_34769,N_34525);
or U35427 (N_35427,N_34580,N_34295);
nand U35428 (N_35428,N_34755,N_34510);
and U35429 (N_35429,N_34448,N_34313);
nor U35430 (N_35430,N_34040,N_34659);
or U35431 (N_35431,N_34913,N_34543);
or U35432 (N_35432,N_34645,N_34966);
and U35433 (N_35433,N_34400,N_34497);
or U35434 (N_35434,N_34860,N_34957);
xnor U35435 (N_35435,N_34605,N_34784);
nor U35436 (N_35436,N_34722,N_34263);
and U35437 (N_35437,N_34078,N_34125);
and U35438 (N_35438,N_34891,N_34117);
and U35439 (N_35439,N_34827,N_34156);
xnor U35440 (N_35440,N_34440,N_34315);
and U35441 (N_35441,N_34601,N_34907);
or U35442 (N_35442,N_34811,N_34141);
and U35443 (N_35443,N_34231,N_34471);
nand U35444 (N_35444,N_34558,N_34903);
and U35445 (N_35445,N_34410,N_34635);
nand U35446 (N_35446,N_34540,N_34093);
xnor U35447 (N_35447,N_34511,N_34465);
xor U35448 (N_35448,N_34080,N_34180);
nor U35449 (N_35449,N_34391,N_34564);
xor U35450 (N_35450,N_34292,N_34905);
xnor U35451 (N_35451,N_34061,N_34949);
and U35452 (N_35452,N_34257,N_34973);
nand U35453 (N_35453,N_34590,N_34626);
xnor U35454 (N_35454,N_34977,N_34819);
or U35455 (N_35455,N_34415,N_34892);
nand U35456 (N_35456,N_34235,N_34809);
xor U35457 (N_35457,N_34173,N_34102);
and U35458 (N_35458,N_34157,N_34594);
nor U35459 (N_35459,N_34833,N_34326);
nand U35460 (N_35460,N_34028,N_34816);
xor U35461 (N_35461,N_34921,N_34899);
and U35462 (N_35462,N_34397,N_34067);
nand U35463 (N_35463,N_34637,N_34697);
and U35464 (N_35464,N_34925,N_34426);
nor U35465 (N_35465,N_34782,N_34271);
nand U35466 (N_35466,N_34279,N_34593);
or U35467 (N_35467,N_34451,N_34989);
xor U35468 (N_35468,N_34177,N_34535);
or U35469 (N_35469,N_34344,N_34197);
or U35470 (N_35470,N_34434,N_34095);
nor U35471 (N_35471,N_34928,N_34701);
xor U35472 (N_35472,N_34948,N_34476);
nor U35473 (N_35473,N_34135,N_34134);
and U35474 (N_35474,N_34041,N_34461);
nor U35475 (N_35475,N_34861,N_34711);
xnor U35476 (N_35476,N_34524,N_34109);
or U35477 (N_35477,N_34099,N_34984);
xnor U35478 (N_35478,N_34421,N_34570);
nand U35479 (N_35479,N_34599,N_34803);
or U35480 (N_35480,N_34725,N_34143);
and U35481 (N_35481,N_34020,N_34480);
nor U35482 (N_35482,N_34298,N_34236);
nor U35483 (N_35483,N_34724,N_34193);
nand U35484 (N_35484,N_34472,N_34660);
xor U35485 (N_35485,N_34739,N_34772);
or U35486 (N_35486,N_34737,N_34106);
xor U35487 (N_35487,N_34442,N_34874);
nand U35488 (N_35488,N_34975,N_34699);
or U35489 (N_35489,N_34409,N_34556);
and U35490 (N_35490,N_34455,N_34246);
or U35491 (N_35491,N_34337,N_34201);
and U35492 (N_35492,N_34915,N_34532);
or U35493 (N_35493,N_34531,N_34047);
or U35494 (N_35494,N_34192,N_34012);
nand U35495 (N_35495,N_34709,N_34436);
and U35496 (N_35496,N_34303,N_34266);
nor U35497 (N_35497,N_34275,N_34343);
or U35498 (N_35498,N_34142,N_34876);
or U35499 (N_35499,N_34700,N_34799);
and U35500 (N_35500,N_34468,N_34245);
nand U35501 (N_35501,N_34129,N_34494);
and U35502 (N_35502,N_34473,N_34168);
xor U35503 (N_35503,N_34596,N_34802);
xor U35504 (N_35504,N_34723,N_34820);
or U35505 (N_35505,N_34279,N_34883);
nand U35506 (N_35506,N_34415,N_34345);
xor U35507 (N_35507,N_34526,N_34734);
or U35508 (N_35508,N_34473,N_34183);
xor U35509 (N_35509,N_34257,N_34210);
nand U35510 (N_35510,N_34640,N_34654);
nand U35511 (N_35511,N_34866,N_34414);
nand U35512 (N_35512,N_34340,N_34317);
nand U35513 (N_35513,N_34239,N_34454);
xor U35514 (N_35514,N_34131,N_34739);
nor U35515 (N_35515,N_34628,N_34543);
nand U35516 (N_35516,N_34911,N_34694);
nand U35517 (N_35517,N_34212,N_34238);
nand U35518 (N_35518,N_34768,N_34969);
nor U35519 (N_35519,N_34611,N_34354);
and U35520 (N_35520,N_34061,N_34817);
and U35521 (N_35521,N_34142,N_34412);
xnor U35522 (N_35522,N_34938,N_34254);
xnor U35523 (N_35523,N_34798,N_34291);
or U35524 (N_35524,N_34100,N_34901);
or U35525 (N_35525,N_34382,N_34634);
nor U35526 (N_35526,N_34170,N_34376);
xor U35527 (N_35527,N_34879,N_34784);
nor U35528 (N_35528,N_34373,N_34274);
xor U35529 (N_35529,N_34602,N_34538);
nor U35530 (N_35530,N_34795,N_34391);
and U35531 (N_35531,N_34386,N_34628);
nor U35532 (N_35532,N_34376,N_34011);
xor U35533 (N_35533,N_34865,N_34436);
xor U35534 (N_35534,N_34825,N_34281);
xnor U35535 (N_35535,N_34872,N_34056);
and U35536 (N_35536,N_34377,N_34321);
nand U35537 (N_35537,N_34468,N_34209);
xor U35538 (N_35538,N_34549,N_34917);
nand U35539 (N_35539,N_34872,N_34754);
xnor U35540 (N_35540,N_34478,N_34534);
xor U35541 (N_35541,N_34979,N_34696);
xor U35542 (N_35542,N_34047,N_34180);
or U35543 (N_35543,N_34208,N_34065);
nand U35544 (N_35544,N_34709,N_34987);
nand U35545 (N_35545,N_34423,N_34768);
nor U35546 (N_35546,N_34868,N_34731);
nand U35547 (N_35547,N_34010,N_34444);
xor U35548 (N_35548,N_34672,N_34679);
nand U35549 (N_35549,N_34598,N_34053);
xnor U35550 (N_35550,N_34754,N_34976);
nor U35551 (N_35551,N_34176,N_34875);
xor U35552 (N_35552,N_34305,N_34509);
nand U35553 (N_35553,N_34218,N_34961);
nor U35554 (N_35554,N_34848,N_34929);
xor U35555 (N_35555,N_34322,N_34825);
nor U35556 (N_35556,N_34467,N_34034);
nor U35557 (N_35557,N_34480,N_34885);
nor U35558 (N_35558,N_34896,N_34460);
or U35559 (N_35559,N_34672,N_34393);
and U35560 (N_35560,N_34566,N_34158);
or U35561 (N_35561,N_34070,N_34450);
nor U35562 (N_35562,N_34369,N_34579);
or U35563 (N_35563,N_34814,N_34298);
and U35564 (N_35564,N_34967,N_34181);
xnor U35565 (N_35565,N_34285,N_34877);
and U35566 (N_35566,N_34118,N_34125);
and U35567 (N_35567,N_34217,N_34851);
xor U35568 (N_35568,N_34517,N_34791);
and U35569 (N_35569,N_34838,N_34267);
nand U35570 (N_35570,N_34691,N_34172);
xnor U35571 (N_35571,N_34389,N_34579);
nor U35572 (N_35572,N_34366,N_34344);
xnor U35573 (N_35573,N_34914,N_34780);
and U35574 (N_35574,N_34651,N_34467);
nand U35575 (N_35575,N_34050,N_34186);
and U35576 (N_35576,N_34184,N_34174);
and U35577 (N_35577,N_34961,N_34476);
nor U35578 (N_35578,N_34685,N_34885);
nor U35579 (N_35579,N_34058,N_34517);
and U35580 (N_35580,N_34655,N_34241);
nand U35581 (N_35581,N_34874,N_34942);
nand U35582 (N_35582,N_34253,N_34468);
xor U35583 (N_35583,N_34201,N_34999);
xor U35584 (N_35584,N_34354,N_34239);
or U35585 (N_35585,N_34088,N_34421);
or U35586 (N_35586,N_34092,N_34444);
nor U35587 (N_35587,N_34986,N_34025);
nor U35588 (N_35588,N_34166,N_34650);
and U35589 (N_35589,N_34232,N_34625);
xor U35590 (N_35590,N_34713,N_34008);
nand U35591 (N_35591,N_34251,N_34631);
xor U35592 (N_35592,N_34424,N_34927);
and U35593 (N_35593,N_34651,N_34205);
xor U35594 (N_35594,N_34077,N_34614);
nor U35595 (N_35595,N_34455,N_34475);
nor U35596 (N_35596,N_34773,N_34891);
nor U35597 (N_35597,N_34138,N_34953);
and U35598 (N_35598,N_34760,N_34863);
or U35599 (N_35599,N_34991,N_34009);
nand U35600 (N_35600,N_34990,N_34212);
or U35601 (N_35601,N_34443,N_34189);
xnor U35602 (N_35602,N_34880,N_34239);
xnor U35603 (N_35603,N_34075,N_34366);
xnor U35604 (N_35604,N_34237,N_34608);
or U35605 (N_35605,N_34449,N_34895);
and U35606 (N_35606,N_34229,N_34371);
xor U35607 (N_35607,N_34935,N_34528);
and U35608 (N_35608,N_34238,N_34053);
and U35609 (N_35609,N_34276,N_34680);
xor U35610 (N_35610,N_34582,N_34740);
nand U35611 (N_35611,N_34659,N_34052);
and U35612 (N_35612,N_34819,N_34868);
and U35613 (N_35613,N_34426,N_34040);
xnor U35614 (N_35614,N_34554,N_34325);
nor U35615 (N_35615,N_34147,N_34419);
nand U35616 (N_35616,N_34805,N_34192);
nor U35617 (N_35617,N_34963,N_34388);
and U35618 (N_35618,N_34861,N_34897);
or U35619 (N_35619,N_34168,N_34680);
nor U35620 (N_35620,N_34618,N_34783);
nor U35621 (N_35621,N_34042,N_34559);
nand U35622 (N_35622,N_34705,N_34832);
xor U35623 (N_35623,N_34009,N_34003);
and U35624 (N_35624,N_34402,N_34598);
or U35625 (N_35625,N_34514,N_34493);
nor U35626 (N_35626,N_34017,N_34045);
xor U35627 (N_35627,N_34998,N_34746);
nand U35628 (N_35628,N_34725,N_34726);
nor U35629 (N_35629,N_34684,N_34981);
nor U35630 (N_35630,N_34157,N_34895);
xor U35631 (N_35631,N_34740,N_34284);
and U35632 (N_35632,N_34706,N_34458);
nand U35633 (N_35633,N_34168,N_34019);
nand U35634 (N_35634,N_34754,N_34752);
or U35635 (N_35635,N_34091,N_34664);
nand U35636 (N_35636,N_34941,N_34665);
xnor U35637 (N_35637,N_34543,N_34734);
and U35638 (N_35638,N_34579,N_34966);
nand U35639 (N_35639,N_34742,N_34976);
or U35640 (N_35640,N_34879,N_34466);
and U35641 (N_35641,N_34509,N_34130);
nor U35642 (N_35642,N_34682,N_34910);
or U35643 (N_35643,N_34988,N_34725);
xor U35644 (N_35644,N_34395,N_34110);
xnor U35645 (N_35645,N_34364,N_34907);
xnor U35646 (N_35646,N_34716,N_34894);
and U35647 (N_35647,N_34316,N_34109);
xor U35648 (N_35648,N_34245,N_34898);
xor U35649 (N_35649,N_34819,N_34691);
xnor U35650 (N_35650,N_34497,N_34853);
xor U35651 (N_35651,N_34081,N_34299);
or U35652 (N_35652,N_34405,N_34509);
nand U35653 (N_35653,N_34357,N_34214);
nor U35654 (N_35654,N_34102,N_34826);
nand U35655 (N_35655,N_34074,N_34342);
nand U35656 (N_35656,N_34526,N_34906);
xor U35657 (N_35657,N_34856,N_34859);
or U35658 (N_35658,N_34202,N_34578);
and U35659 (N_35659,N_34775,N_34147);
and U35660 (N_35660,N_34139,N_34917);
xor U35661 (N_35661,N_34312,N_34848);
nor U35662 (N_35662,N_34799,N_34849);
and U35663 (N_35663,N_34015,N_34249);
or U35664 (N_35664,N_34597,N_34311);
nor U35665 (N_35665,N_34482,N_34271);
nand U35666 (N_35666,N_34968,N_34913);
or U35667 (N_35667,N_34704,N_34383);
or U35668 (N_35668,N_34293,N_34597);
nor U35669 (N_35669,N_34260,N_34983);
xnor U35670 (N_35670,N_34804,N_34553);
or U35671 (N_35671,N_34228,N_34852);
and U35672 (N_35672,N_34403,N_34619);
or U35673 (N_35673,N_34071,N_34810);
or U35674 (N_35674,N_34582,N_34462);
nand U35675 (N_35675,N_34526,N_34267);
and U35676 (N_35676,N_34938,N_34746);
nor U35677 (N_35677,N_34335,N_34497);
or U35678 (N_35678,N_34948,N_34609);
nor U35679 (N_35679,N_34918,N_34602);
nand U35680 (N_35680,N_34546,N_34073);
or U35681 (N_35681,N_34710,N_34962);
xor U35682 (N_35682,N_34293,N_34515);
and U35683 (N_35683,N_34179,N_34393);
nand U35684 (N_35684,N_34869,N_34042);
xor U35685 (N_35685,N_34368,N_34109);
nand U35686 (N_35686,N_34293,N_34363);
nor U35687 (N_35687,N_34426,N_34421);
xor U35688 (N_35688,N_34159,N_34389);
nand U35689 (N_35689,N_34135,N_34187);
and U35690 (N_35690,N_34154,N_34758);
or U35691 (N_35691,N_34180,N_34569);
nor U35692 (N_35692,N_34044,N_34400);
nand U35693 (N_35693,N_34225,N_34926);
and U35694 (N_35694,N_34390,N_34779);
and U35695 (N_35695,N_34439,N_34361);
nor U35696 (N_35696,N_34232,N_34792);
nor U35697 (N_35697,N_34438,N_34346);
nor U35698 (N_35698,N_34866,N_34771);
and U35699 (N_35699,N_34100,N_34011);
and U35700 (N_35700,N_34805,N_34591);
nand U35701 (N_35701,N_34658,N_34853);
nand U35702 (N_35702,N_34093,N_34909);
nor U35703 (N_35703,N_34371,N_34777);
xor U35704 (N_35704,N_34331,N_34182);
or U35705 (N_35705,N_34037,N_34314);
nor U35706 (N_35706,N_34151,N_34378);
or U35707 (N_35707,N_34125,N_34154);
xor U35708 (N_35708,N_34122,N_34316);
or U35709 (N_35709,N_34563,N_34743);
nor U35710 (N_35710,N_34857,N_34518);
and U35711 (N_35711,N_34040,N_34515);
nand U35712 (N_35712,N_34767,N_34857);
nand U35713 (N_35713,N_34823,N_34962);
xnor U35714 (N_35714,N_34407,N_34485);
and U35715 (N_35715,N_34683,N_34194);
nand U35716 (N_35716,N_34256,N_34966);
nand U35717 (N_35717,N_34908,N_34248);
nor U35718 (N_35718,N_34922,N_34737);
nand U35719 (N_35719,N_34642,N_34626);
or U35720 (N_35720,N_34272,N_34997);
nor U35721 (N_35721,N_34597,N_34358);
xor U35722 (N_35722,N_34174,N_34958);
and U35723 (N_35723,N_34466,N_34309);
xor U35724 (N_35724,N_34091,N_34940);
nor U35725 (N_35725,N_34513,N_34307);
and U35726 (N_35726,N_34182,N_34513);
xnor U35727 (N_35727,N_34594,N_34295);
nand U35728 (N_35728,N_34986,N_34479);
xor U35729 (N_35729,N_34029,N_34416);
or U35730 (N_35730,N_34322,N_34262);
or U35731 (N_35731,N_34918,N_34536);
or U35732 (N_35732,N_34557,N_34613);
or U35733 (N_35733,N_34573,N_34097);
xnor U35734 (N_35734,N_34886,N_34033);
nand U35735 (N_35735,N_34485,N_34260);
and U35736 (N_35736,N_34623,N_34532);
nor U35737 (N_35737,N_34954,N_34117);
and U35738 (N_35738,N_34805,N_34173);
and U35739 (N_35739,N_34534,N_34588);
nand U35740 (N_35740,N_34402,N_34758);
nor U35741 (N_35741,N_34434,N_34340);
nand U35742 (N_35742,N_34840,N_34701);
nor U35743 (N_35743,N_34766,N_34814);
or U35744 (N_35744,N_34647,N_34188);
nand U35745 (N_35745,N_34843,N_34378);
xnor U35746 (N_35746,N_34092,N_34760);
or U35747 (N_35747,N_34078,N_34753);
or U35748 (N_35748,N_34061,N_34870);
or U35749 (N_35749,N_34696,N_34703);
and U35750 (N_35750,N_34129,N_34680);
and U35751 (N_35751,N_34608,N_34585);
or U35752 (N_35752,N_34875,N_34463);
or U35753 (N_35753,N_34218,N_34318);
nand U35754 (N_35754,N_34578,N_34348);
xor U35755 (N_35755,N_34875,N_34103);
nor U35756 (N_35756,N_34566,N_34472);
xor U35757 (N_35757,N_34685,N_34814);
nand U35758 (N_35758,N_34594,N_34361);
or U35759 (N_35759,N_34619,N_34406);
nor U35760 (N_35760,N_34361,N_34176);
nand U35761 (N_35761,N_34900,N_34942);
and U35762 (N_35762,N_34251,N_34958);
and U35763 (N_35763,N_34980,N_34852);
nor U35764 (N_35764,N_34658,N_34371);
nand U35765 (N_35765,N_34166,N_34211);
xor U35766 (N_35766,N_34933,N_34145);
nand U35767 (N_35767,N_34573,N_34826);
xnor U35768 (N_35768,N_34773,N_34249);
or U35769 (N_35769,N_34126,N_34502);
or U35770 (N_35770,N_34297,N_34354);
nor U35771 (N_35771,N_34134,N_34039);
nor U35772 (N_35772,N_34948,N_34112);
xor U35773 (N_35773,N_34409,N_34530);
nand U35774 (N_35774,N_34119,N_34723);
xnor U35775 (N_35775,N_34649,N_34511);
xor U35776 (N_35776,N_34292,N_34906);
or U35777 (N_35777,N_34252,N_34732);
nand U35778 (N_35778,N_34959,N_34557);
or U35779 (N_35779,N_34727,N_34316);
or U35780 (N_35780,N_34450,N_34379);
xor U35781 (N_35781,N_34406,N_34981);
nand U35782 (N_35782,N_34184,N_34026);
nand U35783 (N_35783,N_34739,N_34176);
and U35784 (N_35784,N_34393,N_34572);
nand U35785 (N_35785,N_34775,N_34596);
nor U35786 (N_35786,N_34558,N_34901);
nor U35787 (N_35787,N_34269,N_34391);
and U35788 (N_35788,N_34750,N_34845);
or U35789 (N_35789,N_34900,N_34153);
or U35790 (N_35790,N_34283,N_34756);
and U35791 (N_35791,N_34470,N_34926);
xnor U35792 (N_35792,N_34706,N_34159);
nor U35793 (N_35793,N_34166,N_34834);
nand U35794 (N_35794,N_34075,N_34557);
nand U35795 (N_35795,N_34687,N_34992);
and U35796 (N_35796,N_34767,N_34999);
nand U35797 (N_35797,N_34755,N_34631);
and U35798 (N_35798,N_34749,N_34425);
xor U35799 (N_35799,N_34517,N_34897);
xor U35800 (N_35800,N_34117,N_34282);
nor U35801 (N_35801,N_34368,N_34351);
nor U35802 (N_35802,N_34796,N_34733);
or U35803 (N_35803,N_34623,N_34193);
xor U35804 (N_35804,N_34896,N_34181);
or U35805 (N_35805,N_34357,N_34137);
and U35806 (N_35806,N_34237,N_34983);
xnor U35807 (N_35807,N_34853,N_34542);
nand U35808 (N_35808,N_34417,N_34682);
and U35809 (N_35809,N_34804,N_34544);
nor U35810 (N_35810,N_34243,N_34790);
xor U35811 (N_35811,N_34055,N_34634);
xnor U35812 (N_35812,N_34913,N_34338);
nand U35813 (N_35813,N_34969,N_34588);
xnor U35814 (N_35814,N_34882,N_34690);
or U35815 (N_35815,N_34600,N_34981);
or U35816 (N_35816,N_34096,N_34289);
or U35817 (N_35817,N_34418,N_34030);
or U35818 (N_35818,N_34461,N_34653);
and U35819 (N_35819,N_34157,N_34723);
or U35820 (N_35820,N_34360,N_34251);
nor U35821 (N_35821,N_34483,N_34291);
or U35822 (N_35822,N_34576,N_34104);
xor U35823 (N_35823,N_34043,N_34592);
and U35824 (N_35824,N_34446,N_34773);
nor U35825 (N_35825,N_34729,N_34834);
nand U35826 (N_35826,N_34901,N_34809);
nor U35827 (N_35827,N_34969,N_34981);
xnor U35828 (N_35828,N_34193,N_34497);
or U35829 (N_35829,N_34068,N_34036);
nor U35830 (N_35830,N_34539,N_34966);
xnor U35831 (N_35831,N_34542,N_34619);
nor U35832 (N_35832,N_34257,N_34511);
or U35833 (N_35833,N_34154,N_34053);
xnor U35834 (N_35834,N_34413,N_34699);
and U35835 (N_35835,N_34116,N_34017);
and U35836 (N_35836,N_34831,N_34447);
or U35837 (N_35837,N_34316,N_34575);
and U35838 (N_35838,N_34128,N_34460);
or U35839 (N_35839,N_34475,N_34079);
nor U35840 (N_35840,N_34123,N_34431);
or U35841 (N_35841,N_34681,N_34271);
or U35842 (N_35842,N_34990,N_34486);
or U35843 (N_35843,N_34608,N_34193);
nor U35844 (N_35844,N_34417,N_34985);
xor U35845 (N_35845,N_34404,N_34838);
xor U35846 (N_35846,N_34800,N_34846);
and U35847 (N_35847,N_34190,N_34718);
and U35848 (N_35848,N_34300,N_34025);
and U35849 (N_35849,N_34597,N_34099);
nand U35850 (N_35850,N_34743,N_34956);
and U35851 (N_35851,N_34907,N_34889);
or U35852 (N_35852,N_34582,N_34314);
nor U35853 (N_35853,N_34782,N_34057);
nand U35854 (N_35854,N_34535,N_34704);
or U35855 (N_35855,N_34707,N_34622);
nor U35856 (N_35856,N_34491,N_34275);
and U35857 (N_35857,N_34569,N_34920);
or U35858 (N_35858,N_34699,N_34436);
or U35859 (N_35859,N_34459,N_34641);
or U35860 (N_35860,N_34458,N_34143);
or U35861 (N_35861,N_34148,N_34758);
and U35862 (N_35862,N_34846,N_34377);
or U35863 (N_35863,N_34000,N_34831);
and U35864 (N_35864,N_34563,N_34859);
nor U35865 (N_35865,N_34580,N_34826);
or U35866 (N_35866,N_34601,N_34395);
and U35867 (N_35867,N_34142,N_34586);
xnor U35868 (N_35868,N_34227,N_34449);
nor U35869 (N_35869,N_34019,N_34956);
and U35870 (N_35870,N_34912,N_34588);
xnor U35871 (N_35871,N_34232,N_34789);
nand U35872 (N_35872,N_34967,N_34478);
xnor U35873 (N_35873,N_34947,N_34287);
xnor U35874 (N_35874,N_34479,N_34100);
nor U35875 (N_35875,N_34547,N_34699);
nand U35876 (N_35876,N_34931,N_34379);
and U35877 (N_35877,N_34369,N_34870);
xor U35878 (N_35878,N_34508,N_34190);
and U35879 (N_35879,N_34499,N_34449);
xor U35880 (N_35880,N_34963,N_34945);
nor U35881 (N_35881,N_34079,N_34493);
xnor U35882 (N_35882,N_34883,N_34754);
nand U35883 (N_35883,N_34577,N_34559);
nand U35884 (N_35884,N_34386,N_34504);
and U35885 (N_35885,N_34600,N_34588);
nor U35886 (N_35886,N_34091,N_34827);
and U35887 (N_35887,N_34425,N_34678);
nand U35888 (N_35888,N_34103,N_34370);
xnor U35889 (N_35889,N_34055,N_34551);
and U35890 (N_35890,N_34615,N_34447);
nor U35891 (N_35891,N_34270,N_34615);
nor U35892 (N_35892,N_34957,N_34068);
or U35893 (N_35893,N_34719,N_34168);
nand U35894 (N_35894,N_34892,N_34318);
xor U35895 (N_35895,N_34225,N_34718);
or U35896 (N_35896,N_34069,N_34583);
nand U35897 (N_35897,N_34470,N_34127);
nor U35898 (N_35898,N_34235,N_34291);
and U35899 (N_35899,N_34128,N_34568);
nand U35900 (N_35900,N_34670,N_34697);
xnor U35901 (N_35901,N_34863,N_34085);
or U35902 (N_35902,N_34590,N_34441);
and U35903 (N_35903,N_34870,N_34950);
nor U35904 (N_35904,N_34120,N_34742);
nor U35905 (N_35905,N_34702,N_34857);
and U35906 (N_35906,N_34039,N_34771);
nor U35907 (N_35907,N_34931,N_34014);
nor U35908 (N_35908,N_34655,N_34528);
xor U35909 (N_35909,N_34530,N_34231);
nand U35910 (N_35910,N_34608,N_34200);
xor U35911 (N_35911,N_34932,N_34548);
nand U35912 (N_35912,N_34274,N_34051);
nand U35913 (N_35913,N_34096,N_34299);
xor U35914 (N_35914,N_34567,N_34873);
nor U35915 (N_35915,N_34083,N_34431);
or U35916 (N_35916,N_34602,N_34941);
and U35917 (N_35917,N_34335,N_34283);
and U35918 (N_35918,N_34095,N_34747);
or U35919 (N_35919,N_34197,N_34940);
or U35920 (N_35920,N_34384,N_34193);
nand U35921 (N_35921,N_34315,N_34010);
or U35922 (N_35922,N_34719,N_34129);
or U35923 (N_35923,N_34598,N_34336);
nor U35924 (N_35924,N_34773,N_34422);
and U35925 (N_35925,N_34323,N_34609);
nor U35926 (N_35926,N_34046,N_34181);
and U35927 (N_35927,N_34503,N_34378);
xor U35928 (N_35928,N_34732,N_34168);
nor U35929 (N_35929,N_34726,N_34499);
nor U35930 (N_35930,N_34936,N_34896);
nor U35931 (N_35931,N_34668,N_34514);
nor U35932 (N_35932,N_34050,N_34070);
nand U35933 (N_35933,N_34638,N_34419);
nand U35934 (N_35934,N_34500,N_34637);
xnor U35935 (N_35935,N_34414,N_34996);
xnor U35936 (N_35936,N_34162,N_34618);
nor U35937 (N_35937,N_34657,N_34989);
nand U35938 (N_35938,N_34972,N_34659);
nand U35939 (N_35939,N_34198,N_34230);
or U35940 (N_35940,N_34925,N_34765);
and U35941 (N_35941,N_34729,N_34860);
xor U35942 (N_35942,N_34507,N_34574);
xor U35943 (N_35943,N_34890,N_34949);
nor U35944 (N_35944,N_34155,N_34372);
and U35945 (N_35945,N_34680,N_34883);
xor U35946 (N_35946,N_34996,N_34032);
xor U35947 (N_35947,N_34177,N_34281);
xnor U35948 (N_35948,N_34263,N_34900);
xor U35949 (N_35949,N_34457,N_34213);
xnor U35950 (N_35950,N_34981,N_34420);
and U35951 (N_35951,N_34067,N_34122);
and U35952 (N_35952,N_34950,N_34400);
nor U35953 (N_35953,N_34872,N_34937);
and U35954 (N_35954,N_34335,N_34644);
or U35955 (N_35955,N_34591,N_34113);
and U35956 (N_35956,N_34147,N_34148);
and U35957 (N_35957,N_34699,N_34677);
or U35958 (N_35958,N_34075,N_34118);
and U35959 (N_35959,N_34770,N_34128);
nand U35960 (N_35960,N_34480,N_34631);
or U35961 (N_35961,N_34958,N_34141);
or U35962 (N_35962,N_34681,N_34294);
and U35963 (N_35963,N_34340,N_34636);
nor U35964 (N_35964,N_34726,N_34802);
and U35965 (N_35965,N_34947,N_34723);
nor U35966 (N_35966,N_34426,N_34807);
xor U35967 (N_35967,N_34066,N_34752);
or U35968 (N_35968,N_34577,N_34320);
nor U35969 (N_35969,N_34291,N_34639);
nor U35970 (N_35970,N_34347,N_34279);
nor U35971 (N_35971,N_34145,N_34910);
xnor U35972 (N_35972,N_34346,N_34388);
xor U35973 (N_35973,N_34654,N_34139);
or U35974 (N_35974,N_34164,N_34476);
nand U35975 (N_35975,N_34607,N_34307);
xnor U35976 (N_35976,N_34931,N_34353);
and U35977 (N_35977,N_34683,N_34103);
nand U35978 (N_35978,N_34803,N_34128);
nor U35979 (N_35979,N_34335,N_34214);
or U35980 (N_35980,N_34612,N_34207);
nand U35981 (N_35981,N_34018,N_34482);
xor U35982 (N_35982,N_34780,N_34432);
and U35983 (N_35983,N_34926,N_34456);
nor U35984 (N_35984,N_34323,N_34512);
xnor U35985 (N_35985,N_34250,N_34629);
and U35986 (N_35986,N_34965,N_34463);
xor U35987 (N_35987,N_34317,N_34663);
or U35988 (N_35988,N_34850,N_34817);
nand U35989 (N_35989,N_34338,N_34493);
and U35990 (N_35990,N_34042,N_34352);
xnor U35991 (N_35991,N_34910,N_34092);
xnor U35992 (N_35992,N_34724,N_34085);
nand U35993 (N_35993,N_34230,N_34307);
xor U35994 (N_35994,N_34672,N_34490);
and U35995 (N_35995,N_34502,N_34960);
nand U35996 (N_35996,N_34530,N_34523);
or U35997 (N_35997,N_34010,N_34193);
nand U35998 (N_35998,N_34236,N_34426);
nand U35999 (N_35999,N_34420,N_34337);
xnor U36000 (N_36000,N_35862,N_35975);
nand U36001 (N_36001,N_35620,N_35530);
nand U36002 (N_36002,N_35427,N_35450);
nand U36003 (N_36003,N_35008,N_35354);
nand U36004 (N_36004,N_35646,N_35472);
xor U36005 (N_36005,N_35150,N_35383);
nand U36006 (N_36006,N_35602,N_35384);
or U36007 (N_36007,N_35020,N_35915);
or U36008 (N_36008,N_35909,N_35159);
xor U36009 (N_36009,N_35072,N_35837);
nand U36010 (N_36010,N_35274,N_35235);
nand U36011 (N_36011,N_35737,N_35347);
nand U36012 (N_36012,N_35258,N_35393);
nor U36013 (N_36013,N_35764,N_35865);
xnor U36014 (N_36014,N_35942,N_35057);
nor U36015 (N_36015,N_35894,N_35316);
nor U36016 (N_36016,N_35838,N_35046);
nand U36017 (N_36017,N_35937,N_35167);
xor U36018 (N_36018,N_35553,N_35994);
nand U36019 (N_36019,N_35705,N_35310);
xnor U36020 (N_36020,N_35702,N_35355);
or U36021 (N_36021,N_35052,N_35125);
nand U36022 (N_36022,N_35924,N_35630);
or U36023 (N_36023,N_35219,N_35993);
nor U36024 (N_36024,N_35759,N_35058);
or U36025 (N_36025,N_35950,N_35366);
and U36026 (N_36026,N_35350,N_35431);
and U36027 (N_36027,N_35189,N_35585);
nand U36028 (N_36028,N_35406,N_35890);
and U36029 (N_36029,N_35628,N_35673);
xor U36030 (N_36030,N_35752,N_35974);
nor U36031 (N_36031,N_35115,N_35076);
nor U36032 (N_36032,N_35417,N_35322);
and U36033 (N_36033,N_35809,N_35439);
or U36034 (N_36034,N_35246,N_35408);
and U36035 (N_36035,N_35889,N_35490);
nor U36036 (N_36036,N_35850,N_35588);
nand U36037 (N_36037,N_35014,N_35063);
xnor U36038 (N_36038,N_35841,N_35044);
or U36039 (N_36039,N_35556,N_35584);
and U36040 (N_36040,N_35469,N_35681);
xnor U36041 (N_36041,N_35527,N_35970);
nand U36042 (N_36042,N_35626,N_35342);
xnor U36043 (N_36043,N_35707,N_35543);
xnor U36044 (N_36044,N_35339,N_35065);
nand U36045 (N_36045,N_35908,N_35664);
xnor U36046 (N_36046,N_35639,N_35882);
or U36047 (N_36047,N_35242,N_35257);
xor U36048 (N_36048,N_35097,N_35564);
nand U36049 (N_36049,N_35031,N_35933);
nand U36050 (N_36050,N_35206,N_35305);
xnor U36051 (N_36051,N_35609,N_35738);
and U36052 (N_36052,N_35212,N_35188);
nand U36053 (N_36053,N_35625,N_35565);
nor U36054 (N_36054,N_35874,N_35656);
or U36055 (N_36055,N_35094,N_35581);
xnor U36056 (N_36056,N_35800,N_35567);
or U36057 (N_36057,N_35208,N_35637);
xor U36058 (N_36058,N_35353,N_35158);
or U36059 (N_36059,N_35215,N_35443);
nand U36060 (N_36060,N_35716,N_35884);
xor U36061 (N_36061,N_35574,N_35592);
nand U36062 (N_36062,N_35317,N_35922);
or U36063 (N_36063,N_35859,N_35757);
xor U36064 (N_36064,N_35613,N_35096);
or U36065 (N_36065,N_35533,N_35444);
or U36066 (N_36066,N_35708,N_35419);
and U36067 (N_36067,N_35436,N_35943);
xor U36068 (N_36068,N_35591,N_35677);
nor U36069 (N_36069,N_35853,N_35328);
nor U36070 (N_36070,N_35216,N_35260);
nand U36071 (N_36071,N_35992,N_35712);
nand U36072 (N_36072,N_35061,N_35765);
nor U36073 (N_36073,N_35109,N_35751);
nand U36074 (N_36074,N_35135,N_35121);
nor U36075 (N_36075,N_35418,N_35524);
xor U36076 (N_36076,N_35615,N_35810);
nand U36077 (N_36077,N_35866,N_35801);
xnor U36078 (N_36078,N_35166,N_35228);
and U36079 (N_36079,N_35079,N_35641);
nor U36080 (N_36080,N_35648,N_35006);
and U36081 (N_36081,N_35936,N_35197);
nor U36082 (N_36082,N_35341,N_35666);
or U36083 (N_36083,N_35761,N_35259);
or U36084 (N_36084,N_35361,N_35817);
nand U36085 (N_36085,N_35217,N_35042);
and U36086 (N_36086,N_35678,N_35023);
nor U36087 (N_36087,N_35939,N_35163);
and U36088 (N_36088,N_35461,N_35119);
or U36089 (N_36089,N_35780,N_35411);
and U36090 (N_36090,N_35221,N_35794);
or U36091 (N_36091,N_35855,N_35149);
and U36092 (N_36092,N_35458,N_35851);
or U36093 (N_36093,N_35644,N_35518);
nand U36094 (N_36094,N_35815,N_35991);
or U36095 (N_36095,N_35398,N_35498);
or U36096 (N_36096,N_35263,N_35231);
or U36097 (N_36097,N_35016,N_35289);
or U36098 (N_36098,N_35802,N_35364);
nor U36099 (N_36099,N_35291,N_35665);
and U36100 (N_36100,N_35004,N_35110);
xor U36101 (N_36101,N_35963,N_35025);
or U36102 (N_36102,N_35961,N_35966);
nand U36103 (N_36103,N_35368,N_35725);
xnor U36104 (N_36104,N_35488,N_35912);
and U36105 (N_36105,N_35396,N_35831);
and U36106 (N_36106,N_35168,N_35252);
and U36107 (N_36107,N_35338,N_35485);
and U36108 (N_36108,N_35179,N_35248);
nand U36109 (N_36109,N_35336,N_35139);
nor U36110 (N_36110,N_35938,N_35494);
or U36111 (N_36111,N_35561,N_35595);
xor U36112 (N_36112,N_35845,N_35369);
nand U36113 (N_36113,N_35710,N_35477);
xor U36114 (N_36114,N_35551,N_35027);
or U36115 (N_36115,N_35714,N_35978);
and U36116 (N_36116,N_35806,N_35886);
or U36117 (N_36117,N_35798,N_35253);
xor U36118 (N_36118,N_35534,N_35753);
or U36119 (N_36119,N_35539,N_35165);
nand U36120 (N_36120,N_35335,N_35946);
or U36121 (N_36121,N_35391,N_35367);
nor U36122 (N_36122,N_35271,N_35050);
or U36123 (N_36123,N_35875,N_35337);
nand U36124 (N_36124,N_35969,N_35222);
and U36125 (N_36125,N_35812,N_35241);
nand U36126 (N_36126,N_35460,N_35797);
and U36127 (N_36127,N_35985,N_35173);
nor U36128 (N_36128,N_35990,N_35586);
nor U36129 (N_36129,N_35559,N_35114);
nor U36130 (N_36130,N_35500,N_35577);
or U36131 (N_36131,N_35261,N_35399);
xnor U36132 (N_36132,N_35605,N_35611);
nand U36133 (N_36133,N_35086,N_35190);
nor U36134 (N_36134,N_35566,N_35388);
nand U36135 (N_36135,N_35148,N_35576);
xnor U36136 (N_36136,N_35486,N_35186);
nor U36137 (N_36137,N_35295,N_35447);
xnor U36138 (N_36138,N_35734,N_35784);
xnor U36139 (N_36139,N_35402,N_35818);
nor U36140 (N_36140,N_35923,N_35684);
nor U36141 (N_36141,N_35251,N_35315);
or U36142 (N_36142,N_35124,N_35122);
or U36143 (N_36143,N_35285,N_35001);
xor U36144 (N_36144,N_35021,N_35715);
or U36145 (N_36145,N_35441,N_35624);
xor U36146 (N_36146,N_35713,N_35918);
nor U36147 (N_36147,N_35863,N_35265);
xor U36148 (N_36148,N_35778,N_35579);
and U36149 (N_36149,N_35767,N_35535);
nor U36150 (N_36150,N_35421,N_35662);
and U36151 (N_36151,N_35839,N_35789);
xnor U36152 (N_36152,N_35857,N_35155);
nor U36153 (N_36153,N_35298,N_35313);
nand U36154 (N_36154,N_35704,N_35196);
or U36155 (N_36155,N_35520,N_35594);
and U36156 (N_36156,N_35073,N_35379);
nand U36157 (N_36157,N_35226,N_35404);
and U36158 (N_36158,N_35523,N_35203);
or U36159 (N_36159,N_35998,N_35776);
and U36160 (N_36160,N_35876,N_35960);
or U36161 (N_36161,N_35358,N_35528);
and U36162 (N_36162,N_35348,N_35959);
or U36163 (N_36163,N_35371,N_35468);
or U36164 (N_36164,N_35452,N_35036);
xor U36165 (N_36165,N_35980,N_35955);
and U36166 (N_36166,N_35779,N_35278);
and U36167 (N_36167,N_35878,N_35239);
nand U36168 (N_36168,N_35948,N_35842);
nand U36169 (N_36169,N_35092,N_35957);
xor U36170 (N_36170,N_35682,N_35464);
or U36171 (N_36171,N_35746,N_35049);
nor U36172 (N_36172,N_35964,N_35056);
xor U36173 (N_36173,N_35563,N_35277);
xnor U36174 (N_36174,N_35113,N_35899);
nor U36175 (N_36175,N_35038,N_35123);
nand U36176 (N_36176,N_35293,N_35634);
xor U36177 (N_36177,N_35223,N_35856);
nor U36178 (N_36178,N_35496,N_35552);
nor U36179 (N_36179,N_35652,N_35267);
nand U36180 (N_36180,N_35499,N_35996);
nor U36181 (N_36181,N_35803,N_35299);
and U36182 (N_36182,N_35238,N_35141);
nand U36183 (N_36183,N_35733,N_35679);
nor U36184 (N_36184,N_35562,N_35078);
xor U36185 (N_36185,N_35438,N_35979);
nor U36186 (N_36186,N_35037,N_35510);
and U36187 (N_36187,N_35583,N_35034);
or U36188 (N_36188,N_35053,N_35157);
nor U36189 (N_36189,N_35844,N_35146);
nor U36190 (N_36190,N_35651,N_35758);
nand U36191 (N_36191,N_35156,N_35516);
and U36192 (N_36192,N_35944,N_35827);
xnor U36193 (N_36193,N_35284,N_35007);
or U36194 (N_36194,N_35470,N_35286);
nor U36195 (N_36195,N_35687,N_35300);
or U36196 (N_36196,N_35296,N_35781);
nand U36197 (N_36197,N_35442,N_35871);
or U36198 (N_36198,N_35608,N_35280);
nand U36199 (N_36199,N_35279,N_35306);
and U36200 (N_36200,N_35133,N_35127);
and U36201 (N_36201,N_35329,N_35422);
nand U36202 (N_36202,N_35319,N_35549);
xnor U36203 (N_36203,N_35104,N_35653);
and U36204 (N_36204,N_35169,N_35675);
nor U36205 (N_36205,N_35249,N_35836);
nor U36206 (N_36206,N_35193,N_35770);
xor U36207 (N_36207,N_35420,N_35088);
xnor U36208 (N_36208,N_35308,N_35268);
or U36209 (N_36209,N_35723,N_35640);
or U36210 (N_36210,N_35578,N_35795);
or U36211 (N_36211,N_35103,N_35914);
xnor U36212 (N_36212,N_35935,N_35791);
and U36213 (N_36213,N_35917,N_35724);
nand U36214 (N_36214,N_35198,N_35105);
nor U36215 (N_36215,N_35854,N_35243);
or U36216 (N_36216,N_35101,N_35976);
nor U36217 (N_36217,N_35731,N_35895);
or U36218 (N_36218,N_35082,N_35349);
nor U36219 (N_36219,N_35112,N_35068);
or U36220 (N_36220,N_35275,N_35126);
or U36221 (N_36221,N_35823,N_35668);
and U36222 (N_36222,N_35230,N_35987);
or U36223 (N_36223,N_35320,N_35927);
nor U36224 (N_36224,N_35560,N_35425);
or U36225 (N_36225,N_35476,N_35968);
nor U36226 (N_36226,N_35493,N_35698);
and U36227 (N_36227,N_35254,N_35748);
nand U36228 (N_36228,N_35352,N_35544);
and U36229 (N_36229,N_35389,N_35849);
nor U36230 (N_36230,N_35692,N_35981);
or U36231 (N_36231,N_35686,N_35497);
and U36232 (N_36232,N_35192,N_35582);
and U36233 (N_36233,N_35432,N_35603);
nor U36234 (N_36234,N_35487,N_35676);
or U36235 (N_36235,N_35846,N_35290);
and U36236 (N_36236,N_35106,N_35433);
nand U36237 (N_36237,N_35210,N_35786);
nor U36238 (N_36238,N_35473,N_35318);
nor U36239 (N_36239,N_35897,N_35184);
and U36240 (N_36240,N_35906,N_35934);
and U36241 (N_36241,N_35722,N_35995);
xor U36242 (N_36242,N_35330,N_35085);
xnor U36243 (N_36243,N_35726,N_35018);
and U36244 (N_36244,N_35357,N_35180);
and U36245 (N_36245,N_35736,N_35554);
nor U36246 (N_36246,N_35550,N_35202);
nor U36247 (N_36247,N_35382,N_35256);
nor U36248 (N_36248,N_35824,N_35598);
xor U36249 (N_36249,N_35587,N_35893);
nor U36250 (N_36250,N_35035,N_35743);
nor U36251 (N_36251,N_35233,N_35521);
nor U36252 (N_36252,N_35898,N_35907);
nor U36253 (N_36253,N_35445,N_35401);
and U36254 (N_36254,N_35825,N_35182);
xnor U36255 (N_36255,N_35919,N_35526);
nor U36256 (N_36256,N_35170,N_35941);
or U36257 (N_36257,N_35448,N_35953);
nand U36258 (N_36258,N_35091,N_35136);
xor U36259 (N_36259,N_35858,N_35482);
xor U36260 (N_36260,N_35301,N_35397);
and U36261 (N_36261,N_35245,N_35606);
or U36262 (N_36262,N_35504,N_35083);
or U36263 (N_36263,N_35129,N_35832);
nand U36264 (N_36264,N_35973,N_35346);
and U36265 (N_36265,N_35931,N_35896);
or U36266 (N_36266,N_35428,N_35360);
or U36267 (N_36267,N_35947,N_35162);
nor U36268 (N_36268,N_35808,N_35555);
xor U36269 (N_36269,N_35024,N_35569);
xor U36270 (N_36270,N_35775,N_35672);
and U36271 (N_36271,N_35390,N_35616);
nor U36272 (N_36272,N_35478,N_35449);
and U36273 (N_36273,N_35822,N_35392);
nand U36274 (N_36274,N_35660,N_35735);
and U36275 (N_36275,N_35654,N_35745);
xor U36276 (N_36276,N_35043,N_35719);
nor U36277 (N_36277,N_35793,N_35062);
and U36278 (N_36278,N_35940,N_35272);
nand U36279 (N_36279,N_35760,N_35099);
or U36280 (N_36280,N_35374,N_35536);
and U36281 (N_36281,N_35787,N_35029);
or U36282 (N_36282,N_35040,N_35153);
nand U36283 (N_36283,N_35607,N_35768);
nand U36284 (N_36284,N_35811,N_35191);
and U36285 (N_36285,N_35887,N_35281);
xor U36286 (N_36286,N_35209,N_35694);
and U36287 (N_36287,N_35828,N_35773);
nand U36288 (N_36288,N_35227,N_35790);
xnor U36289 (N_36289,N_35814,N_35171);
and U36290 (N_36290,N_35632,N_35711);
nand U36291 (N_36291,N_35385,N_35459);
nor U36292 (N_36292,N_35325,N_35636);
xor U36293 (N_36293,N_35376,N_35916);
xor U36294 (N_36294,N_35883,N_35028);
nand U36295 (N_36295,N_35143,N_35604);
nand U36296 (N_36296,N_35843,N_35309);
xnor U36297 (N_36297,N_35701,N_35690);
or U36298 (N_36298,N_35984,N_35932);
nand U36299 (N_36299,N_35283,N_35834);
or U36300 (N_36300,N_35766,N_35532);
xor U36301 (N_36301,N_35334,N_35455);
nor U36302 (N_36302,N_35982,N_35807);
or U36303 (N_36303,N_35292,N_35517);
and U36304 (N_36304,N_35152,N_35059);
nor U36305 (N_36305,N_35650,N_35688);
xor U36306 (N_36306,N_35276,N_35580);
or U36307 (N_36307,N_35395,N_35160);
xor U36308 (N_36308,N_35323,N_35066);
and U36309 (N_36309,N_35548,N_35945);
nand U36310 (N_36310,N_35891,N_35879);
xnor U36311 (N_36311,N_35225,N_35833);
nand U36312 (N_36312,N_35304,N_35363);
nand U36313 (N_36313,N_35718,N_35120);
nand U36314 (N_36314,N_35989,N_35479);
xor U36315 (N_36315,N_35728,N_35176);
and U36316 (N_36316,N_35645,N_35804);
nand U36317 (N_36317,N_35375,N_35491);
nand U36318 (N_36318,N_35207,N_35199);
xnor U36319 (N_36319,N_35282,N_35589);
and U36320 (N_36320,N_35905,N_35568);
or U36321 (N_36321,N_35703,N_35172);
or U36322 (N_36322,N_35696,N_35695);
and U36323 (N_36323,N_35032,N_35819);
nor U36324 (N_36324,N_35343,N_35685);
and U36325 (N_36325,N_35080,N_35740);
or U36326 (N_36326,N_35739,N_35416);
and U36327 (N_36327,N_35506,N_35920);
and U36328 (N_36328,N_35467,N_35185);
nand U36329 (N_36329,N_35456,N_35400);
nand U36330 (N_36330,N_35255,N_35394);
or U36331 (N_36331,N_35671,N_35505);
or U36332 (N_36332,N_35312,N_35900);
xnor U36333 (N_36333,N_35847,N_35003);
nand U36334 (N_36334,N_35132,N_35010);
xnor U36335 (N_36335,N_35659,N_35575);
nand U36336 (N_36336,N_35547,N_35314);
and U36337 (N_36337,N_35674,N_35638);
nor U36338 (N_36338,N_35087,N_35509);
or U36339 (N_36339,N_35426,N_35596);
and U36340 (N_36340,N_35297,N_35952);
and U36341 (N_36341,N_35002,N_35423);
nor U36342 (N_36342,N_35649,N_35055);
or U36343 (N_36343,N_35623,N_35415);
or U36344 (N_36344,N_35084,N_35511);
or U36345 (N_36345,N_35631,N_35244);
nor U36346 (N_36346,N_35144,N_35741);
nor U36347 (N_36347,N_35039,N_35434);
and U36348 (N_36348,N_35011,N_35888);
nor U36349 (N_36349,N_35796,N_35457);
nand U36350 (N_36350,N_35820,N_35570);
nor U36351 (N_36351,N_35344,N_35345);
xor U36352 (N_36352,N_35558,N_35204);
and U36353 (N_36353,N_35700,N_35921);
and U36354 (N_36354,N_35977,N_35747);
or U36355 (N_36355,N_35151,N_35287);
or U36356 (N_36356,N_35545,N_35669);
or U36357 (N_36357,N_35154,N_35930);
xnor U36358 (N_36358,N_35147,N_35194);
nand U36359 (N_36359,N_35880,N_35840);
nand U36360 (N_36360,N_35601,N_35481);
or U36361 (N_36361,N_35904,N_35512);
or U36362 (N_36362,N_35093,N_35502);
and U36363 (N_36363,N_35872,N_35060);
nand U36364 (N_36364,N_35689,N_35326);
nand U36365 (N_36365,N_35627,N_35128);
xor U36366 (N_36366,N_35683,N_35546);
xor U36367 (N_36367,N_35373,N_35514);
nand U36368 (N_36368,N_35064,N_35492);
nor U36369 (N_36369,N_35174,N_35635);
xnor U36370 (N_36370,N_35463,N_35999);
xor U36371 (N_36371,N_35612,N_35100);
nor U36372 (N_36372,N_35471,N_35250);
and U36373 (N_36373,N_35030,N_35571);
and U36374 (N_36374,N_35962,N_35372);
nor U36375 (N_36375,N_35015,N_35264);
nand U36376 (N_36376,N_35706,N_35540);
nand U36377 (N_36377,N_35911,N_35680);
xnor U36378 (N_36378,N_35116,N_35717);
or U36379 (N_36379,N_35177,N_35307);
or U36380 (N_36380,N_35381,N_35538);
xnor U36381 (N_36381,N_35663,N_35183);
xnor U36382 (N_36382,N_35466,N_35699);
and U36383 (N_36383,N_35885,N_35519);
nand U36384 (N_36384,N_35232,N_35410);
and U36385 (N_36385,N_35691,N_35597);
xor U36386 (N_36386,N_35513,N_35214);
nor U36387 (N_36387,N_35118,N_35067);
and U36388 (N_36388,N_35860,N_35573);
nor U36389 (N_36389,N_35483,N_35412);
xnor U36390 (N_36390,N_35075,N_35771);
and U36391 (N_36391,N_35387,N_35529);
xnor U36392 (N_36392,N_35359,N_35413);
and U36393 (N_36393,N_35835,N_35266);
or U36394 (N_36394,N_35829,N_35769);
or U36395 (N_36395,N_35218,N_35137);
nor U36396 (N_36396,N_35774,N_35095);
nand U36397 (N_36397,N_35629,N_35848);
nor U36398 (N_36398,N_35403,N_35557);
or U36399 (N_36399,N_35220,N_35967);
nor U36400 (N_36400,N_35142,N_35508);
nand U36401 (N_36401,N_35195,N_35537);
or U36402 (N_36402,N_35792,N_35187);
and U36403 (N_36403,N_35910,N_35600);
and U36404 (N_36404,N_35356,N_35622);
and U36405 (N_36405,N_35542,N_35019);
and U36406 (N_36406,N_35785,N_35643);
nor U36407 (N_36407,N_35777,N_35958);
nand U36408 (N_36408,N_35409,N_35380);
or U36409 (N_36409,N_35045,N_35178);
xor U36410 (N_36410,N_35805,N_35236);
nor U36411 (N_36411,N_35429,N_35224);
and U36412 (N_36412,N_35107,N_35211);
and U36413 (N_36413,N_35017,N_35756);
nand U36414 (N_36414,N_35435,N_35614);
or U36415 (N_36415,N_35599,N_35997);
and U36416 (N_36416,N_35852,N_35971);
or U36417 (N_36417,N_35619,N_35437);
and U36418 (N_36418,N_35200,N_35503);
xnor U36419 (N_36419,N_35873,N_35269);
or U36420 (N_36420,N_35414,N_35424);
or U36421 (N_36421,N_35054,N_35134);
nand U36422 (N_36422,N_35729,N_35005);
nand U36423 (N_36423,N_35454,N_35321);
xnor U36424 (N_36424,N_35929,N_35140);
nand U36425 (N_36425,N_35730,N_35090);
or U36426 (N_36426,N_35440,N_35720);
nor U36427 (N_36427,N_35864,N_35181);
or U36428 (N_36428,N_35572,N_35446);
nand U36429 (N_36429,N_35928,N_35288);
xor U36430 (N_36430,N_35138,N_35262);
and U36431 (N_36431,N_35877,N_35525);
nand U36432 (N_36432,N_35332,N_35130);
or U36433 (N_36433,N_35826,N_35324);
xnor U36434 (N_36434,N_35727,N_35378);
nand U36435 (N_36435,N_35453,N_35495);
or U36436 (N_36436,N_35522,N_35175);
and U36437 (N_36437,N_35273,N_35229);
and U36438 (N_36438,N_35489,N_35772);
and U36439 (N_36439,N_35047,N_35697);
nor U36440 (N_36440,N_35145,N_35237);
and U36441 (N_36441,N_35213,N_35474);
or U36442 (N_36442,N_35762,N_35642);
or U36443 (N_36443,N_35507,N_35407);
or U36444 (N_36444,N_35484,N_35658);
or U36445 (N_36445,N_35867,N_35670);
or U36446 (N_36446,N_35541,N_35161);
xnor U36447 (N_36447,N_35881,N_35340);
xnor U36448 (N_36448,N_35531,N_35972);
nor U36449 (N_36449,N_35041,N_35475);
or U36450 (N_36450,N_35012,N_35633);
nor U36451 (N_36451,N_35618,N_35164);
and U36452 (N_36452,N_35647,N_35732);
nor U36453 (N_36453,N_35763,N_35013);
nand U36454 (N_36454,N_35892,N_35755);
nor U36455 (N_36455,N_35026,N_35870);
nand U36456 (N_36456,N_35365,N_35081);
xor U36457 (N_36457,N_35926,N_35988);
or U36458 (N_36458,N_35131,N_35754);
nand U36459 (N_36459,N_35102,N_35515);
or U36460 (N_36460,N_35377,N_35000);
and U36461 (N_36461,N_35362,N_35386);
or U36462 (N_36462,N_35783,N_35721);
and U36463 (N_36463,N_35693,N_35048);
xnor U36464 (N_36464,N_35901,N_35830);
and U36465 (N_36465,N_35351,N_35480);
and U36466 (N_36466,N_35465,N_35709);
xor U36467 (N_36467,N_35451,N_35861);
xnor U36468 (N_36468,N_35744,N_35667);
xnor U36469 (N_36469,N_35333,N_35621);
and U36470 (N_36470,N_35108,N_35077);
nor U36471 (N_36471,N_35240,N_35370);
nand U36472 (N_36472,N_35098,N_35590);
nor U36473 (N_36473,N_35022,N_35247);
nor U36474 (N_36474,N_35902,N_35799);
and U36475 (N_36475,N_35813,N_35788);
and U36476 (N_36476,N_35593,N_35951);
and U36477 (N_36477,N_35986,N_35617);
or U36478 (N_36478,N_35331,N_35327);
nor U36479 (N_36479,N_35009,N_35965);
nor U36480 (N_36480,N_35205,N_35954);
or U36481 (N_36481,N_35869,N_35956);
nand U36482 (N_36482,N_35816,N_35913);
and U36483 (N_36483,N_35405,N_35983);
nor U36484 (N_36484,N_35302,N_35462);
xor U36485 (N_36485,N_35117,N_35657);
or U36486 (N_36486,N_35270,N_35742);
nand U36487 (N_36487,N_35821,N_35089);
nand U36488 (N_36488,N_35071,N_35655);
or U36489 (N_36489,N_35430,N_35111);
or U36490 (N_36490,N_35234,N_35074);
nand U36491 (N_36491,N_35868,N_35925);
nand U36492 (N_36492,N_35782,N_35749);
nand U36493 (N_36493,N_35051,N_35750);
or U36494 (N_36494,N_35070,N_35501);
nand U36495 (N_36495,N_35303,N_35610);
nor U36496 (N_36496,N_35294,N_35311);
nor U36497 (N_36497,N_35661,N_35069);
xor U36498 (N_36498,N_35903,N_35949);
nor U36499 (N_36499,N_35201,N_35033);
nor U36500 (N_36500,N_35267,N_35285);
and U36501 (N_36501,N_35719,N_35414);
nor U36502 (N_36502,N_35143,N_35165);
and U36503 (N_36503,N_35178,N_35984);
or U36504 (N_36504,N_35756,N_35370);
or U36505 (N_36505,N_35262,N_35394);
or U36506 (N_36506,N_35905,N_35951);
or U36507 (N_36507,N_35134,N_35092);
and U36508 (N_36508,N_35466,N_35010);
nor U36509 (N_36509,N_35663,N_35117);
or U36510 (N_36510,N_35301,N_35369);
xnor U36511 (N_36511,N_35029,N_35721);
nor U36512 (N_36512,N_35376,N_35682);
or U36513 (N_36513,N_35103,N_35440);
and U36514 (N_36514,N_35921,N_35387);
xor U36515 (N_36515,N_35245,N_35834);
xnor U36516 (N_36516,N_35502,N_35771);
or U36517 (N_36517,N_35023,N_35473);
xor U36518 (N_36518,N_35778,N_35702);
nor U36519 (N_36519,N_35852,N_35301);
nor U36520 (N_36520,N_35200,N_35339);
nor U36521 (N_36521,N_35008,N_35334);
nor U36522 (N_36522,N_35010,N_35845);
nor U36523 (N_36523,N_35657,N_35550);
or U36524 (N_36524,N_35089,N_35512);
nand U36525 (N_36525,N_35705,N_35394);
xnor U36526 (N_36526,N_35429,N_35423);
nand U36527 (N_36527,N_35445,N_35937);
nor U36528 (N_36528,N_35208,N_35232);
nand U36529 (N_36529,N_35955,N_35075);
nand U36530 (N_36530,N_35776,N_35910);
nor U36531 (N_36531,N_35915,N_35002);
and U36532 (N_36532,N_35632,N_35753);
and U36533 (N_36533,N_35324,N_35674);
and U36534 (N_36534,N_35049,N_35908);
xnor U36535 (N_36535,N_35021,N_35861);
nand U36536 (N_36536,N_35373,N_35161);
nand U36537 (N_36537,N_35696,N_35734);
nand U36538 (N_36538,N_35424,N_35168);
nor U36539 (N_36539,N_35734,N_35490);
xnor U36540 (N_36540,N_35191,N_35711);
xor U36541 (N_36541,N_35865,N_35883);
or U36542 (N_36542,N_35326,N_35340);
and U36543 (N_36543,N_35815,N_35023);
nand U36544 (N_36544,N_35080,N_35539);
xor U36545 (N_36545,N_35086,N_35177);
and U36546 (N_36546,N_35140,N_35755);
nor U36547 (N_36547,N_35650,N_35251);
or U36548 (N_36548,N_35150,N_35125);
and U36549 (N_36549,N_35935,N_35371);
or U36550 (N_36550,N_35235,N_35768);
nand U36551 (N_36551,N_35533,N_35359);
nand U36552 (N_36552,N_35016,N_35758);
xor U36553 (N_36553,N_35217,N_35293);
nand U36554 (N_36554,N_35293,N_35226);
xor U36555 (N_36555,N_35059,N_35355);
or U36556 (N_36556,N_35791,N_35482);
xnor U36557 (N_36557,N_35891,N_35331);
and U36558 (N_36558,N_35727,N_35375);
or U36559 (N_36559,N_35233,N_35600);
xor U36560 (N_36560,N_35691,N_35184);
or U36561 (N_36561,N_35432,N_35563);
xnor U36562 (N_36562,N_35950,N_35407);
and U36563 (N_36563,N_35397,N_35522);
nand U36564 (N_36564,N_35174,N_35837);
and U36565 (N_36565,N_35136,N_35427);
nand U36566 (N_36566,N_35563,N_35859);
nand U36567 (N_36567,N_35153,N_35658);
xnor U36568 (N_36568,N_35568,N_35396);
and U36569 (N_36569,N_35137,N_35751);
nand U36570 (N_36570,N_35216,N_35094);
nor U36571 (N_36571,N_35878,N_35407);
or U36572 (N_36572,N_35366,N_35341);
nor U36573 (N_36573,N_35015,N_35573);
and U36574 (N_36574,N_35886,N_35111);
and U36575 (N_36575,N_35673,N_35900);
nor U36576 (N_36576,N_35846,N_35501);
or U36577 (N_36577,N_35551,N_35773);
nor U36578 (N_36578,N_35567,N_35259);
and U36579 (N_36579,N_35321,N_35709);
or U36580 (N_36580,N_35068,N_35840);
or U36581 (N_36581,N_35342,N_35001);
or U36582 (N_36582,N_35107,N_35904);
and U36583 (N_36583,N_35887,N_35201);
nor U36584 (N_36584,N_35379,N_35462);
xnor U36585 (N_36585,N_35202,N_35206);
nand U36586 (N_36586,N_35663,N_35143);
nor U36587 (N_36587,N_35578,N_35215);
nand U36588 (N_36588,N_35986,N_35316);
and U36589 (N_36589,N_35228,N_35034);
nor U36590 (N_36590,N_35631,N_35569);
and U36591 (N_36591,N_35389,N_35884);
nand U36592 (N_36592,N_35237,N_35347);
nand U36593 (N_36593,N_35460,N_35739);
nor U36594 (N_36594,N_35760,N_35217);
nand U36595 (N_36595,N_35272,N_35276);
or U36596 (N_36596,N_35642,N_35435);
nand U36597 (N_36597,N_35948,N_35626);
nor U36598 (N_36598,N_35118,N_35540);
nand U36599 (N_36599,N_35451,N_35701);
xor U36600 (N_36600,N_35797,N_35384);
or U36601 (N_36601,N_35368,N_35958);
nand U36602 (N_36602,N_35912,N_35561);
nand U36603 (N_36603,N_35517,N_35608);
nand U36604 (N_36604,N_35553,N_35590);
nand U36605 (N_36605,N_35027,N_35329);
nand U36606 (N_36606,N_35098,N_35658);
xor U36607 (N_36607,N_35674,N_35261);
and U36608 (N_36608,N_35775,N_35776);
or U36609 (N_36609,N_35232,N_35671);
and U36610 (N_36610,N_35092,N_35280);
nand U36611 (N_36611,N_35482,N_35911);
xnor U36612 (N_36612,N_35630,N_35348);
nand U36613 (N_36613,N_35216,N_35991);
nand U36614 (N_36614,N_35142,N_35139);
and U36615 (N_36615,N_35927,N_35842);
and U36616 (N_36616,N_35380,N_35316);
nand U36617 (N_36617,N_35449,N_35479);
or U36618 (N_36618,N_35126,N_35774);
nand U36619 (N_36619,N_35242,N_35503);
xor U36620 (N_36620,N_35996,N_35409);
nor U36621 (N_36621,N_35102,N_35174);
and U36622 (N_36622,N_35607,N_35076);
xnor U36623 (N_36623,N_35777,N_35647);
and U36624 (N_36624,N_35859,N_35966);
nor U36625 (N_36625,N_35944,N_35937);
nor U36626 (N_36626,N_35826,N_35676);
or U36627 (N_36627,N_35636,N_35793);
nand U36628 (N_36628,N_35802,N_35607);
or U36629 (N_36629,N_35494,N_35631);
or U36630 (N_36630,N_35319,N_35891);
nor U36631 (N_36631,N_35418,N_35602);
xor U36632 (N_36632,N_35589,N_35881);
nand U36633 (N_36633,N_35613,N_35305);
or U36634 (N_36634,N_35123,N_35448);
xor U36635 (N_36635,N_35567,N_35242);
nor U36636 (N_36636,N_35741,N_35603);
and U36637 (N_36637,N_35352,N_35033);
xor U36638 (N_36638,N_35019,N_35859);
and U36639 (N_36639,N_35926,N_35964);
nand U36640 (N_36640,N_35830,N_35207);
xnor U36641 (N_36641,N_35731,N_35154);
nor U36642 (N_36642,N_35951,N_35612);
xor U36643 (N_36643,N_35868,N_35250);
xor U36644 (N_36644,N_35537,N_35909);
nor U36645 (N_36645,N_35078,N_35340);
and U36646 (N_36646,N_35522,N_35740);
and U36647 (N_36647,N_35806,N_35504);
nand U36648 (N_36648,N_35594,N_35887);
xor U36649 (N_36649,N_35428,N_35180);
nand U36650 (N_36650,N_35172,N_35710);
and U36651 (N_36651,N_35859,N_35167);
nor U36652 (N_36652,N_35784,N_35637);
nand U36653 (N_36653,N_35964,N_35861);
nor U36654 (N_36654,N_35121,N_35727);
and U36655 (N_36655,N_35409,N_35612);
or U36656 (N_36656,N_35330,N_35777);
or U36657 (N_36657,N_35572,N_35401);
or U36658 (N_36658,N_35239,N_35165);
or U36659 (N_36659,N_35495,N_35540);
xor U36660 (N_36660,N_35575,N_35965);
xnor U36661 (N_36661,N_35229,N_35677);
xnor U36662 (N_36662,N_35315,N_35064);
or U36663 (N_36663,N_35089,N_35689);
and U36664 (N_36664,N_35622,N_35837);
or U36665 (N_36665,N_35188,N_35137);
nand U36666 (N_36666,N_35511,N_35052);
and U36667 (N_36667,N_35996,N_35952);
or U36668 (N_36668,N_35990,N_35931);
and U36669 (N_36669,N_35838,N_35117);
xor U36670 (N_36670,N_35822,N_35673);
xnor U36671 (N_36671,N_35540,N_35184);
and U36672 (N_36672,N_35836,N_35073);
xor U36673 (N_36673,N_35733,N_35254);
xor U36674 (N_36674,N_35747,N_35473);
xor U36675 (N_36675,N_35547,N_35430);
xor U36676 (N_36676,N_35244,N_35769);
nand U36677 (N_36677,N_35646,N_35604);
xor U36678 (N_36678,N_35803,N_35915);
xor U36679 (N_36679,N_35219,N_35774);
xnor U36680 (N_36680,N_35129,N_35188);
xnor U36681 (N_36681,N_35768,N_35075);
or U36682 (N_36682,N_35860,N_35299);
and U36683 (N_36683,N_35847,N_35942);
xnor U36684 (N_36684,N_35774,N_35695);
and U36685 (N_36685,N_35171,N_35013);
and U36686 (N_36686,N_35562,N_35437);
nand U36687 (N_36687,N_35878,N_35789);
or U36688 (N_36688,N_35560,N_35000);
or U36689 (N_36689,N_35729,N_35426);
nor U36690 (N_36690,N_35185,N_35629);
or U36691 (N_36691,N_35388,N_35523);
nor U36692 (N_36692,N_35390,N_35145);
and U36693 (N_36693,N_35039,N_35287);
xor U36694 (N_36694,N_35837,N_35537);
nor U36695 (N_36695,N_35915,N_35533);
nand U36696 (N_36696,N_35851,N_35487);
nor U36697 (N_36697,N_35753,N_35019);
xor U36698 (N_36698,N_35695,N_35372);
and U36699 (N_36699,N_35253,N_35032);
xnor U36700 (N_36700,N_35195,N_35275);
or U36701 (N_36701,N_35084,N_35440);
nand U36702 (N_36702,N_35731,N_35583);
and U36703 (N_36703,N_35034,N_35489);
nand U36704 (N_36704,N_35527,N_35508);
nand U36705 (N_36705,N_35510,N_35423);
and U36706 (N_36706,N_35397,N_35155);
and U36707 (N_36707,N_35751,N_35527);
xor U36708 (N_36708,N_35274,N_35998);
and U36709 (N_36709,N_35456,N_35033);
xor U36710 (N_36710,N_35001,N_35480);
xnor U36711 (N_36711,N_35754,N_35592);
xor U36712 (N_36712,N_35214,N_35658);
xnor U36713 (N_36713,N_35321,N_35233);
nor U36714 (N_36714,N_35846,N_35785);
nand U36715 (N_36715,N_35605,N_35220);
nand U36716 (N_36716,N_35862,N_35452);
or U36717 (N_36717,N_35938,N_35829);
and U36718 (N_36718,N_35624,N_35292);
xor U36719 (N_36719,N_35747,N_35484);
and U36720 (N_36720,N_35477,N_35062);
nand U36721 (N_36721,N_35075,N_35284);
nand U36722 (N_36722,N_35628,N_35247);
or U36723 (N_36723,N_35108,N_35397);
nor U36724 (N_36724,N_35282,N_35639);
and U36725 (N_36725,N_35447,N_35336);
nor U36726 (N_36726,N_35582,N_35552);
xor U36727 (N_36727,N_35750,N_35710);
xor U36728 (N_36728,N_35552,N_35056);
xor U36729 (N_36729,N_35544,N_35685);
nor U36730 (N_36730,N_35168,N_35714);
nor U36731 (N_36731,N_35863,N_35277);
nor U36732 (N_36732,N_35897,N_35577);
nor U36733 (N_36733,N_35166,N_35557);
nand U36734 (N_36734,N_35842,N_35894);
and U36735 (N_36735,N_35450,N_35776);
nor U36736 (N_36736,N_35083,N_35716);
or U36737 (N_36737,N_35698,N_35724);
and U36738 (N_36738,N_35407,N_35148);
nand U36739 (N_36739,N_35072,N_35915);
or U36740 (N_36740,N_35753,N_35888);
xor U36741 (N_36741,N_35994,N_35607);
xnor U36742 (N_36742,N_35219,N_35594);
xnor U36743 (N_36743,N_35683,N_35219);
nor U36744 (N_36744,N_35315,N_35437);
and U36745 (N_36745,N_35687,N_35865);
and U36746 (N_36746,N_35766,N_35797);
nor U36747 (N_36747,N_35296,N_35099);
xnor U36748 (N_36748,N_35898,N_35451);
and U36749 (N_36749,N_35631,N_35498);
nand U36750 (N_36750,N_35642,N_35292);
or U36751 (N_36751,N_35218,N_35110);
nand U36752 (N_36752,N_35837,N_35742);
or U36753 (N_36753,N_35759,N_35435);
nor U36754 (N_36754,N_35653,N_35171);
nor U36755 (N_36755,N_35590,N_35606);
nand U36756 (N_36756,N_35492,N_35427);
nor U36757 (N_36757,N_35690,N_35895);
xnor U36758 (N_36758,N_35228,N_35206);
xnor U36759 (N_36759,N_35315,N_35284);
nand U36760 (N_36760,N_35659,N_35385);
nand U36761 (N_36761,N_35306,N_35495);
nor U36762 (N_36762,N_35740,N_35551);
nand U36763 (N_36763,N_35402,N_35447);
nand U36764 (N_36764,N_35121,N_35813);
and U36765 (N_36765,N_35487,N_35371);
xnor U36766 (N_36766,N_35045,N_35786);
or U36767 (N_36767,N_35899,N_35712);
and U36768 (N_36768,N_35967,N_35064);
and U36769 (N_36769,N_35350,N_35107);
xnor U36770 (N_36770,N_35965,N_35579);
xnor U36771 (N_36771,N_35422,N_35882);
and U36772 (N_36772,N_35104,N_35912);
or U36773 (N_36773,N_35729,N_35285);
nand U36774 (N_36774,N_35013,N_35949);
or U36775 (N_36775,N_35335,N_35562);
nor U36776 (N_36776,N_35574,N_35992);
nor U36777 (N_36777,N_35039,N_35342);
xor U36778 (N_36778,N_35743,N_35356);
nand U36779 (N_36779,N_35574,N_35419);
nor U36780 (N_36780,N_35323,N_35985);
and U36781 (N_36781,N_35993,N_35850);
nor U36782 (N_36782,N_35477,N_35709);
nor U36783 (N_36783,N_35857,N_35044);
or U36784 (N_36784,N_35067,N_35601);
and U36785 (N_36785,N_35828,N_35006);
nor U36786 (N_36786,N_35114,N_35014);
and U36787 (N_36787,N_35026,N_35532);
nor U36788 (N_36788,N_35713,N_35395);
nor U36789 (N_36789,N_35925,N_35102);
nor U36790 (N_36790,N_35828,N_35863);
nand U36791 (N_36791,N_35930,N_35947);
and U36792 (N_36792,N_35835,N_35696);
xnor U36793 (N_36793,N_35803,N_35702);
nor U36794 (N_36794,N_35778,N_35522);
and U36795 (N_36795,N_35806,N_35784);
nor U36796 (N_36796,N_35896,N_35595);
xor U36797 (N_36797,N_35249,N_35701);
nand U36798 (N_36798,N_35840,N_35245);
nor U36799 (N_36799,N_35961,N_35725);
nor U36800 (N_36800,N_35026,N_35200);
xor U36801 (N_36801,N_35158,N_35575);
xor U36802 (N_36802,N_35939,N_35848);
and U36803 (N_36803,N_35438,N_35901);
xnor U36804 (N_36804,N_35242,N_35085);
nand U36805 (N_36805,N_35453,N_35587);
xor U36806 (N_36806,N_35042,N_35636);
nor U36807 (N_36807,N_35267,N_35912);
nand U36808 (N_36808,N_35041,N_35102);
or U36809 (N_36809,N_35114,N_35881);
nand U36810 (N_36810,N_35230,N_35228);
and U36811 (N_36811,N_35526,N_35202);
nand U36812 (N_36812,N_35025,N_35183);
and U36813 (N_36813,N_35345,N_35157);
nor U36814 (N_36814,N_35632,N_35084);
nand U36815 (N_36815,N_35421,N_35925);
nand U36816 (N_36816,N_35837,N_35023);
nand U36817 (N_36817,N_35844,N_35301);
or U36818 (N_36818,N_35037,N_35062);
nand U36819 (N_36819,N_35365,N_35785);
or U36820 (N_36820,N_35091,N_35445);
or U36821 (N_36821,N_35269,N_35412);
and U36822 (N_36822,N_35101,N_35201);
and U36823 (N_36823,N_35391,N_35443);
nor U36824 (N_36824,N_35794,N_35743);
or U36825 (N_36825,N_35465,N_35705);
nor U36826 (N_36826,N_35728,N_35265);
or U36827 (N_36827,N_35729,N_35744);
nand U36828 (N_36828,N_35218,N_35922);
nand U36829 (N_36829,N_35642,N_35482);
nand U36830 (N_36830,N_35330,N_35893);
nand U36831 (N_36831,N_35116,N_35881);
nand U36832 (N_36832,N_35853,N_35528);
nand U36833 (N_36833,N_35780,N_35675);
or U36834 (N_36834,N_35513,N_35720);
xor U36835 (N_36835,N_35799,N_35816);
nor U36836 (N_36836,N_35808,N_35222);
nor U36837 (N_36837,N_35539,N_35262);
and U36838 (N_36838,N_35206,N_35218);
nor U36839 (N_36839,N_35514,N_35775);
or U36840 (N_36840,N_35635,N_35433);
and U36841 (N_36841,N_35633,N_35344);
nor U36842 (N_36842,N_35002,N_35470);
and U36843 (N_36843,N_35699,N_35417);
xor U36844 (N_36844,N_35022,N_35974);
and U36845 (N_36845,N_35510,N_35810);
xor U36846 (N_36846,N_35890,N_35803);
xor U36847 (N_36847,N_35729,N_35745);
nor U36848 (N_36848,N_35058,N_35258);
nor U36849 (N_36849,N_35510,N_35222);
nand U36850 (N_36850,N_35803,N_35749);
xor U36851 (N_36851,N_35233,N_35619);
xnor U36852 (N_36852,N_35800,N_35357);
or U36853 (N_36853,N_35799,N_35560);
or U36854 (N_36854,N_35926,N_35139);
and U36855 (N_36855,N_35187,N_35192);
nand U36856 (N_36856,N_35481,N_35321);
nand U36857 (N_36857,N_35875,N_35239);
and U36858 (N_36858,N_35660,N_35734);
nand U36859 (N_36859,N_35617,N_35677);
xor U36860 (N_36860,N_35261,N_35594);
and U36861 (N_36861,N_35253,N_35751);
nor U36862 (N_36862,N_35093,N_35690);
nor U36863 (N_36863,N_35755,N_35105);
xnor U36864 (N_36864,N_35385,N_35533);
xnor U36865 (N_36865,N_35964,N_35921);
nand U36866 (N_36866,N_35598,N_35252);
nor U36867 (N_36867,N_35834,N_35187);
or U36868 (N_36868,N_35352,N_35811);
xnor U36869 (N_36869,N_35672,N_35100);
nor U36870 (N_36870,N_35344,N_35713);
or U36871 (N_36871,N_35249,N_35124);
nand U36872 (N_36872,N_35211,N_35546);
or U36873 (N_36873,N_35536,N_35053);
nand U36874 (N_36874,N_35939,N_35020);
or U36875 (N_36875,N_35470,N_35050);
xnor U36876 (N_36876,N_35012,N_35044);
or U36877 (N_36877,N_35130,N_35885);
nand U36878 (N_36878,N_35948,N_35989);
nand U36879 (N_36879,N_35120,N_35603);
or U36880 (N_36880,N_35258,N_35436);
and U36881 (N_36881,N_35078,N_35109);
or U36882 (N_36882,N_35096,N_35518);
xnor U36883 (N_36883,N_35579,N_35425);
nor U36884 (N_36884,N_35973,N_35671);
nand U36885 (N_36885,N_35624,N_35887);
or U36886 (N_36886,N_35479,N_35638);
or U36887 (N_36887,N_35626,N_35405);
and U36888 (N_36888,N_35944,N_35479);
and U36889 (N_36889,N_35718,N_35398);
or U36890 (N_36890,N_35134,N_35537);
and U36891 (N_36891,N_35513,N_35825);
or U36892 (N_36892,N_35949,N_35506);
or U36893 (N_36893,N_35603,N_35894);
and U36894 (N_36894,N_35070,N_35213);
xor U36895 (N_36895,N_35106,N_35383);
nand U36896 (N_36896,N_35882,N_35116);
xor U36897 (N_36897,N_35548,N_35455);
or U36898 (N_36898,N_35842,N_35670);
xor U36899 (N_36899,N_35022,N_35585);
and U36900 (N_36900,N_35559,N_35883);
or U36901 (N_36901,N_35527,N_35030);
nand U36902 (N_36902,N_35552,N_35786);
xor U36903 (N_36903,N_35595,N_35703);
nand U36904 (N_36904,N_35492,N_35852);
or U36905 (N_36905,N_35047,N_35058);
and U36906 (N_36906,N_35918,N_35108);
nor U36907 (N_36907,N_35987,N_35111);
xnor U36908 (N_36908,N_35077,N_35607);
xor U36909 (N_36909,N_35366,N_35682);
and U36910 (N_36910,N_35819,N_35027);
and U36911 (N_36911,N_35451,N_35506);
or U36912 (N_36912,N_35370,N_35952);
and U36913 (N_36913,N_35024,N_35272);
xnor U36914 (N_36914,N_35888,N_35645);
xor U36915 (N_36915,N_35584,N_35002);
and U36916 (N_36916,N_35145,N_35394);
and U36917 (N_36917,N_35159,N_35623);
or U36918 (N_36918,N_35699,N_35227);
and U36919 (N_36919,N_35585,N_35581);
xor U36920 (N_36920,N_35013,N_35656);
nor U36921 (N_36921,N_35963,N_35576);
nor U36922 (N_36922,N_35381,N_35946);
nor U36923 (N_36923,N_35861,N_35041);
and U36924 (N_36924,N_35411,N_35564);
and U36925 (N_36925,N_35078,N_35234);
and U36926 (N_36926,N_35967,N_35418);
xnor U36927 (N_36927,N_35718,N_35690);
nand U36928 (N_36928,N_35242,N_35582);
xor U36929 (N_36929,N_35603,N_35409);
xnor U36930 (N_36930,N_35617,N_35391);
nand U36931 (N_36931,N_35118,N_35408);
nor U36932 (N_36932,N_35351,N_35826);
nor U36933 (N_36933,N_35797,N_35122);
xor U36934 (N_36934,N_35394,N_35377);
nand U36935 (N_36935,N_35150,N_35877);
nand U36936 (N_36936,N_35770,N_35798);
nand U36937 (N_36937,N_35038,N_35116);
and U36938 (N_36938,N_35891,N_35770);
xnor U36939 (N_36939,N_35051,N_35850);
or U36940 (N_36940,N_35800,N_35607);
or U36941 (N_36941,N_35699,N_35410);
and U36942 (N_36942,N_35551,N_35043);
nor U36943 (N_36943,N_35407,N_35460);
nand U36944 (N_36944,N_35520,N_35673);
nor U36945 (N_36945,N_35831,N_35267);
nor U36946 (N_36946,N_35916,N_35511);
nand U36947 (N_36947,N_35058,N_35036);
nor U36948 (N_36948,N_35489,N_35087);
or U36949 (N_36949,N_35467,N_35162);
nor U36950 (N_36950,N_35369,N_35884);
xnor U36951 (N_36951,N_35343,N_35751);
nor U36952 (N_36952,N_35577,N_35279);
nor U36953 (N_36953,N_35037,N_35084);
nor U36954 (N_36954,N_35550,N_35381);
and U36955 (N_36955,N_35138,N_35657);
nand U36956 (N_36956,N_35417,N_35731);
or U36957 (N_36957,N_35939,N_35502);
xnor U36958 (N_36958,N_35820,N_35289);
xor U36959 (N_36959,N_35568,N_35628);
or U36960 (N_36960,N_35293,N_35691);
xnor U36961 (N_36961,N_35998,N_35035);
nand U36962 (N_36962,N_35740,N_35911);
nand U36963 (N_36963,N_35157,N_35514);
and U36964 (N_36964,N_35456,N_35226);
nand U36965 (N_36965,N_35353,N_35213);
xnor U36966 (N_36966,N_35025,N_35678);
nand U36967 (N_36967,N_35597,N_35813);
nor U36968 (N_36968,N_35657,N_35461);
nor U36969 (N_36969,N_35290,N_35503);
xnor U36970 (N_36970,N_35839,N_35373);
or U36971 (N_36971,N_35678,N_35365);
or U36972 (N_36972,N_35855,N_35113);
and U36973 (N_36973,N_35501,N_35616);
nand U36974 (N_36974,N_35794,N_35459);
nand U36975 (N_36975,N_35239,N_35358);
nor U36976 (N_36976,N_35891,N_35388);
nor U36977 (N_36977,N_35638,N_35395);
or U36978 (N_36978,N_35666,N_35873);
nor U36979 (N_36979,N_35593,N_35552);
and U36980 (N_36980,N_35307,N_35588);
or U36981 (N_36981,N_35379,N_35768);
nor U36982 (N_36982,N_35252,N_35859);
or U36983 (N_36983,N_35768,N_35341);
nand U36984 (N_36984,N_35410,N_35261);
nor U36985 (N_36985,N_35221,N_35140);
xor U36986 (N_36986,N_35849,N_35234);
and U36987 (N_36987,N_35769,N_35594);
nor U36988 (N_36988,N_35770,N_35506);
and U36989 (N_36989,N_35213,N_35130);
nor U36990 (N_36990,N_35892,N_35349);
nand U36991 (N_36991,N_35059,N_35305);
nand U36992 (N_36992,N_35166,N_35460);
nand U36993 (N_36993,N_35754,N_35544);
xnor U36994 (N_36994,N_35243,N_35456);
and U36995 (N_36995,N_35960,N_35918);
xnor U36996 (N_36996,N_35724,N_35249);
or U36997 (N_36997,N_35762,N_35357);
or U36998 (N_36998,N_35241,N_35924);
xor U36999 (N_36999,N_35651,N_35527);
and U37000 (N_37000,N_36506,N_36328);
nor U37001 (N_37001,N_36063,N_36230);
xnor U37002 (N_37002,N_36713,N_36680);
xor U37003 (N_37003,N_36900,N_36019);
nor U37004 (N_37004,N_36465,N_36269);
or U37005 (N_37005,N_36355,N_36586);
or U37006 (N_37006,N_36105,N_36860);
and U37007 (N_37007,N_36255,N_36549);
nor U37008 (N_37008,N_36422,N_36492);
xor U37009 (N_37009,N_36419,N_36681);
or U37010 (N_37010,N_36003,N_36523);
and U37011 (N_37011,N_36353,N_36588);
and U37012 (N_37012,N_36677,N_36849);
and U37013 (N_37013,N_36737,N_36508);
and U37014 (N_37014,N_36342,N_36429);
or U37015 (N_37015,N_36194,N_36780);
and U37016 (N_37016,N_36909,N_36501);
nand U37017 (N_37017,N_36752,N_36314);
or U37018 (N_37018,N_36413,N_36156);
nor U37019 (N_37019,N_36468,N_36042);
xnor U37020 (N_37020,N_36356,N_36482);
nor U37021 (N_37021,N_36620,N_36236);
xor U37022 (N_37022,N_36724,N_36141);
nand U37023 (N_37023,N_36112,N_36293);
nand U37024 (N_37024,N_36814,N_36733);
xor U37025 (N_37025,N_36762,N_36957);
or U37026 (N_37026,N_36801,N_36480);
nand U37027 (N_37027,N_36689,N_36183);
nor U37028 (N_37028,N_36890,N_36216);
nor U37029 (N_37029,N_36440,N_36835);
and U37030 (N_37030,N_36720,N_36545);
or U37031 (N_37031,N_36463,N_36032);
nor U37032 (N_37032,N_36495,N_36007);
or U37033 (N_37033,N_36567,N_36272);
and U37034 (N_37034,N_36197,N_36034);
xnor U37035 (N_37035,N_36300,N_36172);
xor U37036 (N_37036,N_36641,N_36837);
or U37037 (N_37037,N_36329,N_36204);
or U37038 (N_37038,N_36858,N_36327);
nand U37039 (N_37039,N_36180,N_36582);
nand U37040 (N_37040,N_36691,N_36160);
nand U37041 (N_37041,N_36106,N_36539);
or U37042 (N_37042,N_36306,N_36349);
or U37043 (N_37043,N_36601,N_36126);
xnor U37044 (N_37044,N_36098,N_36187);
and U37045 (N_37045,N_36503,N_36690);
or U37046 (N_37046,N_36687,N_36653);
nor U37047 (N_37047,N_36504,N_36088);
nand U37048 (N_37048,N_36916,N_36316);
or U37049 (N_37049,N_36605,N_36064);
and U37050 (N_37050,N_36487,N_36594);
or U37051 (N_37051,N_36763,N_36373);
and U37052 (N_37052,N_36607,N_36921);
nand U37053 (N_37053,N_36371,N_36121);
and U37054 (N_37054,N_36648,N_36873);
or U37055 (N_37055,N_36374,N_36889);
nand U37056 (N_37056,N_36340,N_36627);
xor U37057 (N_37057,N_36838,N_36436);
or U37058 (N_37058,N_36602,N_36922);
nand U37059 (N_37059,N_36417,N_36973);
nor U37060 (N_37060,N_36336,N_36283);
nor U37061 (N_37061,N_36818,N_36745);
or U37062 (N_37062,N_36666,N_36410);
or U37063 (N_37063,N_36553,N_36273);
nand U37064 (N_37064,N_36358,N_36623);
nand U37065 (N_37065,N_36587,N_36531);
and U37066 (N_37066,N_36874,N_36235);
and U37067 (N_37067,N_36335,N_36109);
nand U37068 (N_37068,N_36043,N_36341);
nor U37069 (N_37069,N_36489,N_36507);
and U37070 (N_37070,N_36735,N_36521);
and U37071 (N_37071,N_36882,N_36123);
xor U37072 (N_37072,N_36220,N_36223);
nand U37073 (N_37073,N_36974,N_36920);
nor U37074 (N_37074,N_36161,N_36142);
nor U37075 (N_37075,N_36451,N_36839);
xor U37076 (N_37076,N_36700,N_36093);
xnor U37077 (N_37077,N_36731,N_36954);
nand U37078 (N_37078,N_36815,N_36317);
nor U37079 (N_37079,N_36144,N_36218);
and U37080 (N_37080,N_36879,N_36334);
nand U37081 (N_37081,N_36399,N_36247);
and U37082 (N_37082,N_36092,N_36771);
nor U37083 (N_37083,N_36303,N_36982);
and U37084 (N_37084,N_36449,N_36195);
and U37085 (N_37085,N_36090,N_36536);
xor U37086 (N_37086,N_36716,N_36151);
nand U37087 (N_37087,N_36181,N_36817);
or U37088 (N_37088,N_36357,N_36484);
xor U37089 (N_37089,N_36165,N_36604);
or U37090 (N_37090,N_36391,N_36490);
and U37091 (N_37091,N_36397,N_36229);
or U37092 (N_37092,N_36389,N_36385);
and U37093 (N_37093,N_36411,N_36406);
nor U37094 (N_37094,N_36132,N_36787);
nand U37095 (N_37095,N_36635,N_36932);
xnor U37096 (N_37096,N_36073,N_36499);
and U37097 (N_37097,N_36758,N_36937);
or U37098 (N_37098,N_36201,N_36339);
xnor U37099 (N_37099,N_36946,N_36944);
or U37100 (N_37100,N_36377,N_36853);
or U37101 (N_37101,N_36893,N_36343);
and U37102 (N_37102,N_36829,N_36514);
and U37103 (N_37103,N_36650,N_36538);
and U37104 (N_37104,N_36557,N_36697);
nand U37105 (N_37105,N_36015,N_36759);
xor U37106 (N_37106,N_36592,N_36800);
nand U37107 (N_37107,N_36078,N_36590);
xor U37108 (N_37108,N_36446,N_36452);
nand U37109 (N_37109,N_36625,N_36743);
nor U37110 (N_37110,N_36097,N_36897);
or U37111 (N_37111,N_36943,N_36439);
xnor U37112 (N_37112,N_36797,N_36869);
or U37113 (N_37113,N_36871,N_36200);
nor U37114 (N_37114,N_36703,N_36668);
or U37115 (N_37115,N_36904,N_36091);
or U37116 (N_37116,N_36579,N_36467);
nand U37117 (N_37117,N_36626,N_36387);
xnor U37118 (N_37118,N_36000,N_36732);
or U37119 (N_37119,N_36775,N_36155);
xor U37120 (N_37120,N_36407,N_36584);
nand U37121 (N_37121,N_36622,N_36131);
and U37122 (N_37122,N_36998,N_36840);
and U37123 (N_37123,N_36020,N_36145);
nand U37124 (N_37124,N_36649,N_36393);
or U37125 (N_37125,N_36354,N_36647);
xnor U37126 (N_37126,N_36027,N_36094);
or U37127 (N_37127,N_36896,N_36163);
xor U37128 (N_37128,N_36014,N_36364);
xnor U37129 (N_37129,N_36125,N_36381);
nand U37130 (N_37130,N_36312,N_36778);
or U37131 (N_37131,N_36881,N_36485);
xnor U37132 (N_37132,N_36520,N_36437);
nor U37133 (N_37133,N_36319,N_36662);
or U37134 (N_37134,N_36102,N_36258);
nand U37135 (N_37135,N_36198,N_36908);
nor U37136 (N_37136,N_36863,N_36864);
and U37137 (N_37137,N_36565,N_36834);
and U37138 (N_37138,N_36427,N_36299);
and U37139 (N_37139,N_36718,N_36008);
or U37140 (N_37140,N_36790,N_36256);
xnor U37141 (N_37141,N_36750,N_36192);
nor U37142 (N_37142,N_36722,N_36244);
nand U37143 (N_37143,N_36224,N_36631);
or U37144 (N_37144,N_36940,N_36977);
nor U37145 (N_37145,N_36848,N_36702);
and U37146 (N_37146,N_36456,N_36975);
nor U37147 (N_37147,N_36945,N_36053);
or U37148 (N_37148,N_36108,N_36652);
or U37149 (N_37149,N_36577,N_36799);
nand U37150 (N_37150,N_36210,N_36477);
nor U37151 (N_37151,N_36375,N_36729);
and U37152 (N_37152,N_36331,N_36766);
nor U37153 (N_37153,N_36599,N_36886);
xor U37154 (N_37154,N_36699,N_36136);
xnor U37155 (N_37155,N_36443,N_36395);
nand U37156 (N_37156,N_36157,N_36823);
nor U37157 (N_37157,N_36225,N_36039);
xnor U37158 (N_37158,N_36442,N_36546);
xor U37159 (N_37159,N_36698,N_36177);
nor U37160 (N_37160,N_36332,N_36469);
nand U37161 (N_37161,N_36459,N_36609);
nor U37162 (N_37162,N_36979,N_36017);
nor U37163 (N_37163,N_36241,N_36911);
and U37164 (N_37164,N_36706,N_36645);
or U37165 (N_37165,N_36403,N_36378);
and U37166 (N_37166,N_36827,N_36527);
xnor U37167 (N_37167,N_36770,N_36238);
and U37168 (N_37168,N_36639,N_36392);
nand U37169 (N_37169,N_36617,N_36031);
xnor U37170 (N_37170,N_36040,N_36203);
nor U37171 (N_37171,N_36846,N_36500);
nand U37172 (N_37172,N_36011,N_36862);
or U37173 (N_37173,N_36859,N_36765);
and U37174 (N_37174,N_36473,N_36717);
nor U37175 (N_37175,N_36033,N_36783);
nand U37176 (N_37176,N_36948,N_36453);
and U37177 (N_37177,N_36656,N_36268);
and U37178 (N_37178,N_36928,N_36644);
nor U37179 (N_37179,N_36118,N_36338);
nand U37180 (N_37180,N_36110,N_36426);
and U37181 (N_37181,N_36951,N_36548);
and U37182 (N_37182,N_36372,N_36190);
nand U37183 (N_37183,N_36902,N_36575);
or U37184 (N_37184,N_36619,N_36747);
xnor U37185 (N_37185,N_36832,N_36267);
nor U37186 (N_37186,N_36483,N_36448);
nor U37187 (N_37187,N_36174,N_36528);
nor U37188 (N_37188,N_36791,N_36785);
and U37189 (N_37189,N_36637,N_36021);
or U37190 (N_37190,N_36083,N_36547);
xor U37191 (N_37191,N_36776,N_36866);
or U37192 (N_37192,N_36305,N_36360);
nand U37193 (N_37193,N_36281,N_36980);
nor U37194 (N_37194,N_36628,N_36615);
xor U37195 (N_37195,N_36464,N_36060);
nor U37196 (N_37196,N_36262,N_36741);
and U37197 (N_37197,N_36366,N_36029);
nand U37198 (N_37198,N_36030,N_36746);
nor U37199 (N_37199,N_36825,N_36674);
nand U37200 (N_37200,N_36856,N_36655);
and U37201 (N_37201,N_36414,N_36298);
nor U37202 (N_37202,N_36111,N_36045);
xnor U37203 (N_37203,N_36169,N_36461);
or U37204 (N_37204,N_36868,N_36960);
and U37205 (N_37205,N_36259,N_36854);
nand U37206 (N_37206,N_36277,N_36576);
xor U37207 (N_37207,N_36606,N_36124);
and U37208 (N_37208,N_36404,N_36001);
nand U37209 (N_37209,N_36361,N_36963);
or U37210 (N_37210,N_36153,N_36075);
nor U37211 (N_37211,N_36919,N_36213);
or U37212 (N_37212,N_36719,N_36185);
nand U37213 (N_37213,N_36113,N_36081);
or U37214 (N_37214,N_36905,N_36917);
or U37215 (N_37215,N_36474,N_36792);
and U37216 (N_37216,N_36009,N_36322);
or U37217 (N_37217,N_36738,N_36985);
or U37218 (N_37218,N_36167,N_36250);
and U37219 (N_37219,N_36704,N_36047);
nor U37220 (N_37220,N_36184,N_36274);
xor U37221 (N_37221,N_36209,N_36370);
nand U37222 (N_37222,N_36087,N_36941);
nand U37223 (N_37223,N_36475,N_36543);
or U37224 (N_37224,N_36667,N_36233);
nand U37225 (N_37225,N_36659,N_36784);
xnor U37226 (N_37226,N_36068,N_36898);
and U37227 (N_37227,N_36583,N_36023);
nand U37228 (N_37228,N_36956,N_36050);
nor U37229 (N_37229,N_36611,N_36330);
nand U37230 (N_37230,N_36796,N_36296);
or U37231 (N_37231,N_36526,N_36822);
and U37232 (N_37232,N_36816,N_36457);
nand U37233 (N_37233,N_36510,N_36289);
nand U37234 (N_37234,N_36734,N_36012);
and U37235 (N_37235,N_36875,N_36836);
and U37236 (N_37236,N_36046,N_36679);
and U37237 (N_37237,N_36057,N_36369);
nor U37238 (N_37238,N_36367,N_36261);
xnor U37239 (N_37239,N_36382,N_36754);
xor U37240 (N_37240,N_36935,N_36479);
xor U37241 (N_37241,N_36416,N_36663);
and U37242 (N_37242,N_36753,N_36424);
xor U37243 (N_37243,N_36234,N_36795);
xor U37244 (N_37244,N_36207,N_36175);
xnor U37245 (N_37245,N_36561,N_36772);
xnor U37246 (N_37246,N_36685,N_36143);
xnor U37247 (N_37247,N_36333,N_36560);
nand U37248 (N_37248,N_36950,N_36968);
nor U37249 (N_37249,N_36805,N_36678);
nand U37250 (N_37250,N_36164,N_36037);
nor U37251 (N_37251,N_36925,N_36432);
xor U37252 (N_37252,N_36845,N_36036);
and U37253 (N_37253,N_36170,N_36794);
nand U37254 (N_37254,N_36010,N_36967);
or U37255 (N_37255,N_36253,N_36114);
xor U37256 (N_37256,N_36833,N_36984);
nand U37257 (N_37257,N_36423,N_36598);
or U37258 (N_37258,N_36239,N_36054);
nand U37259 (N_37259,N_36280,N_36673);
and U37260 (N_37260,N_36664,N_36851);
xor U37261 (N_37261,N_36128,N_36646);
xnor U37262 (N_37262,N_36675,N_36297);
nand U37263 (N_37263,N_36292,N_36824);
xnor U37264 (N_37264,N_36512,N_36351);
xor U37265 (N_37265,N_36965,N_36894);
xor U37266 (N_37266,N_36511,N_36251);
or U37267 (N_37267,N_36494,N_36751);
nand U37268 (N_37268,N_36600,N_36970);
nor U37269 (N_37269,N_36242,N_36100);
and U37270 (N_37270,N_36728,N_36642);
or U37271 (N_37271,N_36544,N_36325);
xnor U37272 (N_37272,N_36006,N_36318);
and U37273 (N_37273,N_36994,N_36686);
nor U37274 (N_37274,N_36182,N_36658);
or U37275 (N_37275,N_36742,N_36725);
and U37276 (N_37276,N_36643,N_36913);
nor U37277 (N_37277,N_36566,N_36401);
nand U37278 (N_37278,N_36660,N_36711);
nor U37279 (N_37279,N_36966,N_36537);
or U37280 (N_37280,N_36018,N_36513);
or U37281 (N_37281,N_36555,N_36271);
or U37282 (N_37282,N_36556,N_36542);
xnor U37283 (N_37283,N_36215,N_36807);
and U37284 (N_37284,N_36603,N_36362);
nand U37285 (N_37285,N_36841,N_36107);
nor U37286 (N_37286,N_36257,N_36774);
and U37287 (N_37287,N_36964,N_36518);
nand U37288 (N_37288,N_36263,N_36654);
nand U37289 (N_37289,N_36723,N_36997);
nor U37290 (N_37290,N_36051,N_36912);
nand U37291 (N_37291,N_36564,N_36782);
xor U37292 (N_37292,N_36049,N_36178);
or U37293 (N_37293,N_36552,N_36608);
nor U37294 (N_37294,N_36350,N_36044);
nand U37295 (N_37295,N_36409,N_36249);
or U37296 (N_37296,N_36188,N_36137);
xnor U37297 (N_37297,N_36291,N_36502);
nor U37298 (N_37298,N_36466,N_36883);
and U37299 (N_37299,N_36323,N_36714);
xor U37300 (N_37300,N_36072,N_36802);
and U37301 (N_37301,N_36844,N_36497);
xor U37302 (N_37302,N_36693,N_36450);
xnor U37303 (N_37303,N_36779,N_36384);
and U37304 (N_37304,N_36761,N_36089);
nand U37305 (N_37305,N_36877,N_36880);
and U37306 (N_37306,N_36798,N_36657);
xor U37307 (N_37307,N_36307,N_36004);
nor U37308 (N_37308,N_36744,N_36284);
nand U37309 (N_37309,N_36445,N_36591);
xnor U37310 (N_37310,N_36976,N_36290);
nand U37311 (N_37311,N_36084,N_36129);
nor U37312 (N_37312,N_36872,N_36481);
or U37313 (N_37313,N_36988,N_36831);
xnor U37314 (N_37314,N_36022,N_36804);
nor U37315 (N_37315,N_36788,N_36260);
nand U37316 (N_37316,N_36166,N_36208);
nor U37317 (N_37317,N_36246,N_36359);
nand U37318 (N_37318,N_36270,N_36438);
xnor U37319 (N_37319,N_36135,N_36670);
xor U37320 (N_37320,N_36870,N_36005);
and U37321 (N_37321,N_36884,N_36346);
or U37322 (N_37322,N_36070,N_36630);
nand U37323 (N_37323,N_36024,N_36530);
nor U37324 (N_37324,N_36493,N_36227);
xnor U37325 (N_37325,N_36803,N_36096);
nand U37326 (N_37326,N_36861,N_36154);
or U37327 (N_37327,N_36025,N_36578);
nand U37328 (N_37328,N_36295,N_36572);
nor U37329 (N_37329,N_36936,N_36843);
nand U37330 (N_37330,N_36488,N_36085);
xor U37331 (N_37331,N_36447,N_36808);
nor U37332 (N_37332,N_36961,N_36211);
and U37333 (N_37333,N_36134,N_36739);
nand U37334 (N_37334,N_36610,N_36757);
or U37335 (N_37335,N_36930,N_36554);
nor U37336 (N_37336,N_36162,N_36551);
and U37337 (N_37337,N_36122,N_36388);
xnor U37338 (N_37338,N_36632,N_36597);
nor U37339 (N_37339,N_36688,N_36119);
xor U37340 (N_37340,N_36275,N_36705);
nand U37341 (N_37341,N_36486,N_36265);
nand U37342 (N_37342,N_36321,N_36926);
and U37343 (N_37343,N_36264,N_36962);
nand U37344 (N_37344,N_36458,N_36755);
nor U37345 (N_37345,N_36101,N_36715);
nand U37346 (N_37346,N_36671,N_36232);
xor U37347 (N_37347,N_36568,N_36563);
nor U37348 (N_37348,N_36052,N_36529);
nand U37349 (N_37349,N_36115,N_36756);
and U37350 (N_37350,N_36629,N_36901);
nand U37351 (N_37351,N_36444,N_36949);
and U37352 (N_37352,N_36402,N_36308);
or U37353 (N_37353,N_36953,N_36692);
nand U37354 (N_37354,N_36186,N_36454);
nand U37355 (N_37355,N_36171,N_36809);
xnor U37356 (N_37356,N_36254,N_36365);
nor U37357 (N_37357,N_36159,N_36294);
or U37358 (N_37358,N_36672,N_36947);
nor U37359 (N_37359,N_36286,N_36243);
and U37360 (N_37360,N_36386,N_36683);
nand U37361 (N_37361,N_36337,N_36471);
nand U37362 (N_37362,N_36168,N_36891);
xnor U37363 (N_37363,N_36055,N_36730);
or U37364 (N_37364,N_36472,N_36571);
xnor U37365 (N_37365,N_36769,N_36206);
nand U37366 (N_37366,N_36852,N_36285);
nand U37367 (N_37367,N_36541,N_36158);
or U37368 (N_37368,N_36867,N_36969);
nand U37369 (N_37369,N_36086,N_36707);
or U37370 (N_37370,N_36140,N_36924);
and U37371 (N_37371,N_36038,N_36301);
nor U37372 (N_37372,N_36189,N_36990);
nand U37373 (N_37373,N_36971,N_36661);
or U37374 (N_37374,N_36228,N_36069);
or U37375 (N_37375,N_36491,N_36196);
xnor U37376 (N_37376,N_36179,N_36138);
and U37377 (N_37377,N_36534,N_36139);
or U37378 (N_37378,N_36431,N_36237);
xor U37379 (N_37379,N_36418,N_36080);
or U37380 (N_37380,N_36302,N_36585);
and U37381 (N_37381,N_36996,N_36048);
nor U37382 (N_37382,N_36694,N_36726);
or U37383 (N_37383,N_36279,N_36133);
xnor U37384 (N_37384,N_36222,N_36972);
or U37385 (N_37385,N_36748,N_36721);
or U37386 (N_37386,N_36569,N_36749);
or U37387 (N_37387,N_36918,N_36016);
and U37388 (N_37388,N_36176,N_36435);
and U37389 (N_37389,N_36781,N_36540);
nand U37390 (N_37390,N_36434,N_36887);
nand U37391 (N_37391,N_36640,N_36065);
xor U37392 (N_37392,N_36193,N_36533);
and U37393 (N_37393,N_36116,N_36276);
or U37394 (N_37394,N_36199,N_36383);
and U37395 (N_37395,N_36519,N_36978);
nor U37396 (N_37396,N_36152,N_36959);
xor U37397 (N_37397,N_36056,N_36221);
nor U37398 (N_37398,N_36938,N_36248);
nor U37399 (N_37399,N_36558,N_36226);
nor U37400 (N_37400,N_36266,N_36855);
and U37401 (N_37401,N_36573,N_36310);
or U37402 (N_37402,N_36813,N_36217);
or U37403 (N_37403,N_36214,N_36826);
xnor U37404 (N_37404,N_36740,N_36376);
or U37405 (N_37405,N_36099,N_36104);
or U37406 (N_37406,N_36428,N_36789);
xnor U37407 (N_37407,N_36934,N_36987);
nor U37408 (N_37408,N_36983,N_36103);
or U37409 (N_37409,N_36621,N_36288);
and U37410 (N_37410,N_36379,N_36709);
and U37411 (N_37411,N_36326,N_36895);
nand U37412 (N_37412,N_36614,N_36460);
nor U37413 (N_37413,N_36390,N_36910);
nor U37414 (N_37414,N_36701,N_36793);
xnor U37415 (N_37415,N_36287,N_36550);
nand U37416 (N_37416,N_36535,N_36130);
and U37417 (N_37417,N_36516,N_36712);
or U37418 (N_37418,N_36958,N_36219);
nand U37419 (N_37419,N_36923,N_36074);
nor U37420 (N_37420,N_36992,N_36117);
and U37421 (N_37421,N_36684,N_36915);
nor U37422 (N_37422,N_36311,N_36927);
nand U37423 (N_37423,N_36574,N_36931);
xor U37424 (N_37424,N_36764,N_36150);
and U37425 (N_37425,N_36899,N_36421);
nand U37426 (N_37426,N_36914,N_36624);
or U37427 (N_37427,N_36127,N_36478);
nor U37428 (N_37428,N_36842,N_36616);
and U37429 (N_37429,N_36430,N_36995);
nor U37430 (N_37430,N_36231,N_36524);
nand U37431 (N_37431,N_36363,N_36476);
or U37432 (N_37432,N_36589,N_36821);
nand U37433 (N_37433,N_36313,N_36618);
and U37434 (N_37434,N_36952,N_36522);
nor U37435 (N_37435,N_36061,N_36408);
nor U37436 (N_37436,N_36425,N_36026);
xor U37437 (N_37437,N_36441,N_36282);
xor U37438 (N_37438,N_36191,N_36892);
and U37439 (N_37439,N_36819,N_36278);
nor U37440 (N_37440,N_36532,N_36682);
or U37441 (N_37441,N_36595,N_36768);
or U37442 (N_37442,N_36398,N_36252);
and U37443 (N_37443,N_36939,N_36412);
or U37444 (N_37444,N_36695,N_36580);
nand U37445 (N_37445,N_36828,N_36309);
xor U37446 (N_37446,N_36035,N_36651);
and U37447 (N_37447,N_36955,N_36202);
xor U37448 (N_37448,N_36767,N_36559);
nand U37449 (N_37449,N_36149,N_36173);
nand U37450 (N_37450,N_36760,N_36380);
and U37451 (N_37451,N_36810,N_36633);
and U37452 (N_37452,N_36865,N_36405);
xnor U37453 (N_37453,N_36002,N_36878);
xnor U37454 (N_37454,N_36636,N_36400);
nand U37455 (N_37455,N_36525,N_36498);
xnor U37456 (N_37456,N_36517,N_36028);
and U37457 (N_37457,N_36324,N_36240);
and U37458 (N_37458,N_36071,N_36989);
or U37459 (N_37459,N_36062,N_36876);
nand U37460 (N_37460,N_36907,N_36368);
or U37461 (N_37461,N_36058,N_36515);
and U37462 (N_37462,N_36736,N_36066);
or U37463 (N_37463,N_36986,N_36212);
nand U37464 (N_37464,N_36509,N_36396);
nor U37465 (N_37465,N_36777,N_36727);
or U37466 (N_37466,N_36634,N_36245);
or U37467 (N_37467,N_36773,N_36929);
nor U37468 (N_37468,N_36613,N_36415);
and U37469 (N_37469,N_36347,N_36847);
and U37470 (N_37470,N_36981,N_36067);
nand U37471 (N_37471,N_36999,N_36570);
nor U37472 (N_37472,N_36095,N_36903);
nor U37473 (N_37473,N_36612,N_36665);
xnor U37474 (N_37474,N_36857,N_36786);
and U37475 (N_37475,N_36315,N_36205);
xnor U37476 (N_37476,N_36676,N_36348);
nand U37477 (N_37477,N_36076,N_36470);
nand U37478 (N_37478,N_36811,N_36079);
and U37479 (N_37479,N_36077,N_36708);
xor U37480 (N_37480,N_36320,N_36496);
nand U37481 (N_37481,N_36933,N_36850);
or U37482 (N_37482,N_36885,N_36013);
nand U37483 (N_37483,N_36888,N_36120);
and U37484 (N_37484,N_36820,N_36345);
nor U37485 (N_37485,N_36596,N_36993);
xnor U37486 (N_37486,N_36082,N_36420);
nor U37487 (N_37487,N_36059,N_36806);
xnor U37488 (N_37488,N_36669,N_36812);
nand U37489 (N_37489,N_36505,N_36455);
nor U37490 (N_37490,N_36433,N_36942);
or U37491 (N_37491,N_36041,N_36352);
and U37492 (N_37492,N_36462,N_36991);
nor U37493 (N_37493,N_36638,N_36906);
xor U37494 (N_37494,N_36146,N_36344);
xor U37495 (N_37495,N_36710,N_36696);
and U37496 (N_37496,N_36593,N_36830);
xnor U37497 (N_37497,N_36304,N_36147);
xnor U37498 (N_37498,N_36394,N_36581);
nand U37499 (N_37499,N_36562,N_36148);
and U37500 (N_37500,N_36291,N_36897);
xor U37501 (N_37501,N_36216,N_36449);
nor U37502 (N_37502,N_36268,N_36505);
nand U37503 (N_37503,N_36166,N_36954);
and U37504 (N_37504,N_36119,N_36596);
nor U37505 (N_37505,N_36879,N_36923);
nor U37506 (N_37506,N_36837,N_36267);
nor U37507 (N_37507,N_36376,N_36539);
nor U37508 (N_37508,N_36068,N_36589);
xor U37509 (N_37509,N_36125,N_36447);
nand U37510 (N_37510,N_36384,N_36634);
and U37511 (N_37511,N_36764,N_36658);
xor U37512 (N_37512,N_36066,N_36637);
nand U37513 (N_37513,N_36988,N_36130);
xnor U37514 (N_37514,N_36592,N_36370);
xnor U37515 (N_37515,N_36847,N_36064);
nor U37516 (N_37516,N_36951,N_36364);
and U37517 (N_37517,N_36454,N_36366);
nand U37518 (N_37518,N_36337,N_36685);
and U37519 (N_37519,N_36755,N_36684);
nor U37520 (N_37520,N_36426,N_36276);
and U37521 (N_37521,N_36607,N_36711);
or U37522 (N_37522,N_36613,N_36727);
xor U37523 (N_37523,N_36710,N_36064);
nand U37524 (N_37524,N_36052,N_36584);
nor U37525 (N_37525,N_36159,N_36028);
xnor U37526 (N_37526,N_36057,N_36357);
xor U37527 (N_37527,N_36592,N_36162);
nand U37528 (N_37528,N_36582,N_36698);
and U37529 (N_37529,N_36297,N_36122);
and U37530 (N_37530,N_36947,N_36793);
nor U37531 (N_37531,N_36287,N_36521);
xnor U37532 (N_37532,N_36626,N_36597);
nand U37533 (N_37533,N_36069,N_36445);
xor U37534 (N_37534,N_36460,N_36061);
nand U37535 (N_37535,N_36650,N_36342);
or U37536 (N_37536,N_36965,N_36384);
or U37537 (N_37537,N_36834,N_36724);
or U37538 (N_37538,N_36515,N_36506);
or U37539 (N_37539,N_36068,N_36051);
or U37540 (N_37540,N_36616,N_36321);
or U37541 (N_37541,N_36723,N_36448);
or U37542 (N_37542,N_36589,N_36209);
nand U37543 (N_37543,N_36621,N_36553);
nor U37544 (N_37544,N_36730,N_36257);
nand U37545 (N_37545,N_36826,N_36240);
nand U37546 (N_37546,N_36460,N_36432);
nor U37547 (N_37547,N_36883,N_36058);
nor U37548 (N_37548,N_36634,N_36462);
or U37549 (N_37549,N_36941,N_36624);
nand U37550 (N_37550,N_36548,N_36164);
or U37551 (N_37551,N_36839,N_36460);
nand U37552 (N_37552,N_36552,N_36009);
nand U37553 (N_37553,N_36170,N_36993);
nand U37554 (N_37554,N_36059,N_36496);
nand U37555 (N_37555,N_36967,N_36064);
xor U37556 (N_37556,N_36940,N_36467);
or U37557 (N_37557,N_36744,N_36663);
nor U37558 (N_37558,N_36508,N_36185);
nor U37559 (N_37559,N_36567,N_36154);
and U37560 (N_37560,N_36461,N_36808);
nor U37561 (N_37561,N_36859,N_36800);
nor U37562 (N_37562,N_36915,N_36887);
and U37563 (N_37563,N_36329,N_36830);
nand U37564 (N_37564,N_36915,N_36460);
and U37565 (N_37565,N_36073,N_36861);
nand U37566 (N_37566,N_36717,N_36992);
nor U37567 (N_37567,N_36473,N_36519);
or U37568 (N_37568,N_36676,N_36295);
nand U37569 (N_37569,N_36298,N_36986);
nor U37570 (N_37570,N_36494,N_36104);
and U37571 (N_37571,N_36002,N_36123);
xnor U37572 (N_37572,N_36454,N_36386);
and U37573 (N_37573,N_36325,N_36538);
and U37574 (N_37574,N_36222,N_36338);
nand U37575 (N_37575,N_36443,N_36048);
nor U37576 (N_37576,N_36553,N_36905);
xor U37577 (N_37577,N_36878,N_36523);
xor U37578 (N_37578,N_36540,N_36901);
nor U37579 (N_37579,N_36639,N_36398);
nand U37580 (N_37580,N_36441,N_36838);
or U37581 (N_37581,N_36377,N_36134);
nand U37582 (N_37582,N_36058,N_36907);
nor U37583 (N_37583,N_36465,N_36524);
or U37584 (N_37584,N_36105,N_36592);
nor U37585 (N_37585,N_36895,N_36765);
or U37586 (N_37586,N_36681,N_36986);
and U37587 (N_37587,N_36982,N_36297);
nor U37588 (N_37588,N_36395,N_36983);
nand U37589 (N_37589,N_36393,N_36147);
nor U37590 (N_37590,N_36222,N_36830);
nand U37591 (N_37591,N_36071,N_36966);
nand U37592 (N_37592,N_36803,N_36679);
nor U37593 (N_37593,N_36972,N_36285);
and U37594 (N_37594,N_36257,N_36159);
xor U37595 (N_37595,N_36329,N_36089);
and U37596 (N_37596,N_36292,N_36651);
and U37597 (N_37597,N_36937,N_36493);
nor U37598 (N_37598,N_36419,N_36711);
nand U37599 (N_37599,N_36721,N_36422);
nor U37600 (N_37600,N_36940,N_36950);
and U37601 (N_37601,N_36705,N_36226);
nand U37602 (N_37602,N_36312,N_36761);
xnor U37603 (N_37603,N_36354,N_36565);
xnor U37604 (N_37604,N_36225,N_36275);
nand U37605 (N_37605,N_36533,N_36155);
nand U37606 (N_37606,N_36659,N_36524);
and U37607 (N_37607,N_36995,N_36160);
and U37608 (N_37608,N_36050,N_36811);
nor U37609 (N_37609,N_36305,N_36066);
nor U37610 (N_37610,N_36994,N_36611);
and U37611 (N_37611,N_36664,N_36704);
xor U37612 (N_37612,N_36562,N_36360);
xor U37613 (N_37613,N_36684,N_36349);
nor U37614 (N_37614,N_36559,N_36642);
and U37615 (N_37615,N_36617,N_36604);
nor U37616 (N_37616,N_36749,N_36571);
and U37617 (N_37617,N_36366,N_36231);
and U37618 (N_37618,N_36528,N_36340);
xnor U37619 (N_37619,N_36175,N_36541);
nor U37620 (N_37620,N_36001,N_36541);
xor U37621 (N_37621,N_36457,N_36527);
or U37622 (N_37622,N_36144,N_36308);
nand U37623 (N_37623,N_36153,N_36461);
nor U37624 (N_37624,N_36220,N_36379);
nand U37625 (N_37625,N_36394,N_36883);
and U37626 (N_37626,N_36765,N_36767);
xor U37627 (N_37627,N_36548,N_36401);
and U37628 (N_37628,N_36938,N_36043);
xor U37629 (N_37629,N_36458,N_36524);
nor U37630 (N_37630,N_36446,N_36553);
and U37631 (N_37631,N_36523,N_36694);
nand U37632 (N_37632,N_36201,N_36390);
xnor U37633 (N_37633,N_36739,N_36285);
xnor U37634 (N_37634,N_36201,N_36442);
xnor U37635 (N_37635,N_36188,N_36826);
and U37636 (N_37636,N_36580,N_36854);
nor U37637 (N_37637,N_36289,N_36232);
nor U37638 (N_37638,N_36513,N_36991);
and U37639 (N_37639,N_36899,N_36378);
or U37640 (N_37640,N_36705,N_36626);
nand U37641 (N_37641,N_36448,N_36243);
and U37642 (N_37642,N_36691,N_36085);
nor U37643 (N_37643,N_36453,N_36028);
and U37644 (N_37644,N_36171,N_36467);
nor U37645 (N_37645,N_36134,N_36178);
nor U37646 (N_37646,N_36987,N_36899);
and U37647 (N_37647,N_36132,N_36025);
nor U37648 (N_37648,N_36204,N_36818);
nor U37649 (N_37649,N_36402,N_36647);
nand U37650 (N_37650,N_36552,N_36353);
nand U37651 (N_37651,N_36960,N_36155);
xor U37652 (N_37652,N_36146,N_36663);
and U37653 (N_37653,N_36680,N_36280);
or U37654 (N_37654,N_36574,N_36845);
nor U37655 (N_37655,N_36324,N_36060);
nor U37656 (N_37656,N_36638,N_36988);
nand U37657 (N_37657,N_36619,N_36334);
nor U37658 (N_37658,N_36095,N_36487);
and U37659 (N_37659,N_36969,N_36786);
xor U37660 (N_37660,N_36805,N_36724);
nor U37661 (N_37661,N_36437,N_36583);
nand U37662 (N_37662,N_36579,N_36028);
nor U37663 (N_37663,N_36458,N_36295);
nor U37664 (N_37664,N_36499,N_36254);
and U37665 (N_37665,N_36485,N_36770);
and U37666 (N_37666,N_36806,N_36084);
nor U37667 (N_37667,N_36554,N_36078);
and U37668 (N_37668,N_36181,N_36680);
and U37669 (N_37669,N_36590,N_36250);
nand U37670 (N_37670,N_36474,N_36093);
or U37671 (N_37671,N_36499,N_36385);
or U37672 (N_37672,N_36287,N_36638);
nand U37673 (N_37673,N_36791,N_36407);
xor U37674 (N_37674,N_36988,N_36688);
nor U37675 (N_37675,N_36156,N_36056);
nor U37676 (N_37676,N_36998,N_36047);
nor U37677 (N_37677,N_36771,N_36677);
and U37678 (N_37678,N_36770,N_36021);
or U37679 (N_37679,N_36128,N_36838);
and U37680 (N_37680,N_36377,N_36118);
nor U37681 (N_37681,N_36784,N_36930);
nor U37682 (N_37682,N_36285,N_36110);
nor U37683 (N_37683,N_36470,N_36793);
nand U37684 (N_37684,N_36477,N_36646);
nand U37685 (N_37685,N_36432,N_36874);
and U37686 (N_37686,N_36809,N_36309);
nor U37687 (N_37687,N_36725,N_36935);
xnor U37688 (N_37688,N_36947,N_36749);
xnor U37689 (N_37689,N_36892,N_36160);
and U37690 (N_37690,N_36611,N_36112);
and U37691 (N_37691,N_36951,N_36438);
nor U37692 (N_37692,N_36196,N_36981);
nor U37693 (N_37693,N_36724,N_36979);
or U37694 (N_37694,N_36959,N_36178);
and U37695 (N_37695,N_36739,N_36735);
or U37696 (N_37696,N_36279,N_36176);
nand U37697 (N_37697,N_36260,N_36551);
nor U37698 (N_37698,N_36367,N_36593);
nor U37699 (N_37699,N_36153,N_36997);
nand U37700 (N_37700,N_36595,N_36872);
or U37701 (N_37701,N_36366,N_36737);
and U37702 (N_37702,N_36092,N_36582);
xnor U37703 (N_37703,N_36159,N_36229);
or U37704 (N_37704,N_36205,N_36947);
and U37705 (N_37705,N_36148,N_36926);
nor U37706 (N_37706,N_36983,N_36109);
xnor U37707 (N_37707,N_36370,N_36833);
nor U37708 (N_37708,N_36625,N_36513);
or U37709 (N_37709,N_36264,N_36973);
nor U37710 (N_37710,N_36021,N_36588);
and U37711 (N_37711,N_36347,N_36959);
nor U37712 (N_37712,N_36931,N_36381);
nand U37713 (N_37713,N_36493,N_36047);
xnor U37714 (N_37714,N_36281,N_36548);
xor U37715 (N_37715,N_36304,N_36360);
nor U37716 (N_37716,N_36643,N_36634);
and U37717 (N_37717,N_36158,N_36542);
nand U37718 (N_37718,N_36439,N_36207);
and U37719 (N_37719,N_36183,N_36881);
or U37720 (N_37720,N_36990,N_36083);
nor U37721 (N_37721,N_36867,N_36136);
xnor U37722 (N_37722,N_36744,N_36415);
xor U37723 (N_37723,N_36984,N_36757);
or U37724 (N_37724,N_36010,N_36305);
xnor U37725 (N_37725,N_36956,N_36204);
nand U37726 (N_37726,N_36817,N_36312);
or U37727 (N_37727,N_36707,N_36971);
or U37728 (N_37728,N_36976,N_36309);
nand U37729 (N_37729,N_36401,N_36482);
xnor U37730 (N_37730,N_36229,N_36240);
or U37731 (N_37731,N_36580,N_36331);
nor U37732 (N_37732,N_36486,N_36092);
nand U37733 (N_37733,N_36778,N_36119);
and U37734 (N_37734,N_36959,N_36410);
nor U37735 (N_37735,N_36175,N_36181);
and U37736 (N_37736,N_36879,N_36221);
xnor U37737 (N_37737,N_36619,N_36965);
xor U37738 (N_37738,N_36628,N_36904);
nor U37739 (N_37739,N_36566,N_36690);
nor U37740 (N_37740,N_36292,N_36773);
or U37741 (N_37741,N_36215,N_36404);
xor U37742 (N_37742,N_36651,N_36271);
and U37743 (N_37743,N_36307,N_36298);
nor U37744 (N_37744,N_36379,N_36982);
nand U37745 (N_37745,N_36437,N_36060);
xnor U37746 (N_37746,N_36735,N_36606);
or U37747 (N_37747,N_36182,N_36903);
and U37748 (N_37748,N_36689,N_36271);
xor U37749 (N_37749,N_36728,N_36265);
nor U37750 (N_37750,N_36435,N_36288);
xnor U37751 (N_37751,N_36627,N_36435);
or U37752 (N_37752,N_36382,N_36799);
and U37753 (N_37753,N_36757,N_36527);
xor U37754 (N_37754,N_36542,N_36257);
or U37755 (N_37755,N_36038,N_36833);
nand U37756 (N_37756,N_36990,N_36606);
nor U37757 (N_37757,N_36796,N_36544);
and U37758 (N_37758,N_36977,N_36497);
nand U37759 (N_37759,N_36919,N_36614);
or U37760 (N_37760,N_36816,N_36139);
xor U37761 (N_37761,N_36044,N_36465);
nor U37762 (N_37762,N_36506,N_36425);
or U37763 (N_37763,N_36603,N_36705);
and U37764 (N_37764,N_36401,N_36633);
or U37765 (N_37765,N_36456,N_36378);
or U37766 (N_37766,N_36764,N_36295);
nand U37767 (N_37767,N_36877,N_36149);
nor U37768 (N_37768,N_36266,N_36967);
xor U37769 (N_37769,N_36130,N_36626);
and U37770 (N_37770,N_36901,N_36222);
nor U37771 (N_37771,N_36680,N_36953);
xnor U37772 (N_37772,N_36334,N_36517);
nand U37773 (N_37773,N_36360,N_36872);
and U37774 (N_37774,N_36416,N_36320);
and U37775 (N_37775,N_36564,N_36360);
or U37776 (N_37776,N_36724,N_36484);
nor U37777 (N_37777,N_36893,N_36396);
and U37778 (N_37778,N_36910,N_36903);
xnor U37779 (N_37779,N_36391,N_36913);
nor U37780 (N_37780,N_36609,N_36366);
and U37781 (N_37781,N_36486,N_36294);
nor U37782 (N_37782,N_36649,N_36996);
or U37783 (N_37783,N_36468,N_36075);
nand U37784 (N_37784,N_36554,N_36766);
or U37785 (N_37785,N_36453,N_36742);
nand U37786 (N_37786,N_36293,N_36040);
xnor U37787 (N_37787,N_36021,N_36073);
xor U37788 (N_37788,N_36718,N_36845);
and U37789 (N_37789,N_36372,N_36269);
or U37790 (N_37790,N_36743,N_36977);
or U37791 (N_37791,N_36291,N_36747);
nand U37792 (N_37792,N_36486,N_36145);
or U37793 (N_37793,N_36045,N_36152);
and U37794 (N_37794,N_36058,N_36921);
nand U37795 (N_37795,N_36858,N_36762);
xor U37796 (N_37796,N_36458,N_36669);
nand U37797 (N_37797,N_36996,N_36340);
and U37798 (N_37798,N_36146,N_36072);
or U37799 (N_37799,N_36403,N_36489);
nor U37800 (N_37800,N_36696,N_36077);
or U37801 (N_37801,N_36513,N_36995);
nand U37802 (N_37802,N_36298,N_36698);
or U37803 (N_37803,N_36010,N_36925);
and U37804 (N_37804,N_36061,N_36202);
xor U37805 (N_37805,N_36069,N_36154);
xnor U37806 (N_37806,N_36321,N_36082);
nand U37807 (N_37807,N_36237,N_36501);
xor U37808 (N_37808,N_36084,N_36538);
and U37809 (N_37809,N_36871,N_36114);
xor U37810 (N_37810,N_36993,N_36982);
xnor U37811 (N_37811,N_36832,N_36242);
nand U37812 (N_37812,N_36035,N_36093);
nor U37813 (N_37813,N_36973,N_36843);
xor U37814 (N_37814,N_36092,N_36633);
xor U37815 (N_37815,N_36402,N_36924);
nand U37816 (N_37816,N_36544,N_36837);
nor U37817 (N_37817,N_36498,N_36482);
and U37818 (N_37818,N_36649,N_36804);
and U37819 (N_37819,N_36443,N_36030);
xor U37820 (N_37820,N_36004,N_36592);
xor U37821 (N_37821,N_36476,N_36573);
nor U37822 (N_37822,N_36513,N_36043);
nor U37823 (N_37823,N_36077,N_36135);
and U37824 (N_37824,N_36049,N_36034);
xnor U37825 (N_37825,N_36023,N_36536);
nand U37826 (N_37826,N_36824,N_36571);
or U37827 (N_37827,N_36456,N_36159);
xor U37828 (N_37828,N_36247,N_36274);
xnor U37829 (N_37829,N_36517,N_36627);
nor U37830 (N_37830,N_36001,N_36985);
xor U37831 (N_37831,N_36162,N_36560);
nand U37832 (N_37832,N_36012,N_36447);
or U37833 (N_37833,N_36339,N_36745);
nor U37834 (N_37834,N_36015,N_36472);
or U37835 (N_37835,N_36721,N_36023);
and U37836 (N_37836,N_36618,N_36816);
and U37837 (N_37837,N_36453,N_36444);
and U37838 (N_37838,N_36637,N_36540);
xor U37839 (N_37839,N_36876,N_36768);
xnor U37840 (N_37840,N_36919,N_36338);
xnor U37841 (N_37841,N_36733,N_36405);
and U37842 (N_37842,N_36400,N_36311);
and U37843 (N_37843,N_36493,N_36746);
nor U37844 (N_37844,N_36476,N_36896);
and U37845 (N_37845,N_36193,N_36599);
and U37846 (N_37846,N_36831,N_36248);
nor U37847 (N_37847,N_36331,N_36177);
nor U37848 (N_37848,N_36966,N_36700);
xor U37849 (N_37849,N_36310,N_36894);
xnor U37850 (N_37850,N_36032,N_36779);
or U37851 (N_37851,N_36576,N_36686);
or U37852 (N_37852,N_36094,N_36543);
nand U37853 (N_37853,N_36844,N_36310);
nor U37854 (N_37854,N_36531,N_36476);
or U37855 (N_37855,N_36041,N_36582);
and U37856 (N_37856,N_36186,N_36390);
nor U37857 (N_37857,N_36889,N_36601);
or U37858 (N_37858,N_36306,N_36678);
xor U37859 (N_37859,N_36155,N_36484);
or U37860 (N_37860,N_36189,N_36456);
nor U37861 (N_37861,N_36989,N_36423);
or U37862 (N_37862,N_36565,N_36038);
nand U37863 (N_37863,N_36970,N_36344);
nand U37864 (N_37864,N_36516,N_36382);
nor U37865 (N_37865,N_36316,N_36877);
and U37866 (N_37866,N_36286,N_36467);
and U37867 (N_37867,N_36436,N_36996);
nor U37868 (N_37868,N_36326,N_36231);
xnor U37869 (N_37869,N_36962,N_36793);
nor U37870 (N_37870,N_36972,N_36434);
and U37871 (N_37871,N_36676,N_36941);
xor U37872 (N_37872,N_36611,N_36059);
nor U37873 (N_37873,N_36147,N_36773);
xor U37874 (N_37874,N_36118,N_36437);
or U37875 (N_37875,N_36584,N_36336);
nand U37876 (N_37876,N_36903,N_36501);
nand U37877 (N_37877,N_36762,N_36281);
xor U37878 (N_37878,N_36416,N_36392);
or U37879 (N_37879,N_36059,N_36671);
and U37880 (N_37880,N_36201,N_36039);
and U37881 (N_37881,N_36252,N_36074);
nor U37882 (N_37882,N_36305,N_36730);
nand U37883 (N_37883,N_36394,N_36303);
nor U37884 (N_37884,N_36259,N_36139);
nand U37885 (N_37885,N_36567,N_36348);
or U37886 (N_37886,N_36183,N_36405);
xnor U37887 (N_37887,N_36873,N_36343);
nand U37888 (N_37888,N_36531,N_36511);
nor U37889 (N_37889,N_36239,N_36751);
xor U37890 (N_37890,N_36239,N_36116);
nor U37891 (N_37891,N_36268,N_36716);
or U37892 (N_37892,N_36944,N_36698);
or U37893 (N_37893,N_36608,N_36271);
and U37894 (N_37894,N_36255,N_36233);
and U37895 (N_37895,N_36519,N_36878);
and U37896 (N_37896,N_36826,N_36709);
nand U37897 (N_37897,N_36975,N_36657);
or U37898 (N_37898,N_36819,N_36981);
xnor U37899 (N_37899,N_36504,N_36187);
or U37900 (N_37900,N_36238,N_36955);
nor U37901 (N_37901,N_36910,N_36384);
nand U37902 (N_37902,N_36844,N_36167);
or U37903 (N_37903,N_36786,N_36987);
nor U37904 (N_37904,N_36394,N_36024);
or U37905 (N_37905,N_36834,N_36137);
nand U37906 (N_37906,N_36580,N_36357);
nor U37907 (N_37907,N_36599,N_36596);
and U37908 (N_37908,N_36101,N_36254);
nand U37909 (N_37909,N_36211,N_36224);
xnor U37910 (N_37910,N_36884,N_36419);
nor U37911 (N_37911,N_36461,N_36448);
nor U37912 (N_37912,N_36637,N_36732);
nand U37913 (N_37913,N_36348,N_36975);
or U37914 (N_37914,N_36669,N_36844);
or U37915 (N_37915,N_36475,N_36881);
xnor U37916 (N_37916,N_36192,N_36941);
xor U37917 (N_37917,N_36956,N_36103);
xor U37918 (N_37918,N_36799,N_36757);
or U37919 (N_37919,N_36410,N_36303);
or U37920 (N_37920,N_36761,N_36904);
and U37921 (N_37921,N_36088,N_36643);
xor U37922 (N_37922,N_36020,N_36692);
nor U37923 (N_37923,N_36747,N_36180);
nand U37924 (N_37924,N_36731,N_36533);
xor U37925 (N_37925,N_36279,N_36766);
and U37926 (N_37926,N_36946,N_36134);
nand U37927 (N_37927,N_36306,N_36162);
and U37928 (N_37928,N_36601,N_36028);
and U37929 (N_37929,N_36264,N_36041);
nor U37930 (N_37930,N_36502,N_36973);
nor U37931 (N_37931,N_36138,N_36337);
and U37932 (N_37932,N_36612,N_36636);
and U37933 (N_37933,N_36214,N_36761);
xnor U37934 (N_37934,N_36638,N_36811);
nand U37935 (N_37935,N_36820,N_36688);
nor U37936 (N_37936,N_36590,N_36884);
nand U37937 (N_37937,N_36442,N_36943);
or U37938 (N_37938,N_36779,N_36358);
nor U37939 (N_37939,N_36141,N_36855);
nor U37940 (N_37940,N_36792,N_36315);
nor U37941 (N_37941,N_36067,N_36076);
and U37942 (N_37942,N_36499,N_36112);
or U37943 (N_37943,N_36542,N_36447);
xor U37944 (N_37944,N_36395,N_36348);
and U37945 (N_37945,N_36817,N_36978);
and U37946 (N_37946,N_36313,N_36731);
nor U37947 (N_37947,N_36786,N_36644);
or U37948 (N_37948,N_36424,N_36096);
or U37949 (N_37949,N_36913,N_36023);
xor U37950 (N_37950,N_36300,N_36505);
xor U37951 (N_37951,N_36830,N_36051);
nand U37952 (N_37952,N_36996,N_36858);
nor U37953 (N_37953,N_36134,N_36009);
xor U37954 (N_37954,N_36832,N_36511);
or U37955 (N_37955,N_36642,N_36534);
and U37956 (N_37956,N_36151,N_36170);
and U37957 (N_37957,N_36615,N_36969);
or U37958 (N_37958,N_36912,N_36260);
nor U37959 (N_37959,N_36347,N_36994);
nor U37960 (N_37960,N_36657,N_36743);
or U37961 (N_37961,N_36855,N_36858);
or U37962 (N_37962,N_36167,N_36755);
xor U37963 (N_37963,N_36731,N_36702);
nor U37964 (N_37964,N_36134,N_36780);
nor U37965 (N_37965,N_36539,N_36551);
xnor U37966 (N_37966,N_36356,N_36538);
nand U37967 (N_37967,N_36259,N_36312);
xnor U37968 (N_37968,N_36865,N_36148);
nor U37969 (N_37969,N_36475,N_36906);
nor U37970 (N_37970,N_36224,N_36387);
nor U37971 (N_37971,N_36053,N_36815);
and U37972 (N_37972,N_36493,N_36788);
xnor U37973 (N_37973,N_36168,N_36960);
and U37974 (N_37974,N_36959,N_36492);
nor U37975 (N_37975,N_36973,N_36623);
nand U37976 (N_37976,N_36590,N_36328);
or U37977 (N_37977,N_36368,N_36403);
or U37978 (N_37978,N_36895,N_36672);
nand U37979 (N_37979,N_36584,N_36875);
and U37980 (N_37980,N_36374,N_36810);
xor U37981 (N_37981,N_36352,N_36789);
xor U37982 (N_37982,N_36593,N_36228);
nand U37983 (N_37983,N_36072,N_36380);
nand U37984 (N_37984,N_36279,N_36346);
nor U37985 (N_37985,N_36358,N_36227);
nor U37986 (N_37986,N_36240,N_36679);
nor U37987 (N_37987,N_36984,N_36319);
xnor U37988 (N_37988,N_36487,N_36890);
xnor U37989 (N_37989,N_36736,N_36272);
nor U37990 (N_37990,N_36904,N_36953);
or U37991 (N_37991,N_36367,N_36128);
and U37992 (N_37992,N_36662,N_36507);
xnor U37993 (N_37993,N_36213,N_36963);
or U37994 (N_37994,N_36886,N_36418);
nor U37995 (N_37995,N_36596,N_36924);
nor U37996 (N_37996,N_36475,N_36405);
and U37997 (N_37997,N_36882,N_36802);
nor U37998 (N_37998,N_36560,N_36587);
or U37999 (N_37999,N_36628,N_36838);
nor U38000 (N_38000,N_37508,N_37630);
nor U38001 (N_38001,N_37790,N_37114);
nor U38002 (N_38002,N_37202,N_37561);
or U38003 (N_38003,N_37125,N_37448);
or U38004 (N_38004,N_37690,N_37789);
nand U38005 (N_38005,N_37406,N_37310);
or U38006 (N_38006,N_37287,N_37305);
xor U38007 (N_38007,N_37215,N_37200);
nor U38008 (N_38008,N_37251,N_37421);
and U38009 (N_38009,N_37973,N_37979);
xor U38010 (N_38010,N_37138,N_37405);
xor U38011 (N_38011,N_37375,N_37959);
or U38012 (N_38012,N_37173,N_37850);
nor U38013 (N_38013,N_37218,N_37744);
and U38014 (N_38014,N_37782,N_37890);
nor U38015 (N_38015,N_37052,N_37196);
xor U38016 (N_38016,N_37739,N_37302);
xor U38017 (N_38017,N_37139,N_37460);
nor U38018 (N_38018,N_37669,N_37871);
xor U38019 (N_38019,N_37339,N_37128);
and U38020 (N_38020,N_37045,N_37100);
and U38021 (N_38021,N_37373,N_37926);
nor U38022 (N_38022,N_37293,N_37581);
and U38023 (N_38023,N_37262,N_37543);
and U38024 (N_38024,N_37442,N_37070);
or U38025 (N_38025,N_37802,N_37535);
nand U38026 (N_38026,N_37910,N_37384);
or U38027 (N_38027,N_37320,N_37133);
nor U38028 (N_38028,N_37121,N_37294);
nand U38029 (N_38029,N_37082,N_37837);
xor U38030 (N_38030,N_37076,N_37996);
or U38031 (N_38031,N_37435,N_37658);
xnor U38032 (N_38032,N_37967,N_37360);
or U38033 (N_38033,N_37015,N_37258);
nor U38034 (N_38034,N_37795,N_37368);
or U38035 (N_38035,N_37680,N_37597);
and U38036 (N_38036,N_37720,N_37924);
and U38037 (N_38037,N_37729,N_37160);
or U38038 (N_38038,N_37374,N_37985);
and U38039 (N_38039,N_37388,N_37483);
nand U38040 (N_38040,N_37162,N_37687);
or U38041 (N_38041,N_37370,N_37817);
and U38042 (N_38042,N_37205,N_37291);
nand U38043 (N_38043,N_37799,N_37267);
or U38044 (N_38044,N_37856,N_37638);
xor U38045 (N_38045,N_37635,N_37580);
xor U38046 (N_38046,N_37309,N_37932);
or U38047 (N_38047,N_37278,N_37949);
and U38048 (N_38048,N_37150,N_37812);
xor U38049 (N_38049,N_37351,N_37991);
or U38050 (N_38050,N_37766,N_37645);
nor U38051 (N_38051,N_37920,N_37214);
nor U38052 (N_38052,N_37326,N_37175);
xnor U38053 (N_38053,N_37718,N_37668);
xor U38054 (N_38054,N_37889,N_37145);
nor U38055 (N_38055,N_37292,N_37034);
nand U38056 (N_38056,N_37171,N_37598);
nand U38057 (N_38057,N_37830,N_37422);
and U38058 (N_38058,N_37409,N_37627);
xor U38059 (N_38059,N_37101,N_37230);
nand U38060 (N_38060,N_37964,N_37123);
nor U38061 (N_38061,N_37617,N_37037);
or U38062 (N_38062,N_37783,N_37178);
nand U38063 (N_38063,N_37960,N_37062);
nor U38064 (N_38064,N_37840,N_37747);
nor U38065 (N_38065,N_37445,N_37558);
or U38066 (N_38066,N_37963,N_37616);
or U38067 (N_38067,N_37698,N_37014);
nand U38068 (N_38068,N_37210,N_37024);
or U38069 (N_38069,N_37328,N_37084);
nand U38070 (N_38070,N_37233,N_37290);
nand U38071 (N_38071,N_37283,N_37689);
or U38072 (N_38072,N_37043,N_37134);
xor U38073 (N_38073,N_37023,N_37247);
nor U38074 (N_38074,N_37414,N_37455);
xor U38075 (N_38075,N_37793,N_37754);
xor U38076 (N_38076,N_37716,N_37717);
and U38077 (N_38077,N_37371,N_37877);
nand U38078 (N_38078,N_37000,N_37078);
xor U38079 (N_38079,N_37650,N_37190);
nor U38080 (N_38080,N_37462,N_37402);
or U38081 (N_38081,N_37161,N_37885);
nand U38082 (N_38082,N_37155,N_37059);
xnor U38083 (N_38083,N_37260,N_37018);
and U38084 (N_38084,N_37272,N_37304);
and U38085 (N_38085,N_37700,N_37397);
nor U38086 (N_38086,N_37723,N_37725);
nor U38087 (N_38087,N_37609,N_37987);
xnor U38088 (N_38088,N_37682,N_37343);
or U38089 (N_38089,N_37092,N_37334);
nand U38090 (N_38090,N_37636,N_37531);
or U38091 (N_38091,N_37412,N_37311);
nand U38092 (N_38092,N_37735,N_37324);
and U38093 (N_38093,N_37858,N_37463);
xor U38094 (N_38094,N_37146,N_37363);
nand U38095 (N_38095,N_37839,N_37629);
or U38096 (N_38096,N_37807,N_37358);
nor U38097 (N_38097,N_37095,N_37857);
or U38098 (N_38098,N_37673,N_37007);
nor U38099 (N_38099,N_37653,N_37104);
xor U38100 (N_38100,N_37234,N_37424);
and U38101 (N_38101,N_37042,N_37596);
and U38102 (N_38102,N_37742,N_37403);
or U38103 (N_38103,N_37534,N_37941);
or U38104 (N_38104,N_37117,N_37147);
nor U38105 (N_38105,N_37505,N_37301);
xnor U38106 (N_38106,N_37165,N_37613);
xnor U38107 (N_38107,N_37081,N_37524);
xor U38108 (N_38108,N_37073,N_37229);
nor U38109 (N_38109,N_37679,N_37235);
and U38110 (N_38110,N_37086,N_37168);
xnor U38111 (N_38111,N_37761,N_37903);
and U38112 (N_38112,N_37226,N_37347);
or U38113 (N_38113,N_37225,N_37986);
and U38114 (N_38114,N_37537,N_37096);
xor U38115 (N_38115,N_37437,N_37238);
nand U38116 (N_38116,N_37060,N_37038);
or U38117 (N_38117,N_37553,N_37297);
xnor U38118 (N_38118,N_37588,N_37286);
or U38119 (N_38119,N_37149,N_37240);
and U38120 (N_38120,N_37285,N_37798);
nand U38121 (N_38121,N_37589,N_37148);
and U38122 (N_38122,N_37672,N_37556);
or U38123 (N_38123,N_37900,N_37870);
nand U38124 (N_38124,N_37307,N_37825);
or U38125 (N_38125,N_37449,N_37407);
or U38126 (N_38126,N_37971,N_37352);
or U38127 (N_38127,N_37289,N_37400);
xor U38128 (N_38128,N_37132,N_37459);
and U38129 (N_38129,N_37726,N_37862);
nor U38130 (N_38130,N_37245,N_37264);
nor U38131 (N_38131,N_37486,N_37395);
or U38132 (N_38132,N_37451,N_37241);
nor U38133 (N_38133,N_37475,N_37612);
nand U38134 (N_38134,N_37620,N_37953);
or U38135 (N_38135,N_37333,N_37933);
nand U38136 (N_38136,N_37503,N_37860);
nand U38137 (N_38137,N_37992,N_37608);
and U38138 (N_38138,N_37341,N_37813);
and U38139 (N_38139,N_37622,N_37039);
xor U38140 (N_38140,N_37579,N_37182);
nor U38141 (N_38141,N_37502,N_37458);
xor U38142 (N_38142,N_37595,N_37480);
or U38143 (N_38143,N_37950,N_37053);
and U38144 (N_38144,N_37211,N_37425);
nand U38145 (N_38145,N_37821,N_37049);
nand U38146 (N_38146,N_37377,N_37787);
or U38147 (N_38147,N_37282,N_37509);
and U38148 (N_38148,N_37097,N_37895);
or U38149 (N_38149,N_37444,N_37583);
and U38150 (N_38150,N_37674,N_37863);
nand U38151 (N_38151,N_37441,N_37033);
nand U38152 (N_38152,N_37325,N_37781);
and U38153 (N_38153,N_37657,N_37917);
nand U38154 (N_38154,N_37083,N_37507);
nor U38155 (N_38155,N_37582,N_37186);
and U38156 (N_38156,N_37982,N_37847);
nor U38157 (N_38157,N_37016,N_37276);
nand U38158 (N_38158,N_37281,N_37231);
or U38159 (N_38159,N_37227,N_37841);
nor U38160 (N_38160,N_37521,N_37020);
nor U38161 (N_38161,N_37826,N_37851);
xor U38162 (N_38162,N_37499,N_37077);
nor U38163 (N_38163,N_37923,N_37576);
nand U38164 (N_38164,N_37482,N_37832);
nand U38165 (N_38165,N_37976,N_37506);
nand U38166 (N_38166,N_37275,N_37174);
nand U38167 (N_38167,N_37867,N_37143);
and U38168 (N_38168,N_37894,N_37786);
nor U38169 (N_38169,N_37244,N_37335);
xor U38170 (N_38170,N_37457,N_37488);
nor U38171 (N_38171,N_37124,N_37542);
xnor U38172 (N_38172,N_37193,N_37369);
or U38173 (N_38173,N_37661,N_37879);
or U38174 (N_38174,N_37330,N_37398);
xor U38175 (N_38175,N_37954,N_37257);
nor U38176 (N_38176,N_37731,N_37367);
or U38177 (N_38177,N_37710,N_37216);
and U38178 (N_38178,N_37426,N_37724);
and U38179 (N_38179,N_37965,N_37261);
or U38180 (N_38180,N_37834,N_37712);
or U38181 (N_38181,N_37471,N_37919);
xor U38182 (N_38182,N_37568,N_37207);
nand U38183 (N_38183,N_37329,N_37055);
xnor U38184 (N_38184,N_37899,N_37711);
and U38185 (N_38185,N_37664,N_37005);
xnor U38186 (N_38186,N_37936,N_37602);
or U38187 (N_38187,N_37772,N_37063);
xnor U38188 (N_38188,N_37741,N_37577);
and U38189 (N_38189,N_37896,N_37232);
and U38190 (N_38190,N_37280,N_37915);
xnor U38191 (N_38191,N_37788,N_37935);
and U38192 (N_38192,N_37571,N_37319);
nor U38193 (N_38193,N_37028,N_37852);
xnor U38194 (N_38194,N_37454,N_37494);
nand U38195 (N_38195,N_37088,N_37983);
or U38196 (N_38196,N_37203,N_37818);
nand U38197 (N_38197,N_37469,N_37476);
xor U38198 (N_38198,N_37764,N_37519);
or U38199 (N_38199,N_37662,N_37686);
nand U38200 (N_38200,N_37219,N_37559);
xnor U38201 (N_38201,N_37916,N_37390);
or U38202 (N_38202,N_37520,N_37404);
or U38203 (N_38203,N_37030,N_37771);
and U38204 (N_38204,N_37575,N_37614);
or U38205 (N_38205,N_37794,N_37756);
and U38206 (N_38206,N_37498,N_37237);
nand U38207 (N_38207,N_37431,N_37908);
nand U38208 (N_38208,N_37671,N_37928);
xnor U38209 (N_38209,N_37365,N_37881);
nand U38210 (N_38210,N_37665,N_37943);
nor U38211 (N_38211,N_37995,N_37937);
nor U38212 (N_38212,N_37541,N_37012);
and U38213 (N_38213,N_37882,N_37317);
xnor U38214 (N_38214,N_37906,N_37417);
or U38215 (N_38215,N_37064,N_37532);
or U38216 (N_38216,N_37591,N_37633);
nand U38217 (N_38217,N_37172,N_37872);
or U38218 (N_38218,N_37838,N_37113);
or U38219 (N_38219,N_37270,N_37607);
or U38220 (N_38220,N_37031,N_37530);
nand U38221 (N_38221,N_37001,N_37562);
nor U38222 (N_38222,N_37316,N_37691);
xnor U38223 (N_38223,N_37094,N_37372);
nand U38224 (N_38224,N_37713,N_37255);
or U38225 (N_38225,N_37696,N_37981);
xor U38226 (N_38226,N_37708,N_37643);
nor U38227 (N_38227,N_37748,N_37246);
nand U38228 (N_38228,N_37606,N_37484);
nor U38229 (N_38229,N_37815,N_37808);
xor U38230 (N_38230,N_37224,N_37874);
or U38231 (N_38231,N_37027,N_37056);
and U38232 (N_38232,N_37875,N_37618);
or U38233 (N_38233,N_37141,N_37888);
nand U38234 (N_38234,N_37318,N_37652);
or U38235 (N_38235,N_37169,N_37939);
and U38236 (N_38236,N_37050,N_37192);
or U38237 (N_38237,N_37660,N_37699);
nand U38238 (N_38238,N_37465,N_37675);
or U38239 (N_38239,N_37855,N_37135);
nor U38240 (N_38240,N_37129,N_37925);
xnor U38241 (N_38241,N_37599,N_37099);
nor U38242 (N_38242,N_37468,N_37345);
nor U38243 (N_38243,N_37732,N_37880);
and U38244 (N_38244,N_37719,N_37853);
xnor U38245 (N_38245,N_37416,N_37655);
or U38246 (N_38246,N_37510,N_37762);
xnor U38247 (N_38247,N_37952,N_37470);
xnor U38248 (N_38248,N_37683,N_37144);
nand U38249 (N_38249,N_37479,N_37564);
and U38250 (N_38250,N_37958,N_37298);
nor U38251 (N_38251,N_37868,N_37394);
nand U38252 (N_38252,N_37284,N_37151);
nand U38253 (N_38253,N_37103,N_37355);
and U38254 (N_38254,N_37829,N_37512);
or U38255 (N_38255,N_37946,N_37300);
and U38256 (N_38256,N_37918,N_37977);
or U38257 (N_38257,N_37632,N_37859);
xor U38258 (N_38258,N_37586,N_37566);
and U38259 (N_38259,N_37265,N_37040);
nand U38260 (N_38260,N_37127,N_37998);
xnor U38261 (N_38261,N_37474,N_37640);
and U38262 (N_38262,N_37773,N_37517);
nor U38263 (N_38263,N_37487,N_37697);
and U38264 (N_38264,N_37126,N_37704);
nor U38265 (N_38265,N_37544,N_37107);
xnor U38266 (N_38266,N_37259,N_37277);
and U38267 (N_38267,N_37252,N_37644);
or U38268 (N_38268,N_37934,N_37188);
nand U38269 (N_38269,N_37849,N_37993);
nor U38270 (N_38270,N_37945,N_37051);
xnor U38271 (N_38271,N_37730,N_37760);
nand U38272 (N_38272,N_37728,N_37386);
or U38273 (N_38273,N_37947,N_37538);
xor U38274 (N_38274,N_37864,N_37550);
and U38275 (N_38275,N_37824,N_37770);
xnor U38276 (N_38276,N_37119,N_37041);
nor U38277 (N_38277,N_37912,N_37651);
or U38278 (N_38278,N_37769,N_37274);
or U38279 (N_38279,N_37752,N_37438);
nand U38280 (N_38280,N_37389,N_37180);
nor U38281 (N_38281,N_37466,N_37009);
xnor U38282 (N_38282,N_37288,N_37540);
xor U38283 (N_38283,N_37164,N_37750);
nand U38284 (N_38284,N_37604,N_37670);
xnor U38285 (N_38285,N_37784,N_37927);
xnor U38286 (N_38286,N_37153,N_37740);
xnor U38287 (N_38287,N_37694,N_37376);
xnor U38288 (N_38288,N_37022,N_37842);
nand U38289 (N_38289,N_37554,N_37322);
and U38290 (N_38290,N_37551,N_37066);
and U38291 (N_38291,N_37299,N_37057);
nand U38292 (N_38292,N_37843,N_37380);
nand U38293 (N_38293,N_37089,N_37797);
nor U38294 (N_38294,N_37206,N_37810);
nor U38295 (N_38295,N_37831,N_37156);
and U38296 (N_38296,N_37191,N_37197);
nand U38297 (N_38297,N_37922,N_37387);
or U38298 (N_38298,N_37961,N_37378);
nor U38299 (N_38299,N_37972,N_37044);
xor U38300 (N_38300,N_37481,N_37090);
or U38301 (N_38301,N_37067,N_37514);
and U38302 (N_38302,N_37603,N_37496);
nand U38303 (N_38303,N_37828,N_37243);
nand U38304 (N_38304,N_37570,N_37736);
or U38305 (N_38305,N_37511,N_37080);
and U38306 (N_38306,N_37692,N_37836);
or U38307 (N_38307,N_37108,N_37248);
xnor U38308 (N_38308,N_37295,N_37615);
nor U38309 (N_38309,N_37684,N_37321);
xnor U38310 (N_38310,N_37268,N_37814);
or U38311 (N_38311,N_37199,N_37833);
nor U38312 (N_38312,N_37573,N_37647);
and U38313 (N_38313,N_37179,N_37962);
and U38314 (N_38314,N_37765,N_37228);
or U38315 (N_38315,N_37217,N_37356);
or U38316 (N_38316,N_37883,N_37068);
nand U38317 (N_38317,N_37212,N_37659);
and U38318 (N_38318,N_37379,N_37137);
xnor U38319 (N_38319,N_37796,N_37427);
or U38320 (N_38320,N_37746,N_37048);
and U38321 (N_38321,N_37419,N_37734);
or U38322 (N_38322,N_37637,N_37485);
and U38323 (N_38323,N_37353,N_37625);
and U38324 (N_38324,N_37755,N_37695);
and U38325 (N_38325,N_37102,N_37663);
nor U38326 (N_38326,N_37533,N_37036);
xor U38327 (N_38327,N_37021,N_37118);
nor U38328 (N_38328,N_37213,N_37806);
nand U38329 (N_38329,N_37563,N_37779);
and U38330 (N_38330,N_37715,N_37816);
nor U38331 (N_38331,N_37430,N_37701);
nand U38332 (N_38332,N_37071,N_37970);
or U38333 (N_38333,N_37269,N_37011);
nor U38334 (N_38334,N_37823,N_37029);
xnor U38335 (N_38335,N_37087,N_37768);
or U38336 (N_38336,N_37342,N_37116);
and U38337 (N_38337,N_37504,N_37142);
nor U38338 (N_38338,N_37396,N_37593);
xor U38339 (N_38339,N_37236,N_37536);
nor U38340 (N_38340,N_37477,N_37110);
or U38341 (N_38341,N_37980,N_37529);
and U38342 (N_38342,N_37434,N_37677);
xnor U38343 (N_38343,N_37338,N_37778);
or U38344 (N_38344,N_37428,N_37693);
nand U38345 (N_38345,N_37418,N_37994);
or U38346 (N_38346,N_37239,N_37974);
xnor U38347 (N_38347,N_37938,N_37707);
nand U38348 (N_38348,N_37845,N_37775);
nand U38349 (N_38349,N_37361,N_37767);
or U38350 (N_38350,N_37271,N_37523);
nor U38351 (N_38351,N_37364,N_37822);
and U38352 (N_38352,N_37399,N_37605);
xnor U38353 (N_38353,N_37835,N_37911);
nor U38354 (N_38354,N_37685,N_37515);
nor U38355 (N_38355,N_37120,N_37930);
nand U38356 (N_38356,N_37909,N_37263);
nor U38357 (N_38357,N_37348,N_37303);
or U38358 (N_38358,N_37452,N_37522);
or U38359 (N_38359,N_37641,N_37047);
nor U38360 (N_38360,N_37177,N_37167);
nor U38361 (N_38361,N_37791,N_37619);
nor U38362 (N_38362,N_37446,N_37350);
and U38363 (N_38363,N_37955,N_37774);
and U38364 (N_38364,N_37944,N_37489);
or U38365 (N_38365,N_37914,N_37327);
or U38366 (N_38366,N_37002,N_37032);
and U38367 (N_38367,N_37183,N_37223);
nand U38368 (N_38368,N_37450,N_37978);
nand U38369 (N_38369,N_37065,N_37157);
and U38370 (N_38370,N_37166,N_37743);
and U38371 (N_38371,N_37061,N_37552);
and U38372 (N_38372,N_37600,N_37306);
nand U38373 (N_38373,N_37337,N_37539);
nand U38374 (N_38374,N_37314,N_37194);
or U38375 (N_38375,N_37195,N_37861);
nor U38376 (N_38376,N_37654,N_37869);
nor U38377 (N_38377,N_37130,N_37279);
xnor U38378 (N_38378,N_37344,N_37079);
nor U38379 (N_38379,N_37984,N_37154);
nor U38380 (N_38380,N_37098,N_37359);
and U38381 (N_38381,N_37159,N_37703);
or U38382 (N_38382,N_37560,N_37528);
nor U38383 (N_38383,N_37567,N_37516);
nor U38384 (N_38384,N_37366,N_37313);
nor U38385 (N_38385,N_37093,N_37585);
or U38386 (N_38386,N_37323,N_37545);
nand U38387 (N_38387,N_37006,N_37525);
nor U38388 (N_38388,N_37844,N_37003);
xor U38389 (N_38389,N_37792,N_37131);
nand U38390 (N_38390,N_37158,N_37969);
nand U38391 (N_38391,N_37688,N_37827);
or U38392 (N_38392,N_37546,N_37601);
xor U38393 (N_38393,N_37204,N_37803);
nand U38394 (N_38394,N_37242,N_37315);
or U38395 (N_38395,N_37667,N_37737);
xor U38396 (N_38396,N_37572,N_37420);
nor U38397 (N_38397,N_37758,N_37848);
nor U38398 (N_38398,N_37109,N_37892);
nor U38399 (N_38399,N_37751,N_37383);
and U38400 (N_38400,N_37495,N_37456);
and U38401 (N_38401,N_37745,N_37642);
xor U38402 (N_38402,N_37738,N_37312);
nor U38403 (N_38403,N_37907,N_37902);
nor U38404 (N_38404,N_37501,N_37122);
and U38405 (N_38405,N_37999,N_37163);
nand U38406 (N_38406,N_37631,N_37112);
nor U38407 (N_38407,N_37025,N_37733);
nor U38408 (N_38408,N_37547,N_37819);
nand U38409 (N_38409,N_37187,N_37209);
nand U38410 (N_38410,N_37185,N_37308);
and U38411 (N_38411,N_37478,N_37526);
nand U38412 (N_38412,N_37273,N_37727);
nor U38413 (N_38413,N_37436,N_37492);
nand U38414 (N_38414,N_37921,N_37942);
nor U38415 (N_38415,N_37891,N_37464);
and U38416 (N_38416,N_37336,N_37256);
xor U38417 (N_38417,N_37447,N_37759);
and U38418 (N_38418,N_37249,N_37401);
nand U38419 (N_38419,N_37646,N_37415);
or U38420 (N_38420,N_37574,N_37549);
and U38421 (N_38421,N_37865,N_37811);
nor U38422 (N_38422,N_37220,N_37493);
and U38423 (N_38423,N_37610,N_37809);
xor U38424 (N_38424,N_37777,N_37634);
nor U38425 (N_38425,N_37975,N_37439);
xnor U38426 (N_38426,N_37072,N_37940);
xnor U38427 (N_38427,N_37152,N_37136);
nor U38428 (N_38428,N_37678,N_37931);
nand U38429 (N_38429,N_37461,N_37432);
nor U38430 (N_38430,N_37988,N_37929);
or U38431 (N_38431,N_37221,N_37648);
nor U38432 (N_38432,N_37578,N_37587);
nand U38433 (N_38433,N_37332,N_37354);
and U38434 (N_38434,N_37656,N_37472);
xnor U38435 (N_38435,N_37189,N_37820);
and U38436 (N_38436,N_37990,N_37013);
nand U38437 (N_38437,N_37069,N_37649);
and U38438 (N_38438,N_37413,N_37440);
nand U38439 (N_38439,N_37893,N_37019);
and U38440 (N_38440,N_37391,N_37592);
nor U38441 (N_38441,N_37709,N_37074);
xor U38442 (N_38442,N_37611,N_37250);
nor U38443 (N_38443,N_37091,N_37004);
or U38444 (N_38444,N_37753,N_37548);
and U38445 (N_38445,N_37594,N_37876);
xnor U38446 (N_38446,N_37951,N_37026);
nor U38447 (N_38447,N_37222,N_37898);
nand U38448 (N_38448,N_37046,N_37058);
nor U38449 (N_38449,N_37331,N_37886);
nand U38450 (N_38450,N_37721,N_37854);
xor U38451 (N_38451,N_37557,N_37410);
and U38452 (N_38452,N_37681,N_37757);
and U38453 (N_38453,N_37381,N_37490);
or U38454 (N_38454,N_37968,N_37500);
nor U38455 (N_38455,N_37866,N_37800);
or U38456 (N_38456,N_37702,N_37075);
or U38457 (N_38457,N_37555,N_37513);
or U38458 (N_38458,N_37357,N_37714);
and U38459 (N_38459,N_37846,N_37584);
xor U38460 (N_38460,N_37904,N_37054);
nor U38461 (N_38461,N_37106,N_37997);
nand U38462 (N_38462,N_37010,N_37254);
xor U38463 (N_38463,N_37801,N_37497);
xor U38464 (N_38464,N_37035,N_37623);
xnor U38465 (N_38465,N_37198,N_37749);
nand U38466 (N_38466,N_37362,N_37666);
and U38467 (N_38467,N_37266,N_37780);
nor U38468 (N_38468,N_37349,N_37624);
and U38469 (N_38469,N_37385,N_37411);
and U38470 (N_38470,N_37170,N_37491);
nor U38471 (N_38471,N_37346,N_37392);
nand U38472 (N_38472,N_37966,N_37393);
or U38473 (N_38473,N_37473,N_37296);
nor U38474 (N_38474,N_37467,N_37176);
xnor U38475 (N_38475,N_37706,N_37085);
nor U38476 (N_38476,N_37115,N_37382);
nor U38477 (N_38477,N_37639,N_37776);
xnor U38478 (N_38478,N_37956,N_37340);
and U38479 (N_38479,N_37453,N_37181);
or U38480 (N_38480,N_37008,N_37948);
nor U38481 (N_38481,N_37905,N_37989);
xor U38482 (N_38482,N_37722,N_37111);
or U38483 (N_38483,N_37626,N_37913);
and U38484 (N_38484,N_37804,N_37805);
nand U38485 (N_38485,N_37884,N_37878);
or U38486 (N_38486,N_37201,N_37763);
xor U38487 (N_38487,N_37565,N_37705);
nand U38488 (N_38488,N_37621,N_37590);
and U38489 (N_38489,N_37527,N_37628);
and U38490 (N_38490,N_37208,N_37901);
nand U38491 (N_38491,N_37518,N_37433);
nand U38492 (N_38492,N_37423,N_37443);
nand U38493 (N_38493,N_37887,N_37408);
or U38494 (N_38494,N_37253,N_37429);
and U38495 (N_38495,N_37017,N_37569);
and U38496 (N_38496,N_37140,N_37676);
or U38497 (N_38497,N_37105,N_37184);
or U38498 (N_38498,N_37873,N_37897);
nor U38499 (N_38499,N_37957,N_37785);
nor U38500 (N_38500,N_37502,N_37026);
and U38501 (N_38501,N_37789,N_37539);
and U38502 (N_38502,N_37136,N_37492);
and U38503 (N_38503,N_37580,N_37419);
or U38504 (N_38504,N_37947,N_37893);
nand U38505 (N_38505,N_37085,N_37484);
nor U38506 (N_38506,N_37622,N_37835);
or U38507 (N_38507,N_37714,N_37932);
xor U38508 (N_38508,N_37888,N_37464);
nor U38509 (N_38509,N_37928,N_37164);
xnor U38510 (N_38510,N_37536,N_37430);
nor U38511 (N_38511,N_37709,N_37012);
nor U38512 (N_38512,N_37675,N_37092);
nor U38513 (N_38513,N_37411,N_37484);
nor U38514 (N_38514,N_37076,N_37983);
nand U38515 (N_38515,N_37696,N_37468);
or U38516 (N_38516,N_37617,N_37956);
xor U38517 (N_38517,N_37845,N_37966);
nand U38518 (N_38518,N_37306,N_37216);
or U38519 (N_38519,N_37276,N_37084);
nor U38520 (N_38520,N_37939,N_37280);
or U38521 (N_38521,N_37598,N_37875);
nand U38522 (N_38522,N_37471,N_37309);
nand U38523 (N_38523,N_37890,N_37450);
nand U38524 (N_38524,N_37458,N_37407);
xnor U38525 (N_38525,N_37104,N_37385);
or U38526 (N_38526,N_37704,N_37644);
and U38527 (N_38527,N_37329,N_37758);
and U38528 (N_38528,N_37089,N_37126);
or U38529 (N_38529,N_37017,N_37258);
and U38530 (N_38530,N_37338,N_37805);
nand U38531 (N_38531,N_37072,N_37557);
nand U38532 (N_38532,N_37844,N_37696);
xnor U38533 (N_38533,N_37741,N_37139);
or U38534 (N_38534,N_37923,N_37077);
xor U38535 (N_38535,N_37075,N_37556);
or U38536 (N_38536,N_37559,N_37080);
or U38537 (N_38537,N_37339,N_37436);
and U38538 (N_38538,N_37256,N_37960);
xnor U38539 (N_38539,N_37436,N_37040);
nand U38540 (N_38540,N_37368,N_37019);
xor U38541 (N_38541,N_37253,N_37224);
nand U38542 (N_38542,N_37188,N_37768);
or U38543 (N_38543,N_37174,N_37734);
nand U38544 (N_38544,N_37670,N_37505);
xor U38545 (N_38545,N_37010,N_37850);
xnor U38546 (N_38546,N_37364,N_37488);
nand U38547 (N_38547,N_37560,N_37251);
nand U38548 (N_38548,N_37844,N_37263);
xnor U38549 (N_38549,N_37896,N_37853);
xnor U38550 (N_38550,N_37570,N_37540);
nand U38551 (N_38551,N_37252,N_37648);
nor U38552 (N_38552,N_37207,N_37350);
nor U38553 (N_38553,N_37550,N_37641);
nand U38554 (N_38554,N_37009,N_37489);
or U38555 (N_38555,N_37674,N_37604);
xnor U38556 (N_38556,N_37134,N_37916);
xor U38557 (N_38557,N_37242,N_37786);
nand U38558 (N_38558,N_37305,N_37925);
xor U38559 (N_38559,N_37001,N_37830);
nand U38560 (N_38560,N_37642,N_37713);
or U38561 (N_38561,N_37274,N_37574);
and U38562 (N_38562,N_37313,N_37561);
nor U38563 (N_38563,N_37701,N_37723);
or U38564 (N_38564,N_37847,N_37388);
nor U38565 (N_38565,N_37130,N_37913);
and U38566 (N_38566,N_37081,N_37162);
xnor U38567 (N_38567,N_37091,N_37620);
and U38568 (N_38568,N_37533,N_37563);
nand U38569 (N_38569,N_37313,N_37327);
and U38570 (N_38570,N_37528,N_37439);
or U38571 (N_38571,N_37557,N_37148);
nor U38572 (N_38572,N_37962,N_37564);
or U38573 (N_38573,N_37734,N_37478);
xor U38574 (N_38574,N_37757,N_37875);
nor U38575 (N_38575,N_37459,N_37942);
and U38576 (N_38576,N_37597,N_37939);
or U38577 (N_38577,N_37111,N_37702);
or U38578 (N_38578,N_37579,N_37242);
nand U38579 (N_38579,N_37426,N_37425);
xor U38580 (N_38580,N_37957,N_37379);
nor U38581 (N_38581,N_37055,N_37251);
or U38582 (N_38582,N_37461,N_37439);
and U38583 (N_38583,N_37062,N_37724);
and U38584 (N_38584,N_37689,N_37342);
xor U38585 (N_38585,N_37917,N_37564);
and U38586 (N_38586,N_37189,N_37632);
and U38587 (N_38587,N_37438,N_37173);
nand U38588 (N_38588,N_37228,N_37515);
or U38589 (N_38589,N_37933,N_37266);
and U38590 (N_38590,N_37530,N_37037);
nor U38591 (N_38591,N_37834,N_37655);
or U38592 (N_38592,N_37552,N_37306);
or U38593 (N_38593,N_37076,N_37969);
or U38594 (N_38594,N_37900,N_37246);
and U38595 (N_38595,N_37882,N_37181);
and U38596 (N_38596,N_37992,N_37722);
and U38597 (N_38597,N_37056,N_37757);
nor U38598 (N_38598,N_37382,N_37082);
nand U38599 (N_38599,N_37531,N_37346);
or U38600 (N_38600,N_37627,N_37609);
or U38601 (N_38601,N_37328,N_37771);
xor U38602 (N_38602,N_37664,N_37870);
nor U38603 (N_38603,N_37775,N_37390);
or U38604 (N_38604,N_37511,N_37266);
xnor U38605 (N_38605,N_37192,N_37644);
nor U38606 (N_38606,N_37543,N_37947);
and U38607 (N_38607,N_37211,N_37646);
or U38608 (N_38608,N_37075,N_37186);
and U38609 (N_38609,N_37247,N_37567);
or U38610 (N_38610,N_37089,N_37774);
and U38611 (N_38611,N_37562,N_37302);
xnor U38612 (N_38612,N_37089,N_37983);
nor U38613 (N_38613,N_37367,N_37202);
nor U38614 (N_38614,N_37400,N_37584);
or U38615 (N_38615,N_37245,N_37982);
or U38616 (N_38616,N_37450,N_37918);
nor U38617 (N_38617,N_37887,N_37826);
xor U38618 (N_38618,N_37954,N_37331);
or U38619 (N_38619,N_37295,N_37386);
and U38620 (N_38620,N_37781,N_37490);
nand U38621 (N_38621,N_37494,N_37297);
nand U38622 (N_38622,N_37406,N_37885);
or U38623 (N_38623,N_37990,N_37996);
xor U38624 (N_38624,N_37177,N_37897);
or U38625 (N_38625,N_37252,N_37300);
and U38626 (N_38626,N_37814,N_37656);
nand U38627 (N_38627,N_37396,N_37605);
xor U38628 (N_38628,N_37903,N_37650);
nor U38629 (N_38629,N_37944,N_37316);
nand U38630 (N_38630,N_37351,N_37127);
nor U38631 (N_38631,N_37317,N_37926);
xor U38632 (N_38632,N_37874,N_37475);
xnor U38633 (N_38633,N_37438,N_37561);
xor U38634 (N_38634,N_37156,N_37426);
and U38635 (N_38635,N_37911,N_37791);
or U38636 (N_38636,N_37230,N_37494);
xor U38637 (N_38637,N_37110,N_37832);
or U38638 (N_38638,N_37594,N_37745);
and U38639 (N_38639,N_37059,N_37906);
xnor U38640 (N_38640,N_37079,N_37549);
nand U38641 (N_38641,N_37312,N_37148);
xnor U38642 (N_38642,N_37205,N_37485);
nand U38643 (N_38643,N_37606,N_37337);
nor U38644 (N_38644,N_37572,N_37781);
and U38645 (N_38645,N_37911,N_37590);
or U38646 (N_38646,N_37144,N_37312);
nand U38647 (N_38647,N_37345,N_37600);
nor U38648 (N_38648,N_37417,N_37351);
nand U38649 (N_38649,N_37916,N_37167);
nor U38650 (N_38650,N_37185,N_37677);
and U38651 (N_38651,N_37683,N_37278);
nand U38652 (N_38652,N_37495,N_37378);
nor U38653 (N_38653,N_37094,N_37686);
nand U38654 (N_38654,N_37221,N_37085);
nand U38655 (N_38655,N_37106,N_37315);
and U38656 (N_38656,N_37160,N_37347);
and U38657 (N_38657,N_37669,N_37888);
or U38658 (N_38658,N_37832,N_37935);
and U38659 (N_38659,N_37660,N_37376);
nor U38660 (N_38660,N_37215,N_37169);
nor U38661 (N_38661,N_37555,N_37759);
or U38662 (N_38662,N_37033,N_37891);
xnor U38663 (N_38663,N_37414,N_37578);
nand U38664 (N_38664,N_37958,N_37990);
nor U38665 (N_38665,N_37095,N_37060);
xnor U38666 (N_38666,N_37330,N_37865);
and U38667 (N_38667,N_37914,N_37753);
xor U38668 (N_38668,N_37202,N_37179);
and U38669 (N_38669,N_37729,N_37782);
and U38670 (N_38670,N_37633,N_37733);
nor U38671 (N_38671,N_37049,N_37782);
and U38672 (N_38672,N_37396,N_37194);
and U38673 (N_38673,N_37555,N_37090);
or U38674 (N_38674,N_37661,N_37884);
or U38675 (N_38675,N_37398,N_37214);
xnor U38676 (N_38676,N_37589,N_37057);
xor U38677 (N_38677,N_37040,N_37450);
or U38678 (N_38678,N_37623,N_37040);
or U38679 (N_38679,N_37030,N_37857);
and U38680 (N_38680,N_37915,N_37539);
or U38681 (N_38681,N_37994,N_37781);
nor U38682 (N_38682,N_37597,N_37248);
xnor U38683 (N_38683,N_37608,N_37984);
and U38684 (N_38684,N_37285,N_37384);
nand U38685 (N_38685,N_37802,N_37840);
nor U38686 (N_38686,N_37499,N_37434);
and U38687 (N_38687,N_37508,N_37911);
and U38688 (N_38688,N_37757,N_37703);
nand U38689 (N_38689,N_37852,N_37970);
or U38690 (N_38690,N_37332,N_37878);
xnor U38691 (N_38691,N_37133,N_37977);
and U38692 (N_38692,N_37951,N_37014);
and U38693 (N_38693,N_37336,N_37998);
nand U38694 (N_38694,N_37656,N_37652);
nand U38695 (N_38695,N_37026,N_37662);
xor U38696 (N_38696,N_37398,N_37921);
nand U38697 (N_38697,N_37666,N_37411);
xnor U38698 (N_38698,N_37789,N_37779);
or U38699 (N_38699,N_37675,N_37632);
nand U38700 (N_38700,N_37822,N_37830);
nand U38701 (N_38701,N_37406,N_37984);
nor U38702 (N_38702,N_37992,N_37925);
xnor U38703 (N_38703,N_37476,N_37282);
and U38704 (N_38704,N_37190,N_37003);
and U38705 (N_38705,N_37097,N_37675);
and U38706 (N_38706,N_37786,N_37413);
or U38707 (N_38707,N_37859,N_37608);
xnor U38708 (N_38708,N_37006,N_37614);
nand U38709 (N_38709,N_37838,N_37696);
and U38710 (N_38710,N_37076,N_37992);
xor U38711 (N_38711,N_37624,N_37402);
or U38712 (N_38712,N_37770,N_37345);
nor U38713 (N_38713,N_37192,N_37509);
xnor U38714 (N_38714,N_37648,N_37507);
and U38715 (N_38715,N_37557,N_37011);
nor U38716 (N_38716,N_37219,N_37814);
and U38717 (N_38717,N_37903,N_37505);
and U38718 (N_38718,N_37615,N_37856);
or U38719 (N_38719,N_37468,N_37936);
xnor U38720 (N_38720,N_37454,N_37165);
or U38721 (N_38721,N_37092,N_37155);
xor U38722 (N_38722,N_37450,N_37526);
and U38723 (N_38723,N_37171,N_37523);
nand U38724 (N_38724,N_37111,N_37221);
nand U38725 (N_38725,N_37631,N_37009);
nor U38726 (N_38726,N_37324,N_37082);
or U38727 (N_38727,N_37392,N_37830);
and U38728 (N_38728,N_37806,N_37020);
nor U38729 (N_38729,N_37539,N_37796);
and U38730 (N_38730,N_37805,N_37742);
and U38731 (N_38731,N_37307,N_37701);
xor U38732 (N_38732,N_37260,N_37289);
and U38733 (N_38733,N_37966,N_37354);
nand U38734 (N_38734,N_37732,N_37444);
or U38735 (N_38735,N_37046,N_37397);
nor U38736 (N_38736,N_37173,N_37485);
and U38737 (N_38737,N_37636,N_37199);
xor U38738 (N_38738,N_37898,N_37692);
xor U38739 (N_38739,N_37094,N_37515);
or U38740 (N_38740,N_37745,N_37207);
and U38741 (N_38741,N_37004,N_37448);
xor U38742 (N_38742,N_37545,N_37889);
xnor U38743 (N_38743,N_37662,N_37819);
xnor U38744 (N_38744,N_37749,N_37599);
and U38745 (N_38745,N_37112,N_37733);
nand U38746 (N_38746,N_37103,N_37748);
or U38747 (N_38747,N_37416,N_37262);
and U38748 (N_38748,N_37396,N_37462);
or U38749 (N_38749,N_37301,N_37415);
and U38750 (N_38750,N_37140,N_37993);
and U38751 (N_38751,N_37664,N_37536);
or U38752 (N_38752,N_37352,N_37191);
xor U38753 (N_38753,N_37841,N_37940);
xor U38754 (N_38754,N_37786,N_37303);
xor U38755 (N_38755,N_37541,N_37409);
or U38756 (N_38756,N_37633,N_37738);
or U38757 (N_38757,N_37046,N_37347);
or U38758 (N_38758,N_37154,N_37504);
nand U38759 (N_38759,N_37768,N_37186);
or U38760 (N_38760,N_37613,N_37537);
nand U38761 (N_38761,N_37162,N_37993);
xor U38762 (N_38762,N_37127,N_37937);
nand U38763 (N_38763,N_37521,N_37665);
or U38764 (N_38764,N_37702,N_37078);
and U38765 (N_38765,N_37832,N_37541);
nand U38766 (N_38766,N_37433,N_37460);
nor U38767 (N_38767,N_37665,N_37607);
or U38768 (N_38768,N_37522,N_37416);
xor U38769 (N_38769,N_37010,N_37383);
nand U38770 (N_38770,N_37475,N_37691);
xnor U38771 (N_38771,N_37796,N_37326);
nor U38772 (N_38772,N_37805,N_37836);
nor U38773 (N_38773,N_37992,N_37931);
nand U38774 (N_38774,N_37292,N_37029);
and U38775 (N_38775,N_37300,N_37135);
nor U38776 (N_38776,N_37336,N_37157);
nor U38777 (N_38777,N_37316,N_37180);
nor U38778 (N_38778,N_37654,N_37523);
or U38779 (N_38779,N_37138,N_37665);
nand U38780 (N_38780,N_37159,N_37065);
xnor U38781 (N_38781,N_37674,N_37056);
or U38782 (N_38782,N_37137,N_37850);
and U38783 (N_38783,N_37782,N_37267);
xnor U38784 (N_38784,N_37367,N_37093);
or U38785 (N_38785,N_37493,N_37389);
nor U38786 (N_38786,N_37546,N_37162);
nor U38787 (N_38787,N_37130,N_37982);
xor U38788 (N_38788,N_37895,N_37983);
nor U38789 (N_38789,N_37603,N_37800);
and U38790 (N_38790,N_37428,N_37503);
nor U38791 (N_38791,N_37299,N_37004);
xor U38792 (N_38792,N_37833,N_37115);
or U38793 (N_38793,N_37353,N_37671);
or U38794 (N_38794,N_37240,N_37707);
nand U38795 (N_38795,N_37212,N_37841);
nand U38796 (N_38796,N_37894,N_37576);
nor U38797 (N_38797,N_37913,N_37883);
and U38798 (N_38798,N_37859,N_37604);
or U38799 (N_38799,N_37053,N_37675);
nand U38800 (N_38800,N_37841,N_37584);
nor U38801 (N_38801,N_37837,N_37626);
or U38802 (N_38802,N_37558,N_37903);
or U38803 (N_38803,N_37409,N_37215);
xnor U38804 (N_38804,N_37966,N_37623);
or U38805 (N_38805,N_37204,N_37459);
nor U38806 (N_38806,N_37472,N_37075);
or U38807 (N_38807,N_37572,N_37993);
nor U38808 (N_38808,N_37364,N_37769);
xor U38809 (N_38809,N_37474,N_37176);
xnor U38810 (N_38810,N_37672,N_37294);
and U38811 (N_38811,N_37842,N_37293);
nand U38812 (N_38812,N_37838,N_37426);
and U38813 (N_38813,N_37280,N_37307);
or U38814 (N_38814,N_37446,N_37699);
nor U38815 (N_38815,N_37192,N_37886);
xnor U38816 (N_38816,N_37276,N_37937);
and U38817 (N_38817,N_37508,N_37905);
xor U38818 (N_38818,N_37223,N_37651);
and U38819 (N_38819,N_37825,N_37987);
nor U38820 (N_38820,N_37254,N_37046);
xnor U38821 (N_38821,N_37940,N_37896);
and U38822 (N_38822,N_37470,N_37319);
or U38823 (N_38823,N_37548,N_37211);
and U38824 (N_38824,N_37746,N_37889);
or U38825 (N_38825,N_37868,N_37863);
or U38826 (N_38826,N_37816,N_37183);
and U38827 (N_38827,N_37493,N_37917);
nor U38828 (N_38828,N_37088,N_37581);
or U38829 (N_38829,N_37285,N_37689);
xnor U38830 (N_38830,N_37641,N_37562);
nand U38831 (N_38831,N_37249,N_37326);
or U38832 (N_38832,N_37099,N_37428);
and U38833 (N_38833,N_37739,N_37026);
or U38834 (N_38834,N_37914,N_37890);
nor U38835 (N_38835,N_37960,N_37196);
xor U38836 (N_38836,N_37279,N_37529);
xor U38837 (N_38837,N_37391,N_37540);
or U38838 (N_38838,N_37815,N_37792);
and U38839 (N_38839,N_37040,N_37646);
nor U38840 (N_38840,N_37863,N_37837);
nor U38841 (N_38841,N_37411,N_37984);
nor U38842 (N_38842,N_37891,N_37118);
and U38843 (N_38843,N_37108,N_37147);
nor U38844 (N_38844,N_37958,N_37476);
and U38845 (N_38845,N_37555,N_37929);
and U38846 (N_38846,N_37454,N_37727);
or U38847 (N_38847,N_37231,N_37559);
nor U38848 (N_38848,N_37813,N_37410);
nor U38849 (N_38849,N_37266,N_37363);
xnor U38850 (N_38850,N_37094,N_37236);
xor U38851 (N_38851,N_37610,N_37716);
nand U38852 (N_38852,N_37008,N_37545);
nand U38853 (N_38853,N_37125,N_37251);
nor U38854 (N_38854,N_37165,N_37753);
or U38855 (N_38855,N_37841,N_37695);
and U38856 (N_38856,N_37371,N_37750);
xor U38857 (N_38857,N_37492,N_37595);
or U38858 (N_38858,N_37020,N_37140);
or U38859 (N_38859,N_37801,N_37377);
or U38860 (N_38860,N_37042,N_37359);
or U38861 (N_38861,N_37500,N_37002);
nand U38862 (N_38862,N_37253,N_37487);
and U38863 (N_38863,N_37917,N_37181);
or U38864 (N_38864,N_37494,N_37360);
or U38865 (N_38865,N_37910,N_37908);
nor U38866 (N_38866,N_37903,N_37280);
nor U38867 (N_38867,N_37420,N_37451);
xor U38868 (N_38868,N_37488,N_37919);
and U38869 (N_38869,N_37130,N_37504);
nand U38870 (N_38870,N_37445,N_37758);
or U38871 (N_38871,N_37808,N_37936);
or U38872 (N_38872,N_37132,N_37270);
nand U38873 (N_38873,N_37318,N_37937);
xor U38874 (N_38874,N_37924,N_37514);
nand U38875 (N_38875,N_37332,N_37395);
nor U38876 (N_38876,N_37472,N_37921);
nand U38877 (N_38877,N_37818,N_37479);
or U38878 (N_38878,N_37173,N_37031);
xor U38879 (N_38879,N_37494,N_37217);
or U38880 (N_38880,N_37259,N_37437);
and U38881 (N_38881,N_37825,N_37023);
xor U38882 (N_38882,N_37551,N_37209);
or U38883 (N_38883,N_37142,N_37394);
xor U38884 (N_38884,N_37724,N_37891);
or U38885 (N_38885,N_37947,N_37377);
xor U38886 (N_38886,N_37725,N_37970);
and U38887 (N_38887,N_37585,N_37649);
xnor U38888 (N_38888,N_37245,N_37937);
and U38889 (N_38889,N_37120,N_37587);
and U38890 (N_38890,N_37448,N_37885);
nor U38891 (N_38891,N_37618,N_37793);
or U38892 (N_38892,N_37528,N_37362);
nor U38893 (N_38893,N_37221,N_37828);
nand U38894 (N_38894,N_37072,N_37103);
xnor U38895 (N_38895,N_37206,N_37149);
and U38896 (N_38896,N_37389,N_37540);
or U38897 (N_38897,N_37974,N_37837);
nand U38898 (N_38898,N_37200,N_37918);
and U38899 (N_38899,N_37189,N_37778);
nor U38900 (N_38900,N_37790,N_37690);
xnor U38901 (N_38901,N_37868,N_37583);
xor U38902 (N_38902,N_37930,N_37646);
and U38903 (N_38903,N_37817,N_37830);
nand U38904 (N_38904,N_37279,N_37581);
and U38905 (N_38905,N_37570,N_37755);
or U38906 (N_38906,N_37757,N_37469);
nor U38907 (N_38907,N_37413,N_37659);
nand U38908 (N_38908,N_37749,N_37981);
nand U38909 (N_38909,N_37518,N_37705);
xor U38910 (N_38910,N_37438,N_37884);
nor U38911 (N_38911,N_37403,N_37198);
and U38912 (N_38912,N_37044,N_37537);
nor U38913 (N_38913,N_37664,N_37471);
nand U38914 (N_38914,N_37592,N_37501);
or U38915 (N_38915,N_37269,N_37888);
xnor U38916 (N_38916,N_37420,N_37770);
nand U38917 (N_38917,N_37955,N_37610);
or U38918 (N_38918,N_37184,N_37749);
and U38919 (N_38919,N_37983,N_37090);
nand U38920 (N_38920,N_37268,N_37036);
xnor U38921 (N_38921,N_37100,N_37753);
and U38922 (N_38922,N_37825,N_37539);
nor U38923 (N_38923,N_37346,N_37412);
and U38924 (N_38924,N_37983,N_37418);
and U38925 (N_38925,N_37882,N_37344);
nor U38926 (N_38926,N_37371,N_37253);
and U38927 (N_38927,N_37818,N_37482);
nor U38928 (N_38928,N_37488,N_37030);
nand U38929 (N_38929,N_37528,N_37737);
nand U38930 (N_38930,N_37894,N_37892);
or U38931 (N_38931,N_37423,N_37772);
xnor U38932 (N_38932,N_37360,N_37971);
or U38933 (N_38933,N_37000,N_37714);
and U38934 (N_38934,N_37882,N_37347);
xor U38935 (N_38935,N_37707,N_37350);
and U38936 (N_38936,N_37529,N_37735);
xor U38937 (N_38937,N_37436,N_37283);
and U38938 (N_38938,N_37524,N_37855);
xnor U38939 (N_38939,N_37579,N_37067);
xnor U38940 (N_38940,N_37567,N_37423);
xnor U38941 (N_38941,N_37270,N_37470);
nor U38942 (N_38942,N_37682,N_37635);
nor U38943 (N_38943,N_37015,N_37397);
nor U38944 (N_38944,N_37320,N_37937);
nor U38945 (N_38945,N_37321,N_37754);
xnor U38946 (N_38946,N_37023,N_37499);
and U38947 (N_38947,N_37758,N_37304);
and U38948 (N_38948,N_37523,N_37952);
nor U38949 (N_38949,N_37834,N_37874);
xnor U38950 (N_38950,N_37640,N_37120);
nand U38951 (N_38951,N_37207,N_37697);
nor U38952 (N_38952,N_37584,N_37687);
or U38953 (N_38953,N_37215,N_37602);
xor U38954 (N_38954,N_37579,N_37511);
or U38955 (N_38955,N_37163,N_37338);
xnor U38956 (N_38956,N_37148,N_37240);
or U38957 (N_38957,N_37525,N_37431);
or U38958 (N_38958,N_37620,N_37068);
and U38959 (N_38959,N_37096,N_37668);
or U38960 (N_38960,N_37443,N_37971);
nor U38961 (N_38961,N_37668,N_37477);
and U38962 (N_38962,N_37980,N_37776);
nor U38963 (N_38963,N_37026,N_37011);
nand U38964 (N_38964,N_37320,N_37151);
or U38965 (N_38965,N_37961,N_37030);
xor U38966 (N_38966,N_37773,N_37819);
nand U38967 (N_38967,N_37515,N_37247);
and U38968 (N_38968,N_37746,N_37829);
nand U38969 (N_38969,N_37209,N_37858);
nand U38970 (N_38970,N_37635,N_37575);
nand U38971 (N_38971,N_37785,N_37744);
or U38972 (N_38972,N_37215,N_37760);
and U38973 (N_38973,N_37026,N_37765);
or U38974 (N_38974,N_37574,N_37210);
or U38975 (N_38975,N_37550,N_37159);
xnor U38976 (N_38976,N_37688,N_37340);
xnor U38977 (N_38977,N_37686,N_37907);
nand U38978 (N_38978,N_37913,N_37053);
nand U38979 (N_38979,N_37420,N_37986);
and U38980 (N_38980,N_37398,N_37435);
and U38981 (N_38981,N_37380,N_37584);
or U38982 (N_38982,N_37956,N_37066);
and U38983 (N_38983,N_37696,N_37501);
or U38984 (N_38984,N_37688,N_37760);
nor U38985 (N_38985,N_37456,N_37346);
or U38986 (N_38986,N_37789,N_37805);
nor U38987 (N_38987,N_37603,N_37640);
and U38988 (N_38988,N_37963,N_37113);
nor U38989 (N_38989,N_37066,N_37228);
xnor U38990 (N_38990,N_37458,N_37345);
nor U38991 (N_38991,N_37887,N_37896);
xor U38992 (N_38992,N_37639,N_37050);
nand U38993 (N_38993,N_37765,N_37180);
and U38994 (N_38994,N_37355,N_37654);
xor U38995 (N_38995,N_37521,N_37455);
xor U38996 (N_38996,N_37037,N_37203);
nor U38997 (N_38997,N_37956,N_37910);
and U38998 (N_38998,N_37894,N_37149);
nand U38999 (N_38999,N_37249,N_37430);
nor U39000 (N_39000,N_38526,N_38455);
nand U39001 (N_39001,N_38897,N_38084);
nor U39002 (N_39002,N_38178,N_38549);
nor U39003 (N_39003,N_38152,N_38399);
or U39004 (N_39004,N_38354,N_38102);
nor U39005 (N_39005,N_38690,N_38693);
nand U39006 (N_39006,N_38508,N_38781);
or U39007 (N_39007,N_38763,N_38658);
nor U39008 (N_39008,N_38067,N_38884);
and U39009 (N_39009,N_38050,N_38255);
xnor U39010 (N_39010,N_38671,N_38792);
nor U39011 (N_39011,N_38689,N_38414);
nor U39012 (N_39012,N_38183,N_38976);
xnor U39013 (N_39013,N_38499,N_38972);
nor U39014 (N_39014,N_38638,N_38448);
and U39015 (N_39015,N_38008,N_38584);
or U39016 (N_39016,N_38556,N_38462);
and U39017 (N_39017,N_38900,N_38062);
xnor U39018 (N_39018,N_38465,N_38843);
and U39019 (N_39019,N_38127,N_38100);
xor U39020 (N_39020,N_38487,N_38058);
nand U39021 (N_39021,N_38513,N_38053);
and U39022 (N_39022,N_38672,N_38806);
and U39023 (N_39023,N_38336,N_38847);
and U39024 (N_39024,N_38394,N_38951);
xor U39025 (N_39025,N_38665,N_38735);
and U39026 (N_39026,N_38572,N_38799);
or U39027 (N_39027,N_38630,N_38582);
and U39028 (N_39028,N_38994,N_38683);
nand U39029 (N_39029,N_38870,N_38154);
or U39030 (N_39030,N_38567,N_38576);
and U39031 (N_39031,N_38509,N_38515);
nor U39032 (N_39032,N_38995,N_38385);
or U39033 (N_39033,N_38550,N_38812);
xnor U39034 (N_39034,N_38844,N_38351);
nor U39035 (N_39035,N_38371,N_38089);
or U39036 (N_39036,N_38198,N_38396);
and U39037 (N_39037,N_38500,N_38603);
and U39038 (N_39038,N_38293,N_38025);
nor U39039 (N_39039,N_38544,N_38705);
nor U39040 (N_39040,N_38675,N_38450);
and U39041 (N_39041,N_38047,N_38287);
xor U39042 (N_39042,N_38337,N_38179);
and U39043 (N_39043,N_38194,N_38766);
nor U39044 (N_39044,N_38098,N_38290);
xnor U39045 (N_39045,N_38350,N_38708);
or U39046 (N_39046,N_38483,N_38642);
and U39047 (N_39047,N_38563,N_38277);
nand U39048 (N_39048,N_38626,N_38349);
or U39049 (N_39049,N_38447,N_38876);
xnor U39050 (N_39050,N_38629,N_38326);
nor U39051 (N_39051,N_38566,N_38568);
nor U39052 (N_39052,N_38967,N_38221);
nand U39053 (N_39053,N_38332,N_38871);
nand U39054 (N_39054,N_38219,N_38112);
or U39055 (N_39055,N_38554,N_38898);
nand U39056 (N_39056,N_38969,N_38203);
and U39057 (N_39057,N_38159,N_38535);
or U39058 (N_39058,N_38774,N_38470);
nor U39059 (N_39059,N_38364,N_38751);
or U39060 (N_39060,N_38537,N_38374);
xor U39061 (N_39061,N_38056,N_38055);
and U39062 (N_39062,N_38760,N_38457);
and U39063 (N_39063,N_38920,N_38824);
or U39064 (N_39064,N_38390,N_38041);
nand U39065 (N_39065,N_38264,N_38475);
xor U39066 (N_39066,N_38674,N_38692);
and U39067 (N_39067,N_38542,N_38239);
and U39068 (N_39068,N_38808,N_38668);
xor U39069 (N_39069,N_38966,N_38765);
nand U39070 (N_39070,N_38829,N_38123);
and U39071 (N_39071,N_38181,N_38408);
nor U39072 (N_39072,N_38868,N_38482);
or U39073 (N_39073,N_38771,N_38149);
nand U39074 (N_39074,N_38185,N_38963);
nand U39075 (N_39075,N_38652,N_38360);
xnor U39076 (N_39076,N_38398,N_38661);
nor U39077 (N_39077,N_38384,N_38120);
or U39078 (N_39078,N_38459,N_38511);
or U39079 (N_39079,N_38153,N_38432);
nor U39080 (N_39080,N_38930,N_38233);
nand U39081 (N_39081,N_38212,N_38273);
nand U39082 (N_39082,N_38788,N_38895);
nor U39083 (N_39083,N_38190,N_38862);
or U39084 (N_39084,N_38078,N_38468);
and U39085 (N_39085,N_38421,N_38249);
nand U39086 (N_39086,N_38987,N_38232);
xor U39087 (N_39087,N_38850,N_38315);
nor U39088 (N_39088,N_38655,N_38863);
or U39089 (N_39089,N_38320,N_38775);
nor U39090 (N_39090,N_38131,N_38379);
nand U39091 (N_39091,N_38932,N_38184);
nand U39092 (N_39092,N_38243,N_38126);
xnor U39093 (N_39093,N_38309,N_38659);
and U39094 (N_39094,N_38444,N_38971);
nor U39095 (N_39095,N_38677,N_38024);
nand U39096 (N_39096,N_38237,N_38023);
and U39097 (N_39097,N_38175,N_38193);
or U39098 (N_39098,N_38727,N_38296);
nand U39099 (N_39099,N_38247,N_38540);
xnor U39100 (N_39100,N_38367,N_38722);
and U39101 (N_39101,N_38478,N_38993);
or U39102 (N_39102,N_38142,N_38104);
nand U39103 (N_39103,N_38518,N_38060);
or U39104 (N_39104,N_38541,N_38637);
xor U39105 (N_39105,N_38803,N_38528);
nor U39106 (N_39106,N_38724,N_38947);
xor U39107 (N_39107,N_38064,N_38430);
or U39108 (N_39108,N_38553,N_38136);
and U39109 (N_39109,N_38736,N_38866);
or U39110 (N_39110,N_38321,N_38125);
nor U39111 (N_39111,N_38887,N_38650);
xor U39112 (N_39112,N_38789,N_38191);
and U39113 (N_39113,N_38785,N_38881);
or U39114 (N_39114,N_38501,N_38497);
xor U39115 (N_39115,N_38324,N_38076);
nand U39116 (N_39116,N_38767,N_38837);
or U39117 (N_39117,N_38376,N_38820);
nand U39118 (N_39118,N_38954,N_38935);
and U39119 (N_39119,N_38040,N_38725);
or U39120 (N_39120,N_38507,N_38469);
and U39121 (N_39121,N_38546,N_38797);
and U39122 (N_39122,N_38706,N_38271);
nand U39123 (N_39123,N_38464,N_38691);
or U39124 (N_39124,N_38467,N_38983);
nor U39125 (N_39125,N_38019,N_38519);
nand U39126 (N_39126,N_38344,N_38316);
or U39127 (N_39127,N_38503,N_38739);
nor U39128 (N_39128,N_38527,N_38558);
xor U39129 (N_39129,N_38333,N_38359);
nor U39130 (N_39130,N_38317,N_38624);
or U39131 (N_39131,N_38617,N_38434);
xnor U39132 (N_39132,N_38529,N_38807);
nor U39133 (N_39133,N_38522,N_38890);
xnor U39134 (N_39134,N_38569,N_38817);
or U39135 (N_39135,N_38037,N_38363);
and U39136 (N_39136,N_38801,N_38295);
xor U39137 (N_39137,N_38140,N_38960);
xor U39138 (N_39138,N_38228,N_38646);
nor U39139 (N_39139,N_38709,N_38439);
and U39140 (N_39140,N_38564,N_38283);
and U39141 (N_39141,N_38621,N_38533);
xnor U39142 (N_39142,N_38428,N_38169);
nor U39143 (N_39143,N_38805,N_38044);
and U39144 (N_39144,N_38956,N_38926);
and U39145 (N_39145,N_38049,N_38220);
nand U39146 (N_39146,N_38780,N_38783);
xor U39147 (N_39147,N_38749,N_38458);
xor U39148 (N_39148,N_38451,N_38137);
and U39149 (N_39149,N_38498,N_38919);
nor U39150 (N_39150,N_38991,N_38816);
and U39151 (N_39151,N_38252,N_38051);
nor U39152 (N_39152,N_38073,N_38505);
or U39153 (N_39153,N_38813,N_38453);
or U39154 (N_39154,N_38688,N_38707);
or U39155 (N_39155,N_38686,N_38347);
nor U39156 (N_39156,N_38280,N_38885);
xnor U39157 (N_39157,N_38429,N_38555);
xor U39158 (N_39158,N_38882,N_38004);
nand U39159 (N_39159,N_38879,N_38952);
and U39160 (N_39160,N_38633,N_38562);
xor U39161 (N_39161,N_38086,N_38597);
nand U39162 (N_39162,N_38209,N_38996);
nand U39163 (N_39163,N_38440,N_38188);
nor U39164 (N_39164,N_38640,N_38955);
nand U39165 (N_39165,N_38859,N_38662);
or U39166 (N_39166,N_38445,N_38894);
xor U39167 (N_39167,N_38113,N_38669);
xnor U39168 (N_39168,N_38180,N_38224);
nor U39169 (N_39169,N_38581,N_38045);
xor U39170 (N_39170,N_38605,N_38281);
or U39171 (N_39171,N_38115,N_38609);
nand U39172 (N_39172,N_38305,N_38773);
or U39173 (N_39173,N_38480,N_38857);
nand U39174 (N_39174,N_38422,N_38405);
or U39175 (N_39175,N_38907,N_38227);
nand U39176 (N_39176,N_38201,N_38922);
xor U39177 (N_39177,N_38016,N_38088);
nand U39178 (N_39178,N_38973,N_38740);
xor U39179 (N_39179,N_38075,N_38033);
nor U39180 (N_39180,N_38338,N_38176);
nand U39181 (N_39181,N_38380,N_38716);
and U39182 (N_39182,N_38443,N_38278);
and U39183 (N_39183,N_38061,N_38510);
and U39184 (N_39184,N_38560,N_38391);
nor U39185 (N_39185,N_38006,N_38081);
or U39186 (N_39186,N_38072,N_38578);
nand U39187 (N_39187,N_38306,N_38348);
or U39188 (N_39188,N_38990,N_38046);
nand U39189 (N_39189,N_38158,N_38903);
xor U39190 (N_39190,N_38916,N_38502);
nand U39191 (N_39191,N_38002,N_38710);
nor U39192 (N_39192,N_38342,N_38835);
and U39193 (N_39193,N_38759,N_38551);
xor U39194 (N_39194,N_38752,N_38413);
xnor U39195 (N_39195,N_38595,N_38156);
nand U39196 (N_39196,N_38580,N_38171);
nand U39197 (N_39197,N_38941,N_38848);
or U39198 (N_39198,N_38623,N_38130);
xor U39199 (N_39199,N_38001,N_38852);
or U39200 (N_39200,N_38250,N_38009);
xnor U39201 (N_39201,N_38715,N_38608);
xor U39202 (N_39202,N_38214,N_38998);
and U39203 (N_39203,N_38275,N_38823);
xor U39204 (N_39204,N_38388,N_38641);
xor U39205 (N_39205,N_38625,N_38654);
and U39206 (N_39206,N_38984,N_38636);
or U39207 (N_39207,N_38488,N_38657);
nor U39208 (N_39208,N_38695,N_38777);
nand U39209 (N_39209,N_38694,N_38880);
or U39210 (N_39210,N_38986,N_38815);
or U39211 (N_39211,N_38303,N_38111);
or U39212 (N_39212,N_38036,N_38420);
xor U39213 (N_39213,N_38666,N_38099);
nand U39214 (N_39214,N_38682,N_38375);
or U39215 (N_39215,N_38905,N_38068);
xnor U39216 (N_39216,N_38479,N_38818);
or U39217 (N_39217,N_38370,N_38855);
nand U39218 (N_39218,N_38892,N_38741);
xnor U39219 (N_39219,N_38854,N_38588);
xnor U39220 (N_39220,N_38723,N_38417);
or U39221 (N_39221,N_38079,N_38520);
nand U39222 (N_39222,N_38486,N_38622);
and U39223 (N_39223,N_38474,N_38726);
and U39224 (N_39224,N_38248,N_38970);
nand U39225 (N_39225,N_38231,N_38992);
xnor U39226 (N_39226,N_38254,N_38330);
or U39227 (N_39227,N_38311,N_38210);
nor U39228 (N_39228,N_38085,N_38819);
or U39229 (N_39229,N_38861,N_38128);
nand U39230 (N_39230,N_38092,N_38928);
xor U39231 (N_39231,N_38411,N_38257);
nand U39232 (N_39232,N_38017,N_38943);
nor U39233 (N_39233,N_38034,N_38620);
or U39234 (N_39234,N_38978,N_38719);
and U39235 (N_39235,N_38856,N_38825);
or U39236 (N_39236,N_38832,N_38714);
nor U39237 (N_39237,N_38341,N_38531);
nand U39238 (N_39238,N_38968,N_38794);
xor U39239 (N_39239,N_38313,N_38762);
nor U39240 (N_39240,N_38069,N_38291);
and U39241 (N_39241,N_38242,N_38942);
nor U39242 (N_39242,N_38246,N_38407);
nand U39243 (N_39243,N_38573,N_38548);
nor U39244 (N_39244,N_38702,N_38925);
nor U39245 (N_39245,N_38010,N_38048);
nor U39246 (N_39246,N_38750,N_38754);
xnor U39247 (N_39247,N_38744,N_38020);
nor U39248 (N_39248,N_38961,N_38018);
nor U39249 (N_39249,N_38787,N_38218);
xor U39250 (N_39250,N_38628,N_38891);
nand U39251 (N_39251,N_38981,N_38308);
xnor U39252 (N_39252,N_38322,N_38168);
or U39253 (N_39253,N_38160,N_38600);
nand U39254 (N_39254,N_38071,N_38786);
nor U39255 (N_39255,N_38521,N_38899);
or U39256 (N_39256,N_38733,N_38192);
or U39257 (N_39257,N_38229,N_38957);
nand U39258 (N_39258,N_38696,N_38294);
and U39259 (N_39259,N_38846,N_38979);
and U39260 (N_39260,N_38356,N_38433);
nor U39261 (N_39261,N_38082,N_38331);
nand U39262 (N_39262,N_38343,N_38836);
nand U39263 (N_39263,N_38094,N_38800);
nor U39264 (N_39264,N_38416,N_38393);
or U39265 (N_39265,N_38756,N_38005);
and U39266 (N_39266,N_38423,N_38265);
nand U39267 (N_39267,N_38205,N_38953);
and U39268 (N_39268,N_38743,N_38174);
or U39269 (N_39269,N_38138,N_38599);
xor U39270 (N_39270,N_38012,N_38875);
and U39271 (N_39271,N_38485,N_38980);
xnor U39272 (N_39272,N_38031,N_38093);
xnor U39273 (N_39273,N_38685,N_38262);
and U39274 (N_39274,N_38673,N_38424);
and U39275 (N_39275,N_38177,N_38559);
xnor U39276 (N_39276,N_38245,N_38105);
nand U39277 (N_39277,N_38286,N_38170);
nor U39278 (N_39278,N_38831,N_38684);
nand U39279 (N_39279,N_38858,N_38878);
or U39280 (N_39280,N_38616,N_38590);
nor U39281 (N_39281,N_38680,N_38028);
nand U39282 (N_39282,N_38108,N_38297);
xnor U39283 (N_39283,N_38292,N_38867);
nor U39284 (N_39284,N_38225,N_38575);
nand U39285 (N_39285,N_38030,N_38090);
nor U39286 (N_39286,N_38631,N_38997);
or U39287 (N_39287,N_38366,N_38999);
and U39288 (N_39288,N_38914,N_38604);
and U39289 (N_39289,N_38213,N_38974);
xor U39290 (N_39290,N_38977,N_38570);
nand U39291 (N_39291,N_38770,N_38793);
xor U39292 (N_39292,N_38589,N_38938);
xor U39293 (N_39293,N_38606,N_38934);
nand U39294 (N_39294,N_38378,N_38387);
xor U39295 (N_39295,N_38811,N_38196);
nand U39296 (N_39296,N_38769,N_38267);
and U39297 (N_39297,N_38096,N_38494);
and U39298 (N_39298,N_38784,N_38352);
nor U39299 (N_39299,N_38840,N_38944);
xnor U39300 (N_39300,N_38199,N_38426);
nor U39301 (N_39301,N_38027,N_38216);
xor U39302 (N_39302,N_38207,N_38670);
and U39303 (N_39303,N_38757,N_38755);
nand U39304 (N_39304,N_38516,N_38314);
or U39305 (N_39305,N_38738,N_38574);
and U39306 (N_39306,N_38687,N_38274);
nand U39307 (N_39307,N_38372,N_38368);
or U39308 (N_39308,N_38425,N_38013);
nor U39309 (N_39309,N_38427,N_38155);
and U39310 (N_39310,N_38651,N_38074);
nand U39311 (N_39311,N_38101,N_38007);
xnor U39312 (N_39312,N_38150,N_38300);
nand U39313 (N_39313,N_38596,N_38664);
and U39314 (N_39314,N_38889,N_38463);
nand U39315 (N_39315,N_38054,N_38403);
or U39316 (N_39316,N_38373,N_38461);
xor U39317 (N_39317,N_38235,N_38717);
and U39318 (N_39318,N_38442,N_38946);
nor U39319 (N_39319,N_38285,N_38933);
nor U39320 (N_39320,N_38864,N_38746);
nor U39321 (N_39321,N_38116,N_38798);
xnor U39322 (N_39322,N_38383,N_38489);
xnor U39323 (N_39323,N_38147,N_38206);
nor U39324 (N_39324,N_38734,N_38748);
and U39325 (N_39325,N_38340,N_38985);
or U39326 (N_39326,N_38594,N_38400);
or U39327 (N_39327,N_38392,N_38256);
nand U39328 (N_39328,N_38222,N_38110);
or U39329 (N_39329,N_38240,N_38253);
xnor U39330 (N_39330,N_38648,N_38307);
or U39331 (N_39331,N_38369,N_38276);
xor U39332 (N_39332,N_38197,N_38679);
nor U39333 (N_39333,N_38678,N_38146);
or U39334 (N_39334,N_38833,N_38395);
xor U39335 (N_39335,N_38318,N_38796);
xnor U39336 (N_39336,N_38477,N_38122);
nand U39337 (N_39337,N_38779,N_38543);
or U39338 (N_39338,N_38167,N_38057);
nand U39339 (N_39339,N_38524,N_38676);
nand U39340 (N_39340,N_38720,N_38959);
nand U39341 (N_39341,N_38145,N_38901);
or U39342 (N_39342,N_38304,N_38329);
nor U39343 (N_39343,N_38830,N_38269);
xor U39344 (N_39344,N_38063,N_38157);
nor U39345 (N_39345,N_38139,N_38545);
or U39346 (N_39346,N_38711,N_38591);
xnor U39347 (N_39347,N_38382,N_38189);
nor U39348 (N_39348,N_38215,N_38328);
nor U39349 (N_39349,N_38441,N_38557);
and U39350 (N_39350,N_38910,N_38512);
or U39351 (N_39351,N_38263,N_38842);
nand U39352 (N_39352,N_38618,N_38607);
or U39353 (N_39353,N_38401,N_38107);
and U39354 (N_39354,N_38965,N_38134);
and U39355 (N_39355,N_38187,N_38106);
nor U39356 (N_39356,N_38026,N_38299);
xor U39357 (N_39357,N_38270,N_38460);
or U39358 (N_39358,N_38547,N_38161);
and U39359 (N_39359,N_38230,N_38718);
or U39360 (N_39360,N_38782,N_38473);
xor U39361 (N_39361,N_38525,N_38163);
nand U39362 (N_39362,N_38656,N_38731);
and U39363 (N_39363,N_38135,N_38583);
xor U39364 (N_39364,N_38619,N_38284);
or U39365 (N_39365,N_38663,N_38172);
nand U39366 (N_39366,N_38173,N_38251);
xor U39367 (N_39367,N_38810,N_38059);
nand U39368 (N_39368,N_38319,N_38491);
and U39369 (N_39369,N_38964,N_38923);
nand U39370 (N_39370,N_38517,N_38386);
xor U39371 (N_39371,N_38109,N_38912);
or U39372 (N_39372,N_38182,N_38538);
or U39373 (N_39373,N_38828,N_38896);
nor U39374 (N_39374,N_38790,N_38827);
nor U39375 (N_39375,N_38698,N_38975);
or U39376 (N_39376,N_38087,N_38355);
nand U39377 (N_39377,N_38377,N_38419);
xor U39378 (N_39378,N_38409,N_38472);
xor U39379 (N_39379,N_38449,N_38593);
nor U39380 (N_39380,N_38365,N_38402);
nand U39381 (N_39381,N_38639,N_38795);
or U39382 (N_39382,N_38579,N_38851);
and U39383 (N_39383,N_38883,N_38029);
xnor U39384 (N_39384,N_38758,N_38335);
or U39385 (N_39385,N_38841,N_38612);
or U39386 (N_39386,N_38406,N_38200);
xor U39387 (N_39387,N_38611,N_38141);
nor U39388 (N_39388,N_38021,N_38412);
or U39389 (N_39389,N_38118,N_38471);
nor U39390 (N_39390,N_38312,N_38431);
nor U39391 (N_39391,N_38834,N_38032);
and U39392 (N_39392,N_38989,N_38948);
or U39393 (N_39393,N_38768,N_38083);
and U39394 (N_39394,N_38091,N_38721);
and U39395 (N_39395,N_38838,N_38404);
nand U39396 (N_39396,N_38778,N_38162);
nor U39397 (N_39397,N_38747,N_38732);
or U39398 (N_39398,N_38602,N_38346);
nand U39399 (N_39399,N_38070,N_38492);
nand U39400 (N_39400,N_38598,N_38035);
xor U39401 (N_39401,N_38610,N_38266);
nor U39402 (N_39402,N_38982,N_38904);
nand U39403 (N_39403,N_38217,N_38011);
nor U39404 (N_39404,N_38845,N_38298);
nand U39405 (N_39405,N_38592,N_38647);
xor U39406 (N_39406,N_38909,N_38586);
xnor U39407 (N_39407,N_38334,N_38282);
and U39408 (N_39408,N_38065,N_38117);
xnor U39409 (N_39409,N_38565,N_38761);
nand U39410 (N_39410,N_38700,N_38886);
nand U39411 (N_39411,N_38211,N_38042);
nor U39412 (N_39412,N_38534,N_38446);
or U39413 (N_39413,N_38361,N_38523);
nor U39414 (N_39414,N_38821,N_38077);
or U39415 (N_39415,N_38186,N_38849);
nor U39416 (N_39416,N_38643,N_38259);
and U39417 (N_39417,N_38301,N_38915);
or U39418 (N_39418,N_38802,N_38962);
xor U39419 (N_39419,N_38103,N_38772);
xnor U39420 (N_39420,N_38660,N_38279);
xor U39421 (N_39421,N_38166,N_38052);
or U39422 (N_39422,N_38873,N_38124);
or U39423 (N_39423,N_38937,N_38202);
nand U39424 (N_39424,N_38362,N_38456);
nor U39425 (N_39425,N_38737,N_38791);
xnor U39426 (N_39426,N_38949,N_38437);
or U39427 (N_39427,N_38729,N_38940);
and U39428 (N_39428,N_38151,N_38888);
nor U39429 (N_39429,N_38614,N_38234);
nand U39430 (N_39430,N_38310,N_38260);
nor U39431 (N_39431,N_38902,N_38132);
nand U39432 (N_39432,N_38701,N_38635);
xor U39433 (N_39433,N_38950,N_38381);
and U39434 (N_39434,N_38435,N_38601);
nand U39435 (N_39435,N_38921,N_38357);
or U39436 (N_39436,N_38822,N_38632);
nor U39437 (N_39437,N_38730,N_38418);
nand U39438 (N_39438,N_38804,N_38667);
nand U39439 (N_39439,N_38204,N_38927);
and U39440 (N_39440,N_38587,N_38415);
and U39441 (N_39441,N_38917,N_38258);
and U39442 (N_39442,N_38003,N_38645);
nand U39443 (N_39443,N_38860,N_38649);
xor U39444 (N_39444,N_38764,N_38014);
nor U39445 (N_39445,N_38712,N_38874);
nor U39446 (N_39446,N_38918,N_38809);
xnor U39447 (N_39447,N_38114,N_38261);
nor U39448 (N_39448,N_38452,N_38238);
or U39449 (N_39449,N_38148,N_38530);
nand U39450 (N_39450,N_38877,N_38038);
nor U39451 (N_39451,N_38345,N_38585);
and U39452 (N_39452,N_38484,N_38713);
xor U39453 (N_39453,N_38389,N_38121);
xor U39454 (N_39454,N_38097,N_38129);
nor U39455 (N_39455,N_38839,N_38438);
or U39456 (N_39456,N_38244,N_38144);
nor U39457 (N_39457,N_38945,N_38353);
or U39458 (N_39458,N_38043,N_38703);
nor U39459 (N_39459,N_38325,N_38165);
nand U39460 (N_39460,N_38911,N_38358);
or U39461 (N_39461,N_38697,N_38095);
xor U39462 (N_39462,N_38865,N_38699);
nand U39463 (N_39463,N_38704,N_38133);
nor U39464 (N_39464,N_38561,N_38924);
xnor U39465 (N_39465,N_38195,N_38577);
nor U39466 (N_39466,N_38143,N_38022);
xnor U39467 (N_39467,N_38644,N_38000);
nand U39468 (N_39468,N_38634,N_38536);
or U39469 (N_39469,N_38853,N_38514);
nand U39470 (N_39470,N_38241,N_38268);
nand U39471 (N_39471,N_38613,N_38504);
nand U39472 (N_39472,N_38066,N_38681);
nor U39473 (N_39473,N_38039,N_38236);
nand U39474 (N_39474,N_38931,N_38490);
or U39475 (N_39475,N_38627,N_38552);
nor U39476 (N_39476,N_38288,N_38302);
nor U39477 (N_39477,N_38476,N_38936);
or U39478 (N_39478,N_38742,N_38939);
nor U39479 (N_39479,N_38080,N_38776);
nor U39480 (N_39480,N_38015,N_38869);
or U39481 (N_39481,N_38119,N_38481);
nor U39482 (N_39482,N_38496,N_38745);
or U39483 (N_39483,N_38223,N_38493);
xor U39484 (N_39484,N_38653,N_38327);
nand U39485 (N_39485,N_38615,N_38908);
and U39486 (N_39486,N_38929,N_38466);
and U39487 (N_39487,N_38506,N_38289);
and U39488 (N_39488,N_38913,N_38495);
nand U39489 (N_39489,N_38539,N_38272);
nand U39490 (N_39490,N_38397,N_38208);
nand U39491 (N_39491,N_38339,N_38436);
xnor U39492 (N_39492,N_38893,N_38958);
nor U39493 (N_39493,N_38323,N_38226);
or U39494 (N_39494,N_38410,N_38826);
xor U39495 (N_39495,N_38571,N_38454);
and U39496 (N_39496,N_38814,N_38532);
or U39497 (N_39497,N_38164,N_38872);
nand U39498 (N_39498,N_38906,N_38728);
xnor U39499 (N_39499,N_38988,N_38753);
nand U39500 (N_39500,N_38952,N_38592);
or U39501 (N_39501,N_38786,N_38764);
or U39502 (N_39502,N_38940,N_38046);
and U39503 (N_39503,N_38267,N_38394);
xnor U39504 (N_39504,N_38259,N_38470);
and U39505 (N_39505,N_38702,N_38095);
nor U39506 (N_39506,N_38341,N_38106);
xnor U39507 (N_39507,N_38343,N_38766);
nand U39508 (N_39508,N_38136,N_38681);
nor U39509 (N_39509,N_38303,N_38908);
nor U39510 (N_39510,N_38375,N_38628);
or U39511 (N_39511,N_38625,N_38803);
xnor U39512 (N_39512,N_38136,N_38888);
nor U39513 (N_39513,N_38842,N_38720);
nor U39514 (N_39514,N_38017,N_38406);
or U39515 (N_39515,N_38566,N_38868);
and U39516 (N_39516,N_38899,N_38283);
xor U39517 (N_39517,N_38963,N_38494);
nand U39518 (N_39518,N_38582,N_38626);
and U39519 (N_39519,N_38913,N_38665);
or U39520 (N_39520,N_38293,N_38357);
and U39521 (N_39521,N_38832,N_38221);
xnor U39522 (N_39522,N_38589,N_38088);
xnor U39523 (N_39523,N_38582,N_38510);
or U39524 (N_39524,N_38932,N_38660);
xnor U39525 (N_39525,N_38585,N_38716);
and U39526 (N_39526,N_38013,N_38932);
nor U39527 (N_39527,N_38948,N_38760);
xor U39528 (N_39528,N_38330,N_38118);
nand U39529 (N_39529,N_38211,N_38670);
and U39530 (N_39530,N_38734,N_38238);
or U39531 (N_39531,N_38993,N_38248);
nor U39532 (N_39532,N_38406,N_38107);
or U39533 (N_39533,N_38659,N_38415);
and U39534 (N_39534,N_38357,N_38171);
nor U39535 (N_39535,N_38893,N_38444);
nand U39536 (N_39536,N_38740,N_38719);
nor U39537 (N_39537,N_38816,N_38829);
nor U39538 (N_39538,N_38506,N_38184);
nor U39539 (N_39539,N_38461,N_38014);
nand U39540 (N_39540,N_38075,N_38486);
xor U39541 (N_39541,N_38459,N_38011);
or U39542 (N_39542,N_38521,N_38210);
nand U39543 (N_39543,N_38708,N_38249);
nand U39544 (N_39544,N_38186,N_38188);
xor U39545 (N_39545,N_38718,N_38832);
xnor U39546 (N_39546,N_38495,N_38308);
nand U39547 (N_39547,N_38083,N_38846);
nand U39548 (N_39548,N_38590,N_38015);
and U39549 (N_39549,N_38799,N_38774);
and U39550 (N_39550,N_38883,N_38257);
nand U39551 (N_39551,N_38745,N_38654);
nand U39552 (N_39552,N_38052,N_38382);
xnor U39553 (N_39553,N_38045,N_38833);
xor U39554 (N_39554,N_38110,N_38124);
nand U39555 (N_39555,N_38796,N_38439);
xor U39556 (N_39556,N_38792,N_38143);
xor U39557 (N_39557,N_38164,N_38525);
xor U39558 (N_39558,N_38689,N_38234);
nand U39559 (N_39559,N_38948,N_38581);
or U39560 (N_39560,N_38528,N_38810);
and U39561 (N_39561,N_38350,N_38842);
nand U39562 (N_39562,N_38021,N_38534);
xor U39563 (N_39563,N_38477,N_38181);
or U39564 (N_39564,N_38098,N_38465);
or U39565 (N_39565,N_38422,N_38166);
xnor U39566 (N_39566,N_38608,N_38132);
or U39567 (N_39567,N_38476,N_38062);
nand U39568 (N_39568,N_38698,N_38842);
nor U39569 (N_39569,N_38292,N_38398);
nor U39570 (N_39570,N_38925,N_38596);
nor U39571 (N_39571,N_38122,N_38742);
xnor U39572 (N_39572,N_38287,N_38788);
xor U39573 (N_39573,N_38828,N_38432);
and U39574 (N_39574,N_38526,N_38238);
and U39575 (N_39575,N_38115,N_38822);
and U39576 (N_39576,N_38757,N_38493);
nor U39577 (N_39577,N_38942,N_38199);
nor U39578 (N_39578,N_38922,N_38756);
nor U39579 (N_39579,N_38920,N_38535);
xor U39580 (N_39580,N_38568,N_38677);
xnor U39581 (N_39581,N_38395,N_38420);
nand U39582 (N_39582,N_38128,N_38708);
or U39583 (N_39583,N_38687,N_38442);
nor U39584 (N_39584,N_38560,N_38608);
nand U39585 (N_39585,N_38582,N_38145);
or U39586 (N_39586,N_38915,N_38676);
xnor U39587 (N_39587,N_38095,N_38790);
nand U39588 (N_39588,N_38926,N_38184);
and U39589 (N_39589,N_38691,N_38750);
xnor U39590 (N_39590,N_38338,N_38040);
and U39591 (N_39591,N_38582,N_38222);
nor U39592 (N_39592,N_38761,N_38070);
xor U39593 (N_39593,N_38219,N_38804);
or U39594 (N_39594,N_38146,N_38039);
and U39595 (N_39595,N_38554,N_38288);
nand U39596 (N_39596,N_38969,N_38711);
or U39597 (N_39597,N_38374,N_38984);
and U39598 (N_39598,N_38166,N_38276);
and U39599 (N_39599,N_38722,N_38956);
xnor U39600 (N_39600,N_38903,N_38001);
nor U39601 (N_39601,N_38259,N_38034);
and U39602 (N_39602,N_38014,N_38996);
or U39603 (N_39603,N_38893,N_38401);
xnor U39604 (N_39604,N_38346,N_38645);
xnor U39605 (N_39605,N_38542,N_38257);
and U39606 (N_39606,N_38132,N_38568);
nor U39607 (N_39607,N_38179,N_38823);
or U39608 (N_39608,N_38736,N_38733);
or U39609 (N_39609,N_38080,N_38862);
and U39610 (N_39610,N_38072,N_38643);
xnor U39611 (N_39611,N_38986,N_38602);
xnor U39612 (N_39612,N_38246,N_38103);
or U39613 (N_39613,N_38543,N_38437);
or U39614 (N_39614,N_38776,N_38026);
or U39615 (N_39615,N_38260,N_38391);
or U39616 (N_39616,N_38414,N_38043);
xnor U39617 (N_39617,N_38674,N_38113);
and U39618 (N_39618,N_38413,N_38093);
nand U39619 (N_39619,N_38263,N_38138);
or U39620 (N_39620,N_38070,N_38573);
nand U39621 (N_39621,N_38436,N_38551);
nand U39622 (N_39622,N_38354,N_38208);
nand U39623 (N_39623,N_38860,N_38898);
or U39624 (N_39624,N_38992,N_38595);
xnor U39625 (N_39625,N_38416,N_38562);
and U39626 (N_39626,N_38931,N_38000);
nand U39627 (N_39627,N_38399,N_38149);
nor U39628 (N_39628,N_38841,N_38833);
or U39629 (N_39629,N_38130,N_38147);
nor U39630 (N_39630,N_38173,N_38320);
and U39631 (N_39631,N_38423,N_38127);
nor U39632 (N_39632,N_38373,N_38813);
and U39633 (N_39633,N_38407,N_38577);
nor U39634 (N_39634,N_38994,N_38478);
or U39635 (N_39635,N_38126,N_38147);
or U39636 (N_39636,N_38759,N_38069);
nor U39637 (N_39637,N_38095,N_38224);
and U39638 (N_39638,N_38081,N_38933);
xor U39639 (N_39639,N_38475,N_38918);
nor U39640 (N_39640,N_38067,N_38035);
and U39641 (N_39641,N_38763,N_38408);
nand U39642 (N_39642,N_38346,N_38335);
or U39643 (N_39643,N_38376,N_38385);
xnor U39644 (N_39644,N_38365,N_38500);
or U39645 (N_39645,N_38258,N_38728);
or U39646 (N_39646,N_38135,N_38052);
nand U39647 (N_39647,N_38806,N_38224);
xor U39648 (N_39648,N_38250,N_38713);
xnor U39649 (N_39649,N_38134,N_38819);
or U39650 (N_39650,N_38388,N_38032);
and U39651 (N_39651,N_38088,N_38683);
nor U39652 (N_39652,N_38445,N_38374);
nor U39653 (N_39653,N_38878,N_38189);
nor U39654 (N_39654,N_38051,N_38231);
xor U39655 (N_39655,N_38048,N_38209);
nor U39656 (N_39656,N_38407,N_38174);
and U39657 (N_39657,N_38196,N_38404);
or U39658 (N_39658,N_38221,N_38627);
xor U39659 (N_39659,N_38617,N_38275);
and U39660 (N_39660,N_38224,N_38326);
nor U39661 (N_39661,N_38335,N_38928);
or U39662 (N_39662,N_38128,N_38782);
xnor U39663 (N_39663,N_38017,N_38136);
nand U39664 (N_39664,N_38563,N_38965);
nand U39665 (N_39665,N_38117,N_38244);
nor U39666 (N_39666,N_38127,N_38319);
or U39667 (N_39667,N_38748,N_38076);
or U39668 (N_39668,N_38934,N_38207);
nor U39669 (N_39669,N_38871,N_38151);
and U39670 (N_39670,N_38519,N_38155);
nand U39671 (N_39671,N_38449,N_38766);
or U39672 (N_39672,N_38050,N_38975);
and U39673 (N_39673,N_38913,N_38279);
and U39674 (N_39674,N_38326,N_38790);
and U39675 (N_39675,N_38054,N_38900);
and U39676 (N_39676,N_38809,N_38307);
xor U39677 (N_39677,N_38318,N_38870);
and U39678 (N_39678,N_38019,N_38966);
or U39679 (N_39679,N_38521,N_38492);
xnor U39680 (N_39680,N_38714,N_38393);
or U39681 (N_39681,N_38508,N_38684);
nand U39682 (N_39682,N_38721,N_38355);
nand U39683 (N_39683,N_38369,N_38227);
nand U39684 (N_39684,N_38705,N_38416);
nor U39685 (N_39685,N_38274,N_38427);
and U39686 (N_39686,N_38780,N_38218);
xor U39687 (N_39687,N_38836,N_38750);
and U39688 (N_39688,N_38812,N_38535);
nand U39689 (N_39689,N_38491,N_38710);
nand U39690 (N_39690,N_38594,N_38101);
nand U39691 (N_39691,N_38241,N_38959);
or U39692 (N_39692,N_38475,N_38265);
nand U39693 (N_39693,N_38239,N_38652);
nor U39694 (N_39694,N_38963,N_38413);
nor U39695 (N_39695,N_38707,N_38000);
nor U39696 (N_39696,N_38419,N_38901);
and U39697 (N_39697,N_38923,N_38235);
nor U39698 (N_39698,N_38472,N_38192);
and U39699 (N_39699,N_38925,N_38794);
and U39700 (N_39700,N_38192,N_38289);
nor U39701 (N_39701,N_38424,N_38889);
nor U39702 (N_39702,N_38481,N_38355);
or U39703 (N_39703,N_38289,N_38004);
nand U39704 (N_39704,N_38315,N_38434);
or U39705 (N_39705,N_38760,N_38110);
nand U39706 (N_39706,N_38066,N_38571);
nor U39707 (N_39707,N_38767,N_38214);
or U39708 (N_39708,N_38987,N_38420);
or U39709 (N_39709,N_38878,N_38843);
nor U39710 (N_39710,N_38047,N_38675);
xor U39711 (N_39711,N_38383,N_38163);
xnor U39712 (N_39712,N_38011,N_38461);
or U39713 (N_39713,N_38566,N_38591);
or U39714 (N_39714,N_38656,N_38023);
nor U39715 (N_39715,N_38206,N_38160);
nor U39716 (N_39716,N_38939,N_38884);
nand U39717 (N_39717,N_38899,N_38564);
xor U39718 (N_39718,N_38912,N_38491);
xnor U39719 (N_39719,N_38129,N_38879);
and U39720 (N_39720,N_38800,N_38270);
and U39721 (N_39721,N_38498,N_38521);
or U39722 (N_39722,N_38558,N_38754);
and U39723 (N_39723,N_38699,N_38317);
and U39724 (N_39724,N_38622,N_38645);
nand U39725 (N_39725,N_38900,N_38263);
nor U39726 (N_39726,N_38521,N_38756);
or U39727 (N_39727,N_38773,N_38674);
nand U39728 (N_39728,N_38550,N_38299);
nor U39729 (N_39729,N_38610,N_38202);
nand U39730 (N_39730,N_38258,N_38866);
or U39731 (N_39731,N_38849,N_38729);
nor U39732 (N_39732,N_38412,N_38785);
nor U39733 (N_39733,N_38754,N_38380);
and U39734 (N_39734,N_38221,N_38982);
nor U39735 (N_39735,N_38127,N_38814);
and U39736 (N_39736,N_38392,N_38730);
and U39737 (N_39737,N_38848,N_38254);
and U39738 (N_39738,N_38890,N_38072);
xnor U39739 (N_39739,N_38679,N_38462);
and U39740 (N_39740,N_38634,N_38492);
nand U39741 (N_39741,N_38806,N_38747);
xnor U39742 (N_39742,N_38729,N_38063);
nand U39743 (N_39743,N_38988,N_38773);
and U39744 (N_39744,N_38443,N_38871);
and U39745 (N_39745,N_38826,N_38395);
xnor U39746 (N_39746,N_38853,N_38360);
xor U39747 (N_39747,N_38248,N_38017);
nor U39748 (N_39748,N_38823,N_38967);
nand U39749 (N_39749,N_38673,N_38771);
or U39750 (N_39750,N_38106,N_38091);
or U39751 (N_39751,N_38443,N_38147);
xnor U39752 (N_39752,N_38278,N_38496);
nor U39753 (N_39753,N_38409,N_38418);
and U39754 (N_39754,N_38483,N_38972);
or U39755 (N_39755,N_38598,N_38705);
and U39756 (N_39756,N_38971,N_38499);
and U39757 (N_39757,N_38092,N_38311);
and U39758 (N_39758,N_38316,N_38787);
nor U39759 (N_39759,N_38250,N_38257);
xnor U39760 (N_39760,N_38677,N_38037);
or U39761 (N_39761,N_38565,N_38630);
nand U39762 (N_39762,N_38044,N_38726);
and U39763 (N_39763,N_38024,N_38574);
xor U39764 (N_39764,N_38844,N_38784);
and U39765 (N_39765,N_38250,N_38408);
nand U39766 (N_39766,N_38361,N_38447);
nand U39767 (N_39767,N_38401,N_38238);
nor U39768 (N_39768,N_38503,N_38894);
xor U39769 (N_39769,N_38541,N_38890);
xor U39770 (N_39770,N_38169,N_38760);
xor U39771 (N_39771,N_38358,N_38022);
nand U39772 (N_39772,N_38077,N_38986);
and U39773 (N_39773,N_38907,N_38248);
nor U39774 (N_39774,N_38151,N_38254);
or U39775 (N_39775,N_38105,N_38269);
and U39776 (N_39776,N_38202,N_38340);
xnor U39777 (N_39777,N_38923,N_38085);
or U39778 (N_39778,N_38726,N_38448);
and U39779 (N_39779,N_38671,N_38769);
nand U39780 (N_39780,N_38816,N_38253);
nand U39781 (N_39781,N_38441,N_38136);
nand U39782 (N_39782,N_38395,N_38676);
or U39783 (N_39783,N_38524,N_38768);
xnor U39784 (N_39784,N_38150,N_38851);
or U39785 (N_39785,N_38234,N_38284);
nand U39786 (N_39786,N_38961,N_38727);
xor U39787 (N_39787,N_38281,N_38781);
nand U39788 (N_39788,N_38757,N_38240);
and U39789 (N_39789,N_38309,N_38588);
xnor U39790 (N_39790,N_38713,N_38139);
nor U39791 (N_39791,N_38418,N_38142);
xnor U39792 (N_39792,N_38332,N_38665);
and U39793 (N_39793,N_38822,N_38813);
nand U39794 (N_39794,N_38347,N_38536);
nand U39795 (N_39795,N_38667,N_38246);
nand U39796 (N_39796,N_38267,N_38375);
or U39797 (N_39797,N_38944,N_38207);
nand U39798 (N_39798,N_38970,N_38136);
xnor U39799 (N_39799,N_38585,N_38945);
and U39800 (N_39800,N_38159,N_38569);
or U39801 (N_39801,N_38252,N_38936);
nand U39802 (N_39802,N_38995,N_38761);
nand U39803 (N_39803,N_38945,N_38371);
and U39804 (N_39804,N_38001,N_38918);
nor U39805 (N_39805,N_38903,N_38929);
and U39806 (N_39806,N_38303,N_38919);
and U39807 (N_39807,N_38234,N_38348);
nand U39808 (N_39808,N_38724,N_38589);
nor U39809 (N_39809,N_38381,N_38502);
and U39810 (N_39810,N_38896,N_38086);
nor U39811 (N_39811,N_38514,N_38957);
nand U39812 (N_39812,N_38279,N_38770);
xnor U39813 (N_39813,N_38152,N_38420);
xor U39814 (N_39814,N_38623,N_38771);
and U39815 (N_39815,N_38936,N_38050);
nor U39816 (N_39816,N_38224,N_38256);
nand U39817 (N_39817,N_38118,N_38094);
and U39818 (N_39818,N_38712,N_38154);
nand U39819 (N_39819,N_38108,N_38389);
nand U39820 (N_39820,N_38927,N_38601);
and U39821 (N_39821,N_38667,N_38714);
nor U39822 (N_39822,N_38980,N_38200);
xor U39823 (N_39823,N_38939,N_38188);
nand U39824 (N_39824,N_38005,N_38596);
nor U39825 (N_39825,N_38417,N_38429);
and U39826 (N_39826,N_38521,N_38067);
and U39827 (N_39827,N_38897,N_38031);
nand U39828 (N_39828,N_38033,N_38700);
nand U39829 (N_39829,N_38756,N_38745);
xor U39830 (N_39830,N_38082,N_38462);
nand U39831 (N_39831,N_38861,N_38330);
xnor U39832 (N_39832,N_38910,N_38357);
and U39833 (N_39833,N_38206,N_38990);
xor U39834 (N_39834,N_38450,N_38826);
nand U39835 (N_39835,N_38805,N_38902);
nor U39836 (N_39836,N_38762,N_38182);
and U39837 (N_39837,N_38890,N_38851);
nand U39838 (N_39838,N_38608,N_38103);
nand U39839 (N_39839,N_38960,N_38569);
nor U39840 (N_39840,N_38284,N_38884);
nor U39841 (N_39841,N_38107,N_38669);
xor U39842 (N_39842,N_38411,N_38413);
nand U39843 (N_39843,N_38170,N_38863);
xnor U39844 (N_39844,N_38209,N_38829);
xor U39845 (N_39845,N_38156,N_38032);
or U39846 (N_39846,N_38054,N_38037);
xnor U39847 (N_39847,N_38785,N_38847);
xnor U39848 (N_39848,N_38215,N_38559);
nand U39849 (N_39849,N_38345,N_38224);
nand U39850 (N_39850,N_38344,N_38887);
or U39851 (N_39851,N_38416,N_38052);
and U39852 (N_39852,N_38987,N_38773);
or U39853 (N_39853,N_38403,N_38511);
xor U39854 (N_39854,N_38138,N_38845);
and U39855 (N_39855,N_38226,N_38088);
nor U39856 (N_39856,N_38556,N_38495);
and U39857 (N_39857,N_38103,N_38757);
xor U39858 (N_39858,N_38118,N_38592);
xor U39859 (N_39859,N_38525,N_38376);
or U39860 (N_39860,N_38982,N_38532);
nor U39861 (N_39861,N_38215,N_38214);
or U39862 (N_39862,N_38311,N_38831);
xor U39863 (N_39863,N_38615,N_38816);
nand U39864 (N_39864,N_38985,N_38877);
xnor U39865 (N_39865,N_38214,N_38703);
nand U39866 (N_39866,N_38848,N_38008);
or U39867 (N_39867,N_38033,N_38508);
xnor U39868 (N_39868,N_38497,N_38384);
and U39869 (N_39869,N_38722,N_38928);
xnor U39870 (N_39870,N_38923,N_38383);
nor U39871 (N_39871,N_38723,N_38819);
xnor U39872 (N_39872,N_38252,N_38654);
or U39873 (N_39873,N_38365,N_38205);
nor U39874 (N_39874,N_38755,N_38205);
nor U39875 (N_39875,N_38000,N_38039);
and U39876 (N_39876,N_38416,N_38466);
or U39877 (N_39877,N_38015,N_38859);
xnor U39878 (N_39878,N_38513,N_38358);
nand U39879 (N_39879,N_38106,N_38527);
or U39880 (N_39880,N_38992,N_38616);
nand U39881 (N_39881,N_38519,N_38982);
and U39882 (N_39882,N_38621,N_38728);
nand U39883 (N_39883,N_38673,N_38332);
xor U39884 (N_39884,N_38527,N_38516);
nor U39885 (N_39885,N_38712,N_38864);
nand U39886 (N_39886,N_38427,N_38782);
and U39887 (N_39887,N_38237,N_38222);
xor U39888 (N_39888,N_38511,N_38614);
nor U39889 (N_39889,N_38834,N_38117);
nand U39890 (N_39890,N_38303,N_38923);
nor U39891 (N_39891,N_38668,N_38736);
or U39892 (N_39892,N_38307,N_38003);
and U39893 (N_39893,N_38012,N_38053);
and U39894 (N_39894,N_38434,N_38396);
nand U39895 (N_39895,N_38684,N_38118);
or U39896 (N_39896,N_38968,N_38133);
nand U39897 (N_39897,N_38183,N_38636);
or U39898 (N_39898,N_38989,N_38384);
and U39899 (N_39899,N_38785,N_38296);
nor U39900 (N_39900,N_38216,N_38497);
or U39901 (N_39901,N_38080,N_38460);
or U39902 (N_39902,N_38814,N_38935);
and U39903 (N_39903,N_38625,N_38355);
nand U39904 (N_39904,N_38205,N_38207);
and U39905 (N_39905,N_38282,N_38164);
nand U39906 (N_39906,N_38022,N_38566);
nor U39907 (N_39907,N_38318,N_38601);
xor U39908 (N_39908,N_38926,N_38783);
or U39909 (N_39909,N_38173,N_38295);
nor U39910 (N_39910,N_38606,N_38533);
nand U39911 (N_39911,N_38475,N_38757);
nand U39912 (N_39912,N_38611,N_38374);
or U39913 (N_39913,N_38286,N_38646);
nor U39914 (N_39914,N_38681,N_38618);
and U39915 (N_39915,N_38500,N_38708);
nor U39916 (N_39916,N_38977,N_38794);
xor U39917 (N_39917,N_38669,N_38174);
nor U39918 (N_39918,N_38302,N_38473);
nor U39919 (N_39919,N_38716,N_38654);
and U39920 (N_39920,N_38811,N_38115);
or U39921 (N_39921,N_38715,N_38360);
xor U39922 (N_39922,N_38204,N_38562);
or U39923 (N_39923,N_38767,N_38925);
or U39924 (N_39924,N_38338,N_38420);
or U39925 (N_39925,N_38173,N_38776);
nand U39926 (N_39926,N_38098,N_38731);
or U39927 (N_39927,N_38997,N_38892);
nand U39928 (N_39928,N_38245,N_38421);
nand U39929 (N_39929,N_38564,N_38060);
nor U39930 (N_39930,N_38297,N_38665);
or U39931 (N_39931,N_38500,N_38378);
xor U39932 (N_39932,N_38586,N_38249);
and U39933 (N_39933,N_38261,N_38400);
nor U39934 (N_39934,N_38482,N_38088);
nand U39935 (N_39935,N_38423,N_38269);
and U39936 (N_39936,N_38636,N_38055);
nand U39937 (N_39937,N_38378,N_38152);
nand U39938 (N_39938,N_38279,N_38443);
and U39939 (N_39939,N_38931,N_38172);
and U39940 (N_39940,N_38212,N_38682);
nor U39941 (N_39941,N_38905,N_38581);
or U39942 (N_39942,N_38417,N_38676);
or U39943 (N_39943,N_38742,N_38310);
or U39944 (N_39944,N_38196,N_38867);
or U39945 (N_39945,N_38394,N_38051);
nor U39946 (N_39946,N_38595,N_38308);
nand U39947 (N_39947,N_38305,N_38034);
and U39948 (N_39948,N_38727,N_38284);
nor U39949 (N_39949,N_38315,N_38418);
nand U39950 (N_39950,N_38192,N_38477);
xor U39951 (N_39951,N_38418,N_38484);
nor U39952 (N_39952,N_38268,N_38078);
xnor U39953 (N_39953,N_38190,N_38516);
or U39954 (N_39954,N_38622,N_38964);
xor U39955 (N_39955,N_38352,N_38895);
or U39956 (N_39956,N_38989,N_38628);
xnor U39957 (N_39957,N_38156,N_38652);
and U39958 (N_39958,N_38865,N_38198);
and U39959 (N_39959,N_38793,N_38679);
and U39960 (N_39960,N_38063,N_38487);
or U39961 (N_39961,N_38845,N_38434);
xnor U39962 (N_39962,N_38420,N_38486);
xnor U39963 (N_39963,N_38208,N_38325);
nand U39964 (N_39964,N_38302,N_38275);
nand U39965 (N_39965,N_38063,N_38932);
and U39966 (N_39966,N_38967,N_38765);
and U39967 (N_39967,N_38328,N_38460);
nand U39968 (N_39968,N_38752,N_38924);
xor U39969 (N_39969,N_38195,N_38887);
xor U39970 (N_39970,N_38612,N_38622);
or U39971 (N_39971,N_38703,N_38436);
nor U39972 (N_39972,N_38614,N_38393);
and U39973 (N_39973,N_38028,N_38150);
or U39974 (N_39974,N_38071,N_38871);
nor U39975 (N_39975,N_38766,N_38966);
or U39976 (N_39976,N_38413,N_38924);
and U39977 (N_39977,N_38211,N_38712);
nand U39978 (N_39978,N_38226,N_38018);
nor U39979 (N_39979,N_38408,N_38313);
xor U39980 (N_39980,N_38877,N_38335);
nand U39981 (N_39981,N_38199,N_38948);
and U39982 (N_39982,N_38828,N_38486);
nand U39983 (N_39983,N_38955,N_38708);
nor U39984 (N_39984,N_38756,N_38517);
and U39985 (N_39985,N_38495,N_38001);
and U39986 (N_39986,N_38261,N_38310);
xnor U39987 (N_39987,N_38441,N_38122);
xnor U39988 (N_39988,N_38260,N_38168);
xor U39989 (N_39989,N_38732,N_38786);
or U39990 (N_39990,N_38220,N_38567);
nor U39991 (N_39991,N_38508,N_38649);
and U39992 (N_39992,N_38120,N_38797);
and U39993 (N_39993,N_38967,N_38876);
nor U39994 (N_39994,N_38789,N_38994);
nand U39995 (N_39995,N_38972,N_38801);
and U39996 (N_39996,N_38271,N_38736);
nand U39997 (N_39997,N_38175,N_38802);
nand U39998 (N_39998,N_38904,N_38028);
or U39999 (N_39999,N_38329,N_38106);
nand U40000 (N_40000,N_39485,N_39273);
nor U40001 (N_40001,N_39839,N_39393);
nand U40002 (N_40002,N_39910,N_39780);
and U40003 (N_40003,N_39755,N_39879);
nor U40004 (N_40004,N_39191,N_39529);
and U40005 (N_40005,N_39306,N_39739);
nand U40006 (N_40006,N_39475,N_39614);
or U40007 (N_40007,N_39868,N_39387);
or U40008 (N_40008,N_39491,N_39501);
and U40009 (N_40009,N_39092,N_39415);
nor U40010 (N_40010,N_39824,N_39423);
and U40011 (N_40011,N_39747,N_39625);
xnor U40012 (N_40012,N_39714,N_39634);
or U40013 (N_40013,N_39935,N_39914);
and U40014 (N_40014,N_39198,N_39759);
or U40015 (N_40015,N_39336,N_39401);
nor U40016 (N_40016,N_39568,N_39972);
and U40017 (N_40017,N_39892,N_39621);
or U40018 (N_40018,N_39608,N_39451);
and U40019 (N_40019,N_39495,N_39037);
xor U40020 (N_40020,N_39808,N_39090);
or U40021 (N_40021,N_39407,N_39158);
nand U40022 (N_40022,N_39321,N_39885);
nor U40023 (N_40023,N_39760,N_39711);
xnor U40024 (N_40024,N_39968,N_39999);
nor U40025 (N_40025,N_39987,N_39442);
and U40026 (N_40026,N_39834,N_39362);
and U40027 (N_40027,N_39317,N_39623);
nor U40028 (N_40028,N_39505,N_39943);
xnor U40029 (N_40029,N_39278,N_39216);
nor U40030 (N_40030,N_39514,N_39984);
nor U40031 (N_40031,N_39311,N_39165);
and U40032 (N_40032,N_39603,N_39752);
nor U40033 (N_40033,N_39229,N_39671);
nand U40034 (N_40034,N_39499,N_39771);
nand U40035 (N_40035,N_39497,N_39453);
or U40036 (N_40036,N_39595,N_39384);
xor U40037 (N_40037,N_39590,N_39955);
xnor U40038 (N_40038,N_39633,N_39537);
xnor U40039 (N_40039,N_39149,N_39325);
nand U40040 (N_40040,N_39443,N_39316);
nor U40041 (N_40041,N_39861,N_39378);
and U40042 (N_40042,N_39795,N_39333);
xor U40043 (N_40043,N_39836,N_39656);
xor U40044 (N_40044,N_39267,N_39779);
nand U40045 (N_40045,N_39255,N_39772);
nor U40046 (N_40046,N_39648,N_39166);
nor U40047 (N_40047,N_39732,N_39129);
and U40048 (N_40048,N_39519,N_39189);
nor U40049 (N_40049,N_39891,N_39706);
nor U40050 (N_40050,N_39734,N_39439);
and U40051 (N_40051,N_39469,N_39234);
or U40052 (N_40052,N_39111,N_39061);
nand U40053 (N_40053,N_39350,N_39639);
or U40054 (N_40054,N_39328,N_39632);
or U40055 (N_40055,N_39337,N_39877);
nor U40056 (N_40056,N_39339,N_39026);
and U40057 (N_40057,N_39182,N_39421);
xnor U40058 (N_40058,N_39658,N_39146);
and U40059 (N_40059,N_39109,N_39853);
and U40060 (N_40060,N_39054,N_39629);
nand U40061 (N_40061,N_39386,N_39847);
or U40062 (N_40062,N_39265,N_39017);
nor U40063 (N_40063,N_39813,N_39410);
and U40064 (N_40064,N_39526,N_39638);
or U40065 (N_40065,N_39480,N_39425);
and U40066 (N_40066,N_39087,N_39261);
or U40067 (N_40067,N_39684,N_39073);
nor U40068 (N_40068,N_39967,N_39918);
xor U40069 (N_40069,N_39607,N_39749);
or U40070 (N_40070,N_39997,N_39327);
xnor U40071 (N_40071,N_39677,N_39498);
xor U40072 (N_40072,N_39855,N_39019);
and U40073 (N_40073,N_39996,N_39721);
nor U40074 (N_40074,N_39377,N_39516);
xnor U40075 (N_40075,N_39181,N_39678);
nor U40076 (N_40076,N_39144,N_39399);
nor U40077 (N_40077,N_39823,N_39245);
xnor U40078 (N_40078,N_39252,N_39820);
xnor U40079 (N_40079,N_39150,N_39661);
or U40080 (N_40080,N_39581,N_39496);
xnor U40081 (N_40081,N_39919,N_39707);
and U40082 (N_40082,N_39976,N_39123);
nor U40083 (N_40083,N_39735,N_39110);
and U40084 (N_40084,N_39553,N_39483);
and U40085 (N_40085,N_39571,N_39986);
nand U40086 (N_40086,N_39010,N_39942);
nor U40087 (N_40087,N_39578,N_39355);
xnor U40088 (N_40088,N_39689,N_39507);
xor U40089 (N_40089,N_39356,N_39064);
and U40090 (N_40090,N_39322,N_39540);
or U40091 (N_40091,N_39047,N_39596);
or U40092 (N_40092,N_39254,N_39107);
nand U40093 (N_40093,N_39650,N_39391);
nor U40094 (N_40094,N_39601,N_39418);
nand U40095 (N_40095,N_39988,N_39736);
and U40096 (N_40096,N_39725,N_39408);
and U40097 (N_40097,N_39978,N_39295);
xor U40098 (N_40098,N_39679,N_39081);
and U40099 (N_40099,N_39330,N_39115);
nand U40100 (N_40100,N_39890,N_39610);
xnor U40101 (N_40101,N_39645,N_39649);
nor U40102 (N_40102,N_39782,N_39096);
nand U40103 (N_40103,N_39164,N_39600);
xnor U40104 (N_40104,N_39703,N_39214);
or U40105 (N_40105,N_39863,N_39354);
and U40106 (N_40106,N_39768,N_39597);
and U40107 (N_40107,N_39412,N_39687);
nand U40108 (N_40108,N_39750,N_39361);
or U40109 (N_40109,N_39402,N_39758);
or U40110 (N_40110,N_39702,N_39484);
xor U40111 (N_40111,N_39358,N_39205);
xor U40112 (N_40112,N_39113,N_39641);
xor U40113 (N_40113,N_39127,N_39449);
nor U40114 (N_40114,N_39085,N_39077);
nand U40115 (N_40115,N_39023,N_39559);
or U40116 (N_40116,N_39913,N_39681);
xor U40117 (N_40117,N_39331,N_39697);
nand U40118 (N_40118,N_39688,N_39811);
nand U40119 (N_40119,N_39288,N_39618);
or U40120 (N_40120,N_39270,N_39959);
and U40121 (N_40121,N_39276,N_39635);
xor U40122 (N_40122,N_39414,N_39977);
nand U40123 (N_40123,N_39664,N_39277);
nor U40124 (N_40124,N_39659,N_39598);
nand U40125 (N_40125,N_39726,N_39227);
nand U40126 (N_40126,N_39131,N_39285);
or U40127 (N_40127,N_39550,N_39046);
or U40128 (N_40128,N_39852,N_39945);
or U40129 (N_40129,N_39141,N_39134);
and U40130 (N_40130,N_39669,N_39920);
nand U40131 (N_40131,N_39944,N_39591);
nor U40132 (N_40132,N_39695,N_39041);
nor U40133 (N_40133,N_39366,N_39178);
and U40134 (N_40134,N_39812,N_39546);
xor U40135 (N_40135,N_39124,N_39825);
nor U40136 (N_40136,N_39236,N_39381);
or U40137 (N_40137,N_39843,N_39062);
nand U40138 (N_40138,N_39922,N_39156);
or U40139 (N_40139,N_39136,N_39477);
nor U40140 (N_40140,N_39209,N_39512);
nor U40141 (N_40141,N_39912,N_39076);
nand U40142 (N_40142,N_39867,N_39958);
or U40143 (N_40143,N_39733,N_39045);
xor U40144 (N_40144,N_39617,N_39347);
xor U40145 (N_40145,N_39120,N_39441);
or U40146 (N_40146,N_39523,N_39798);
and U40147 (N_40147,N_39098,N_39508);
and U40148 (N_40148,N_39201,N_39130);
nor U40149 (N_40149,N_39057,N_39175);
and U40150 (N_40150,N_39646,N_39338);
nand U40151 (N_40151,N_39332,N_39173);
and U40152 (N_40152,N_39493,N_39564);
or U40153 (N_40153,N_39615,N_39520);
nand U40154 (N_40154,N_39187,N_39280);
or U40155 (N_40155,N_39970,N_39680);
nor U40156 (N_40156,N_39713,N_39864);
or U40157 (N_40157,N_39690,N_39653);
or U40158 (N_40158,N_39940,N_39761);
nand U40159 (N_40159,N_39777,N_39886);
xor U40160 (N_40160,N_39655,N_39799);
or U40161 (N_40161,N_39313,N_39670);
nor U40162 (N_40162,N_39791,N_39217);
nor U40163 (N_40163,N_39506,N_39434);
or U40164 (N_40164,N_39230,N_39872);
and U40165 (N_40165,N_39095,N_39479);
nor U40166 (N_40166,N_39049,N_39374);
nand U40167 (N_40167,N_39592,N_39562);
and U40168 (N_40168,N_39902,N_39800);
and U40169 (N_40169,N_39905,N_39125);
nor U40170 (N_40170,N_39642,N_39140);
and U40171 (N_40171,N_39396,N_39938);
and U40172 (N_40172,N_39203,N_39478);
and U40173 (N_40173,N_39993,N_39998);
xor U40174 (N_40174,N_39962,N_39226);
and U40175 (N_40175,N_39360,N_39079);
and U40176 (N_40176,N_39666,N_39225);
xnor U40177 (N_40177,N_39427,N_39348);
nor U40178 (N_40178,N_39792,N_39405);
xnor U40179 (N_40179,N_39980,N_39168);
xor U40180 (N_40180,N_39574,N_39583);
nor U40181 (N_40181,N_39738,N_39424);
or U40182 (N_40182,N_39860,N_39193);
and U40183 (N_40183,N_39036,N_39207);
and U40184 (N_40184,N_39024,N_39841);
nor U40185 (N_40185,N_39246,N_39630);
nor U40186 (N_40186,N_39065,N_39161);
and U40187 (N_40187,N_39253,N_39712);
or U40188 (N_40188,N_39139,N_39627);
and U40189 (N_40189,N_39305,N_39807);
xnor U40190 (N_40190,N_39232,N_39137);
and U40191 (N_40191,N_39152,N_39740);
or U40192 (N_40192,N_39455,N_39199);
or U40193 (N_40193,N_39731,N_39138);
and U40194 (N_40194,N_39882,N_39809);
nor U40195 (N_40195,N_39119,N_39832);
and U40196 (N_40196,N_39566,N_39221);
xor U40197 (N_40197,N_39488,N_39513);
or U40198 (N_40198,N_39774,N_39174);
or U40199 (N_40199,N_39981,N_39042);
nor U40200 (N_40200,N_39710,N_39558);
or U40201 (N_40201,N_39014,N_39929);
or U40202 (N_40202,N_39547,N_39835);
xnor U40203 (N_40203,N_39476,N_39619);
and U40204 (N_40204,N_39510,N_39640);
or U40205 (N_40205,N_39925,N_39783);
nand U40206 (N_40206,N_39793,N_39934);
or U40207 (N_40207,N_39030,N_39050);
nand U40208 (N_40208,N_39091,N_39541);
and U40209 (N_40209,N_39694,N_39300);
or U40210 (N_40210,N_39404,N_39856);
xor U40211 (N_40211,N_39433,N_39428);
or U40212 (N_40212,N_39818,N_39237);
or U40213 (N_40213,N_39326,N_39373);
and U40214 (N_40214,N_39921,N_39586);
and U40215 (N_40215,N_39185,N_39816);
xor U40216 (N_40216,N_39257,N_39580);
nand U40217 (N_40217,N_39100,N_39027);
or U40218 (N_40218,N_39375,N_39685);
and U40219 (N_40219,N_39471,N_39522);
xor U40220 (N_40220,N_39069,N_39924);
nor U40221 (N_40221,N_39588,N_39419);
nor U40222 (N_40222,N_39930,N_39440);
xnor U40223 (N_40223,N_39990,N_39622);
or U40224 (N_40224,N_39991,N_39197);
or U40225 (N_40225,N_39275,N_39299);
xnor U40226 (N_40226,N_39570,N_39624);
nor U40227 (N_40227,N_39298,N_39936);
and U40228 (N_40228,N_39579,N_39143);
nor U40229 (N_40229,N_39416,N_39587);
nand U40230 (N_40230,N_39437,N_39775);
and U40231 (N_40231,N_39517,N_39033);
and U40232 (N_40232,N_39163,N_39492);
nor U40233 (N_40233,N_39662,N_39866);
nand U40234 (N_40234,N_39481,N_39859);
xnor U40235 (N_40235,N_39542,N_39900);
xnor U40236 (N_40236,N_39371,N_39390);
nor U40237 (N_40237,N_39838,N_39605);
xor U40238 (N_40238,N_39911,N_39701);
nor U40239 (N_40239,N_39281,N_39950);
nor U40240 (N_40240,N_39211,N_39643);
nand U40241 (N_40241,N_39693,N_39154);
nand U40242 (N_40242,N_39284,N_39457);
or U40243 (N_40243,N_39323,N_39948);
nor U40244 (N_40244,N_39611,N_39956);
or U40245 (N_40245,N_39059,N_39781);
and U40246 (N_40246,N_39392,N_39283);
nor U40247 (N_40247,N_39487,N_39367);
or U40248 (N_40248,N_39654,N_39682);
nand U40249 (N_40249,N_39828,N_39094);
or U40250 (N_40250,N_39698,N_39887);
nor U40251 (N_40251,N_39363,N_39353);
nand U40252 (N_40252,N_39088,N_39031);
nand U40253 (N_40253,N_39575,N_39233);
nand U40254 (N_40254,N_39531,N_39224);
nand U40255 (N_40255,N_39420,N_39906);
xor U40256 (N_40256,N_39829,N_39121);
or U40257 (N_40257,N_39965,N_39982);
nand U40258 (N_40258,N_39971,N_39345);
or U40259 (N_40259,N_39446,N_39683);
and U40260 (N_40260,N_39573,N_39901);
nand U40261 (N_40261,N_39709,N_39204);
nand U40262 (N_40262,N_39222,N_39889);
nand U40263 (N_40263,N_39845,N_39857);
nor U40264 (N_40264,N_39370,N_39025);
xnor U40265 (N_40265,N_39745,N_39368);
or U40266 (N_40266,N_39286,N_39552);
nor U40267 (N_40267,N_39862,N_39894);
nor U40268 (N_40268,N_39179,N_39636);
xnor U40269 (N_40269,N_39034,N_39274);
or U40270 (N_40270,N_39456,N_39751);
nor U40271 (N_40271,N_39258,N_39803);
xor U40272 (N_40272,N_39533,N_39675);
nand U40273 (N_40273,N_39310,N_39794);
and U40274 (N_40274,N_39715,N_39383);
or U40275 (N_40275,N_39118,N_39318);
and U40276 (N_40276,N_39644,N_39206);
nor U40277 (N_40277,N_39490,N_39068);
nand U40278 (N_40278,N_39078,N_39448);
nand U40279 (N_40279,N_39931,N_39369);
and U40280 (N_40280,N_39122,N_39917);
xor U40281 (N_40281,N_39320,N_39251);
nand U40282 (N_40282,N_39303,N_39953);
or U40283 (N_40283,N_39567,N_39035);
xor U40284 (N_40284,N_39007,N_39947);
and U40285 (N_40285,N_39022,N_39223);
or U40286 (N_40286,N_39831,N_39409);
nor U40287 (N_40287,N_39389,N_39458);
xnor U40288 (N_40288,N_39473,N_39244);
nor U40289 (N_40289,N_39296,N_39021);
nor U40290 (N_40290,N_39974,N_39932);
xor U40291 (N_40291,N_39171,N_39904);
nor U40292 (N_40292,N_39543,N_39874);
nand U40293 (N_40293,N_39840,N_39302);
nor U40294 (N_40294,N_39005,N_39279);
nor U40295 (N_40295,N_39915,N_39815);
and U40296 (N_40296,N_39786,N_39470);
and U40297 (N_40297,N_39833,N_39202);
or U40298 (N_40298,N_39927,N_39013);
nand U40299 (N_40299,N_39663,N_39534);
nand U40300 (N_40300,N_39003,N_39742);
or U40301 (N_40301,N_39242,N_39044);
or U40302 (N_40302,N_39063,N_39875);
nor U40303 (N_40303,N_39612,N_39511);
nor U40304 (N_40304,N_39213,N_39746);
nor U40305 (N_40305,N_39324,N_39357);
or U40306 (N_40306,N_39268,N_39674);
or U40307 (N_40307,N_39099,N_39071);
nand U40308 (N_40308,N_39952,N_39103);
nor U40309 (N_40309,N_39756,N_39992);
xor U40310 (N_40310,N_39235,N_39018);
nor U40311 (N_40311,N_39960,N_39528);
or U40312 (N_40312,N_39557,N_39183);
or U40313 (N_40313,N_39444,N_39292);
nand U40314 (N_40314,N_39873,N_39002);
nor U40315 (N_40315,N_39153,N_39822);
or U40316 (N_40316,N_39728,N_39926);
nor U40317 (N_40317,N_39604,N_39814);
or U40318 (N_40318,N_39539,N_39380);
or U40319 (N_40319,N_39504,N_39436);
nand U40320 (N_40320,N_39538,N_39723);
nand U40321 (N_40321,N_39784,N_39716);
xnor U40322 (N_40322,N_39072,N_39720);
and U40323 (N_40323,N_39946,N_39148);
nand U40324 (N_40324,N_39613,N_39340);
nand U40325 (N_40325,N_39544,N_39105);
xnor U40326 (N_40326,N_39264,N_39341);
and U40327 (N_40327,N_39382,N_39256);
xor U40328 (N_40328,N_39351,N_39397);
xnor U40329 (N_40329,N_39097,N_39116);
or U40330 (N_40330,N_39015,N_39773);
nor U40331 (N_40331,N_39385,N_39754);
and U40332 (N_40332,N_39626,N_39797);
and U40333 (N_40333,N_39527,N_39218);
nand U40334 (N_40334,N_39142,N_39718);
or U40335 (N_40335,N_39837,N_39447);
or U40336 (N_40336,N_39432,N_39169);
or U40337 (N_40337,N_39101,N_39854);
nor U40338 (N_40338,N_39923,N_39190);
nor U40339 (N_40339,N_39472,N_39796);
nor U40340 (N_40340,N_39609,N_39177);
xor U40341 (N_40341,N_39764,N_39194);
xnor U40342 (N_40342,N_39766,N_39880);
or U40343 (N_40343,N_39135,N_39727);
nand U40344 (N_40344,N_39114,N_39240);
xor U40345 (N_40345,N_39060,N_39494);
or U40346 (N_40346,N_39459,N_39200);
or U40347 (N_40347,N_39430,N_39212);
nand U40348 (N_40348,N_39994,N_39851);
or U40349 (N_40349,N_39266,N_39093);
nand U40350 (N_40350,N_39665,N_39975);
or U40351 (N_40351,N_39561,N_39569);
or U40352 (N_40352,N_39802,N_39309);
xor U40353 (N_40353,N_39565,N_39184);
xnor U40354 (N_40354,N_39445,N_39667);
nand U40355 (N_40355,N_39028,N_39673);
xor U40356 (N_40356,N_39220,N_39787);
or U40357 (N_40357,N_39038,N_39770);
nor U40358 (N_40358,N_39379,N_39941);
nor U40359 (N_40359,N_39672,N_39536);
or U40360 (N_40360,N_39343,N_39884);
or U40361 (N_40361,N_39730,N_39269);
nor U40362 (N_40362,N_39067,N_39112);
or U40363 (N_40363,N_39468,N_39810);
nand U40364 (N_40364,N_39817,N_39388);
nand U40365 (N_40365,N_39250,N_39188);
and U40366 (N_40366,N_39249,N_39006);
nand U40367 (N_40367,N_39949,N_39748);
nand U40368 (N_40368,N_39084,N_39830);
and U40369 (N_40369,N_39785,N_39668);
or U40370 (N_40370,N_39502,N_39599);
nor U40371 (N_40371,N_39753,N_39699);
nand U40372 (N_40372,N_39957,N_39145);
xnor U40373 (N_40373,N_39403,N_39287);
and U40374 (N_40374,N_39554,N_39602);
or U40375 (N_40375,N_39372,N_39461);
and U40376 (N_40376,N_39460,N_39263);
and U40377 (N_40377,N_39637,N_39208);
xnor U40378 (N_40378,N_39040,N_39176);
nand U40379 (N_40379,N_39053,N_39951);
or U40380 (N_40380,N_39308,N_39705);
and U40381 (N_40381,N_39763,N_39966);
xor U40382 (N_40382,N_39429,N_39744);
xnor U40383 (N_40383,N_39294,N_39083);
xor U40384 (N_40384,N_39307,N_39524);
xor U40385 (N_40385,N_39192,N_39104);
nor U40386 (N_40386,N_39417,N_39954);
nand U40387 (N_40387,N_39589,N_39692);
nor U40388 (N_40388,N_39102,N_39908);
xnor U40389 (N_40389,N_39011,N_39248);
nand U40390 (N_40390,N_39535,N_39909);
xnor U40391 (N_40391,N_39086,N_39651);
nand U40392 (N_40392,N_39743,N_39172);
or U40393 (N_40393,N_39963,N_39961);
nand U40394 (N_40394,N_39757,N_39319);
xnor U40395 (N_40395,N_39969,N_39532);
nand U40396 (N_40396,N_39160,N_39686);
and U40397 (N_40397,N_39907,N_39406);
nor U40398 (N_40398,N_39676,N_39474);
and U40399 (N_40399,N_39074,N_39349);
and U40400 (N_40400,N_39515,N_39876);
nor U40401 (N_40401,N_39708,N_39259);
nor U40402 (N_40402,N_39582,N_39241);
or U40403 (N_40403,N_39620,N_39549);
xor U40404 (N_40404,N_39821,N_39555);
and U40405 (N_40405,N_39466,N_39260);
nor U40406 (N_40406,N_39467,N_39973);
nand U40407 (N_40407,N_39008,N_39228);
nand U40408 (N_40408,N_39186,N_39422);
nand U40409 (N_40409,N_39334,N_39762);
xor U40410 (N_40410,N_39717,N_39411);
or U40411 (N_40411,N_39767,N_39395);
nand U40412 (N_40412,N_39584,N_39219);
nand U40413 (N_40413,N_39737,N_39858);
nor U40414 (N_40414,N_39070,N_39039);
and U40415 (N_40415,N_39126,N_39147);
and U40416 (N_40416,N_39431,N_39167);
nor U40417 (N_40417,N_39765,N_39525);
nand U40418 (N_40418,N_39000,N_39464);
and U40419 (N_40419,N_39572,N_39870);
or U40420 (N_40420,N_39365,N_39700);
or U40421 (N_40421,N_39089,N_39180);
or U40422 (N_40422,N_39315,N_39359);
or U40423 (N_40423,N_39056,N_39462);
or U40424 (N_40424,N_39196,N_39652);
or U40425 (N_40425,N_39082,N_39724);
xor U40426 (N_40426,N_39329,N_39314);
nor U40427 (N_40427,N_39210,N_39157);
or U40428 (N_40428,N_39729,N_39593);
nand U40429 (N_40429,N_39983,N_39577);
and U40430 (N_40430,N_39801,N_39848);
nand U40431 (N_40431,N_39398,N_39606);
nand U40432 (N_40432,N_39342,N_39151);
nor U40433 (N_40433,N_39482,N_39238);
nand U40434 (N_40434,N_39438,N_39413);
nand U40435 (N_40435,N_39790,N_39888);
nand U40436 (N_40436,N_39048,N_39108);
xnor U40437 (N_40437,N_39696,N_39043);
and U40438 (N_40438,N_39304,N_39290);
or U40439 (N_40439,N_39871,N_39806);
or U40440 (N_40440,N_39080,N_39297);
nand U40441 (N_40441,N_39691,N_39301);
and U40442 (N_40442,N_39647,N_39895);
and U40443 (N_40443,N_39776,N_39995);
nor U40444 (N_40444,N_39530,N_39521);
nand U40445 (N_40445,N_39881,N_39159);
nand U40446 (N_40446,N_39016,N_39452);
xnor U40447 (N_40447,N_39400,N_39789);
and U40448 (N_40448,N_39518,N_39029);
nand U40449 (N_40449,N_39075,N_39020);
xor U40450 (N_40450,N_39560,N_39545);
and U40451 (N_40451,N_39939,N_39293);
and U40452 (N_40452,N_39247,N_39704);
or U40453 (N_40453,N_39271,N_39576);
nor U40454 (N_40454,N_39878,N_39660);
nand U40455 (N_40455,N_39231,N_39933);
nor U40456 (N_40456,N_39500,N_39722);
xor U40457 (N_40457,N_39051,N_39869);
nand U40458 (N_40458,N_39117,N_39364);
nor U40459 (N_40459,N_39376,N_39548);
nand U40460 (N_40460,N_39985,N_39465);
and U40461 (N_40461,N_39804,N_39594);
nand U40462 (N_40462,N_39291,N_39195);
xor U40463 (N_40463,N_39897,N_39503);
or U40464 (N_40464,N_39032,N_39162);
and U40465 (N_40465,N_39898,N_39842);
nand U40466 (N_40466,N_39155,N_39964);
nand U40467 (N_40467,N_39058,N_39896);
nor U40468 (N_40468,N_39616,N_39631);
nand U40469 (N_40469,N_39883,N_39335);
xnor U40470 (N_40470,N_39312,N_39979);
nand U40471 (N_40471,N_39551,N_39585);
xnor U40472 (N_40472,N_39657,N_39489);
nand U40473 (N_40473,N_39628,N_39805);
and U40474 (N_40474,N_39004,N_39066);
xor U40475 (N_40475,N_39450,N_39719);
nor U40476 (N_40476,N_39106,N_39128);
nand U40477 (N_40477,N_39394,N_39819);
or U40478 (N_40478,N_39132,N_39903);
nand U40479 (N_40479,N_39769,N_39170);
nor U40480 (N_40480,N_39741,N_39001);
xnor U40481 (N_40481,N_39989,N_39937);
xor U40482 (N_40482,N_39272,N_39849);
or U40483 (N_40483,N_39509,N_39262);
nor U40484 (N_40484,N_39916,N_39844);
xor U40485 (N_40485,N_39352,N_39788);
nor U40486 (N_40486,N_39055,N_39893);
nor U40487 (N_40487,N_39463,N_39865);
nor U40488 (N_40488,N_39009,N_39239);
nand U40489 (N_40489,N_39846,N_39928);
nor U40490 (N_40490,N_39346,N_39827);
xnor U40491 (N_40491,N_39243,N_39850);
xnor U40492 (N_40492,N_39435,N_39289);
nor U40493 (N_40493,N_39563,N_39778);
and U40494 (N_40494,N_39133,N_39426);
nand U40495 (N_40495,N_39012,N_39282);
nor U40496 (N_40496,N_39486,N_39826);
and U40497 (N_40497,N_39454,N_39556);
xnor U40498 (N_40498,N_39215,N_39344);
nand U40499 (N_40499,N_39052,N_39899);
xnor U40500 (N_40500,N_39573,N_39738);
nor U40501 (N_40501,N_39405,N_39461);
xnor U40502 (N_40502,N_39855,N_39659);
nor U40503 (N_40503,N_39849,N_39579);
and U40504 (N_40504,N_39926,N_39474);
xnor U40505 (N_40505,N_39425,N_39346);
nor U40506 (N_40506,N_39600,N_39921);
or U40507 (N_40507,N_39308,N_39530);
and U40508 (N_40508,N_39929,N_39698);
nor U40509 (N_40509,N_39287,N_39484);
or U40510 (N_40510,N_39184,N_39400);
nand U40511 (N_40511,N_39804,N_39785);
nand U40512 (N_40512,N_39655,N_39337);
or U40513 (N_40513,N_39761,N_39309);
or U40514 (N_40514,N_39953,N_39925);
xor U40515 (N_40515,N_39423,N_39082);
xnor U40516 (N_40516,N_39813,N_39661);
and U40517 (N_40517,N_39171,N_39696);
xor U40518 (N_40518,N_39021,N_39614);
nor U40519 (N_40519,N_39554,N_39864);
and U40520 (N_40520,N_39621,N_39125);
nor U40521 (N_40521,N_39119,N_39724);
nor U40522 (N_40522,N_39801,N_39850);
xnor U40523 (N_40523,N_39669,N_39413);
and U40524 (N_40524,N_39533,N_39288);
and U40525 (N_40525,N_39461,N_39035);
and U40526 (N_40526,N_39199,N_39809);
nand U40527 (N_40527,N_39371,N_39521);
nor U40528 (N_40528,N_39374,N_39655);
xnor U40529 (N_40529,N_39083,N_39754);
xnor U40530 (N_40530,N_39744,N_39509);
xor U40531 (N_40531,N_39544,N_39629);
nand U40532 (N_40532,N_39483,N_39343);
and U40533 (N_40533,N_39388,N_39527);
and U40534 (N_40534,N_39408,N_39809);
xnor U40535 (N_40535,N_39550,N_39077);
or U40536 (N_40536,N_39860,N_39375);
and U40537 (N_40537,N_39283,N_39282);
xnor U40538 (N_40538,N_39005,N_39579);
nor U40539 (N_40539,N_39356,N_39032);
nor U40540 (N_40540,N_39374,N_39502);
nand U40541 (N_40541,N_39894,N_39472);
and U40542 (N_40542,N_39046,N_39852);
and U40543 (N_40543,N_39792,N_39546);
or U40544 (N_40544,N_39142,N_39923);
and U40545 (N_40545,N_39509,N_39865);
nor U40546 (N_40546,N_39875,N_39664);
and U40547 (N_40547,N_39039,N_39625);
xor U40548 (N_40548,N_39364,N_39890);
nor U40549 (N_40549,N_39456,N_39397);
xnor U40550 (N_40550,N_39353,N_39921);
and U40551 (N_40551,N_39286,N_39371);
xor U40552 (N_40552,N_39464,N_39141);
nor U40553 (N_40553,N_39614,N_39332);
xor U40554 (N_40554,N_39292,N_39116);
nand U40555 (N_40555,N_39234,N_39637);
nand U40556 (N_40556,N_39450,N_39096);
nor U40557 (N_40557,N_39773,N_39131);
xor U40558 (N_40558,N_39983,N_39338);
and U40559 (N_40559,N_39450,N_39031);
xnor U40560 (N_40560,N_39055,N_39789);
nor U40561 (N_40561,N_39319,N_39104);
and U40562 (N_40562,N_39185,N_39768);
xnor U40563 (N_40563,N_39268,N_39898);
and U40564 (N_40564,N_39577,N_39419);
nand U40565 (N_40565,N_39172,N_39204);
nor U40566 (N_40566,N_39720,N_39631);
xnor U40567 (N_40567,N_39747,N_39888);
nand U40568 (N_40568,N_39044,N_39990);
nor U40569 (N_40569,N_39902,N_39639);
or U40570 (N_40570,N_39660,N_39390);
xnor U40571 (N_40571,N_39852,N_39228);
or U40572 (N_40572,N_39345,N_39659);
nor U40573 (N_40573,N_39590,N_39313);
or U40574 (N_40574,N_39408,N_39148);
or U40575 (N_40575,N_39381,N_39476);
nor U40576 (N_40576,N_39464,N_39439);
nor U40577 (N_40577,N_39498,N_39361);
or U40578 (N_40578,N_39975,N_39846);
or U40579 (N_40579,N_39723,N_39993);
nand U40580 (N_40580,N_39170,N_39258);
or U40581 (N_40581,N_39500,N_39286);
and U40582 (N_40582,N_39076,N_39131);
xnor U40583 (N_40583,N_39206,N_39339);
or U40584 (N_40584,N_39487,N_39973);
or U40585 (N_40585,N_39982,N_39352);
or U40586 (N_40586,N_39758,N_39018);
and U40587 (N_40587,N_39818,N_39210);
or U40588 (N_40588,N_39205,N_39118);
or U40589 (N_40589,N_39349,N_39508);
nand U40590 (N_40590,N_39591,N_39455);
nor U40591 (N_40591,N_39291,N_39215);
or U40592 (N_40592,N_39684,N_39818);
nor U40593 (N_40593,N_39722,N_39355);
nor U40594 (N_40594,N_39596,N_39321);
xor U40595 (N_40595,N_39788,N_39612);
and U40596 (N_40596,N_39825,N_39813);
xnor U40597 (N_40597,N_39561,N_39321);
and U40598 (N_40598,N_39305,N_39231);
and U40599 (N_40599,N_39156,N_39653);
nor U40600 (N_40600,N_39121,N_39953);
or U40601 (N_40601,N_39481,N_39813);
and U40602 (N_40602,N_39420,N_39242);
or U40603 (N_40603,N_39394,N_39747);
or U40604 (N_40604,N_39730,N_39616);
nand U40605 (N_40605,N_39002,N_39578);
nor U40606 (N_40606,N_39648,N_39535);
nor U40607 (N_40607,N_39395,N_39503);
or U40608 (N_40608,N_39591,N_39385);
xnor U40609 (N_40609,N_39568,N_39015);
xor U40610 (N_40610,N_39445,N_39923);
nand U40611 (N_40611,N_39313,N_39911);
nor U40612 (N_40612,N_39015,N_39825);
xnor U40613 (N_40613,N_39769,N_39254);
and U40614 (N_40614,N_39359,N_39113);
nand U40615 (N_40615,N_39750,N_39820);
or U40616 (N_40616,N_39730,N_39747);
and U40617 (N_40617,N_39422,N_39776);
or U40618 (N_40618,N_39069,N_39769);
nor U40619 (N_40619,N_39016,N_39479);
and U40620 (N_40620,N_39206,N_39944);
or U40621 (N_40621,N_39630,N_39395);
and U40622 (N_40622,N_39043,N_39937);
xor U40623 (N_40623,N_39001,N_39495);
nor U40624 (N_40624,N_39245,N_39098);
nor U40625 (N_40625,N_39949,N_39696);
and U40626 (N_40626,N_39974,N_39674);
nor U40627 (N_40627,N_39805,N_39557);
nor U40628 (N_40628,N_39335,N_39948);
xor U40629 (N_40629,N_39863,N_39406);
nand U40630 (N_40630,N_39948,N_39502);
nor U40631 (N_40631,N_39019,N_39675);
nor U40632 (N_40632,N_39999,N_39259);
xnor U40633 (N_40633,N_39548,N_39540);
xnor U40634 (N_40634,N_39582,N_39650);
nor U40635 (N_40635,N_39679,N_39391);
and U40636 (N_40636,N_39999,N_39398);
nand U40637 (N_40637,N_39373,N_39566);
and U40638 (N_40638,N_39644,N_39394);
and U40639 (N_40639,N_39470,N_39774);
xor U40640 (N_40640,N_39268,N_39127);
nand U40641 (N_40641,N_39719,N_39751);
and U40642 (N_40642,N_39068,N_39365);
or U40643 (N_40643,N_39467,N_39413);
nand U40644 (N_40644,N_39970,N_39582);
or U40645 (N_40645,N_39593,N_39697);
nand U40646 (N_40646,N_39025,N_39380);
xnor U40647 (N_40647,N_39327,N_39538);
or U40648 (N_40648,N_39041,N_39076);
and U40649 (N_40649,N_39187,N_39196);
nand U40650 (N_40650,N_39437,N_39564);
nand U40651 (N_40651,N_39938,N_39535);
xnor U40652 (N_40652,N_39637,N_39084);
or U40653 (N_40653,N_39325,N_39397);
nor U40654 (N_40654,N_39411,N_39336);
nor U40655 (N_40655,N_39370,N_39827);
nand U40656 (N_40656,N_39342,N_39648);
nand U40657 (N_40657,N_39989,N_39745);
xnor U40658 (N_40658,N_39168,N_39649);
nand U40659 (N_40659,N_39571,N_39758);
and U40660 (N_40660,N_39476,N_39311);
xnor U40661 (N_40661,N_39652,N_39825);
nor U40662 (N_40662,N_39540,N_39272);
and U40663 (N_40663,N_39279,N_39566);
nor U40664 (N_40664,N_39839,N_39015);
xor U40665 (N_40665,N_39685,N_39580);
nor U40666 (N_40666,N_39045,N_39714);
and U40667 (N_40667,N_39178,N_39530);
and U40668 (N_40668,N_39640,N_39549);
nor U40669 (N_40669,N_39609,N_39673);
nand U40670 (N_40670,N_39983,N_39297);
xor U40671 (N_40671,N_39277,N_39862);
xor U40672 (N_40672,N_39115,N_39287);
nand U40673 (N_40673,N_39084,N_39319);
or U40674 (N_40674,N_39283,N_39015);
and U40675 (N_40675,N_39930,N_39887);
xnor U40676 (N_40676,N_39724,N_39125);
and U40677 (N_40677,N_39314,N_39239);
or U40678 (N_40678,N_39463,N_39587);
nor U40679 (N_40679,N_39316,N_39685);
nor U40680 (N_40680,N_39012,N_39764);
nand U40681 (N_40681,N_39285,N_39314);
and U40682 (N_40682,N_39153,N_39814);
nand U40683 (N_40683,N_39271,N_39353);
nand U40684 (N_40684,N_39870,N_39230);
nor U40685 (N_40685,N_39642,N_39371);
or U40686 (N_40686,N_39741,N_39077);
xor U40687 (N_40687,N_39737,N_39109);
and U40688 (N_40688,N_39778,N_39575);
nor U40689 (N_40689,N_39390,N_39002);
and U40690 (N_40690,N_39319,N_39297);
or U40691 (N_40691,N_39345,N_39913);
and U40692 (N_40692,N_39517,N_39472);
or U40693 (N_40693,N_39369,N_39235);
and U40694 (N_40694,N_39054,N_39033);
nand U40695 (N_40695,N_39064,N_39757);
or U40696 (N_40696,N_39925,N_39962);
nor U40697 (N_40697,N_39770,N_39351);
nand U40698 (N_40698,N_39681,N_39043);
nor U40699 (N_40699,N_39668,N_39927);
nand U40700 (N_40700,N_39501,N_39952);
xor U40701 (N_40701,N_39002,N_39196);
and U40702 (N_40702,N_39141,N_39595);
nand U40703 (N_40703,N_39637,N_39909);
or U40704 (N_40704,N_39428,N_39268);
nand U40705 (N_40705,N_39215,N_39033);
nand U40706 (N_40706,N_39773,N_39108);
and U40707 (N_40707,N_39962,N_39062);
nand U40708 (N_40708,N_39352,N_39357);
or U40709 (N_40709,N_39070,N_39051);
and U40710 (N_40710,N_39786,N_39755);
nor U40711 (N_40711,N_39923,N_39715);
nand U40712 (N_40712,N_39000,N_39684);
nor U40713 (N_40713,N_39098,N_39213);
or U40714 (N_40714,N_39979,N_39107);
or U40715 (N_40715,N_39262,N_39427);
or U40716 (N_40716,N_39133,N_39981);
xnor U40717 (N_40717,N_39284,N_39839);
nor U40718 (N_40718,N_39410,N_39804);
nand U40719 (N_40719,N_39121,N_39032);
xor U40720 (N_40720,N_39511,N_39282);
or U40721 (N_40721,N_39956,N_39068);
or U40722 (N_40722,N_39837,N_39559);
nand U40723 (N_40723,N_39311,N_39671);
and U40724 (N_40724,N_39377,N_39281);
and U40725 (N_40725,N_39917,N_39193);
nand U40726 (N_40726,N_39712,N_39440);
nand U40727 (N_40727,N_39279,N_39781);
and U40728 (N_40728,N_39249,N_39382);
nand U40729 (N_40729,N_39296,N_39363);
nor U40730 (N_40730,N_39154,N_39131);
nand U40731 (N_40731,N_39936,N_39048);
xor U40732 (N_40732,N_39997,N_39592);
or U40733 (N_40733,N_39209,N_39758);
nor U40734 (N_40734,N_39401,N_39984);
xor U40735 (N_40735,N_39754,N_39808);
xor U40736 (N_40736,N_39437,N_39459);
nand U40737 (N_40737,N_39738,N_39081);
nand U40738 (N_40738,N_39362,N_39583);
xnor U40739 (N_40739,N_39162,N_39133);
nor U40740 (N_40740,N_39347,N_39291);
xor U40741 (N_40741,N_39066,N_39058);
xnor U40742 (N_40742,N_39885,N_39005);
and U40743 (N_40743,N_39057,N_39247);
or U40744 (N_40744,N_39536,N_39644);
and U40745 (N_40745,N_39287,N_39007);
nand U40746 (N_40746,N_39099,N_39888);
nand U40747 (N_40747,N_39746,N_39871);
xnor U40748 (N_40748,N_39155,N_39259);
and U40749 (N_40749,N_39103,N_39567);
and U40750 (N_40750,N_39341,N_39038);
nand U40751 (N_40751,N_39670,N_39189);
nor U40752 (N_40752,N_39810,N_39084);
nor U40753 (N_40753,N_39917,N_39001);
or U40754 (N_40754,N_39810,N_39103);
and U40755 (N_40755,N_39988,N_39419);
nand U40756 (N_40756,N_39219,N_39100);
nor U40757 (N_40757,N_39474,N_39322);
nor U40758 (N_40758,N_39339,N_39177);
xnor U40759 (N_40759,N_39726,N_39459);
and U40760 (N_40760,N_39487,N_39418);
nand U40761 (N_40761,N_39018,N_39698);
xor U40762 (N_40762,N_39559,N_39470);
or U40763 (N_40763,N_39879,N_39938);
or U40764 (N_40764,N_39204,N_39759);
xor U40765 (N_40765,N_39936,N_39766);
nand U40766 (N_40766,N_39630,N_39996);
xnor U40767 (N_40767,N_39969,N_39881);
and U40768 (N_40768,N_39453,N_39482);
nand U40769 (N_40769,N_39823,N_39575);
nor U40770 (N_40770,N_39549,N_39258);
and U40771 (N_40771,N_39985,N_39059);
and U40772 (N_40772,N_39421,N_39870);
and U40773 (N_40773,N_39896,N_39101);
or U40774 (N_40774,N_39750,N_39901);
nor U40775 (N_40775,N_39066,N_39049);
or U40776 (N_40776,N_39098,N_39543);
nand U40777 (N_40777,N_39097,N_39433);
and U40778 (N_40778,N_39687,N_39801);
xnor U40779 (N_40779,N_39522,N_39364);
or U40780 (N_40780,N_39710,N_39095);
or U40781 (N_40781,N_39698,N_39758);
nor U40782 (N_40782,N_39996,N_39537);
xnor U40783 (N_40783,N_39798,N_39734);
xnor U40784 (N_40784,N_39621,N_39803);
xor U40785 (N_40785,N_39576,N_39443);
nand U40786 (N_40786,N_39344,N_39389);
and U40787 (N_40787,N_39656,N_39463);
nor U40788 (N_40788,N_39687,N_39065);
or U40789 (N_40789,N_39117,N_39451);
nand U40790 (N_40790,N_39373,N_39659);
and U40791 (N_40791,N_39503,N_39217);
xor U40792 (N_40792,N_39018,N_39537);
nor U40793 (N_40793,N_39412,N_39275);
and U40794 (N_40794,N_39564,N_39294);
and U40795 (N_40795,N_39265,N_39007);
or U40796 (N_40796,N_39330,N_39548);
or U40797 (N_40797,N_39514,N_39216);
nand U40798 (N_40798,N_39324,N_39204);
nor U40799 (N_40799,N_39179,N_39933);
or U40800 (N_40800,N_39622,N_39288);
xor U40801 (N_40801,N_39481,N_39062);
nand U40802 (N_40802,N_39038,N_39795);
nor U40803 (N_40803,N_39459,N_39324);
nand U40804 (N_40804,N_39725,N_39306);
and U40805 (N_40805,N_39590,N_39051);
or U40806 (N_40806,N_39139,N_39281);
or U40807 (N_40807,N_39524,N_39363);
or U40808 (N_40808,N_39364,N_39042);
xnor U40809 (N_40809,N_39667,N_39618);
and U40810 (N_40810,N_39429,N_39817);
xnor U40811 (N_40811,N_39848,N_39049);
nand U40812 (N_40812,N_39860,N_39097);
nor U40813 (N_40813,N_39639,N_39486);
or U40814 (N_40814,N_39894,N_39913);
or U40815 (N_40815,N_39407,N_39125);
and U40816 (N_40816,N_39966,N_39257);
xor U40817 (N_40817,N_39915,N_39687);
or U40818 (N_40818,N_39259,N_39158);
nor U40819 (N_40819,N_39881,N_39156);
or U40820 (N_40820,N_39746,N_39607);
nor U40821 (N_40821,N_39414,N_39206);
xnor U40822 (N_40822,N_39748,N_39281);
and U40823 (N_40823,N_39595,N_39429);
nand U40824 (N_40824,N_39473,N_39030);
xor U40825 (N_40825,N_39049,N_39575);
xnor U40826 (N_40826,N_39162,N_39100);
and U40827 (N_40827,N_39361,N_39748);
nor U40828 (N_40828,N_39069,N_39849);
xor U40829 (N_40829,N_39753,N_39283);
and U40830 (N_40830,N_39211,N_39814);
nand U40831 (N_40831,N_39422,N_39519);
or U40832 (N_40832,N_39536,N_39343);
or U40833 (N_40833,N_39114,N_39600);
and U40834 (N_40834,N_39209,N_39075);
xnor U40835 (N_40835,N_39678,N_39486);
and U40836 (N_40836,N_39772,N_39909);
or U40837 (N_40837,N_39238,N_39449);
xor U40838 (N_40838,N_39207,N_39440);
nor U40839 (N_40839,N_39539,N_39132);
xor U40840 (N_40840,N_39234,N_39763);
or U40841 (N_40841,N_39022,N_39055);
xor U40842 (N_40842,N_39824,N_39149);
nand U40843 (N_40843,N_39121,N_39970);
nand U40844 (N_40844,N_39017,N_39427);
nor U40845 (N_40845,N_39850,N_39989);
and U40846 (N_40846,N_39273,N_39904);
xnor U40847 (N_40847,N_39445,N_39327);
nor U40848 (N_40848,N_39938,N_39105);
and U40849 (N_40849,N_39600,N_39516);
or U40850 (N_40850,N_39472,N_39745);
nand U40851 (N_40851,N_39054,N_39060);
nor U40852 (N_40852,N_39526,N_39313);
xnor U40853 (N_40853,N_39706,N_39879);
nand U40854 (N_40854,N_39535,N_39861);
nor U40855 (N_40855,N_39159,N_39126);
nor U40856 (N_40856,N_39278,N_39833);
nand U40857 (N_40857,N_39201,N_39962);
xor U40858 (N_40858,N_39417,N_39934);
and U40859 (N_40859,N_39309,N_39866);
nand U40860 (N_40860,N_39511,N_39085);
and U40861 (N_40861,N_39732,N_39041);
nand U40862 (N_40862,N_39460,N_39408);
nor U40863 (N_40863,N_39056,N_39097);
xnor U40864 (N_40864,N_39792,N_39225);
or U40865 (N_40865,N_39613,N_39122);
nor U40866 (N_40866,N_39709,N_39894);
xnor U40867 (N_40867,N_39679,N_39263);
nor U40868 (N_40868,N_39488,N_39072);
nand U40869 (N_40869,N_39897,N_39383);
or U40870 (N_40870,N_39945,N_39633);
or U40871 (N_40871,N_39907,N_39745);
nand U40872 (N_40872,N_39402,N_39028);
nor U40873 (N_40873,N_39361,N_39863);
nor U40874 (N_40874,N_39607,N_39097);
or U40875 (N_40875,N_39012,N_39051);
or U40876 (N_40876,N_39444,N_39546);
nor U40877 (N_40877,N_39979,N_39805);
and U40878 (N_40878,N_39839,N_39381);
xor U40879 (N_40879,N_39303,N_39683);
nor U40880 (N_40880,N_39973,N_39703);
or U40881 (N_40881,N_39128,N_39195);
and U40882 (N_40882,N_39069,N_39938);
xnor U40883 (N_40883,N_39753,N_39710);
nand U40884 (N_40884,N_39550,N_39869);
or U40885 (N_40885,N_39486,N_39535);
or U40886 (N_40886,N_39935,N_39598);
nor U40887 (N_40887,N_39067,N_39272);
and U40888 (N_40888,N_39011,N_39351);
or U40889 (N_40889,N_39143,N_39058);
nor U40890 (N_40890,N_39084,N_39115);
nor U40891 (N_40891,N_39396,N_39128);
nor U40892 (N_40892,N_39039,N_39282);
nor U40893 (N_40893,N_39421,N_39335);
xor U40894 (N_40894,N_39700,N_39145);
nor U40895 (N_40895,N_39984,N_39894);
or U40896 (N_40896,N_39371,N_39558);
nor U40897 (N_40897,N_39706,N_39571);
or U40898 (N_40898,N_39507,N_39920);
or U40899 (N_40899,N_39581,N_39544);
nor U40900 (N_40900,N_39629,N_39660);
and U40901 (N_40901,N_39689,N_39640);
xor U40902 (N_40902,N_39703,N_39459);
or U40903 (N_40903,N_39871,N_39427);
nand U40904 (N_40904,N_39510,N_39245);
or U40905 (N_40905,N_39836,N_39057);
or U40906 (N_40906,N_39850,N_39118);
nor U40907 (N_40907,N_39045,N_39375);
nand U40908 (N_40908,N_39700,N_39676);
xor U40909 (N_40909,N_39161,N_39105);
nor U40910 (N_40910,N_39193,N_39566);
or U40911 (N_40911,N_39206,N_39928);
nor U40912 (N_40912,N_39483,N_39645);
xor U40913 (N_40913,N_39962,N_39705);
or U40914 (N_40914,N_39859,N_39549);
nor U40915 (N_40915,N_39066,N_39138);
or U40916 (N_40916,N_39404,N_39499);
nor U40917 (N_40917,N_39759,N_39556);
xor U40918 (N_40918,N_39199,N_39487);
or U40919 (N_40919,N_39289,N_39246);
and U40920 (N_40920,N_39750,N_39727);
xor U40921 (N_40921,N_39014,N_39086);
xor U40922 (N_40922,N_39446,N_39144);
or U40923 (N_40923,N_39569,N_39496);
nand U40924 (N_40924,N_39209,N_39018);
or U40925 (N_40925,N_39999,N_39988);
xnor U40926 (N_40926,N_39333,N_39933);
xor U40927 (N_40927,N_39610,N_39679);
nand U40928 (N_40928,N_39812,N_39921);
nand U40929 (N_40929,N_39173,N_39077);
nand U40930 (N_40930,N_39361,N_39724);
and U40931 (N_40931,N_39350,N_39028);
and U40932 (N_40932,N_39576,N_39816);
nor U40933 (N_40933,N_39159,N_39117);
nor U40934 (N_40934,N_39585,N_39498);
nor U40935 (N_40935,N_39978,N_39708);
and U40936 (N_40936,N_39160,N_39088);
or U40937 (N_40937,N_39295,N_39027);
xor U40938 (N_40938,N_39672,N_39214);
xor U40939 (N_40939,N_39252,N_39151);
nand U40940 (N_40940,N_39705,N_39141);
xor U40941 (N_40941,N_39930,N_39173);
nand U40942 (N_40942,N_39027,N_39583);
nand U40943 (N_40943,N_39408,N_39280);
or U40944 (N_40944,N_39460,N_39700);
xor U40945 (N_40945,N_39133,N_39141);
and U40946 (N_40946,N_39590,N_39904);
and U40947 (N_40947,N_39097,N_39713);
or U40948 (N_40948,N_39592,N_39832);
nand U40949 (N_40949,N_39711,N_39333);
nand U40950 (N_40950,N_39292,N_39906);
and U40951 (N_40951,N_39195,N_39427);
nor U40952 (N_40952,N_39400,N_39240);
nand U40953 (N_40953,N_39721,N_39073);
nor U40954 (N_40954,N_39043,N_39477);
nor U40955 (N_40955,N_39411,N_39878);
and U40956 (N_40956,N_39613,N_39912);
nand U40957 (N_40957,N_39878,N_39708);
nor U40958 (N_40958,N_39972,N_39434);
and U40959 (N_40959,N_39385,N_39776);
xor U40960 (N_40960,N_39913,N_39202);
nand U40961 (N_40961,N_39720,N_39481);
or U40962 (N_40962,N_39044,N_39930);
nor U40963 (N_40963,N_39767,N_39074);
xor U40964 (N_40964,N_39530,N_39926);
or U40965 (N_40965,N_39930,N_39978);
xor U40966 (N_40966,N_39025,N_39281);
xnor U40967 (N_40967,N_39767,N_39942);
nor U40968 (N_40968,N_39968,N_39599);
or U40969 (N_40969,N_39385,N_39587);
nand U40970 (N_40970,N_39948,N_39124);
and U40971 (N_40971,N_39549,N_39118);
or U40972 (N_40972,N_39510,N_39933);
and U40973 (N_40973,N_39409,N_39497);
or U40974 (N_40974,N_39868,N_39851);
and U40975 (N_40975,N_39307,N_39756);
xor U40976 (N_40976,N_39359,N_39485);
xor U40977 (N_40977,N_39693,N_39325);
xnor U40978 (N_40978,N_39655,N_39102);
nand U40979 (N_40979,N_39620,N_39616);
nor U40980 (N_40980,N_39163,N_39400);
nand U40981 (N_40981,N_39470,N_39793);
and U40982 (N_40982,N_39938,N_39010);
nor U40983 (N_40983,N_39543,N_39009);
and U40984 (N_40984,N_39228,N_39472);
nand U40985 (N_40985,N_39739,N_39408);
xnor U40986 (N_40986,N_39664,N_39336);
and U40987 (N_40987,N_39329,N_39014);
nand U40988 (N_40988,N_39058,N_39256);
and U40989 (N_40989,N_39259,N_39852);
or U40990 (N_40990,N_39721,N_39848);
xor U40991 (N_40991,N_39211,N_39447);
or U40992 (N_40992,N_39467,N_39485);
and U40993 (N_40993,N_39453,N_39712);
nand U40994 (N_40994,N_39827,N_39470);
and U40995 (N_40995,N_39911,N_39378);
xnor U40996 (N_40996,N_39403,N_39784);
or U40997 (N_40997,N_39195,N_39550);
nand U40998 (N_40998,N_39800,N_39981);
nor U40999 (N_40999,N_39125,N_39456);
nor U41000 (N_41000,N_40082,N_40285);
xnor U41001 (N_41001,N_40958,N_40736);
nor U41002 (N_41002,N_40591,N_40734);
and U41003 (N_41003,N_40050,N_40257);
or U41004 (N_41004,N_40998,N_40897);
nand U41005 (N_41005,N_40858,N_40363);
or U41006 (N_41006,N_40777,N_40494);
and U41007 (N_41007,N_40551,N_40772);
nand U41008 (N_41008,N_40864,N_40417);
nand U41009 (N_41009,N_40751,N_40236);
nand U41010 (N_41010,N_40240,N_40879);
and U41011 (N_41011,N_40126,N_40439);
or U41012 (N_41012,N_40112,N_40818);
nor U41013 (N_41013,N_40607,N_40606);
or U41014 (N_41014,N_40825,N_40183);
nand U41015 (N_41015,N_40553,N_40048);
or U41016 (N_41016,N_40447,N_40182);
and U41017 (N_41017,N_40326,N_40731);
or U41018 (N_41018,N_40654,N_40749);
and U41019 (N_41019,N_40881,N_40402);
or U41020 (N_41020,N_40484,N_40910);
nand U41021 (N_41021,N_40718,N_40332);
and U41022 (N_41022,N_40700,N_40632);
and U41023 (N_41023,N_40275,N_40918);
or U41024 (N_41024,N_40692,N_40672);
nor U41025 (N_41025,N_40199,N_40260);
and U41026 (N_41026,N_40284,N_40537);
and U41027 (N_41027,N_40250,N_40265);
xor U41028 (N_41028,N_40656,N_40255);
nand U41029 (N_41029,N_40440,N_40811);
nor U41030 (N_41030,N_40624,N_40648);
nand U41031 (N_41031,N_40241,N_40015);
nand U41032 (N_41032,N_40376,N_40037);
and U41033 (N_41033,N_40391,N_40878);
xnor U41034 (N_41034,N_40708,N_40165);
nand U41035 (N_41035,N_40456,N_40572);
or U41036 (N_41036,N_40324,N_40486);
or U41037 (N_41037,N_40630,N_40667);
xnor U41038 (N_41038,N_40721,N_40244);
nand U41039 (N_41039,N_40857,N_40823);
or U41040 (N_41040,N_40095,N_40690);
xor U41041 (N_41041,N_40438,N_40931);
and U41042 (N_41042,N_40807,N_40173);
nor U41043 (N_41043,N_40849,N_40306);
nor U41044 (N_41044,N_40441,N_40990);
or U41045 (N_41045,N_40780,N_40481);
or U41046 (N_41046,N_40058,N_40688);
or U41047 (N_41047,N_40033,N_40418);
nor U41048 (N_41048,N_40345,N_40600);
nor U41049 (N_41049,N_40270,N_40188);
and U41050 (N_41050,N_40365,N_40548);
nand U41051 (N_41051,N_40406,N_40530);
nor U41052 (N_41052,N_40087,N_40121);
and U41053 (N_41053,N_40571,N_40940);
nor U41054 (N_41054,N_40018,N_40791);
or U41055 (N_41055,N_40171,N_40198);
xnor U41056 (N_41056,N_40576,N_40492);
nand U41057 (N_41057,N_40827,N_40601);
xor U41058 (N_41058,N_40951,N_40725);
nand U41059 (N_41059,N_40068,N_40505);
xnor U41060 (N_41060,N_40894,N_40097);
and U41061 (N_41061,N_40153,N_40853);
nor U41062 (N_41062,N_40582,N_40099);
nand U41063 (N_41063,N_40869,N_40666);
nor U41064 (N_41064,N_40542,N_40681);
nand U41065 (N_41065,N_40683,N_40920);
nand U41066 (N_41066,N_40806,N_40761);
xnor U41067 (N_41067,N_40249,N_40215);
or U41068 (N_41068,N_40549,N_40522);
nor U41069 (N_41069,N_40049,N_40384);
and U41070 (N_41070,N_40541,N_40320);
xor U41071 (N_41071,N_40676,N_40006);
nand U41072 (N_41072,N_40730,N_40679);
nor U41073 (N_41073,N_40615,N_40354);
nand U41074 (N_41074,N_40014,N_40637);
xor U41075 (N_41075,N_40580,N_40403);
nand U41076 (N_41076,N_40593,N_40740);
and U41077 (N_41077,N_40955,N_40562);
nor U41078 (N_41078,N_40538,N_40273);
and U41079 (N_41079,N_40358,N_40883);
or U41080 (N_41080,N_40079,N_40638);
nand U41081 (N_41081,N_40525,N_40093);
and U41082 (N_41082,N_40642,N_40355);
and U41083 (N_41083,N_40297,N_40797);
nand U41084 (N_41084,N_40763,N_40178);
or U41085 (N_41085,N_40616,N_40599);
and U41086 (N_41086,N_40206,N_40259);
nand U41087 (N_41087,N_40875,N_40096);
nand U41088 (N_41088,N_40308,N_40929);
nor U41089 (N_41089,N_40794,N_40474);
nor U41090 (N_41090,N_40115,N_40063);
and U41091 (N_41091,N_40392,N_40620);
nor U41092 (N_41092,N_40043,N_40304);
nor U41093 (N_41093,N_40557,N_40129);
nor U41094 (N_41094,N_40733,N_40532);
and U41095 (N_41095,N_40922,N_40911);
nand U41096 (N_41096,N_40127,N_40816);
or U41097 (N_41097,N_40561,N_40021);
xor U41098 (N_41098,N_40135,N_40521);
nor U41099 (N_41099,N_40221,N_40437);
and U41100 (N_41100,N_40975,N_40661);
and U41101 (N_41101,N_40458,N_40223);
xor U41102 (N_41102,N_40871,N_40231);
and U41103 (N_41103,N_40983,N_40070);
xor U41104 (N_41104,N_40232,N_40469);
nor U41105 (N_41105,N_40578,N_40060);
nor U41106 (N_41106,N_40674,N_40042);
nand U41107 (N_41107,N_40841,N_40077);
or U41108 (N_41108,N_40934,N_40116);
xnor U41109 (N_41109,N_40776,N_40587);
and U41110 (N_41110,N_40832,N_40076);
xor U41111 (N_41111,N_40109,N_40432);
and U41112 (N_41112,N_40067,N_40737);
nor U41113 (N_41113,N_40602,N_40640);
xnor U41114 (N_41114,N_40583,N_40919);
nor U41115 (N_41115,N_40010,N_40985);
xnor U41116 (N_41116,N_40820,N_40787);
or U41117 (N_41117,N_40194,N_40248);
nor U41118 (N_41118,N_40367,N_40208);
nor U41119 (N_41119,N_40274,N_40298);
xnor U41120 (N_41120,N_40810,N_40765);
xnor U41121 (N_41121,N_40086,N_40888);
nand U41122 (N_41122,N_40992,N_40565);
nor U41123 (N_41123,N_40370,N_40344);
xnor U41124 (N_41124,N_40608,N_40670);
or U41125 (N_41125,N_40146,N_40817);
or U41126 (N_41126,N_40848,N_40967);
or U41127 (N_41127,N_40125,N_40426);
xnor U41128 (N_41128,N_40533,N_40137);
and U41129 (N_41129,N_40999,N_40907);
xnor U41130 (N_41130,N_40352,N_40547);
or U41131 (N_41131,N_40094,N_40760);
nand U41132 (N_41132,N_40479,N_40891);
and U41133 (N_41133,N_40176,N_40472);
nor U41134 (N_41134,N_40979,N_40162);
and U41135 (N_41135,N_40812,N_40696);
nand U41136 (N_41136,N_40187,N_40768);
and U41137 (N_41137,N_40246,N_40263);
or U41138 (N_41138,N_40313,N_40405);
nor U41139 (N_41139,N_40005,N_40477);
nor U41140 (N_41140,N_40655,N_40483);
or U41141 (N_41141,N_40108,N_40793);
and U41142 (N_41142,N_40673,N_40660);
nor U41143 (N_41143,N_40353,N_40658);
nor U41144 (N_41144,N_40711,N_40379);
nor U41145 (N_41145,N_40467,N_40119);
nor U41146 (N_41146,N_40166,N_40824);
or U41147 (N_41147,N_40963,N_40289);
nor U41148 (N_41148,N_40210,N_40154);
and U41149 (N_41149,N_40161,N_40719);
xnor U41150 (N_41150,N_40948,N_40366);
nand U41151 (N_41151,N_40829,N_40536);
nand U41152 (N_41152,N_40909,N_40444);
xnor U41153 (N_41153,N_40335,N_40327);
nor U41154 (N_41154,N_40359,N_40429);
and U41155 (N_41155,N_40603,N_40933);
and U41156 (N_41156,N_40083,N_40938);
or U41157 (N_41157,N_40585,N_40433);
and U41158 (N_41158,N_40779,N_40895);
nand U41159 (N_41159,N_40588,N_40974);
or U41160 (N_41160,N_40570,N_40579);
and U41161 (N_41161,N_40527,N_40105);
or U41162 (N_41162,N_40464,N_40380);
and U41163 (N_41163,N_40431,N_40942);
nand U41164 (N_41164,N_40502,N_40993);
nand U41165 (N_41165,N_40148,N_40267);
xor U41166 (N_41166,N_40051,N_40266);
xor U41167 (N_41167,N_40678,N_40937);
or U41168 (N_41168,N_40026,N_40446);
or U41169 (N_41169,N_40234,N_40283);
and U41170 (N_41170,N_40128,N_40168);
xnor U41171 (N_41171,N_40949,N_40921);
and U41172 (N_41172,N_40971,N_40722);
or U41173 (N_41173,N_40987,N_40253);
and U41174 (N_41174,N_40214,N_40061);
nand U41175 (N_41175,N_40716,N_40511);
nand U41176 (N_41176,N_40174,N_40185);
and U41177 (N_41177,N_40350,N_40509);
or U41178 (N_41178,N_40717,N_40381);
nor U41179 (N_41179,N_40302,N_40752);
xor U41180 (N_41180,N_40926,N_40118);
nand U41181 (N_41181,N_40321,N_40150);
xnor U41182 (N_41182,N_40643,N_40027);
or U41183 (N_41183,N_40568,N_40314);
nor U41184 (N_41184,N_40212,N_40695);
or U41185 (N_41185,N_40802,N_40045);
nand U41186 (N_41186,N_40664,N_40325);
or U41187 (N_41187,N_40633,N_40575);
xnor U41188 (N_41188,N_40924,N_40743);
or U41189 (N_41189,N_40550,N_40790);
and U41190 (N_41190,N_40268,N_40395);
and U41191 (N_41191,N_40339,N_40139);
and U41192 (N_41192,N_40629,N_40651);
nand U41193 (N_41193,N_40745,N_40342);
and U41194 (N_41194,N_40281,N_40254);
xor U41195 (N_41195,N_40517,N_40855);
nand U41196 (N_41196,N_40396,N_40997);
nand U41197 (N_41197,N_40338,N_40706);
nand U41198 (N_41198,N_40104,N_40282);
or U41199 (N_41199,N_40235,N_40497);
and U41200 (N_41200,N_40216,N_40053);
nand U41201 (N_41201,N_40175,N_40362);
or U41202 (N_41202,N_40555,N_40621);
or U41203 (N_41203,N_40594,N_40300);
xnor U41204 (N_41204,N_40224,N_40543);
nor U41205 (N_41205,N_40969,N_40710);
or U41206 (N_41206,N_40876,N_40767);
nor U41207 (N_41207,N_40896,N_40506);
nor U41208 (N_41208,N_40619,N_40330);
and U41209 (N_41209,N_40647,N_40778);
or U41210 (N_41210,N_40455,N_40170);
nand U41211 (N_41211,N_40288,N_40230);
nor U41212 (N_41212,N_40310,N_40377);
xor U41213 (N_41213,N_40155,N_40276);
nor U41214 (N_41214,N_40754,N_40930);
or U41215 (N_41215,N_40668,N_40197);
nor U41216 (N_41216,N_40833,N_40687);
nor U41217 (N_41217,N_40556,N_40465);
nand U41218 (N_41218,N_40085,N_40982);
xor U41219 (N_41219,N_40540,N_40613);
and U41220 (N_41220,N_40928,N_40203);
xnor U41221 (N_41221,N_40419,N_40775);
and U41222 (N_41222,N_40393,N_40389);
nor U41223 (N_41223,N_40387,N_40813);
xnor U41224 (N_41224,N_40205,N_40084);
nor U41225 (N_41225,N_40445,N_40074);
nand U41226 (N_41226,N_40184,N_40322);
nand U41227 (N_41227,N_40346,N_40880);
xnor U41228 (N_41228,N_40507,N_40073);
xnor U41229 (N_41229,N_40410,N_40177);
and U41230 (N_41230,N_40623,N_40892);
and U41231 (N_41231,N_40424,N_40336);
and U41232 (N_41232,N_40172,N_40480);
xor U41233 (N_41233,N_40500,N_40762);
or U41234 (N_41234,N_40685,N_40493);
and U41235 (N_41235,N_40054,N_40757);
nor U41236 (N_41236,N_40586,N_40329);
nand U41237 (N_41237,N_40792,N_40657);
xor U41238 (N_41238,N_40834,N_40461);
xnor U41239 (N_41239,N_40133,N_40916);
or U41240 (N_41240,N_40519,N_40986);
or U41241 (N_41241,N_40596,N_40013);
xor U41242 (N_41242,N_40645,N_40913);
nand U41243 (N_41243,N_40914,N_40499);
or U41244 (N_41244,N_40059,N_40031);
and U41245 (N_41245,N_40195,N_40134);
xnor U41246 (N_41246,N_40341,N_40373);
xnor U41247 (N_41247,N_40022,N_40167);
and U41248 (N_41248,N_40451,N_40644);
nor U41249 (N_41249,N_40625,N_40808);
nand U41250 (N_41250,N_40251,N_40627);
nor U41251 (N_41251,N_40147,N_40663);
nand U41252 (N_41252,N_40866,N_40753);
or U41253 (N_41253,N_40123,N_40835);
or U41254 (N_41254,N_40091,N_40039);
xor U41255 (N_41255,N_40628,N_40783);
and U41256 (N_41256,N_40652,N_40498);
or U41257 (N_41257,N_40523,N_40140);
nor U41258 (N_41258,N_40795,N_40219);
nor U41259 (N_41259,N_40434,N_40905);
and U41260 (N_41260,N_40798,N_40747);
nor U41261 (N_41261,N_40893,N_40901);
nor U41262 (N_41262,N_40293,N_40066);
nor U41263 (N_41263,N_40524,N_40741);
xor U41264 (N_41264,N_40520,N_40636);
nor U41265 (N_41265,N_40025,N_40028);
nand U41266 (N_41266,N_40351,N_40544);
nor U41267 (N_41267,N_40252,N_40965);
or U41268 (N_41268,N_40292,N_40149);
nand U41269 (N_41269,N_40796,N_40279);
and U41270 (N_41270,N_40694,N_40904);
and U41271 (N_41271,N_40945,N_40296);
xor U41272 (N_41272,N_40229,N_40756);
nand U41273 (N_41273,N_40781,N_40732);
xnor U41274 (N_41274,N_40641,N_40539);
and U41275 (N_41275,N_40152,N_40689);
and U41276 (N_41276,N_40269,N_40390);
nand U41277 (N_41277,N_40944,N_40144);
xor U41278 (N_41278,N_40407,N_40114);
or U41279 (N_41279,N_40181,N_40072);
nand U41280 (N_41280,N_40960,N_40805);
and U41281 (N_41281,N_40495,N_40041);
xor U41282 (N_41282,N_40131,N_40038);
or U41283 (N_41283,N_40449,N_40882);
or U41284 (N_41284,N_40157,N_40782);
xor U41285 (N_41285,N_40192,N_40766);
and U41286 (N_41286,N_40868,N_40845);
nor U41287 (N_41287,N_40699,N_40132);
xnor U41288 (N_41288,N_40515,N_40744);
nor U41289 (N_41289,N_40707,N_40017);
xnor U41290 (N_41290,N_40785,N_40057);
and U41291 (N_41291,N_40592,N_40428);
nor U41292 (N_41292,N_40436,N_40473);
nand U41293 (N_41293,N_40081,N_40190);
xor U41294 (N_41294,N_40397,N_40264);
nor U41295 (N_41295,N_40245,N_40156);
or U41296 (N_41296,N_40563,N_40755);
and U41297 (N_41297,N_40315,N_40906);
nand U41298 (N_41298,N_40145,N_40023);
nand U41299 (N_41299,N_40340,N_40122);
and U41300 (N_41300,N_40902,N_40090);
or U41301 (N_41301,N_40925,N_40200);
or U41302 (N_41302,N_40416,N_40008);
and U41303 (N_41303,N_40318,N_40489);
nand U41304 (N_41304,N_40598,N_40243);
xor U41305 (N_41305,N_40052,N_40605);
or U41306 (N_41306,N_40334,N_40080);
nor U41307 (N_41307,N_40225,N_40294);
xor U41308 (N_41308,N_40107,N_40671);
nand U41309 (N_41309,N_40317,N_40004);
and U41310 (N_41310,N_40742,N_40261);
and U41311 (N_41311,N_40784,N_40972);
and U41312 (N_41312,N_40287,N_40138);
nand U41313 (N_41313,N_40475,N_40226);
and U41314 (N_41314,N_40814,N_40801);
nor U41315 (N_41315,N_40650,N_40062);
nor U41316 (N_41316,N_40535,N_40899);
nand U41317 (N_41317,N_40078,N_40724);
or U41318 (N_41318,N_40356,N_40847);
xnor U41319 (N_41319,N_40941,N_40682);
nor U41320 (N_41320,N_40189,N_40295);
or U41321 (N_41321,N_40452,N_40398);
and U41322 (N_41322,N_40516,N_40774);
nor U41323 (N_41323,N_40211,N_40799);
xnor U41324 (N_41324,N_40485,N_40610);
nand U41325 (N_41325,N_40531,N_40204);
and U41326 (N_41326,N_40691,N_40915);
xnor U41327 (N_41327,N_40697,N_40482);
xor U41328 (N_41328,N_40089,N_40003);
and U41329 (N_41329,N_40618,N_40030);
xor U41330 (N_41330,N_40343,N_40769);
or U41331 (N_41331,N_40560,N_40712);
nand U41332 (N_41332,N_40512,N_40262);
xor U41333 (N_41333,N_40976,N_40371);
and U41334 (N_41334,N_40337,N_40964);
nor U41335 (N_41335,N_40382,N_40513);
and U41336 (N_41336,N_40994,N_40552);
nand U41337 (N_41337,N_40164,N_40349);
nand U41338 (N_41338,N_40970,N_40316);
or U41339 (N_41339,N_40009,N_40614);
or U41340 (N_41340,N_40202,N_40714);
nand U41341 (N_41341,N_40328,N_40748);
and U41342 (N_41342,N_40545,N_40980);
xor U41343 (N_41343,N_40885,N_40912);
nor U41344 (N_41344,N_40071,N_40856);
nor U41345 (N_41345,N_40374,N_40369);
or U41346 (N_41346,N_40534,N_40846);
nor U41347 (N_41347,N_40256,N_40238);
or U41348 (N_41348,N_40935,N_40388);
or U41349 (N_41349,N_40111,N_40305);
nand U41350 (N_41350,N_40303,N_40786);
and U41351 (N_41351,N_40401,N_40822);
nor U41352 (N_41352,N_40457,N_40375);
or U41353 (N_41353,N_40961,N_40842);
or U41354 (N_41354,N_40491,N_40634);
or U41355 (N_41355,N_40649,N_40011);
or U41356 (N_41356,N_40143,N_40839);
nand U41357 (N_41357,N_40943,N_40988);
or U41358 (N_41358,N_40903,N_40577);
nor U41359 (N_41359,N_40237,N_40514);
xnor U41360 (N_41360,N_40106,N_40946);
or U41361 (N_41361,N_40867,N_40889);
nand U41362 (N_41362,N_40704,N_40981);
and U41363 (N_41363,N_40917,N_40012);
and U41364 (N_41364,N_40597,N_40669);
nor U41365 (N_41365,N_40984,N_40900);
and U41366 (N_41366,N_40415,N_40488);
nand U41367 (N_41367,N_40333,N_40662);
nand U41368 (N_41368,N_40860,N_40877);
and U41369 (N_41369,N_40065,N_40450);
xnor U41370 (N_41370,N_40686,N_40665);
nor U41371 (N_41371,N_40404,N_40510);
xor U41372 (N_41372,N_40954,N_40851);
xnor U41373 (N_41373,N_40047,N_40764);
and U41374 (N_41374,N_40908,N_40454);
nor U41375 (N_41375,N_40639,N_40277);
nand U41376 (N_41376,N_40462,N_40151);
xnor U41377 (N_41377,N_40529,N_40227);
or U41378 (N_41378,N_40258,N_40209);
nand U41379 (N_41379,N_40826,N_40290);
xor U41380 (N_41380,N_40101,N_40968);
and U41381 (N_41381,N_40055,N_40383);
and U41382 (N_41382,N_40991,N_40569);
nand U41383 (N_41383,N_40400,N_40684);
and U41384 (N_41384,N_40421,N_40098);
or U41385 (N_41385,N_40723,N_40069);
nand U41386 (N_41386,N_40361,N_40617);
and U41387 (N_41387,N_40932,N_40311);
and U41388 (N_41388,N_40872,N_40966);
and U41389 (N_41389,N_40564,N_40035);
or U41390 (N_41390,N_40854,N_40466);
or U41391 (N_41391,N_40977,N_40448);
nor U41392 (N_41392,N_40584,N_40959);
or U41393 (N_41393,N_40828,N_40113);
nand U41394 (N_41394,N_40459,N_40193);
or U41395 (N_41395,N_40978,N_40088);
nand U41396 (N_41396,N_40950,N_40709);
and U41397 (N_41397,N_40819,N_40962);
or U41398 (N_41398,N_40136,N_40180);
and U41399 (N_41399,N_40863,N_40307);
and U41400 (N_41400,N_40233,N_40546);
nand U41401 (N_41401,N_40032,N_40413);
or U41402 (N_41402,N_40727,N_40471);
and U41403 (N_41403,N_40423,N_40927);
or U41404 (N_41404,N_40201,N_40442);
nor U41405 (N_41405,N_40836,N_40843);
nand U41406 (N_41406,N_40728,N_40286);
and U41407 (N_41407,N_40635,N_40453);
xnor U41408 (N_41408,N_40228,N_40470);
xor U41409 (N_41409,N_40581,N_40862);
xnor U41410 (N_41410,N_40102,N_40729);
nand U41411 (N_41411,N_40000,N_40715);
and U41412 (N_41412,N_40936,N_40815);
xor U41413 (N_41413,N_40103,N_40773);
nand U41414 (N_41414,N_40859,N_40064);
nor U41415 (N_41415,N_40701,N_40693);
xnor U41416 (N_41416,N_40789,N_40898);
and U41417 (N_41417,N_40476,N_40890);
and U41418 (N_41418,N_40443,N_40220);
and U41419 (N_41419,N_40411,N_40213);
nor U41420 (N_41420,N_40271,N_40110);
or U41421 (N_41421,N_40357,N_40726);
or U41422 (N_41422,N_40278,N_40299);
or U41423 (N_41423,N_40056,N_40364);
and U41424 (N_41424,N_40559,N_40844);
nor U41425 (N_41425,N_40422,N_40414);
nand U41426 (N_41426,N_40957,N_40399);
xor U41427 (N_41427,N_40360,N_40196);
nor U41428 (N_41428,N_40323,N_40850);
or U41429 (N_41429,N_40653,N_40368);
nor U41430 (N_41430,N_40016,N_40750);
xnor U41431 (N_41431,N_40590,N_40738);
nand U41432 (N_41432,N_40567,N_40720);
nand U41433 (N_41433,N_40837,N_40996);
or U41434 (N_41434,N_40120,N_40759);
and U41435 (N_41435,N_40622,N_40372);
and U41436 (N_41436,N_40490,N_40034);
and U41437 (N_41437,N_40046,N_40973);
xnor U41438 (N_41438,N_40141,N_40830);
xnor U41439 (N_41439,N_40508,N_40952);
xnor U41440 (N_41440,N_40040,N_40788);
nor U41441 (N_41441,N_40029,N_40631);
nand U41442 (N_41442,N_40217,N_40840);
nor U41443 (N_41443,N_40409,N_40207);
and U41444 (N_41444,N_40408,N_40558);
nand U41445 (N_41445,N_40412,N_40075);
or U41446 (N_41446,N_40804,N_40478);
and U41447 (N_41447,N_40589,N_40487);
and U41448 (N_41448,N_40394,N_40953);
nand U41449 (N_41449,N_40002,N_40528);
nand U41450 (N_41450,N_40160,N_40609);
or U41451 (N_41451,N_40646,N_40865);
and U41452 (N_41452,N_40705,N_40612);
nor U41453 (N_41453,N_40626,N_40886);
nor U41454 (N_41454,N_40020,N_40703);
or U41455 (N_41455,N_40242,N_40611);
nor U41456 (N_41456,N_40386,N_40809);
nand U41457 (N_41457,N_40378,N_40001);
xnor U41458 (N_41458,N_40874,N_40158);
and U41459 (N_41459,N_40501,N_40771);
and U41460 (N_41460,N_40870,N_40247);
xnor U41461 (N_41461,N_40887,N_40179);
or U41462 (N_41462,N_40130,N_40554);
or U41463 (N_41463,N_40117,N_40319);
and U41464 (N_41464,N_40677,N_40947);
or U41465 (N_41465,N_40758,N_40770);
or U41466 (N_41466,N_40100,N_40526);
and U41467 (N_41467,N_40861,N_40884);
xor U41468 (N_41468,N_40331,N_40169);
nand U41469 (N_41469,N_40739,N_40873);
nor U41470 (N_41470,N_40159,N_40124);
xnor U41471 (N_41471,N_40659,N_40191);
nand U41472 (N_41472,N_40142,N_40019);
or U41473 (N_41473,N_40496,N_40956);
or U41474 (N_41474,N_40430,N_40347);
and U41475 (N_41475,N_40222,N_40291);
nand U41476 (N_41476,N_40427,N_40800);
nand U41477 (N_41477,N_40923,N_40821);
and U41478 (N_41478,N_40435,N_40385);
xor U41479 (N_41479,N_40735,N_40995);
nor U41480 (N_41480,N_40675,N_40939);
and U41481 (N_41481,N_40468,N_40852);
nor U41482 (N_41482,N_40301,N_40746);
nand U41483 (N_41483,N_40574,N_40007);
and U41484 (N_41484,N_40218,N_40280);
and U41485 (N_41485,N_40425,N_40698);
xor U41486 (N_41486,N_40420,N_40595);
xor U41487 (N_41487,N_40309,N_40566);
xnor U41488 (N_41488,N_40503,N_40044);
and U41489 (N_41489,N_40573,N_40604);
and U41490 (N_41490,N_40463,N_40024);
or U41491 (N_41491,N_40518,N_40460);
nand U41492 (N_41492,N_40163,N_40831);
nor U41493 (N_41493,N_40803,N_40504);
nor U41494 (N_41494,N_40838,N_40312);
xor U41495 (N_41495,N_40680,N_40702);
nand U41496 (N_41496,N_40239,N_40713);
nand U41497 (N_41497,N_40092,N_40272);
or U41498 (N_41498,N_40036,N_40186);
and U41499 (N_41499,N_40989,N_40348);
and U41500 (N_41500,N_40219,N_40059);
xor U41501 (N_41501,N_40585,N_40640);
nor U41502 (N_41502,N_40108,N_40236);
or U41503 (N_41503,N_40587,N_40170);
and U41504 (N_41504,N_40849,N_40130);
or U41505 (N_41505,N_40135,N_40275);
nand U41506 (N_41506,N_40857,N_40237);
xor U41507 (N_41507,N_40310,N_40151);
nor U41508 (N_41508,N_40569,N_40504);
nand U41509 (N_41509,N_40305,N_40225);
and U41510 (N_41510,N_40404,N_40791);
and U41511 (N_41511,N_40243,N_40499);
and U41512 (N_41512,N_40010,N_40923);
nor U41513 (N_41513,N_40340,N_40380);
nor U41514 (N_41514,N_40568,N_40024);
nor U41515 (N_41515,N_40889,N_40835);
xor U41516 (N_41516,N_40088,N_40676);
or U41517 (N_41517,N_40881,N_40595);
nand U41518 (N_41518,N_40921,N_40628);
nand U41519 (N_41519,N_40389,N_40512);
xor U41520 (N_41520,N_40687,N_40428);
nand U41521 (N_41521,N_40116,N_40844);
nor U41522 (N_41522,N_40509,N_40425);
or U41523 (N_41523,N_40531,N_40217);
nand U41524 (N_41524,N_40750,N_40968);
and U41525 (N_41525,N_40845,N_40383);
and U41526 (N_41526,N_40035,N_40239);
or U41527 (N_41527,N_40968,N_40944);
and U41528 (N_41528,N_40547,N_40124);
nor U41529 (N_41529,N_40775,N_40772);
or U41530 (N_41530,N_40485,N_40707);
xnor U41531 (N_41531,N_40664,N_40931);
xnor U41532 (N_41532,N_40590,N_40639);
xnor U41533 (N_41533,N_40295,N_40576);
or U41534 (N_41534,N_40939,N_40318);
or U41535 (N_41535,N_40180,N_40573);
nand U41536 (N_41536,N_40363,N_40180);
xnor U41537 (N_41537,N_40136,N_40871);
and U41538 (N_41538,N_40509,N_40004);
or U41539 (N_41539,N_40056,N_40960);
nor U41540 (N_41540,N_40767,N_40396);
nor U41541 (N_41541,N_40086,N_40329);
nor U41542 (N_41542,N_40336,N_40922);
and U41543 (N_41543,N_40990,N_40214);
nand U41544 (N_41544,N_40357,N_40260);
or U41545 (N_41545,N_40658,N_40268);
and U41546 (N_41546,N_40235,N_40163);
nor U41547 (N_41547,N_40357,N_40177);
or U41548 (N_41548,N_40572,N_40893);
nor U41549 (N_41549,N_40596,N_40578);
nor U41550 (N_41550,N_40412,N_40419);
xor U41551 (N_41551,N_40195,N_40220);
and U41552 (N_41552,N_40285,N_40452);
xor U41553 (N_41553,N_40363,N_40614);
nor U41554 (N_41554,N_40184,N_40082);
nor U41555 (N_41555,N_40347,N_40425);
xor U41556 (N_41556,N_40702,N_40143);
or U41557 (N_41557,N_40677,N_40692);
or U41558 (N_41558,N_40078,N_40876);
or U41559 (N_41559,N_40083,N_40717);
nand U41560 (N_41560,N_40887,N_40189);
or U41561 (N_41561,N_40554,N_40298);
nor U41562 (N_41562,N_40476,N_40346);
and U41563 (N_41563,N_40709,N_40719);
and U41564 (N_41564,N_40458,N_40592);
xor U41565 (N_41565,N_40559,N_40275);
or U41566 (N_41566,N_40988,N_40100);
xnor U41567 (N_41567,N_40679,N_40359);
and U41568 (N_41568,N_40894,N_40565);
and U41569 (N_41569,N_40928,N_40828);
and U41570 (N_41570,N_40375,N_40554);
nand U41571 (N_41571,N_40861,N_40469);
nand U41572 (N_41572,N_40492,N_40108);
nor U41573 (N_41573,N_40894,N_40077);
nand U41574 (N_41574,N_40605,N_40810);
xnor U41575 (N_41575,N_40947,N_40413);
and U41576 (N_41576,N_40206,N_40313);
nor U41577 (N_41577,N_40444,N_40849);
nor U41578 (N_41578,N_40133,N_40832);
and U41579 (N_41579,N_40754,N_40198);
nand U41580 (N_41580,N_40540,N_40411);
nand U41581 (N_41581,N_40191,N_40390);
xor U41582 (N_41582,N_40120,N_40121);
nand U41583 (N_41583,N_40940,N_40805);
nor U41584 (N_41584,N_40921,N_40662);
or U41585 (N_41585,N_40759,N_40801);
and U41586 (N_41586,N_40974,N_40752);
and U41587 (N_41587,N_40245,N_40149);
nor U41588 (N_41588,N_40172,N_40149);
or U41589 (N_41589,N_40235,N_40387);
nand U41590 (N_41590,N_40596,N_40169);
and U41591 (N_41591,N_40394,N_40343);
and U41592 (N_41592,N_40981,N_40312);
nor U41593 (N_41593,N_40469,N_40238);
xnor U41594 (N_41594,N_40458,N_40365);
xor U41595 (N_41595,N_40239,N_40500);
nand U41596 (N_41596,N_40699,N_40394);
or U41597 (N_41597,N_40937,N_40761);
nand U41598 (N_41598,N_40993,N_40301);
nand U41599 (N_41599,N_40495,N_40951);
or U41600 (N_41600,N_40477,N_40380);
nor U41601 (N_41601,N_40275,N_40381);
or U41602 (N_41602,N_40340,N_40554);
and U41603 (N_41603,N_40823,N_40405);
nand U41604 (N_41604,N_40157,N_40014);
or U41605 (N_41605,N_40349,N_40526);
nor U41606 (N_41606,N_40230,N_40760);
nor U41607 (N_41607,N_40517,N_40901);
nand U41608 (N_41608,N_40276,N_40121);
and U41609 (N_41609,N_40450,N_40522);
or U41610 (N_41610,N_40174,N_40457);
nand U41611 (N_41611,N_40948,N_40286);
nor U41612 (N_41612,N_40147,N_40526);
nor U41613 (N_41613,N_40769,N_40392);
nand U41614 (N_41614,N_40281,N_40087);
and U41615 (N_41615,N_40738,N_40080);
xnor U41616 (N_41616,N_40521,N_40435);
or U41617 (N_41617,N_40885,N_40222);
and U41618 (N_41618,N_40415,N_40193);
or U41619 (N_41619,N_40795,N_40460);
or U41620 (N_41620,N_40387,N_40779);
and U41621 (N_41621,N_40621,N_40896);
or U41622 (N_41622,N_40329,N_40409);
nand U41623 (N_41623,N_40131,N_40403);
and U41624 (N_41624,N_40340,N_40980);
and U41625 (N_41625,N_40905,N_40079);
and U41626 (N_41626,N_40174,N_40302);
nand U41627 (N_41627,N_40994,N_40918);
nor U41628 (N_41628,N_40959,N_40382);
nand U41629 (N_41629,N_40010,N_40649);
nand U41630 (N_41630,N_40621,N_40771);
xor U41631 (N_41631,N_40656,N_40264);
and U41632 (N_41632,N_40435,N_40789);
nand U41633 (N_41633,N_40635,N_40022);
or U41634 (N_41634,N_40945,N_40442);
xnor U41635 (N_41635,N_40900,N_40870);
nand U41636 (N_41636,N_40412,N_40039);
nand U41637 (N_41637,N_40706,N_40451);
nor U41638 (N_41638,N_40800,N_40187);
or U41639 (N_41639,N_40910,N_40409);
xnor U41640 (N_41640,N_40423,N_40072);
and U41641 (N_41641,N_40451,N_40897);
nand U41642 (N_41642,N_40691,N_40166);
xor U41643 (N_41643,N_40031,N_40585);
and U41644 (N_41644,N_40565,N_40568);
nand U41645 (N_41645,N_40483,N_40298);
or U41646 (N_41646,N_40660,N_40478);
and U41647 (N_41647,N_40557,N_40828);
or U41648 (N_41648,N_40906,N_40629);
nand U41649 (N_41649,N_40108,N_40237);
nand U41650 (N_41650,N_40193,N_40665);
nand U41651 (N_41651,N_40395,N_40426);
xnor U41652 (N_41652,N_40612,N_40281);
and U41653 (N_41653,N_40275,N_40663);
nor U41654 (N_41654,N_40741,N_40721);
nor U41655 (N_41655,N_40715,N_40436);
nor U41656 (N_41656,N_40632,N_40565);
nor U41657 (N_41657,N_40105,N_40257);
or U41658 (N_41658,N_40886,N_40053);
and U41659 (N_41659,N_40905,N_40126);
xnor U41660 (N_41660,N_40833,N_40800);
nand U41661 (N_41661,N_40033,N_40879);
nand U41662 (N_41662,N_40596,N_40203);
nand U41663 (N_41663,N_40677,N_40660);
or U41664 (N_41664,N_40847,N_40772);
and U41665 (N_41665,N_40721,N_40871);
and U41666 (N_41666,N_40989,N_40120);
nand U41667 (N_41667,N_40470,N_40248);
nor U41668 (N_41668,N_40295,N_40588);
xnor U41669 (N_41669,N_40957,N_40149);
or U41670 (N_41670,N_40756,N_40876);
xnor U41671 (N_41671,N_40496,N_40765);
or U41672 (N_41672,N_40615,N_40219);
xnor U41673 (N_41673,N_40692,N_40319);
and U41674 (N_41674,N_40787,N_40927);
and U41675 (N_41675,N_40886,N_40558);
or U41676 (N_41676,N_40824,N_40743);
and U41677 (N_41677,N_40466,N_40068);
or U41678 (N_41678,N_40815,N_40545);
or U41679 (N_41679,N_40892,N_40108);
and U41680 (N_41680,N_40165,N_40963);
and U41681 (N_41681,N_40963,N_40659);
nor U41682 (N_41682,N_40907,N_40581);
or U41683 (N_41683,N_40496,N_40382);
xor U41684 (N_41684,N_40417,N_40693);
or U41685 (N_41685,N_40001,N_40115);
nand U41686 (N_41686,N_40335,N_40169);
xnor U41687 (N_41687,N_40173,N_40379);
and U41688 (N_41688,N_40360,N_40882);
nor U41689 (N_41689,N_40891,N_40315);
nor U41690 (N_41690,N_40076,N_40662);
and U41691 (N_41691,N_40422,N_40063);
or U41692 (N_41692,N_40074,N_40472);
nand U41693 (N_41693,N_40119,N_40578);
and U41694 (N_41694,N_40314,N_40647);
nor U41695 (N_41695,N_40812,N_40792);
nand U41696 (N_41696,N_40212,N_40687);
xnor U41697 (N_41697,N_40054,N_40717);
nand U41698 (N_41698,N_40405,N_40780);
or U41699 (N_41699,N_40413,N_40509);
or U41700 (N_41700,N_40849,N_40019);
nand U41701 (N_41701,N_40355,N_40204);
xnor U41702 (N_41702,N_40302,N_40401);
nor U41703 (N_41703,N_40389,N_40247);
nand U41704 (N_41704,N_40525,N_40165);
xor U41705 (N_41705,N_40047,N_40834);
nor U41706 (N_41706,N_40753,N_40693);
xor U41707 (N_41707,N_40322,N_40439);
xor U41708 (N_41708,N_40968,N_40150);
and U41709 (N_41709,N_40821,N_40406);
xnor U41710 (N_41710,N_40317,N_40748);
nor U41711 (N_41711,N_40689,N_40176);
nor U41712 (N_41712,N_40096,N_40258);
xnor U41713 (N_41713,N_40399,N_40299);
xor U41714 (N_41714,N_40352,N_40926);
xor U41715 (N_41715,N_40652,N_40302);
nand U41716 (N_41716,N_40549,N_40559);
nand U41717 (N_41717,N_40900,N_40817);
or U41718 (N_41718,N_40492,N_40921);
xor U41719 (N_41719,N_40641,N_40592);
and U41720 (N_41720,N_40978,N_40329);
nor U41721 (N_41721,N_40366,N_40263);
nand U41722 (N_41722,N_40047,N_40463);
and U41723 (N_41723,N_40271,N_40590);
nor U41724 (N_41724,N_40039,N_40642);
or U41725 (N_41725,N_40585,N_40174);
xor U41726 (N_41726,N_40404,N_40163);
and U41727 (N_41727,N_40586,N_40019);
nor U41728 (N_41728,N_40014,N_40581);
or U41729 (N_41729,N_40856,N_40838);
nand U41730 (N_41730,N_40083,N_40952);
or U41731 (N_41731,N_40081,N_40507);
and U41732 (N_41732,N_40278,N_40857);
nor U41733 (N_41733,N_40875,N_40291);
nor U41734 (N_41734,N_40668,N_40596);
and U41735 (N_41735,N_40180,N_40104);
or U41736 (N_41736,N_40747,N_40972);
xnor U41737 (N_41737,N_40576,N_40222);
nand U41738 (N_41738,N_40952,N_40981);
xor U41739 (N_41739,N_40317,N_40078);
xor U41740 (N_41740,N_40997,N_40706);
nand U41741 (N_41741,N_40369,N_40400);
xor U41742 (N_41742,N_40183,N_40489);
nand U41743 (N_41743,N_40095,N_40592);
nor U41744 (N_41744,N_40260,N_40818);
xor U41745 (N_41745,N_40137,N_40866);
or U41746 (N_41746,N_40543,N_40517);
xor U41747 (N_41747,N_40346,N_40594);
or U41748 (N_41748,N_40350,N_40701);
or U41749 (N_41749,N_40753,N_40909);
or U41750 (N_41750,N_40486,N_40106);
or U41751 (N_41751,N_40627,N_40488);
or U41752 (N_41752,N_40121,N_40716);
and U41753 (N_41753,N_40465,N_40224);
nand U41754 (N_41754,N_40160,N_40716);
nand U41755 (N_41755,N_40529,N_40242);
xnor U41756 (N_41756,N_40154,N_40920);
or U41757 (N_41757,N_40094,N_40383);
nor U41758 (N_41758,N_40982,N_40625);
nand U41759 (N_41759,N_40399,N_40517);
and U41760 (N_41760,N_40359,N_40969);
and U41761 (N_41761,N_40366,N_40353);
nor U41762 (N_41762,N_40317,N_40745);
xor U41763 (N_41763,N_40110,N_40213);
nor U41764 (N_41764,N_40815,N_40475);
or U41765 (N_41765,N_40582,N_40879);
or U41766 (N_41766,N_40044,N_40312);
and U41767 (N_41767,N_40116,N_40180);
nand U41768 (N_41768,N_40764,N_40312);
or U41769 (N_41769,N_40198,N_40216);
nand U41770 (N_41770,N_40048,N_40350);
or U41771 (N_41771,N_40012,N_40212);
nand U41772 (N_41772,N_40818,N_40314);
nor U41773 (N_41773,N_40846,N_40543);
nor U41774 (N_41774,N_40169,N_40106);
nor U41775 (N_41775,N_40509,N_40511);
and U41776 (N_41776,N_40396,N_40497);
nor U41777 (N_41777,N_40621,N_40326);
nor U41778 (N_41778,N_40000,N_40325);
nand U41779 (N_41779,N_40410,N_40005);
nand U41780 (N_41780,N_40368,N_40524);
nand U41781 (N_41781,N_40058,N_40351);
xor U41782 (N_41782,N_40726,N_40392);
xnor U41783 (N_41783,N_40207,N_40387);
xor U41784 (N_41784,N_40165,N_40628);
or U41785 (N_41785,N_40873,N_40077);
nor U41786 (N_41786,N_40002,N_40504);
nor U41787 (N_41787,N_40225,N_40391);
xor U41788 (N_41788,N_40178,N_40100);
xnor U41789 (N_41789,N_40907,N_40816);
xor U41790 (N_41790,N_40264,N_40914);
or U41791 (N_41791,N_40023,N_40204);
nor U41792 (N_41792,N_40527,N_40784);
or U41793 (N_41793,N_40537,N_40751);
nor U41794 (N_41794,N_40225,N_40339);
or U41795 (N_41795,N_40889,N_40340);
and U41796 (N_41796,N_40387,N_40565);
nand U41797 (N_41797,N_40040,N_40000);
nor U41798 (N_41798,N_40276,N_40307);
xor U41799 (N_41799,N_40165,N_40541);
and U41800 (N_41800,N_40568,N_40148);
nor U41801 (N_41801,N_40983,N_40923);
nor U41802 (N_41802,N_40070,N_40746);
and U41803 (N_41803,N_40418,N_40521);
nor U41804 (N_41804,N_40085,N_40436);
xor U41805 (N_41805,N_40911,N_40178);
nor U41806 (N_41806,N_40288,N_40831);
and U41807 (N_41807,N_40869,N_40684);
nor U41808 (N_41808,N_40147,N_40375);
xnor U41809 (N_41809,N_40906,N_40851);
nor U41810 (N_41810,N_40493,N_40833);
xor U41811 (N_41811,N_40794,N_40710);
or U41812 (N_41812,N_40409,N_40392);
nand U41813 (N_41813,N_40537,N_40349);
nor U41814 (N_41814,N_40764,N_40899);
and U41815 (N_41815,N_40712,N_40812);
xor U41816 (N_41816,N_40478,N_40598);
nand U41817 (N_41817,N_40034,N_40666);
and U41818 (N_41818,N_40809,N_40365);
or U41819 (N_41819,N_40395,N_40070);
nand U41820 (N_41820,N_40545,N_40886);
nand U41821 (N_41821,N_40792,N_40150);
nor U41822 (N_41822,N_40157,N_40426);
xor U41823 (N_41823,N_40675,N_40480);
or U41824 (N_41824,N_40806,N_40116);
or U41825 (N_41825,N_40640,N_40873);
nand U41826 (N_41826,N_40629,N_40337);
and U41827 (N_41827,N_40188,N_40076);
or U41828 (N_41828,N_40528,N_40092);
and U41829 (N_41829,N_40272,N_40343);
nand U41830 (N_41830,N_40249,N_40278);
nor U41831 (N_41831,N_40571,N_40558);
and U41832 (N_41832,N_40857,N_40116);
nand U41833 (N_41833,N_40712,N_40562);
nand U41834 (N_41834,N_40524,N_40615);
xnor U41835 (N_41835,N_40319,N_40625);
xor U41836 (N_41836,N_40156,N_40669);
and U41837 (N_41837,N_40103,N_40393);
xnor U41838 (N_41838,N_40281,N_40481);
nand U41839 (N_41839,N_40292,N_40803);
or U41840 (N_41840,N_40422,N_40056);
and U41841 (N_41841,N_40988,N_40139);
xnor U41842 (N_41842,N_40516,N_40926);
and U41843 (N_41843,N_40059,N_40798);
xor U41844 (N_41844,N_40478,N_40177);
nand U41845 (N_41845,N_40174,N_40540);
or U41846 (N_41846,N_40423,N_40320);
or U41847 (N_41847,N_40624,N_40056);
and U41848 (N_41848,N_40310,N_40636);
xnor U41849 (N_41849,N_40951,N_40297);
nand U41850 (N_41850,N_40769,N_40359);
xnor U41851 (N_41851,N_40472,N_40498);
and U41852 (N_41852,N_40849,N_40384);
or U41853 (N_41853,N_40209,N_40803);
xor U41854 (N_41854,N_40308,N_40529);
or U41855 (N_41855,N_40854,N_40978);
xnor U41856 (N_41856,N_40930,N_40132);
or U41857 (N_41857,N_40856,N_40775);
or U41858 (N_41858,N_40175,N_40170);
and U41859 (N_41859,N_40490,N_40768);
nand U41860 (N_41860,N_40732,N_40113);
and U41861 (N_41861,N_40515,N_40570);
or U41862 (N_41862,N_40971,N_40630);
nand U41863 (N_41863,N_40731,N_40809);
and U41864 (N_41864,N_40247,N_40028);
or U41865 (N_41865,N_40368,N_40985);
and U41866 (N_41866,N_40048,N_40016);
xor U41867 (N_41867,N_40146,N_40244);
xnor U41868 (N_41868,N_40922,N_40258);
or U41869 (N_41869,N_40724,N_40207);
or U41870 (N_41870,N_40203,N_40839);
xnor U41871 (N_41871,N_40149,N_40176);
and U41872 (N_41872,N_40380,N_40782);
or U41873 (N_41873,N_40264,N_40828);
and U41874 (N_41874,N_40266,N_40190);
nand U41875 (N_41875,N_40457,N_40580);
nor U41876 (N_41876,N_40152,N_40092);
nor U41877 (N_41877,N_40781,N_40993);
nor U41878 (N_41878,N_40213,N_40602);
nor U41879 (N_41879,N_40197,N_40146);
and U41880 (N_41880,N_40747,N_40000);
xor U41881 (N_41881,N_40690,N_40807);
nor U41882 (N_41882,N_40853,N_40326);
xnor U41883 (N_41883,N_40911,N_40062);
nand U41884 (N_41884,N_40397,N_40171);
nand U41885 (N_41885,N_40580,N_40991);
or U41886 (N_41886,N_40077,N_40901);
xor U41887 (N_41887,N_40186,N_40339);
nand U41888 (N_41888,N_40901,N_40267);
and U41889 (N_41889,N_40162,N_40363);
or U41890 (N_41890,N_40805,N_40156);
nand U41891 (N_41891,N_40004,N_40098);
nor U41892 (N_41892,N_40913,N_40745);
nand U41893 (N_41893,N_40981,N_40294);
or U41894 (N_41894,N_40658,N_40527);
xnor U41895 (N_41895,N_40509,N_40646);
or U41896 (N_41896,N_40527,N_40018);
and U41897 (N_41897,N_40462,N_40572);
and U41898 (N_41898,N_40893,N_40990);
and U41899 (N_41899,N_40135,N_40447);
nand U41900 (N_41900,N_40865,N_40248);
and U41901 (N_41901,N_40110,N_40333);
nand U41902 (N_41902,N_40448,N_40761);
xor U41903 (N_41903,N_40320,N_40461);
nor U41904 (N_41904,N_40127,N_40284);
nor U41905 (N_41905,N_40406,N_40549);
nor U41906 (N_41906,N_40984,N_40761);
and U41907 (N_41907,N_40699,N_40763);
and U41908 (N_41908,N_40995,N_40092);
or U41909 (N_41909,N_40580,N_40273);
and U41910 (N_41910,N_40872,N_40768);
or U41911 (N_41911,N_40948,N_40670);
xnor U41912 (N_41912,N_40201,N_40746);
nand U41913 (N_41913,N_40377,N_40691);
xor U41914 (N_41914,N_40331,N_40629);
nor U41915 (N_41915,N_40902,N_40844);
and U41916 (N_41916,N_40746,N_40589);
nand U41917 (N_41917,N_40855,N_40399);
xor U41918 (N_41918,N_40936,N_40385);
and U41919 (N_41919,N_40452,N_40457);
nor U41920 (N_41920,N_40556,N_40111);
or U41921 (N_41921,N_40445,N_40878);
or U41922 (N_41922,N_40500,N_40517);
nor U41923 (N_41923,N_40402,N_40306);
and U41924 (N_41924,N_40937,N_40777);
nor U41925 (N_41925,N_40425,N_40422);
xnor U41926 (N_41926,N_40511,N_40922);
xor U41927 (N_41927,N_40632,N_40395);
xor U41928 (N_41928,N_40943,N_40069);
nand U41929 (N_41929,N_40413,N_40404);
nor U41930 (N_41930,N_40549,N_40099);
and U41931 (N_41931,N_40265,N_40617);
or U41932 (N_41932,N_40222,N_40481);
xnor U41933 (N_41933,N_40364,N_40176);
and U41934 (N_41934,N_40362,N_40404);
nor U41935 (N_41935,N_40870,N_40430);
and U41936 (N_41936,N_40701,N_40580);
nand U41937 (N_41937,N_40243,N_40612);
or U41938 (N_41938,N_40089,N_40158);
or U41939 (N_41939,N_40159,N_40600);
nand U41940 (N_41940,N_40655,N_40697);
nor U41941 (N_41941,N_40116,N_40765);
or U41942 (N_41942,N_40066,N_40208);
xor U41943 (N_41943,N_40274,N_40635);
xor U41944 (N_41944,N_40630,N_40967);
and U41945 (N_41945,N_40951,N_40185);
or U41946 (N_41946,N_40666,N_40000);
or U41947 (N_41947,N_40982,N_40033);
and U41948 (N_41948,N_40035,N_40396);
or U41949 (N_41949,N_40211,N_40573);
or U41950 (N_41950,N_40614,N_40524);
and U41951 (N_41951,N_40862,N_40956);
xor U41952 (N_41952,N_40715,N_40581);
xor U41953 (N_41953,N_40222,N_40876);
nor U41954 (N_41954,N_40910,N_40334);
nor U41955 (N_41955,N_40392,N_40559);
xor U41956 (N_41956,N_40276,N_40254);
and U41957 (N_41957,N_40640,N_40295);
and U41958 (N_41958,N_40783,N_40942);
or U41959 (N_41959,N_40986,N_40140);
and U41960 (N_41960,N_40267,N_40171);
and U41961 (N_41961,N_40069,N_40679);
and U41962 (N_41962,N_40894,N_40533);
nand U41963 (N_41963,N_40169,N_40614);
and U41964 (N_41964,N_40141,N_40823);
nor U41965 (N_41965,N_40554,N_40741);
or U41966 (N_41966,N_40149,N_40145);
or U41967 (N_41967,N_40370,N_40603);
nor U41968 (N_41968,N_40145,N_40283);
nand U41969 (N_41969,N_40958,N_40611);
nor U41970 (N_41970,N_40000,N_40457);
or U41971 (N_41971,N_40628,N_40607);
xor U41972 (N_41972,N_40846,N_40547);
and U41973 (N_41973,N_40965,N_40340);
or U41974 (N_41974,N_40723,N_40181);
and U41975 (N_41975,N_40299,N_40908);
or U41976 (N_41976,N_40644,N_40466);
or U41977 (N_41977,N_40761,N_40466);
xor U41978 (N_41978,N_40071,N_40553);
and U41979 (N_41979,N_40727,N_40021);
or U41980 (N_41980,N_40382,N_40129);
nand U41981 (N_41981,N_40952,N_40333);
nor U41982 (N_41982,N_40908,N_40318);
nor U41983 (N_41983,N_40990,N_40229);
and U41984 (N_41984,N_40918,N_40125);
or U41985 (N_41985,N_40408,N_40911);
and U41986 (N_41986,N_40938,N_40907);
nand U41987 (N_41987,N_40565,N_40647);
nand U41988 (N_41988,N_40101,N_40453);
xnor U41989 (N_41989,N_40666,N_40092);
nor U41990 (N_41990,N_40422,N_40858);
or U41991 (N_41991,N_40881,N_40986);
nand U41992 (N_41992,N_40016,N_40222);
nor U41993 (N_41993,N_40278,N_40775);
xor U41994 (N_41994,N_40865,N_40394);
or U41995 (N_41995,N_40164,N_40524);
and U41996 (N_41996,N_40522,N_40684);
xor U41997 (N_41997,N_40165,N_40714);
or U41998 (N_41998,N_40772,N_40802);
and U41999 (N_41999,N_40296,N_40733);
and U42000 (N_42000,N_41466,N_41139);
and U42001 (N_42001,N_41358,N_41828);
nand U42002 (N_42002,N_41720,N_41025);
nand U42003 (N_42003,N_41729,N_41245);
xor U42004 (N_42004,N_41799,N_41768);
or U42005 (N_42005,N_41052,N_41334);
nand U42006 (N_42006,N_41685,N_41581);
xor U42007 (N_42007,N_41123,N_41375);
xnor U42008 (N_42008,N_41457,N_41817);
or U42009 (N_42009,N_41395,N_41340);
and U42010 (N_42010,N_41699,N_41028);
xor U42011 (N_42011,N_41985,N_41066);
xnor U42012 (N_42012,N_41006,N_41185);
nor U42013 (N_42013,N_41343,N_41984);
or U42014 (N_42014,N_41109,N_41550);
and U42015 (N_42015,N_41670,N_41210);
and U42016 (N_42016,N_41121,N_41382);
or U42017 (N_42017,N_41861,N_41671);
nand U42018 (N_42018,N_41976,N_41418);
nor U42019 (N_42019,N_41273,N_41863);
xnor U42020 (N_42020,N_41240,N_41002);
and U42021 (N_42021,N_41431,N_41763);
nand U42022 (N_42022,N_41308,N_41300);
nand U42023 (N_42023,N_41241,N_41362);
xor U42024 (N_42024,N_41355,N_41184);
xor U42025 (N_42025,N_41281,N_41790);
and U42026 (N_42026,N_41713,N_41331);
nand U42027 (N_42027,N_41305,N_41092);
xor U42028 (N_42028,N_41909,N_41638);
nand U42029 (N_42029,N_41607,N_41392);
nor U42030 (N_42030,N_41858,N_41596);
or U42031 (N_42031,N_41757,N_41136);
xor U42032 (N_42032,N_41841,N_41654);
nand U42033 (N_42033,N_41243,N_41318);
and U42034 (N_42034,N_41405,N_41045);
nand U42035 (N_42035,N_41107,N_41467);
nand U42036 (N_42036,N_41950,N_41055);
and U42037 (N_42037,N_41365,N_41862);
xor U42038 (N_42038,N_41703,N_41625);
and U42039 (N_42039,N_41824,N_41187);
nand U42040 (N_42040,N_41738,N_41851);
nor U42041 (N_42041,N_41421,N_41250);
and U42042 (N_42042,N_41260,N_41887);
nor U42043 (N_42043,N_41749,N_41366);
nand U42044 (N_42044,N_41016,N_41856);
nor U42045 (N_42045,N_41419,N_41777);
nand U42046 (N_42046,N_41577,N_41645);
nand U42047 (N_42047,N_41113,N_41403);
nor U42048 (N_42048,N_41428,N_41277);
and U42049 (N_42049,N_41439,N_41193);
nand U42050 (N_42050,N_41056,N_41259);
and U42051 (N_42051,N_41849,N_41748);
or U42052 (N_42052,N_41708,N_41565);
or U42053 (N_42053,N_41662,N_41915);
nand U42054 (N_42054,N_41425,N_41486);
nand U42055 (N_42055,N_41021,N_41942);
and U42056 (N_42056,N_41935,N_41735);
or U42057 (N_42057,N_41682,N_41034);
and U42058 (N_42058,N_41474,N_41829);
or U42059 (N_42059,N_41339,N_41093);
nor U42060 (N_42060,N_41619,N_41801);
or U42061 (N_42061,N_41301,N_41188);
and U42062 (N_42062,N_41000,N_41320);
and U42063 (N_42063,N_41914,N_41992);
and U42064 (N_42064,N_41541,N_41401);
and U42065 (N_42065,N_41153,N_41632);
nand U42066 (N_42066,N_41999,N_41356);
nor U42067 (N_42067,N_41567,N_41981);
nand U42068 (N_42068,N_41499,N_41520);
nor U42069 (N_42069,N_41787,N_41737);
nor U42070 (N_42070,N_41222,N_41916);
xor U42071 (N_42071,N_41227,N_41733);
nand U42072 (N_42072,N_41866,N_41328);
and U42073 (N_42073,N_41716,N_41007);
xor U42074 (N_42074,N_41588,N_41404);
or U42075 (N_42075,N_41201,N_41566);
nor U42076 (N_42076,N_41623,N_41324);
or U42077 (N_42077,N_41551,N_41678);
nand U42078 (N_42078,N_41722,N_41746);
nand U42079 (N_42079,N_41199,N_41159);
nor U42080 (N_42080,N_41723,N_41311);
nor U42081 (N_42081,N_41693,N_41770);
nand U42082 (N_42082,N_41811,N_41399);
nand U42083 (N_42083,N_41162,N_41473);
or U42084 (N_42084,N_41297,N_41264);
or U42085 (N_42085,N_41037,N_41884);
nor U42086 (N_42086,N_41043,N_41456);
xor U42087 (N_42087,N_41017,N_41253);
and U42088 (N_42088,N_41701,N_41569);
or U42089 (N_42089,N_41561,N_41830);
xnor U42090 (N_42090,N_41195,N_41144);
nand U42091 (N_42091,N_41917,N_41774);
nand U42092 (N_42092,N_41954,N_41333);
nand U42093 (N_42093,N_41600,N_41203);
or U42094 (N_42094,N_41986,N_41628);
nand U42095 (N_42095,N_41657,N_41562);
or U42096 (N_42096,N_41347,N_41026);
or U42097 (N_42097,N_41674,N_41249);
and U42098 (N_42098,N_41510,N_41911);
nor U42099 (N_42099,N_41819,N_41663);
and U42100 (N_42100,N_41163,N_41758);
nor U42101 (N_42101,N_41272,N_41364);
or U42102 (N_42102,N_41476,N_41594);
and U42103 (N_42103,N_41357,N_41317);
xor U42104 (N_42104,N_41635,N_41953);
nand U42105 (N_42105,N_41627,N_41462);
and U42106 (N_42106,N_41665,N_41642);
nand U42107 (N_42107,N_41054,N_41238);
or U42108 (N_42108,N_41212,N_41711);
or U42109 (N_42109,N_41445,N_41501);
xor U42110 (N_42110,N_41725,N_41079);
nor U42111 (N_42111,N_41962,N_41689);
xor U42112 (N_42112,N_41387,N_41621);
and U42113 (N_42113,N_41995,N_41389);
nor U42114 (N_42114,N_41837,N_41527);
nand U42115 (N_42115,N_41064,N_41891);
nand U42116 (N_42116,N_41480,N_41289);
nor U42117 (N_42117,N_41767,N_41102);
and U42118 (N_42118,N_41591,N_41046);
or U42119 (N_42119,N_41142,N_41815);
nor U42120 (N_42120,N_41233,N_41951);
nand U42121 (N_42121,N_41108,N_41704);
xor U42122 (N_42122,N_41570,N_41279);
or U42123 (N_42123,N_41743,N_41785);
nor U42124 (N_42124,N_41971,N_41047);
xor U42125 (N_42125,N_41280,N_41420);
nor U42126 (N_42126,N_41417,N_41434);
xnor U42127 (N_42127,N_41410,N_41881);
xnor U42128 (N_42128,N_41922,N_41666);
nand U42129 (N_42129,N_41702,N_41393);
or U42130 (N_42130,N_41274,N_41105);
xor U42131 (N_42131,N_41945,N_41798);
or U42132 (N_42132,N_41397,N_41530);
and U42133 (N_42133,N_41948,N_41468);
nor U42134 (N_42134,N_41342,N_41230);
or U42135 (N_42135,N_41062,N_41788);
nor U42136 (N_42136,N_41871,N_41656);
and U42137 (N_42137,N_41802,N_41049);
nand U42138 (N_42138,N_41870,N_41744);
and U42139 (N_42139,N_41571,N_41460);
or U42140 (N_42140,N_41526,N_41269);
and U42141 (N_42141,N_41218,N_41011);
and U42142 (N_42142,N_41997,N_41082);
nand U42143 (N_42143,N_41680,N_41578);
nand U42144 (N_42144,N_41469,N_41634);
xor U42145 (N_42145,N_41112,N_41327);
nor U42146 (N_42146,N_41030,N_41033);
nand U42147 (N_42147,N_41545,N_41715);
or U42148 (N_42148,N_41736,N_41537);
nor U42149 (N_42149,N_41974,N_41923);
and U42150 (N_42150,N_41424,N_41455);
and U42151 (N_42151,N_41536,N_41487);
and U42152 (N_42152,N_41321,N_41001);
or U42153 (N_42153,N_41146,N_41225);
and U42154 (N_42154,N_41560,N_41038);
nand U42155 (N_42155,N_41549,N_41574);
nor U42156 (N_42156,N_41521,N_41080);
nor U42157 (N_42157,N_41073,N_41061);
nand U42158 (N_42158,N_41874,N_41989);
nor U42159 (N_42159,N_41831,N_41104);
and U42160 (N_42160,N_41765,N_41888);
nor U42161 (N_42161,N_41676,N_41544);
nand U42162 (N_42162,N_41009,N_41067);
or U42163 (N_42163,N_41370,N_41369);
or U42164 (N_42164,N_41019,N_41620);
or U42165 (N_42165,N_41091,N_41247);
or U42166 (N_42166,N_41805,N_41004);
and U42167 (N_42167,N_41940,N_41673);
nor U42168 (N_42168,N_41859,N_41122);
xor U42169 (N_42169,N_41116,N_41630);
xnor U42170 (N_42170,N_41154,N_41813);
or U42171 (N_42171,N_41015,N_41883);
and U42172 (N_42172,N_41616,N_41117);
nor U42173 (N_42173,N_41132,N_41934);
and U42174 (N_42174,N_41111,N_41381);
and U42175 (N_42175,N_41338,N_41406);
and U42176 (N_42176,N_41794,N_41414);
xor U42177 (N_42177,N_41453,N_41552);
or U42178 (N_42178,N_41438,N_41857);
nand U42179 (N_42179,N_41939,N_41470);
or U42180 (N_42180,N_41543,N_41659);
nand U42181 (N_42181,N_41961,N_41533);
xnor U42182 (N_42182,N_41088,N_41416);
or U42183 (N_42183,N_41285,N_41609);
nand U42184 (N_42184,N_41826,N_41959);
or U42185 (N_42185,N_41584,N_41221);
nor U42186 (N_42186,N_41148,N_41895);
nor U42187 (N_42187,N_41361,N_41430);
or U42188 (N_42188,N_41205,N_41189);
or U42189 (N_42189,N_41529,N_41993);
nand U42190 (N_42190,N_41484,N_41374);
xor U42191 (N_42191,N_41947,N_41683);
and U42192 (N_42192,N_41714,N_41293);
or U42193 (N_42193,N_41070,N_41523);
xor U42194 (N_42194,N_41252,N_41348);
or U42195 (N_42195,N_41335,N_41766);
nand U42196 (N_42196,N_41795,N_41119);
or U42197 (N_42197,N_41603,N_41178);
or U42198 (N_42198,N_41782,N_41991);
and U42199 (N_42199,N_41488,N_41576);
or U42200 (N_42200,N_41727,N_41898);
nand U42201 (N_42201,N_41039,N_41675);
nor U42202 (N_42202,N_41215,N_41394);
xor U42203 (N_42203,N_41265,N_41681);
or U42204 (N_42204,N_41482,N_41943);
xor U42205 (N_42205,N_41402,N_41161);
xnor U42206 (N_42206,N_41970,N_41373);
xor U42207 (N_42207,N_41595,N_41204);
xor U42208 (N_42208,N_41155,N_41865);
nand U42209 (N_42209,N_41302,N_41003);
and U42210 (N_42210,N_41496,N_41459);
and U42211 (N_42211,N_41847,N_41156);
and U42212 (N_42212,N_41312,N_41332);
nand U42213 (N_42213,N_41429,N_41775);
or U42214 (N_42214,N_41979,N_41756);
nor U42215 (N_42215,N_41937,N_41839);
xnor U42216 (N_42216,N_41843,N_41877);
and U42217 (N_42217,N_41718,N_41446);
or U42218 (N_42218,N_41465,N_41008);
and U42219 (N_42219,N_41987,N_41602);
xnor U42220 (N_42220,N_41170,N_41691);
nor U42221 (N_42221,N_41441,N_41214);
or U42222 (N_42222,N_41388,N_41919);
nor U42223 (N_42223,N_41747,N_41506);
or U42224 (N_42224,N_41792,N_41236);
nor U42225 (N_42225,N_41294,N_41651);
and U42226 (N_42226,N_41918,N_41341);
xor U42227 (N_42227,N_41739,N_41282);
nand U42228 (N_42228,N_41885,N_41140);
xor U42229 (N_42229,N_41485,N_41427);
nand U42230 (N_42230,N_41936,N_41271);
nand U42231 (N_42231,N_41946,N_41323);
nor U42232 (N_42232,N_41700,N_41372);
nor U42233 (N_42233,N_41071,N_41029);
nand U42234 (N_42234,N_41044,N_41622);
nor U42235 (N_42235,N_41653,N_41901);
or U42236 (N_42236,N_41069,N_41612);
or U42237 (N_42237,N_41207,N_41315);
or U42238 (N_42238,N_41796,N_41791);
nor U42239 (N_42239,N_41228,N_41237);
or U42240 (N_42240,N_41579,N_41745);
or U42241 (N_42241,N_41732,N_41614);
nor U42242 (N_42242,N_41165,N_41631);
nor U42243 (N_42243,N_41712,N_41076);
or U42244 (N_42244,N_41169,N_41921);
nor U42245 (N_42245,N_41152,N_41353);
nor U42246 (N_42246,N_41085,N_41930);
xnor U42247 (N_42247,N_41505,N_41449);
xor U42248 (N_42248,N_41647,N_41310);
xnor U42249 (N_42249,N_41513,N_41068);
and U42250 (N_42250,N_41514,N_41927);
xor U42251 (N_42251,N_41896,N_41672);
nand U42252 (N_42252,N_41980,N_41160);
and U42253 (N_42253,N_41925,N_41040);
or U42254 (N_42254,N_41229,N_41624);
xnor U42255 (N_42255,N_41778,N_41721);
and U42256 (N_42256,N_41127,N_41296);
xnor U42257 (N_42257,N_41090,N_41451);
or U42258 (N_42258,N_41910,N_41955);
xnor U42259 (N_42259,N_41907,N_41728);
or U42260 (N_42260,N_41875,N_41211);
nor U42261 (N_42261,N_41330,N_41924);
nor U42262 (N_42262,N_41409,N_41359);
and U42263 (N_42263,N_41141,N_41844);
nor U42264 (N_42264,N_41626,N_41966);
and U42265 (N_42265,N_41741,N_41268);
xor U42266 (N_42266,N_41809,N_41690);
xnor U42267 (N_42267,N_41816,N_41679);
xnor U42268 (N_42268,N_41423,N_41650);
nand U42269 (N_42269,N_41180,N_41027);
xnor U42270 (N_42270,N_41542,N_41564);
nor U42271 (N_42271,N_41575,N_41894);
or U42272 (N_42272,N_41035,N_41825);
or U42273 (N_42273,N_41590,N_41483);
xnor U42274 (N_42274,N_41692,N_41806);
nor U42275 (N_42275,N_41608,N_41492);
xor U42276 (N_42276,N_41903,N_41978);
or U42277 (N_42277,N_41440,N_41316);
nor U42278 (N_42278,N_41695,N_41171);
nor U42279 (N_42279,N_41648,N_41617);
nor U42280 (N_42280,N_41437,N_41705);
xnor U42281 (N_42281,N_41593,N_41539);
or U42282 (N_42282,N_41175,N_41827);
or U42283 (N_42283,N_41511,N_41649);
nand U42284 (N_42284,N_41731,N_41823);
nand U42285 (N_42285,N_41208,N_41100);
xnor U42286 (N_42286,N_41835,N_41196);
or U42287 (N_42287,N_41833,N_41640);
and U42288 (N_42288,N_41504,N_41597);
or U42289 (N_42289,N_41125,N_41753);
nand U42290 (N_42290,N_41257,N_41478);
or U42291 (N_42291,N_41181,N_41773);
or U42292 (N_42292,N_41426,N_41760);
nand U42293 (N_42293,N_41652,N_41251);
and U42294 (N_42294,N_41754,N_41036);
nand U42295 (N_42295,N_41458,N_41326);
nand U42296 (N_42296,N_41868,N_41051);
and U42297 (N_42297,N_41598,N_41694);
and U42298 (N_42298,N_41442,N_41479);
or U42299 (N_42299,N_41309,N_41968);
nand U42300 (N_42300,N_41965,N_41495);
nand U42301 (N_42301,N_41838,N_41179);
and U42302 (N_42302,N_41717,N_41698);
or U42303 (N_42303,N_41078,N_41912);
xor U42304 (N_42304,N_41752,N_41553);
xor U42305 (N_42305,N_41267,N_41547);
and U42306 (N_42306,N_41548,N_41899);
nor U42307 (N_42307,N_41696,N_41147);
nor U42308 (N_42308,N_41385,N_41314);
and U42309 (N_42309,N_41836,N_41292);
or U42310 (N_42310,N_41655,N_41095);
nor U42311 (N_42311,N_41135,N_41502);
xor U42312 (N_42312,N_41941,N_41854);
and U42313 (N_42313,N_41878,N_41779);
xnor U42314 (N_42314,N_41531,N_41256);
nor U42315 (N_42315,N_41599,N_41065);
xor U42316 (N_42316,N_41083,N_41246);
and U42317 (N_42317,N_41099,N_41262);
nand U42318 (N_42318,N_41337,N_41783);
nand U42319 (N_42319,N_41503,N_41284);
nor U42320 (N_42320,N_41604,N_41150);
xnor U42321 (N_42321,N_41500,N_41557);
nand U42322 (N_42322,N_41890,N_41508);
nor U42323 (N_42323,N_41846,N_41512);
or U42324 (N_42324,N_41772,N_41864);
nor U42325 (N_42325,N_41448,N_41920);
nand U42326 (N_42326,N_41464,N_41053);
nor U42327 (N_42327,N_41166,N_41586);
xor U42328 (N_42328,N_41050,N_41759);
nor U42329 (N_42329,N_41516,N_41850);
or U42330 (N_42330,N_41018,N_41130);
nor U42331 (N_42331,N_41601,N_41475);
or U42332 (N_42332,N_41618,N_41555);
nand U42333 (N_42333,N_41780,N_41658);
or U42334 (N_42334,N_41730,N_41220);
or U42335 (N_42335,N_41967,N_41519);
and U42336 (N_42336,N_41288,N_41048);
nand U42337 (N_42337,N_41145,N_41063);
and U42338 (N_42338,N_41244,N_41589);
or U42339 (N_42339,N_41810,N_41764);
xor U42340 (N_42340,N_41287,N_41568);
and U42341 (N_42341,N_41734,N_41190);
and U42342 (N_42342,N_41223,N_41643);
or U42343 (N_42343,N_41538,N_41074);
xor U42344 (N_42344,N_41808,N_41855);
and U42345 (N_42345,N_41615,N_41688);
or U42346 (N_42346,N_41014,N_41477);
nor U42347 (N_42347,N_41020,N_41969);
nand U42348 (N_42348,N_41192,N_41303);
xor U42349 (N_42349,N_41814,N_41345);
xor U42350 (N_42350,N_41902,N_41174);
xor U42351 (N_42351,N_41173,N_41452);
or U42352 (N_42352,N_41224,N_41972);
xor U42353 (N_42353,N_41086,N_41128);
xor U42354 (N_42354,N_41270,N_41528);
nor U42355 (N_42355,N_41194,N_41234);
and U42356 (N_42356,N_41908,N_41217);
xnor U42357 (N_42357,N_41306,N_41637);
nand U42358 (N_42358,N_41024,N_41592);
nor U42359 (N_42359,N_41834,N_41059);
and U42360 (N_42360,N_41167,N_41023);
or U42361 (N_42361,N_41186,N_41411);
and U42362 (N_42362,N_41860,N_41363);
or U42363 (N_42363,N_41143,N_41384);
nor U42364 (N_42364,N_41761,N_41360);
nor U42365 (N_42365,N_41278,N_41867);
and U42366 (N_42366,N_41060,N_41820);
nor U42367 (N_42367,N_41707,N_41376);
and U42368 (N_42368,N_41115,N_41325);
xor U42369 (N_42369,N_41789,N_41371);
or U42370 (N_42370,N_41821,N_41304);
nand U42371 (N_42371,N_41982,N_41202);
or U42372 (N_42372,N_41182,N_41087);
nor U42373 (N_42373,N_41793,N_41398);
nand U42374 (N_42374,N_41509,N_41491);
and U42375 (N_42375,N_41963,N_41042);
xor U42376 (N_42376,N_41216,N_41436);
nor U42377 (N_42377,N_41075,N_41176);
and U42378 (N_42378,N_41351,N_41893);
and U42379 (N_42379,N_41769,N_41299);
xor U42380 (N_42380,N_41904,N_41498);
xnor U42381 (N_42381,N_41724,N_41797);
xor U42382 (N_42382,N_41905,N_41964);
xnor U42383 (N_42383,N_41879,N_41886);
and U42384 (N_42384,N_41261,N_41869);
nand U42385 (N_42385,N_41507,N_41582);
nor U42386 (N_42386,N_41077,N_41433);
nor U42387 (N_42387,N_41956,N_41022);
nor U42388 (N_42388,N_41726,N_41913);
and U42389 (N_42389,N_41636,N_41290);
and U42390 (N_42390,N_41977,N_41800);
and U42391 (N_42391,N_41669,N_41149);
and U42392 (N_42392,N_41784,N_41686);
xor U42393 (N_42393,N_41832,N_41771);
xnor U42394 (N_42394,N_41933,N_41239);
or U42395 (N_42395,N_41641,N_41276);
or U42396 (N_42396,N_41629,N_41639);
or U42397 (N_42397,N_41413,N_41706);
or U42398 (N_42398,N_41710,N_41081);
xor U42399 (N_42399,N_41200,N_41750);
or U42400 (N_42400,N_41709,N_41957);
and U42401 (N_42401,N_41412,N_41687);
xor U42402 (N_42402,N_41131,N_41906);
nor U42403 (N_42403,N_41329,N_41248);
xor U42404 (N_42404,N_41872,N_41900);
or U42405 (N_42405,N_41546,N_41447);
or U42406 (N_42406,N_41336,N_41646);
and U42407 (N_42407,N_41120,N_41103);
nor U42408 (N_42408,N_41283,N_41892);
and U42409 (N_42409,N_41454,N_41880);
nand U42410 (N_42410,N_41667,N_41522);
nor U42411 (N_42411,N_41661,N_41461);
xnor U42412 (N_42412,N_41344,N_41932);
or U42413 (N_42413,N_41041,N_41400);
nand U42414 (N_42414,N_41138,N_41534);
xnor U42415 (N_42415,N_41380,N_41379);
nor U42416 (N_42416,N_41209,N_41346);
and U42417 (N_42417,N_41390,N_41463);
xor U42418 (N_42418,N_41151,N_41101);
xnor U42419 (N_42419,N_41213,N_41852);
nand U42420 (N_42420,N_41254,N_41298);
or U42421 (N_42421,N_41089,N_41032);
and U42422 (N_42422,N_41383,N_41106);
nand U42423 (N_42423,N_41354,N_41515);
xnor U42424 (N_42424,N_41494,N_41481);
and U42425 (N_42425,N_41096,N_41391);
and U42426 (N_42426,N_41818,N_41191);
nor U42427 (N_42427,N_41559,N_41206);
xnor U42428 (N_42428,N_41133,N_41563);
nor U42429 (N_42429,N_41263,N_41804);
xor U42430 (N_42430,N_41554,N_41408);
or U42431 (N_42431,N_41926,N_41944);
or U42432 (N_42432,N_41605,N_41422);
and U42433 (N_42433,N_41235,N_41938);
or U42434 (N_42434,N_41580,N_41803);
nor U42435 (N_42435,N_41958,N_41988);
nor U42436 (N_42436,N_41435,N_41084);
xor U42437 (N_42437,N_41443,N_41882);
nand U42438 (N_42438,N_41489,N_41848);
and U42439 (N_42439,N_41097,N_41010);
nand U42440 (N_42440,N_41493,N_41258);
nor U42441 (N_42441,N_41172,N_41057);
or U42442 (N_42442,N_41517,N_41996);
nor U42443 (N_42443,N_41668,N_41322);
nor U42444 (N_42444,N_41158,N_41558);
or U42445 (N_42445,N_41168,N_41232);
or U42446 (N_42446,N_41197,N_41853);
nand U42447 (N_42447,N_41889,N_41129);
xnor U42448 (N_42448,N_41928,N_41177);
nor U42449 (N_42449,N_41762,N_41013);
nand U42450 (N_42450,N_41242,N_41525);
and U42451 (N_42451,N_41684,N_41291);
xnor U42452 (N_42452,N_41994,N_41518);
or U42453 (N_42453,N_41873,N_41307);
nand U42454 (N_42454,N_41876,N_41350);
xor U42455 (N_42455,N_41098,N_41137);
nand U42456 (N_42456,N_41275,N_41124);
xor U42457 (N_42457,N_41407,N_41664);
or U42458 (N_42458,N_41633,N_41644);
xnor U42459 (N_42459,N_41931,N_41532);
xnor U42460 (N_42460,N_41058,N_41929);
nand U42461 (N_42461,N_41610,N_41349);
nor U42462 (N_42462,N_41432,N_41497);
nor U42463 (N_42463,N_41755,N_41807);
xnor U42464 (N_42464,N_41198,N_41572);
and U42465 (N_42465,N_41444,N_41983);
xor U42466 (N_42466,N_41973,N_41377);
or U42467 (N_42467,N_41697,N_41157);
nand U42468 (N_42468,N_41781,N_41255);
and U42469 (N_42469,N_41386,N_41573);
xor U42470 (N_42470,N_41114,N_41118);
and U42471 (N_42471,N_41660,N_41535);
nand U42472 (N_42472,N_41845,N_41319);
xor U42473 (N_42473,N_41998,N_41471);
xor U42474 (N_42474,N_41812,N_41134);
and U42475 (N_42475,N_41367,N_41990);
xor U42476 (N_42476,N_41072,N_41613);
and U42477 (N_42477,N_41110,N_41677);
and U42478 (N_42478,N_41164,N_41012);
nand U42479 (N_42479,N_41556,N_41415);
xor U42480 (N_42480,N_41583,N_41975);
and U42481 (N_42481,N_41960,N_41952);
nand U42482 (N_42482,N_41295,N_41949);
nand U42483 (N_42483,N_41126,N_41352);
xor U42484 (N_42484,N_41611,N_41822);
nand U42485 (N_42485,N_41226,N_41524);
xor U42486 (N_42486,N_41183,N_41450);
nor U42487 (N_42487,N_41368,N_41490);
nand U42488 (N_42488,N_41840,N_41472);
xnor U42489 (N_42489,N_41396,N_41231);
or U42490 (N_42490,N_41031,N_41094);
and U42491 (N_42491,N_41005,N_41266);
nand U42492 (N_42492,N_41897,N_41740);
xor U42493 (N_42493,N_41742,N_41540);
and U42494 (N_42494,N_41842,N_41606);
or U42495 (N_42495,N_41219,N_41786);
nor U42496 (N_42496,N_41776,N_41313);
and U42497 (N_42497,N_41587,N_41286);
nor U42498 (N_42498,N_41751,N_41719);
or U42499 (N_42499,N_41585,N_41378);
or U42500 (N_42500,N_41737,N_41868);
nor U42501 (N_42501,N_41277,N_41592);
nor U42502 (N_42502,N_41908,N_41700);
nand U42503 (N_42503,N_41928,N_41776);
nor U42504 (N_42504,N_41705,N_41710);
nor U42505 (N_42505,N_41356,N_41103);
xor U42506 (N_42506,N_41526,N_41313);
nand U42507 (N_42507,N_41442,N_41475);
nand U42508 (N_42508,N_41311,N_41101);
xnor U42509 (N_42509,N_41555,N_41571);
nor U42510 (N_42510,N_41655,N_41656);
or U42511 (N_42511,N_41730,N_41992);
and U42512 (N_42512,N_41350,N_41326);
nor U42513 (N_42513,N_41934,N_41884);
xor U42514 (N_42514,N_41885,N_41912);
xnor U42515 (N_42515,N_41525,N_41267);
nor U42516 (N_42516,N_41286,N_41802);
nor U42517 (N_42517,N_41461,N_41007);
or U42518 (N_42518,N_41216,N_41482);
nand U42519 (N_42519,N_41373,N_41485);
and U42520 (N_42520,N_41569,N_41796);
nand U42521 (N_42521,N_41163,N_41577);
nor U42522 (N_42522,N_41358,N_41732);
xnor U42523 (N_42523,N_41522,N_41432);
nor U42524 (N_42524,N_41321,N_41628);
nand U42525 (N_42525,N_41983,N_41541);
or U42526 (N_42526,N_41240,N_41687);
nor U42527 (N_42527,N_41236,N_41485);
and U42528 (N_42528,N_41101,N_41276);
and U42529 (N_42529,N_41942,N_41900);
and U42530 (N_42530,N_41158,N_41732);
nand U42531 (N_42531,N_41228,N_41669);
or U42532 (N_42532,N_41136,N_41420);
nand U42533 (N_42533,N_41077,N_41696);
nand U42534 (N_42534,N_41150,N_41670);
nor U42535 (N_42535,N_41596,N_41435);
nand U42536 (N_42536,N_41298,N_41840);
nand U42537 (N_42537,N_41280,N_41259);
xnor U42538 (N_42538,N_41902,N_41203);
nor U42539 (N_42539,N_41877,N_41624);
nor U42540 (N_42540,N_41979,N_41699);
xnor U42541 (N_42541,N_41394,N_41444);
nor U42542 (N_42542,N_41728,N_41568);
xor U42543 (N_42543,N_41138,N_41475);
nand U42544 (N_42544,N_41940,N_41510);
nand U42545 (N_42545,N_41479,N_41043);
nand U42546 (N_42546,N_41301,N_41498);
nor U42547 (N_42547,N_41303,N_41080);
and U42548 (N_42548,N_41991,N_41068);
nor U42549 (N_42549,N_41948,N_41543);
xor U42550 (N_42550,N_41683,N_41327);
nor U42551 (N_42551,N_41028,N_41723);
nor U42552 (N_42552,N_41503,N_41864);
xnor U42553 (N_42553,N_41597,N_41244);
nor U42554 (N_42554,N_41408,N_41452);
or U42555 (N_42555,N_41688,N_41679);
and U42556 (N_42556,N_41906,N_41316);
and U42557 (N_42557,N_41379,N_41820);
or U42558 (N_42558,N_41955,N_41673);
and U42559 (N_42559,N_41037,N_41626);
nor U42560 (N_42560,N_41533,N_41462);
and U42561 (N_42561,N_41117,N_41718);
nand U42562 (N_42562,N_41176,N_41959);
or U42563 (N_42563,N_41452,N_41933);
nand U42564 (N_42564,N_41226,N_41642);
xnor U42565 (N_42565,N_41821,N_41529);
and U42566 (N_42566,N_41973,N_41125);
and U42567 (N_42567,N_41447,N_41370);
or U42568 (N_42568,N_41506,N_41654);
nor U42569 (N_42569,N_41052,N_41225);
xnor U42570 (N_42570,N_41000,N_41526);
nor U42571 (N_42571,N_41936,N_41779);
nand U42572 (N_42572,N_41047,N_41037);
or U42573 (N_42573,N_41757,N_41093);
nor U42574 (N_42574,N_41433,N_41261);
and U42575 (N_42575,N_41919,N_41484);
nand U42576 (N_42576,N_41688,N_41183);
nor U42577 (N_42577,N_41572,N_41535);
nor U42578 (N_42578,N_41889,N_41714);
nand U42579 (N_42579,N_41697,N_41812);
nor U42580 (N_42580,N_41104,N_41958);
and U42581 (N_42581,N_41205,N_41671);
xor U42582 (N_42582,N_41150,N_41727);
and U42583 (N_42583,N_41637,N_41804);
nor U42584 (N_42584,N_41327,N_41393);
xor U42585 (N_42585,N_41808,N_41432);
nor U42586 (N_42586,N_41858,N_41754);
and U42587 (N_42587,N_41341,N_41954);
xor U42588 (N_42588,N_41021,N_41546);
xnor U42589 (N_42589,N_41817,N_41772);
and U42590 (N_42590,N_41015,N_41632);
or U42591 (N_42591,N_41698,N_41513);
or U42592 (N_42592,N_41952,N_41654);
and U42593 (N_42593,N_41416,N_41238);
and U42594 (N_42594,N_41171,N_41616);
and U42595 (N_42595,N_41027,N_41491);
nand U42596 (N_42596,N_41804,N_41579);
nand U42597 (N_42597,N_41056,N_41057);
xor U42598 (N_42598,N_41458,N_41992);
and U42599 (N_42599,N_41364,N_41965);
nand U42600 (N_42600,N_41959,N_41513);
nor U42601 (N_42601,N_41818,N_41956);
or U42602 (N_42602,N_41626,N_41492);
nand U42603 (N_42603,N_41541,N_41036);
or U42604 (N_42604,N_41778,N_41511);
and U42605 (N_42605,N_41900,N_41821);
and U42606 (N_42606,N_41271,N_41373);
nor U42607 (N_42607,N_41183,N_41212);
nand U42608 (N_42608,N_41531,N_41837);
and U42609 (N_42609,N_41173,N_41328);
nand U42610 (N_42610,N_41927,N_41509);
nor U42611 (N_42611,N_41710,N_41313);
nor U42612 (N_42612,N_41180,N_41124);
nand U42613 (N_42613,N_41507,N_41762);
nor U42614 (N_42614,N_41788,N_41443);
xnor U42615 (N_42615,N_41898,N_41017);
nor U42616 (N_42616,N_41058,N_41719);
and U42617 (N_42617,N_41290,N_41355);
or U42618 (N_42618,N_41876,N_41017);
and U42619 (N_42619,N_41529,N_41017);
and U42620 (N_42620,N_41090,N_41871);
nand U42621 (N_42621,N_41431,N_41594);
and U42622 (N_42622,N_41621,N_41511);
or U42623 (N_42623,N_41444,N_41975);
nor U42624 (N_42624,N_41941,N_41984);
xor U42625 (N_42625,N_41798,N_41045);
nor U42626 (N_42626,N_41964,N_41217);
and U42627 (N_42627,N_41189,N_41197);
and U42628 (N_42628,N_41250,N_41682);
or U42629 (N_42629,N_41791,N_41068);
or U42630 (N_42630,N_41289,N_41240);
or U42631 (N_42631,N_41940,N_41115);
and U42632 (N_42632,N_41768,N_41186);
xor U42633 (N_42633,N_41945,N_41932);
nand U42634 (N_42634,N_41676,N_41633);
and U42635 (N_42635,N_41372,N_41038);
and U42636 (N_42636,N_41718,N_41301);
and U42637 (N_42637,N_41329,N_41972);
nand U42638 (N_42638,N_41765,N_41810);
xnor U42639 (N_42639,N_41676,N_41640);
and U42640 (N_42640,N_41863,N_41059);
or U42641 (N_42641,N_41847,N_41070);
or U42642 (N_42642,N_41512,N_41734);
and U42643 (N_42643,N_41474,N_41336);
and U42644 (N_42644,N_41168,N_41824);
or U42645 (N_42645,N_41256,N_41818);
nor U42646 (N_42646,N_41685,N_41274);
xor U42647 (N_42647,N_41188,N_41877);
and U42648 (N_42648,N_41815,N_41650);
nand U42649 (N_42649,N_41769,N_41013);
nand U42650 (N_42650,N_41492,N_41618);
nand U42651 (N_42651,N_41264,N_41510);
nand U42652 (N_42652,N_41674,N_41595);
xor U42653 (N_42653,N_41841,N_41151);
xor U42654 (N_42654,N_41803,N_41030);
or U42655 (N_42655,N_41308,N_41522);
nor U42656 (N_42656,N_41430,N_41990);
nand U42657 (N_42657,N_41695,N_41006);
and U42658 (N_42658,N_41607,N_41931);
or U42659 (N_42659,N_41040,N_41049);
or U42660 (N_42660,N_41652,N_41567);
and U42661 (N_42661,N_41186,N_41249);
nand U42662 (N_42662,N_41825,N_41109);
and U42663 (N_42663,N_41946,N_41003);
and U42664 (N_42664,N_41457,N_41806);
nand U42665 (N_42665,N_41983,N_41041);
xor U42666 (N_42666,N_41200,N_41952);
xnor U42667 (N_42667,N_41060,N_41942);
or U42668 (N_42668,N_41108,N_41021);
xnor U42669 (N_42669,N_41214,N_41891);
and U42670 (N_42670,N_41898,N_41416);
nor U42671 (N_42671,N_41210,N_41666);
or U42672 (N_42672,N_41771,N_41691);
and U42673 (N_42673,N_41314,N_41883);
or U42674 (N_42674,N_41974,N_41724);
and U42675 (N_42675,N_41161,N_41959);
xnor U42676 (N_42676,N_41564,N_41581);
nor U42677 (N_42677,N_41772,N_41303);
xnor U42678 (N_42678,N_41810,N_41897);
and U42679 (N_42679,N_41709,N_41155);
nand U42680 (N_42680,N_41071,N_41845);
and U42681 (N_42681,N_41597,N_41290);
nand U42682 (N_42682,N_41377,N_41893);
nand U42683 (N_42683,N_41828,N_41417);
nand U42684 (N_42684,N_41374,N_41483);
nor U42685 (N_42685,N_41188,N_41369);
or U42686 (N_42686,N_41835,N_41645);
nor U42687 (N_42687,N_41214,N_41108);
nor U42688 (N_42688,N_41376,N_41862);
nand U42689 (N_42689,N_41218,N_41001);
or U42690 (N_42690,N_41973,N_41245);
xnor U42691 (N_42691,N_41648,N_41644);
and U42692 (N_42692,N_41237,N_41251);
xnor U42693 (N_42693,N_41885,N_41345);
xnor U42694 (N_42694,N_41474,N_41882);
and U42695 (N_42695,N_41270,N_41973);
xnor U42696 (N_42696,N_41806,N_41771);
xnor U42697 (N_42697,N_41169,N_41545);
nor U42698 (N_42698,N_41810,N_41544);
nor U42699 (N_42699,N_41622,N_41591);
nor U42700 (N_42700,N_41836,N_41970);
and U42701 (N_42701,N_41517,N_41674);
nand U42702 (N_42702,N_41596,N_41053);
xnor U42703 (N_42703,N_41269,N_41241);
nor U42704 (N_42704,N_41040,N_41707);
nor U42705 (N_42705,N_41951,N_41181);
nor U42706 (N_42706,N_41498,N_41228);
nor U42707 (N_42707,N_41226,N_41824);
nand U42708 (N_42708,N_41803,N_41365);
and U42709 (N_42709,N_41285,N_41123);
nor U42710 (N_42710,N_41866,N_41960);
xor U42711 (N_42711,N_41947,N_41890);
nand U42712 (N_42712,N_41410,N_41320);
and U42713 (N_42713,N_41683,N_41276);
and U42714 (N_42714,N_41016,N_41066);
nor U42715 (N_42715,N_41223,N_41168);
xnor U42716 (N_42716,N_41356,N_41179);
and U42717 (N_42717,N_41862,N_41727);
nand U42718 (N_42718,N_41886,N_41613);
xor U42719 (N_42719,N_41793,N_41751);
nor U42720 (N_42720,N_41274,N_41259);
xnor U42721 (N_42721,N_41652,N_41553);
and U42722 (N_42722,N_41049,N_41894);
nor U42723 (N_42723,N_41759,N_41259);
xor U42724 (N_42724,N_41165,N_41122);
or U42725 (N_42725,N_41382,N_41651);
nor U42726 (N_42726,N_41522,N_41379);
or U42727 (N_42727,N_41152,N_41237);
or U42728 (N_42728,N_41973,N_41707);
or U42729 (N_42729,N_41385,N_41958);
and U42730 (N_42730,N_41019,N_41926);
or U42731 (N_42731,N_41087,N_41593);
nor U42732 (N_42732,N_41686,N_41604);
or U42733 (N_42733,N_41784,N_41494);
and U42734 (N_42734,N_41472,N_41112);
nor U42735 (N_42735,N_41207,N_41205);
or U42736 (N_42736,N_41563,N_41375);
nand U42737 (N_42737,N_41058,N_41134);
xnor U42738 (N_42738,N_41747,N_41472);
or U42739 (N_42739,N_41068,N_41631);
and U42740 (N_42740,N_41739,N_41755);
or U42741 (N_42741,N_41167,N_41171);
xor U42742 (N_42742,N_41608,N_41491);
and U42743 (N_42743,N_41994,N_41863);
or U42744 (N_42744,N_41586,N_41728);
or U42745 (N_42745,N_41196,N_41814);
nand U42746 (N_42746,N_41585,N_41986);
nor U42747 (N_42747,N_41434,N_41973);
and U42748 (N_42748,N_41221,N_41807);
nor U42749 (N_42749,N_41252,N_41391);
and U42750 (N_42750,N_41789,N_41571);
xor U42751 (N_42751,N_41698,N_41581);
nand U42752 (N_42752,N_41300,N_41744);
or U42753 (N_42753,N_41201,N_41612);
xnor U42754 (N_42754,N_41295,N_41951);
or U42755 (N_42755,N_41722,N_41224);
nand U42756 (N_42756,N_41269,N_41331);
xor U42757 (N_42757,N_41645,N_41284);
and U42758 (N_42758,N_41656,N_41446);
and U42759 (N_42759,N_41632,N_41566);
nand U42760 (N_42760,N_41272,N_41887);
and U42761 (N_42761,N_41645,N_41339);
nand U42762 (N_42762,N_41423,N_41402);
or U42763 (N_42763,N_41512,N_41968);
nand U42764 (N_42764,N_41781,N_41344);
nand U42765 (N_42765,N_41687,N_41702);
or U42766 (N_42766,N_41303,N_41523);
xnor U42767 (N_42767,N_41850,N_41283);
nand U42768 (N_42768,N_41503,N_41463);
xor U42769 (N_42769,N_41415,N_41337);
xnor U42770 (N_42770,N_41660,N_41945);
nor U42771 (N_42771,N_41548,N_41648);
and U42772 (N_42772,N_41417,N_41480);
nand U42773 (N_42773,N_41214,N_41348);
and U42774 (N_42774,N_41792,N_41599);
or U42775 (N_42775,N_41291,N_41666);
nand U42776 (N_42776,N_41827,N_41069);
xnor U42777 (N_42777,N_41618,N_41327);
and U42778 (N_42778,N_41994,N_41178);
and U42779 (N_42779,N_41170,N_41607);
and U42780 (N_42780,N_41036,N_41903);
xor U42781 (N_42781,N_41089,N_41057);
or U42782 (N_42782,N_41730,N_41044);
xnor U42783 (N_42783,N_41768,N_41526);
nor U42784 (N_42784,N_41562,N_41794);
and U42785 (N_42785,N_41705,N_41381);
nand U42786 (N_42786,N_41374,N_41683);
nand U42787 (N_42787,N_41114,N_41919);
and U42788 (N_42788,N_41823,N_41622);
xnor U42789 (N_42789,N_41981,N_41531);
nor U42790 (N_42790,N_41464,N_41324);
or U42791 (N_42791,N_41689,N_41731);
and U42792 (N_42792,N_41007,N_41888);
xnor U42793 (N_42793,N_41733,N_41215);
and U42794 (N_42794,N_41580,N_41459);
xor U42795 (N_42795,N_41743,N_41056);
nand U42796 (N_42796,N_41489,N_41394);
nor U42797 (N_42797,N_41131,N_41583);
xor U42798 (N_42798,N_41976,N_41417);
and U42799 (N_42799,N_41776,N_41018);
and U42800 (N_42800,N_41605,N_41579);
xnor U42801 (N_42801,N_41065,N_41962);
and U42802 (N_42802,N_41563,N_41715);
nor U42803 (N_42803,N_41456,N_41256);
xor U42804 (N_42804,N_41503,N_41466);
nor U42805 (N_42805,N_41558,N_41930);
xor U42806 (N_42806,N_41888,N_41621);
nor U42807 (N_42807,N_41784,N_41999);
nand U42808 (N_42808,N_41670,N_41818);
xnor U42809 (N_42809,N_41643,N_41475);
nor U42810 (N_42810,N_41098,N_41677);
and U42811 (N_42811,N_41410,N_41584);
xor U42812 (N_42812,N_41435,N_41212);
or U42813 (N_42813,N_41991,N_41453);
nor U42814 (N_42814,N_41413,N_41552);
or U42815 (N_42815,N_41591,N_41389);
and U42816 (N_42816,N_41564,N_41761);
nand U42817 (N_42817,N_41503,N_41879);
and U42818 (N_42818,N_41667,N_41558);
xor U42819 (N_42819,N_41698,N_41177);
nand U42820 (N_42820,N_41770,N_41582);
nand U42821 (N_42821,N_41623,N_41074);
and U42822 (N_42822,N_41826,N_41691);
or U42823 (N_42823,N_41553,N_41596);
xnor U42824 (N_42824,N_41704,N_41896);
and U42825 (N_42825,N_41967,N_41790);
nand U42826 (N_42826,N_41872,N_41779);
or U42827 (N_42827,N_41314,N_41900);
nand U42828 (N_42828,N_41294,N_41094);
nand U42829 (N_42829,N_41653,N_41077);
xor U42830 (N_42830,N_41788,N_41757);
xor U42831 (N_42831,N_41580,N_41369);
or U42832 (N_42832,N_41278,N_41387);
and U42833 (N_42833,N_41432,N_41026);
nand U42834 (N_42834,N_41758,N_41812);
and U42835 (N_42835,N_41537,N_41013);
or U42836 (N_42836,N_41346,N_41581);
nor U42837 (N_42837,N_41793,N_41828);
nor U42838 (N_42838,N_41576,N_41378);
nand U42839 (N_42839,N_41244,N_41365);
or U42840 (N_42840,N_41346,N_41774);
xnor U42841 (N_42841,N_41341,N_41640);
nand U42842 (N_42842,N_41702,N_41860);
and U42843 (N_42843,N_41166,N_41488);
or U42844 (N_42844,N_41714,N_41171);
nor U42845 (N_42845,N_41644,N_41609);
nand U42846 (N_42846,N_41368,N_41399);
nor U42847 (N_42847,N_41634,N_41953);
and U42848 (N_42848,N_41902,N_41150);
nand U42849 (N_42849,N_41113,N_41437);
or U42850 (N_42850,N_41301,N_41601);
and U42851 (N_42851,N_41460,N_41114);
and U42852 (N_42852,N_41902,N_41659);
xor U42853 (N_42853,N_41118,N_41868);
xor U42854 (N_42854,N_41397,N_41078);
nand U42855 (N_42855,N_41317,N_41587);
xnor U42856 (N_42856,N_41805,N_41996);
nor U42857 (N_42857,N_41912,N_41853);
nand U42858 (N_42858,N_41179,N_41813);
nand U42859 (N_42859,N_41887,N_41691);
nand U42860 (N_42860,N_41566,N_41613);
nand U42861 (N_42861,N_41218,N_41000);
nor U42862 (N_42862,N_41048,N_41196);
nand U42863 (N_42863,N_41417,N_41655);
xor U42864 (N_42864,N_41722,N_41195);
or U42865 (N_42865,N_41645,N_41431);
nor U42866 (N_42866,N_41202,N_41824);
xor U42867 (N_42867,N_41356,N_41157);
nand U42868 (N_42868,N_41694,N_41501);
or U42869 (N_42869,N_41872,N_41348);
and U42870 (N_42870,N_41250,N_41048);
or U42871 (N_42871,N_41413,N_41862);
nor U42872 (N_42872,N_41369,N_41502);
and U42873 (N_42873,N_41671,N_41281);
nor U42874 (N_42874,N_41400,N_41343);
nand U42875 (N_42875,N_41203,N_41601);
and U42876 (N_42876,N_41402,N_41435);
nor U42877 (N_42877,N_41203,N_41709);
xor U42878 (N_42878,N_41553,N_41620);
or U42879 (N_42879,N_41788,N_41028);
nor U42880 (N_42880,N_41347,N_41720);
nor U42881 (N_42881,N_41513,N_41941);
nand U42882 (N_42882,N_41777,N_41757);
xnor U42883 (N_42883,N_41632,N_41912);
and U42884 (N_42884,N_41986,N_41229);
xnor U42885 (N_42885,N_41366,N_41054);
xnor U42886 (N_42886,N_41040,N_41470);
nand U42887 (N_42887,N_41237,N_41334);
nand U42888 (N_42888,N_41413,N_41207);
or U42889 (N_42889,N_41898,N_41118);
xor U42890 (N_42890,N_41671,N_41498);
and U42891 (N_42891,N_41431,N_41928);
and U42892 (N_42892,N_41984,N_41172);
and U42893 (N_42893,N_41459,N_41058);
nand U42894 (N_42894,N_41980,N_41617);
nor U42895 (N_42895,N_41962,N_41609);
nor U42896 (N_42896,N_41491,N_41578);
and U42897 (N_42897,N_41048,N_41280);
and U42898 (N_42898,N_41724,N_41371);
nand U42899 (N_42899,N_41319,N_41347);
nand U42900 (N_42900,N_41551,N_41766);
or U42901 (N_42901,N_41954,N_41355);
nand U42902 (N_42902,N_41116,N_41780);
nor U42903 (N_42903,N_41657,N_41186);
nor U42904 (N_42904,N_41217,N_41607);
xnor U42905 (N_42905,N_41374,N_41848);
and U42906 (N_42906,N_41505,N_41883);
or U42907 (N_42907,N_41265,N_41916);
nor U42908 (N_42908,N_41009,N_41659);
xor U42909 (N_42909,N_41022,N_41052);
nand U42910 (N_42910,N_41310,N_41510);
or U42911 (N_42911,N_41024,N_41591);
nand U42912 (N_42912,N_41141,N_41574);
or U42913 (N_42913,N_41410,N_41909);
xor U42914 (N_42914,N_41537,N_41090);
or U42915 (N_42915,N_41908,N_41127);
or U42916 (N_42916,N_41820,N_41935);
and U42917 (N_42917,N_41220,N_41790);
or U42918 (N_42918,N_41997,N_41021);
or U42919 (N_42919,N_41335,N_41207);
or U42920 (N_42920,N_41092,N_41165);
nor U42921 (N_42921,N_41694,N_41508);
nand U42922 (N_42922,N_41214,N_41987);
nand U42923 (N_42923,N_41625,N_41056);
nor U42924 (N_42924,N_41508,N_41953);
xnor U42925 (N_42925,N_41856,N_41177);
nor U42926 (N_42926,N_41181,N_41674);
and U42927 (N_42927,N_41734,N_41272);
and U42928 (N_42928,N_41704,N_41009);
nand U42929 (N_42929,N_41220,N_41044);
and U42930 (N_42930,N_41266,N_41527);
and U42931 (N_42931,N_41557,N_41188);
nand U42932 (N_42932,N_41633,N_41092);
xnor U42933 (N_42933,N_41311,N_41918);
xor U42934 (N_42934,N_41310,N_41786);
or U42935 (N_42935,N_41397,N_41879);
or U42936 (N_42936,N_41471,N_41938);
nand U42937 (N_42937,N_41690,N_41619);
nor U42938 (N_42938,N_41543,N_41068);
xnor U42939 (N_42939,N_41798,N_41038);
nor U42940 (N_42940,N_41176,N_41593);
or U42941 (N_42941,N_41123,N_41645);
nor U42942 (N_42942,N_41451,N_41022);
or U42943 (N_42943,N_41904,N_41283);
and U42944 (N_42944,N_41082,N_41727);
xor U42945 (N_42945,N_41865,N_41729);
nor U42946 (N_42946,N_41456,N_41224);
and U42947 (N_42947,N_41123,N_41996);
nor U42948 (N_42948,N_41255,N_41991);
or U42949 (N_42949,N_41662,N_41181);
and U42950 (N_42950,N_41314,N_41784);
or U42951 (N_42951,N_41900,N_41965);
nand U42952 (N_42952,N_41003,N_41566);
or U42953 (N_42953,N_41976,N_41613);
nand U42954 (N_42954,N_41724,N_41538);
and U42955 (N_42955,N_41939,N_41116);
nor U42956 (N_42956,N_41833,N_41391);
xor U42957 (N_42957,N_41480,N_41754);
nand U42958 (N_42958,N_41389,N_41442);
xor U42959 (N_42959,N_41197,N_41720);
xnor U42960 (N_42960,N_41529,N_41738);
and U42961 (N_42961,N_41380,N_41807);
and U42962 (N_42962,N_41194,N_41645);
nor U42963 (N_42963,N_41027,N_41053);
nand U42964 (N_42964,N_41745,N_41333);
nand U42965 (N_42965,N_41014,N_41884);
or U42966 (N_42966,N_41788,N_41546);
nor U42967 (N_42967,N_41157,N_41519);
and U42968 (N_42968,N_41710,N_41299);
xor U42969 (N_42969,N_41759,N_41865);
xnor U42970 (N_42970,N_41979,N_41854);
nor U42971 (N_42971,N_41514,N_41266);
or U42972 (N_42972,N_41507,N_41766);
and U42973 (N_42973,N_41659,N_41126);
and U42974 (N_42974,N_41714,N_41008);
nor U42975 (N_42975,N_41833,N_41933);
nand U42976 (N_42976,N_41471,N_41146);
and U42977 (N_42977,N_41858,N_41606);
nor U42978 (N_42978,N_41910,N_41206);
xor U42979 (N_42979,N_41410,N_41745);
or U42980 (N_42980,N_41916,N_41960);
nand U42981 (N_42981,N_41333,N_41588);
nor U42982 (N_42982,N_41693,N_41139);
xnor U42983 (N_42983,N_41130,N_41947);
or U42984 (N_42984,N_41101,N_41467);
xnor U42985 (N_42985,N_41415,N_41582);
xnor U42986 (N_42986,N_41060,N_41171);
xor U42987 (N_42987,N_41580,N_41154);
nor U42988 (N_42988,N_41289,N_41840);
and U42989 (N_42989,N_41955,N_41138);
and U42990 (N_42990,N_41807,N_41438);
or U42991 (N_42991,N_41722,N_41031);
nand U42992 (N_42992,N_41046,N_41407);
and U42993 (N_42993,N_41705,N_41978);
nor U42994 (N_42994,N_41409,N_41436);
and U42995 (N_42995,N_41819,N_41308);
nor U42996 (N_42996,N_41528,N_41402);
nand U42997 (N_42997,N_41043,N_41020);
xnor U42998 (N_42998,N_41118,N_41595);
nand U42999 (N_42999,N_41300,N_41702);
nor U43000 (N_43000,N_42485,N_42583);
xnor U43001 (N_43001,N_42584,N_42338);
nand U43002 (N_43002,N_42650,N_42088);
nand U43003 (N_43003,N_42502,N_42100);
xor U43004 (N_43004,N_42531,N_42856);
xnor U43005 (N_43005,N_42169,N_42077);
or U43006 (N_43006,N_42179,N_42678);
xor U43007 (N_43007,N_42075,N_42599);
xor U43008 (N_43008,N_42807,N_42339);
and U43009 (N_43009,N_42649,N_42398);
or U43010 (N_43010,N_42023,N_42539);
nor U43011 (N_43011,N_42285,N_42298);
or U43012 (N_43012,N_42775,N_42747);
xor U43013 (N_43013,N_42853,N_42358);
nand U43014 (N_43014,N_42361,N_42598);
nor U43015 (N_43015,N_42756,N_42282);
nor U43016 (N_43016,N_42306,N_42659);
nand U43017 (N_43017,N_42810,N_42034);
nor U43018 (N_43018,N_42102,N_42990);
nand U43019 (N_43019,N_42039,N_42803);
and U43020 (N_43020,N_42692,N_42363);
and U43021 (N_43021,N_42580,N_42195);
xnor U43022 (N_43022,N_42537,N_42800);
nand U43023 (N_43023,N_42593,N_42629);
xor U43024 (N_43024,N_42001,N_42210);
nand U43025 (N_43025,N_42809,N_42496);
nand U43026 (N_43026,N_42595,N_42746);
and U43027 (N_43027,N_42569,N_42574);
nor U43028 (N_43028,N_42324,N_42229);
xnor U43029 (N_43029,N_42737,N_42357);
and U43030 (N_43030,N_42846,N_42707);
and U43031 (N_43031,N_42082,N_42283);
or U43032 (N_43032,N_42095,N_42049);
or U43033 (N_43033,N_42070,N_42880);
xor U43034 (N_43034,N_42723,N_42474);
xor U43035 (N_43035,N_42771,N_42783);
nand U43036 (N_43036,N_42196,N_42187);
and U43037 (N_43037,N_42867,N_42011);
xnor U43038 (N_43038,N_42828,N_42063);
nand U43039 (N_43039,N_42612,N_42287);
nand U43040 (N_43040,N_42183,N_42958);
xnor U43041 (N_43041,N_42036,N_42774);
xor U43042 (N_43042,N_42142,N_42256);
nor U43043 (N_43043,N_42516,N_42206);
and U43044 (N_43044,N_42136,N_42762);
or U43045 (N_43045,N_42244,N_42547);
and U43046 (N_43046,N_42526,N_42207);
or U43047 (N_43047,N_42676,N_42121);
nand U43048 (N_43048,N_42727,N_42975);
nand U43049 (N_43049,N_42223,N_42441);
nor U43050 (N_43050,N_42850,N_42632);
xor U43051 (N_43051,N_42563,N_42590);
xor U43052 (N_43052,N_42277,N_42482);
nor U43053 (N_43053,N_42388,N_42909);
xor U43054 (N_43054,N_42211,N_42227);
xor U43055 (N_43055,N_42717,N_42232);
and U43056 (N_43056,N_42438,N_42863);
and U43057 (N_43057,N_42180,N_42240);
xnor U43058 (N_43058,N_42213,N_42585);
or U43059 (N_43059,N_42830,N_42381);
xor U43060 (N_43060,N_42926,N_42416);
xnor U43061 (N_43061,N_42780,N_42307);
nor U43062 (N_43062,N_42760,N_42146);
nor U43063 (N_43063,N_42950,N_42076);
xor U43064 (N_43064,N_42586,N_42564);
and U43065 (N_43065,N_42041,N_42020);
or U43066 (N_43066,N_42899,N_42665);
xor U43067 (N_43067,N_42607,N_42739);
nor U43068 (N_43068,N_42512,N_42645);
xnor U43069 (N_43069,N_42522,N_42708);
xnor U43070 (N_43070,N_42370,N_42423);
and U43071 (N_43071,N_42006,N_42059);
nand U43072 (N_43072,N_42888,N_42552);
nand U43073 (N_43073,N_42509,N_42394);
nor U43074 (N_43074,N_42241,N_42004);
xor U43075 (N_43075,N_42166,N_42107);
nand U43076 (N_43076,N_42966,N_42532);
or U43077 (N_43077,N_42353,N_42060);
nand U43078 (N_43078,N_42015,N_42410);
xor U43079 (N_43079,N_42905,N_42725);
xnor U43080 (N_43080,N_42029,N_42164);
nand U43081 (N_43081,N_42677,N_42731);
xnor U43082 (N_43082,N_42127,N_42979);
or U43083 (N_43083,N_42745,N_42973);
or U43084 (N_43084,N_42843,N_42981);
xor U43085 (N_43085,N_42911,N_42631);
and U43086 (N_43086,N_42705,N_42500);
or U43087 (N_43087,N_42231,N_42667);
and U43088 (N_43088,N_42953,N_42640);
xor U43089 (N_43089,N_42845,N_42663);
xnor U43090 (N_43090,N_42831,N_42654);
and U43091 (N_43091,N_42889,N_42009);
or U43092 (N_43092,N_42835,N_42691);
nand U43093 (N_43093,N_42426,N_42260);
nand U43094 (N_43094,N_42616,N_42092);
or U43095 (N_43095,N_42924,N_42093);
and U43096 (N_43096,N_42556,N_42327);
or U43097 (N_43097,N_42212,N_42468);
nand U43098 (N_43098,N_42804,N_42073);
nand U43099 (N_43099,N_42637,N_42085);
or U43100 (N_43100,N_42523,N_42711);
or U43101 (N_43101,N_42340,N_42840);
and U43102 (N_43102,N_42550,N_42842);
xnor U43103 (N_43103,N_42535,N_42790);
xnor U43104 (N_43104,N_42252,N_42996);
nor U43105 (N_43105,N_42238,N_42904);
nor U43106 (N_43106,N_42561,N_42209);
or U43107 (N_43107,N_42787,N_42669);
xnor U43108 (N_43108,N_42626,N_42396);
nor U43109 (N_43109,N_42744,N_42837);
xor U43110 (N_43110,N_42280,N_42754);
xor U43111 (N_43111,N_42977,N_42215);
and U43112 (N_43112,N_42995,N_42314);
and U43113 (N_43113,N_42581,N_42055);
and U43114 (N_43114,N_42163,N_42944);
and U43115 (N_43115,N_42883,N_42477);
nor U43116 (N_43116,N_42302,N_42980);
and U43117 (N_43117,N_42778,N_42999);
nor U43118 (N_43118,N_42310,N_42934);
and U43119 (N_43119,N_42942,N_42655);
or U43120 (N_43120,N_42801,N_42770);
and U43121 (N_43121,N_42673,N_42434);
and U43122 (N_43122,N_42890,N_42696);
or U43123 (N_43123,N_42978,N_42007);
or U43124 (N_43124,N_42894,N_42040);
and U43125 (N_43125,N_42334,N_42752);
and U43126 (N_43126,N_42408,N_42750);
nor U43127 (N_43127,N_42317,N_42923);
nand U43128 (N_43128,N_42554,N_42194);
nor U43129 (N_43129,N_42757,N_42635);
xor U43130 (N_43130,N_42902,N_42335);
and U43131 (N_43131,N_42177,N_42559);
or U43132 (N_43132,N_42106,N_42524);
nor U43133 (N_43133,N_42562,N_42829);
and U43134 (N_43134,N_42299,N_42788);
nor U43135 (N_43135,N_42415,N_42019);
or U43136 (N_43136,N_42946,N_42495);
nand U43137 (N_43137,N_42724,N_42542);
nor U43138 (N_43138,N_42138,N_42797);
nor U43139 (N_43139,N_42035,N_42466);
or U43140 (N_43140,N_42808,N_42083);
or U43141 (N_43141,N_42568,N_42697);
or U43142 (N_43142,N_42638,N_42704);
xnor U43143 (N_43143,N_42687,N_42439);
nor U43144 (N_43144,N_42813,N_42467);
nor U43145 (N_43145,N_42453,N_42794);
and U43146 (N_43146,N_42118,N_42749);
xnor U43147 (N_43147,N_42816,N_42472);
or U43148 (N_43148,N_42375,N_42191);
nand U43149 (N_43149,N_42269,N_42938);
nor U43150 (N_43150,N_42008,N_42470);
nor U43151 (N_43151,N_42447,N_42651);
nand U43152 (N_43152,N_42906,N_42940);
xnor U43153 (N_43153,N_42090,N_42618);
or U43154 (N_43154,N_42119,N_42898);
and U43155 (N_43155,N_42456,N_42200);
or U43156 (N_43156,N_42819,N_42617);
and U43157 (N_43157,N_42917,N_42450);
or U43158 (N_43158,N_42235,N_42570);
and U43159 (N_43159,N_42189,N_42346);
or U43160 (N_43160,N_42862,N_42714);
and U43161 (N_43161,N_42684,N_42489);
xnor U43162 (N_43162,N_42887,N_42120);
xnor U43163 (N_43163,N_42814,N_42817);
and U43164 (N_43164,N_42219,N_42175);
nor U43165 (N_43165,N_42476,N_42367);
xor U43166 (N_43166,N_42094,N_42147);
xor U43167 (N_43167,N_42478,N_42767);
or U43168 (N_43168,N_42290,N_42185);
and U43169 (N_43169,N_42374,N_42379);
or U43170 (N_43170,N_42551,N_42326);
or U43171 (N_43171,N_42879,N_42462);
nand U43172 (N_43172,N_42832,N_42233);
nand U43173 (N_43173,N_42356,N_42251);
and U43174 (N_43174,N_42553,N_42544);
xnor U43175 (N_43175,N_42281,N_42258);
and U43176 (N_43176,N_42135,N_42224);
nor U43177 (N_43177,N_42857,N_42132);
xor U43178 (N_43178,N_42087,N_42647);
nor U43179 (N_43179,N_42504,N_42546);
nand U43180 (N_43180,N_42949,N_42886);
or U43181 (N_43181,N_42125,N_42855);
nor U43182 (N_43182,N_42877,N_42170);
nand U43183 (N_43183,N_42249,N_42266);
xor U43184 (N_43184,N_42936,N_42733);
or U43185 (N_43185,N_42974,N_42572);
or U43186 (N_43186,N_42262,N_42791);
nor U43187 (N_43187,N_42858,N_42261);
and U43188 (N_43188,N_42592,N_42751);
nand U43189 (N_43189,N_42080,N_42028);
nand U43190 (N_43190,N_42295,N_42014);
and U43191 (N_43191,N_42172,N_42997);
xor U43192 (N_43192,N_42480,N_42716);
nor U43193 (N_43193,N_42428,N_42989);
nand U43194 (N_43194,N_42141,N_42920);
xor U43195 (N_43195,N_42699,N_42452);
xnor U43196 (N_43196,N_42376,N_42168);
or U43197 (N_43197,N_42425,N_42827);
xnor U43198 (N_43198,N_42644,N_42518);
nor U43199 (N_43199,N_42341,N_42159);
or U43200 (N_43200,N_42613,N_42881);
xor U43201 (N_43201,N_42519,N_42893);
or U43202 (N_43202,N_42892,N_42962);
nor U43203 (N_43203,N_42648,N_42722);
or U43204 (N_43204,N_42854,N_42460);
or U43205 (N_43205,N_42037,N_42498);
xor U43206 (N_43206,N_42305,N_42225);
nand U43207 (N_43207,N_42091,N_42543);
xor U43208 (N_43208,N_42123,N_42250);
nand U43209 (N_43209,N_42027,N_42915);
or U43210 (N_43210,N_42994,N_42377);
nor U43211 (N_43211,N_42160,N_42510);
or U43212 (N_43212,N_42430,N_42401);
xnor U43213 (N_43213,N_42359,N_42329);
xnor U43214 (N_43214,N_42263,N_42922);
nor U43215 (N_43215,N_42397,N_42131);
nand U43216 (N_43216,N_42321,N_42276);
xor U43217 (N_43217,N_42018,N_42955);
nor U43218 (N_43218,N_42521,N_42758);
xnor U43219 (N_43219,N_42264,N_42390);
xnor U43220 (N_43220,N_42322,N_42411);
or U43221 (N_43221,N_42448,N_42735);
nand U43222 (N_43222,N_42391,N_42908);
nor U43223 (N_43223,N_42101,N_42715);
xor U43224 (N_43224,N_42957,N_42429);
nand U43225 (N_43225,N_42961,N_42424);
or U43226 (N_43226,N_42875,N_42186);
nand U43227 (N_43227,N_42952,N_42116);
and U43228 (N_43228,N_42701,N_42089);
xor U43229 (N_43229,N_42491,N_42308);
nor U43230 (N_43230,N_42935,N_42105);
xor U43231 (N_43231,N_42963,N_42151);
nand U43232 (N_43232,N_42442,N_42002);
nor U43233 (N_43233,N_42350,N_42702);
and U43234 (N_43234,N_42833,N_42078);
xor U43235 (N_43235,N_42668,N_42972);
and U43236 (N_43236,N_42712,N_42604);
and U43237 (N_43237,N_42108,N_42372);
and U43238 (N_43238,N_42721,N_42293);
or U43239 (N_43239,N_42204,N_42157);
and U43240 (N_43240,N_42245,N_42013);
or U43241 (N_43241,N_42203,N_42689);
nand U43242 (N_43242,N_42623,N_42565);
or U43243 (N_43243,N_42220,N_42865);
nand U43244 (N_43244,N_42181,N_42662);
or U43245 (N_43245,N_42190,N_42956);
and U43246 (N_43246,N_42866,N_42071);
nor U43247 (N_43247,N_42954,N_42440);
xnor U43248 (N_43248,N_42736,N_42560);
or U43249 (N_43249,N_42475,N_42919);
nand U43250 (N_43250,N_42992,N_42826);
and U43251 (N_43251,N_42382,N_42483);
or U43252 (N_43252,N_42624,N_42000);
xor U43253 (N_43253,N_42615,N_42834);
nor U43254 (N_43254,N_42536,N_42901);
nand U43255 (N_43255,N_42825,N_42571);
nor U43256 (N_43256,N_42362,N_42921);
or U43257 (N_43257,N_42449,N_42230);
and U43258 (N_43258,N_42603,N_42948);
and U43259 (N_43259,N_42349,N_42084);
nor U43260 (N_43260,N_42386,N_42454);
or U43261 (N_43261,N_42680,N_42109);
or U43262 (N_43262,N_42968,N_42548);
and U43263 (N_43263,N_42741,N_42383);
or U43264 (N_43264,N_42032,N_42418);
nand U43265 (N_43265,N_42369,N_42311);
xor U43266 (N_43266,N_42520,N_42690);
nor U43267 (N_43267,N_42998,N_42218);
nand U43268 (N_43268,N_42812,N_42871);
xor U43269 (N_43269,N_42884,N_42785);
nand U43270 (N_43270,N_42636,N_42026);
nand U43271 (N_43271,N_42852,N_42066);
and U43272 (N_43272,N_42103,N_42214);
xor U43273 (N_43273,N_42967,N_42044);
xnor U43274 (N_43274,N_42755,N_42567);
nand U43275 (N_43275,N_42288,N_42294);
xnor U43276 (N_43276,N_42621,N_42471);
nand U43277 (N_43277,N_42903,N_42822);
or U43278 (N_43278,N_42844,N_42096);
and U43279 (N_43279,N_42399,N_42937);
or U43280 (N_43280,N_42303,N_42683);
nand U43281 (N_43281,N_42660,N_42487);
or U43282 (N_43282,N_42664,N_42117);
nand U43283 (N_43283,N_42505,N_42301);
nor U43284 (N_43284,N_42533,N_42336);
xnor U43285 (N_43285,N_42389,N_42300);
nand U43286 (N_43286,N_42291,N_42703);
xnor U43287 (N_43287,N_42575,N_42150);
xor U43288 (N_43288,N_42777,N_42464);
nor U43289 (N_43289,N_42184,N_42010);
nand U43290 (N_43290,N_42639,N_42292);
xor U43291 (N_43291,N_42182,N_42868);
nor U43292 (N_43292,N_42304,N_42201);
xor U43293 (N_43293,N_42134,N_42404);
and U43294 (N_43294,N_42316,N_42422);
or U43295 (N_43295,N_42759,N_42538);
or U43296 (N_43296,N_42016,N_42473);
nand U43297 (N_43297,N_42602,N_42786);
and U43298 (N_43298,N_42985,N_42065);
nand U43299 (N_43299,N_42368,N_42588);
nor U43300 (N_43300,N_42236,N_42895);
xor U43301 (N_43301,N_42242,N_42685);
nor U43302 (N_43302,N_42156,N_42445);
and U43303 (N_43303,N_42743,N_42634);
nand U43304 (N_43304,N_42419,N_42969);
and U43305 (N_43305,N_42661,N_42870);
nor U43306 (N_43306,N_42038,N_42821);
and U43307 (N_43307,N_42221,N_42130);
nor U43308 (N_43308,N_42666,N_42074);
xor U43309 (N_43309,N_42140,N_42900);
xnor U43310 (N_43310,N_42882,N_42497);
nand U43311 (N_43311,N_42319,N_42328);
nor U43312 (N_43312,N_42433,N_42713);
or U43313 (N_43313,N_42932,N_42686);
xnor U43314 (N_43314,N_42848,N_42628);
or U43315 (N_43315,N_42400,N_42601);
or U43316 (N_43316,N_42481,N_42597);
and U43317 (N_43317,N_42270,N_42811);
nand U43318 (N_43318,N_42799,N_42492);
nand U43319 (N_43319,N_42838,N_42005);
xor U43320 (N_43320,N_42081,N_42987);
or U43321 (N_43321,N_42594,N_42048);
or U43322 (N_43322,N_42403,N_42047);
xor U43323 (N_43323,N_42323,N_42407);
xor U43324 (N_43324,N_42630,N_42124);
nand U43325 (N_43325,N_42046,N_42499);
or U43326 (N_43326,N_42941,N_42247);
xor U43327 (N_43327,N_42534,N_42062);
xnor U43328 (N_43328,N_42022,N_42337);
and U43329 (N_43329,N_42494,N_42729);
nand U43330 (N_43330,N_42781,N_42289);
xnor U43331 (N_43331,N_42993,N_42782);
nor U43332 (N_43332,N_42054,N_42061);
xnor U43333 (N_43333,N_42351,N_42173);
and U43334 (N_43334,N_42576,N_42625);
and U43335 (N_43335,N_42947,N_42162);
nand U43336 (N_43336,N_42964,N_42058);
xnor U43337 (N_43337,N_42874,N_42086);
xor U43338 (N_43338,N_42508,N_42600);
or U43339 (N_43339,N_42573,N_42710);
and U43340 (N_43340,N_42675,N_42943);
xor U43341 (N_43341,N_42525,N_42719);
or U43342 (N_43342,N_42239,N_42610);
xor U43343 (N_43343,N_42860,N_42682);
or U43344 (N_43344,N_42951,N_42414);
nand U43345 (N_43345,N_42851,N_42587);
or U43346 (N_43346,N_42405,N_42158);
and U43347 (N_43347,N_42469,N_42620);
or U43348 (N_43348,N_42929,N_42726);
nor U43349 (N_43349,N_42412,N_42017);
or U43350 (N_43350,N_42769,N_42693);
xnor U43351 (N_43351,N_42313,N_42137);
and U43352 (N_43352,N_42861,N_42393);
xor U43353 (N_43353,N_42067,N_42557);
nor U43354 (N_43354,N_42272,N_42217);
and U43355 (N_43355,N_42273,N_42366);
or U43356 (N_43356,N_42776,N_42384);
and U43357 (N_43357,N_42872,N_42965);
xnor U43358 (N_43358,N_42694,N_42152);
or U43359 (N_43359,N_42823,N_42795);
or U43360 (N_43360,N_42171,N_42789);
or U43361 (N_43361,N_42918,N_42344);
and U43362 (N_43362,N_42216,N_42873);
nand U43363 (N_43363,N_42596,N_42188);
xor U43364 (N_43364,N_42064,N_42925);
or U43365 (N_43365,N_42458,N_42698);
and U43366 (N_43366,N_42145,N_42939);
or U43367 (N_43367,N_42154,N_42761);
xnor U43368 (N_43368,N_42488,N_42378);
and U43369 (N_43369,N_42199,N_42354);
nand U43370 (N_43370,N_42982,N_42578);
and U43371 (N_43371,N_42459,N_42540);
and U43372 (N_43372,N_42779,N_42228);
nor U43373 (N_43373,N_42332,N_42527);
nor U43374 (N_43374,N_42253,N_42237);
nand U43375 (N_43375,N_42988,N_42633);
xor U43376 (N_43376,N_42406,N_42766);
or U43377 (N_43377,N_42461,N_42435);
nor U43378 (N_43378,N_42971,N_42312);
xor U43379 (N_43379,N_42333,N_42099);
and U43380 (N_43380,N_42457,N_42446);
nor U43381 (N_43381,N_42348,N_42805);
nor U43382 (N_43382,N_42986,N_42806);
and U43383 (N_43383,N_42773,N_42984);
nand U43384 (N_43384,N_42222,N_42202);
nand U43385 (N_43385,N_42342,N_42234);
or U43386 (N_43386,N_42068,N_42345);
and U43387 (N_43387,N_42279,N_42197);
nor U43388 (N_43388,N_42748,N_42591);
nand U43389 (N_43389,N_42174,N_42579);
nand U43390 (N_43390,N_42796,N_42331);
nand U43391 (N_43391,N_42318,N_42490);
nand U43392 (N_43392,N_42364,N_42432);
xor U43393 (N_43393,N_42259,N_42128);
or U43394 (N_43394,N_42133,N_42529);
xnor U43395 (N_43395,N_42891,N_42515);
or U43396 (N_43396,N_42657,N_42143);
nand U43397 (N_43397,N_42149,N_42614);
nand U43398 (N_43398,N_42056,N_42286);
nor U43399 (N_43399,N_42097,N_42802);
nor U43400 (N_43400,N_42330,N_42641);
nor U43401 (N_43401,N_42878,N_42841);
nand U43402 (N_43402,N_42025,N_42864);
or U43403 (N_43403,N_42511,N_42609);
nand U43404 (N_43404,N_42153,N_42051);
nor U43405 (N_43405,N_42380,N_42465);
xor U43406 (N_43406,N_42869,N_42024);
nor U43407 (N_43407,N_42325,N_42320);
nor U43408 (N_43408,N_42192,N_42126);
nor U43409 (N_43409,N_42976,N_42420);
nor U43410 (N_43410,N_42653,N_42764);
xor U43411 (N_43411,N_42528,N_42437);
and U43412 (N_43412,N_42385,N_42730);
xor U43413 (N_43413,N_42114,N_42658);
xnor U43414 (N_43414,N_42387,N_42506);
xnor U43415 (N_43415,N_42355,N_42672);
nand U43416 (N_43416,N_42818,N_42820);
nand U43417 (N_43417,N_42392,N_42983);
nor U43418 (N_43418,N_42144,N_42098);
xor U43419 (N_43419,N_42836,N_42611);
or U43420 (N_43420,N_42274,N_42254);
and U43421 (N_43421,N_42413,N_42284);
nor U43422 (N_43422,N_42267,N_42815);
xor U43423 (N_43423,N_42343,N_42265);
nand U43424 (N_43424,N_42960,N_42003);
xnor U43425 (N_43425,N_42656,N_42139);
xnor U43426 (N_43426,N_42930,N_42679);
nand U43427 (N_43427,N_42052,N_42031);
nor U43428 (N_43428,N_42627,N_42912);
nand U43429 (N_43429,N_42431,N_42129);
nand U43430 (N_43430,N_42352,N_42451);
nand U43431 (N_43431,N_42309,N_42885);
nand U43432 (N_43432,N_42057,N_42371);
and U43433 (N_43433,N_42582,N_42021);
xnor U43434 (N_43434,N_42069,N_42530);
nand U43435 (N_43435,N_42257,N_42916);
or U43436 (N_43436,N_42738,N_42155);
or U43437 (N_43437,N_42928,N_42360);
and U43438 (N_43438,N_42931,N_42275);
and U43439 (N_43439,N_42688,N_42577);
xnor U43440 (N_43440,N_42566,N_42501);
nor U43441 (N_43441,N_42896,N_42765);
and U43442 (N_43442,N_42053,N_42718);
nand U43443 (N_43443,N_42167,N_42112);
nor U43444 (N_43444,N_42670,N_42549);
nor U43445 (N_43445,N_42945,N_42763);
nor U43446 (N_43446,N_42728,N_42734);
nand U43447 (N_43447,N_42148,N_42178);
and U43448 (N_43448,N_42246,N_42605);
xnor U43449 (N_43449,N_42297,N_42784);
and U43450 (N_43450,N_42113,N_42910);
nand U43451 (N_43451,N_42296,N_42793);
nand U43452 (N_43452,N_42824,N_42427);
nor U43453 (N_43453,N_42643,N_42395);
nand U43454 (N_43454,N_42176,N_42111);
nor U43455 (N_43455,N_42205,N_42622);
nand U43456 (N_43456,N_42243,N_42674);
or U43457 (N_43457,N_42122,N_42161);
xor U43458 (N_43458,N_42507,N_42030);
xor U43459 (N_43459,N_42365,N_42646);
nor U43460 (N_43460,N_42642,N_42876);
nand U43461 (N_43461,N_42681,N_42991);
xnor U43462 (N_43462,N_42402,N_42315);
nor U43463 (N_43463,N_42706,N_42720);
or U43464 (N_43464,N_42732,N_42700);
nor U43465 (N_43465,N_42198,N_42619);
xor U43466 (N_43466,N_42479,N_42072);
nor U43467 (N_43467,N_42558,N_42042);
and U43468 (N_43468,N_42271,N_42859);
nor U43469 (N_43469,N_42933,N_42455);
or U43470 (N_43470,N_42045,N_42839);
nor U43471 (N_43471,N_42927,N_42493);
nor U43472 (N_43472,N_42347,N_42555);
nor U43473 (N_43473,N_42652,N_42268);
nand U43474 (N_43474,N_42443,N_42110);
or U43475 (N_43475,N_42671,N_42792);
nor U43476 (N_43476,N_42165,N_42104);
xnor U43477 (N_43477,N_42421,N_42849);
or U43478 (N_43478,N_42740,N_42248);
nor U43479 (N_43479,N_42514,N_42589);
xnor U43480 (N_43480,N_42417,N_42959);
or U43481 (N_43481,N_42772,N_42012);
nand U43482 (N_43482,N_42768,N_42517);
or U43483 (N_43483,N_42847,N_42050);
and U43484 (N_43484,N_42798,N_42115);
or U43485 (N_43485,N_42484,N_42914);
or U43486 (N_43486,N_42742,N_42913);
nor U43487 (N_43487,N_42463,N_42444);
nand U43488 (N_43488,N_42278,N_42436);
nor U43489 (N_43489,N_42970,N_42193);
or U43490 (N_43490,N_42907,N_42753);
nor U43491 (N_43491,N_42079,N_42695);
nand U43492 (N_43492,N_42541,N_42373);
nor U43493 (N_43493,N_42208,N_42608);
xor U43494 (N_43494,N_42226,N_42255);
nor U43495 (N_43495,N_42709,N_42606);
xor U43496 (N_43496,N_42897,N_42033);
nand U43497 (N_43497,N_42043,N_42486);
or U43498 (N_43498,N_42545,N_42503);
and U43499 (N_43499,N_42513,N_42409);
or U43500 (N_43500,N_42755,N_42558);
xor U43501 (N_43501,N_42883,N_42175);
nand U43502 (N_43502,N_42895,N_42625);
or U43503 (N_43503,N_42544,N_42898);
or U43504 (N_43504,N_42358,N_42413);
nor U43505 (N_43505,N_42910,N_42337);
xor U43506 (N_43506,N_42463,N_42541);
xor U43507 (N_43507,N_42491,N_42083);
and U43508 (N_43508,N_42105,N_42186);
xor U43509 (N_43509,N_42346,N_42671);
and U43510 (N_43510,N_42855,N_42549);
or U43511 (N_43511,N_42243,N_42941);
xor U43512 (N_43512,N_42190,N_42200);
or U43513 (N_43513,N_42727,N_42206);
or U43514 (N_43514,N_42370,N_42340);
and U43515 (N_43515,N_42536,N_42962);
and U43516 (N_43516,N_42266,N_42412);
or U43517 (N_43517,N_42234,N_42892);
nand U43518 (N_43518,N_42974,N_42118);
nor U43519 (N_43519,N_42145,N_42650);
nor U43520 (N_43520,N_42879,N_42436);
nand U43521 (N_43521,N_42202,N_42398);
nor U43522 (N_43522,N_42554,N_42519);
nand U43523 (N_43523,N_42633,N_42865);
xor U43524 (N_43524,N_42451,N_42344);
nand U43525 (N_43525,N_42418,N_42755);
nand U43526 (N_43526,N_42116,N_42769);
xor U43527 (N_43527,N_42482,N_42481);
and U43528 (N_43528,N_42542,N_42860);
nand U43529 (N_43529,N_42266,N_42885);
xor U43530 (N_43530,N_42174,N_42782);
nand U43531 (N_43531,N_42212,N_42324);
xor U43532 (N_43532,N_42999,N_42752);
or U43533 (N_43533,N_42189,N_42879);
and U43534 (N_43534,N_42774,N_42167);
and U43535 (N_43535,N_42435,N_42764);
and U43536 (N_43536,N_42187,N_42960);
and U43537 (N_43537,N_42924,N_42497);
nand U43538 (N_43538,N_42808,N_42980);
nor U43539 (N_43539,N_42936,N_42860);
nor U43540 (N_43540,N_42788,N_42759);
and U43541 (N_43541,N_42196,N_42986);
nor U43542 (N_43542,N_42618,N_42458);
xor U43543 (N_43543,N_42814,N_42919);
nor U43544 (N_43544,N_42054,N_42907);
xor U43545 (N_43545,N_42243,N_42196);
or U43546 (N_43546,N_42935,N_42752);
or U43547 (N_43547,N_42638,N_42199);
nand U43548 (N_43548,N_42219,N_42462);
nor U43549 (N_43549,N_42140,N_42068);
or U43550 (N_43550,N_42012,N_42144);
nor U43551 (N_43551,N_42263,N_42292);
or U43552 (N_43552,N_42751,N_42811);
or U43553 (N_43553,N_42423,N_42683);
or U43554 (N_43554,N_42651,N_42746);
nand U43555 (N_43555,N_42420,N_42741);
and U43556 (N_43556,N_42816,N_42296);
and U43557 (N_43557,N_42589,N_42342);
nor U43558 (N_43558,N_42074,N_42536);
xnor U43559 (N_43559,N_42032,N_42097);
nand U43560 (N_43560,N_42311,N_42716);
xnor U43561 (N_43561,N_42527,N_42725);
nor U43562 (N_43562,N_42871,N_42022);
nor U43563 (N_43563,N_42542,N_42157);
and U43564 (N_43564,N_42490,N_42822);
nand U43565 (N_43565,N_42197,N_42164);
xor U43566 (N_43566,N_42188,N_42168);
xor U43567 (N_43567,N_42168,N_42400);
xnor U43568 (N_43568,N_42583,N_42575);
nor U43569 (N_43569,N_42718,N_42512);
or U43570 (N_43570,N_42443,N_42475);
or U43571 (N_43571,N_42522,N_42091);
xor U43572 (N_43572,N_42121,N_42165);
or U43573 (N_43573,N_42638,N_42706);
and U43574 (N_43574,N_42640,N_42186);
and U43575 (N_43575,N_42384,N_42072);
nand U43576 (N_43576,N_42185,N_42131);
or U43577 (N_43577,N_42203,N_42327);
and U43578 (N_43578,N_42904,N_42938);
nor U43579 (N_43579,N_42883,N_42307);
and U43580 (N_43580,N_42928,N_42856);
xnor U43581 (N_43581,N_42524,N_42339);
or U43582 (N_43582,N_42300,N_42385);
and U43583 (N_43583,N_42747,N_42942);
nor U43584 (N_43584,N_42730,N_42097);
or U43585 (N_43585,N_42890,N_42374);
and U43586 (N_43586,N_42775,N_42748);
nand U43587 (N_43587,N_42327,N_42863);
xor U43588 (N_43588,N_42741,N_42629);
nand U43589 (N_43589,N_42246,N_42414);
or U43590 (N_43590,N_42559,N_42585);
or U43591 (N_43591,N_42931,N_42968);
nand U43592 (N_43592,N_42586,N_42512);
and U43593 (N_43593,N_42178,N_42447);
or U43594 (N_43594,N_42267,N_42036);
xnor U43595 (N_43595,N_42390,N_42270);
and U43596 (N_43596,N_42968,N_42825);
nor U43597 (N_43597,N_42399,N_42825);
nand U43598 (N_43598,N_42349,N_42970);
and U43599 (N_43599,N_42026,N_42295);
and U43600 (N_43600,N_42780,N_42525);
and U43601 (N_43601,N_42336,N_42452);
nand U43602 (N_43602,N_42369,N_42898);
and U43603 (N_43603,N_42521,N_42399);
nor U43604 (N_43604,N_42547,N_42768);
nor U43605 (N_43605,N_42683,N_42620);
or U43606 (N_43606,N_42596,N_42017);
nor U43607 (N_43607,N_42298,N_42618);
xnor U43608 (N_43608,N_42826,N_42303);
or U43609 (N_43609,N_42438,N_42857);
or U43610 (N_43610,N_42189,N_42562);
xor U43611 (N_43611,N_42007,N_42423);
or U43612 (N_43612,N_42806,N_42368);
nand U43613 (N_43613,N_42548,N_42470);
and U43614 (N_43614,N_42885,N_42045);
and U43615 (N_43615,N_42770,N_42214);
nor U43616 (N_43616,N_42924,N_42399);
and U43617 (N_43617,N_42621,N_42940);
xnor U43618 (N_43618,N_42719,N_42805);
and U43619 (N_43619,N_42289,N_42953);
and U43620 (N_43620,N_42228,N_42259);
nor U43621 (N_43621,N_42032,N_42525);
or U43622 (N_43622,N_42033,N_42458);
or U43623 (N_43623,N_42397,N_42702);
nand U43624 (N_43624,N_42081,N_42036);
or U43625 (N_43625,N_42168,N_42672);
nor U43626 (N_43626,N_42706,N_42508);
nor U43627 (N_43627,N_42021,N_42405);
xnor U43628 (N_43628,N_42155,N_42884);
and U43629 (N_43629,N_42590,N_42223);
or U43630 (N_43630,N_42676,N_42356);
nor U43631 (N_43631,N_42410,N_42436);
xnor U43632 (N_43632,N_42727,N_42676);
nor U43633 (N_43633,N_42881,N_42635);
xnor U43634 (N_43634,N_42765,N_42832);
nor U43635 (N_43635,N_42165,N_42687);
nor U43636 (N_43636,N_42060,N_42330);
or U43637 (N_43637,N_42147,N_42343);
nor U43638 (N_43638,N_42222,N_42961);
and U43639 (N_43639,N_42431,N_42972);
nor U43640 (N_43640,N_42601,N_42361);
nor U43641 (N_43641,N_42246,N_42864);
xor U43642 (N_43642,N_42728,N_42169);
xor U43643 (N_43643,N_42320,N_42931);
nand U43644 (N_43644,N_42613,N_42841);
xor U43645 (N_43645,N_42691,N_42565);
nand U43646 (N_43646,N_42278,N_42734);
or U43647 (N_43647,N_42101,N_42813);
xnor U43648 (N_43648,N_42857,N_42113);
or U43649 (N_43649,N_42296,N_42051);
xnor U43650 (N_43650,N_42345,N_42161);
xnor U43651 (N_43651,N_42016,N_42407);
nand U43652 (N_43652,N_42878,N_42127);
nand U43653 (N_43653,N_42797,N_42300);
or U43654 (N_43654,N_42832,N_42227);
nor U43655 (N_43655,N_42621,N_42270);
and U43656 (N_43656,N_42317,N_42680);
nor U43657 (N_43657,N_42522,N_42369);
or U43658 (N_43658,N_42128,N_42860);
xnor U43659 (N_43659,N_42672,N_42119);
nor U43660 (N_43660,N_42812,N_42635);
or U43661 (N_43661,N_42722,N_42059);
nor U43662 (N_43662,N_42149,N_42832);
nor U43663 (N_43663,N_42668,N_42855);
xnor U43664 (N_43664,N_42694,N_42484);
and U43665 (N_43665,N_42257,N_42979);
nor U43666 (N_43666,N_42446,N_42609);
and U43667 (N_43667,N_42300,N_42903);
or U43668 (N_43668,N_42429,N_42083);
xnor U43669 (N_43669,N_42312,N_42750);
or U43670 (N_43670,N_42021,N_42592);
and U43671 (N_43671,N_42176,N_42651);
nand U43672 (N_43672,N_42975,N_42441);
nand U43673 (N_43673,N_42515,N_42244);
xnor U43674 (N_43674,N_42365,N_42974);
nand U43675 (N_43675,N_42089,N_42975);
and U43676 (N_43676,N_42048,N_42467);
or U43677 (N_43677,N_42926,N_42913);
nor U43678 (N_43678,N_42352,N_42023);
or U43679 (N_43679,N_42127,N_42411);
and U43680 (N_43680,N_42088,N_42293);
xnor U43681 (N_43681,N_42718,N_42995);
or U43682 (N_43682,N_42054,N_42900);
nand U43683 (N_43683,N_42991,N_42574);
nand U43684 (N_43684,N_42846,N_42636);
or U43685 (N_43685,N_42611,N_42772);
or U43686 (N_43686,N_42110,N_42991);
or U43687 (N_43687,N_42872,N_42241);
nand U43688 (N_43688,N_42377,N_42568);
nor U43689 (N_43689,N_42526,N_42663);
nor U43690 (N_43690,N_42941,N_42426);
nand U43691 (N_43691,N_42091,N_42191);
or U43692 (N_43692,N_42998,N_42854);
and U43693 (N_43693,N_42898,N_42687);
xor U43694 (N_43694,N_42250,N_42033);
nor U43695 (N_43695,N_42920,N_42170);
nor U43696 (N_43696,N_42115,N_42052);
or U43697 (N_43697,N_42858,N_42922);
xnor U43698 (N_43698,N_42116,N_42579);
and U43699 (N_43699,N_42037,N_42405);
nand U43700 (N_43700,N_42424,N_42406);
xor U43701 (N_43701,N_42724,N_42645);
and U43702 (N_43702,N_42562,N_42319);
and U43703 (N_43703,N_42857,N_42740);
xnor U43704 (N_43704,N_42122,N_42649);
or U43705 (N_43705,N_42192,N_42151);
xnor U43706 (N_43706,N_42746,N_42034);
nand U43707 (N_43707,N_42740,N_42373);
xor U43708 (N_43708,N_42753,N_42672);
and U43709 (N_43709,N_42533,N_42622);
nor U43710 (N_43710,N_42593,N_42643);
nor U43711 (N_43711,N_42664,N_42427);
nor U43712 (N_43712,N_42725,N_42846);
nand U43713 (N_43713,N_42727,N_42890);
and U43714 (N_43714,N_42648,N_42530);
xnor U43715 (N_43715,N_42123,N_42542);
nand U43716 (N_43716,N_42704,N_42840);
or U43717 (N_43717,N_42697,N_42878);
nor U43718 (N_43718,N_42196,N_42391);
or U43719 (N_43719,N_42758,N_42994);
or U43720 (N_43720,N_42480,N_42545);
and U43721 (N_43721,N_42678,N_42039);
xnor U43722 (N_43722,N_42335,N_42520);
and U43723 (N_43723,N_42611,N_42302);
or U43724 (N_43724,N_42786,N_42222);
nand U43725 (N_43725,N_42104,N_42089);
nor U43726 (N_43726,N_42655,N_42003);
xnor U43727 (N_43727,N_42645,N_42080);
xnor U43728 (N_43728,N_42306,N_42593);
xor U43729 (N_43729,N_42474,N_42188);
or U43730 (N_43730,N_42590,N_42060);
and U43731 (N_43731,N_42429,N_42523);
and U43732 (N_43732,N_42289,N_42593);
nand U43733 (N_43733,N_42520,N_42534);
nand U43734 (N_43734,N_42964,N_42458);
nor U43735 (N_43735,N_42518,N_42640);
nand U43736 (N_43736,N_42418,N_42958);
nor U43737 (N_43737,N_42378,N_42229);
xnor U43738 (N_43738,N_42712,N_42977);
xor U43739 (N_43739,N_42409,N_42704);
nand U43740 (N_43740,N_42772,N_42409);
nor U43741 (N_43741,N_42581,N_42605);
and U43742 (N_43742,N_42293,N_42799);
nor U43743 (N_43743,N_42575,N_42306);
xnor U43744 (N_43744,N_42306,N_42051);
nor U43745 (N_43745,N_42724,N_42225);
or U43746 (N_43746,N_42247,N_42666);
or U43747 (N_43747,N_42090,N_42511);
nand U43748 (N_43748,N_42222,N_42317);
or U43749 (N_43749,N_42729,N_42877);
and U43750 (N_43750,N_42464,N_42532);
and U43751 (N_43751,N_42854,N_42424);
or U43752 (N_43752,N_42584,N_42450);
and U43753 (N_43753,N_42229,N_42464);
and U43754 (N_43754,N_42437,N_42842);
nand U43755 (N_43755,N_42928,N_42083);
or U43756 (N_43756,N_42858,N_42423);
xnor U43757 (N_43757,N_42219,N_42562);
nor U43758 (N_43758,N_42107,N_42025);
nor U43759 (N_43759,N_42689,N_42634);
xnor U43760 (N_43760,N_42435,N_42534);
xnor U43761 (N_43761,N_42032,N_42763);
nand U43762 (N_43762,N_42349,N_42386);
xor U43763 (N_43763,N_42986,N_42162);
nor U43764 (N_43764,N_42314,N_42467);
and U43765 (N_43765,N_42733,N_42389);
nor U43766 (N_43766,N_42709,N_42976);
xnor U43767 (N_43767,N_42626,N_42045);
and U43768 (N_43768,N_42674,N_42826);
nand U43769 (N_43769,N_42129,N_42534);
xnor U43770 (N_43770,N_42982,N_42981);
and U43771 (N_43771,N_42539,N_42607);
and U43772 (N_43772,N_42175,N_42740);
nor U43773 (N_43773,N_42278,N_42135);
or U43774 (N_43774,N_42108,N_42161);
or U43775 (N_43775,N_42131,N_42874);
and U43776 (N_43776,N_42885,N_42291);
nor U43777 (N_43777,N_42114,N_42322);
and U43778 (N_43778,N_42314,N_42034);
nand U43779 (N_43779,N_42213,N_42485);
nor U43780 (N_43780,N_42924,N_42964);
nand U43781 (N_43781,N_42219,N_42372);
and U43782 (N_43782,N_42206,N_42219);
xor U43783 (N_43783,N_42404,N_42542);
xor U43784 (N_43784,N_42684,N_42917);
xnor U43785 (N_43785,N_42582,N_42303);
nor U43786 (N_43786,N_42581,N_42914);
nand U43787 (N_43787,N_42137,N_42105);
xnor U43788 (N_43788,N_42310,N_42155);
or U43789 (N_43789,N_42440,N_42890);
nor U43790 (N_43790,N_42746,N_42998);
xor U43791 (N_43791,N_42334,N_42557);
nand U43792 (N_43792,N_42414,N_42343);
nor U43793 (N_43793,N_42506,N_42021);
nor U43794 (N_43794,N_42877,N_42589);
nor U43795 (N_43795,N_42962,N_42384);
and U43796 (N_43796,N_42629,N_42636);
nand U43797 (N_43797,N_42390,N_42978);
and U43798 (N_43798,N_42024,N_42752);
xnor U43799 (N_43799,N_42231,N_42949);
or U43800 (N_43800,N_42414,N_42701);
xnor U43801 (N_43801,N_42518,N_42732);
nand U43802 (N_43802,N_42233,N_42371);
or U43803 (N_43803,N_42656,N_42357);
and U43804 (N_43804,N_42335,N_42626);
xor U43805 (N_43805,N_42991,N_42441);
nor U43806 (N_43806,N_42288,N_42502);
or U43807 (N_43807,N_42536,N_42198);
nor U43808 (N_43808,N_42460,N_42654);
or U43809 (N_43809,N_42117,N_42542);
or U43810 (N_43810,N_42704,N_42108);
or U43811 (N_43811,N_42662,N_42875);
or U43812 (N_43812,N_42229,N_42723);
or U43813 (N_43813,N_42615,N_42583);
xor U43814 (N_43814,N_42024,N_42044);
nor U43815 (N_43815,N_42908,N_42053);
xor U43816 (N_43816,N_42753,N_42023);
nand U43817 (N_43817,N_42105,N_42668);
and U43818 (N_43818,N_42004,N_42564);
or U43819 (N_43819,N_42388,N_42503);
nand U43820 (N_43820,N_42349,N_42582);
xor U43821 (N_43821,N_42222,N_42419);
nand U43822 (N_43822,N_42122,N_42656);
nand U43823 (N_43823,N_42385,N_42196);
xnor U43824 (N_43824,N_42105,N_42097);
xor U43825 (N_43825,N_42061,N_42825);
nor U43826 (N_43826,N_42642,N_42255);
xnor U43827 (N_43827,N_42670,N_42799);
or U43828 (N_43828,N_42985,N_42820);
and U43829 (N_43829,N_42247,N_42953);
or U43830 (N_43830,N_42211,N_42831);
xor U43831 (N_43831,N_42125,N_42049);
and U43832 (N_43832,N_42773,N_42586);
or U43833 (N_43833,N_42844,N_42396);
and U43834 (N_43834,N_42334,N_42798);
xor U43835 (N_43835,N_42165,N_42634);
nand U43836 (N_43836,N_42904,N_42734);
xor U43837 (N_43837,N_42640,N_42117);
nor U43838 (N_43838,N_42055,N_42969);
or U43839 (N_43839,N_42382,N_42719);
xor U43840 (N_43840,N_42788,N_42587);
nor U43841 (N_43841,N_42459,N_42639);
or U43842 (N_43842,N_42808,N_42389);
xnor U43843 (N_43843,N_42881,N_42458);
or U43844 (N_43844,N_42552,N_42909);
nand U43845 (N_43845,N_42747,N_42318);
and U43846 (N_43846,N_42387,N_42688);
nand U43847 (N_43847,N_42211,N_42835);
or U43848 (N_43848,N_42798,N_42892);
xor U43849 (N_43849,N_42321,N_42055);
or U43850 (N_43850,N_42573,N_42220);
and U43851 (N_43851,N_42753,N_42054);
nand U43852 (N_43852,N_42883,N_42796);
nand U43853 (N_43853,N_42331,N_42743);
nand U43854 (N_43854,N_42217,N_42831);
or U43855 (N_43855,N_42757,N_42043);
and U43856 (N_43856,N_42189,N_42205);
nand U43857 (N_43857,N_42566,N_42264);
or U43858 (N_43858,N_42986,N_42683);
nand U43859 (N_43859,N_42146,N_42717);
xnor U43860 (N_43860,N_42323,N_42111);
and U43861 (N_43861,N_42823,N_42651);
or U43862 (N_43862,N_42628,N_42438);
or U43863 (N_43863,N_42635,N_42980);
nor U43864 (N_43864,N_42373,N_42856);
nor U43865 (N_43865,N_42325,N_42227);
nor U43866 (N_43866,N_42566,N_42784);
xor U43867 (N_43867,N_42224,N_42560);
or U43868 (N_43868,N_42612,N_42740);
or U43869 (N_43869,N_42336,N_42345);
nor U43870 (N_43870,N_42128,N_42953);
nand U43871 (N_43871,N_42568,N_42018);
nor U43872 (N_43872,N_42414,N_42818);
and U43873 (N_43873,N_42687,N_42702);
and U43874 (N_43874,N_42006,N_42536);
nor U43875 (N_43875,N_42344,N_42535);
xnor U43876 (N_43876,N_42699,N_42338);
or U43877 (N_43877,N_42879,N_42928);
and U43878 (N_43878,N_42844,N_42969);
or U43879 (N_43879,N_42643,N_42569);
xor U43880 (N_43880,N_42230,N_42787);
nand U43881 (N_43881,N_42833,N_42396);
nand U43882 (N_43882,N_42865,N_42666);
nor U43883 (N_43883,N_42064,N_42191);
or U43884 (N_43884,N_42108,N_42956);
nor U43885 (N_43885,N_42840,N_42218);
nand U43886 (N_43886,N_42579,N_42943);
nand U43887 (N_43887,N_42970,N_42488);
nor U43888 (N_43888,N_42144,N_42475);
or U43889 (N_43889,N_42760,N_42868);
nor U43890 (N_43890,N_42234,N_42190);
and U43891 (N_43891,N_42128,N_42359);
nand U43892 (N_43892,N_42034,N_42615);
or U43893 (N_43893,N_42763,N_42906);
nand U43894 (N_43894,N_42820,N_42345);
and U43895 (N_43895,N_42100,N_42706);
nor U43896 (N_43896,N_42265,N_42658);
xnor U43897 (N_43897,N_42545,N_42306);
or U43898 (N_43898,N_42066,N_42046);
nor U43899 (N_43899,N_42347,N_42664);
xor U43900 (N_43900,N_42600,N_42900);
nor U43901 (N_43901,N_42435,N_42123);
nand U43902 (N_43902,N_42906,N_42336);
nor U43903 (N_43903,N_42064,N_42483);
nor U43904 (N_43904,N_42522,N_42404);
and U43905 (N_43905,N_42917,N_42821);
nand U43906 (N_43906,N_42961,N_42187);
xnor U43907 (N_43907,N_42270,N_42028);
nand U43908 (N_43908,N_42485,N_42064);
xor U43909 (N_43909,N_42131,N_42986);
xor U43910 (N_43910,N_42873,N_42548);
and U43911 (N_43911,N_42196,N_42387);
or U43912 (N_43912,N_42177,N_42469);
or U43913 (N_43913,N_42745,N_42574);
nor U43914 (N_43914,N_42702,N_42278);
nor U43915 (N_43915,N_42696,N_42356);
and U43916 (N_43916,N_42070,N_42571);
nor U43917 (N_43917,N_42425,N_42312);
xnor U43918 (N_43918,N_42719,N_42730);
nand U43919 (N_43919,N_42154,N_42000);
xnor U43920 (N_43920,N_42983,N_42749);
xnor U43921 (N_43921,N_42858,N_42448);
nor U43922 (N_43922,N_42298,N_42953);
nor U43923 (N_43923,N_42392,N_42402);
and U43924 (N_43924,N_42122,N_42744);
nand U43925 (N_43925,N_42595,N_42516);
nor U43926 (N_43926,N_42774,N_42984);
nor U43927 (N_43927,N_42070,N_42405);
or U43928 (N_43928,N_42571,N_42801);
nor U43929 (N_43929,N_42098,N_42916);
or U43930 (N_43930,N_42965,N_42469);
or U43931 (N_43931,N_42340,N_42998);
nor U43932 (N_43932,N_42943,N_42500);
nor U43933 (N_43933,N_42088,N_42455);
xor U43934 (N_43934,N_42239,N_42695);
nor U43935 (N_43935,N_42789,N_42886);
nand U43936 (N_43936,N_42780,N_42046);
nand U43937 (N_43937,N_42348,N_42293);
and U43938 (N_43938,N_42752,N_42050);
xor U43939 (N_43939,N_42669,N_42463);
or U43940 (N_43940,N_42833,N_42456);
or U43941 (N_43941,N_42855,N_42124);
nand U43942 (N_43942,N_42126,N_42094);
nor U43943 (N_43943,N_42251,N_42920);
nor U43944 (N_43944,N_42451,N_42746);
xor U43945 (N_43945,N_42174,N_42702);
or U43946 (N_43946,N_42233,N_42061);
or U43947 (N_43947,N_42441,N_42906);
nand U43948 (N_43948,N_42994,N_42773);
nand U43949 (N_43949,N_42569,N_42449);
and U43950 (N_43950,N_42006,N_42937);
xor U43951 (N_43951,N_42504,N_42984);
or U43952 (N_43952,N_42005,N_42103);
nand U43953 (N_43953,N_42843,N_42839);
and U43954 (N_43954,N_42499,N_42511);
nor U43955 (N_43955,N_42446,N_42852);
and U43956 (N_43956,N_42797,N_42176);
xor U43957 (N_43957,N_42386,N_42306);
nor U43958 (N_43958,N_42332,N_42121);
or U43959 (N_43959,N_42661,N_42025);
nor U43960 (N_43960,N_42189,N_42650);
nor U43961 (N_43961,N_42492,N_42043);
nor U43962 (N_43962,N_42760,N_42078);
nor U43963 (N_43963,N_42364,N_42750);
and U43964 (N_43964,N_42776,N_42730);
nand U43965 (N_43965,N_42697,N_42816);
xnor U43966 (N_43966,N_42501,N_42468);
or U43967 (N_43967,N_42118,N_42263);
and U43968 (N_43968,N_42209,N_42085);
or U43969 (N_43969,N_42446,N_42589);
or U43970 (N_43970,N_42238,N_42492);
or U43971 (N_43971,N_42415,N_42985);
nor U43972 (N_43972,N_42088,N_42435);
nand U43973 (N_43973,N_42532,N_42172);
or U43974 (N_43974,N_42750,N_42145);
or U43975 (N_43975,N_42265,N_42968);
nor U43976 (N_43976,N_42748,N_42779);
and U43977 (N_43977,N_42175,N_42326);
xnor U43978 (N_43978,N_42063,N_42485);
and U43979 (N_43979,N_42301,N_42050);
xnor U43980 (N_43980,N_42382,N_42610);
nor U43981 (N_43981,N_42757,N_42151);
and U43982 (N_43982,N_42885,N_42656);
and U43983 (N_43983,N_42559,N_42185);
or U43984 (N_43984,N_42850,N_42969);
xor U43985 (N_43985,N_42428,N_42903);
nor U43986 (N_43986,N_42008,N_42746);
and U43987 (N_43987,N_42265,N_42332);
xor U43988 (N_43988,N_42644,N_42969);
or U43989 (N_43989,N_42191,N_42837);
nor U43990 (N_43990,N_42035,N_42438);
or U43991 (N_43991,N_42228,N_42718);
nor U43992 (N_43992,N_42476,N_42995);
xnor U43993 (N_43993,N_42262,N_42154);
or U43994 (N_43994,N_42897,N_42010);
xor U43995 (N_43995,N_42358,N_42682);
xor U43996 (N_43996,N_42089,N_42549);
xor U43997 (N_43997,N_42742,N_42650);
nand U43998 (N_43998,N_42796,N_42747);
xor U43999 (N_43999,N_42042,N_42035);
or U44000 (N_44000,N_43047,N_43228);
or U44001 (N_44001,N_43596,N_43694);
xnor U44002 (N_44002,N_43203,N_43490);
and U44003 (N_44003,N_43450,N_43400);
and U44004 (N_44004,N_43572,N_43365);
or U44005 (N_44005,N_43724,N_43292);
xor U44006 (N_44006,N_43139,N_43125);
or U44007 (N_44007,N_43967,N_43735);
xor U44008 (N_44008,N_43373,N_43609);
nand U44009 (N_44009,N_43117,N_43612);
nor U44010 (N_44010,N_43987,N_43314);
nand U44011 (N_44011,N_43994,N_43944);
nor U44012 (N_44012,N_43178,N_43091);
or U44013 (N_44013,N_43981,N_43827);
nor U44014 (N_44014,N_43273,N_43756);
xnor U44015 (N_44015,N_43169,N_43798);
nor U44016 (N_44016,N_43473,N_43386);
xor U44017 (N_44017,N_43749,N_43915);
nor U44018 (N_44018,N_43281,N_43330);
xor U44019 (N_44019,N_43313,N_43343);
nor U44020 (N_44020,N_43268,N_43076);
or U44021 (N_44021,N_43719,N_43112);
and U44022 (N_44022,N_43776,N_43498);
or U44023 (N_44023,N_43843,N_43005);
xor U44024 (N_44024,N_43451,N_43437);
nor U44025 (N_44025,N_43443,N_43555);
nor U44026 (N_44026,N_43906,N_43908);
and U44027 (N_44027,N_43895,N_43767);
and U44028 (N_44028,N_43624,N_43298);
nand U44029 (N_44029,N_43684,N_43757);
and U44030 (N_44030,N_43050,N_43833);
and U44031 (N_44031,N_43340,N_43030);
nor U44032 (N_44032,N_43722,N_43529);
and U44033 (N_44033,N_43739,N_43222);
nand U44034 (N_44034,N_43607,N_43920);
and U44035 (N_44035,N_43973,N_43114);
xor U44036 (N_44036,N_43699,N_43935);
or U44037 (N_44037,N_43802,N_43662);
nor U44038 (N_44038,N_43746,N_43872);
nor U44039 (N_44039,N_43301,N_43744);
xor U44040 (N_44040,N_43462,N_43209);
nand U44041 (N_44041,N_43962,N_43177);
xnor U44042 (N_44042,N_43457,N_43339);
nand U44043 (N_44043,N_43602,N_43140);
nor U44044 (N_44044,N_43585,N_43149);
nor U44045 (N_44045,N_43069,N_43928);
or U44046 (N_44046,N_43784,N_43970);
or U44047 (N_44047,N_43007,N_43870);
and U44048 (N_44048,N_43295,N_43493);
nand U44049 (N_44049,N_43098,N_43708);
or U44050 (N_44050,N_43816,N_43315);
or U44051 (N_44051,N_43855,N_43977);
nand U44052 (N_44052,N_43147,N_43282);
xnor U44053 (N_44053,N_43564,N_43865);
or U44054 (N_44054,N_43530,N_43310);
and U44055 (N_44055,N_43914,N_43847);
nand U44056 (N_44056,N_43955,N_43853);
xor U44057 (N_44057,N_43041,N_43760);
and U44058 (N_44058,N_43425,N_43848);
or U44059 (N_44059,N_43943,N_43531);
nor U44060 (N_44060,N_43033,N_43308);
nand U44061 (N_44061,N_43629,N_43038);
nor U44062 (N_44062,N_43547,N_43590);
nand U44063 (N_44063,N_43185,N_43689);
or U44064 (N_44064,N_43604,N_43353);
or U44065 (N_44065,N_43211,N_43900);
xnor U44066 (N_44066,N_43247,N_43413);
nand U44067 (N_44067,N_43713,N_43415);
xnor U44068 (N_44068,N_43186,N_43674);
xor U44069 (N_44069,N_43960,N_43912);
and U44070 (N_44070,N_43219,N_43600);
xnor U44071 (N_44071,N_43785,N_43893);
or U44072 (N_44072,N_43902,N_43601);
xor U44073 (N_44073,N_43773,N_43469);
nor U44074 (N_44074,N_43546,N_43525);
or U44075 (N_44075,N_43747,N_43840);
nor U44076 (N_44076,N_43874,N_43532);
and U44077 (N_44077,N_43367,N_43333);
xor U44078 (N_44078,N_43284,N_43477);
and U44079 (N_44079,N_43288,N_43143);
nand U44080 (N_44080,N_43605,N_43402);
and U44081 (N_44081,N_43653,N_43334);
xnor U44082 (N_44082,N_43535,N_43946);
nor U44083 (N_44083,N_43412,N_43082);
xnor U44084 (N_44084,N_43976,N_43107);
nand U44085 (N_44085,N_43740,N_43225);
or U44086 (N_44086,N_43834,N_43048);
nand U44087 (N_44087,N_43787,N_43841);
xnor U44088 (N_44088,N_43763,N_43283);
or U44089 (N_44089,N_43108,N_43709);
and U44090 (N_44090,N_43949,N_43495);
and U44091 (N_44091,N_43680,N_43028);
xor U44092 (N_44092,N_43509,N_43697);
xor U44093 (N_44093,N_43817,N_43964);
nor U44094 (N_44094,N_43475,N_43064);
and U44095 (N_44095,N_43020,N_43641);
xor U44096 (N_44096,N_43772,N_43622);
nor U44097 (N_44097,N_43542,N_43877);
nand U44098 (N_44098,N_43644,N_43356);
xor U44099 (N_44099,N_43594,N_43441);
nor U44100 (N_44100,N_43974,N_43246);
xor U44101 (N_44101,N_43300,N_43510);
and U44102 (N_44102,N_43567,N_43545);
nand U44103 (N_44103,N_43901,N_43579);
nor U44104 (N_44104,N_43319,N_43860);
or U44105 (N_44105,N_43677,N_43102);
or U44106 (N_44106,N_43471,N_43382);
and U44107 (N_44107,N_43696,N_43921);
and U44108 (N_44108,N_43364,N_43253);
and U44109 (N_44109,N_43716,N_43474);
xor U44110 (N_44110,N_43170,N_43686);
or U44111 (N_44111,N_43878,N_43968);
or U44112 (N_44112,N_43200,N_43110);
xnor U44113 (N_44113,N_43565,N_43312);
and U44114 (N_44114,N_43801,N_43769);
xnor U44115 (N_44115,N_43807,N_43371);
nand U44116 (N_44116,N_43737,N_43500);
or U44117 (N_44117,N_43990,N_43428);
xnor U44118 (N_44118,N_43839,N_43741);
or U44119 (N_44119,N_43327,N_43232);
nor U44120 (N_44120,N_43942,N_43698);
nor U44121 (N_44121,N_43911,N_43099);
nand U44122 (N_44122,N_43499,N_43933);
nor U44123 (N_44123,N_43182,N_43126);
nand U44124 (N_44124,N_43925,N_43771);
and U44125 (N_44125,N_43562,N_43775);
and U44126 (N_44126,N_43966,N_43006);
or U44127 (N_44127,N_43369,N_43777);
nand U44128 (N_44128,N_43589,N_43844);
and U44129 (N_44129,N_43276,N_43389);
nor U44130 (N_44130,N_43941,N_43057);
xnor U44131 (N_44131,N_43591,N_43891);
xor U44132 (N_44132,N_43507,N_43431);
xor U44133 (N_44133,N_43536,N_43266);
and U44134 (N_44134,N_43146,N_43279);
and U44135 (N_44135,N_43213,N_43285);
xor U44136 (N_44136,N_43461,N_43808);
nor U44137 (N_44137,N_43448,N_43537);
or U44138 (N_44138,N_43486,N_43963);
nand U44139 (N_44139,N_43951,N_43027);
or U44140 (N_44140,N_43275,N_43189);
nor U44141 (N_44141,N_43634,N_43732);
nand U44142 (N_44142,N_43692,N_43916);
or U44143 (N_44143,N_43818,N_43615);
nor U44144 (N_44144,N_43411,N_43418);
xor U44145 (N_44145,N_43274,N_43676);
or U44146 (N_44146,N_43265,N_43804);
xnor U44147 (N_44147,N_43354,N_43563);
and U44148 (N_44148,N_43937,N_43826);
or U44149 (N_44149,N_43693,N_43049);
or U44150 (N_44150,N_43145,N_43237);
or U44151 (N_44151,N_43574,N_43329);
or U44152 (N_44152,N_43183,N_43986);
or U44153 (N_44153,N_43433,N_43635);
and U44154 (N_44154,N_43121,N_43861);
nand U44155 (N_44155,N_43637,N_43578);
and U44156 (N_44156,N_43081,N_43142);
nor U44157 (N_44157,N_43190,N_43862);
or U44158 (N_44158,N_43561,N_43181);
or U44159 (N_44159,N_43559,N_43240);
nand U44160 (N_44160,N_43399,N_43950);
and U44161 (N_44161,N_43290,N_43945);
nor U44162 (N_44162,N_43257,N_43666);
nor U44163 (N_44163,N_43780,N_43639);
or U44164 (N_44164,N_43056,N_43938);
or U44165 (N_44165,N_43717,N_43224);
nand U44166 (N_44166,N_43053,N_43096);
nand U44167 (N_44167,N_43813,N_43882);
or U44168 (N_44168,N_43445,N_43791);
nor U44169 (N_44169,N_43851,N_43318);
xor U44170 (N_44170,N_43161,N_43258);
nor U44171 (N_44171,N_43518,N_43023);
and U44172 (N_44172,N_43360,N_43778);
xnor U44173 (N_44173,N_43001,N_43800);
nand U44174 (N_44174,N_43338,N_43971);
nand U44175 (N_44175,N_43095,N_43370);
nor U44176 (N_44176,N_43859,N_43100);
nand U44177 (N_44177,N_43188,N_43707);
xor U44178 (N_44178,N_43191,N_43830);
or U44179 (N_44179,N_43077,N_43505);
nor U44180 (N_44180,N_43018,N_43180);
and U44181 (N_44181,N_43278,N_43723);
xor U44182 (N_44182,N_43299,N_43452);
nor U44183 (N_44183,N_43144,N_43435);
or U44184 (N_44184,N_43393,N_43460);
and U44185 (N_44185,N_43195,N_43598);
xor U44186 (N_44186,N_43204,N_43754);
nor U44187 (N_44187,N_43133,N_43062);
or U44188 (N_44188,N_43588,N_43384);
nor U44189 (N_44189,N_43194,N_43811);
or U44190 (N_44190,N_43829,N_43538);
nand U44191 (N_44191,N_43710,N_43026);
nor U44192 (N_44192,N_43328,N_43658);
xor U44193 (N_44193,N_43132,N_43700);
nand U44194 (N_44194,N_43845,N_43199);
nor U44195 (N_44195,N_43372,N_43036);
nand U44196 (N_44196,N_43106,N_43506);
or U44197 (N_44197,N_43280,N_43712);
nor U44198 (N_44198,N_43051,N_43002);
or U44199 (N_44199,N_43119,N_43704);
and U44200 (N_44200,N_43972,N_43094);
and U44201 (N_44201,N_43464,N_43439);
or U44202 (N_44202,N_43230,N_43640);
and U44203 (N_44203,N_43683,N_43163);
or U44204 (N_44204,N_43482,N_43122);
or U44205 (N_44205,N_43101,N_43856);
and U44206 (N_44206,N_43823,N_43032);
xnor U44207 (N_44207,N_43066,N_43380);
and U44208 (N_44208,N_43993,N_43297);
xor U44209 (N_44209,N_43476,N_43000);
nand U44210 (N_44210,N_43919,N_43991);
nor U44211 (N_44211,N_43999,N_43489);
or U44212 (N_44212,N_43446,N_43502);
or U44213 (N_44213,N_43430,N_43034);
nand U44214 (N_44214,N_43260,N_43271);
or U44215 (N_44215,N_43690,N_43376);
xor U44216 (N_44216,N_43383,N_43786);
and U44217 (N_44217,N_43294,N_43515);
or U44218 (N_44218,N_43206,N_43646);
or U44219 (N_44219,N_43391,N_43670);
nor U44220 (N_44220,N_43892,N_43158);
or U44221 (N_44221,N_43401,N_43654);
nor U44222 (N_44222,N_43350,N_43819);
nand U44223 (N_44223,N_43332,N_43262);
or U44224 (N_44224,N_43521,N_43961);
xor U44225 (N_44225,N_43837,N_43661);
nor U44226 (N_44226,N_43029,N_43608);
or U44227 (N_44227,N_43583,N_43358);
xor U44228 (N_44228,N_43603,N_43336);
nor U44229 (N_44229,N_43820,N_43141);
or U44230 (N_44230,N_43085,N_43116);
or U44231 (N_44231,N_43959,N_43742);
or U44232 (N_44232,N_43011,N_43909);
xor U44233 (N_44233,N_43725,N_43035);
nor U44234 (N_44234,N_43166,N_43571);
or U44235 (N_44235,N_43207,N_43753);
or U44236 (N_44236,N_43058,N_43998);
or U44237 (N_44237,N_43037,N_43361);
and U44238 (N_44238,N_43947,N_43174);
or U44239 (N_44239,N_43846,N_43688);
nand U44240 (N_44240,N_43377,N_43884);
nor U44241 (N_44241,N_43514,N_43215);
and U44242 (N_44242,N_43347,N_43470);
or U44243 (N_44243,N_43508,N_43927);
and U44244 (N_44244,N_43014,N_43304);
nand U44245 (N_44245,N_43645,N_43783);
xnor U44246 (N_44246,N_43325,N_43135);
xnor U44247 (N_44247,N_43003,N_43952);
nand U44248 (N_44248,N_43889,N_43750);
and U44249 (N_44249,N_43824,N_43012);
or U44250 (N_44250,N_43067,N_43396);
or U44251 (N_44251,N_43187,N_43782);
nor U44252 (N_44252,N_43019,N_43581);
and U44253 (N_44253,N_43103,N_43828);
nand U44254 (N_44254,N_43766,N_43429);
nor U44255 (N_44255,N_43903,N_43236);
nand U44256 (N_44256,N_43503,N_43617);
and U44257 (N_44257,N_43394,N_43072);
nor U44258 (N_44258,N_43426,N_43483);
xor U44259 (N_44259,N_43478,N_43256);
or U44260 (N_44260,N_43447,N_43229);
nor U44261 (N_44261,N_43918,N_43625);
xor U44262 (N_44262,N_43434,N_43907);
or U44263 (N_44263,N_43613,N_43910);
and U44264 (N_44264,N_43423,N_43835);
and U44265 (N_44265,N_43168,N_43930);
nand U44266 (N_44266,N_43650,N_43541);
or U44267 (N_44267,N_43992,N_43796);
and U44268 (N_44268,N_43831,N_43042);
and U44269 (N_44269,N_43931,N_43701);
and U44270 (N_44270,N_43836,N_43205);
xnor U44271 (N_44271,N_43729,N_43794);
or U44272 (N_44272,N_43522,N_43795);
nand U44273 (N_44273,N_43592,N_43071);
xnor U44274 (N_44274,N_43210,N_43044);
nand U44275 (N_44275,N_43586,N_43235);
and U44276 (N_44276,N_43458,N_43454);
and U44277 (N_44277,N_43934,N_43533);
xnor U44278 (N_44278,N_43351,N_43449);
nor U44279 (N_44279,N_43517,N_43455);
or U44280 (N_44280,N_43414,N_43636);
nor U44281 (N_44281,N_43984,N_43788);
or U44282 (N_44282,N_43736,N_43160);
xor U44283 (N_44283,N_43223,N_43733);
nand U44284 (N_44284,N_43929,N_43936);
nor U44285 (N_44285,N_43953,N_43638);
or U44286 (N_44286,N_43277,N_43619);
nand U44287 (N_44287,N_43528,N_43492);
nand U44288 (N_44288,N_43326,N_43004);
xnor U44289 (N_44289,N_43876,N_43869);
nor U44290 (N_44290,N_43375,N_43021);
or U44291 (N_44291,N_43346,N_43385);
and U44292 (N_44292,N_43025,N_43109);
and U44293 (N_44293,N_43024,N_43263);
nor U44294 (N_44294,N_43648,N_43453);
nor U44295 (N_44295,N_43381,N_43444);
and U44296 (N_44296,N_43179,N_43923);
or U44297 (N_44297,N_43989,N_43173);
xor U44298 (N_44298,N_43924,N_43789);
nor U44299 (N_44299,N_43996,N_43587);
and U44300 (N_44300,N_43797,N_43781);
and U44301 (N_44301,N_43196,N_43259);
and U44302 (N_44302,N_43995,N_43269);
nand U44303 (N_44303,N_43255,N_43087);
nand U44304 (N_44304,N_43342,N_43496);
xnor U44305 (N_44305,N_43118,N_43467);
and U44306 (N_44306,N_43193,N_43123);
nor U44307 (N_44307,N_43084,N_43374);
nand U44308 (N_44308,N_43864,N_43761);
and U44309 (N_44309,N_43046,N_43850);
or U44310 (N_44310,N_43504,N_43616);
or U44311 (N_44311,N_43097,N_43129);
xnor U44312 (N_44312,N_43480,N_43655);
and U44313 (N_44313,N_43417,N_43664);
and U44314 (N_44314,N_43582,N_43218);
and U44315 (N_44315,N_43679,N_43809);
nand U44316 (N_44316,N_43408,N_43731);
or U44317 (N_44317,N_43242,N_43956);
nand U44318 (N_44318,N_43045,N_43352);
nor U44319 (N_44319,N_43089,N_43932);
nor U44320 (N_44320,N_43212,N_43172);
and U44321 (N_44321,N_43405,N_43523);
nor U44322 (N_44322,N_43849,N_43880);
nor U44323 (N_44323,N_43164,N_43896);
or U44324 (N_44324,N_43948,N_43569);
and U44325 (N_44325,N_43234,N_43863);
nand U44326 (N_44326,N_43551,N_43321);
and U44327 (N_44327,N_43153,N_43184);
and U44328 (N_44328,N_43887,N_43822);
nor U44329 (N_44329,N_43345,N_43286);
xnor U44330 (N_44330,N_43202,N_43244);
and U44331 (N_44331,N_43392,N_43980);
xor U44332 (N_44332,N_43303,N_43543);
and U44333 (N_44333,N_43770,N_43558);
nor U44334 (N_44334,N_43063,N_43815);
and U44335 (N_44335,N_43387,N_43759);
or U44336 (N_44336,N_43871,N_43104);
nand U44337 (N_44337,N_43468,N_43080);
nand U44338 (N_44338,N_43054,N_43768);
xnor U44339 (N_44339,N_43867,N_43293);
nor U44340 (N_44340,N_43440,N_43366);
or U44341 (N_44341,N_43151,N_43810);
or U44342 (N_44342,N_43337,N_43208);
nand U44343 (N_44343,N_43969,N_43611);
nand U44344 (N_44344,N_43243,N_43359);
xnor U44345 (N_44345,N_43652,N_43703);
or U44346 (N_44346,N_43883,N_43171);
nor U44347 (N_44347,N_43068,N_43721);
nand U44348 (N_44348,N_43702,N_43497);
nand U44349 (N_44349,N_43628,N_43407);
nor U44350 (N_44350,N_43630,N_43554);
nor U44351 (N_44351,N_43390,N_43623);
nand U44352 (N_44352,N_43881,N_43610);
xnor U44353 (N_44353,N_43040,N_43362);
or U44354 (N_44354,N_43074,N_43227);
or U44355 (N_44355,N_43159,N_43552);
xnor U44356 (N_44356,N_43251,N_43306);
nand U44357 (N_44357,N_43627,N_43894);
nand U44358 (N_44358,N_43241,N_43073);
nand U44359 (N_44359,N_43136,N_43484);
xnor U44360 (N_44360,N_43316,N_43534);
nor U44361 (N_44361,N_43805,N_43879);
or U44362 (N_44362,N_43706,N_43904);
and U44363 (N_44363,N_43649,N_43857);
or U44364 (N_44364,N_43519,N_43511);
nor U44365 (N_44365,N_43745,N_43442);
nand U44366 (N_44366,N_43570,N_43250);
and U44367 (N_44367,N_43656,N_43093);
nand U44368 (N_44368,N_43568,N_43672);
nor U44369 (N_44369,N_43762,N_43513);
nand U44370 (N_44370,N_43978,N_43388);
xnor U44371 (N_44371,N_43913,N_43165);
xnor U44372 (N_44372,N_43854,N_43403);
xor U44373 (N_44373,N_43105,N_43618);
nor U44374 (N_44374,N_43705,N_43010);
or U44375 (N_44375,N_43792,N_43065);
or U44376 (N_44376,N_43803,N_43682);
or U44377 (N_44377,N_43905,N_43621);
xnor U44378 (N_44378,N_43245,N_43852);
and U44379 (N_44379,N_43738,N_43566);
xnor U44380 (N_44380,N_43459,N_43039);
nand U44381 (N_44381,N_43549,N_43357);
nor U44382 (N_44382,N_43524,N_43432);
nor U44383 (N_44383,N_43424,N_43687);
nor U44384 (N_44384,N_43553,N_43083);
and U44385 (N_44385,N_43642,N_43217);
or U44386 (N_44386,N_43728,N_43660);
xnor U44387 (N_44387,N_43544,N_43331);
nor U44388 (N_44388,N_43291,N_43890);
and U44389 (N_44389,N_43626,N_43127);
xor U44390 (N_44390,N_43886,N_43550);
or U44391 (N_44391,N_43917,N_43985);
nor U44392 (N_44392,N_43481,N_43317);
and U44393 (N_44393,N_43556,N_43527);
xnor U44394 (N_44394,N_43821,N_43975);
nand U44395 (N_44395,N_43368,N_43577);
nor U44396 (N_44396,N_43214,N_43404);
and U44397 (N_44397,N_43718,N_43226);
and U44398 (N_44398,N_43957,N_43311);
nand U44399 (N_44399,N_43557,N_43156);
and U44400 (N_44400,N_43111,N_43239);
nand U44401 (N_44401,N_43363,N_43115);
nor U44402 (N_44402,N_43070,N_43814);
xnor U44403 (N_44403,N_43620,N_43120);
and U44404 (N_44404,N_43086,N_43485);
nor U44405 (N_44405,N_43599,N_43309);
nand U44406 (N_44406,N_43669,N_43885);
and U44407 (N_44407,N_43866,N_43261);
or U44408 (N_44408,N_43665,N_43052);
xor U44409 (N_44409,N_43264,N_43939);
and U44410 (N_44410,N_43320,N_43092);
nand U44411 (N_44411,N_43516,N_43595);
nand U44412 (N_44412,N_43580,N_43897);
and U44413 (N_44413,N_43015,N_43651);
or U44414 (N_44414,N_43305,N_43526);
nand U44415 (N_44415,N_43838,N_43075);
and U44416 (N_44416,N_43548,N_43422);
or U44417 (N_44417,N_43678,N_43248);
xor U44418 (N_44418,N_43162,N_43233);
nand U44419 (N_44419,N_43520,N_43465);
and U44420 (N_44420,N_43267,N_43270);
xor U44421 (N_44421,N_43958,N_43659);
and U44422 (N_44422,N_43512,N_43576);
or U44423 (N_44423,N_43965,N_43926);
nand U44424 (N_44424,N_43997,N_43249);
xnor U44425 (N_44425,N_43061,N_43888);
nand U44426 (N_44426,N_43079,N_43150);
xor U44427 (N_44427,N_43479,N_43197);
nor U44428 (N_44428,N_43220,N_43715);
or U44429 (N_44429,N_43631,N_43755);
xnor U44430 (N_44430,N_43922,N_43420);
nand U44431 (N_44431,N_43335,N_43008);
and U44432 (N_44432,N_43176,N_43988);
or U44433 (N_44433,N_43031,N_43501);
nand U44434 (N_44434,N_43216,N_43720);
and U44435 (N_44435,N_43379,N_43055);
or U44436 (N_44436,N_43348,N_43416);
and U44437 (N_44437,N_43875,N_43560);
and U44438 (N_44438,N_43765,N_43192);
nand U44439 (N_44439,N_43287,N_43137);
and U44440 (N_44440,N_43491,N_43983);
xor U44441 (N_44441,N_43472,N_43349);
or U44442 (N_44442,N_43302,N_43675);
nand U44443 (N_44443,N_43289,N_43427);
and U44444 (N_44444,N_43131,N_43378);
or U44445 (N_44445,N_43633,N_43774);
nor U44446 (N_44446,N_43438,N_43663);
nor U44447 (N_44447,N_43090,N_43494);
or U44448 (N_44448,N_43979,N_43231);
nand U44449 (N_44449,N_43940,N_43734);
and U44450 (N_44450,N_43790,N_43421);
or U44451 (N_44451,N_43647,N_43130);
or U44452 (N_44452,N_43398,N_43982);
or U44453 (N_44453,N_43017,N_43410);
or U44454 (N_44454,N_43307,N_43009);
nand U44455 (N_44455,N_43409,N_43606);
and U44456 (N_44456,N_43436,N_43873);
xor U44457 (N_44457,N_43272,N_43113);
nor U44458 (N_44458,N_43842,N_43463);
xor U44459 (N_44459,N_43730,N_43711);
nand U44460 (N_44460,N_43673,N_43751);
xor U44461 (N_44461,N_43825,N_43681);
and U44462 (N_44462,N_43016,N_43575);
or U44463 (N_44463,N_43355,N_43487);
nor U44464 (N_44464,N_43152,N_43078);
or U44465 (N_44465,N_43858,N_43323);
nand U44466 (N_44466,N_43344,N_43154);
xor U44467 (N_44467,N_43138,N_43198);
and U44468 (N_44468,N_43726,N_43668);
and U44469 (N_44469,N_43748,N_43322);
and U44470 (N_44470,N_43614,N_43124);
nand U44471 (N_44471,N_43657,N_43691);
nand U44472 (N_44472,N_43406,N_43812);
and U44473 (N_44473,N_43593,N_43201);
or U44474 (N_44474,N_43799,N_43743);
nor U44475 (N_44475,N_43296,N_43167);
nand U44476 (N_44476,N_43584,N_43540);
or U44477 (N_44477,N_43088,N_43148);
nor U44478 (N_44478,N_43128,N_43155);
or U44479 (N_44479,N_43254,N_43727);
and U44480 (N_44480,N_43341,N_43868);
xor U44481 (N_44481,N_43252,N_43806);
nand U44482 (N_44482,N_43779,N_43752);
and U44483 (N_44483,N_43013,N_43632);
and U44484 (N_44484,N_43395,N_43175);
xor U44485 (N_44485,N_43324,N_43832);
nor U44486 (N_44486,N_43134,N_43764);
nor U44487 (N_44487,N_43714,N_43954);
nand U44488 (N_44488,N_43456,N_43667);
nand U44489 (N_44489,N_43060,N_43793);
or U44490 (N_44490,N_43539,N_43397);
and U44491 (N_44491,N_43043,N_43597);
xor U44492 (N_44492,N_43466,N_43238);
xor U44493 (N_44493,N_43898,N_43059);
xnor U44494 (N_44494,N_43221,N_43643);
or U44495 (N_44495,N_43695,N_43022);
nor U44496 (N_44496,N_43157,N_43758);
nor U44497 (N_44497,N_43419,N_43488);
nand U44498 (N_44498,N_43685,N_43671);
nand U44499 (N_44499,N_43573,N_43899);
nor U44500 (N_44500,N_43204,N_43055);
and U44501 (N_44501,N_43750,N_43340);
nand U44502 (N_44502,N_43266,N_43211);
nor U44503 (N_44503,N_43604,N_43289);
nor U44504 (N_44504,N_43732,N_43525);
nand U44505 (N_44505,N_43774,N_43986);
nand U44506 (N_44506,N_43991,N_43471);
nand U44507 (N_44507,N_43687,N_43757);
nor U44508 (N_44508,N_43312,N_43421);
nor U44509 (N_44509,N_43313,N_43485);
and U44510 (N_44510,N_43537,N_43405);
nor U44511 (N_44511,N_43160,N_43589);
xor U44512 (N_44512,N_43822,N_43753);
xor U44513 (N_44513,N_43963,N_43336);
or U44514 (N_44514,N_43714,N_43669);
nor U44515 (N_44515,N_43770,N_43537);
nor U44516 (N_44516,N_43276,N_43030);
or U44517 (N_44517,N_43673,N_43194);
or U44518 (N_44518,N_43577,N_43633);
xnor U44519 (N_44519,N_43367,N_43085);
nor U44520 (N_44520,N_43119,N_43062);
nand U44521 (N_44521,N_43057,N_43531);
nand U44522 (N_44522,N_43622,N_43519);
xnor U44523 (N_44523,N_43581,N_43592);
or U44524 (N_44524,N_43319,N_43800);
nor U44525 (N_44525,N_43299,N_43226);
or U44526 (N_44526,N_43434,N_43379);
nor U44527 (N_44527,N_43420,N_43605);
nor U44528 (N_44528,N_43740,N_43191);
and U44529 (N_44529,N_43617,N_43943);
xnor U44530 (N_44530,N_43523,N_43031);
xor U44531 (N_44531,N_43927,N_43870);
or U44532 (N_44532,N_43229,N_43953);
nor U44533 (N_44533,N_43647,N_43345);
nor U44534 (N_44534,N_43650,N_43977);
and U44535 (N_44535,N_43667,N_43721);
and U44536 (N_44536,N_43053,N_43362);
and U44537 (N_44537,N_43612,N_43235);
xnor U44538 (N_44538,N_43696,N_43946);
xnor U44539 (N_44539,N_43635,N_43123);
xnor U44540 (N_44540,N_43162,N_43853);
nor U44541 (N_44541,N_43162,N_43604);
xnor U44542 (N_44542,N_43999,N_43044);
xnor U44543 (N_44543,N_43806,N_43053);
nor U44544 (N_44544,N_43819,N_43338);
and U44545 (N_44545,N_43007,N_43471);
or U44546 (N_44546,N_43541,N_43226);
or U44547 (N_44547,N_43420,N_43920);
and U44548 (N_44548,N_43298,N_43626);
xnor U44549 (N_44549,N_43772,N_43251);
and U44550 (N_44550,N_43024,N_43571);
nor U44551 (N_44551,N_43876,N_43966);
nor U44552 (N_44552,N_43471,N_43054);
xor U44553 (N_44553,N_43381,N_43732);
nor U44554 (N_44554,N_43932,N_43434);
xnor U44555 (N_44555,N_43681,N_43229);
or U44556 (N_44556,N_43432,N_43740);
nand U44557 (N_44557,N_43668,N_43977);
nand U44558 (N_44558,N_43130,N_43291);
xnor U44559 (N_44559,N_43550,N_43015);
xnor U44560 (N_44560,N_43540,N_43141);
nor U44561 (N_44561,N_43333,N_43656);
and U44562 (N_44562,N_43023,N_43323);
xnor U44563 (N_44563,N_43268,N_43566);
and U44564 (N_44564,N_43227,N_43786);
nand U44565 (N_44565,N_43379,N_43121);
nand U44566 (N_44566,N_43887,N_43906);
or U44567 (N_44567,N_43688,N_43120);
xor U44568 (N_44568,N_43536,N_43343);
nand U44569 (N_44569,N_43463,N_43107);
nand U44570 (N_44570,N_43076,N_43808);
nor U44571 (N_44571,N_43923,N_43142);
and U44572 (N_44572,N_43126,N_43244);
or U44573 (N_44573,N_43512,N_43491);
and U44574 (N_44574,N_43463,N_43960);
and U44575 (N_44575,N_43455,N_43539);
xor U44576 (N_44576,N_43952,N_43199);
xor U44577 (N_44577,N_43612,N_43043);
or U44578 (N_44578,N_43130,N_43808);
and U44579 (N_44579,N_43989,N_43788);
nor U44580 (N_44580,N_43391,N_43416);
nand U44581 (N_44581,N_43885,N_43098);
xor U44582 (N_44582,N_43008,N_43156);
xnor U44583 (N_44583,N_43063,N_43378);
or U44584 (N_44584,N_43666,N_43131);
or U44585 (N_44585,N_43712,N_43671);
and U44586 (N_44586,N_43773,N_43075);
or U44587 (N_44587,N_43714,N_43288);
nor U44588 (N_44588,N_43128,N_43644);
or U44589 (N_44589,N_43850,N_43796);
xnor U44590 (N_44590,N_43901,N_43101);
nand U44591 (N_44591,N_43334,N_43565);
nand U44592 (N_44592,N_43428,N_43568);
nand U44593 (N_44593,N_43502,N_43972);
and U44594 (N_44594,N_43067,N_43937);
xor U44595 (N_44595,N_43144,N_43107);
nor U44596 (N_44596,N_43102,N_43254);
xor U44597 (N_44597,N_43802,N_43171);
nor U44598 (N_44598,N_43305,N_43923);
nor U44599 (N_44599,N_43880,N_43274);
or U44600 (N_44600,N_43579,N_43955);
nand U44601 (N_44601,N_43359,N_43611);
or U44602 (N_44602,N_43380,N_43400);
and U44603 (N_44603,N_43890,N_43217);
or U44604 (N_44604,N_43899,N_43601);
and U44605 (N_44605,N_43537,N_43474);
xnor U44606 (N_44606,N_43905,N_43355);
and U44607 (N_44607,N_43121,N_43882);
and U44608 (N_44608,N_43446,N_43851);
and U44609 (N_44609,N_43244,N_43430);
or U44610 (N_44610,N_43112,N_43981);
xor U44611 (N_44611,N_43885,N_43533);
nand U44612 (N_44612,N_43488,N_43873);
and U44613 (N_44613,N_43900,N_43053);
xor U44614 (N_44614,N_43857,N_43459);
or U44615 (N_44615,N_43915,N_43954);
xnor U44616 (N_44616,N_43800,N_43851);
nand U44617 (N_44617,N_43593,N_43646);
and U44618 (N_44618,N_43377,N_43319);
xnor U44619 (N_44619,N_43767,N_43070);
nor U44620 (N_44620,N_43143,N_43392);
nand U44621 (N_44621,N_43222,N_43322);
nand U44622 (N_44622,N_43404,N_43066);
xnor U44623 (N_44623,N_43586,N_43871);
or U44624 (N_44624,N_43707,N_43977);
or U44625 (N_44625,N_43601,N_43130);
xor U44626 (N_44626,N_43448,N_43109);
and U44627 (N_44627,N_43733,N_43714);
xor U44628 (N_44628,N_43408,N_43285);
xor U44629 (N_44629,N_43363,N_43234);
and U44630 (N_44630,N_43314,N_43592);
nor U44631 (N_44631,N_43038,N_43741);
nor U44632 (N_44632,N_43584,N_43649);
nor U44633 (N_44633,N_43504,N_43263);
nand U44634 (N_44634,N_43138,N_43169);
nor U44635 (N_44635,N_43774,N_43918);
nor U44636 (N_44636,N_43437,N_43745);
nand U44637 (N_44637,N_43034,N_43180);
nor U44638 (N_44638,N_43661,N_43569);
and U44639 (N_44639,N_43554,N_43228);
nor U44640 (N_44640,N_43101,N_43558);
xor U44641 (N_44641,N_43050,N_43646);
nand U44642 (N_44642,N_43644,N_43332);
or U44643 (N_44643,N_43230,N_43292);
nor U44644 (N_44644,N_43842,N_43627);
xor U44645 (N_44645,N_43090,N_43324);
or U44646 (N_44646,N_43236,N_43168);
or U44647 (N_44647,N_43627,N_43512);
nand U44648 (N_44648,N_43448,N_43283);
and U44649 (N_44649,N_43281,N_43823);
and U44650 (N_44650,N_43014,N_43567);
nor U44651 (N_44651,N_43239,N_43560);
or U44652 (N_44652,N_43870,N_43803);
nor U44653 (N_44653,N_43022,N_43219);
nor U44654 (N_44654,N_43798,N_43709);
or U44655 (N_44655,N_43919,N_43825);
xor U44656 (N_44656,N_43688,N_43443);
or U44657 (N_44657,N_43881,N_43870);
nor U44658 (N_44658,N_43521,N_43702);
or U44659 (N_44659,N_43453,N_43697);
xnor U44660 (N_44660,N_43355,N_43753);
or U44661 (N_44661,N_43602,N_43290);
or U44662 (N_44662,N_43521,N_43298);
or U44663 (N_44663,N_43415,N_43243);
and U44664 (N_44664,N_43057,N_43807);
nor U44665 (N_44665,N_43554,N_43768);
or U44666 (N_44666,N_43917,N_43117);
xor U44667 (N_44667,N_43673,N_43149);
xor U44668 (N_44668,N_43783,N_43449);
nor U44669 (N_44669,N_43561,N_43761);
xnor U44670 (N_44670,N_43509,N_43880);
or U44671 (N_44671,N_43823,N_43756);
nand U44672 (N_44672,N_43758,N_43757);
nand U44673 (N_44673,N_43445,N_43618);
and U44674 (N_44674,N_43879,N_43388);
or U44675 (N_44675,N_43955,N_43328);
or U44676 (N_44676,N_43742,N_43652);
xnor U44677 (N_44677,N_43231,N_43453);
nor U44678 (N_44678,N_43526,N_43465);
xor U44679 (N_44679,N_43117,N_43176);
or U44680 (N_44680,N_43599,N_43838);
or U44681 (N_44681,N_43366,N_43663);
nor U44682 (N_44682,N_43584,N_43884);
or U44683 (N_44683,N_43379,N_43160);
or U44684 (N_44684,N_43632,N_43896);
and U44685 (N_44685,N_43548,N_43268);
nand U44686 (N_44686,N_43807,N_43605);
nor U44687 (N_44687,N_43944,N_43940);
nand U44688 (N_44688,N_43350,N_43007);
or U44689 (N_44689,N_43956,N_43967);
xnor U44690 (N_44690,N_43524,N_43653);
or U44691 (N_44691,N_43540,N_43415);
xor U44692 (N_44692,N_43690,N_43523);
nand U44693 (N_44693,N_43980,N_43669);
or U44694 (N_44694,N_43418,N_43783);
nand U44695 (N_44695,N_43137,N_43609);
nand U44696 (N_44696,N_43342,N_43484);
xnor U44697 (N_44697,N_43796,N_43910);
nand U44698 (N_44698,N_43535,N_43980);
or U44699 (N_44699,N_43030,N_43209);
or U44700 (N_44700,N_43064,N_43354);
and U44701 (N_44701,N_43819,N_43321);
xnor U44702 (N_44702,N_43893,N_43458);
xnor U44703 (N_44703,N_43422,N_43186);
or U44704 (N_44704,N_43058,N_43300);
nand U44705 (N_44705,N_43573,N_43023);
and U44706 (N_44706,N_43584,N_43277);
or U44707 (N_44707,N_43888,N_43718);
nand U44708 (N_44708,N_43467,N_43255);
or U44709 (N_44709,N_43484,N_43523);
and U44710 (N_44710,N_43082,N_43984);
nor U44711 (N_44711,N_43512,N_43855);
and U44712 (N_44712,N_43166,N_43297);
and U44713 (N_44713,N_43154,N_43911);
xnor U44714 (N_44714,N_43728,N_43754);
nand U44715 (N_44715,N_43854,N_43400);
nand U44716 (N_44716,N_43100,N_43068);
or U44717 (N_44717,N_43623,N_43868);
nand U44718 (N_44718,N_43591,N_43821);
xnor U44719 (N_44719,N_43417,N_43996);
xnor U44720 (N_44720,N_43898,N_43151);
nand U44721 (N_44721,N_43516,N_43119);
and U44722 (N_44722,N_43794,N_43342);
and U44723 (N_44723,N_43732,N_43270);
and U44724 (N_44724,N_43962,N_43470);
nand U44725 (N_44725,N_43306,N_43598);
xnor U44726 (N_44726,N_43267,N_43241);
xor U44727 (N_44727,N_43634,N_43528);
and U44728 (N_44728,N_43702,N_43159);
or U44729 (N_44729,N_43585,N_43852);
nor U44730 (N_44730,N_43759,N_43458);
nor U44731 (N_44731,N_43559,N_43442);
and U44732 (N_44732,N_43056,N_43387);
nand U44733 (N_44733,N_43983,N_43570);
xnor U44734 (N_44734,N_43984,N_43646);
and U44735 (N_44735,N_43419,N_43996);
nor U44736 (N_44736,N_43237,N_43182);
or U44737 (N_44737,N_43351,N_43390);
nand U44738 (N_44738,N_43859,N_43233);
and U44739 (N_44739,N_43120,N_43891);
nor U44740 (N_44740,N_43981,N_43464);
nor U44741 (N_44741,N_43557,N_43522);
nand U44742 (N_44742,N_43052,N_43518);
nand U44743 (N_44743,N_43717,N_43712);
nand U44744 (N_44744,N_43328,N_43078);
xor U44745 (N_44745,N_43447,N_43136);
or U44746 (N_44746,N_43162,N_43616);
and U44747 (N_44747,N_43449,N_43612);
nand U44748 (N_44748,N_43221,N_43316);
xor U44749 (N_44749,N_43452,N_43729);
xor U44750 (N_44750,N_43976,N_43272);
nor U44751 (N_44751,N_43648,N_43128);
and U44752 (N_44752,N_43490,N_43377);
xnor U44753 (N_44753,N_43093,N_43925);
nor U44754 (N_44754,N_43349,N_43154);
nand U44755 (N_44755,N_43211,N_43880);
nor U44756 (N_44756,N_43921,N_43023);
or U44757 (N_44757,N_43903,N_43339);
nand U44758 (N_44758,N_43895,N_43973);
or U44759 (N_44759,N_43279,N_43627);
nand U44760 (N_44760,N_43717,N_43533);
xnor U44761 (N_44761,N_43883,N_43754);
nor U44762 (N_44762,N_43234,N_43354);
nor U44763 (N_44763,N_43809,N_43413);
or U44764 (N_44764,N_43148,N_43403);
nor U44765 (N_44765,N_43269,N_43468);
or U44766 (N_44766,N_43368,N_43312);
and U44767 (N_44767,N_43658,N_43345);
nor U44768 (N_44768,N_43688,N_43249);
nand U44769 (N_44769,N_43440,N_43846);
or U44770 (N_44770,N_43462,N_43984);
xnor U44771 (N_44771,N_43943,N_43791);
nand U44772 (N_44772,N_43856,N_43845);
or U44773 (N_44773,N_43367,N_43170);
nand U44774 (N_44774,N_43113,N_43173);
xnor U44775 (N_44775,N_43217,N_43345);
xor U44776 (N_44776,N_43890,N_43541);
or U44777 (N_44777,N_43871,N_43428);
and U44778 (N_44778,N_43903,N_43219);
nand U44779 (N_44779,N_43434,N_43137);
and U44780 (N_44780,N_43821,N_43076);
xnor U44781 (N_44781,N_43599,N_43004);
and U44782 (N_44782,N_43328,N_43574);
xor U44783 (N_44783,N_43751,N_43481);
and U44784 (N_44784,N_43994,N_43029);
and U44785 (N_44785,N_43874,N_43990);
nand U44786 (N_44786,N_43889,N_43625);
and U44787 (N_44787,N_43795,N_43033);
xor U44788 (N_44788,N_43020,N_43094);
nand U44789 (N_44789,N_43137,N_43971);
nand U44790 (N_44790,N_43909,N_43142);
nand U44791 (N_44791,N_43593,N_43008);
nand U44792 (N_44792,N_43358,N_43855);
and U44793 (N_44793,N_43355,N_43698);
and U44794 (N_44794,N_43740,N_43842);
xor U44795 (N_44795,N_43530,N_43384);
nand U44796 (N_44796,N_43493,N_43408);
nand U44797 (N_44797,N_43334,N_43255);
or U44798 (N_44798,N_43130,N_43178);
or U44799 (N_44799,N_43976,N_43668);
xor U44800 (N_44800,N_43088,N_43202);
or U44801 (N_44801,N_43581,N_43373);
nand U44802 (N_44802,N_43787,N_43293);
nor U44803 (N_44803,N_43341,N_43477);
or U44804 (N_44804,N_43650,N_43027);
nand U44805 (N_44805,N_43885,N_43455);
nor U44806 (N_44806,N_43605,N_43077);
and U44807 (N_44807,N_43559,N_43392);
xnor U44808 (N_44808,N_43901,N_43096);
nor U44809 (N_44809,N_43547,N_43069);
nand U44810 (N_44810,N_43233,N_43451);
and U44811 (N_44811,N_43505,N_43160);
nand U44812 (N_44812,N_43977,N_43576);
or U44813 (N_44813,N_43958,N_43014);
or U44814 (N_44814,N_43182,N_43932);
xor U44815 (N_44815,N_43596,N_43328);
and U44816 (N_44816,N_43244,N_43663);
xor U44817 (N_44817,N_43601,N_43705);
nor U44818 (N_44818,N_43413,N_43009);
and U44819 (N_44819,N_43309,N_43936);
xnor U44820 (N_44820,N_43990,N_43219);
xnor U44821 (N_44821,N_43318,N_43579);
nor U44822 (N_44822,N_43431,N_43252);
or U44823 (N_44823,N_43671,N_43914);
nor U44824 (N_44824,N_43703,N_43078);
nor U44825 (N_44825,N_43920,N_43834);
xor U44826 (N_44826,N_43684,N_43793);
nor U44827 (N_44827,N_43649,N_43645);
nor U44828 (N_44828,N_43723,N_43192);
and U44829 (N_44829,N_43331,N_43657);
nor U44830 (N_44830,N_43665,N_43930);
nor U44831 (N_44831,N_43569,N_43440);
or U44832 (N_44832,N_43981,N_43973);
nand U44833 (N_44833,N_43144,N_43206);
and U44834 (N_44834,N_43324,N_43934);
nand U44835 (N_44835,N_43444,N_43278);
or U44836 (N_44836,N_43902,N_43767);
nand U44837 (N_44837,N_43326,N_43042);
nor U44838 (N_44838,N_43315,N_43123);
or U44839 (N_44839,N_43697,N_43269);
and U44840 (N_44840,N_43705,N_43225);
or U44841 (N_44841,N_43582,N_43067);
nand U44842 (N_44842,N_43816,N_43553);
or U44843 (N_44843,N_43740,N_43080);
xor U44844 (N_44844,N_43245,N_43085);
xor U44845 (N_44845,N_43495,N_43349);
or U44846 (N_44846,N_43363,N_43865);
and U44847 (N_44847,N_43357,N_43023);
nand U44848 (N_44848,N_43498,N_43016);
nand U44849 (N_44849,N_43020,N_43469);
xor U44850 (N_44850,N_43588,N_43849);
nor U44851 (N_44851,N_43458,N_43070);
xor U44852 (N_44852,N_43227,N_43416);
or U44853 (N_44853,N_43998,N_43249);
and U44854 (N_44854,N_43317,N_43237);
and U44855 (N_44855,N_43565,N_43865);
or U44856 (N_44856,N_43183,N_43515);
or U44857 (N_44857,N_43682,N_43448);
nand U44858 (N_44858,N_43949,N_43434);
xnor U44859 (N_44859,N_43372,N_43779);
xnor U44860 (N_44860,N_43490,N_43359);
or U44861 (N_44861,N_43209,N_43119);
and U44862 (N_44862,N_43430,N_43916);
xor U44863 (N_44863,N_43732,N_43485);
nor U44864 (N_44864,N_43852,N_43804);
xnor U44865 (N_44865,N_43965,N_43811);
nor U44866 (N_44866,N_43084,N_43801);
xor U44867 (N_44867,N_43937,N_43617);
xnor U44868 (N_44868,N_43217,N_43675);
nor U44869 (N_44869,N_43085,N_43061);
xnor U44870 (N_44870,N_43592,N_43890);
or U44871 (N_44871,N_43491,N_43755);
and U44872 (N_44872,N_43052,N_43384);
or U44873 (N_44873,N_43852,N_43868);
nand U44874 (N_44874,N_43893,N_43025);
nand U44875 (N_44875,N_43077,N_43596);
nand U44876 (N_44876,N_43186,N_43353);
or U44877 (N_44877,N_43132,N_43883);
and U44878 (N_44878,N_43314,N_43146);
nand U44879 (N_44879,N_43726,N_43437);
nor U44880 (N_44880,N_43388,N_43581);
xor U44881 (N_44881,N_43792,N_43428);
and U44882 (N_44882,N_43869,N_43264);
nand U44883 (N_44883,N_43956,N_43811);
nor U44884 (N_44884,N_43147,N_43273);
or U44885 (N_44885,N_43087,N_43128);
and U44886 (N_44886,N_43264,N_43500);
nor U44887 (N_44887,N_43452,N_43283);
xnor U44888 (N_44888,N_43349,N_43049);
and U44889 (N_44889,N_43140,N_43168);
or U44890 (N_44890,N_43976,N_43439);
and U44891 (N_44891,N_43640,N_43735);
xor U44892 (N_44892,N_43083,N_43836);
or U44893 (N_44893,N_43736,N_43860);
and U44894 (N_44894,N_43086,N_43854);
xor U44895 (N_44895,N_43477,N_43114);
nand U44896 (N_44896,N_43437,N_43325);
or U44897 (N_44897,N_43236,N_43862);
xor U44898 (N_44898,N_43435,N_43085);
and U44899 (N_44899,N_43851,N_43793);
nor U44900 (N_44900,N_43422,N_43358);
xor U44901 (N_44901,N_43537,N_43425);
nor U44902 (N_44902,N_43489,N_43198);
nor U44903 (N_44903,N_43836,N_43812);
and U44904 (N_44904,N_43827,N_43599);
xnor U44905 (N_44905,N_43610,N_43335);
nor U44906 (N_44906,N_43173,N_43181);
and U44907 (N_44907,N_43885,N_43627);
nand U44908 (N_44908,N_43857,N_43885);
nand U44909 (N_44909,N_43288,N_43590);
and U44910 (N_44910,N_43759,N_43324);
nor U44911 (N_44911,N_43547,N_43458);
or U44912 (N_44912,N_43958,N_43498);
nor U44913 (N_44913,N_43801,N_43577);
and U44914 (N_44914,N_43574,N_43608);
and U44915 (N_44915,N_43485,N_43770);
or U44916 (N_44916,N_43820,N_43694);
nand U44917 (N_44917,N_43354,N_43734);
nor U44918 (N_44918,N_43809,N_43767);
nor U44919 (N_44919,N_43130,N_43743);
nor U44920 (N_44920,N_43939,N_43779);
or U44921 (N_44921,N_43442,N_43377);
or U44922 (N_44922,N_43197,N_43549);
or U44923 (N_44923,N_43370,N_43380);
or U44924 (N_44924,N_43839,N_43076);
nor U44925 (N_44925,N_43632,N_43052);
nand U44926 (N_44926,N_43317,N_43592);
nor U44927 (N_44927,N_43922,N_43602);
and U44928 (N_44928,N_43809,N_43541);
nand U44929 (N_44929,N_43488,N_43428);
xnor U44930 (N_44930,N_43431,N_43934);
nand U44931 (N_44931,N_43417,N_43724);
nor U44932 (N_44932,N_43316,N_43107);
and U44933 (N_44933,N_43370,N_43566);
nand U44934 (N_44934,N_43419,N_43379);
nor U44935 (N_44935,N_43239,N_43041);
or U44936 (N_44936,N_43595,N_43175);
or U44937 (N_44937,N_43177,N_43557);
and U44938 (N_44938,N_43622,N_43486);
and U44939 (N_44939,N_43309,N_43289);
xor U44940 (N_44940,N_43709,N_43663);
nor U44941 (N_44941,N_43204,N_43508);
nor U44942 (N_44942,N_43722,N_43614);
or U44943 (N_44943,N_43580,N_43913);
or U44944 (N_44944,N_43715,N_43386);
xnor U44945 (N_44945,N_43326,N_43389);
and U44946 (N_44946,N_43756,N_43634);
nor U44947 (N_44947,N_43162,N_43606);
nand U44948 (N_44948,N_43101,N_43594);
and U44949 (N_44949,N_43732,N_43328);
and U44950 (N_44950,N_43558,N_43274);
nor U44951 (N_44951,N_43450,N_43553);
xnor U44952 (N_44952,N_43422,N_43372);
nand U44953 (N_44953,N_43922,N_43234);
and U44954 (N_44954,N_43689,N_43087);
nand U44955 (N_44955,N_43082,N_43446);
xnor U44956 (N_44956,N_43582,N_43321);
nand U44957 (N_44957,N_43874,N_43124);
xor U44958 (N_44958,N_43167,N_43401);
xnor U44959 (N_44959,N_43460,N_43933);
or U44960 (N_44960,N_43988,N_43824);
nor U44961 (N_44961,N_43518,N_43608);
nand U44962 (N_44962,N_43302,N_43358);
nor U44963 (N_44963,N_43957,N_43314);
and U44964 (N_44964,N_43275,N_43928);
or U44965 (N_44965,N_43362,N_43431);
or U44966 (N_44966,N_43721,N_43445);
xnor U44967 (N_44967,N_43093,N_43419);
xnor U44968 (N_44968,N_43360,N_43245);
or U44969 (N_44969,N_43684,N_43909);
or U44970 (N_44970,N_43910,N_43524);
and U44971 (N_44971,N_43850,N_43494);
nor U44972 (N_44972,N_43108,N_43010);
nand U44973 (N_44973,N_43141,N_43850);
or U44974 (N_44974,N_43195,N_43985);
nand U44975 (N_44975,N_43743,N_43183);
and U44976 (N_44976,N_43627,N_43113);
or U44977 (N_44977,N_43729,N_43980);
nand U44978 (N_44978,N_43552,N_43170);
or U44979 (N_44979,N_43193,N_43358);
xor U44980 (N_44980,N_43598,N_43765);
nor U44981 (N_44981,N_43104,N_43685);
and U44982 (N_44982,N_43995,N_43979);
and U44983 (N_44983,N_43863,N_43697);
nand U44984 (N_44984,N_43637,N_43358);
nand U44985 (N_44985,N_43506,N_43233);
nand U44986 (N_44986,N_43601,N_43875);
and U44987 (N_44987,N_43389,N_43317);
nor U44988 (N_44988,N_43773,N_43874);
or U44989 (N_44989,N_43127,N_43934);
and U44990 (N_44990,N_43327,N_43520);
or U44991 (N_44991,N_43133,N_43538);
xor U44992 (N_44992,N_43646,N_43820);
and U44993 (N_44993,N_43037,N_43506);
nand U44994 (N_44994,N_43490,N_43829);
xor U44995 (N_44995,N_43357,N_43328);
xor U44996 (N_44996,N_43392,N_43740);
nand U44997 (N_44997,N_43172,N_43433);
nor U44998 (N_44998,N_43424,N_43294);
nor U44999 (N_44999,N_43842,N_43157);
nand U45000 (N_45000,N_44842,N_44128);
nor U45001 (N_45001,N_44661,N_44628);
nand U45002 (N_45002,N_44277,N_44237);
or U45003 (N_45003,N_44226,N_44660);
nor U45004 (N_45004,N_44245,N_44504);
nand U45005 (N_45005,N_44167,N_44190);
or U45006 (N_45006,N_44044,N_44750);
nor U45007 (N_45007,N_44940,N_44895);
or U45008 (N_45008,N_44869,N_44333);
and U45009 (N_45009,N_44995,N_44948);
xor U45010 (N_45010,N_44028,N_44191);
and U45011 (N_45011,N_44789,N_44259);
or U45012 (N_45012,N_44486,N_44740);
and U45013 (N_45013,N_44032,N_44319);
nand U45014 (N_45014,N_44240,N_44563);
or U45015 (N_45015,N_44142,N_44324);
and U45016 (N_45016,N_44703,N_44357);
nor U45017 (N_45017,N_44623,N_44129);
nor U45018 (N_45018,N_44604,N_44217);
xnor U45019 (N_45019,N_44288,N_44861);
nand U45020 (N_45020,N_44805,N_44967);
nor U45021 (N_45021,N_44784,N_44701);
or U45022 (N_45022,N_44335,N_44408);
xnor U45023 (N_45023,N_44154,N_44951);
or U45024 (N_45024,N_44433,N_44111);
nor U45025 (N_45025,N_44689,N_44183);
and U45026 (N_45026,N_44531,N_44395);
nor U45027 (N_45027,N_44270,N_44428);
xor U45028 (N_45028,N_44492,N_44562);
nand U45029 (N_45029,N_44620,N_44204);
and U45030 (N_45030,N_44975,N_44748);
xnor U45031 (N_45031,N_44762,N_44373);
or U45032 (N_45032,N_44123,N_44530);
xor U45033 (N_45033,N_44806,N_44309);
nand U45034 (N_45034,N_44558,N_44077);
or U45035 (N_45035,N_44220,N_44688);
nor U45036 (N_45036,N_44365,N_44120);
and U45037 (N_45037,N_44591,N_44903);
xnor U45038 (N_45038,N_44389,N_44673);
nand U45039 (N_45039,N_44089,N_44606);
and U45040 (N_45040,N_44521,N_44051);
nand U45041 (N_45041,N_44140,N_44932);
and U45042 (N_45042,N_44300,N_44523);
or U45043 (N_45043,N_44043,N_44609);
nor U45044 (N_45044,N_44276,N_44117);
and U45045 (N_45045,N_44810,N_44901);
nor U45046 (N_45046,N_44543,N_44564);
xnor U45047 (N_45047,N_44060,N_44872);
xor U45048 (N_45048,N_44314,N_44105);
nand U45049 (N_45049,N_44496,N_44133);
nor U45050 (N_45050,N_44273,N_44616);
or U45051 (N_45051,N_44261,N_44739);
nor U45052 (N_45052,N_44802,N_44993);
xor U45053 (N_45053,N_44985,N_44144);
or U45054 (N_45054,N_44476,N_44378);
nor U45055 (N_45055,N_44159,N_44990);
nor U45056 (N_45056,N_44513,N_44196);
or U45057 (N_45057,N_44706,N_44090);
nand U45058 (N_45058,N_44075,N_44672);
nor U45059 (N_45059,N_44539,N_44532);
or U45060 (N_45060,N_44011,N_44691);
nand U45061 (N_45061,N_44526,N_44247);
nor U45062 (N_45062,N_44453,N_44037);
or U45063 (N_45063,N_44198,N_44731);
or U45064 (N_45064,N_44279,N_44393);
nor U45065 (N_45065,N_44696,N_44339);
or U45066 (N_45066,N_44832,N_44617);
or U45067 (N_45067,N_44738,N_44186);
xnor U45068 (N_45068,N_44219,N_44505);
or U45069 (N_45069,N_44960,N_44354);
and U45070 (N_45070,N_44836,N_44008);
or U45071 (N_45071,N_44329,N_44299);
nor U45072 (N_45072,N_44875,N_44068);
or U45073 (N_45073,N_44494,N_44886);
nand U45074 (N_45074,N_44094,N_44390);
nand U45075 (N_45075,N_44643,N_44361);
nand U45076 (N_45076,N_44624,N_44657);
nand U45077 (N_45077,N_44468,N_44902);
xor U45078 (N_45078,N_44430,N_44265);
and U45079 (N_45079,N_44405,N_44106);
nand U45080 (N_45080,N_44796,N_44537);
or U45081 (N_45081,N_44340,N_44404);
nand U45082 (N_45082,N_44423,N_44976);
and U45083 (N_45083,N_44596,N_44814);
and U45084 (N_45084,N_44500,N_44507);
nor U45085 (N_45085,N_44857,N_44310);
and U45086 (N_45086,N_44173,N_44846);
xor U45087 (N_45087,N_44798,N_44294);
nor U45088 (N_45088,N_44765,N_44388);
or U45089 (N_45089,N_44599,N_44027);
or U45090 (N_45090,N_44369,N_44344);
or U45091 (N_45091,N_44045,N_44488);
xor U45092 (N_45092,N_44171,N_44454);
nor U45093 (N_45093,N_44080,N_44004);
and U45094 (N_45094,N_44225,N_44224);
and U45095 (N_45095,N_44595,N_44029);
nand U45096 (N_45096,N_44398,N_44025);
nand U45097 (N_45097,N_44317,N_44269);
nor U45098 (N_45098,N_44356,N_44718);
nand U45099 (N_45099,N_44865,N_44401);
nor U45100 (N_45100,N_44293,N_44195);
and U45101 (N_45101,N_44939,N_44727);
and U45102 (N_45102,N_44424,N_44457);
nor U45103 (N_45103,N_44809,N_44947);
or U45104 (N_45104,N_44355,N_44753);
nor U45105 (N_45105,N_44728,N_44851);
and U45106 (N_45106,N_44502,N_44435);
or U45107 (N_45107,N_44193,N_44127);
and U45108 (N_45108,N_44399,N_44046);
or U45109 (N_45109,N_44296,N_44282);
nor U45110 (N_45110,N_44963,N_44916);
nand U45111 (N_45111,N_44443,N_44268);
xor U45112 (N_45112,N_44945,N_44135);
xnor U45113 (N_45113,N_44297,N_44066);
or U45114 (N_45114,N_44059,N_44612);
xnor U45115 (N_45115,N_44061,N_44725);
nand U45116 (N_45116,N_44954,N_44911);
or U45117 (N_45117,N_44803,N_44671);
nand U45118 (N_45118,N_44311,N_44455);
nor U45119 (N_45119,N_44113,N_44306);
or U45120 (N_45120,N_44284,N_44603);
nand U45121 (N_45121,N_44250,N_44848);
or U45122 (N_45122,N_44015,N_44651);
or U45123 (N_45123,N_44576,N_44447);
nor U45124 (N_45124,N_44347,N_44257);
nand U45125 (N_45125,N_44087,N_44464);
and U45126 (N_45126,N_44098,N_44376);
and U45127 (N_45127,N_44555,N_44790);
xnor U45128 (N_45128,N_44065,N_44601);
and U45129 (N_45129,N_44605,N_44438);
nand U45130 (N_45130,N_44209,N_44588);
and U45131 (N_45131,N_44574,N_44837);
xor U45132 (N_45132,N_44481,N_44808);
xnor U45133 (N_45133,N_44618,N_44637);
xor U45134 (N_45134,N_44343,N_44205);
nand U45135 (N_45135,N_44131,N_44763);
xor U45136 (N_45136,N_44002,N_44516);
or U45137 (N_45137,N_44881,N_44565);
nor U45138 (N_45138,N_44092,N_44999);
nand U45139 (N_45139,N_44348,N_44069);
nand U45140 (N_45140,N_44174,N_44958);
nor U45141 (N_45141,N_44473,N_44160);
or U45142 (N_45142,N_44503,N_44511);
xnor U45143 (N_45143,N_44444,N_44179);
nor U45144 (N_45144,N_44501,N_44049);
and U45145 (N_45145,N_44182,N_44654);
nor U45146 (N_45146,N_44082,N_44410);
nor U45147 (N_45147,N_44491,N_44716);
and U45148 (N_45148,N_44441,N_44286);
and U45149 (N_45149,N_44074,N_44017);
nand U45150 (N_45150,N_44819,N_44462);
and U45151 (N_45151,N_44560,N_44322);
nand U45152 (N_45152,N_44387,N_44783);
nor U45153 (N_45153,N_44943,N_44684);
nand U45154 (N_45154,N_44242,N_44307);
xnor U45155 (N_45155,N_44658,N_44996);
xnor U45156 (N_45156,N_44047,N_44134);
xnor U45157 (N_45157,N_44845,N_44546);
nand U45158 (N_45158,N_44368,N_44704);
or U45159 (N_45159,N_44289,N_44631);
and U45160 (N_45160,N_44328,N_44371);
nand U45161 (N_45161,N_44914,N_44550);
nand U45162 (N_45162,N_44165,N_44579);
xor U45163 (N_45163,N_44917,N_44653);
or U45164 (N_45164,N_44717,N_44295);
and U45165 (N_45165,N_44811,N_44692);
or U45166 (N_45166,N_44450,N_44417);
nor U45167 (N_45167,N_44570,N_44807);
or U45168 (N_45168,N_44013,N_44830);
xor U45169 (N_45169,N_44332,N_44681);
nor U45170 (N_45170,N_44346,N_44619);
nand U45171 (N_45171,N_44484,N_44122);
or U45172 (N_45172,N_44222,N_44206);
nor U45173 (N_45173,N_44164,N_44924);
nor U45174 (N_45174,N_44705,N_44714);
nor U45175 (N_45175,N_44583,N_44918);
nor U45176 (N_45176,N_44263,N_44062);
nand U45177 (N_45177,N_44452,N_44915);
or U45178 (N_45178,N_44909,N_44327);
nor U45179 (N_45179,N_44635,N_44093);
nand U45180 (N_45180,N_44187,N_44126);
xnor U45181 (N_45181,N_44936,N_44732);
nor U45182 (N_45182,N_44018,N_44253);
nor U45183 (N_45183,N_44866,N_44058);
or U45184 (N_45184,N_44774,N_44556);
nand U45185 (N_45185,N_44952,N_44188);
and U45186 (N_45186,N_44003,N_44412);
xnor U45187 (N_45187,N_44862,N_44192);
xor U45188 (N_45188,N_44370,N_44236);
nand U45189 (N_45189,N_44997,N_44634);
nand U45190 (N_45190,N_44930,N_44734);
or U45191 (N_45191,N_44971,N_44385);
nor U45192 (N_45192,N_44415,N_44359);
and U45193 (N_45193,N_44493,N_44034);
xnor U45194 (N_45194,N_44274,N_44112);
or U45195 (N_45195,N_44518,N_44463);
nor U45196 (N_45196,N_44699,N_44852);
xnor U45197 (N_45197,N_44019,N_44228);
or U45198 (N_45198,N_44573,N_44755);
xnor U45199 (N_45199,N_44031,N_44888);
and U45200 (N_45200,N_44650,N_44258);
nor U45201 (N_45201,N_44035,N_44229);
xor U45202 (N_45202,N_44157,N_44533);
xor U45203 (N_45203,N_44152,N_44207);
nand U45204 (N_45204,N_44668,N_44538);
and U45205 (N_45205,N_44337,N_44950);
nand U45206 (N_45206,N_44897,N_44782);
or U45207 (N_45207,N_44239,N_44168);
xnor U45208 (N_45208,N_44477,N_44694);
xor U45209 (N_45209,N_44384,N_44610);
xor U45210 (N_45210,N_44715,N_44214);
xor U45211 (N_45211,N_44325,N_44334);
nor U45212 (N_45212,N_44419,N_44956);
xor U45213 (N_45213,N_44038,N_44535);
or U45214 (N_45214,N_44291,N_44366);
or U45215 (N_45215,N_44099,N_44431);
nand U45216 (N_45216,N_44893,N_44422);
and U45217 (N_45217,N_44100,N_44965);
xnor U45218 (N_45218,N_44621,N_44854);
xor U45219 (N_45219,N_44115,N_44281);
and U45220 (N_45220,N_44891,N_44264);
and U45221 (N_45221,N_44267,N_44244);
xnor U45222 (N_45222,N_44665,N_44478);
xor U45223 (N_45223,N_44301,N_44973);
and U45224 (N_45224,N_44076,N_44949);
nor U45225 (N_45225,N_44998,N_44829);
nand U45226 (N_45226,N_44121,N_44780);
nor U45227 (N_45227,N_44561,N_44697);
and U45228 (N_45228,N_44552,N_44303);
nand U45229 (N_45229,N_44440,N_44312);
xor U45230 (N_45230,N_44858,N_44786);
nor U45231 (N_45231,N_44132,N_44735);
xor U45232 (N_45232,N_44839,N_44986);
xnor U45233 (N_45233,N_44683,N_44107);
or U45234 (N_45234,N_44506,N_44804);
and U45235 (N_45235,N_44772,N_44778);
and U45236 (N_45236,N_44921,N_44005);
and U45237 (N_45237,N_44828,N_44818);
and U45238 (N_45238,N_44754,N_44469);
nand U45239 (N_45239,N_44553,N_44156);
nand U45240 (N_45240,N_44906,N_44266);
nand U45241 (N_45241,N_44801,N_44280);
and U45242 (N_45242,N_44271,N_44073);
nand U45243 (N_45243,N_44372,N_44713);
xor U45244 (N_45244,N_44899,N_44146);
nor U45245 (N_45245,N_44109,N_44437);
and U45246 (N_45246,N_44812,N_44834);
nor U45247 (N_45247,N_44983,N_44172);
or U45248 (N_45248,N_44088,N_44639);
and U45249 (N_45249,N_44794,N_44321);
nand U45250 (N_45250,N_44770,N_44987);
nor U45251 (N_45251,N_44208,N_44912);
xor U45252 (N_45252,N_44232,N_44474);
xnor U45253 (N_45253,N_44544,N_44644);
xnor U45254 (N_45254,N_44568,N_44479);
nand U45255 (N_45255,N_44629,N_44036);
nor U45256 (N_45256,N_44012,N_44235);
and U45257 (N_45257,N_44723,N_44813);
and U45258 (N_45258,N_44498,N_44097);
xor U45259 (N_45259,N_44908,N_44425);
and U45260 (N_45260,N_44756,N_44730);
and U45261 (N_45261,N_44210,N_44680);
and U45262 (N_45262,N_44380,N_44542);
nand U45263 (N_45263,N_44548,N_44039);
nor U45264 (N_45264,N_44868,N_44460);
nand U45265 (N_45265,N_44984,N_44929);
xnor U45266 (N_45266,N_44085,N_44255);
nand U45267 (N_45267,N_44968,N_44181);
xnor U45268 (N_45268,N_44470,N_44592);
xor U45269 (N_45269,N_44040,N_44071);
or U45270 (N_45270,N_44345,N_44835);
xor U45271 (N_45271,N_44231,N_44323);
or U45272 (N_45272,N_44349,N_44305);
and U45273 (N_45273,N_44907,N_44508);
nor U45274 (N_45274,N_44519,N_44180);
nand U45275 (N_45275,N_44358,N_44178);
nor U45276 (N_45276,N_44795,N_44737);
nand U45277 (N_45277,N_44955,N_44449);
and U45278 (N_45278,N_44000,N_44820);
or U45279 (N_45279,N_44522,N_44840);
nand U45280 (N_45280,N_44655,N_44148);
xor U45281 (N_45281,N_44664,N_44988);
xnor U45282 (N_45282,N_44722,N_44104);
xnor U45283 (N_45283,N_44878,N_44768);
nand U45284 (N_45284,N_44981,N_44292);
and U45285 (N_45285,N_44095,N_44330);
or U45286 (N_45286,N_44194,N_44063);
and U45287 (N_45287,N_44625,N_44030);
nand U45288 (N_45288,N_44016,N_44429);
xnor U45289 (N_45289,N_44302,N_44145);
or U45290 (N_45290,N_44147,N_44243);
xor U45291 (N_45291,N_44760,N_44230);
xnor U45292 (N_45292,N_44776,N_44659);
nand U45293 (N_45293,N_44607,N_44557);
xor U45294 (N_45294,N_44890,N_44184);
and U45295 (N_45295,N_44248,N_44108);
nor U45296 (N_45296,N_44363,N_44517);
xnor U45297 (N_45297,N_44409,N_44992);
or U45298 (N_45298,N_44636,N_44793);
nand U45299 (N_45299,N_44042,N_44577);
or U45300 (N_45300,N_44392,N_44396);
xor U45301 (N_45301,N_44567,N_44391);
nor U45302 (N_45302,N_44685,N_44241);
nand U45303 (N_45303,N_44663,N_44726);
xnor U45304 (N_45304,N_44549,N_44767);
or U45305 (N_45305,N_44966,N_44456);
and U45306 (N_45306,N_44056,N_44054);
nand U45307 (N_45307,N_44375,N_44114);
xor U45308 (N_45308,N_44202,N_44642);
or U45309 (N_45309,N_44941,N_44448);
nor U45310 (N_45310,N_44761,N_44402);
nand U45311 (N_45311,N_44931,N_44033);
nand U45312 (N_45312,N_44649,N_44136);
nor U45313 (N_45313,N_44600,N_44843);
xnor U45314 (N_45314,N_44407,N_44926);
nor U45315 (N_45315,N_44693,N_44744);
nor U45316 (N_45316,N_44304,N_44024);
or U45317 (N_45317,N_44499,N_44101);
or U45318 (N_45318,N_44674,N_44153);
or U45319 (N_45319,N_44362,N_44969);
nand U45320 (N_45320,N_44510,N_44964);
nand U45321 (N_45321,N_44439,N_44382);
and U45322 (N_45322,N_44959,N_44775);
and U45323 (N_45323,N_44896,N_44850);
or U45324 (N_45324,N_44528,N_44887);
nor U45325 (N_45325,N_44260,N_44166);
or U45326 (N_45326,N_44615,N_44199);
xor U45327 (N_45327,N_44838,N_44551);
and U45328 (N_45328,N_44189,N_44442);
nor U45329 (N_45329,N_44055,N_44646);
or U45330 (N_45330,N_44495,N_44320);
or U45331 (N_45331,N_44158,N_44290);
and U45332 (N_45332,N_44471,N_44928);
nand U45333 (N_45333,N_44883,N_44072);
and U45334 (N_45334,N_44197,N_44420);
nor U45335 (N_45335,N_44249,N_44855);
nor U45336 (N_45336,N_44070,N_44877);
nor U45337 (N_45337,N_44844,N_44078);
xnor U45338 (N_45338,N_44707,N_44622);
nor U45339 (N_45339,N_44515,N_44386);
nor U45340 (N_45340,N_44451,N_44527);
or U45341 (N_45341,N_44894,N_44580);
and U45342 (N_45342,N_44741,N_44831);
or U45343 (N_45343,N_44406,N_44594);
nand U45344 (N_45344,N_44982,N_44991);
or U45345 (N_45345,N_44787,N_44006);
or U45346 (N_45346,N_44238,N_44566);
nand U45347 (N_45347,N_44149,N_44547);
nand U45348 (N_45348,N_44138,N_44632);
xor U45349 (N_45349,N_44213,N_44020);
and U45350 (N_45350,N_44298,N_44285);
nor U45351 (N_45351,N_44590,N_44151);
and U45352 (N_45352,N_44223,N_44934);
nand U45353 (N_45353,N_44514,N_44426);
or U45354 (N_45354,N_44667,N_44096);
or U45355 (N_45355,N_44125,N_44326);
nand U45356 (N_45356,N_44856,N_44185);
nor U45357 (N_45357,N_44743,N_44678);
and U45358 (N_45358,N_44086,N_44757);
nand U45359 (N_45359,N_44472,N_44081);
xnor U45360 (N_45360,N_44745,N_44638);
or U45361 (N_45361,N_44418,N_44962);
or U45362 (N_45362,N_44022,N_44010);
nor U45363 (N_45363,N_44816,N_44227);
or U45364 (N_45364,N_44690,N_44823);
and U45365 (N_45365,N_44394,N_44746);
xnor U45366 (N_45366,N_44175,N_44827);
and U45367 (N_45367,N_44880,N_44709);
nand U45368 (N_45368,N_44919,N_44465);
or U45369 (N_45369,N_44898,N_44920);
or U45370 (N_45370,N_44913,N_44432);
nor U45371 (N_45371,N_44489,N_44791);
nand U45372 (N_45372,N_44799,N_44524);
nand U45373 (N_45373,N_44825,N_44251);
and U45374 (N_45374,N_44377,N_44970);
nor U45375 (N_45375,N_44733,N_44262);
nand U45376 (N_45376,N_44053,N_44677);
or U45377 (N_45377,N_44884,N_44711);
nand U45378 (N_45378,N_44785,N_44233);
nor U45379 (N_45379,N_44067,N_44416);
nor U45380 (N_45380,N_44841,N_44922);
xnor U45381 (N_45381,N_44721,N_44421);
nor U45382 (N_45382,N_44118,N_44381);
xor U45383 (N_45383,N_44758,N_44467);
and U45384 (N_45384,N_44686,N_44788);
and U45385 (N_45385,N_44602,N_44598);
nor U45386 (N_45386,N_44720,N_44859);
xor U45387 (N_45387,N_44177,N_44860);
nand U45388 (N_45388,N_44079,N_44771);
nor U45389 (N_45389,N_44863,N_44352);
xor U45390 (N_45390,N_44351,N_44647);
nand U45391 (N_45391,N_44670,N_44490);
or U45392 (N_45392,N_44482,N_44218);
and U45393 (N_45393,N_44708,N_44091);
nand U45394 (N_45394,N_44041,N_44350);
nand U45395 (N_45395,N_44994,N_44162);
or U45396 (N_45396,N_44892,N_44800);
or U45397 (N_45397,N_44882,N_44139);
or U45398 (N_45398,N_44413,N_44001);
and U45399 (N_45399,N_44287,N_44545);
xor U45400 (N_45400,N_44626,N_44572);
and U45401 (N_45401,N_44700,N_44446);
nor U45402 (N_45402,N_44933,N_44586);
xnor U45403 (N_45403,N_44534,N_44459);
or U45404 (N_45404,N_44445,N_44752);
or U45405 (N_45405,N_44170,N_44978);
nor U45406 (N_45406,N_44614,N_44946);
xnor U45407 (N_45407,N_44211,N_44980);
xnor U45408 (N_45408,N_44215,N_44826);
and U45409 (N_45409,N_44052,N_44853);
and U45410 (N_45410,N_44427,N_44797);
or U45411 (N_45411,N_44318,N_44512);
and U45412 (N_45412,N_44953,N_44163);
or U45413 (N_45413,N_44742,N_44904);
nor U45414 (N_45414,N_44536,N_44710);
or U45415 (N_45415,N_44283,N_44736);
and U45416 (N_45416,N_44910,N_44316);
nand U45417 (N_45417,N_44766,N_44611);
nand U45418 (N_45418,N_44541,N_44870);
or U45419 (N_45419,N_44702,N_44308);
or U45420 (N_45420,N_44509,N_44341);
xor U45421 (N_45421,N_44749,N_44203);
and U45422 (N_45422,N_44083,N_44662);
nor U45423 (N_45423,N_44822,N_44792);
nor U45424 (N_45424,N_44379,N_44436);
or U45425 (N_45425,N_44764,N_44587);
and U45426 (N_45426,N_44821,N_44124);
or U45427 (N_45427,N_44695,N_44400);
and U45428 (N_45428,N_44905,N_44252);
nand U45429 (N_45429,N_44026,N_44064);
xnor U45430 (N_45430,N_44585,N_44169);
or U45431 (N_45431,N_44116,N_44640);
xnor U45432 (N_45432,N_44414,N_44777);
nand U45433 (N_45433,N_44216,N_44007);
xor U45434 (N_45434,N_44781,N_44925);
nor U45435 (N_45435,N_44497,N_44712);
and U45436 (N_45436,N_44889,N_44103);
and U45437 (N_45437,N_44937,N_44974);
or U45438 (N_45438,N_44682,N_44584);
nor U45439 (N_45439,N_44698,N_44520);
or U45440 (N_45440,N_44613,N_44155);
and U45441 (N_45441,N_44176,N_44212);
and U45442 (N_45442,N_44833,N_44961);
nor U45443 (N_45443,N_44221,N_44593);
xor U45444 (N_45444,N_44942,N_44687);
or U45445 (N_45445,N_44575,N_44719);
and U45446 (N_45446,N_44315,N_44729);
nand U45447 (N_45447,N_44938,N_44666);
or U45448 (N_45448,N_44525,N_44342);
or U45449 (N_45449,N_44589,N_44675);
nor U45450 (N_45450,N_44608,N_44989);
xnor U45451 (N_45451,N_44141,N_44669);
or U45452 (N_45452,N_44313,N_44272);
and U45453 (N_45453,N_44540,N_44057);
nand U45454 (N_45454,N_44254,N_44397);
xnor U45455 (N_45455,N_44652,N_44630);
nand U45456 (N_45456,N_44724,N_44201);
and U45457 (N_45457,N_44374,N_44403);
xnor U45458 (N_45458,N_44084,N_44234);
nor U45459 (N_45459,N_44871,N_44773);
and U45460 (N_45460,N_44256,N_44648);
nor U45461 (N_45461,N_44367,N_44466);
and U45462 (N_45462,N_44014,N_44458);
nand U45463 (N_45463,N_44383,N_44483);
nor U45464 (N_45464,N_44487,N_44867);
or U45465 (N_45465,N_44885,N_44627);
xnor U45466 (N_45466,N_44353,N_44569);
nor U45467 (N_45467,N_44102,N_44246);
and U45468 (N_45468,N_44009,N_44864);
xor U45469 (N_45469,N_44957,N_44360);
and U45470 (N_45470,N_44559,N_44150);
or U45471 (N_45471,N_44048,N_44137);
or U45472 (N_45472,N_44571,N_44977);
nor U45473 (N_45473,N_44847,N_44923);
or U45474 (N_45474,N_44751,N_44597);
or U45475 (N_45475,N_44050,N_44879);
xor U45476 (N_45476,N_44769,N_44900);
xor U45477 (N_45477,N_44759,N_44434);
xor U45478 (N_45478,N_44979,N_44200);
nand U45479 (N_45479,N_44972,N_44656);
nand U45480 (N_45480,N_44161,N_44935);
nor U45481 (N_45481,N_44475,N_44278);
nor U45482 (N_45482,N_44143,N_44824);
nor U45483 (N_45483,N_44336,N_44581);
xnor U45484 (N_45484,N_44633,N_44331);
or U45485 (N_45485,N_44461,N_44817);
nor U45486 (N_45486,N_44338,N_44876);
xor U45487 (N_45487,N_44021,N_44944);
and U45488 (N_45488,N_44485,N_44873);
nor U45489 (N_45489,N_44676,N_44582);
and U45490 (N_45490,N_44779,N_44874);
or U45491 (N_45491,N_44849,N_44023);
and U45492 (N_45492,N_44815,N_44130);
xor U45493 (N_45493,N_44110,N_44641);
or U45494 (N_45494,N_44364,N_44679);
nor U45495 (N_45495,N_44554,N_44480);
xnor U45496 (N_45496,N_44275,N_44747);
and U45497 (N_45497,N_44119,N_44927);
or U45498 (N_45498,N_44578,N_44529);
and U45499 (N_45499,N_44645,N_44411);
and U45500 (N_45500,N_44240,N_44302);
nand U45501 (N_45501,N_44992,N_44035);
nor U45502 (N_45502,N_44347,N_44268);
or U45503 (N_45503,N_44057,N_44551);
and U45504 (N_45504,N_44650,N_44914);
and U45505 (N_45505,N_44420,N_44918);
or U45506 (N_45506,N_44714,N_44414);
nor U45507 (N_45507,N_44620,N_44744);
and U45508 (N_45508,N_44746,N_44188);
xnor U45509 (N_45509,N_44151,N_44155);
xor U45510 (N_45510,N_44658,N_44735);
and U45511 (N_45511,N_44633,N_44693);
nor U45512 (N_45512,N_44428,N_44702);
or U45513 (N_45513,N_44309,N_44294);
nor U45514 (N_45514,N_44176,N_44963);
xnor U45515 (N_45515,N_44210,N_44609);
nand U45516 (N_45516,N_44825,N_44252);
nor U45517 (N_45517,N_44686,N_44571);
nor U45518 (N_45518,N_44546,N_44745);
xor U45519 (N_45519,N_44244,N_44154);
or U45520 (N_45520,N_44015,N_44437);
xnor U45521 (N_45521,N_44153,N_44114);
nand U45522 (N_45522,N_44740,N_44016);
nor U45523 (N_45523,N_44952,N_44895);
or U45524 (N_45524,N_44695,N_44117);
or U45525 (N_45525,N_44999,N_44459);
and U45526 (N_45526,N_44133,N_44583);
xor U45527 (N_45527,N_44922,N_44335);
xor U45528 (N_45528,N_44329,N_44523);
xnor U45529 (N_45529,N_44438,N_44582);
xor U45530 (N_45530,N_44329,N_44951);
nand U45531 (N_45531,N_44713,N_44615);
or U45532 (N_45532,N_44926,N_44176);
xnor U45533 (N_45533,N_44658,N_44742);
or U45534 (N_45534,N_44823,N_44434);
and U45535 (N_45535,N_44530,N_44458);
nand U45536 (N_45536,N_44450,N_44277);
or U45537 (N_45537,N_44698,N_44982);
nor U45538 (N_45538,N_44183,N_44312);
or U45539 (N_45539,N_44113,N_44906);
nor U45540 (N_45540,N_44219,N_44962);
nor U45541 (N_45541,N_44434,N_44089);
nor U45542 (N_45542,N_44049,N_44334);
nand U45543 (N_45543,N_44976,N_44213);
or U45544 (N_45544,N_44047,N_44556);
and U45545 (N_45545,N_44089,N_44608);
nor U45546 (N_45546,N_44952,N_44230);
nor U45547 (N_45547,N_44588,N_44384);
xor U45548 (N_45548,N_44281,N_44357);
nand U45549 (N_45549,N_44787,N_44798);
or U45550 (N_45550,N_44117,N_44465);
nor U45551 (N_45551,N_44766,N_44244);
nor U45552 (N_45552,N_44921,N_44606);
nand U45553 (N_45553,N_44238,N_44612);
nand U45554 (N_45554,N_44421,N_44176);
and U45555 (N_45555,N_44195,N_44689);
or U45556 (N_45556,N_44842,N_44340);
and U45557 (N_45557,N_44592,N_44058);
nand U45558 (N_45558,N_44191,N_44217);
and U45559 (N_45559,N_44835,N_44715);
nand U45560 (N_45560,N_44399,N_44587);
nor U45561 (N_45561,N_44489,N_44229);
nor U45562 (N_45562,N_44580,N_44453);
xor U45563 (N_45563,N_44617,N_44035);
xnor U45564 (N_45564,N_44914,N_44947);
or U45565 (N_45565,N_44993,N_44510);
nand U45566 (N_45566,N_44850,N_44468);
nand U45567 (N_45567,N_44600,N_44154);
nor U45568 (N_45568,N_44902,N_44257);
or U45569 (N_45569,N_44350,N_44665);
nor U45570 (N_45570,N_44949,N_44540);
nand U45571 (N_45571,N_44437,N_44356);
and U45572 (N_45572,N_44491,N_44477);
nor U45573 (N_45573,N_44306,N_44942);
and U45574 (N_45574,N_44312,N_44434);
nand U45575 (N_45575,N_44560,N_44957);
and U45576 (N_45576,N_44360,N_44231);
nor U45577 (N_45577,N_44469,N_44659);
and U45578 (N_45578,N_44742,N_44385);
and U45579 (N_45579,N_44066,N_44342);
nand U45580 (N_45580,N_44502,N_44633);
nor U45581 (N_45581,N_44807,N_44688);
or U45582 (N_45582,N_44351,N_44944);
xnor U45583 (N_45583,N_44278,N_44793);
or U45584 (N_45584,N_44652,N_44486);
xnor U45585 (N_45585,N_44798,N_44429);
nand U45586 (N_45586,N_44646,N_44822);
nand U45587 (N_45587,N_44528,N_44714);
xnor U45588 (N_45588,N_44580,N_44224);
nor U45589 (N_45589,N_44781,N_44470);
xor U45590 (N_45590,N_44866,N_44476);
and U45591 (N_45591,N_44266,N_44419);
or U45592 (N_45592,N_44078,N_44104);
or U45593 (N_45593,N_44148,N_44881);
and U45594 (N_45594,N_44874,N_44574);
xor U45595 (N_45595,N_44147,N_44142);
or U45596 (N_45596,N_44970,N_44922);
nor U45597 (N_45597,N_44566,N_44283);
or U45598 (N_45598,N_44782,N_44478);
or U45599 (N_45599,N_44090,N_44967);
and U45600 (N_45600,N_44971,N_44300);
or U45601 (N_45601,N_44572,N_44691);
nor U45602 (N_45602,N_44337,N_44298);
nor U45603 (N_45603,N_44499,N_44765);
nand U45604 (N_45604,N_44135,N_44143);
or U45605 (N_45605,N_44470,N_44964);
nor U45606 (N_45606,N_44622,N_44384);
and U45607 (N_45607,N_44060,N_44963);
nor U45608 (N_45608,N_44794,N_44332);
nor U45609 (N_45609,N_44891,N_44827);
or U45610 (N_45610,N_44664,N_44317);
nand U45611 (N_45611,N_44476,N_44916);
nand U45612 (N_45612,N_44817,N_44929);
xor U45613 (N_45613,N_44005,N_44261);
nor U45614 (N_45614,N_44726,N_44201);
and U45615 (N_45615,N_44956,N_44641);
or U45616 (N_45616,N_44868,N_44262);
xor U45617 (N_45617,N_44288,N_44939);
or U45618 (N_45618,N_44705,N_44538);
xor U45619 (N_45619,N_44066,N_44370);
or U45620 (N_45620,N_44094,N_44541);
nor U45621 (N_45621,N_44734,N_44988);
xor U45622 (N_45622,N_44129,N_44848);
nand U45623 (N_45623,N_44894,N_44688);
nor U45624 (N_45624,N_44215,N_44985);
xnor U45625 (N_45625,N_44626,N_44595);
nor U45626 (N_45626,N_44703,N_44272);
and U45627 (N_45627,N_44121,N_44877);
nor U45628 (N_45628,N_44206,N_44194);
nor U45629 (N_45629,N_44180,N_44382);
and U45630 (N_45630,N_44399,N_44979);
nor U45631 (N_45631,N_44388,N_44984);
or U45632 (N_45632,N_44938,N_44974);
nand U45633 (N_45633,N_44650,N_44719);
xnor U45634 (N_45634,N_44933,N_44629);
xor U45635 (N_45635,N_44838,N_44427);
nor U45636 (N_45636,N_44161,N_44715);
or U45637 (N_45637,N_44058,N_44999);
or U45638 (N_45638,N_44132,N_44533);
nor U45639 (N_45639,N_44798,N_44805);
nor U45640 (N_45640,N_44443,N_44936);
nand U45641 (N_45641,N_44785,N_44407);
or U45642 (N_45642,N_44345,N_44453);
and U45643 (N_45643,N_44878,N_44092);
nor U45644 (N_45644,N_44894,N_44576);
or U45645 (N_45645,N_44414,N_44513);
and U45646 (N_45646,N_44554,N_44985);
and U45647 (N_45647,N_44845,N_44437);
or U45648 (N_45648,N_44363,N_44665);
nor U45649 (N_45649,N_44298,N_44720);
and U45650 (N_45650,N_44803,N_44055);
or U45651 (N_45651,N_44935,N_44060);
or U45652 (N_45652,N_44111,N_44465);
xor U45653 (N_45653,N_44121,N_44879);
xor U45654 (N_45654,N_44923,N_44415);
and U45655 (N_45655,N_44681,N_44771);
and U45656 (N_45656,N_44957,N_44998);
xnor U45657 (N_45657,N_44128,N_44392);
or U45658 (N_45658,N_44139,N_44723);
and U45659 (N_45659,N_44966,N_44057);
nand U45660 (N_45660,N_44219,N_44690);
xor U45661 (N_45661,N_44063,N_44825);
xor U45662 (N_45662,N_44995,N_44562);
nor U45663 (N_45663,N_44902,N_44807);
or U45664 (N_45664,N_44355,N_44295);
nand U45665 (N_45665,N_44320,N_44477);
nor U45666 (N_45666,N_44938,N_44018);
xor U45667 (N_45667,N_44073,N_44952);
xnor U45668 (N_45668,N_44723,N_44049);
and U45669 (N_45669,N_44701,N_44697);
nand U45670 (N_45670,N_44649,N_44233);
or U45671 (N_45671,N_44457,N_44228);
and U45672 (N_45672,N_44802,N_44424);
nor U45673 (N_45673,N_44050,N_44854);
xor U45674 (N_45674,N_44364,N_44627);
and U45675 (N_45675,N_44747,N_44386);
and U45676 (N_45676,N_44508,N_44999);
or U45677 (N_45677,N_44453,N_44576);
nand U45678 (N_45678,N_44046,N_44606);
and U45679 (N_45679,N_44464,N_44397);
or U45680 (N_45680,N_44904,N_44937);
nor U45681 (N_45681,N_44123,N_44926);
and U45682 (N_45682,N_44901,N_44052);
and U45683 (N_45683,N_44006,N_44916);
xnor U45684 (N_45684,N_44173,N_44888);
xnor U45685 (N_45685,N_44060,N_44094);
and U45686 (N_45686,N_44819,N_44321);
nand U45687 (N_45687,N_44894,N_44572);
xnor U45688 (N_45688,N_44805,N_44244);
xnor U45689 (N_45689,N_44344,N_44803);
or U45690 (N_45690,N_44543,N_44082);
and U45691 (N_45691,N_44373,N_44090);
xnor U45692 (N_45692,N_44314,N_44950);
or U45693 (N_45693,N_44440,N_44547);
or U45694 (N_45694,N_44348,N_44365);
xnor U45695 (N_45695,N_44086,N_44977);
nand U45696 (N_45696,N_44052,N_44632);
or U45697 (N_45697,N_44228,N_44100);
nor U45698 (N_45698,N_44079,N_44927);
and U45699 (N_45699,N_44689,N_44009);
and U45700 (N_45700,N_44764,N_44773);
xor U45701 (N_45701,N_44045,N_44054);
nor U45702 (N_45702,N_44339,N_44757);
nor U45703 (N_45703,N_44535,N_44721);
nor U45704 (N_45704,N_44816,N_44942);
nand U45705 (N_45705,N_44307,N_44068);
and U45706 (N_45706,N_44396,N_44815);
or U45707 (N_45707,N_44655,N_44220);
and U45708 (N_45708,N_44559,N_44711);
xor U45709 (N_45709,N_44065,N_44747);
or U45710 (N_45710,N_44507,N_44064);
or U45711 (N_45711,N_44385,N_44520);
or U45712 (N_45712,N_44112,N_44549);
xor U45713 (N_45713,N_44581,N_44181);
nand U45714 (N_45714,N_44666,N_44095);
nand U45715 (N_45715,N_44115,N_44652);
or U45716 (N_45716,N_44072,N_44704);
nor U45717 (N_45717,N_44648,N_44972);
or U45718 (N_45718,N_44023,N_44337);
nor U45719 (N_45719,N_44623,N_44890);
nand U45720 (N_45720,N_44804,N_44057);
and U45721 (N_45721,N_44463,N_44118);
xor U45722 (N_45722,N_44373,N_44503);
or U45723 (N_45723,N_44978,N_44224);
xnor U45724 (N_45724,N_44749,N_44272);
xnor U45725 (N_45725,N_44767,N_44132);
and U45726 (N_45726,N_44765,N_44877);
nor U45727 (N_45727,N_44236,N_44320);
nor U45728 (N_45728,N_44717,N_44948);
and U45729 (N_45729,N_44707,N_44647);
nand U45730 (N_45730,N_44462,N_44761);
xnor U45731 (N_45731,N_44227,N_44394);
nand U45732 (N_45732,N_44129,N_44488);
nor U45733 (N_45733,N_44711,N_44802);
and U45734 (N_45734,N_44293,N_44058);
or U45735 (N_45735,N_44503,N_44743);
nor U45736 (N_45736,N_44860,N_44675);
or U45737 (N_45737,N_44844,N_44676);
nand U45738 (N_45738,N_44467,N_44340);
or U45739 (N_45739,N_44477,N_44447);
xnor U45740 (N_45740,N_44642,N_44491);
and U45741 (N_45741,N_44543,N_44815);
nor U45742 (N_45742,N_44577,N_44730);
xnor U45743 (N_45743,N_44201,N_44477);
or U45744 (N_45744,N_44519,N_44824);
nor U45745 (N_45745,N_44095,N_44721);
nand U45746 (N_45746,N_44672,N_44933);
or U45747 (N_45747,N_44092,N_44720);
or U45748 (N_45748,N_44459,N_44508);
and U45749 (N_45749,N_44196,N_44874);
nor U45750 (N_45750,N_44040,N_44658);
and U45751 (N_45751,N_44743,N_44032);
nand U45752 (N_45752,N_44523,N_44395);
nor U45753 (N_45753,N_44862,N_44565);
xnor U45754 (N_45754,N_44195,N_44187);
nor U45755 (N_45755,N_44841,N_44021);
nand U45756 (N_45756,N_44450,N_44727);
xnor U45757 (N_45757,N_44484,N_44780);
xnor U45758 (N_45758,N_44120,N_44805);
xor U45759 (N_45759,N_44750,N_44117);
xnor U45760 (N_45760,N_44367,N_44138);
nand U45761 (N_45761,N_44647,N_44501);
and U45762 (N_45762,N_44234,N_44514);
or U45763 (N_45763,N_44308,N_44850);
nand U45764 (N_45764,N_44721,N_44747);
or U45765 (N_45765,N_44620,N_44267);
xor U45766 (N_45766,N_44624,N_44868);
nand U45767 (N_45767,N_44622,N_44059);
and U45768 (N_45768,N_44907,N_44906);
nor U45769 (N_45769,N_44228,N_44832);
nand U45770 (N_45770,N_44183,N_44650);
xor U45771 (N_45771,N_44971,N_44170);
nand U45772 (N_45772,N_44576,N_44031);
or U45773 (N_45773,N_44593,N_44650);
and U45774 (N_45774,N_44432,N_44063);
xnor U45775 (N_45775,N_44487,N_44052);
xor U45776 (N_45776,N_44086,N_44947);
nor U45777 (N_45777,N_44049,N_44777);
or U45778 (N_45778,N_44975,N_44114);
nor U45779 (N_45779,N_44450,N_44053);
or U45780 (N_45780,N_44450,N_44939);
and U45781 (N_45781,N_44666,N_44561);
nor U45782 (N_45782,N_44693,N_44968);
xor U45783 (N_45783,N_44273,N_44810);
or U45784 (N_45784,N_44112,N_44982);
nand U45785 (N_45785,N_44461,N_44276);
nand U45786 (N_45786,N_44842,N_44519);
and U45787 (N_45787,N_44287,N_44726);
or U45788 (N_45788,N_44908,N_44409);
nor U45789 (N_45789,N_44171,N_44722);
or U45790 (N_45790,N_44958,N_44847);
xor U45791 (N_45791,N_44295,N_44065);
or U45792 (N_45792,N_44247,N_44749);
and U45793 (N_45793,N_44986,N_44793);
nand U45794 (N_45794,N_44268,N_44875);
or U45795 (N_45795,N_44745,N_44901);
xor U45796 (N_45796,N_44124,N_44084);
nand U45797 (N_45797,N_44946,N_44468);
or U45798 (N_45798,N_44008,N_44943);
or U45799 (N_45799,N_44286,N_44256);
or U45800 (N_45800,N_44329,N_44774);
xnor U45801 (N_45801,N_44947,N_44759);
nor U45802 (N_45802,N_44714,N_44387);
or U45803 (N_45803,N_44960,N_44099);
nand U45804 (N_45804,N_44083,N_44837);
and U45805 (N_45805,N_44801,N_44445);
and U45806 (N_45806,N_44882,N_44342);
or U45807 (N_45807,N_44560,N_44833);
nand U45808 (N_45808,N_44162,N_44039);
nor U45809 (N_45809,N_44975,N_44858);
xnor U45810 (N_45810,N_44100,N_44422);
nor U45811 (N_45811,N_44509,N_44609);
xor U45812 (N_45812,N_44849,N_44856);
xor U45813 (N_45813,N_44721,N_44976);
and U45814 (N_45814,N_44548,N_44679);
nor U45815 (N_45815,N_44395,N_44833);
nor U45816 (N_45816,N_44897,N_44091);
xor U45817 (N_45817,N_44409,N_44895);
nor U45818 (N_45818,N_44293,N_44324);
or U45819 (N_45819,N_44070,N_44853);
and U45820 (N_45820,N_44322,N_44627);
nor U45821 (N_45821,N_44254,N_44512);
xor U45822 (N_45822,N_44659,N_44493);
xnor U45823 (N_45823,N_44179,N_44883);
nor U45824 (N_45824,N_44084,N_44205);
nand U45825 (N_45825,N_44778,N_44301);
and U45826 (N_45826,N_44776,N_44974);
and U45827 (N_45827,N_44873,N_44769);
and U45828 (N_45828,N_44716,N_44058);
nand U45829 (N_45829,N_44481,N_44320);
nor U45830 (N_45830,N_44579,N_44005);
and U45831 (N_45831,N_44971,N_44830);
nor U45832 (N_45832,N_44479,N_44021);
xnor U45833 (N_45833,N_44344,N_44200);
xnor U45834 (N_45834,N_44738,N_44278);
nor U45835 (N_45835,N_44810,N_44281);
nand U45836 (N_45836,N_44588,N_44284);
nand U45837 (N_45837,N_44997,N_44945);
nor U45838 (N_45838,N_44292,N_44603);
xor U45839 (N_45839,N_44072,N_44810);
nor U45840 (N_45840,N_44326,N_44914);
or U45841 (N_45841,N_44168,N_44559);
or U45842 (N_45842,N_44025,N_44530);
nor U45843 (N_45843,N_44369,N_44676);
nand U45844 (N_45844,N_44703,N_44096);
nand U45845 (N_45845,N_44301,N_44172);
or U45846 (N_45846,N_44914,N_44653);
nor U45847 (N_45847,N_44863,N_44913);
xnor U45848 (N_45848,N_44359,N_44715);
or U45849 (N_45849,N_44873,N_44621);
xnor U45850 (N_45850,N_44786,N_44641);
xor U45851 (N_45851,N_44928,N_44733);
or U45852 (N_45852,N_44320,N_44737);
xnor U45853 (N_45853,N_44625,N_44469);
xnor U45854 (N_45854,N_44791,N_44616);
xnor U45855 (N_45855,N_44156,N_44619);
nor U45856 (N_45856,N_44015,N_44186);
nand U45857 (N_45857,N_44199,N_44396);
nor U45858 (N_45858,N_44016,N_44561);
and U45859 (N_45859,N_44622,N_44029);
or U45860 (N_45860,N_44450,N_44684);
nor U45861 (N_45861,N_44108,N_44267);
xnor U45862 (N_45862,N_44731,N_44085);
xnor U45863 (N_45863,N_44685,N_44476);
and U45864 (N_45864,N_44972,N_44216);
nand U45865 (N_45865,N_44757,N_44122);
nor U45866 (N_45866,N_44813,N_44852);
nor U45867 (N_45867,N_44708,N_44579);
nand U45868 (N_45868,N_44111,N_44374);
nand U45869 (N_45869,N_44752,N_44075);
xor U45870 (N_45870,N_44956,N_44729);
nand U45871 (N_45871,N_44171,N_44063);
xnor U45872 (N_45872,N_44018,N_44614);
xnor U45873 (N_45873,N_44904,N_44706);
and U45874 (N_45874,N_44905,N_44069);
xnor U45875 (N_45875,N_44892,N_44345);
and U45876 (N_45876,N_44570,N_44160);
and U45877 (N_45877,N_44773,N_44201);
nor U45878 (N_45878,N_44648,N_44824);
xnor U45879 (N_45879,N_44396,N_44783);
or U45880 (N_45880,N_44518,N_44742);
or U45881 (N_45881,N_44967,N_44530);
and U45882 (N_45882,N_44295,N_44689);
or U45883 (N_45883,N_44307,N_44837);
xnor U45884 (N_45884,N_44397,N_44181);
xor U45885 (N_45885,N_44988,N_44306);
xnor U45886 (N_45886,N_44359,N_44548);
xor U45887 (N_45887,N_44993,N_44883);
xnor U45888 (N_45888,N_44340,N_44978);
xor U45889 (N_45889,N_44950,N_44014);
and U45890 (N_45890,N_44294,N_44856);
nor U45891 (N_45891,N_44928,N_44432);
xor U45892 (N_45892,N_44920,N_44582);
and U45893 (N_45893,N_44376,N_44219);
nor U45894 (N_45894,N_44383,N_44318);
and U45895 (N_45895,N_44082,N_44701);
xor U45896 (N_45896,N_44109,N_44965);
xnor U45897 (N_45897,N_44705,N_44629);
nand U45898 (N_45898,N_44189,N_44124);
or U45899 (N_45899,N_44818,N_44181);
and U45900 (N_45900,N_44271,N_44316);
or U45901 (N_45901,N_44020,N_44065);
xor U45902 (N_45902,N_44662,N_44345);
and U45903 (N_45903,N_44833,N_44250);
nor U45904 (N_45904,N_44724,N_44424);
xor U45905 (N_45905,N_44116,N_44282);
xor U45906 (N_45906,N_44678,N_44000);
nand U45907 (N_45907,N_44097,N_44739);
nor U45908 (N_45908,N_44626,N_44593);
and U45909 (N_45909,N_44131,N_44486);
xnor U45910 (N_45910,N_44422,N_44202);
nor U45911 (N_45911,N_44799,N_44641);
and U45912 (N_45912,N_44239,N_44091);
and U45913 (N_45913,N_44653,N_44380);
xnor U45914 (N_45914,N_44291,N_44167);
or U45915 (N_45915,N_44254,N_44878);
or U45916 (N_45916,N_44709,N_44083);
nand U45917 (N_45917,N_44441,N_44926);
xnor U45918 (N_45918,N_44730,N_44293);
nand U45919 (N_45919,N_44129,N_44291);
or U45920 (N_45920,N_44633,N_44893);
nor U45921 (N_45921,N_44372,N_44339);
nor U45922 (N_45922,N_44078,N_44724);
or U45923 (N_45923,N_44636,N_44271);
xnor U45924 (N_45924,N_44970,N_44186);
and U45925 (N_45925,N_44067,N_44841);
nand U45926 (N_45926,N_44844,N_44477);
or U45927 (N_45927,N_44106,N_44179);
nand U45928 (N_45928,N_44108,N_44041);
or U45929 (N_45929,N_44683,N_44928);
nand U45930 (N_45930,N_44267,N_44854);
nand U45931 (N_45931,N_44257,N_44416);
nand U45932 (N_45932,N_44933,N_44126);
or U45933 (N_45933,N_44350,N_44391);
xor U45934 (N_45934,N_44946,N_44400);
or U45935 (N_45935,N_44821,N_44541);
nor U45936 (N_45936,N_44817,N_44853);
nand U45937 (N_45937,N_44769,N_44824);
or U45938 (N_45938,N_44620,N_44294);
and U45939 (N_45939,N_44540,N_44891);
nand U45940 (N_45940,N_44780,N_44538);
and U45941 (N_45941,N_44528,N_44795);
nor U45942 (N_45942,N_44211,N_44633);
and U45943 (N_45943,N_44335,N_44708);
and U45944 (N_45944,N_44091,N_44749);
or U45945 (N_45945,N_44504,N_44630);
and U45946 (N_45946,N_44877,N_44253);
nor U45947 (N_45947,N_44669,N_44749);
xor U45948 (N_45948,N_44773,N_44666);
and U45949 (N_45949,N_44618,N_44231);
or U45950 (N_45950,N_44371,N_44690);
xnor U45951 (N_45951,N_44228,N_44315);
nor U45952 (N_45952,N_44610,N_44432);
xor U45953 (N_45953,N_44355,N_44259);
or U45954 (N_45954,N_44961,N_44097);
xnor U45955 (N_45955,N_44172,N_44554);
or U45956 (N_45956,N_44994,N_44958);
or U45957 (N_45957,N_44648,N_44436);
and U45958 (N_45958,N_44378,N_44794);
nor U45959 (N_45959,N_44098,N_44166);
or U45960 (N_45960,N_44336,N_44978);
nand U45961 (N_45961,N_44327,N_44444);
nand U45962 (N_45962,N_44697,N_44092);
xnor U45963 (N_45963,N_44075,N_44446);
xor U45964 (N_45964,N_44870,N_44558);
nor U45965 (N_45965,N_44779,N_44348);
or U45966 (N_45966,N_44718,N_44615);
xor U45967 (N_45967,N_44185,N_44024);
or U45968 (N_45968,N_44745,N_44478);
nand U45969 (N_45969,N_44469,N_44551);
or U45970 (N_45970,N_44762,N_44455);
and U45971 (N_45971,N_44037,N_44169);
or U45972 (N_45972,N_44605,N_44198);
or U45973 (N_45973,N_44021,N_44984);
or U45974 (N_45974,N_44220,N_44609);
nand U45975 (N_45975,N_44527,N_44184);
nor U45976 (N_45976,N_44970,N_44613);
xnor U45977 (N_45977,N_44045,N_44111);
nor U45978 (N_45978,N_44818,N_44971);
or U45979 (N_45979,N_44583,N_44326);
and U45980 (N_45980,N_44027,N_44389);
nand U45981 (N_45981,N_44667,N_44333);
and U45982 (N_45982,N_44372,N_44165);
or U45983 (N_45983,N_44800,N_44885);
nand U45984 (N_45984,N_44427,N_44280);
nand U45985 (N_45985,N_44776,N_44996);
nor U45986 (N_45986,N_44889,N_44788);
xnor U45987 (N_45987,N_44257,N_44497);
xor U45988 (N_45988,N_44236,N_44323);
and U45989 (N_45989,N_44012,N_44126);
nand U45990 (N_45990,N_44873,N_44681);
nand U45991 (N_45991,N_44396,N_44882);
nand U45992 (N_45992,N_44053,N_44424);
and U45993 (N_45993,N_44648,N_44670);
nor U45994 (N_45994,N_44459,N_44978);
nor U45995 (N_45995,N_44294,N_44631);
xor U45996 (N_45996,N_44447,N_44930);
nor U45997 (N_45997,N_44425,N_44851);
xor U45998 (N_45998,N_44896,N_44800);
or U45999 (N_45999,N_44871,N_44499);
and U46000 (N_46000,N_45619,N_45296);
and U46001 (N_46001,N_45160,N_45212);
xnor U46002 (N_46002,N_45912,N_45740);
nand U46003 (N_46003,N_45468,N_45193);
and U46004 (N_46004,N_45030,N_45424);
nor U46005 (N_46005,N_45475,N_45811);
and U46006 (N_46006,N_45666,N_45171);
and U46007 (N_46007,N_45636,N_45023);
and U46008 (N_46008,N_45727,N_45991);
nand U46009 (N_46009,N_45051,N_45122);
and U46010 (N_46010,N_45606,N_45530);
nor U46011 (N_46011,N_45058,N_45478);
nand U46012 (N_46012,N_45040,N_45162);
or U46013 (N_46013,N_45192,N_45954);
nor U46014 (N_46014,N_45346,N_45258);
or U46015 (N_46015,N_45379,N_45820);
nand U46016 (N_46016,N_45118,N_45190);
nand U46017 (N_46017,N_45084,N_45265);
or U46018 (N_46018,N_45573,N_45618);
and U46019 (N_46019,N_45797,N_45067);
or U46020 (N_46020,N_45673,N_45929);
or U46021 (N_46021,N_45589,N_45043);
and U46022 (N_46022,N_45514,N_45286);
and U46023 (N_46023,N_45541,N_45235);
or U46024 (N_46024,N_45560,N_45466);
or U46025 (N_46025,N_45056,N_45986);
and U46026 (N_46026,N_45378,N_45388);
and U46027 (N_46027,N_45683,N_45342);
or U46028 (N_46028,N_45768,N_45998);
nand U46029 (N_46029,N_45832,N_45052);
nor U46030 (N_46030,N_45248,N_45882);
nand U46031 (N_46031,N_45874,N_45777);
and U46032 (N_46032,N_45701,N_45967);
nand U46033 (N_46033,N_45690,N_45668);
or U46034 (N_46034,N_45965,N_45376);
and U46035 (N_46035,N_45276,N_45574);
and U46036 (N_46036,N_45593,N_45999);
or U46037 (N_46037,N_45571,N_45840);
xor U46038 (N_46038,N_45729,N_45665);
nand U46039 (N_46039,N_45305,N_45521);
or U46040 (N_46040,N_45760,N_45936);
and U46041 (N_46041,N_45922,N_45973);
xor U46042 (N_46042,N_45269,N_45578);
and U46043 (N_46043,N_45138,N_45303);
nor U46044 (N_46044,N_45713,N_45498);
nor U46045 (N_46045,N_45195,N_45615);
nor U46046 (N_46046,N_45037,N_45282);
nor U46047 (N_46047,N_45370,N_45399);
xnor U46048 (N_46048,N_45351,N_45858);
xor U46049 (N_46049,N_45057,N_45823);
and U46050 (N_46050,N_45497,N_45904);
nor U46051 (N_46051,N_45396,N_45487);
nor U46052 (N_46052,N_45557,N_45054);
nor U46053 (N_46053,N_45790,N_45073);
or U46054 (N_46054,N_45640,N_45100);
and U46055 (N_46055,N_45253,N_45460);
nor U46056 (N_46056,N_45712,N_45580);
and U46057 (N_46057,N_45196,N_45005);
or U46058 (N_46058,N_45504,N_45720);
xor U46059 (N_46059,N_45816,N_45564);
nand U46060 (N_46060,N_45069,N_45523);
nor U46061 (N_46061,N_45128,N_45168);
nand U46062 (N_46062,N_45637,N_45358);
or U46063 (N_46063,N_45219,N_45545);
nand U46064 (N_46064,N_45135,N_45208);
and U46065 (N_46065,N_45825,N_45472);
nor U46066 (N_46066,N_45060,N_45794);
xnor U46067 (N_46067,N_45739,N_45170);
and U46068 (N_46068,N_45588,N_45716);
or U46069 (N_46069,N_45203,N_45380);
nand U46070 (N_46070,N_45134,N_45698);
nand U46071 (N_46071,N_45315,N_45048);
and U46072 (N_46072,N_45322,N_45743);
or U46073 (N_46073,N_45941,N_45481);
nand U46074 (N_46074,N_45446,N_45031);
nor U46075 (N_46075,N_45624,N_45479);
nand U46076 (N_46076,N_45584,N_45008);
xor U46077 (N_46077,N_45197,N_45995);
nand U46078 (N_46078,N_45719,N_45651);
or U46079 (N_46079,N_45232,N_45937);
nand U46080 (N_46080,N_45951,N_45393);
or U46081 (N_46081,N_45340,N_45722);
nand U46082 (N_46082,N_45707,N_45136);
or U46083 (N_46083,N_45792,N_45293);
and U46084 (N_46084,N_45141,N_45220);
nor U46085 (N_46085,N_45458,N_45164);
xor U46086 (N_46086,N_45471,N_45394);
or U46087 (N_46087,N_45610,N_45486);
nor U46088 (N_46088,N_45109,N_45205);
xor U46089 (N_46089,N_45670,N_45997);
or U46090 (N_46090,N_45550,N_45125);
nand U46091 (N_46091,N_45959,N_45845);
or U46092 (N_46092,N_45107,N_45279);
or U46093 (N_46093,N_45178,N_45254);
and U46094 (N_46094,N_45108,N_45085);
or U46095 (N_46095,N_45605,N_45184);
nand U46096 (N_46096,N_45968,N_45587);
nand U46097 (N_46097,N_45207,N_45749);
nand U46098 (N_46098,N_45309,N_45464);
or U46099 (N_46099,N_45508,N_45601);
nand U46100 (N_46100,N_45076,N_45176);
xnor U46101 (N_46101,N_45417,N_45274);
and U46102 (N_46102,N_45061,N_45510);
and U46103 (N_46103,N_45694,N_45019);
or U46104 (N_46104,N_45103,N_45744);
xnor U46105 (N_46105,N_45449,N_45524);
nand U46106 (N_46106,N_45570,N_45635);
or U46107 (N_46107,N_45865,N_45110);
xnor U46108 (N_46108,N_45401,N_45021);
nor U46109 (N_46109,N_45405,N_45717);
and U46110 (N_46110,N_45554,N_45714);
and U46111 (N_46111,N_45301,N_45256);
nand U46112 (N_46112,N_45117,N_45325);
or U46113 (N_46113,N_45803,N_45266);
nand U46114 (N_46114,N_45526,N_45402);
nor U46115 (N_46115,N_45724,N_45907);
and U46116 (N_46116,N_45983,N_45503);
and U46117 (N_46117,N_45243,N_45596);
xnor U46118 (N_46118,N_45038,N_45230);
or U46119 (N_46119,N_45201,N_45369);
xor U46120 (N_46120,N_45600,N_45906);
nand U46121 (N_46121,N_45864,N_45373);
nor U46122 (N_46122,N_45834,N_45774);
and U46123 (N_46123,N_45897,N_45147);
and U46124 (N_46124,N_45577,N_45533);
nor U46125 (N_46125,N_45347,N_45330);
and U46126 (N_46126,N_45980,N_45518);
nand U46127 (N_46127,N_45808,N_45126);
or U46128 (N_46128,N_45028,N_45231);
nand U46129 (N_46129,N_45708,N_45689);
nand U46130 (N_46130,N_45535,N_45101);
nor U46131 (N_46131,N_45154,N_45785);
nor U46132 (N_46132,N_45529,N_45960);
nor U46133 (N_46133,N_45151,N_45211);
nand U46134 (N_46134,N_45075,N_45338);
xnor U46135 (N_46135,N_45260,N_45320);
or U46136 (N_46136,N_45591,N_45956);
and U46137 (N_46137,N_45415,N_45661);
xnor U46138 (N_46138,N_45461,N_45306);
nor U46139 (N_46139,N_45447,N_45224);
xor U46140 (N_46140,N_45699,N_45324);
or U46141 (N_46141,N_45507,N_45344);
nand U46142 (N_46142,N_45940,N_45970);
nand U46143 (N_46143,N_45971,N_45121);
xor U46144 (N_46144,N_45767,N_45115);
or U46145 (N_46145,N_45066,N_45642);
xor U46146 (N_46146,N_45942,N_45801);
xnor U46147 (N_46147,N_45660,N_45490);
nand U46148 (N_46148,N_45569,N_45307);
and U46149 (N_46149,N_45050,N_45511);
nor U46150 (N_46150,N_45543,N_45658);
xnor U46151 (N_46151,N_45400,N_45945);
or U46152 (N_46152,N_45444,N_45844);
nand U46153 (N_46153,N_45992,N_45285);
xor U46154 (N_46154,N_45068,N_45887);
and U46155 (N_46155,N_45289,N_45988);
or U46156 (N_46156,N_45482,N_45742);
nor U46157 (N_46157,N_45657,N_45901);
xor U46158 (N_46158,N_45181,N_45806);
and U46159 (N_46159,N_45617,N_45867);
nor U46160 (N_46160,N_45982,N_45830);
and U46161 (N_46161,N_45757,N_45928);
or U46162 (N_46162,N_45693,N_45140);
xnor U46163 (N_46163,N_45563,N_45562);
and U46164 (N_46164,N_45902,N_45985);
nand U46165 (N_46165,N_45963,N_45202);
nor U46166 (N_46166,N_45159,N_45723);
xnor U46167 (N_46167,N_45528,N_45662);
xnor U46168 (N_46168,N_45218,N_45080);
nand U46169 (N_46169,N_45969,N_45442);
nand U46170 (N_46170,N_45851,N_45221);
nand U46171 (N_46171,N_45782,N_45431);
or U46172 (N_46172,N_45352,N_45798);
xor U46173 (N_46173,N_45656,N_45416);
and U46174 (N_46174,N_45020,N_45924);
and U46175 (N_46175,N_45977,N_45311);
nor U46176 (N_46176,N_45775,N_45946);
nor U46177 (N_46177,N_45515,N_45145);
or U46178 (N_46178,N_45372,N_45927);
nand U46179 (N_46179,N_45161,N_45480);
or U46180 (N_46180,N_45731,N_45228);
xnor U46181 (N_46181,N_45632,N_45227);
or U46182 (N_46182,N_45104,N_45718);
xnor U46183 (N_46183,N_45055,N_45634);
and U46184 (N_46184,N_45966,N_45007);
or U46185 (N_46185,N_45185,N_45839);
or U46186 (N_46186,N_45249,N_45456);
or U46187 (N_46187,N_45488,N_45500);
nand U46188 (N_46188,N_45931,N_45900);
xnor U46189 (N_46189,N_45548,N_45106);
nor U46190 (N_46190,N_45214,N_45863);
nor U46191 (N_46191,N_45403,N_45264);
nand U46192 (N_46192,N_45827,N_45169);
or U46193 (N_46193,N_45413,N_45143);
nand U46194 (N_46194,N_45703,N_45200);
xnor U46195 (N_46195,N_45215,N_45063);
nor U46196 (N_46196,N_45331,N_45327);
xnor U46197 (N_46197,N_45566,N_45793);
nand U46198 (N_46198,N_45654,N_45861);
nor U46199 (N_46199,N_45333,N_45981);
nor U46200 (N_46200,N_45011,N_45278);
nor U46201 (N_46201,N_45631,N_45319);
or U46202 (N_46202,N_45871,N_45706);
and U46203 (N_46203,N_45321,N_45217);
and U46204 (N_46204,N_45824,N_45462);
xor U46205 (N_46205,N_45738,N_45923);
xnor U46206 (N_46206,N_45873,N_45835);
xor U46207 (N_46207,N_45741,N_45586);
nand U46208 (N_46208,N_45990,N_45065);
or U46209 (N_46209,N_45492,N_45819);
nor U46210 (N_46210,N_45152,N_45407);
and U46211 (N_46211,N_45086,N_45594);
nor U46212 (N_46212,N_45229,N_45158);
and U46213 (N_46213,N_45129,N_45189);
and U46214 (N_46214,N_45764,N_45565);
nand U46215 (N_46215,N_45263,N_45209);
or U46216 (N_46216,N_45418,N_45916);
or U46217 (N_46217,N_45697,N_45355);
and U46218 (N_46218,N_45626,N_45172);
nand U46219 (N_46219,N_45976,N_45261);
nor U46220 (N_46220,N_45167,N_45093);
or U46221 (N_46221,N_45889,N_45377);
xnor U46222 (N_46222,N_45572,N_45705);
and U46223 (N_46223,N_45025,N_45896);
and U46224 (N_46224,N_45341,N_45875);
xor U46225 (N_46225,N_45427,N_45750);
and U46226 (N_46226,N_45675,N_45520);
nor U46227 (N_46227,N_45421,N_45292);
nor U46228 (N_46228,N_45318,N_45892);
or U46229 (N_46229,N_45733,N_45879);
or U46230 (N_46230,N_45602,N_45919);
nand U46231 (N_46231,N_45495,N_45911);
and U46232 (N_46232,N_45206,N_45317);
nor U46233 (N_46233,N_45244,N_45392);
xnor U46234 (N_46234,N_45555,N_45072);
or U46235 (N_46235,N_45818,N_45046);
xnor U46236 (N_46236,N_45860,N_45805);
nand U46237 (N_46237,N_45575,N_45312);
and U46238 (N_46238,N_45842,N_45348);
nor U46239 (N_46239,N_45888,N_45337);
or U46240 (N_46240,N_45387,N_45288);
nand U46241 (N_46241,N_45002,N_45608);
xnor U46242 (N_46242,N_45807,N_45033);
nand U46243 (N_46243,N_45385,N_45964);
nor U46244 (N_46244,N_45519,N_45450);
or U46245 (N_46245,N_45778,N_45756);
xor U46246 (N_46246,N_45237,N_45763);
or U46247 (N_46247,N_45383,N_45137);
or U46248 (N_46248,N_45938,N_45150);
or U46249 (N_46249,N_45979,N_45246);
nand U46250 (N_46250,N_45509,N_45696);
xor U46251 (N_46251,N_45680,N_45843);
nand U46252 (N_46252,N_45796,N_45664);
xnor U46253 (N_46253,N_45975,N_45921);
nand U46254 (N_46254,N_45006,N_45531);
and U46255 (N_46255,N_45083,N_45188);
or U46256 (N_46256,N_45667,N_45925);
or U46257 (N_46257,N_45438,N_45210);
xor U46258 (N_46258,N_45485,N_45859);
and U46259 (N_46259,N_45334,N_45003);
xor U46260 (N_46260,N_45962,N_45009);
or U46261 (N_46261,N_45476,N_45627);
nand U46262 (N_46262,N_45895,N_45585);
and U46263 (N_46263,N_45730,N_45786);
nor U46264 (N_46264,N_45079,N_45684);
or U46265 (N_46265,N_45166,N_45240);
nor U46266 (N_46266,N_45360,N_45926);
nor U46267 (N_46267,N_45721,N_45391);
nand U46268 (N_46268,N_45802,N_45645);
or U46269 (N_46269,N_45609,N_45633);
and U46270 (N_46270,N_45153,N_45119);
and U46271 (N_46271,N_45641,N_45536);
nor U46272 (N_46272,N_45898,N_45769);
nand U46273 (N_46273,N_45583,N_45247);
nor U46274 (N_46274,N_45855,N_45746);
xnor U46275 (N_46275,N_45682,N_45692);
and U46276 (N_46276,N_45643,N_45809);
nand U46277 (N_46277,N_45182,N_45275);
or U46278 (N_46278,N_45148,N_45653);
nor U46279 (N_46279,N_45499,N_45457);
or U46280 (N_46280,N_45089,N_45629);
and U46281 (N_46281,N_45647,N_45287);
nand U46282 (N_46282,N_45259,N_45071);
and U46283 (N_46283,N_45493,N_45551);
or U46284 (N_46284,N_45512,N_45903);
nor U46285 (N_46285,N_45174,N_45886);
nor U46286 (N_46286,N_45544,N_45542);
nor U46287 (N_46287,N_45622,N_45078);
or U46288 (N_46288,N_45027,N_45198);
nor U46289 (N_46289,N_45828,N_45821);
and U46290 (N_46290,N_45612,N_45869);
xnor U46291 (N_46291,N_45426,N_45893);
nor U46292 (N_46292,N_45621,N_45398);
xor U46293 (N_46293,N_45862,N_45491);
xnor U46294 (N_46294,N_45677,N_45425);
or U46295 (N_46295,N_45681,N_45817);
or U46296 (N_46296,N_45905,N_45179);
xnor U46297 (N_46297,N_45866,N_45620);
nor U46298 (N_46298,N_45894,N_45779);
xor U46299 (N_46299,N_45868,N_45336);
nand U46300 (N_46300,N_45726,N_45099);
nand U46301 (N_46301,N_45017,N_45024);
or U46302 (N_46302,N_45582,N_45384);
xnor U46303 (N_46303,N_45463,N_45077);
nand U46304 (N_46304,N_45111,N_45517);
and U46305 (N_46305,N_45113,N_45395);
and U46306 (N_46306,N_45271,N_45829);
nand U46307 (N_46307,N_45298,N_45381);
nand U46308 (N_46308,N_45592,N_45004);
xor U46309 (N_46309,N_45097,N_45857);
or U46310 (N_46310,N_45314,N_45837);
and U46311 (N_46311,N_45909,N_45302);
nor U46312 (N_46312,N_45300,N_45870);
and U46313 (N_46313,N_45590,N_45496);
xnor U46314 (N_46314,N_45725,N_45532);
xnor U46315 (N_46315,N_45236,N_45933);
nor U46316 (N_46316,N_45546,N_45241);
nor U46317 (N_46317,N_45112,N_45155);
xnor U46318 (N_46318,N_45053,N_45935);
xor U46319 (N_46319,N_45081,N_45669);
nor U46320 (N_46320,N_45049,N_45538);
and U46321 (N_46321,N_45273,N_45652);
or U46322 (N_46322,N_45294,N_45978);
nor U46323 (N_46323,N_45428,N_45146);
or U46324 (N_46324,N_45091,N_45087);
or U46325 (N_46325,N_45678,N_45368);
or U46326 (N_46326,N_45761,N_45556);
nand U46327 (N_46327,N_45194,N_45993);
or U46328 (N_46328,N_45445,N_45382);
and U46329 (N_46329,N_45124,N_45412);
nand U46330 (N_46330,N_45386,N_45501);
or U46331 (N_46331,N_45223,N_45453);
nand U46332 (N_46332,N_45568,N_45949);
xor U46333 (N_46333,N_45534,N_45848);
nand U46334 (N_46334,N_45186,N_45687);
xor U46335 (N_46335,N_45751,N_45216);
and U46336 (N_46336,N_45180,N_45173);
and U46337 (N_46337,N_45788,N_45772);
or U46338 (N_46338,N_45452,N_45597);
nor U46339 (N_46339,N_45308,N_45070);
and U46340 (N_46340,N_45120,N_45789);
nor U46341 (N_46341,N_45540,N_45748);
or U46342 (N_46342,N_45525,N_45679);
nor U46343 (N_46343,N_45252,N_45088);
nor U46344 (N_46344,N_45813,N_45953);
nand U46345 (N_46345,N_45233,N_45156);
or U46346 (N_46346,N_45847,N_45822);
xnor U46347 (N_46347,N_45422,N_45074);
nand U46348 (N_46348,N_45947,N_45611);
nor U46349 (N_46349,N_45345,N_45251);
or U46350 (N_46350,N_45225,N_45934);
and U46351 (N_46351,N_45362,N_45350);
and U46352 (N_46352,N_45144,N_45814);
nand U46353 (N_46353,N_45695,N_45715);
nor U46354 (N_46354,N_45709,N_45361);
xnor U46355 (N_46355,N_45434,N_45989);
nand U46356 (N_46356,N_45132,N_45957);
and U46357 (N_46357,N_45354,N_45604);
xnor U46358 (N_46358,N_45773,N_45357);
nand U46359 (N_46359,N_45872,N_45854);
xor U46360 (N_46360,N_45776,N_45436);
xor U46361 (N_46361,N_45810,N_45752);
and U46362 (N_46362,N_45036,N_45000);
or U46363 (N_46363,N_45559,N_45408);
or U46364 (N_46364,N_45467,N_45257);
or U46365 (N_46365,N_45766,N_45952);
nand U46366 (N_46366,N_45853,N_45477);
or U46367 (N_46367,N_45187,N_45014);
nor U46368 (N_46368,N_45239,N_45270);
or U46369 (N_46369,N_45414,N_45026);
or U46370 (N_46370,N_45042,N_45437);
nor U46371 (N_46371,N_45579,N_45943);
nand U46372 (N_46372,N_45625,N_45116);
or U46373 (N_46373,N_45780,N_45672);
or U46374 (N_46374,N_45759,N_45163);
nor U46375 (N_46375,N_45800,N_45238);
nor U46376 (N_46376,N_45096,N_45890);
and U46377 (N_46377,N_45595,N_45771);
nor U46378 (N_46378,N_45671,N_45812);
xor U46379 (N_46379,N_45932,N_45603);
or U46380 (N_46380,N_45638,N_45044);
nand U46381 (N_46381,N_45432,N_45908);
or U46382 (N_46382,N_45753,N_45581);
and U46383 (N_46383,N_45255,N_45440);
nand U46384 (N_46384,N_45527,N_45473);
nor U46385 (N_46385,N_45469,N_45039);
nor U46386 (N_46386,N_45277,N_45349);
nand U46387 (N_46387,N_45397,N_45297);
and U46388 (N_46388,N_45419,N_45326);
or U46389 (N_46389,N_45799,N_45364);
nand U46390 (N_46390,N_45737,N_45429);
nor U46391 (N_46391,N_45663,N_45918);
nand U46392 (N_46392,N_45082,N_45836);
and U46393 (N_46393,N_45765,N_45323);
xnor U46394 (N_46394,N_45213,N_45272);
nor U46395 (N_46395,N_45313,N_45961);
nor U46396 (N_46396,N_45390,N_45423);
nand U46397 (N_46397,N_45262,N_45280);
or U46398 (N_46398,N_45987,N_45114);
and U46399 (N_46399,N_45646,N_45599);
nand U46400 (N_46400,N_45833,N_45770);
xnor U46401 (N_46401,N_45374,N_45018);
xnor U46402 (N_46402,N_45804,N_45245);
and U46403 (N_46403,N_45537,N_45506);
and U46404 (N_46404,N_45328,N_45758);
xnor U46405 (N_46405,N_45704,N_45996);
xor U46406 (N_46406,N_45650,N_45826);
or U46407 (N_46407,N_45371,N_45441);
and U46408 (N_46408,N_45558,N_45686);
nor U46409 (N_46409,N_45489,N_45359);
and U46410 (N_46410,N_45710,N_45948);
or U46411 (N_46411,N_45950,N_45105);
or U46412 (N_46412,N_45702,N_45310);
nor U46413 (N_46413,N_45883,N_45064);
nor U46414 (N_46414,N_45972,N_45142);
and U46415 (N_46415,N_45850,N_45041);
or U46416 (N_46416,N_45013,N_45910);
or U46417 (N_46417,N_45539,N_45877);
or U46418 (N_46418,N_45420,N_45045);
xor U46419 (N_46419,N_45955,N_45881);
nand U46420 (N_46420,N_45149,N_45516);
nand U46421 (N_46421,N_45455,N_45891);
nand U46422 (N_46422,N_45856,N_45204);
nand U46423 (N_46423,N_45483,N_45284);
nor U46424 (N_46424,N_45846,N_45685);
xor U46425 (N_46425,N_45513,N_45831);
xnor U46426 (N_46426,N_45676,N_45130);
xor U46427 (N_46427,N_45165,N_45688);
nor U46428 (N_46428,N_45505,N_45430);
nor U46429 (N_46429,N_45443,N_45914);
and U46430 (N_46430,N_45290,N_45884);
nand U46431 (N_46431,N_45411,N_45994);
and U46432 (N_46432,N_45878,N_45459);
or U46433 (N_46433,N_45127,N_45332);
or U46434 (N_46434,N_45465,N_45090);
xnor U46435 (N_46435,N_45448,N_45494);
xnor U46436 (N_46436,N_45711,N_45920);
or U46437 (N_46437,N_45781,N_45522);
nand U46438 (N_46438,N_45001,N_45630);
xnor U46439 (N_46439,N_45304,N_45291);
nor U46440 (N_46440,N_45183,N_45366);
and U46441 (N_46441,N_45451,N_45316);
nor U46442 (N_46442,N_45029,N_45267);
or U46443 (N_46443,N_45022,N_45648);
xnor U46444 (N_46444,N_45561,N_45102);
and U46445 (N_46445,N_45783,N_45841);
and U46446 (N_46446,N_45639,N_45607);
and U46447 (N_46447,N_45404,N_45092);
nand U46448 (N_46448,N_45123,N_45614);
nand U46449 (N_46449,N_45700,N_45736);
nand U46450 (N_46450,N_45410,N_45032);
or U46451 (N_46451,N_45177,N_45283);
nor U46452 (N_46452,N_45944,N_45062);
xor U46453 (N_46453,N_45885,N_45226);
xor U46454 (N_46454,N_45734,N_45015);
xnor U46455 (N_46455,N_45365,N_45010);
nand U46456 (N_46456,N_45439,N_45917);
nor U46457 (N_46457,N_45474,N_45470);
nand U46458 (N_46458,N_45762,N_45547);
xnor U46459 (N_46459,N_45367,N_45016);
nor U46460 (N_46460,N_45958,N_45375);
nor U46461 (N_46461,N_45502,N_45649);
and U46462 (N_46462,N_45454,N_45974);
nor U46463 (N_46463,N_45849,N_45242);
nor U46464 (N_46464,N_45389,N_45281);
xor U46465 (N_46465,N_45623,N_45250);
xor U46466 (N_46466,N_45655,N_45343);
nor U46467 (N_46467,N_45435,N_45915);
and U46468 (N_46468,N_45175,N_45728);
or U46469 (N_46469,N_45047,N_45930);
xor U46470 (N_46470,N_45133,N_45747);
nor U46471 (N_46471,N_45553,N_45234);
nor U46472 (N_46472,N_45598,N_45406);
nand U46473 (N_46473,N_45335,N_45939);
or U46474 (N_46474,N_45567,N_45484);
nor U46475 (N_46475,N_45059,N_45012);
or U46476 (N_46476,N_45295,N_45222);
nand U46477 (N_46477,N_45409,N_45755);
nand U46478 (N_46478,N_45549,N_45745);
nor U46479 (N_46479,N_45784,N_45576);
xnor U46480 (N_46480,N_45353,N_45795);
xnor U46481 (N_46481,N_45268,N_45098);
nand U46482 (N_46482,N_45984,N_45095);
xor U46483 (N_46483,N_45299,N_45329);
or U46484 (N_46484,N_45613,N_45732);
nand U46485 (N_46485,N_45674,N_45787);
and U46486 (N_46486,N_45094,N_45691);
and U46487 (N_46487,N_45754,N_45876);
xor U46488 (N_46488,N_45735,N_45034);
nand U46489 (N_46489,N_45791,N_45433);
or U46490 (N_46490,N_45191,N_45199);
nand U46491 (N_46491,N_45880,N_45157);
or U46492 (N_46492,N_45644,N_45356);
or U46493 (N_46493,N_45659,N_45139);
nor U46494 (N_46494,N_45131,N_45899);
and U46495 (N_46495,N_45815,N_45913);
xor U46496 (N_46496,N_45339,N_45838);
or U46497 (N_46497,N_45363,N_45852);
and U46498 (N_46498,N_45616,N_45035);
or U46499 (N_46499,N_45552,N_45628);
xor U46500 (N_46500,N_45143,N_45723);
xor U46501 (N_46501,N_45279,N_45396);
nand U46502 (N_46502,N_45427,N_45912);
and U46503 (N_46503,N_45147,N_45255);
nand U46504 (N_46504,N_45420,N_45594);
nor U46505 (N_46505,N_45631,N_45718);
nor U46506 (N_46506,N_45799,N_45851);
xor U46507 (N_46507,N_45400,N_45810);
nand U46508 (N_46508,N_45793,N_45406);
or U46509 (N_46509,N_45213,N_45823);
or U46510 (N_46510,N_45578,N_45063);
nand U46511 (N_46511,N_45433,N_45601);
nand U46512 (N_46512,N_45192,N_45203);
nand U46513 (N_46513,N_45777,N_45794);
or U46514 (N_46514,N_45065,N_45604);
or U46515 (N_46515,N_45180,N_45896);
xnor U46516 (N_46516,N_45383,N_45836);
or U46517 (N_46517,N_45077,N_45453);
and U46518 (N_46518,N_45999,N_45287);
xnor U46519 (N_46519,N_45881,N_45751);
nor U46520 (N_46520,N_45391,N_45650);
nor U46521 (N_46521,N_45978,N_45116);
or U46522 (N_46522,N_45222,N_45547);
nand U46523 (N_46523,N_45777,N_45464);
xor U46524 (N_46524,N_45377,N_45683);
nor U46525 (N_46525,N_45816,N_45721);
nor U46526 (N_46526,N_45824,N_45381);
nor U46527 (N_46527,N_45977,N_45479);
and U46528 (N_46528,N_45845,N_45627);
nand U46529 (N_46529,N_45564,N_45481);
and U46530 (N_46530,N_45343,N_45018);
nand U46531 (N_46531,N_45872,N_45477);
xor U46532 (N_46532,N_45070,N_45528);
and U46533 (N_46533,N_45443,N_45141);
xor U46534 (N_46534,N_45681,N_45584);
or U46535 (N_46535,N_45376,N_45209);
or U46536 (N_46536,N_45430,N_45777);
and U46537 (N_46537,N_45673,N_45838);
nor U46538 (N_46538,N_45374,N_45759);
or U46539 (N_46539,N_45509,N_45549);
nand U46540 (N_46540,N_45603,N_45983);
xor U46541 (N_46541,N_45243,N_45401);
nand U46542 (N_46542,N_45830,N_45790);
or U46543 (N_46543,N_45246,N_45815);
nand U46544 (N_46544,N_45402,N_45474);
xnor U46545 (N_46545,N_45912,N_45569);
xnor U46546 (N_46546,N_45993,N_45350);
xor U46547 (N_46547,N_45224,N_45997);
xor U46548 (N_46548,N_45436,N_45734);
or U46549 (N_46549,N_45483,N_45734);
and U46550 (N_46550,N_45376,N_45596);
and U46551 (N_46551,N_45088,N_45648);
and U46552 (N_46552,N_45645,N_45119);
xnor U46553 (N_46553,N_45059,N_45486);
or U46554 (N_46554,N_45651,N_45659);
nor U46555 (N_46555,N_45040,N_45388);
nor U46556 (N_46556,N_45482,N_45145);
nand U46557 (N_46557,N_45937,N_45471);
nor U46558 (N_46558,N_45194,N_45761);
and U46559 (N_46559,N_45781,N_45950);
xor U46560 (N_46560,N_45695,N_45940);
or U46561 (N_46561,N_45045,N_45150);
or U46562 (N_46562,N_45375,N_45767);
or U46563 (N_46563,N_45115,N_45726);
nor U46564 (N_46564,N_45792,N_45495);
or U46565 (N_46565,N_45337,N_45785);
xnor U46566 (N_46566,N_45299,N_45828);
nand U46567 (N_46567,N_45228,N_45813);
or U46568 (N_46568,N_45742,N_45993);
xor U46569 (N_46569,N_45868,N_45422);
nand U46570 (N_46570,N_45835,N_45294);
xor U46571 (N_46571,N_45248,N_45753);
xor U46572 (N_46572,N_45037,N_45252);
and U46573 (N_46573,N_45256,N_45524);
nand U46574 (N_46574,N_45193,N_45411);
or U46575 (N_46575,N_45761,N_45021);
xnor U46576 (N_46576,N_45817,N_45149);
nand U46577 (N_46577,N_45428,N_45266);
or U46578 (N_46578,N_45969,N_45131);
xor U46579 (N_46579,N_45304,N_45917);
or U46580 (N_46580,N_45807,N_45080);
nand U46581 (N_46581,N_45377,N_45577);
nand U46582 (N_46582,N_45473,N_45418);
xnor U46583 (N_46583,N_45252,N_45755);
nand U46584 (N_46584,N_45230,N_45733);
nand U46585 (N_46585,N_45997,N_45334);
or U46586 (N_46586,N_45971,N_45120);
xnor U46587 (N_46587,N_45634,N_45445);
nor U46588 (N_46588,N_45254,N_45951);
nor U46589 (N_46589,N_45789,N_45716);
xnor U46590 (N_46590,N_45259,N_45574);
nor U46591 (N_46591,N_45434,N_45216);
and U46592 (N_46592,N_45050,N_45531);
and U46593 (N_46593,N_45308,N_45772);
xor U46594 (N_46594,N_45705,N_45535);
nand U46595 (N_46595,N_45482,N_45286);
nand U46596 (N_46596,N_45405,N_45851);
nor U46597 (N_46597,N_45754,N_45270);
and U46598 (N_46598,N_45722,N_45472);
xnor U46599 (N_46599,N_45171,N_45419);
xor U46600 (N_46600,N_45310,N_45939);
xor U46601 (N_46601,N_45255,N_45525);
or U46602 (N_46602,N_45760,N_45437);
and U46603 (N_46603,N_45064,N_45190);
and U46604 (N_46604,N_45012,N_45950);
or U46605 (N_46605,N_45116,N_45310);
nand U46606 (N_46606,N_45025,N_45547);
or U46607 (N_46607,N_45798,N_45334);
xnor U46608 (N_46608,N_45116,N_45364);
and U46609 (N_46609,N_45658,N_45749);
and U46610 (N_46610,N_45741,N_45861);
or U46611 (N_46611,N_45772,N_45955);
or U46612 (N_46612,N_45382,N_45704);
xor U46613 (N_46613,N_45018,N_45669);
nand U46614 (N_46614,N_45590,N_45033);
and U46615 (N_46615,N_45017,N_45306);
xor U46616 (N_46616,N_45711,N_45571);
nor U46617 (N_46617,N_45910,N_45006);
xor U46618 (N_46618,N_45354,N_45881);
or U46619 (N_46619,N_45977,N_45606);
nand U46620 (N_46620,N_45020,N_45413);
xor U46621 (N_46621,N_45352,N_45902);
xor U46622 (N_46622,N_45273,N_45799);
nand U46623 (N_46623,N_45540,N_45617);
or U46624 (N_46624,N_45870,N_45325);
or U46625 (N_46625,N_45864,N_45746);
nor U46626 (N_46626,N_45504,N_45546);
xnor U46627 (N_46627,N_45347,N_45288);
xor U46628 (N_46628,N_45722,N_45178);
and U46629 (N_46629,N_45594,N_45020);
or U46630 (N_46630,N_45727,N_45939);
nand U46631 (N_46631,N_45964,N_45729);
or U46632 (N_46632,N_45010,N_45765);
or U46633 (N_46633,N_45981,N_45797);
nor U46634 (N_46634,N_45317,N_45791);
nand U46635 (N_46635,N_45543,N_45665);
nor U46636 (N_46636,N_45436,N_45937);
nand U46637 (N_46637,N_45227,N_45119);
and U46638 (N_46638,N_45924,N_45917);
and U46639 (N_46639,N_45771,N_45677);
and U46640 (N_46640,N_45254,N_45329);
and U46641 (N_46641,N_45640,N_45656);
xnor U46642 (N_46642,N_45469,N_45320);
nor U46643 (N_46643,N_45470,N_45031);
nor U46644 (N_46644,N_45465,N_45114);
or U46645 (N_46645,N_45965,N_45997);
nand U46646 (N_46646,N_45527,N_45779);
nand U46647 (N_46647,N_45159,N_45807);
and U46648 (N_46648,N_45685,N_45419);
and U46649 (N_46649,N_45748,N_45403);
xor U46650 (N_46650,N_45519,N_45168);
or U46651 (N_46651,N_45155,N_45168);
and U46652 (N_46652,N_45731,N_45615);
nor U46653 (N_46653,N_45221,N_45344);
xnor U46654 (N_46654,N_45387,N_45310);
nand U46655 (N_46655,N_45782,N_45668);
nand U46656 (N_46656,N_45832,N_45649);
or U46657 (N_46657,N_45698,N_45979);
and U46658 (N_46658,N_45506,N_45647);
and U46659 (N_46659,N_45748,N_45926);
xnor U46660 (N_46660,N_45465,N_45444);
nor U46661 (N_46661,N_45810,N_45483);
nand U46662 (N_46662,N_45726,N_45772);
or U46663 (N_46663,N_45377,N_45469);
or U46664 (N_46664,N_45489,N_45874);
and U46665 (N_46665,N_45006,N_45876);
and U46666 (N_46666,N_45418,N_45336);
or U46667 (N_46667,N_45609,N_45946);
and U46668 (N_46668,N_45747,N_45997);
or U46669 (N_46669,N_45956,N_45370);
and U46670 (N_46670,N_45494,N_45774);
nor U46671 (N_46671,N_45953,N_45418);
or U46672 (N_46672,N_45209,N_45222);
nor U46673 (N_46673,N_45894,N_45997);
and U46674 (N_46674,N_45084,N_45438);
xor U46675 (N_46675,N_45346,N_45498);
nor U46676 (N_46676,N_45655,N_45819);
nand U46677 (N_46677,N_45603,N_45449);
or U46678 (N_46678,N_45160,N_45383);
and U46679 (N_46679,N_45450,N_45632);
xor U46680 (N_46680,N_45702,N_45601);
and U46681 (N_46681,N_45126,N_45422);
and U46682 (N_46682,N_45017,N_45112);
or U46683 (N_46683,N_45508,N_45265);
nor U46684 (N_46684,N_45561,N_45341);
nand U46685 (N_46685,N_45382,N_45338);
nor U46686 (N_46686,N_45281,N_45357);
xor U46687 (N_46687,N_45111,N_45653);
and U46688 (N_46688,N_45001,N_45775);
or U46689 (N_46689,N_45533,N_45807);
nand U46690 (N_46690,N_45598,N_45992);
and U46691 (N_46691,N_45852,N_45539);
and U46692 (N_46692,N_45010,N_45410);
and U46693 (N_46693,N_45398,N_45719);
xor U46694 (N_46694,N_45488,N_45855);
nand U46695 (N_46695,N_45402,N_45756);
nor U46696 (N_46696,N_45857,N_45008);
or U46697 (N_46697,N_45573,N_45690);
and U46698 (N_46698,N_45747,N_45696);
nand U46699 (N_46699,N_45259,N_45867);
nor U46700 (N_46700,N_45575,N_45492);
nand U46701 (N_46701,N_45145,N_45302);
or U46702 (N_46702,N_45471,N_45795);
xor U46703 (N_46703,N_45906,N_45280);
and U46704 (N_46704,N_45125,N_45592);
and U46705 (N_46705,N_45018,N_45698);
or U46706 (N_46706,N_45932,N_45709);
xnor U46707 (N_46707,N_45136,N_45339);
or U46708 (N_46708,N_45718,N_45603);
and U46709 (N_46709,N_45115,N_45260);
xor U46710 (N_46710,N_45279,N_45015);
nand U46711 (N_46711,N_45940,N_45233);
nand U46712 (N_46712,N_45233,N_45505);
and U46713 (N_46713,N_45128,N_45964);
xnor U46714 (N_46714,N_45850,N_45061);
xor U46715 (N_46715,N_45825,N_45471);
or U46716 (N_46716,N_45627,N_45262);
and U46717 (N_46717,N_45072,N_45998);
nor U46718 (N_46718,N_45249,N_45192);
nand U46719 (N_46719,N_45025,N_45358);
and U46720 (N_46720,N_45119,N_45097);
nor U46721 (N_46721,N_45818,N_45358);
nand U46722 (N_46722,N_45897,N_45892);
and U46723 (N_46723,N_45356,N_45007);
or U46724 (N_46724,N_45991,N_45041);
nand U46725 (N_46725,N_45392,N_45130);
and U46726 (N_46726,N_45445,N_45101);
nor U46727 (N_46727,N_45162,N_45502);
nor U46728 (N_46728,N_45112,N_45277);
and U46729 (N_46729,N_45631,N_45503);
and U46730 (N_46730,N_45640,N_45723);
nor U46731 (N_46731,N_45079,N_45784);
and U46732 (N_46732,N_45674,N_45948);
or U46733 (N_46733,N_45151,N_45758);
xor U46734 (N_46734,N_45831,N_45492);
xor U46735 (N_46735,N_45649,N_45161);
or U46736 (N_46736,N_45805,N_45496);
nor U46737 (N_46737,N_45741,N_45494);
and U46738 (N_46738,N_45652,N_45255);
and U46739 (N_46739,N_45231,N_45001);
nor U46740 (N_46740,N_45425,N_45705);
or U46741 (N_46741,N_45937,N_45423);
and U46742 (N_46742,N_45699,N_45950);
and U46743 (N_46743,N_45044,N_45614);
or U46744 (N_46744,N_45490,N_45201);
nor U46745 (N_46745,N_45569,N_45930);
or U46746 (N_46746,N_45219,N_45817);
nand U46747 (N_46747,N_45155,N_45820);
and U46748 (N_46748,N_45042,N_45568);
nand U46749 (N_46749,N_45603,N_45172);
nand U46750 (N_46750,N_45183,N_45884);
or U46751 (N_46751,N_45907,N_45948);
or U46752 (N_46752,N_45668,N_45620);
or U46753 (N_46753,N_45862,N_45231);
and U46754 (N_46754,N_45584,N_45600);
and U46755 (N_46755,N_45754,N_45981);
xnor U46756 (N_46756,N_45026,N_45872);
nand U46757 (N_46757,N_45643,N_45123);
xor U46758 (N_46758,N_45841,N_45728);
nor U46759 (N_46759,N_45186,N_45989);
nand U46760 (N_46760,N_45234,N_45437);
xnor U46761 (N_46761,N_45154,N_45449);
xnor U46762 (N_46762,N_45447,N_45401);
nor U46763 (N_46763,N_45482,N_45299);
nor U46764 (N_46764,N_45411,N_45983);
nor U46765 (N_46765,N_45743,N_45883);
nand U46766 (N_46766,N_45606,N_45451);
nor U46767 (N_46767,N_45889,N_45081);
nand U46768 (N_46768,N_45368,N_45967);
nor U46769 (N_46769,N_45915,N_45793);
nand U46770 (N_46770,N_45030,N_45757);
nor U46771 (N_46771,N_45065,N_45862);
nand U46772 (N_46772,N_45693,N_45238);
or U46773 (N_46773,N_45739,N_45059);
or U46774 (N_46774,N_45273,N_45727);
xnor U46775 (N_46775,N_45343,N_45708);
nor U46776 (N_46776,N_45967,N_45791);
xnor U46777 (N_46777,N_45675,N_45034);
and U46778 (N_46778,N_45258,N_45544);
xnor U46779 (N_46779,N_45690,N_45466);
xor U46780 (N_46780,N_45314,N_45529);
nand U46781 (N_46781,N_45861,N_45473);
or U46782 (N_46782,N_45467,N_45363);
or U46783 (N_46783,N_45511,N_45352);
or U46784 (N_46784,N_45360,N_45049);
and U46785 (N_46785,N_45048,N_45112);
nand U46786 (N_46786,N_45494,N_45046);
nand U46787 (N_46787,N_45990,N_45514);
and U46788 (N_46788,N_45952,N_45263);
or U46789 (N_46789,N_45940,N_45254);
or U46790 (N_46790,N_45596,N_45603);
nand U46791 (N_46791,N_45149,N_45594);
and U46792 (N_46792,N_45997,N_45451);
nand U46793 (N_46793,N_45079,N_45387);
nand U46794 (N_46794,N_45426,N_45843);
xnor U46795 (N_46795,N_45215,N_45392);
nor U46796 (N_46796,N_45211,N_45941);
xnor U46797 (N_46797,N_45157,N_45184);
nor U46798 (N_46798,N_45311,N_45501);
or U46799 (N_46799,N_45432,N_45485);
or U46800 (N_46800,N_45822,N_45620);
or U46801 (N_46801,N_45897,N_45960);
and U46802 (N_46802,N_45704,N_45760);
nor U46803 (N_46803,N_45222,N_45142);
or U46804 (N_46804,N_45843,N_45313);
xor U46805 (N_46805,N_45961,N_45822);
or U46806 (N_46806,N_45733,N_45658);
and U46807 (N_46807,N_45075,N_45950);
nor U46808 (N_46808,N_45062,N_45750);
nand U46809 (N_46809,N_45489,N_45484);
nor U46810 (N_46810,N_45395,N_45327);
or U46811 (N_46811,N_45830,N_45138);
nor U46812 (N_46812,N_45516,N_45131);
or U46813 (N_46813,N_45082,N_45319);
xor U46814 (N_46814,N_45827,N_45754);
and U46815 (N_46815,N_45332,N_45348);
or U46816 (N_46816,N_45816,N_45024);
nand U46817 (N_46817,N_45358,N_45787);
or U46818 (N_46818,N_45137,N_45142);
and U46819 (N_46819,N_45480,N_45060);
and U46820 (N_46820,N_45093,N_45117);
xor U46821 (N_46821,N_45304,N_45575);
nor U46822 (N_46822,N_45538,N_45249);
or U46823 (N_46823,N_45648,N_45819);
xor U46824 (N_46824,N_45054,N_45363);
nand U46825 (N_46825,N_45801,N_45881);
nor U46826 (N_46826,N_45102,N_45729);
nand U46827 (N_46827,N_45558,N_45409);
nand U46828 (N_46828,N_45864,N_45673);
xor U46829 (N_46829,N_45945,N_45647);
and U46830 (N_46830,N_45827,N_45220);
xnor U46831 (N_46831,N_45298,N_45299);
xnor U46832 (N_46832,N_45288,N_45683);
and U46833 (N_46833,N_45270,N_45646);
and U46834 (N_46834,N_45407,N_45260);
nor U46835 (N_46835,N_45796,N_45498);
or U46836 (N_46836,N_45829,N_45530);
nand U46837 (N_46837,N_45385,N_45947);
nor U46838 (N_46838,N_45975,N_45762);
xnor U46839 (N_46839,N_45627,N_45393);
or U46840 (N_46840,N_45603,N_45602);
xnor U46841 (N_46841,N_45662,N_45742);
nor U46842 (N_46842,N_45116,N_45536);
or U46843 (N_46843,N_45720,N_45003);
nor U46844 (N_46844,N_45587,N_45189);
xor U46845 (N_46845,N_45892,N_45495);
nand U46846 (N_46846,N_45607,N_45979);
and U46847 (N_46847,N_45241,N_45240);
and U46848 (N_46848,N_45624,N_45923);
nand U46849 (N_46849,N_45346,N_45971);
and U46850 (N_46850,N_45354,N_45519);
nor U46851 (N_46851,N_45147,N_45037);
and U46852 (N_46852,N_45551,N_45514);
nand U46853 (N_46853,N_45763,N_45920);
and U46854 (N_46854,N_45639,N_45633);
nand U46855 (N_46855,N_45947,N_45136);
nor U46856 (N_46856,N_45843,N_45350);
nor U46857 (N_46857,N_45874,N_45467);
xor U46858 (N_46858,N_45516,N_45388);
nor U46859 (N_46859,N_45326,N_45630);
nor U46860 (N_46860,N_45126,N_45161);
nor U46861 (N_46861,N_45257,N_45490);
xnor U46862 (N_46862,N_45905,N_45434);
and U46863 (N_46863,N_45476,N_45999);
nor U46864 (N_46864,N_45139,N_45176);
and U46865 (N_46865,N_45149,N_45592);
xor U46866 (N_46866,N_45282,N_45967);
xor U46867 (N_46867,N_45826,N_45130);
and U46868 (N_46868,N_45910,N_45188);
nor U46869 (N_46869,N_45691,N_45650);
or U46870 (N_46870,N_45094,N_45328);
nand U46871 (N_46871,N_45488,N_45139);
nand U46872 (N_46872,N_45267,N_45975);
nor U46873 (N_46873,N_45011,N_45417);
or U46874 (N_46874,N_45888,N_45729);
xor U46875 (N_46875,N_45196,N_45323);
xor U46876 (N_46876,N_45038,N_45628);
nor U46877 (N_46877,N_45641,N_45407);
and U46878 (N_46878,N_45626,N_45394);
xor U46879 (N_46879,N_45959,N_45886);
nor U46880 (N_46880,N_45205,N_45879);
nand U46881 (N_46881,N_45887,N_45049);
xor U46882 (N_46882,N_45315,N_45160);
and U46883 (N_46883,N_45820,N_45228);
nor U46884 (N_46884,N_45573,N_45915);
and U46885 (N_46885,N_45272,N_45199);
xor U46886 (N_46886,N_45121,N_45410);
and U46887 (N_46887,N_45037,N_45755);
and U46888 (N_46888,N_45495,N_45683);
nand U46889 (N_46889,N_45216,N_45457);
and U46890 (N_46890,N_45323,N_45758);
and U46891 (N_46891,N_45248,N_45588);
and U46892 (N_46892,N_45535,N_45542);
xnor U46893 (N_46893,N_45304,N_45615);
nand U46894 (N_46894,N_45585,N_45929);
and U46895 (N_46895,N_45830,N_45760);
xnor U46896 (N_46896,N_45994,N_45503);
and U46897 (N_46897,N_45487,N_45140);
nand U46898 (N_46898,N_45977,N_45351);
nor U46899 (N_46899,N_45228,N_45257);
nor U46900 (N_46900,N_45965,N_45767);
or U46901 (N_46901,N_45177,N_45581);
xnor U46902 (N_46902,N_45472,N_45333);
or U46903 (N_46903,N_45807,N_45256);
and U46904 (N_46904,N_45243,N_45199);
nand U46905 (N_46905,N_45137,N_45244);
or U46906 (N_46906,N_45245,N_45401);
nor U46907 (N_46907,N_45204,N_45828);
nand U46908 (N_46908,N_45958,N_45641);
and U46909 (N_46909,N_45632,N_45625);
and U46910 (N_46910,N_45138,N_45597);
nand U46911 (N_46911,N_45254,N_45949);
xor U46912 (N_46912,N_45116,N_45650);
nand U46913 (N_46913,N_45727,N_45594);
xor U46914 (N_46914,N_45742,N_45182);
or U46915 (N_46915,N_45042,N_45255);
xor U46916 (N_46916,N_45756,N_45980);
and U46917 (N_46917,N_45755,N_45138);
and U46918 (N_46918,N_45417,N_45690);
nand U46919 (N_46919,N_45275,N_45141);
nand U46920 (N_46920,N_45799,N_45344);
and U46921 (N_46921,N_45835,N_45154);
and U46922 (N_46922,N_45357,N_45538);
nand U46923 (N_46923,N_45899,N_45451);
xnor U46924 (N_46924,N_45072,N_45000);
xnor U46925 (N_46925,N_45152,N_45276);
nand U46926 (N_46926,N_45423,N_45717);
nand U46927 (N_46927,N_45820,N_45482);
or U46928 (N_46928,N_45198,N_45345);
nor U46929 (N_46929,N_45508,N_45667);
nor U46930 (N_46930,N_45361,N_45972);
xnor U46931 (N_46931,N_45724,N_45875);
xor U46932 (N_46932,N_45386,N_45607);
nand U46933 (N_46933,N_45084,N_45316);
nand U46934 (N_46934,N_45653,N_45412);
nor U46935 (N_46935,N_45479,N_45979);
xor U46936 (N_46936,N_45249,N_45225);
xor U46937 (N_46937,N_45292,N_45236);
and U46938 (N_46938,N_45187,N_45496);
xnor U46939 (N_46939,N_45963,N_45956);
or U46940 (N_46940,N_45341,N_45433);
or U46941 (N_46941,N_45674,N_45973);
nand U46942 (N_46942,N_45178,N_45409);
xor U46943 (N_46943,N_45648,N_45236);
nor U46944 (N_46944,N_45221,N_45004);
nor U46945 (N_46945,N_45019,N_45937);
xor U46946 (N_46946,N_45174,N_45337);
and U46947 (N_46947,N_45309,N_45009);
nand U46948 (N_46948,N_45299,N_45843);
or U46949 (N_46949,N_45539,N_45614);
xor U46950 (N_46950,N_45874,N_45115);
or U46951 (N_46951,N_45423,N_45271);
or U46952 (N_46952,N_45774,N_45083);
and U46953 (N_46953,N_45632,N_45432);
and U46954 (N_46954,N_45105,N_45886);
nand U46955 (N_46955,N_45662,N_45012);
nor U46956 (N_46956,N_45145,N_45035);
nand U46957 (N_46957,N_45605,N_45183);
xnor U46958 (N_46958,N_45186,N_45510);
or U46959 (N_46959,N_45937,N_45739);
nand U46960 (N_46960,N_45925,N_45100);
nand U46961 (N_46961,N_45525,N_45635);
nor U46962 (N_46962,N_45856,N_45462);
nor U46963 (N_46963,N_45243,N_45642);
xnor U46964 (N_46964,N_45836,N_45604);
xor U46965 (N_46965,N_45085,N_45790);
nand U46966 (N_46966,N_45148,N_45923);
nor U46967 (N_46967,N_45808,N_45240);
or U46968 (N_46968,N_45479,N_45530);
nor U46969 (N_46969,N_45038,N_45659);
nand U46970 (N_46970,N_45627,N_45928);
nor U46971 (N_46971,N_45468,N_45148);
and U46972 (N_46972,N_45319,N_45636);
nand U46973 (N_46973,N_45606,N_45085);
or U46974 (N_46974,N_45030,N_45609);
xnor U46975 (N_46975,N_45900,N_45165);
and U46976 (N_46976,N_45652,N_45610);
xor U46977 (N_46977,N_45261,N_45254);
nand U46978 (N_46978,N_45188,N_45106);
nand U46979 (N_46979,N_45486,N_45500);
or U46980 (N_46980,N_45263,N_45521);
xnor U46981 (N_46981,N_45315,N_45000);
or U46982 (N_46982,N_45027,N_45036);
nor U46983 (N_46983,N_45183,N_45075);
and U46984 (N_46984,N_45041,N_45642);
nand U46985 (N_46985,N_45206,N_45396);
or U46986 (N_46986,N_45433,N_45178);
nor U46987 (N_46987,N_45937,N_45744);
or U46988 (N_46988,N_45125,N_45427);
and U46989 (N_46989,N_45691,N_45505);
nand U46990 (N_46990,N_45388,N_45798);
nor U46991 (N_46991,N_45895,N_45357);
and U46992 (N_46992,N_45327,N_45584);
and U46993 (N_46993,N_45202,N_45391);
nor U46994 (N_46994,N_45853,N_45770);
and U46995 (N_46995,N_45768,N_45600);
xnor U46996 (N_46996,N_45038,N_45029);
or U46997 (N_46997,N_45469,N_45772);
nand U46998 (N_46998,N_45136,N_45520);
nand U46999 (N_46999,N_45067,N_45828);
nand U47000 (N_47000,N_46189,N_46088);
and U47001 (N_47001,N_46466,N_46473);
nor U47002 (N_47002,N_46073,N_46153);
and U47003 (N_47003,N_46076,N_46729);
or U47004 (N_47004,N_46870,N_46106);
nor U47005 (N_47005,N_46269,N_46639);
nor U47006 (N_47006,N_46130,N_46908);
nor U47007 (N_47007,N_46480,N_46867);
xnor U47008 (N_47008,N_46333,N_46818);
nand U47009 (N_47009,N_46450,N_46880);
or U47010 (N_47010,N_46795,N_46471);
or U47011 (N_47011,N_46810,N_46652);
nand U47012 (N_47012,N_46525,N_46435);
or U47013 (N_47013,N_46537,N_46503);
or U47014 (N_47014,N_46474,N_46558);
or U47015 (N_47015,N_46118,N_46135);
nor U47016 (N_47016,N_46006,N_46846);
nand U47017 (N_47017,N_46332,N_46402);
or U47018 (N_47018,N_46311,N_46221);
or U47019 (N_47019,N_46266,N_46562);
and U47020 (N_47020,N_46711,N_46233);
or U47021 (N_47021,N_46369,N_46097);
xor U47022 (N_47022,N_46085,N_46938);
nor U47023 (N_47023,N_46581,N_46806);
xor U47024 (N_47024,N_46033,N_46296);
xor U47025 (N_47025,N_46984,N_46678);
or U47026 (N_47026,N_46164,N_46860);
or U47027 (N_47027,N_46023,N_46143);
xor U47028 (N_47028,N_46363,N_46765);
or U47029 (N_47029,N_46357,N_46007);
xnor U47030 (N_47030,N_46655,N_46965);
nor U47031 (N_47031,N_46102,N_46874);
xnor U47032 (N_47032,N_46513,N_46326);
or U47033 (N_47033,N_46848,N_46213);
xnor U47034 (N_47034,N_46578,N_46775);
nand U47035 (N_47035,N_46351,N_46918);
and U47036 (N_47036,N_46434,N_46975);
and U47037 (N_47037,N_46421,N_46585);
nor U47038 (N_47038,N_46543,N_46358);
and U47039 (N_47039,N_46069,N_46350);
or U47040 (N_47040,N_46997,N_46425);
xor U47041 (N_47041,N_46500,N_46361);
nor U47042 (N_47042,N_46445,N_46321);
nor U47043 (N_47043,N_46641,N_46868);
nand U47044 (N_47044,N_46961,N_46178);
nand U47045 (N_47045,N_46013,N_46527);
nand U47046 (N_47046,N_46408,N_46077);
nor U47047 (N_47047,N_46339,N_46574);
xor U47048 (N_47048,N_46442,N_46043);
and U47049 (N_47049,N_46851,N_46891);
xnor U47050 (N_47050,N_46624,N_46760);
or U47051 (N_47051,N_46032,N_46053);
or U47052 (N_47052,N_46991,N_46092);
nor U47053 (N_47053,N_46941,N_46458);
nor U47054 (N_47054,N_46741,N_46451);
nand U47055 (N_47055,N_46298,N_46968);
xnor U47056 (N_47056,N_46909,N_46847);
and U47057 (N_47057,N_46637,N_46012);
and U47058 (N_47058,N_46969,N_46075);
nor U47059 (N_47059,N_46668,N_46418);
or U47060 (N_47060,N_46956,N_46622);
or U47061 (N_47061,N_46716,N_46696);
nand U47062 (N_47062,N_46057,N_46228);
xnor U47063 (N_47063,N_46763,N_46936);
xnor U47064 (N_47064,N_46808,N_46879);
or U47065 (N_47065,N_46823,N_46087);
or U47066 (N_47066,N_46548,N_46258);
nor U47067 (N_47067,N_46319,N_46971);
nand U47068 (N_47068,N_46125,N_46694);
or U47069 (N_47069,N_46252,N_46105);
xor U47070 (N_47070,N_46920,N_46272);
xnor U47071 (N_47071,N_46551,N_46403);
nand U47072 (N_47072,N_46432,N_46833);
nand U47073 (N_47073,N_46573,N_46003);
nor U47074 (N_47074,N_46841,N_46376);
or U47075 (N_47075,N_46204,N_46174);
nand U47076 (N_47076,N_46009,N_46690);
nand U47077 (N_47077,N_46120,N_46507);
or U47078 (N_47078,N_46169,N_46828);
nor U47079 (N_47079,N_46727,N_46519);
nand U47080 (N_47080,N_46188,N_46770);
xor U47081 (N_47081,N_46196,N_46560);
xor U47082 (N_47082,N_46669,N_46029);
xnor U47083 (N_47083,N_46303,N_46406);
or U47084 (N_47084,N_46923,N_46510);
and U47085 (N_47085,N_46697,N_46985);
or U47086 (N_47086,N_46972,N_46888);
and U47087 (N_47087,N_46679,N_46264);
xnor U47088 (N_47088,N_46355,N_46022);
xnor U47089 (N_47089,N_46515,N_46225);
and U47090 (N_47090,N_46448,N_46268);
xor U47091 (N_47091,N_46664,N_46988);
or U47092 (N_47092,N_46773,N_46005);
nand U47093 (N_47093,N_46235,N_46116);
and U47094 (N_47094,N_46890,N_46516);
nor U47095 (N_47095,N_46996,N_46147);
xnor U47096 (N_47096,N_46994,N_46942);
or U47097 (N_47097,N_46020,N_46356);
xor U47098 (N_47098,N_46602,N_46774);
or U47099 (N_47099,N_46460,N_46577);
nand U47100 (N_47100,N_46101,N_46325);
and U47101 (N_47101,N_46865,N_46001);
nor U47102 (N_47102,N_46200,N_46963);
nor U47103 (N_47103,N_46935,N_46504);
xnor U47104 (N_47104,N_46108,N_46417);
nor U47105 (N_47105,N_46839,N_46820);
nor U47106 (N_47106,N_46384,N_46485);
nor U47107 (N_47107,N_46394,N_46202);
or U47108 (N_47108,N_46280,N_46826);
nor U47109 (N_47109,N_46559,N_46615);
or U47110 (N_47110,N_46712,N_46732);
xnor U47111 (N_47111,N_46365,N_46083);
or U47112 (N_47112,N_46522,N_46031);
xnor U47113 (N_47113,N_46216,N_46227);
nand U47114 (N_47114,N_46966,N_46912);
nand U47115 (N_47115,N_46995,N_46541);
nand U47116 (N_47116,N_46486,N_46079);
or U47117 (N_47117,N_46205,N_46084);
or U47118 (N_47118,N_46008,N_46433);
xor U47119 (N_47119,N_46149,N_46575);
xor U47120 (N_47120,N_46190,N_46010);
or U47121 (N_47121,N_46929,N_46334);
and U47122 (N_47122,N_46282,N_46671);
xor U47123 (N_47123,N_46062,N_46858);
or U47124 (N_47124,N_46722,N_46761);
nand U47125 (N_47125,N_46784,N_46107);
and U47126 (N_47126,N_46337,N_46000);
xnor U47127 (N_47127,N_46064,N_46903);
xnor U47128 (N_47128,N_46786,N_46887);
or U47129 (N_47129,N_46387,N_46281);
nand U47130 (N_47130,N_46497,N_46875);
nor U47131 (N_47131,N_46980,N_46374);
xnor U47132 (N_47132,N_46998,N_46398);
nand U47133 (N_47133,N_46462,N_46547);
nor U47134 (N_47134,N_46168,N_46301);
or U47135 (N_47135,N_46951,N_46185);
xor U47136 (N_47136,N_46844,N_46166);
nand U47137 (N_47137,N_46159,N_46857);
or U47138 (N_47138,N_46199,N_46372);
and U47139 (N_47139,N_46048,N_46928);
and U47140 (N_47140,N_46654,N_46663);
or U47141 (N_47141,N_46790,N_46608);
nand U47142 (N_47142,N_46501,N_46699);
and U47143 (N_47143,N_46892,N_46250);
and U47144 (N_47144,N_46530,N_46505);
and U47145 (N_47145,N_46569,N_46489);
xor U47146 (N_47146,N_46067,N_46813);
xnor U47147 (N_47147,N_46491,N_46977);
xor U47148 (N_47148,N_46026,N_46197);
xor U47149 (N_47149,N_46127,N_46142);
or U47150 (N_47150,N_46152,N_46508);
nor U47151 (N_47151,N_46014,N_46348);
or U47152 (N_47152,N_46482,N_46593);
nor U47153 (N_47153,N_46222,N_46499);
nor U47154 (N_47154,N_46068,N_46091);
nor U47155 (N_47155,N_46566,N_46647);
nor U47156 (N_47156,N_46934,N_46628);
nor U47157 (N_47157,N_46124,N_46978);
nor U47158 (N_47158,N_46302,N_46039);
nand U47159 (N_47159,N_46950,N_46836);
xnor U47160 (N_47160,N_46255,N_46646);
and U47161 (N_47161,N_46295,N_46733);
nand U47162 (N_47162,N_46603,N_46554);
nor U47163 (N_47163,N_46044,N_46805);
nand U47164 (N_47164,N_46484,N_46572);
or U47165 (N_47165,N_46958,N_46821);
nor U47166 (N_47166,N_46932,N_46568);
nor U47167 (N_47167,N_46446,N_46247);
or U47168 (N_47168,N_46873,N_46257);
and U47169 (N_47169,N_46894,N_46390);
xnor U47170 (N_47170,N_46481,N_46090);
or U47171 (N_47171,N_46900,N_46714);
or U47172 (N_47172,N_46443,N_46380);
nand U47173 (N_47173,N_46287,N_46842);
and U47174 (N_47174,N_46160,N_46957);
or U47175 (N_47175,N_46322,N_46399);
or U47176 (N_47176,N_46156,N_46122);
nor U47177 (N_47177,N_46276,N_46538);
nand U47178 (N_47178,N_46744,N_46953);
nor U47179 (N_47179,N_46708,N_46521);
nand U47180 (N_47180,N_46134,N_46742);
and U47181 (N_47181,N_46316,N_46586);
and U47182 (N_47182,N_46126,N_46834);
xnor U47183 (N_47183,N_46772,N_46452);
nand U47184 (N_47184,N_46625,N_46277);
and U47185 (N_47185,N_46922,N_46465);
nand U47186 (N_47186,N_46278,N_46373);
nand U47187 (N_47187,N_46518,N_46871);
xnor U47188 (N_47188,N_46587,N_46050);
or U47189 (N_47189,N_46952,N_46240);
nand U47190 (N_47190,N_46198,N_46747);
or U47191 (N_47191,N_46056,N_46035);
xnor U47192 (N_47192,N_46753,N_46927);
nor U47193 (N_47193,N_46036,N_46184);
nor U47194 (N_47194,N_46674,N_46970);
and U47195 (N_47195,N_46219,N_46746);
xor U47196 (N_47196,N_46893,N_46074);
nor U47197 (N_47197,N_46931,N_46439);
and U47198 (N_47198,N_46379,N_46297);
xor U47199 (N_47199,N_46803,N_46370);
and U47200 (N_47200,N_46565,N_46414);
nor U47201 (N_47201,N_46306,N_46511);
nand U47202 (N_47202,N_46274,N_46705);
nor U47203 (N_47203,N_46150,N_46740);
nand U47204 (N_47204,N_46634,N_46488);
nor U47205 (N_47205,N_46317,N_46176);
or U47206 (N_47206,N_46237,N_46905);
xor U47207 (N_47207,N_46165,N_46299);
and U47208 (N_47208,N_46864,N_46644);
or U47209 (N_47209,N_46901,N_46889);
nand U47210 (N_47210,N_46065,N_46094);
or U47211 (N_47211,N_46218,N_46632);
xor U47212 (N_47212,N_46183,N_46990);
or U47213 (N_47213,N_46144,N_46393);
xor U47214 (N_47214,N_46241,N_46463);
nor U47215 (N_47215,N_46114,N_46328);
xnor U47216 (N_47216,N_46955,N_46430);
or U47217 (N_47217,N_46059,N_46588);
nor U47218 (N_47218,N_46535,N_46146);
xor U47219 (N_47219,N_46726,N_46234);
xnor U47220 (N_47220,N_46086,N_46692);
xor U47221 (N_47221,N_46382,N_46613);
xnor U47222 (N_47222,N_46724,N_46738);
nand U47223 (N_47223,N_46532,N_46080);
xnor U47224 (N_47224,N_46308,N_46171);
nand U47225 (N_47225,N_46040,N_46579);
and U47226 (N_47226,N_46231,N_46420);
nor U47227 (N_47227,N_46881,N_46401);
nor U47228 (N_47228,N_46832,N_46855);
nor U47229 (N_47229,N_46270,N_46464);
nor U47230 (N_47230,N_46940,N_46098);
nor U47231 (N_47231,N_46493,N_46170);
nor U47232 (N_47232,N_46730,N_46095);
and U47233 (N_47233,N_46749,N_46754);
and U47234 (N_47234,N_46476,N_46054);
and U47235 (N_47235,N_46404,N_46686);
xor U47236 (N_47236,N_46827,N_46208);
xnor U47237 (N_47237,N_46631,N_46536);
and U47238 (N_47238,N_46273,N_46071);
xor U47239 (N_47239,N_46709,N_46426);
and U47240 (N_47240,N_46206,N_46666);
nor U47241 (N_47241,N_46158,N_46078);
or U47242 (N_47242,N_46843,N_46226);
nor U47243 (N_47243,N_46155,N_46524);
and U47244 (N_47244,N_46391,N_46695);
and U47245 (N_47245,N_46954,N_46752);
xor U47246 (N_47246,N_46028,N_46590);
or U47247 (N_47247,N_46896,N_46362);
xor U47248 (N_47248,N_46267,N_46019);
and U47249 (N_47249,N_46807,N_46556);
or U47250 (N_47250,N_46025,N_46653);
or U47251 (N_47251,N_46878,N_46148);
and U47252 (N_47252,N_46992,N_46045);
and U47253 (N_47253,N_46378,N_46531);
nand U47254 (N_47254,N_46546,N_46468);
or U47255 (N_47255,N_46520,N_46151);
nand U47256 (N_47256,N_46413,N_46261);
nand U47257 (N_47257,N_46495,N_46093);
and U47258 (N_47258,N_46346,N_46869);
and U47259 (N_47259,N_46735,N_46061);
or U47260 (N_47260,N_46719,N_46478);
and U47261 (N_47261,N_46787,N_46771);
nand U47262 (N_47262,N_46620,N_46591);
and U47263 (N_47263,N_46801,N_46700);
nand U47264 (N_47264,N_46314,N_46849);
xor U47265 (N_47265,N_46852,N_46816);
nor U47266 (N_47266,N_46070,N_46780);
and U47267 (N_47267,N_46410,N_46338);
and U47268 (N_47268,N_46989,N_46825);
nand U47269 (N_47269,N_46910,N_46862);
nand U47270 (N_47270,N_46769,N_46112);
nand U47271 (N_47271,N_46283,N_46656);
xor U47272 (N_47272,N_46163,N_46411);
nand U47273 (N_47273,N_46534,N_46230);
nor U47274 (N_47274,N_46580,N_46438);
nand U47275 (N_47275,N_46186,N_46902);
nand U47276 (N_47276,N_46072,N_46982);
nor U47277 (N_47277,N_46814,N_46089);
or U47278 (N_47278,N_46141,N_46294);
xor U47279 (N_47279,N_46330,N_46377);
xor U47280 (N_47280,N_46837,N_46440);
nand U47281 (N_47281,N_46717,N_46110);
xor U47282 (N_47282,N_46611,N_46099);
xnor U47283 (N_47283,N_46979,N_46528);
nand U47284 (N_47284,N_46244,N_46265);
xor U47285 (N_47285,N_46002,N_46802);
and U47286 (N_47286,N_46509,N_46824);
and U47287 (N_47287,N_46756,N_46215);
and U47288 (N_47288,N_46037,N_46549);
nand U47289 (N_47289,N_46423,N_46907);
or U47290 (N_47290,N_46115,N_46193);
xnor U47291 (N_47291,N_46352,N_46757);
or U47292 (N_47292,N_46245,N_46051);
and U47293 (N_47293,N_46343,N_46854);
or U47294 (N_47294,N_46623,N_46687);
nand U47295 (N_47295,N_46444,N_46016);
or U47296 (N_47296,N_46897,N_46180);
nor U47297 (N_47297,N_46604,N_46781);
xnor U47298 (N_47298,N_46422,N_46861);
nand U47299 (N_47299,N_46454,N_46472);
xor U47300 (N_47300,N_46455,N_46467);
nor U47301 (N_47301,N_46305,N_46456);
nand U47302 (N_47302,N_46947,N_46926);
or U47303 (N_47303,N_46342,N_46610);
nor U47304 (N_47304,N_46618,N_46713);
nand U47305 (N_47305,N_46424,N_46917);
nand U47306 (N_47306,N_46798,N_46260);
or U47307 (N_47307,N_46331,N_46293);
xor U47308 (N_47308,N_46866,N_46042);
nor U47309 (N_47309,N_46436,N_46024);
xnor U47310 (N_47310,N_46412,N_46976);
nand U47311 (N_47311,N_46389,N_46494);
nand U47312 (N_47312,N_46041,N_46981);
and U47313 (N_47313,N_46138,N_46517);
nand U47314 (N_47314,N_46318,N_46038);
nand U47315 (N_47315,N_46648,N_46212);
and U47316 (N_47316,N_46490,N_46529);
and U47317 (N_47317,N_46598,N_46289);
or U47318 (N_47318,N_46487,N_46640);
or U47319 (N_47319,N_46173,N_46220);
nor U47320 (N_47320,N_46492,N_46211);
nor U47321 (N_47321,N_46831,N_46395);
and U47322 (N_47322,N_46884,N_46223);
nand U47323 (N_47323,N_46930,N_46983);
or U47324 (N_47324,N_46986,N_46238);
nand U47325 (N_47325,N_46437,N_46312);
or U47326 (N_47326,N_46665,N_46253);
nand U47327 (N_47327,N_46285,N_46916);
nand U47328 (N_47328,N_46397,N_46948);
and U47329 (N_47329,N_46111,N_46661);
or U47330 (N_47330,N_46320,N_46811);
xnor U47331 (N_47331,N_46662,N_46767);
nor U47332 (N_47332,N_46539,N_46658);
nor U47333 (N_47333,N_46309,N_46431);
and U47334 (N_47334,N_46502,N_46725);
nand U47335 (N_47335,N_46596,N_46104);
nor U47336 (N_47336,N_46052,N_46616);
nand U47337 (N_47337,N_46419,N_46162);
or U47338 (N_47338,N_46021,N_46514);
nor U47339 (N_47339,N_46693,N_46645);
xor U47340 (N_47340,N_46046,N_46592);
xnor U47341 (N_47341,N_46876,N_46636);
or U47342 (N_47342,N_46737,N_46845);
nor U47343 (N_47343,N_46937,N_46385);
or U47344 (N_47344,N_46249,N_46745);
nor U47345 (N_47345,N_46307,N_46919);
xor U47346 (N_47346,N_46791,N_46676);
or U47347 (N_47347,N_46288,N_46673);
and U47348 (N_47348,N_46914,N_46545);
nand U47349 (N_47349,N_46766,N_46405);
or U47350 (N_47350,N_46667,N_46882);
and U47351 (N_47351,N_46792,N_46315);
xor U47352 (N_47352,N_46796,N_46207);
xor U47353 (N_47353,N_46286,N_46939);
or U47354 (N_47354,N_46096,N_46232);
or U47355 (N_47355,N_46386,N_46913);
or U47356 (N_47356,N_46915,N_46049);
and U47357 (N_47357,N_46718,N_46210);
and U47358 (N_47358,N_46248,N_46540);
or U47359 (N_47359,N_46300,N_46856);
nor U47360 (N_47360,N_46477,N_46133);
nand U47361 (N_47361,N_46182,N_46710);
or U47362 (N_47362,N_46682,N_46263);
and U47363 (N_47363,N_46128,N_46121);
and U47364 (N_47364,N_46428,N_46911);
xor U47365 (N_47365,N_46600,N_46310);
nor U47366 (N_47366,N_46945,N_46739);
or U47367 (N_47367,N_46279,N_46782);
and U47368 (N_47368,N_46161,N_46154);
and U47369 (N_47369,N_46704,N_46734);
xor U47370 (N_47370,N_46768,N_46819);
and U47371 (N_47371,N_46553,N_46723);
and U47372 (N_47372,N_46840,N_46872);
nor U47373 (N_47373,N_46584,N_46371);
and U47374 (N_47374,N_46651,N_46817);
xor U47375 (N_47375,N_46132,N_46140);
and U47376 (N_47376,N_46621,N_46364);
or U47377 (N_47377,N_46347,N_46179);
nor U47378 (N_47378,N_46681,N_46381);
xor U47379 (N_47379,N_46703,N_46899);
or U47380 (N_47380,N_46571,N_46944);
xnor U47381 (N_47381,N_46762,N_46542);
nor U47382 (N_47382,N_46275,N_46683);
nor U47383 (N_47383,N_46933,N_46526);
xnor U47384 (N_47384,N_46360,N_46030);
and U47385 (N_47385,N_46779,N_46396);
xor U47386 (N_47386,N_46034,N_46400);
nor U47387 (N_47387,N_46720,N_46353);
nor U47388 (N_47388,N_46649,N_46271);
xnor U47389 (N_47389,N_46366,N_46672);
nor U47390 (N_47390,N_46292,N_46512);
nand U47391 (N_47391,N_46925,N_46850);
nand U47392 (N_47392,N_46479,N_46224);
nand U47393 (N_47393,N_46863,N_46217);
xnor U47394 (N_47394,N_46764,N_46469);
nor U47395 (N_47395,N_46194,N_46789);
nand U47396 (N_47396,N_46946,N_46552);
or U47397 (N_47397,N_46670,N_46885);
xnor U47398 (N_47398,N_46457,N_46027);
nor U47399 (N_47399,N_46557,N_46838);
xnor U47400 (N_47400,N_46131,N_46058);
xor U47401 (N_47401,N_46383,N_46607);
xnor U47402 (N_47402,N_46685,N_46329);
or U47403 (N_47403,N_46109,N_46066);
and U47404 (N_47404,N_46594,N_46776);
xnor U47405 (N_47405,N_46113,N_46139);
or U47406 (N_47406,N_46192,N_46612);
or U47407 (N_47407,N_46254,N_46987);
or U47408 (N_47408,N_46721,N_46407);
nand U47409 (N_47409,N_46633,N_46172);
nand U47410 (N_47410,N_46354,N_46453);
nor U47411 (N_47411,N_46251,N_46582);
nor U47412 (N_47412,N_46689,N_46236);
nand U47413 (N_47413,N_46429,N_46367);
and U47414 (N_47414,N_46063,N_46447);
and U47415 (N_47415,N_46175,N_46943);
or U47416 (N_47416,N_46470,N_46691);
nor U47417 (N_47417,N_46191,N_46145);
or U47418 (N_47418,N_46659,N_46544);
and U47419 (N_47419,N_46209,N_46345);
xnor U47420 (N_47420,N_46809,N_46246);
xor U47421 (N_47421,N_46627,N_46017);
xnor U47422 (N_47422,N_46555,N_46688);
and U47423 (N_47423,N_46924,N_46751);
and U47424 (N_47424,N_46822,N_46959);
nor U47425 (N_47425,N_46181,N_46340);
nand U47426 (N_47426,N_46728,N_46341);
xor U47427 (N_47427,N_46830,N_46256);
xnor U47428 (N_47428,N_46313,N_46777);
nor U47429 (N_47429,N_46793,N_46614);
or U47430 (N_47430,N_46259,N_46015);
and U47431 (N_47431,N_46388,N_46677);
or U47432 (N_47432,N_46599,N_46788);
or U47433 (N_47433,N_46324,N_46657);
xnor U47434 (N_47434,N_46629,N_46815);
or U47435 (N_47435,N_46736,N_46157);
and U47436 (N_47436,N_46291,N_46701);
xnor U47437 (N_47437,N_46706,N_46523);
nor U47438 (N_47438,N_46415,N_46103);
or U47439 (N_47439,N_46284,N_46055);
xor U47440 (N_47440,N_46921,N_46617);
or U47441 (N_47441,N_46778,N_46853);
xor U47442 (N_47442,N_46595,N_46835);
or U47443 (N_47443,N_46047,N_46583);
nor U47444 (N_47444,N_46336,N_46609);
nor U47445 (N_47445,N_46323,N_46550);
nand U47446 (N_47446,N_46794,N_46576);
nor U47447 (N_47447,N_46392,N_46187);
and U47448 (N_47448,N_46496,N_46698);
xnor U47449 (N_47449,N_46137,N_46886);
xnor U47450 (N_47450,N_46167,N_46974);
xor U47451 (N_47451,N_46004,N_46123);
nand U47452 (N_47452,N_46349,N_46117);
and U47453 (N_47453,N_46785,N_46335);
nand U47454 (N_47454,N_46597,N_46635);
xnor U47455 (N_47455,N_46606,N_46859);
or U47456 (N_47456,N_46906,N_46660);
xnor U47457 (N_47457,N_46506,N_46895);
xnor U47458 (N_47458,N_46898,N_46327);
and U47459 (N_47459,N_46883,N_46748);
nand U47460 (N_47460,N_46702,N_46804);
nand U47461 (N_47461,N_46011,N_46427);
and U47462 (N_47462,N_46626,N_46797);
and U47463 (N_47463,N_46759,N_46081);
or U47464 (N_47464,N_46290,N_46563);
nand U47465 (N_47465,N_46812,N_46018);
xnor U47466 (N_47466,N_46758,N_46449);
xnor U47467 (N_47467,N_46409,N_46783);
or U47468 (N_47468,N_46877,N_46214);
nand U47469 (N_47469,N_46650,N_46262);
xnor U47470 (N_47470,N_46973,N_46642);
and U47471 (N_47471,N_46304,N_46750);
and U47472 (N_47472,N_46368,N_46755);
nand U47473 (N_47473,N_46203,N_46561);
and U47474 (N_47474,N_46060,N_46475);
nor U47475 (N_47475,N_46483,N_46242);
nor U47476 (N_47476,N_46993,N_46829);
nor U47477 (N_47477,N_46177,N_46461);
and U47478 (N_47478,N_46800,N_46589);
nand U47479 (N_47479,N_46100,N_46229);
or U47480 (N_47480,N_46533,N_46416);
and U47481 (N_47481,N_46601,N_46999);
xnor U47482 (N_47482,N_46731,N_46605);
xnor U47483 (N_47483,N_46459,N_46359);
and U47484 (N_47484,N_46243,N_46195);
nor U47485 (N_47485,N_46441,N_46129);
and U47486 (N_47486,N_46239,N_46201);
xnor U47487 (N_47487,N_46799,N_46619);
nand U47488 (N_47488,N_46119,N_46743);
or U47489 (N_47489,N_46675,N_46630);
and U47490 (N_47490,N_46904,N_46684);
xnor U47491 (N_47491,N_46082,N_46564);
or U47492 (N_47492,N_46344,N_46570);
or U47493 (N_47493,N_46949,N_46567);
xnor U47494 (N_47494,N_46707,N_46964);
and U47495 (N_47495,N_46375,N_46136);
xnor U47496 (N_47496,N_46638,N_46967);
nor U47497 (N_47497,N_46962,N_46680);
xor U47498 (N_47498,N_46498,N_46960);
and U47499 (N_47499,N_46715,N_46643);
xor U47500 (N_47500,N_46072,N_46192);
or U47501 (N_47501,N_46089,N_46389);
and U47502 (N_47502,N_46465,N_46610);
and U47503 (N_47503,N_46951,N_46756);
xor U47504 (N_47504,N_46233,N_46037);
or U47505 (N_47505,N_46011,N_46924);
or U47506 (N_47506,N_46161,N_46376);
xnor U47507 (N_47507,N_46063,N_46635);
nor U47508 (N_47508,N_46815,N_46235);
or U47509 (N_47509,N_46541,N_46764);
nand U47510 (N_47510,N_46647,N_46720);
or U47511 (N_47511,N_46807,N_46686);
nor U47512 (N_47512,N_46130,N_46735);
xnor U47513 (N_47513,N_46250,N_46023);
or U47514 (N_47514,N_46169,N_46060);
nand U47515 (N_47515,N_46765,N_46601);
nor U47516 (N_47516,N_46960,N_46779);
nor U47517 (N_47517,N_46177,N_46615);
or U47518 (N_47518,N_46309,N_46841);
and U47519 (N_47519,N_46411,N_46429);
nand U47520 (N_47520,N_46626,N_46806);
or U47521 (N_47521,N_46005,N_46584);
or U47522 (N_47522,N_46893,N_46506);
xor U47523 (N_47523,N_46781,N_46497);
xnor U47524 (N_47524,N_46668,N_46904);
or U47525 (N_47525,N_46318,N_46965);
xor U47526 (N_47526,N_46341,N_46532);
nor U47527 (N_47527,N_46863,N_46053);
or U47528 (N_47528,N_46734,N_46173);
nor U47529 (N_47529,N_46240,N_46476);
nand U47530 (N_47530,N_46675,N_46347);
nand U47531 (N_47531,N_46047,N_46985);
nor U47532 (N_47532,N_46759,N_46196);
xnor U47533 (N_47533,N_46186,N_46497);
xor U47534 (N_47534,N_46397,N_46936);
nand U47535 (N_47535,N_46829,N_46894);
nand U47536 (N_47536,N_46720,N_46985);
and U47537 (N_47537,N_46709,N_46919);
nand U47538 (N_47538,N_46393,N_46118);
nand U47539 (N_47539,N_46476,N_46813);
nor U47540 (N_47540,N_46132,N_46929);
xnor U47541 (N_47541,N_46816,N_46966);
and U47542 (N_47542,N_46491,N_46554);
or U47543 (N_47543,N_46987,N_46677);
xor U47544 (N_47544,N_46027,N_46321);
nand U47545 (N_47545,N_46210,N_46418);
xor U47546 (N_47546,N_46371,N_46380);
or U47547 (N_47547,N_46440,N_46474);
nor U47548 (N_47548,N_46530,N_46498);
or U47549 (N_47549,N_46969,N_46123);
nand U47550 (N_47550,N_46931,N_46608);
xor U47551 (N_47551,N_46697,N_46471);
xnor U47552 (N_47552,N_46948,N_46597);
and U47553 (N_47553,N_46771,N_46090);
or U47554 (N_47554,N_46981,N_46768);
nor U47555 (N_47555,N_46928,N_46808);
nor U47556 (N_47556,N_46952,N_46177);
nor U47557 (N_47557,N_46119,N_46840);
or U47558 (N_47558,N_46999,N_46327);
xnor U47559 (N_47559,N_46432,N_46084);
or U47560 (N_47560,N_46407,N_46055);
and U47561 (N_47561,N_46251,N_46819);
nand U47562 (N_47562,N_46038,N_46093);
nor U47563 (N_47563,N_46440,N_46277);
nor U47564 (N_47564,N_46453,N_46046);
nor U47565 (N_47565,N_46359,N_46907);
nor U47566 (N_47566,N_46933,N_46579);
xor U47567 (N_47567,N_46347,N_46311);
nand U47568 (N_47568,N_46166,N_46524);
or U47569 (N_47569,N_46419,N_46066);
and U47570 (N_47570,N_46646,N_46393);
or U47571 (N_47571,N_46344,N_46723);
nor U47572 (N_47572,N_46968,N_46428);
nand U47573 (N_47573,N_46293,N_46903);
and U47574 (N_47574,N_46445,N_46156);
or U47575 (N_47575,N_46590,N_46541);
or U47576 (N_47576,N_46258,N_46100);
nor U47577 (N_47577,N_46530,N_46515);
xor U47578 (N_47578,N_46877,N_46335);
or U47579 (N_47579,N_46152,N_46675);
or U47580 (N_47580,N_46742,N_46064);
xnor U47581 (N_47581,N_46955,N_46100);
nor U47582 (N_47582,N_46518,N_46988);
and U47583 (N_47583,N_46000,N_46396);
or U47584 (N_47584,N_46720,N_46042);
nor U47585 (N_47585,N_46561,N_46407);
and U47586 (N_47586,N_46589,N_46486);
or U47587 (N_47587,N_46898,N_46536);
or U47588 (N_47588,N_46651,N_46338);
or U47589 (N_47589,N_46817,N_46621);
xnor U47590 (N_47590,N_46812,N_46688);
and U47591 (N_47591,N_46012,N_46459);
nor U47592 (N_47592,N_46686,N_46800);
and U47593 (N_47593,N_46199,N_46271);
and U47594 (N_47594,N_46399,N_46564);
or U47595 (N_47595,N_46506,N_46897);
and U47596 (N_47596,N_46916,N_46583);
xor U47597 (N_47597,N_46030,N_46897);
or U47598 (N_47598,N_46728,N_46936);
nand U47599 (N_47599,N_46691,N_46044);
and U47600 (N_47600,N_46315,N_46195);
and U47601 (N_47601,N_46931,N_46136);
nand U47602 (N_47602,N_46073,N_46749);
and U47603 (N_47603,N_46689,N_46417);
and U47604 (N_47604,N_46642,N_46214);
xor U47605 (N_47605,N_46887,N_46199);
or U47606 (N_47606,N_46223,N_46338);
nand U47607 (N_47607,N_46880,N_46353);
nand U47608 (N_47608,N_46584,N_46099);
nand U47609 (N_47609,N_46964,N_46158);
nor U47610 (N_47610,N_46863,N_46613);
or U47611 (N_47611,N_46876,N_46762);
xnor U47612 (N_47612,N_46910,N_46387);
nand U47613 (N_47613,N_46003,N_46322);
or U47614 (N_47614,N_46310,N_46622);
xnor U47615 (N_47615,N_46766,N_46228);
or U47616 (N_47616,N_46967,N_46044);
nand U47617 (N_47617,N_46172,N_46515);
and U47618 (N_47618,N_46175,N_46450);
nor U47619 (N_47619,N_46599,N_46393);
or U47620 (N_47620,N_46536,N_46552);
nor U47621 (N_47621,N_46785,N_46761);
nand U47622 (N_47622,N_46106,N_46114);
and U47623 (N_47623,N_46819,N_46561);
nor U47624 (N_47624,N_46434,N_46187);
or U47625 (N_47625,N_46766,N_46283);
and U47626 (N_47626,N_46815,N_46573);
and U47627 (N_47627,N_46303,N_46997);
and U47628 (N_47628,N_46798,N_46849);
and U47629 (N_47629,N_46546,N_46323);
or U47630 (N_47630,N_46528,N_46049);
nor U47631 (N_47631,N_46687,N_46733);
and U47632 (N_47632,N_46460,N_46532);
or U47633 (N_47633,N_46761,N_46932);
nand U47634 (N_47634,N_46921,N_46416);
nor U47635 (N_47635,N_46390,N_46252);
or U47636 (N_47636,N_46322,N_46406);
nor U47637 (N_47637,N_46907,N_46815);
nor U47638 (N_47638,N_46454,N_46783);
and U47639 (N_47639,N_46784,N_46774);
nor U47640 (N_47640,N_46464,N_46696);
nor U47641 (N_47641,N_46695,N_46735);
and U47642 (N_47642,N_46809,N_46440);
xnor U47643 (N_47643,N_46793,N_46847);
xnor U47644 (N_47644,N_46555,N_46395);
nor U47645 (N_47645,N_46425,N_46672);
and U47646 (N_47646,N_46947,N_46045);
or U47647 (N_47647,N_46817,N_46352);
and U47648 (N_47648,N_46483,N_46620);
or U47649 (N_47649,N_46499,N_46521);
nor U47650 (N_47650,N_46662,N_46191);
nor U47651 (N_47651,N_46569,N_46485);
or U47652 (N_47652,N_46108,N_46879);
nand U47653 (N_47653,N_46450,N_46768);
and U47654 (N_47654,N_46084,N_46504);
or U47655 (N_47655,N_46942,N_46080);
nor U47656 (N_47656,N_46429,N_46131);
and U47657 (N_47657,N_46481,N_46044);
or U47658 (N_47658,N_46002,N_46390);
nand U47659 (N_47659,N_46015,N_46675);
and U47660 (N_47660,N_46588,N_46399);
nor U47661 (N_47661,N_46010,N_46743);
nor U47662 (N_47662,N_46436,N_46819);
xnor U47663 (N_47663,N_46708,N_46567);
or U47664 (N_47664,N_46328,N_46370);
or U47665 (N_47665,N_46392,N_46934);
and U47666 (N_47666,N_46233,N_46897);
and U47667 (N_47667,N_46031,N_46817);
nor U47668 (N_47668,N_46925,N_46400);
nor U47669 (N_47669,N_46967,N_46124);
xor U47670 (N_47670,N_46676,N_46819);
nor U47671 (N_47671,N_46242,N_46780);
nor U47672 (N_47672,N_46389,N_46187);
or U47673 (N_47673,N_46494,N_46522);
and U47674 (N_47674,N_46209,N_46279);
and U47675 (N_47675,N_46272,N_46167);
and U47676 (N_47676,N_46817,N_46719);
nor U47677 (N_47677,N_46032,N_46931);
and U47678 (N_47678,N_46000,N_46100);
nand U47679 (N_47679,N_46412,N_46201);
xor U47680 (N_47680,N_46596,N_46611);
xor U47681 (N_47681,N_46638,N_46106);
nand U47682 (N_47682,N_46720,N_46500);
or U47683 (N_47683,N_46466,N_46580);
and U47684 (N_47684,N_46519,N_46952);
nand U47685 (N_47685,N_46768,N_46623);
or U47686 (N_47686,N_46556,N_46337);
and U47687 (N_47687,N_46308,N_46179);
xor U47688 (N_47688,N_46273,N_46396);
or U47689 (N_47689,N_46070,N_46189);
nor U47690 (N_47690,N_46891,N_46754);
nor U47691 (N_47691,N_46077,N_46592);
nor U47692 (N_47692,N_46020,N_46645);
nand U47693 (N_47693,N_46153,N_46545);
xnor U47694 (N_47694,N_46030,N_46135);
or U47695 (N_47695,N_46538,N_46777);
and U47696 (N_47696,N_46237,N_46173);
nand U47697 (N_47697,N_46010,N_46593);
or U47698 (N_47698,N_46134,N_46468);
nand U47699 (N_47699,N_46529,N_46391);
nand U47700 (N_47700,N_46957,N_46024);
nor U47701 (N_47701,N_46928,N_46271);
xnor U47702 (N_47702,N_46088,N_46804);
nor U47703 (N_47703,N_46468,N_46617);
or U47704 (N_47704,N_46230,N_46704);
and U47705 (N_47705,N_46706,N_46367);
nand U47706 (N_47706,N_46795,N_46640);
and U47707 (N_47707,N_46160,N_46876);
or U47708 (N_47708,N_46979,N_46223);
or U47709 (N_47709,N_46865,N_46888);
and U47710 (N_47710,N_46575,N_46998);
and U47711 (N_47711,N_46649,N_46006);
or U47712 (N_47712,N_46238,N_46239);
xnor U47713 (N_47713,N_46066,N_46442);
nand U47714 (N_47714,N_46619,N_46992);
and U47715 (N_47715,N_46182,N_46009);
or U47716 (N_47716,N_46312,N_46953);
xnor U47717 (N_47717,N_46061,N_46060);
xor U47718 (N_47718,N_46640,N_46268);
nand U47719 (N_47719,N_46399,N_46488);
xnor U47720 (N_47720,N_46804,N_46707);
nand U47721 (N_47721,N_46671,N_46573);
xnor U47722 (N_47722,N_46204,N_46212);
nor U47723 (N_47723,N_46021,N_46700);
xor U47724 (N_47724,N_46334,N_46877);
nand U47725 (N_47725,N_46750,N_46348);
xor U47726 (N_47726,N_46016,N_46416);
or U47727 (N_47727,N_46047,N_46388);
or U47728 (N_47728,N_46866,N_46046);
nor U47729 (N_47729,N_46700,N_46743);
xor U47730 (N_47730,N_46691,N_46737);
xnor U47731 (N_47731,N_46543,N_46415);
nor U47732 (N_47732,N_46923,N_46867);
or U47733 (N_47733,N_46233,N_46368);
xor U47734 (N_47734,N_46479,N_46999);
nor U47735 (N_47735,N_46636,N_46906);
xnor U47736 (N_47736,N_46872,N_46181);
xor U47737 (N_47737,N_46791,N_46669);
or U47738 (N_47738,N_46078,N_46705);
nand U47739 (N_47739,N_46866,N_46779);
or U47740 (N_47740,N_46980,N_46619);
and U47741 (N_47741,N_46310,N_46479);
or U47742 (N_47742,N_46775,N_46802);
nand U47743 (N_47743,N_46967,N_46217);
nand U47744 (N_47744,N_46002,N_46358);
nand U47745 (N_47745,N_46991,N_46014);
nor U47746 (N_47746,N_46488,N_46734);
or U47747 (N_47747,N_46931,N_46895);
or U47748 (N_47748,N_46573,N_46983);
nor U47749 (N_47749,N_46884,N_46147);
or U47750 (N_47750,N_46094,N_46250);
and U47751 (N_47751,N_46487,N_46854);
nor U47752 (N_47752,N_46886,N_46991);
xor U47753 (N_47753,N_46952,N_46655);
nand U47754 (N_47754,N_46429,N_46943);
nand U47755 (N_47755,N_46888,N_46605);
and U47756 (N_47756,N_46224,N_46042);
nor U47757 (N_47757,N_46255,N_46410);
nor U47758 (N_47758,N_46872,N_46395);
nand U47759 (N_47759,N_46951,N_46531);
or U47760 (N_47760,N_46755,N_46383);
nand U47761 (N_47761,N_46751,N_46166);
xor U47762 (N_47762,N_46705,N_46068);
and U47763 (N_47763,N_46059,N_46648);
and U47764 (N_47764,N_46686,N_46541);
and U47765 (N_47765,N_46779,N_46965);
and U47766 (N_47766,N_46222,N_46093);
and U47767 (N_47767,N_46886,N_46371);
and U47768 (N_47768,N_46956,N_46413);
nor U47769 (N_47769,N_46777,N_46200);
or U47770 (N_47770,N_46310,N_46617);
or U47771 (N_47771,N_46059,N_46667);
or U47772 (N_47772,N_46011,N_46358);
xnor U47773 (N_47773,N_46314,N_46357);
or U47774 (N_47774,N_46310,N_46004);
and U47775 (N_47775,N_46860,N_46036);
xor U47776 (N_47776,N_46545,N_46895);
xor U47777 (N_47777,N_46637,N_46872);
xor U47778 (N_47778,N_46318,N_46020);
or U47779 (N_47779,N_46893,N_46001);
xor U47780 (N_47780,N_46286,N_46910);
nand U47781 (N_47781,N_46770,N_46759);
xor U47782 (N_47782,N_46921,N_46430);
nand U47783 (N_47783,N_46165,N_46399);
or U47784 (N_47784,N_46466,N_46993);
nand U47785 (N_47785,N_46562,N_46652);
xor U47786 (N_47786,N_46017,N_46596);
or U47787 (N_47787,N_46497,N_46924);
nor U47788 (N_47788,N_46573,N_46668);
and U47789 (N_47789,N_46529,N_46880);
nor U47790 (N_47790,N_46434,N_46336);
nor U47791 (N_47791,N_46608,N_46923);
or U47792 (N_47792,N_46641,N_46989);
nor U47793 (N_47793,N_46908,N_46146);
and U47794 (N_47794,N_46869,N_46435);
and U47795 (N_47795,N_46343,N_46920);
and U47796 (N_47796,N_46798,N_46539);
nor U47797 (N_47797,N_46649,N_46202);
nand U47798 (N_47798,N_46813,N_46388);
and U47799 (N_47799,N_46246,N_46695);
or U47800 (N_47800,N_46460,N_46439);
xnor U47801 (N_47801,N_46800,N_46105);
or U47802 (N_47802,N_46976,N_46033);
xor U47803 (N_47803,N_46006,N_46018);
xnor U47804 (N_47804,N_46994,N_46513);
nor U47805 (N_47805,N_46754,N_46262);
xnor U47806 (N_47806,N_46044,N_46550);
nand U47807 (N_47807,N_46387,N_46902);
nor U47808 (N_47808,N_46551,N_46481);
xnor U47809 (N_47809,N_46133,N_46687);
nand U47810 (N_47810,N_46341,N_46706);
nor U47811 (N_47811,N_46526,N_46914);
xnor U47812 (N_47812,N_46999,N_46929);
xor U47813 (N_47813,N_46938,N_46419);
xnor U47814 (N_47814,N_46862,N_46922);
nor U47815 (N_47815,N_46864,N_46072);
or U47816 (N_47816,N_46683,N_46680);
nand U47817 (N_47817,N_46318,N_46139);
nand U47818 (N_47818,N_46600,N_46645);
xnor U47819 (N_47819,N_46498,N_46077);
nand U47820 (N_47820,N_46316,N_46860);
xnor U47821 (N_47821,N_46234,N_46434);
and U47822 (N_47822,N_46239,N_46322);
and U47823 (N_47823,N_46860,N_46732);
or U47824 (N_47824,N_46280,N_46954);
nor U47825 (N_47825,N_46078,N_46457);
nor U47826 (N_47826,N_46706,N_46841);
xor U47827 (N_47827,N_46222,N_46563);
xor U47828 (N_47828,N_46540,N_46780);
xor U47829 (N_47829,N_46557,N_46275);
xnor U47830 (N_47830,N_46257,N_46285);
nor U47831 (N_47831,N_46357,N_46292);
xnor U47832 (N_47832,N_46266,N_46094);
or U47833 (N_47833,N_46745,N_46861);
and U47834 (N_47834,N_46378,N_46079);
and U47835 (N_47835,N_46976,N_46184);
nor U47836 (N_47836,N_46644,N_46271);
xnor U47837 (N_47837,N_46730,N_46172);
nand U47838 (N_47838,N_46243,N_46585);
nor U47839 (N_47839,N_46539,N_46383);
nand U47840 (N_47840,N_46251,N_46026);
xnor U47841 (N_47841,N_46527,N_46847);
nor U47842 (N_47842,N_46281,N_46515);
and U47843 (N_47843,N_46511,N_46588);
and U47844 (N_47844,N_46205,N_46193);
and U47845 (N_47845,N_46547,N_46824);
nand U47846 (N_47846,N_46047,N_46837);
or U47847 (N_47847,N_46114,N_46644);
xnor U47848 (N_47848,N_46015,N_46551);
nand U47849 (N_47849,N_46806,N_46247);
and U47850 (N_47850,N_46541,N_46458);
or U47851 (N_47851,N_46276,N_46061);
nand U47852 (N_47852,N_46711,N_46509);
and U47853 (N_47853,N_46287,N_46771);
and U47854 (N_47854,N_46170,N_46544);
and U47855 (N_47855,N_46554,N_46900);
nor U47856 (N_47856,N_46188,N_46881);
xor U47857 (N_47857,N_46415,N_46069);
nand U47858 (N_47858,N_46647,N_46266);
or U47859 (N_47859,N_46194,N_46978);
and U47860 (N_47860,N_46928,N_46619);
xor U47861 (N_47861,N_46828,N_46130);
nor U47862 (N_47862,N_46003,N_46993);
nand U47863 (N_47863,N_46315,N_46303);
or U47864 (N_47864,N_46247,N_46980);
nor U47865 (N_47865,N_46667,N_46185);
nand U47866 (N_47866,N_46267,N_46707);
or U47867 (N_47867,N_46505,N_46866);
and U47868 (N_47868,N_46266,N_46439);
or U47869 (N_47869,N_46562,N_46242);
nand U47870 (N_47870,N_46940,N_46117);
xnor U47871 (N_47871,N_46615,N_46664);
nor U47872 (N_47872,N_46847,N_46595);
and U47873 (N_47873,N_46126,N_46674);
xnor U47874 (N_47874,N_46929,N_46996);
xnor U47875 (N_47875,N_46362,N_46467);
nor U47876 (N_47876,N_46503,N_46632);
xnor U47877 (N_47877,N_46012,N_46600);
or U47878 (N_47878,N_46037,N_46411);
xnor U47879 (N_47879,N_46376,N_46699);
or U47880 (N_47880,N_46459,N_46268);
and U47881 (N_47881,N_46174,N_46548);
nand U47882 (N_47882,N_46429,N_46986);
or U47883 (N_47883,N_46874,N_46548);
xor U47884 (N_47884,N_46463,N_46033);
xor U47885 (N_47885,N_46342,N_46028);
nand U47886 (N_47886,N_46652,N_46251);
xor U47887 (N_47887,N_46504,N_46842);
nand U47888 (N_47888,N_46601,N_46764);
and U47889 (N_47889,N_46451,N_46648);
nor U47890 (N_47890,N_46102,N_46566);
and U47891 (N_47891,N_46104,N_46887);
and U47892 (N_47892,N_46955,N_46305);
and U47893 (N_47893,N_46069,N_46227);
nor U47894 (N_47894,N_46227,N_46853);
xor U47895 (N_47895,N_46470,N_46642);
nor U47896 (N_47896,N_46595,N_46592);
nor U47897 (N_47897,N_46111,N_46585);
or U47898 (N_47898,N_46769,N_46113);
xor U47899 (N_47899,N_46999,N_46749);
xor U47900 (N_47900,N_46918,N_46292);
or U47901 (N_47901,N_46070,N_46280);
and U47902 (N_47902,N_46435,N_46150);
or U47903 (N_47903,N_46874,N_46390);
and U47904 (N_47904,N_46058,N_46088);
and U47905 (N_47905,N_46207,N_46321);
nor U47906 (N_47906,N_46809,N_46761);
nand U47907 (N_47907,N_46244,N_46805);
or U47908 (N_47908,N_46123,N_46272);
and U47909 (N_47909,N_46361,N_46594);
nor U47910 (N_47910,N_46302,N_46865);
nand U47911 (N_47911,N_46128,N_46462);
or U47912 (N_47912,N_46948,N_46059);
and U47913 (N_47913,N_46819,N_46213);
nor U47914 (N_47914,N_46688,N_46609);
xnor U47915 (N_47915,N_46641,N_46946);
and U47916 (N_47916,N_46353,N_46691);
and U47917 (N_47917,N_46286,N_46434);
nor U47918 (N_47918,N_46745,N_46437);
xnor U47919 (N_47919,N_46863,N_46501);
nor U47920 (N_47920,N_46899,N_46510);
nand U47921 (N_47921,N_46312,N_46676);
and U47922 (N_47922,N_46813,N_46174);
nor U47923 (N_47923,N_46057,N_46061);
or U47924 (N_47924,N_46582,N_46513);
nor U47925 (N_47925,N_46193,N_46726);
nor U47926 (N_47926,N_46003,N_46109);
nor U47927 (N_47927,N_46921,N_46131);
nand U47928 (N_47928,N_46463,N_46935);
and U47929 (N_47929,N_46409,N_46416);
nor U47930 (N_47930,N_46028,N_46585);
and U47931 (N_47931,N_46595,N_46205);
and U47932 (N_47932,N_46847,N_46720);
nor U47933 (N_47933,N_46868,N_46736);
xnor U47934 (N_47934,N_46467,N_46570);
nand U47935 (N_47935,N_46650,N_46965);
xor U47936 (N_47936,N_46618,N_46174);
or U47937 (N_47937,N_46836,N_46212);
nor U47938 (N_47938,N_46090,N_46311);
xor U47939 (N_47939,N_46644,N_46303);
nor U47940 (N_47940,N_46473,N_46328);
nor U47941 (N_47941,N_46742,N_46684);
nand U47942 (N_47942,N_46814,N_46633);
nand U47943 (N_47943,N_46177,N_46395);
xor U47944 (N_47944,N_46458,N_46938);
xnor U47945 (N_47945,N_46391,N_46592);
or U47946 (N_47946,N_46033,N_46080);
and U47947 (N_47947,N_46843,N_46955);
xor U47948 (N_47948,N_46575,N_46569);
and U47949 (N_47949,N_46455,N_46496);
or U47950 (N_47950,N_46540,N_46790);
nand U47951 (N_47951,N_46262,N_46120);
nand U47952 (N_47952,N_46474,N_46368);
xor U47953 (N_47953,N_46608,N_46963);
or U47954 (N_47954,N_46106,N_46585);
or U47955 (N_47955,N_46608,N_46916);
and U47956 (N_47956,N_46475,N_46977);
xnor U47957 (N_47957,N_46465,N_46938);
nor U47958 (N_47958,N_46423,N_46931);
or U47959 (N_47959,N_46927,N_46182);
nor U47960 (N_47960,N_46690,N_46922);
nand U47961 (N_47961,N_46993,N_46158);
and U47962 (N_47962,N_46419,N_46192);
or U47963 (N_47963,N_46400,N_46710);
and U47964 (N_47964,N_46418,N_46965);
or U47965 (N_47965,N_46631,N_46932);
xor U47966 (N_47966,N_46418,N_46389);
nand U47967 (N_47967,N_46188,N_46452);
nor U47968 (N_47968,N_46306,N_46856);
or U47969 (N_47969,N_46947,N_46601);
nor U47970 (N_47970,N_46376,N_46824);
nand U47971 (N_47971,N_46927,N_46190);
xnor U47972 (N_47972,N_46141,N_46662);
and U47973 (N_47973,N_46165,N_46659);
and U47974 (N_47974,N_46318,N_46541);
nand U47975 (N_47975,N_46467,N_46292);
xor U47976 (N_47976,N_46832,N_46724);
or U47977 (N_47977,N_46721,N_46864);
nand U47978 (N_47978,N_46909,N_46645);
or U47979 (N_47979,N_46637,N_46576);
nand U47980 (N_47980,N_46929,N_46135);
nand U47981 (N_47981,N_46271,N_46277);
nor U47982 (N_47982,N_46577,N_46771);
nand U47983 (N_47983,N_46811,N_46318);
nand U47984 (N_47984,N_46055,N_46063);
and U47985 (N_47985,N_46440,N_46476);
nor U47986 (N_47986,N_46644,N_46214);
nor U47987 (N_47987,N_46346,N_46900);
nor U47988 (N_47988,N_46516,N_46178);
xor U47989 (N_47989,N_46534,N_46258);
nor U47990 (N_47990,N_46073,N_46459);
and U47991 (N_47991,N_46446,N_46060);
and U47992 (N_47992,N_46261,N_46990);
and U47993 (N_47993,N_46057,N_46371);
nand U47994 (N_47994,N_46437,N_46176);
nor U47995 (N_47995,N_46068,N_46361);
or U47996 (N_47996,N_46665,N_46794);
xnor U47997 (N_47997,N_46045,N_46174);
xor U47998 (N_47998,N_46661,N_46159);
nand U47999 (N_47999,N_46290,N_46301);
xor U48000 (N_48000,N_47100,N_47113);
and U48001 (N_48001,N_47845,N_47711);
nor U48002 (N_48002,N_47124,N_47508);
nor U48003 (N_48003,N_47268,N_47614);
and U48004 (N_48004,N_47252,N_47768);
or U48005 (N_48005,N_47696,N_47609);
nor U48006 (N_48006,N_47802,N_47451);
xor U48007 (N_48007,N_47267,N_47161);
or U48008 (N_48008,N_47803,N_47649);
or U48009 (N_48009,N_47436,N_47042);
nor U48010 (N_48010,N_47652,N_47262);
or U48011 (N_48011,N_47815,N_47705);
nand U48012 (N_48012,N_47779,N_47567);
nor U48013 (N_48013,N_47141,N_47187);
xor U48014 (N_48014,N_47559,N_47443);
or U48015 (N_48015,N_47002,N_47008);
nor U48016 (N_48016,N_47497,N_47441);
nor U48017 (N_48017,N_47704,N_47073);
nor U48018 (N_48018,N_47055,N_47307);
and U48019 (N_48019,N_47345,N_47112);
nor U48020 (N_48020,N_47931,N_47438);
xor U48021 (N_48021,N_47994,N_47261);
and U48022 (N_48022,N_47388,N_47725);
nand U48023 (N_48023,N_47525,N_47374);
nor U48024 (N_48024,N_47843,N_47075);
and U48025 (N_48025,N_47203,N_47738);
or U48026 (N_48026,N_47852,N_47185);
and U48027 (N_48027,N_47901,N_47592);
nor U48028 (N_48028,N_47353,N_47236);
xnor U48029 (N_48029,N_47360,N_47174);
xor U48030 (N_48030,N_47624,N_47882);
xor U48031 (N_48031,N_47357,N_47908);
and U48032 (N_48032,N_47076,N_47708);
nand U48033 (N_48033,N_47201,N_47766);
and U48034 (N_48034,N_47283,N_47759);
and U48035 (N_48035,N_47937,N_47190);
xnor U48036 (N_48036,N_47968,N_47538);
xor U48037 (N_48037,N_47133,N_47256);
nor U48038 (N_48038,N_47051,N_47965);
nor U48039 (N_48039,N_47933,N_47814);
and U48040 (N_48040,N_47390,N_47707);
xnor U48041 (N_48041,N_47912,N_47665);
nor U48042 (N_48042,N_47993,N_47231);
nor U48043 (N_48043,N_47499,N_47688);
or U48044 (N_48044,N_47160,N_47461);
or U48045 (N_48045,N_47217,N_47315);
xnor U48046 (N_48046,N_47640,N_47781);
and U48047 (N_48047,N_47975,N_47167);
or U48048 (N_48048,N_47524,N_47849);
or U48049 (N_48049,N_47054,N_47862);
xnor U48050 (N_48050,N_47980,N_47930);
nor U48051 (N_48051,N_47566,N_47023);
nor U48052 (N_48052,N_47039,N_47173);
xor U48053 (N_48053,N_47215,N_47188);
and U48054 (N_48054,N_47924,N_47335);
or U48055 (N_48055,N_47093,N_47864);
xnor U48056 (N_48056,N_47354,N_47402);
nor U48057 (N_48057,N_47134,N_47506);
nand U48058 (N_48058,N_47312,N_47774);
nand U48059 (N_48059,N_47898,N_47367);
and U48060 (N_48060,N_47229,N_47954);
xor U48061 (N_48061,N_47866,N_47128);
and U48062 (N_48062,N_47899,N_47208);
nand U48063 (N_48063,N_47721,N_47736);
or U48064 (N_48064,N_47029,N_47309);
nand U48065 (N_48065,N_47485,N_47507);
or U48066 (N_48066,N_47484,N_47286);
nor U48067 (N_48067,N_47305,N_47597);
xor U48068 (N_48068,N_47383,N_47145);
nor U48069 (N_48069,N_47021,N_47394);
nor U48070 (N_48070,N_47162,N_47593);
nand U48071 (N_48071,N_47751,N_47847);
xnor U48072 (N_48072,N_47590,N_47154);
nand U48073 (N_48073,N_47637,N_47384);
nor U48074 (N_48074,N_47366,N_47272);
or U48075 (N_48075,N_47420,N_47522);
nand U48076 (N_48076,N_47311,N_47660);
nor U48077 (N_48077,N_47427,N_47944);
nor U48078 (N_48078,N_47156,N_47210);
nor U48079 (N_48079,N_47453,N_47433);
xor U48080 (N_48080,N_47765,N_47961);
nor U48081 (N_48081,N_47728,N_47428);
or U48082 (N_48082,N_47547,N_47004);
and U48083 (N_48083,N_47958,N_47121);
and U48084 (N_48084,N_47117,N_47581);
xnor U48085 (N_48085,N_47056,N_47998);
and U48086 (N_48086,N_47532,N_47411);
and U48087 (N_48087,N_47419,N_47615);
or U48088 (N_48088,N_47977,N_47118);
xnor U48089 (N_48089,N_47046,N_47047);
nor U48090 (N_48090,N_47656,N_47602);
xor U48091 (N_48091,N_47697,N_47372);
nand U48092 (N_48092,N_47209,N_47601);
nand U48093 (N_48093,N_47833,N_47137);
nor U48094 (N_48094,N_47646,N_47359);
nor U48095 (N_48095,N_47698,N_47009);
nor U48096 (N_48096,N_47491,N_47891);
nand U48097 (N_48097,N_47139,N_47713);
nand U48098 (N_48098,N_47196,N_47037);
xor U48099 (N_48099,N_47942,N_47683);
and U48100 (N_48100,N_47483,N_47985);
xnor U48101 (N_48101,N_47929,N_47594);
and U48102 (N_48102,N_47786,N_47396);
xnor U48103 (N_48103,N_47885,N_47537);
and U48104 (N_48104,N_47099,N_47407);
and U48105 (N_48105,N_47745,N_47880);
nand U48106 (N_48106,N_47923,N_47595);
or U48107 (N_48107,N_47867,N_47049);
and U48108 (N_48108,N_47431,N_47111);
nor U48109 (N_48109,N_47316,N_47621);
nor U48110 (N_48110,N_47990,N_47691);
nand U48111 (N_48111,N_47747,N_47775);
or U48112 (N_48112,N_47276,N_47278);
or U48113 (N_48113,N_47523,N_47176);
and U48114 (N_48114,N_47169,N_47290);
and U48115 (N_48115,N_47531,N_47519);
xnor U48116 (N_48116,N_47580,N_47545);
or U48117 (N_48117,N_47680,N_47999);
or U48118 (N_48118,N_47025,N_47148);
xor U48119 (N_48119,N_47031,N_47772);
nand U48120 (N_48120,N_47586,N_47058);
or U48121 (N_48121,N_47344,N_47067);
and U48122 (N_48122,N_47719,N_47887);
xnor U48123 (N_48123,N_47064,N_47274);
and U48124 (N_48124,N_47540,N_47446);
or U48125 (N_48125,N_47604,N_47082);
or U48126 (N_48126,N_47466,N_47724);
or U48127 (N_48127,N_47239,N_47655);
nand U48128 (N_48128,N_47838,N_47414);
nor U48129 (N_48129,N_47295,N_47304);
and U48130 (N_48130,N_47598,N_47098);
nand U48131 (N_48131,N_47735,N_47501);
xor U48132 (N_48132,N_47269,N_47789);
nor U48133 (N_48133,N_47914,N_47103);
and U48134 (N_48134,N_47184,N_47462);
or U48135 (N_48135,N_47654,N_47753);
and U48136 (N_48136,N_47643,N_47539);
xor U48137 (N_48137,N_47478,N_47007);
nor U48138 (N_48138,N_47079,N_47000);
nor U48139 (N_48139,N_47279,N_47518);
or U48140 (N_48140,N_47489,N_47906);
xor U48141 (N_48141,N_47458,N_47569);
and U48142 (N_48142,N_47417,N_47361);
nor U48143 (N_48143,N_47758,N_47257);
and U48144 (N_48144,N_47066,N_47243);
xor U48145 (N_48145,N_47676,N_47636);
xnor U48146 (N_48146,N_47945,N_47726);
nor U48147 (N_48147,N_47535,N_47213);
nand U48148 (N_48148,N_47149,N_47627);
nor U48149 (N_48149,N_47780,N_47626);
nand U48150 (N_48150,N_47342,N_47541);
nor U48151 (N_48151,N_47973,N_47858);
or U48152 (N_48152,N_47808,N_47432);
nand U48153 (N_48153,N_47425,N_47130);
nand U48154 (N_48154,N_47495,N_47804);
and U48155 (N_48155,N_47953,N_47920);
or U48156 (N_48156,N_47633,N_47378);
and U48157 (N_48157,N_47555,N_47763);
nor U48158 (N_48158,N_47138,N_47952);
nor U48159 (N_48159,N_47827,N_47258);
and U48160 (N_48160,N_47327,N_47116);
nand U48161 (N_48161,N_47526,N_47101);
or U48162 (N_48162,N_47024,N_47895);
xnor U48163 (N_48163,N_47785,N_47505);
nand U48164 (N_48164,N_47632,N_47080);
nand U48165 (N_48165,N_47907,N_47041);
nor U48166 (N_48166,N_47421,N_47510);
nand U48167 (N_48167,N_47227,N_47668);
xnor U48168 (N_48168,N_47608,N_47260);
nand U48169 (N_48169,N_47065,N_47313);
xor U48170 (N_48170,N_47369,N_47232);
xnor U48171 (N_48171,N_47835,N_47701);
or U48172 (N_48172,N_47589,N_47338);
nor U48173 (N_48173,N_47872,N_47142);
nor U48174 (N_48174,N_47574,N_47317);
nor U48175 (N_48175,N_47797,N_47163);
xor U48176 (N_48176,N_47890,N_47465);
or U48177 (N_48177,N_47870,N_47198);
or U48178 (N_48178,N_47795,N_47669);
and U48179 (N_48179,N_47812,N_47263);
xor U48180 (N_48180,N_47909,N_47081);
nor U48181 (N_48181,N_47346,N_47500);
nor U48182 (N_48182,N_47410,N_47036);
nor U48183 (N_48183,N_47405,N_47424);
xor U48184 (N_48184,N_47333,N_47886);
and U48185 (N_48185,N_47140,N_47913);
nand U48186 (N_48186,N_47230,N_47463);
xor U48187 (N_48187,N_47219,N_47622);
xnor U48188 (N_48188,N_47385,N_47810);
and U48189 (N_48189,N_47972,N_47693);
nand U48190 (N_48190,N_47387,N_47509);
nand U48191 (N_48191,N_47755,N_47828);
and U48192 (N_48192,N_47107,N_47984);
nor U48193 (N_48193,N_47306,N_47528);
xnor U48194 (N_48194,N_47962,N_47634);
and U48195 (N_48195,N_47404,N_47964);
or U48196 (N_48196,N_47105,N_47271);
nor U48197 (N_48197,N_47259,N_47587);
xor U48198 (N_48198,N_47800,N_47741);
or U48199 (N_48199,N_47266,N_47444);
nand U48200 (N_48200,N_47712,N_47090);
xor U48201 (N_48201,N_47254,N_47883);
and U48202 (N_48202,N_47855,N_47158);
nor U48203 (N_48203,N_47896,N_47784);
nor U48204 (N_48204,N_47350,N_47771);
xor U48205 (N_48205,N_47293,N_47514);
or U48206 (N_48206,N_47381,N_47343);
xnor U48207 (N_48207,N_47299,N_47692);
nor U48208 (N_48208,N_47440,N_47644);
and U48209 (N_48209,N_47413,N_47332);
and U48210 (N_48210,N_47610,N_47147);
and U48211 (N_48211,N_47034,N_47694);
nor U48212 (N_48212,N_47430,N_47481);
nand U48213 (N_48213,N_47416,N_47600);
nand U48214 (N_48214,N_47630,N_47238);
xnor U48215 (N_48215,N_47275,N_47233);
and U48216 (N_48216,N_47328,N_47948);
and U48217 (N_48217,N_47207,N_47578);
nor U48218 (N_48218,N_47799,N_47879);
nor U48219 (N_48219,N_47482,N_47546);
nand U48220 (N_48220,N_47474,N_47470);
and U48221 (N_48221,N_47194,N_47679);
xor U48222 (N_48222,N_47788,N_47352);
and U48223 (N_48223,N_47645,N_47573);
xnor U48224 (N_48224,N_47435,N_47934);
nand U48225 (N_48225,N_47302,N_47502);
and U48226 (N_48226,N_47010,N_47926);
and U48227 (N_48227,N_47992,N_47770);
nand U48228 (N_48228,N_47853,N_47830);
nand U48229 (N_48229,N_47143,N_47368);
and U48230 (N_48230,N_47480,N_47681);
nand U48231 (N_48231,N_47826,N_47938);
xnor U48232 (N_48232,N_47337,N_47362);
xor U48233 (N_48233,N_47068,N_47617);
nor U48234 (N_48234,N_47970,N_47748);
nor U48235 (N_48235,N_47949,N_47153);
and U48236 (N_48236,N_47556,N_47991);
and U48237 (N_48237,N_47186,N_47022);
nor U48238 (N_48238,N_47677,N_47277);
and U48239 (N_48239,N_47695,N_47248);
and U48240 (N_48240,N_47550,N_47400);
nor U48241 (N_48241,N_47603,N_47863);
nor U48242 (N_48242,N_47324,N_47019);
nor U48243 (N_48243,N_47494,N_47742);
and U48244 (N_48244,N_47119,N_47840);
and U48245 (N_48245,N_47191,N_47135);
and U48246 (N_48246,N_47012,N_47083);
and U48247 (N_48247,N_47832,N_47061);
nand U48248 (N_48248,N_47809,N_47796);
xnor U48249 (N_48249,N_47776,N_47310);
xnor U48250 (N_48250,N_47287,N_47653);
nand U48251 (N_48251,N_47270,N_47534);
nor U48252 (N_48252,N_47437,N_47146);
or U48253 (N_48253,N_47875,N_47422);
xnor U48254 (N_48254,N_47925,N_47513);
nor U48255 (N_48255,N_47816,N_47997);
nand U48256 (N_48256,N_47897,N_47894);
or U48257 (N_48257,N_47222,N_47571);
nor U48258 (N_48258,N_47418,N_47957);
nor U48259 (N_48259,N_47941,N_47445);
nor U48260 (N_48260,N_47635,N_47631);
nand U48261 (N_48261,N_47108,N_47792);
or U48262 (N_48262,N_47981,N_47322);
and U48263 (N_48263,N_47658,N_47159);
or U48264 (N_48264,N_47006,N_47249);
or U48265 (N_48265,N_47983,N_47666);
and U48266 (N_48266,N_47710,N_47314);
xnor U48267 (N_48267,N_47206,N_47746);
and U48268 (N_48268,N_47558,N_47166);
nor U48269 (N_48269,N_47490,N_47469);
or U48270 (N_48270,N_47717,N_47996);
xnor U48271 (N_48271,N_47729,N_47439);
nor U48272 (N_48272,N_47043,N_47399);
nand U48273 (N_48273,N_47091,N_47503);
nor U48274 (N_48274,N_47044,N_47177);
or U48275 (N_48275,N_47364,N_47122);
xor U48276 (N_48276,N_47255,N_47211);
or U48277 (N_48277,N_47641,N_47181);
and U48278 (N_48278,N_47479,N_47805);
xor U48279 (N_48279,N_47686,N_47842);
xnor U48280 (N_48280,N_47892,N_47069);
xnor U48281 (N_48281,N_47251,N_47195);
or U48282 (N_48282,N_47752,N_47092);
xnor U48283 (N_48283,N_47987,N_47690);
xor U48284 (N_48284,N_47038,N_47123);
or U48285 (N_48285,N_47356,N_47449);
xor U48286 (N_48286,N_47200,N_47951);
or U48287 (N_48287,N_47563,N_47020);
and U48288 (N_48288,N_47955,N_47672);
or U48289 (N_48289,N_47801,N_47459);
nand U48290 (N_48290,N_47492,N_47819);
nand U48291 (N_48291,N_47171,N_47591);
and U48292 (N_48292,N_47976,N_47409);
xor U48293 (N_48293,N_47865,N_47454);
nor U48294 (N_48294,N_47115,N_47289);
nor U48295 (N_48295,N_47613,N_47193);
or U48296 (N_48296,N_47189,N_47831);
nand U48297 (N_48297,N_47226,N_47429);
or U48298 (N_48298,N_47033,N_47183);
or U48299 (N_48299,N_47172,N_47442);
or U48300 (N_48300,N_47423,N_47723);
xor U48301 (N_48301,N_47979,N_47915);
xnor U48302 (N_48302,N_47859,N_47778);
xnor U48303 (N_48303,N_47301,N_47889);
and U48304 (N_48304,N_47253,N_47638);
nor U48305 (N_48305,N_47486,N_47678);
and U48306 (N_48306,N_47235,N_47401);
nand U48307 (N_48307,N_47448,N_47918);
nor U48308 (N_48308,N_47861,N_47087);
nor U48309 (N_48309,N_47165,N_47062);
nand U48310 (N_48310,N_47032,N_47319);
and U48311 (N_48311,N_47877,N_47702);
xnor U48312 (N_48312,N_47714,N_47016);
nor U48313 (N_48313,N_47553,N_47671);
nor U48314 (N_48314,N_47294,N_47959);
or U48315 (N_48315,N_47850,N_47089);
nand U48316 (N_48316,N_47699,N_47732);
nor U48317 (N_48317,N_47308,N_47406);
xor U48318 (N_48318,N_47291,N_47722);
and U48319 (N_48319,N_47709,N_47205);
and U48320 (N_48320,N_47572,N_47986);
nand U48321 (N_48321,N_47989,N_47504);
or U48322 (N_48322,N_47472,N_47329);
nand U48323 (N_48323,N_47059,N_47922);
and U48324 (N_48324,N_47052,N_47839);
or U48325 (N_48325,N_47131,N_47647);
and U48326 (N_48326,N_47223,N_47182);
or U48327 (N_48327,N_47393,N_47214);
nand U48328 (N_48328,N_47351,N_47946);
xnor U48329 (N_48329,N_47689,N_47876);
xor U48330 (N_48330,N_47136,N_47086);
nor U48331 (N_48331,N_47579,N_47928);
nand U48332 (N_48332,N_47794,N_47860);
or U48333 (N_48333,N_47734,N_47325);
xor U48334 (N_48334,N_47575,N_47365);
nand U48335 (N_48335,N_47242,N_47629);
and U48336 (N_48336,N_47434,N_47077);
nor U48337 (N_48337,N_47910,N_47074);
nor U48338 (N_48338,N_47102,N_47667);
xnor U48339 (N_48339,N_47028,N_47533);
nor U48340 (N_48340,N_47341,N_47282);
or U48341 (N_48341,N_47935,N_47040);
xor U48342 (N_48342,N_47408,N_47857);
or U48343 (N_48343,N_47212,N_47822);
xnor U48344 (N_48344,N_47967,N_47783);
and U48345 (N_48345,N_47403,N_47129);
nor U48346 (N_48346,N_47936,N_47498);
or U48347 (N_48347,N_47927,N_47767);
nor U48348 (N_48348,N_47588,N_47718);
nor U48349 (N_48349,N_47648,N_47798);
nor U48350 (N_48350,N_47095,N_47884);
or U48351 (N_48351,N_47829,N_47460);
xor U48352 (N_48352,N_47782,N_47557);
nand U48353 (N_48353,N_47577,N_47197);
or U48354 (N_48354,N_47568,N_47670);
nand U48355 (N_48355,N_47339,N_47905);
or U48356 (N_48356,N_47921,N_47806);
xnor U48357 (N_48357,N_47625,N_47606);
or U48358 (N_48358,N_47764,N_47731);
nand U48359 (N_48359,N_47974,N_47228);
xnor U48360 (N_48360,N_47218,N_47720);
xnor U48361 (N_48361,N_47576,N_47285);
xnor U48362 (N_48362,N_47811,N_47412);
and U48363 (N_48363,N_47334,N_47488);
nor U48364 (N_48364,N_47902,N_47246);
xor U48365 (N_48365,N_47241,N_47072);
nor U48366 (N_48366,N_47003,N_47216);
nand U48367 (N_48367,N_47358,N_47088);
xor U48368 (N_48368,N_47841,N_47966);
or U48369 (N_48369,N_47265,N_47762);
and U48370 (N_48370,N_47940,N_47045);
and U48371 (N_48371,N_47084,N_47565);
nor U48372 (N_48372,N_47094,N_47303);
nor U48373 (N_48373,N_47097,N_47114);
or U48374 (N_48374,N_47754,N_47326);
and U48375 (N_48375,N_47150,N_47628);
nand U48376 (N_48376,N_47126,N_47180);
nor U48377 (N_48377,N_47749,N_47706);
nor U48378 (N_48378,N_47247,N_47464);
xor U48379 (N_48379,N_47280,N_47684);
or U48380 (N_48380,N_47297,N_47225);
nor U48381 (N_48381,N_47818,N_47371);
nand U48382 (N_48382,N_47960,N_47727);
nor U48383 (N_48383,N_47001,N_47529);
nor U48384 (N_48384,N_47456,N_47426);
nor U48385 (N_48385,N_47651,N_47817);
nand U48386 (N_48386,N_47292,N_47607);
nand U48387 (N_48387,N_47616,N_47048);
and U48388 (N_48388,N_47455,N_47769);
or U48389 (N_48389,N_47823,N_47564);
or U48390 (N_48390,N_47947,N_47836);
nand U48391 (N_48391,N_47281,N_47825);
xor U48392 (N_48392,N_47750,N_47848);
xnor U48393 (N_48393,N_47932,N_47380);
nand U48394 (N_48394,N_47675,N_47834);
and U48395 (N_48395,N_47982,N_47548);
and U48396 (N_48396,N_47026,N_47813);
xnor U48397 (N_48397,N_47851,N_47544);
xor U48398 (N_48398,N_47300,N_47168);
and U48399 (N_48399,N_47496,N_47447);
xor U48400 (N_48400,N_47321,N_47582);
xor U48401 (N_48401,N_47737,N_47791);
xor U48402 (N_48402,N_47662,N_47674);
and U48403 (N_48403,N_47642,N_47554);
nor U48404 (N_48404,N_47599,N_47323);
xor U48405 (N_48405,N_47175,N_47583);
nand U48406 (N_48406,N_47030,N_47618);
and U48407 (N_48407,N_47790,N_47296);
or U48408 (N_48408,N_47473,N_47916);
xnor U48409 (N_48409,N_47096,N_47386);
or U48410 (N_48410,N_47733,N_47663);
nand U48411 (N_48411,N_47050,N_47661);
xor U48412 (N_48412,N_47549,N_47620);
xor U48413 (N_48413,N_47740,N_47888);
or U48414 (N_48414,N_47893,N_47739);
nand U48415 (N_48415,N_47650,N_47657);
nand U48416 (N_48416,N_47398,N_47837);
xnor U48417 (N_48417,N_47060,N_47487);
nor U48418 (N_48418,N_47716,N_47700);
nor U48419 (N_48419,N_47298,N_47373);
or U48420 (N_48420,N_47005,N_47871);
or U48421 (N_48421,N_47685,N_47170);
or U48422 (N_48422,N_47475,N_47078);
nor U48423 (N_48423,N_47284,N_47273);
or U48424 (N_48424,N_47527,N_47164);
xor U48425 (N_48425,N_47515,N_47516);
and U48426 (N_48426,N_47471,N_47376);
nor U48427 (N_48427,N_47264,N_47063);
or U48428 (N_48428,N_47536,N_47109);
and U48429 (N_48429,N_47584,N_47450);
or U48430 (N_48430,N_47157,N_47120);
or U48431 (N_48431,N_47106,N_47057);
nand U48432 (N_48432,N_47363,N_47512);
and U48433 (N_48433,N_47151,N_47744);
nor U48434 (N_48434,N_47415,N_47659);
nor U48435 (N_48435,N_47551,N_47240);
nand U48436 (N_48436,N_47939,N_47035);
and U48437 (N_48437,N_47015,N_47017);
xor U48438 (N_48438,N_47234,N_47071);
or U48439 (N_48439,N_47395,N_47682);
nand U48440 (N_48440,N_47760,N_47521);
or U48441 (N_48441,N_47389,N_47347);
and U48442 (N_48442,N_47152,N_47943);
xnor U48443 (N_48443,N_47868,N_47856);
nor U48444 (N_48444,N_47027,N_47144);
nor U48445 (N_48445,N_47673,N_47336);
or U48446 (N_48446,N_47543,N_47018);
xnor U48447 (N_48447,N_47605,N_47331);
and U48448 (N_48448,N_47493,N_47623);
xnor U48449 (N_48449,N_47639,N_47777);
xnor U48450 (N_48450,N_47820,N_47397);
xor U48451 (N_48451,N_47014,N_47382);
or U48452 (N_48452,N_47245,N_47969);
nor U48453 (N_48453,N_47237,N_47995);
nor U48454 (N_48454,N_47476,N_47950);
and U48455 (N_48455,N_47664,N_47199);
and U48456 (N_48456,N_47192,N_47391);
or U48457 (N_48457,N_47318,N_47869);
nand U48458 (N_48458,N_47561,N_47703);
or U48459 (N_48459,N_47375,N_47756);
nor U48460 (N_48460,N_47125,N_47178);
xor U48461 (N_48461,N_47773,N_47919);
and U48462 (N_48462,N_47085,N_47202);
nor U48463 (N_48463,N_47900,N_47348);
nor U48464 (N_48464,N_47467,N_47956);
or U48465 (N_48465,N_47687,N_47743);
nor U48466 (N_48466,N_47340,N_47585);
or U48467 (N_48467,N_47220,N_47807);
nand U48468 (N_48468,N_47179,N_47224);
nand U48469 (N_48469,N_47204,N_47377);
xor U48470 (N_48470,N_47457,N_47349);
nor U48471 (N_48471,N_47787,N_47978);
xor U48472 (N_48472,N_47619,N_47132);
nor U48473 (N_48473,N_47874,N_47878);
or U48474 (N_48474,N_47288,N_47221);
and U48475 (N_48475,N_47715,N_47854);
nand U48476 (N_48476,N_47468,N_47988);
and U48477 (N_48477,N_47562,N_47070);
and U48478 (N_48478,N_47530,N_47011);
nand U48479 (N_48479,N_47517,N_47013);
and U48480 (N_48480,N_47596,N_47053);
or U48481 (N_48481,N_47761,N_47320);
and U48482 (N_48482,N_47392,N_47250);
nand U48483 (N_48483,N_47127,N_47824);
nor U48484 (N_48484,N_47570,N_47971);
or U48485 (N_48485,N_47730,N_47477);
or U48486 (N_48486,N_47844,N_47370);
xnor U48487 (N_48487,N_47903,N_47104);
nor U48488 (N_48488,N_47873,N_47330);
or U48489 (N_48489,N_47511,N_47155);
nor U48490 (N_48490,N_47904,N_47244);
or U48491 (N_48491,N_47452,N_47963);
nand U48492 (N_48492,N_47560,N_47612);
nand U48493 (N_48493,N_47757,N_47542);
nor U48494 (N_48494,N_47552,N_47881);
and U48495 (N_48495,N_47355,N_47846);
and U48496 (N_48496,N_47821,N_47520);
nand U48497 (N_48497,N_47911,N_47793);
or U48498 (N_48498,N_47110,N_47917);
nand U48499 (N_48499,N_47379,N_47611);
or U48500 (N_48500,N_47914,N_47743);
or U48501 (N_48501,N_47718,N_47753);
and U48502 (N_48502,N_47345,N_47518);
or U48503 (N_48503,N_47666,N_47960);
nand U48504 (N_48504,N_47678,N_47393);
nor U48505 (N_48505,N_47351,N_47435);
xor U48506 (N_48506,N_47458,N_47316);
nor U48507 (N_48507,N_47176,N_47883);
or U48508 (N_48508,N_47891,N_47205);
nor U48509 (N_48509,N_47052,N_47510);
nand U48510 (N_48510,N_47835,N_47473);
nor U48511 (N_48511,N_47411,N_47636);
and U48512 (N_48512,N_47934,N_47570);
nand U48513 (N_48513,N_47998,N_47527);
xnor U48514 (N_48514,N_47163,N_47355);
or U48515 (N_48515,N_47098,N_47380);
or U48516 (N_48516,N_47614,N_47818);
xor U48517 (N_48517,N_47268,N_47930);
and U48518 (N_48518,N_47350,N_47577);
or U48519 (N_48519,N_47391,N_47445);
and U48520 (N_48520,N_47503,N_47110);
xor U48521 (N_48521,N_47153,N_47809);
and U48522 (N_48522,N_47934,N_47087);
and U48523 (N_48523,N_47324,N_47275);
nor U48524 (N_48524,N_47641,N_47030);
or U48525 (N_48525,N_47948,N_47773);
and U48526 (N_48526,N_47581,N_47154);
nand U48527 (N_48527,N_47745,N_47456);
xor U48528 (N_48528,N_47562,N_47065);
or U48529 (N_48529,N_47545,N_47570);
or U48530 (N_48530,N_47355,N_47848);
or U48531 (N_48531,N_47850,N_47326);
or U48532 (N_48532,N_47171,N_47272);
nand U48533 (N_48533,N_47094,N_47273);
nand U48534 (N_48534,N_47530,N_47928);
nand U48535 (N_48535,N_47575,N_47833);
nand U48536 (N_48536,N_47277,N_47158);
xor U48537 (N_48537,N_47260,N_47444);
or U48538 (N_48538,N_47507,N_47233);
and U48539 (N_48539,N_47762,N_47571);
or U48540 (N_48540,N_47357,N_47512);
xnor U48541 (N_48541,N_47718,N_47721);
or U48542 (N_48542,N_47946,N_47871);
xnor U48543 (N_48543,N_47807,N_47678);
or U48544 (N_48544,N_47639,N_47994);
and U48545 (N_48545,N_47169,N_47014);
and U48546 (N_48546,N_47772,N_47679);
nor U48547 (N_48547,N_47262,N_47020);
nor U48548 (N_48548,N_47776,N_47151);
xnor U48549 (N_48549,N_47632,N_47825);
nor U48550 (N_48550,N_47611,N_47262);
nor U48551 (N_48551,N_47898,N_47082);
or U48552 (N_48552,N_47821,N_47350);
nor U48553 (N_48553,N_47660,N_47249);
xor U48554 (N_48554,N_47406,N_47480);
nand U48555 (N_48555,N_47301,N_47119);
xnor U48556 (N_48556,N_47675,N_47639);
and U48557 (N_48557,N_47618,N_47971);
nor U48558 (N_48558,N_47648,N_47261);
and U48559 (N_48559,N_47046,N_47182);
or U48560 (N_48560,N_47384,N_47503);
nor U48561 (N_48561,N_47580,N_47451);
and U48562 (N_48562,N_47237,N_47351);
xnor U48563 (N_48563,N_47484,N_47423);
and U48564 (N_48564,N_47663,N_47023);
xor U48565 (N_48565,N_47548,N_47117);
and U48566 (N_48566,N_47874,N_47197);
nor U48567 (N_48567,N_47525,N_47050);
or U48568 (N_48568,N_47235,N_47222);
and U48569 (N_48569,N_47309,N_47124);
nor U48570 (N_48570,N_47405,N_47728);
or U48571 (N_48571,N_47178,N_47407);
nor U48572 (N_48572,N_47174,N_47611);
or U48573 (N_48573,N_47029,N_47076);
nand U48574 (N_48574,N_47913,N_47688);
or U48575 (N_48575,N_47850,N_47196);
xor U48576 (N_48576,N_47191,N_47440);
xnor U48577 (N_48577,N_47446,N_47013);
xnor U48578 (N_48578,N_47259,N_47006);
xnor U48579 (N_48579,N_47440,N_47419);
nor U48580 (N_48580,N_47849,N_47746);
xor U48581 (N_48581,N_47700,N_47622);
nand U48582 (N_48582,N_47312,N_47775);
nor U48583 (N_48583,N_47329,N_47845);
nor U48584 (N_48584,N_47544,N_47473);
xnor U48585 (N_48585,N_47545,N_47592);
nor U48586 (N_48586,N_47695,N_47841);
nor U48587 (N_48587,N_47457,N_47689);
xor U48588 (N_48588,N_47443,N_47670);
nor U48589 (N_48589,N_47158,N_47878);
nand U48590 (N_48590,N_47803,N_47996);
nand U48591 (N_48591,N_47207,N_47977);
nor U48592 (N_48592,N_47112,N_47698);
xnor U48593 (N_48593,N_47159,N_47377);
nor U48594 (N_48594,N_47327,N_47639);
or U48595 (N_48595,N_47243,N_47127);
nand U48596 (N_48596,N_47700,N_47058);
xor U48597 (N_48597,N_47951,N_47495);
nor U48598 (N_48598,N_47086,N_47287);
or U48599 (N_48599,N_47792,N_47505);
nand U48600 (N_48600,N_47291,N_47429);
nand U48601 (N_48601,N_47650,N_47717);
and U48602 (N_48602,N_47848,N_47436);
and U48603 (N_48603,N_47350,N_47571);
nand U48604 (N_48604,N_47695,N_47789);
nand U48605 (N_48605,N_47727,N_47886);
nand U48606 (N_48606,N_47371,N_47367);
and U48607 (N_48607,N_47012,N_47111);
xnor U48608 (N_48608,N_47631,N_47603);
xnor U48609 (N_48609,N_47070,N_47833);
nand U48610 (N_48610,N_47923,N_47015);
xor U48611 (N_48611,N_47223,N_47318);
nor U48612 (N_48612,N_47367,N_47796);
or U48613 (N_48613,N_47902,N_47580);
nand U48614 (N_48614,N_47309,N_47847);
nor U48615 (N_48615,N_47530,N_47489);
nand U48616 (N_48616,N_47831,N_47234);
nor U48617 (N_48617,N_47965,N_47446);
xnor U48618 (N_48618,N_47902,N_47735);
or U48619 (N_48619,N_47336,N_47637);
and U48620 (N_48620,N_47847,N_47554);
nand U48621 (N_48621,N_47632,N_47901);
or U48622 (N_48622,N_47920,N_47990);
and U48623 (N_48623,N_47401,N_47059);
xor U48624 (N_48624,N_47694,N_47227);
nand U48625 (N_48625,N_47626,N_47848);
nand U48626 (N_48626,N_47302,N_47499);
xnor U48627 (N_48627,N_47134,N_47406);
nand U48628 (N_48628,N_47332,N_47213);
xor U48629 (N_48629,N_47681,N_47653);
or U48630 (N_48630,N_47357,N_47463);
and U48631 (N_48631,N_47702,N_47690);
or U48632 (N_48632,N_47471,N_47624);
nand U48633 (N_48633,N_47154,N_47831);
nand U48634 (N_48634,N_47404,N_47159);
or U48635 (N_48635,N_47390,N_47871);
and U48636 (N_48636,N_47257,N_47549);
nor U48637 (N_48637,N_47486,N_47661);
nor U48638 (N_48638,N_47929,N_47821);
nor U48639 (N_48639,N_47049,N_47952);
nand U48640 (N_48640,N_47051,N_47370);
xnor U48641 (N_48641,N_47928,N_47678);
xnor U48642 (N_48642,N_47335,N_47913);
and U48643 (N_48643,N_47913,N_47377);
or U48644 (N_48644,N_47237,N_47993);
nand U48645 (N_48645,N_47590,N_47179);
or U48646 (N_48646,N_47158,N_47316);
or U48647 (N_48647,N_47550,N_47347);
and U48648 (N_48648,N_47818,N_47976);
or U48649 (N_48649,N_47719,N_47235);
or U48650 (N_48650,N_47052,N_47516);
nor U48651 (N_48651,N_47930,N_47707);
and U48652 (N_48652,N_47582,N_47141);
xnor U48653 (N_48653,N_47047,N_47020);
nand U48654 (N_48654,N_47428,N_47463);
nand U48655 (N_48655,N_47301,N_47133);
nand U48656 (N_48656,N_47514,N_47640);
xnor U48657 (N_48657,N_47455,N_47062);
and U48658 (N_48658,N_47697,N_47111);
nor U48659 (N_48659,N_47036,N_47210);
xor U48660 (N_48660,N_47327,N_47576);
xor U48661 (N_48661,N_47119,N_47344);
or U48662 (N_48662,N_47592,N_47989);
nor U48663 (N_48663,N_47352,N_47987);
and U48664 (N_48664,N_47234,N_47724);
nand U48665 (N_48665,N_47758,N_47278);
and U48666 (N_48666,N_47001,N_47312);
or U48667 (N_48667,N_47443,N_47128);
nand U48668 (N_48668,N_47937,N_47815);
nor U48669 (N_48669,N_47302,N_47185);
nor U48670 (N_48670,N_47994,N_47093);
or U48671 (N_48671,N_47320,N_47702);
and U48672 (N_48672,N_47799,N_47953);
and U48673 (N_48673,N_47930,N_47419);
nor U48674 (N_48674,N_47523,N_47656);
xnor U48675 (N_48675,N_47901,N_47820);
and U48676 (N_48676,N_47125,N_47923);
and U48677 (N_48677,N_47245,N_47273);
xnor U48678 (N_48678,N_47504,N_47441);
or U48679 (N_48679,N_47079,N_47790);
xor U48680 (N_48680,N_47636,N_47435);
nor U48681 (N_48681,N_47056,N_47486);
or U48682 (N_48682,N_47942,N_47316);
nand U48683 (N_48683,N_47754,N_47039);
or U48684 (N_48684,N_47039,N_47290);
nand U48685 (N_48685,N_47421,N_47368);
xor U48686 (N_48686,N_47371,N_47783);
xor U48687 (N_48687,N_47595,N_47694);
nand U48688 (N_48688,N_47795,N_47043);
or U48689 (N_48689,N_47856,N_47150);
nand U48690 (N_48690,N_47852,N_47805);
or U48691 (N_48691,N_47199,N_47261);
and U48692 (N_48692,N_47067,N_47729);
nor U48693 (N_48693,N_47147,N_47911);
and U48694 (N_48694,N_47693,N_47654);
or U48695 (N_48695,N_47853,N_47344);
nand U48696 (N_48696,N_47431,N_47630);
and U48697 (N_48697,N_47301,N_47031);
and U48698 (N_48698,N_47067,N_47221);
xor U48699 (N_48699,N_47629,N_47216);
nand U48700 (N_48700,N_47727,N_47883);
nand U48701 (N_48701,N_47014,N_47271);
xor U48702 (N_48702,N_47168,N_47431);
nand U48703 (N_48703,N_47419,N_47037);
or U48704 (N_48704,N_47488,N_47899);
or U48705 (N_48705,N_47090,N_47501);
xnor U48706 (N_48706,N_47688,N_47968);
nor U48707 (N_48707,N_47594,N_47513);
and U48708 (N_48708,N_47057,N_47584);
or U48709 (N_48709,N_47479,N_47714);
or U48710 (N_48710,N_47650,N_47442);
nand U48711 (N_48711,N_47057,N_47210);
nor U48712 (N_48712,N_47347,N_47485);
or U48713 (N_48713,N_47116,N_47068);
nand U48714 (N_48714,N_47339,N_47712);
and U48715 (N_48715,N_47033,N_47079);
nor U48716 (N_48716,N_47855,N_47672);
xnor U48717 (N_48717,N_47602,N_47655);
and U48718 (N_48718,N_47997,N_47192);
xor U48719 (N_48719,N_47559,N_47539);
nand U48720 (N_48720,N_47678,N_47933);
and U48721 (N_48721,N_47018,N_47562);
nor U48722 (N_48722,N_47965,N_47052);
nand U48723 (N_48723,N_47518,N_47218);
nand U48724 (N_48724,N_47909,N_47219);
and U48725 (N_48725,N_47175,N_47613);
nand U48726 (N_48726,N_47082,N_47500);
or U48727 (N_48727,N_47560,N_47509);
and U48728 (N_48728,N_47469,N_47216);
and U48729 (N_48729,N_47852,N_47677);
and U48730 (N_48730,N_47949,N_47198);
or U48731 (N_48731,N_47324,N_47805);
and U48732 (N_48732,N_47055,N_47236);
nor U48733 (N_48733,N_47216,N_47354);
nor U48734 (N_48734,N_47608,N_47154);
or U48735 (N_48735,N_47069,N_47019);
or U48736 (N_48736,N_47141,N_47012);
nor U48737 (N_48737,N_47674,N_47494);
nand U48738 (N_48738,N_47408,N_47024);
nand U48739 (N_48739,N_47563,N_47497);
and U48740 (N_48740,N_47929,N_47749);
or U48741 (N_48741,N_47345,N_47379);
and U48742 (N_48742,N_47598,N_47676);
or U48743 (N_48743,N_47422,N_47922);
nand U48744 (N_48744,N_47113,N_47938);
nor U48745 (N_48745,N_47203,N_47638);
xnor U48746 (N_48746,N_47233,N_47661);
xnor U48747 (N_48747,N_47453,N_47249);
nand U48748 (N_48748,N_47245,N_47297);
nand U48749 (N_48749,N_47144,N_47383);
nor U48750 (N_48750,N_47836,N_47768);
and U48751 (N_48751,N_47867,N_47537);
nor U48752 (N_48752,N_47051,N_47963);
and U48753 (N_48753,N_47821,N_47630);
xor U48754 (N_48754,N_47643,N_47784);
or U48755 (N_48755,N_47208,N_47212);
nor U48756 (N_48756,N_47438,N_47953);
or U48757 (N_48757,N_47246,N_47156);
and U48758 (N_48758,N_47670,N_47522);
nand U48759 (N_48759,N_47858,N_47751);
xnor U48760 (N_48760,N_47754,N_47834);
or U48761 (N_48761,N_47732,N_47141);
and U48762 (N_48762,N_47480,N_47872);
or U48763 (N_48763,N_47470,N_47149);
and U48764 (N_48764,N_47575,N_47433);
xnor U48765 (N_48765,N_47333,N_47589);
or U48766 (N_48766,N_47130,N_47916);
or U48767 (N_48767,N_47071,N_47177);
nand U48768 (N_48768,N_47721,N_47315);
or U48769 (N_48769,N_47876,N_47963);
nand U48770 (N_48770,N_47485,N_47647);
or U48771 (N_48771,N_47121,N_47093);
nand U48772 (N_48772,N_47236,N_47794);
or U48773 (N_48773,N_47785,N_47113);
or U48774 (N_48774,N_47328,N_47412);
xnor U48775 (N_48775,N_47386,N_47020);
and U48776 (N_48776,N_47743,N_47078);
nand U48777 (N_48777,N_47889,N_47173);
and U48778 (N_48778,N_47778,N_47259);
and U48779 (N_48779,N_47055,N_47931);
nor U48780 (N_48780,N_47699,N_47639);
and U48781 (N_48781,N_47701,N_47919);
xor U48782 (N_48782,N_47313,N_47251);
nand U48783 (N_48783,N_47779,N_47778);
nand U48784 (N_48784,N_47648,N_47751);
and U48785 (N_48785,N_47397,N_47480);
and U48786 (N_48786,N_47064,N_47010);
nor U48787 (N_48787,N_47084,N_47881);
nor U48788 (N_48788,N_47865,N_47419);
nor U48789 (N_48789,N_47006,N_47669);
and U48790 (N_48790,N_47798,N_47784);
or U48791 (N_48791,N_47210,N_47230);
or U48792 (N_48792,N_47380,N_47726);
nand U48793 (N_48793,N_47587,N_47085);
nand U48794 (N_48794,N_47183,N_47755);
nand U48795 (N_48795,N_47133,N_47048);
xor U48796 (N_48796,N_47849,N_47022);
nand U48797 (N_48797,N_47011,N_47402);
or U48798 (N_48798,N_47379,N_47707);
and U48799 (N_48799,N_47397,N_47425);
nand U48800 (N_48800,N_47772,N_47165);
nand U48801 (N_48801,N_47284,N_47047);
or U48802 (N_48802,N_47231,N_47267);
nor U48803 (N_48803,N_47626,N_47228);
nand U48804 (N_48804,N_47619,N_47690);
and U48805 (N_48805,N_47649,N_47455);
nand U48806 (N_48806,N_47765,N_47092);
nor U48807 (N_48807,N_47611,N_47920);
or U48808 (N_48808,N_47179,N_47757);
xnor U48809 (N_48809,N_47265,N_47405);
and U48810 (N_48810,N_47902,N_47282);
nand U48811 (N_48811,N_47205,N_47908);
nor U48812 (N_48812,N_47082,N_47484);
xor U48813 (N_48813,N_47800,N_47311);
and U48814 (N_48814,N_47208,N_47441);
nand U48815 (N_48815,N_47586,N_47332);
and U48816 (N_48816,N_47608,N_47411);
nor U48817 (N_48817,N_47436,N_47267);
and U48818 (N_48818,N_47290,N_47122);
nand U48819 (N_48819,N_47701,N_47301);
nand U48820 (N_48820,N_47113,N_47490);
xor U48821 (N_48821,N_47221,N_47834);
and U48822 (N_48822,N_47040,N_47688);
xnor U48823 (N_48823,N_47549,N_47693);
xor U48824 (N_48824,N_47724,N_47040);
nor U48825 (N_48825,N_47445,N_47273);
or U48826 (N_48826,N_47866,N_47475);
xnor U48827 (N_48827,N_47301,N_47860);
and U48828 (N_48828,N_47916,N_47406);
nand U48829 (N_48829,N_47232,N_47591);
xor U48830 (N_48830,N_47525,N_47311);
nor U48831 (N_48831,N_47266,N_47209);
nor U48832 (N_48832,N_47963,N_47955);
nand U48833 (N_48833,N_47513,N_47020);
xor U48834 (N_48834,N_47473,N_47927);
nand U48835 (N_48835,N_47720,N_47071);
nor U48836 (N_48836,N_47049,N_47158);
and U48837 (N_48837,N_47543,N_47053);
nand U48838 (N_48838,N_47639,N_47199);
or U48839 (N_48839,N_47210,N_47794);
nand U48840 (N_48840,N_47552,N_47446);
or U48841 (N_48841,N_47867,N_47590);
or U48842 (N_48842,N_47697,N_47789);
and U48843 (N_48843,N_47103,N_47449);
or U48844 (N_48844,N_47139,N_47597);
and U48845 (N_48845,N_47991,N_47339);
xnor U48846 (N_48846,N_47560,N_47177);
or U48847 (N_48847,N_47775,N_47680);
nor U48848 (N_48848,N_47548,N_47211);
nand U48849 (N_48849,N_47215,N_47050);
and U48850 (N_48850,N_47801,N_47340);
xnor U48851 (N_48851,N_47133,N_47739);
and U48852 (N_48852,N_47698,N_47822);
xnor U48853 (N_48853,N_47079,N_47626);
and U48854 (N_48854,N_47145,N_47884);
or U48855 (N_48855,N_47466,N_47674);
xnor U48856 (N_48856,N_47372,N_47905);
and U48857 (N_48857,N_47803,N_47820);
or U48858 (N_48858,N_47095,N_47059);
and U48859 (N_48859,N_47663,N_47922);
xnor U48860 (N_48860,N_47806,N_47641);
nand U48861 (N_48861,N_47574,N_47234);
nor U48862 (N_48862,N_47958,N_47755);
nand U48863 (N_48863,N_47727,N_47052);
xnor U48864 (N_48864,N_47742,N_47086);
and U48865 (N_48865,N_47334,N_47418);
nor U48866 (N_48866,N_47747,N_47403);
xor U48867 (N_48867,N_47856,N_47852);
nor U48868 (N_48868,N_47071,N_47296);
and U48869 (N_48869,N_47899,N_47486);
or U48870 (N_48870,N_47698,N_47503);
nand U48871 (N_48871,N_47990,N_47461);
and U48872 (N_48872,N_47712,N_47052);
nand U48873 (N_48873,N_47337,N_47348);
xnor U48874 (N_48874,N_47280,N_47725);
nand U48875 (N_48875,N_47187,N_47329);
nand U48876 (N_48876,N_47149,N_47576);
and U48877 (N_48877,N_47552,N_47958);
xor U48878 (N_48878,N_47832,N_47662);
nand U48879 (N_48879,N_47546,N_47624);
and U48880 (N_48880,N_47071,N_47059);
nor U48881 (N_48881,N_47982,N_47892);
nand U48882 (N_48882,N_47300,N_47022);
and U48883 (N_48883,N_47902,N_47896);
xnor U48884 (N_48884,N_47388,N_47943);
or U48885 (N_48885,N_47110,N_47136);
nor U48886 (N_48886,N_47650,N_47794);
xnor U48887 (N_48887,N_47732,N_47299);
xnor U48888 (N_48888,N_47082,N_47900);
xnor U48889 (N_48889,N_47232,N_47354);
nor U48890 (N_48890,N_47836,N_47032);
or U48891 (N_48891,N_47944,N_47253);
or U48892 (N_48892,N_47610,N_47466);
nand U48893 (N_48893,N_47447,N_47561);
xnor U48894 (N_48894,N_47133,N_47297);
or U48895 (N_48895,N_47995,N_47103);
nand U48896 (N_48896,N_47214,N_47654);
nand U48897 (N_48897,N_47623,N_47341);
nand U48898 (N_48898,N_47414,N_47397);
nand U48899 (N_48899,N_47241,N_47841);
and U48900 (N_48900,N_47962,N_47199);
and U48901 (N_48901,N_47385,N_47733);
xnor U48902 (N_48902,N_47776,N_47235);
nor U48903 (N_48903,N_47216,N_47257);
nor U48904 (N_48904,N_47894,N_47542);
xor U48905 (N_48905,N_47889,N_47586);
nand U48906 (N_48906,N_47762,N_47921);
xor U48907 (N_48907,N_47199,N_47280);
nor U48908 (N_48908,N_47748,N_47404);
xnor U48909 (N_48909,N_47438,N_47048);
nand U48910 (N_48910,N_47389,N_47485);
and U48911 (N_48911,N_47931,N_47050);
xnor U48912 (N_48912,N_47872,N_47924);
or U48913 (N_48913,N_47714,N_47524);
nand U48914 (N_48914,N_47786,N_47918);
or U48915 (N_48915,N_47014,N_47547);
and U48916 (N_48916,N_47960,N_47748);
and U48917 (N_48917,N_47752,N_47812);
or U48918 (N_48918,N_47041,N_47129);
nor U48919 (N_48919,N_47927,N_47514);
or U48920 (N_48920,N_47277,N_47670);
nor U48921 (N_48921,N_47629,N_47889);
or U48922 (N_48922,N_47408,N_47190);
xor U48923 (N_48923,N_47800,N_47013);
nand U48924 (N_48924,N_47254,N_47090);
nand U48925 (N_48925,N_47798,N_47376);
nand U48926 (N_48926,N_47203,N_47195);
nand U48927 (N_48927,N_47561,N_47380);
xnor U48928 (N_48928,N_47428,N_47289);
nand U48929 (N_48929,N_47599,N_47548);
nand U48930 (N_48930,N_47749,N_47145);
or U48931 (N_48931,N_47840,N_47602);
and U48932 (N_48932,N_47524,N_47572);
nor U48933 (N_48933,N_47716,N_47513);
xor U48934 (N_48934,N_47250,N_47690);
or U48935 (N_48935,N_47512,N_47881);
or U48936 (N_48936,N_47723,N_47469);
nor U48937 (N_48937,N_47187,N_47966);
nor U48938 (N_48938,N_47015,N_47347);
xnor U48939 (N_48939,N_47249,N_47385);
nand U48940 (N_48940,N_47848,N_47314);
or U48941 (N_48941,N_47195,N_47838);
xor U48942 (N_48942,N_47239,N_47330);
nand U48943 (N_48943,N_47955,N_47477);
xnor U48944 (N_48944,N_47576,N_47975);
nor U48945 (N_48945,N_47024,N_47824);
nand U48946 (N_48946,N_47138,N_47797);
and U48947 (N_48947,N_47644,N_47699);
or U48948 (N_48948,N_47779,N_47638);
or U48949 (N_48949,N_47072,N_47574);
xor U48950 (N_48950,N_47107,N_47229);
nand U48951 (N_48951,N_47884,N_47292);
xnor U48952 (N_48952,N_47114,N_47506);
xor U48953 (N_48953,N_47262,N_47720);
nor U48954 (N_48954,N_47328,N_47022);
and U48955 (N_48955,N_47636,N_47684);
xnor U48956 (N_48956,N_47966,N_47542);
or U48957 (N_48957,N_47595,N_47843);
and U48958 (N_48958,N_47126,N_47218);
or U48959 (N_48959,N_47783,N_47119);
nand U48960 (N_48960,N_47528,N_47080);
or U48961 (N_48961,N_47168,N_47554);
xnor U48962 (N_48962,N_47863,N_47308);
xor U48963 (N_48963,N_47896,N_47336);
or U48964 (N_48964,N_47669,N_47870);
xnor U48965 (N_48965,N_47861,N_47459);
nand U48966 (N_48966,N_47477,N_47209);
xnor U48967 (N_48967,N_47520,N_47665);
nand U48968 (N_48968,N_47823,N_47872);
nor U48969 (N_48969,N_47098,N_47330);
xor U48970 (N_48970,N_47058,N_47359);
or U48971 (N_48971,N_47172,N_47738);
xor U48972 (N_48972,N_47543,N_47314);
nand U48973 (N_48973,N_47250,N_47861);
nor U48974 (N_48974,N_47383,N_47925);
xor U48975 (N_48975,N_47786,N_47077);
nor U48976 (N_48976,N_47504,N_47778);
nand U48977 (N_48977,N_47658,N_47995);
nor U48978 (N_48978,N_47418,N_47890);
xnor U48979 (N_48979,N_47919,N_47534);
or U48980 (N_48980,N_47447,N_47159);
and U48981 (N_48981,N_47698,N_47033);
nor U48982 (N_48982,N_47855,N_47519);
and U48983 (N_48983,N_47886,N_47823);
xor U48984 (N_48984,N_47325,N_47052);
xor U48985 (N_48985,N_47617,N_47248);
or U48986 (N_48986,N_47596,N_47892);
or U48987 (N_48987,N_47165,N_47832);
nor U48988 (N_48988,N_47977,N_47128);
xor U48989 (N_48989,N_47024,N_47324);
nand U48990 (N_48990,N_47287,N_47921);
nor U48991 (N_48991,N_47123,N_47650);
nor U48992 (N_48992,N_47778,N_47172);
xor U48993 (N_48993,N_47618,N_47388);
or U48994 (N_48994,N_47939,N_47777);
or U48995 (N_48995,N_47247,N_47612);
nor U48996 (N_48996,N_47815,N_47203);
nand U48997 (N_48997,N_47754,N_47523);
and U48998 (N_48998,N_47398,N_47812);
xor U48999 (N_48999,N_47882,N_47888);
nor U49000 (N_49000,N_48586,N_48677);
xnor U49001 (N_49001,N_48002,N_48502);
or U49002 (N_49002,N_48132,N_48791);
xor U49003 (N_49003,N_48826,N_48560);
nor U49004 (N_49004,N_48497,N_48816);
xnor U49005 (N_49005,N_48371,N_48590);
or U49006 (N_49006,N_48163,N_48680);
and U49007 (N_49007,N_48164,N_48891);
xnor U49008 (N_49008,N_48366,N_48285);
or U49009 (N_49009,N_48123,N_48667);
and U49010 (N_49010,N_48741,N_48582);
xor U49011 (N_49011,N_48662,N_48925);
and U49012 (N_49012,N_48038,N_48670);
nor U49013 (N_49013,N_48444,N_48706);
xor U49014 (N_49014,N_48997,N_48980);
or U49015 (N_49015,N_48551,N_48776);
or U49016 (N_49016,N_48740,N_48341);
nor U49017 (N_49017,N_48514,N_48346);
nand U49018 (N_49018,N_48759,N_48490);
or U49019 (N_49019,N_48620,N_48781);
or U49020 (N_49020,N_48108,N_48778);
or U49021 (N_49021,N_48295,N_48086);
and U49022 (N_49022,N_48865,N_48562);
nor U49023 (N_49023,N_48316,N_48446);
nor U49024 (N_49024,N_48090,N_48202);
nand U49025 (N_49025,N_48313,N_48613);
and U49026 (N_49026,N_48375,N_48096);
nor U49027 (N_49027,N_48656,N_48325);
nand U49028 (N_49028,N_48665,N_48068);
xor U49029 (N_49029,N_48278,N_48328);
and U49030 (N_49030,N_48718,N_48138);
xnor U49031 (N_49031,N_48238,N_48940);
and U49032 (N_49032,N_48290,N_48877);
nor U49033 (N_49033,N_48728,N_48570);
xnor U49034 (N_49034,N_48326,N_48367);
or U49035 (N_49035,N_48257,N_48355);
or U49036 (N_49036,N_48655,N_48763);
nor U49037 (N_49037,N_48957,N_48974);
xnor U49038 (N_49038,N_48427,N_48978);
nor U49039 (N_49039,N_48401,N_48822);
xnor U49040 (N_49040,N_48516,N_48528);
nand U49041 (N_49041,N_48890,N_48755);
and U49042 (N_49042,N_48291,N_48731);
or U49043 (N_49043,N_48557,N_48664);
nand U49044 (N_49044,N_48000,N_48585);
and U49045 (N_49045,N_48395,N_48615);
nand U49046 (N_49046,N_48266,N_48927);
or U49047 (N_49047,N_48463,N_48150);
and U49048 (N_49048,N_48621,N_48833);
nor U49049 (N_49049,N_48683,N_48811);
and U49050 (N_49050,N_48530,N_48142);
nand U49051 (N_49051,N_48919,N_48795);
and U49052 (N_49052,N_48074,N_48765);
or U49053 (N_49053,N_48353,N_48310);
xor U49054 (N_49054,N_48565,N_48722);
xor U49055 (N_49055,N_48394,N_48179);
nand U49056 (N_49056,N_48724,N_48913);
nand U49057 (N_49057,N_48466,N_48209);
xnor U49058 (N_49058,N_48248,N_48568);
nor U49059 (N_49059,N_48292,N_48631);
xnor U49060 (N_49060,N_48846,N_48647);
and U49061 (N_49061,N_48600,N_48478);
xor U49062 (N_49062,N_48536,N_48032);
and U49063 (N_49063,N_48605,N_48013);
or U49064 (N_49064,N_48732,N_48253);
nor U49065 (N_49065,N_48835,N_48194);
or U49066 (N_49066,N_48244,N_48533);
or U49067 (N_49067,N_48124,N_48028);
xnor U49068 (N_49068,N_48691,N_48524);
and U49069 (N_49069,N_48085,N_48409);
xnor U49070 (N_49070,N_48232,N_48803);
xor U49071 (N_49071,N_48230,N_48505);
and U49072 (N_49072,N_48552,N_48734);
xnor U49073 (N_49073,N_48465,N_48162);
and U49074 (N_49074,N_48348,N_48785);
nor U49075 (N_49075,N_48224,N_48976);
nor U49076 (N_49076,N_48218,N_48454);
xor U49077 (N_49077,N_48007,N_48538);
nor U49078 (N_49078,N_48602,N_48991);
and U49079 (N_49079,N_48284,N_48076);
nand U49080 (N_49080,N_48930,N_48668);
nand U49081 (N_49081,N_48693,N_48413);
nand U49082 (N_49082,N_48223,N_48420);
and U49083 (N_49083,N_48301,N_48770);
nand U49084 (N_49084,N_48589,N_48334);
nand U49085 (N_49085,N_48182,N_48486);
nor U49086 (N_49086,N_48629,N_48003);
xnor U49087 (N_49087,N_48167,N_48452);
and U49088 (N_49088,N_48540,N_48064);
nor U49089 (N_49089,N_48844,N_48738);
nor U49090 (N_49090,N_48424,N_48384);
nand U49091 (N_49091,N_48060,N_48210);
or U49092 (N_49092,N_48416,N_48566);
nand U49093 (N_49093,N_48773,N_48669);
and U49094 (N_49094,N_48513,N_48944);
and U49095 (N_49095,N_48801,N_48360);
nor U49096 (N_49096,N_48131,N_48018);
xnor U49097 (N_49097,N_48507,N_48347);
nand U49098 (N_49098,N_48004,N_48012);
and U49099 (N_49099,N_48775,N_48322);
and U49100 (N_49100,N_48483,N_48817);
nand U49101 (N_49101,N_48658,N_48898);
xnor U49102 (N_49102,N_48343,N_48922);
nand U49103 (N_49103,N_48958,N_48931);
nand U49104 (N_49104,N_48027,N_48461);
nand U49105 (N_49105,N_48354,N_48226);
or U49106 (N_49106,N_48023,N_48410);
nand U49107 (N_49107,N_48742,N_48153);
nand U49108 (N_49108,N_48572,N_48415);
and U49109 (N_49109,N_48399,N_48261);
or U49110 (N_49110,N_48779,N_48159);
and U49111 (N_49111,N_48084,N_48286);
nor U49112 (N_49112,N_48289,N_48640);
or U49113 (N_49113,N_48964,N_48333);
xnor U49114 (N_49114,N_48687,N_48445);
or U49115 (N_49115,N_48715,N_48554);
or U49116 (N_49116,N_48067,N_48556);
xor U49117 (N_49117,N_48821,N_48148);
nand U49118 (N_49118,N_48357,N_48034);
and U49119 (N_49119,N_48686,N_48908);
and U49120 (N_49120,N_48379,N_48033);
xnor U49121 (N_49121,N_48121,N_48361);
and U49122 (N_49122,N_48406,N_48120);
and U49123 (N_49123,N_48443,N_48152);
or U49124 (N_49124,N_48845,N_48783);
nand U49125 (N_49125,N_48708,N_48442);
nand U49126 (N_49126,N_48104,N_48905);
nand U49127 (N_49127,N_48247,N_48176);
or U49128 (N_49128,N_48797,N_48648);
xor U49129 (N_49129,N_48470,N_48591);
nor U49130 (N_49130,N_48933,N_48055);
nor U49131 (N_49131,N_48282,N_48240);
xnor U49132 (N_49132,N_48476,N_48598);
and U49133 (N_49133,N_48082,N_48970);
xnor U49134 (N_49134,N_48807,N_48579);
nor U49135 (N_49135,N_48369,N_48508);
nor U49136 (N_49136,N_48576,N_48187);
nor U49137 (N_49137,N_48504,N_48679);
nor U49138 (N_49138,N_48725,N_48491);
nand U49139 (N_49139,N_48723,N_48743);
nand U49140 (N_49140,N_48362,N_48876);
xor U49141 (N_49141,N_48831,N_48875);
xor U49142 (N_49142,N_48872,N_48986);
and U49143 (N_49143,N_48965,N_48998);
nand U49144 (N_49144,N_48727,N_48269);
nor U49145 (N_49145,N_48404,N_48382);
or U49146 (N_49146,N_48800,N_48711);
nor U49147 (N_49147,N_48365,N_48915);
and U49148 (N_49148,N_48246,N_48947);
nand U49149 (N_49149,N_48690,N_48094);
nor U49150 (N_49150,N_48042,N_48414);
or U49151 (N_49151,N_48848,N_48421);
or U49152 (N_49152,N_48016,N_48926);
nor U49153 (N_49153,N_48544,N_48169);
xor U49154 (N_49154,N_48106,N_48307);
nor U49155 (N_49155,N_48713,N_48485);
and U49156 (N_49156,N_48144,N_48573);
xnor U49157 (N_49157,N_48623,N_48627);
xor U49158 (N_49158,N_48049,N_48903);
and U49159 (N_49159,N_48390,N_48233);
and U49160 (N_49160,N_48345,N_48128);
and U49161 (N_49161,N_48275,N_48789);
xor U49162 (N_49162,N_48564,N_48212);
nand U49163 (N_49163,N_48638,N_48329);
and U49164 (N_49164,N_48274,N_48987);
and U49165 (N_49165,N_48071,N_48061);
or U49166 (N_49166,N_48837,N_48858);
or U49167 (N_49167,N_48617,N_48059);
or U49168 (N_49168,N_48867,N_48852);
or U49169 (N_49169,N_48735,N_48087);
xnor U49170 (N_49170,N_48660,N_48139);
or U49171 (N_49171,N_48961,N_48215);
and U49172 (N_49172,N_48948,N_48651);
and U49173 (N_49173,N_48432,N_48237);
or U49174 (N_49174,N_48784,N_48529);
nand U49175 (N_49175,N_48035,N_48319);
nor U49176 (N_49176,N_48095,N_48641);
xor U49177 (N_49177,N_48851,N_48906);
nor U49178 (N_49178,N_48161,N_48818);
xnor U49179 (N_49179,N_48479,N_48721);
nand U49180 (N_49180,N_48625,N_48039);
nand U49181 (N_49181,N_48356,N_48654);
nor U49182 (N_49182,N_48306,N_48971);
or U49183 (N_49183,N_48263,N_48389);
nor U49184 (N_49184,N_48079,N_48093);
or U49185 (N_49185,N_48841,N_48659);
xnor U49186 (N_49186,N_48772,N_48788);
nor U49187 (N_49187,N_48058,N_48798);
nand U49188 (N_49188,N_48193,N_48955);
and U49189 (N_49189,N_48663,N_48635);
xor U49190 (N_49190,N_48911,N_48448);
or U49191 (N_49191,N_48241,N_48642);
nor U49192 (N_49192,N_48422,N_48920);
xor U49193 (N_49193,N_48607,N_48293);
and U49194 (N_49194,N_48736,N_48489);
xnor U49195 (N_49195,N_48984,N_48323);
and U49196 (N_49196,N_48227,N_48403);
and U49197 (N_49197,N_48030,N_48517);
or U49198 (N_49198,N_48595,N_48726);
nand U49199 (N_49199,N_48695,N_48934);
nand U49200 (N_49200,N_48762,N_48337);
and U49201 (N_49201,N_48151,N_48633);
xor U49202 (N_49202,N_48063,N_48515);
nor U49203 (N_49203,N_48252,N_48692);
and U49204 (N_49204,N_48904,N_48973);
xor U49205 (N_49205,N_48468,N_48653);
xor U49206 (N_49206,N_48405,N_48769);
nand U49207 (N_49207,N_48205,N_48214);
nand U49208 (N_49208,N_48168,N_48231);
nand U49209 (N_49209,N_48879,N_48137);
or U49210 (N_49210,N_48283,N_48939);
nor U49211 (N_49211,N_48666,N_48057);
or U49212 (N_49212,N_48558,N_48459);
and U49213 (N_49213,N_48234,N_48819);
xnor U49214 (N_49214,N_48972,N_48281);
nor U49215 (N_49215,N_48411,N_48881);
nand U49216 (N_49216,N_48160,N_48916);
or U49217 (N_49217,N_48645,N_48989);
or U49218 (N_49218,N_48914,N_48114);
xnor U49219 (N_49219,N_48982,N_48618);
nand U49220 (N_49220,N_48488,N_48988);
or U49221 (N_49221,N_48288,N_48439);
xor U49222 (N_49222,N_48813,N_48184);
or U49223 (N_49223,N_48510,N_48859);
and U49224 (N_49224,N_48563,N_48196);
or U49225 (N_49225,N_48588,N_48207);
or U49226 (N_49226,N_48219,N_48650);
and U49227 (N_49227,N_48496,N_48847);
nor U49228 (N_49228,N_48436,N_48861);
or U49229 (N_49229,N_48764,N_48857);
nand U49230 (N_49230,N_48447,N_48815);
nand U49231 (N_49231,N_48780,N_48799);
nor U49232 (N_49232,N_48043,N_48894);
xor U49233 (N_49233,N_48189,N_48689);
nand U49234 (N_49234,N_48630,N_48419);
xnor U49235 (N_49235,N_48412,N_48499);
xnor U49236 (N_49236,N_48363,N_48046);
nand U49237 (N_49237,N_48705,N_48135);
xnor U49238 (N_49238,N_48019,N_48298);
nand U49239 (N_49239,N_48751,N_48907);
and U49240 (N_49240,N_48397,N_48349);
or U49241 (N_49241,N_48830,N_48155);
xor U49242 (N_49242,N_48036,N_48197);
and U49243 (N_49243,N_48370,N_48228);
or U49244 (N_49244,N_48754,N_48386);
or U49245 (N_49245,N_48601,N_48391);
or U49246 (N_49246,N_48047,N_48099);
and U49247 (N_49247,N_48103,N_48336);
xor U49248 (N_49248,N_48080,N_48398);
xnor U49249 (N_49249,N_48923,N_48512);
xnor U49250 (N_49250,N_48758,N_48511);
or U49251 (N_49251,N_48332,N_48315);
or U49252 (N_49252,N_48632,N_48069);
and U49253 (N_49253,N_48949,N_48456);
nor U49254 (N_49254,N_48477,N_48198);
nand U49255 (N_49255,N_48450,N_48277);
nor U49256 (N_49256,N_48802,N_48025);
xor U49257 (N_49257,N_48746,N_48578);
nor U49258 (N_49258,N_48899,N_48766);
nand U49259 (N_49259,N_48981,N_48242);
xor U49260 (N_49260,N_48583,N_48183);
or U49261 (N_49261,N_48863,N_48475);
nand U49262 (N_49262,N_48714,N_48717);
or U49263 (N_49263,N_48481,N_48967);
and U49264 (N_49264,N_48378,N_48111);
nand U49265 (N_49265,N_48434,N_48075);
nor U49266 (N_49266,N_48239,N_48344);
nor U49267 (N_49267,N_48786,N_48311);
xor U49268 (N_49268,N_48873,N_48200);
or U49269 (N_49269,N_48140,N_48745);
xnor U49270 (N_49270,N_48271,N_48339);
nor U49271 (N_49271,N_48954,N_48935);
or U49272 (N_49272,N_48593,N_48195);
or U49273 (N_49273,N_48340,N_48685);
nor U49274 (N_49274,N_48272,N_48628);
xnor U49275 (N_49275,N_48880,N_48300);
and U49276 (N_49276,N_48804,N_48190);
and U49277 (N_49277,N_48172,N_48888);
or U49278 (N_49278,N_48719,N_48053);
nand U49279 (N_49279,N_48545,N_48960);
xor U49280 (N_49280,N_48338,N_48015);
nand U49281 (N_49281,N_48221,N_48500);
nand U49282 (N_49282,N_48464,N_48608);
nor U49283 (N_49283,N_48887,N_48938);
or U49284 (N_49284,N_48644,N_48321);
nand U49285 (N_49285,N_48175,N_48119);
nor U49286 (N_49286,N_48828,N_48309);
and U49287 (N_49287,N_48387,N_48276);
xnor U49288 (N_49288,N_48441,N_48267);
and U49289 (N_49289,N_48682,N_48614);
or U49290 (N_49290,N_48279,N_48433);
nand U49291 (N_49291,N_48066,N_48985);
and U49292 (N_49292,N_48860,N_48943);
or U49293 (N_49293,N_48048,N_48701);
and U49294 (N_49294,N_48637,N_48426);
xor U49295 (N_49295,N_48118,N_48050);
or U49296 (N_49296,N_48594,N_48710);
xnor U49297 (N_49297,N_48474,N_48553);
and U49298 (N_49298,N_48744,N_48052);
or U49299 (N_49299,N_48262,N_48806);
nor U49300 (N_49300,N_48428,N_48525);
nand U49301 (N_49301,N_48408,N_48400);
or U49302 (N_49302,N_48969,N_48993);
or U49303 (N_49303,N_48924,N_48134);
xor U49304 (N_49304,N_48372,N_48056);
xnor U49305 (N_49305,N_48051,N_48849);
or U49306 (N_49306,N_48342,N_48145);
or U49307 (N_49307,N_48122,N_48739);
or U49308 (N_49308,N_48287,N_48882);
nor U49309 (N_49309,N_48449,N_48519);
xor U49310 (N_49310,N_48136,N_48983);
nor U49311 (N_49311,N_48199,N_48143);
xor U49312 (N_49312,N_48294,N_48975);
nand U49313 (N_49313,N_48805,N_48302);
and U49314 (N_49314,N_48681,N_48259);
nor U49315 (N_49315,N_48078,N_48657);
xor U49316 (N_49316,N_48577,N_48917);
xor U49317 (N_49317,N_48531,N_48225);
nand U49318 (N_49318,N_48928,N_48661);
xor U49319 (N_49319,N_48639,N_48678);
and U49320 (N_49320,N_48381,N_48767);
or U49321 (N_49321,N_48634,N_48280);
nand U49322 (N_49322,N_48855,N_48995);
xor U49323 (N_49323,N_48469,N_48707);
xor U49324 (N_49324,N_48895,N_48181);
and U49325 (N_49325,N_48921,N_48675);
or U49326 (N_49326,N_48597,N_48709);
and U49327 (N_49327,N_48435,N_48102);
nand U49328 (N_49328,N_48953,N_48203);
and U49329 (N_49329,N_48768,N_48037);
xor U49330 (N_49330,N_48946,N_48070);
and U49331 (N_49331,N_48487,N_48902);
xnor U49332 (N_49332,N_48856,N_48116);
or U49333 (N_49333,N_48024,N_48008);
or U49334 (N_49334,N_48388,N_48684);
nor U49335 (N_49335,N_48918,N_48473);
xnor U49336 (N_49336,N_48838,N_48112);
nand U49337 (N_49337,N_48010,N_48810);
and U49338 (N_49338,N_48793,N_48110);
or U49339 (N_49339,N_48945,N_48229);
nand U49340 (N_49340,N_48383,N_48546);
nand U49341 (N_49341,N_48757,N_48157);
nor U49342 (N_49342,N_48866,N_48368);
xnor U49343 (N_49343,N_48178,N_48149);
or U49344 (N_49344,N_48878,N_48688);
and U49345 (N_49345,N_48092,N_48571);
or U49346 (N_49346,N_48484,N_48962);
and U49347 (N_49347,N_48966,N_48787);
and U49348 (N_49348,N_48156,N_48245);
xnor U49349 (N_49349,N_48083,N_48431);
nor U49350 (N_49350,N_48761,N_48418);
and U49351 (N_49351,N_48304,N_48990);
or U49352 (N_49352,N_48587,N_48567);
nor U49353 (N_49353,N_48117,N_48535);
or U49354 (N_49354,N_48451,N_48809);
nand U49355 (N_49355,N_48255,N_48359);
nor U49356 (N_49356,N_48154,N_48113);
or U49357 (N_49357,N_48580,N_48480);
xor U49358 (N_49358,N_48874,N_48825);
nand U49359 (N_49359,N_48592,N_48303);
and U49360 (N_49360,N_48115,N_48699);
or U49361 (N_49361,N_48534,N_48996);
nand U49362 (N_49362,N_48222,N_48886);
nand U49363 (N_49363,N_48457,N_48782);
nand U49364 (N_49364,N_48609,N_48606);
xor U49365 (N_49365,N_48889,N_48824);
xor U49366 (N_49366,N_48129,N_48549);
xnor U49367 (N_49367,N_48760,N_48089);
xor U49368 (N_49368,N_48929,N_48458);
nor U49369 (N_49369,N_48694,N_48377);
and U49370 (N_49370,N_48979,N_48501);
nor U49371 (N_49371,N_48900,N_48130);
nand U49372 (N_49372,N_48652,N_48204);
nor U49373 (N_49373,N_48021,N_48192);
nor U49374 (N_49374,N_48952,N_48584);
nand U49375 (N_49375,N_48720,N_48753);
or U49376 (N_49376,N_48532,N_48729);
or U49377 (N_49377,N_48147,N_48864);
nor U49378 (N_49378,N_48892,N_48737);
nand U49379 (N_49379,N_48305,N_48376);
nor U49380 (N_49380,N_48186,N_48065);
and U49381 (N_49381,N_48909,N_48752);
xnor U49382 (N_49382,N_48559,N_48314);
nand U49383 (N_49383,N_48462,N_48455);
xor U49384 (N_49384,N_48127,N_48520);
and U49385 (N_49385,N_48098,N_48820);
nand U49386 (N_49386,N_48808,N_48862);
nor U49387 (N_49387,N_48109,N_48703);
xnor U49388 (N_49388,N_48671,N_48324);
xor U49389 (N_49389,N_48440,N_48077);
and U49390 (N_49390,N_48054,N_48141);
and U49391 (N_49391,N_48425,N_48506);
xor U49392 (N_49392,N_48884,N_48100);
or U49393 (N_49393,N_48044,N_48853);
and U49394 (N_49394,N_48335,N_48977);
or U49395 (N_49395,N_48208,N_48790);
xnor U49396 (N_49396,N_48697,N_48407);
xor U49397 (N_49397,N_48636,N_48733);
nor U49398 (N_49398,N_48543,N_48031);
nor U49399 (N_49399,N_48561,N_48296);
nor U49400 (N_49400,N_48539,N_48771);
nand U49401 (N_49401,N_48869,N_48268);
and U49402 (N_49402,N_48603,N_48352);
or U49403 (N_49403,N_48188,N_48062);
or U49404 (N_49404,N_48073,N_48358);
nor U49405 (N_49405,N_48471,N_48249);
and U49406 (N_49406,N_48756,N_48467);
nor U49407 (N_49407,N_48393,N_48482);
nand U49408 (N_49408,N_48649,N_48373);
and U49409 (N_49409,N_48616,N_48950);
nand U49410 (N_49410,N_48747,N_48581);
nand U49411 (N_49411,N_48351,N_48430);
or U49412 (N_49412,N_48794,N_48185);
nor U49413 (N_49413,N_48133,N_48270);
nor U49414 (N_49414,N_48088,N_48702);
nand U49415 (N_49415,N_48211,N_48250);
xor U49416 (N_49416,N_48312,N_48827);
nand U49417 (N_49417,N_48236,N_48897);
xnor U49418 (N_49418,N_48963,N_48672);
nor U49419 (N_49419,N_48429,N_48011);
nor U49420 (N_49420,N_48750,N_48017);
or U49421 (N_49421,N_48472,N_48541);
nor U49422 (N_49422,N_48327,N_48385);
xor U49423 (N_49423,N_48550,N_48165);
nor U49424 (N_49424,N_48217,N_48643);
nor U49425 (N_49425,N_48317,N_48942);
nand U49426 (N_49426,N_48774,N_48492);
nor U49427 (N_49427,N_48673,N_48956);
or U49428 (N_49428,N_48870,N_48380);
nand U49429 (N_49429,N_48604,N_48125);
nor U49430 (N_49430,N_48045,N_48001);
and U49431 (N_49431,N_48547,N_48850);
nand U49432 (N_49432,N_48842,N_48814);
xor U49433 (N_49433,N_48213,N_48839);
or U49434 (N_49434,N_48216,N_48438);
or U49435 (N_49435,N_48992,N_48883);
xnor U49436 (N_49436,N_48854,N_48936);
xor U49437 (N_49437,N_48612,N_48460);
or U49438 (N_49438,N_48171,N_48180);
nand U49439 (N_49439,N_48912,N_48868);
or U49440 (N_49440,N_48364,N_48299);
or U49441 (N_49441,N_48777,N_48201);
nor U49442 (N_49442,N_48610,N_48041);
nor U49443 (N_49443,N_48220,N_48318);
nand U49444 (N_49444,N_48166,N_48730);
and U49445 (N_49445,N_48523,N_48437);
and U49446 (N_49446,N_48097,N_48331);
xor U49447 (N_49447,N_48624,N_48146);
nand U49448 (N_49448,N_48107,N_48494);
nand U49449 (N_49449,N_48622,N_48126);
and U49450 (N_49450,N_48843,N_48101);
and U49451 (N_49451,N_48265,N_48792);
and U49452 (N_49452,N_48829,N_48258);
nand U49453 (N_49453,N_48374,N_48308);
and U49454 (N_49454,N_48005,N_48009);
nor U49455 (N_49455,N_48243,N_48256);
xor U49456 (N_49456,N_48968,N_48574);
and U49457 (N_49457,N_48493,N_48646);
xor U49458 (N_49458,N_48498,N_48264);
or U49459 (N_49459,N_48893,N_48840);
and U49460 (N_49460,N_48674,N_48704);
and U49461 (N_49461,N_48330,N_48091);
nor U49462 (N_49462,N_48896,N_48937);
nand U49463 (N_49463,N_48712,N_48832);
and U49464 (N_49464,N_48105,N_48932);
nor U49465 (N_49465,N_48696,N_48417);
nor U49466 (N_49466,N_48575,N_48885);
nor U49467 (N_49467,N_48029,N_48423);
xor U49468 (N_49468,N_48526,N_48548);
and U49469 (N_49469,N_48191,N_48537);
nand U49470 (N_49470,N_48999,N_48812);
or U49471 (N_49471,N_48503,N_48716);
nand U49472 (N_49472,N_48392,N_48698);
and U49473 (N_49473,N_48871,N_48599);
nor U49474 (N_49474,N_48235,N_48836);
nor U49475 (N_49475,N_48951,N_48251);
or U49476 (N_49476,N_48026,N_48453);
or U49477 (N_49477,N_48834,N_48994);
and U49478 (N_49478,N_48081,N_48748);
nor U49479 (N_49479,N_48495,N_48796);
and U49480 (N_49480,N_48749,N_48941);
and U49481 (N_49481,N_48527,N_48260);
or U49482 (N_49482,N_48396,N_48522);
and U49483 (N_49483,N_48676,N_48542);
xor U49484 (N_49484,N_48006,N_48910);
and U49485 (N_49485,N_48040,N_48611);
nand U49486 (N_49486,N_48569,N_48022);
nand U49487 (N_49487,N_48177,N_48020);
or U49488 (N_49488,N_48555,N_48518);
nor U49489 (N_49489,N_48254,N_48350);
nand U49490 (N_49490,N_48402,N_48320);
or U49491 (N_49491,N_48521,N_48619);
or U49492 (N_49492,N_48297,N_48959);
nor U49493 (N_49493,N_48823,N_48072);
xor U49494 (N_49494,N_48901,N_48626);
nor U49495 (N_49495,N_48273,N_48014);
nor U49496 (N_49496,N_48700,N_48158);
xnor U49497 (N_49497,N_48509,N_48173);
and U49498 (N_49498,N_48206,N_48174);
nor U49499 (N_49499,N_48596,N_48170);
or U49500 (N_49500,N_48554,N_48586);
or U49501 (N_49501,N_48895,N_48912);
nor U49502 (N_49502,N_48826,N_48268);
or U49503 (N_49503,N_48475,N_48950);
or U49504 (N_49504,N_48832,N_48635);
and U49505 (N_49505,N_48252,N_48758);
nor U49506 (N_49506,N_48892,N_48031);
xor U49507 (N_49507,N_48779,N_48666);
xnor U49508 (N_49508,N_48339,N_48386);
or U49509 (N_49509,N_48096,N_48979);
or U49510 (N_49510,N_48739,N_48674);
or U49511 (N_49511,N_48994,N_48396);
nand U49512 (N_49512,N_48957,N_48322);
or U49513 (N_49513,N_48842,N_48191);
and U49514 (N_49514,N_48417,N_48381);
and U49515 (N_49515,N_48178,N_48469);
and U49516 (N_49516,N_48921,N_48852);
nand U49517 (N_49517,N_48849,N_48214);
and U49518 (N_49518,N_48334,N_48254);
xor U49519 (N_49519,N_48115,N_48414);
nor U49520 (N_49520,N_48537,N_48894);
nor U49521 (N_49521,N_48326,N_48598);
nand U49522 (N_49522,N_48439,N_48608);
xor U49523 (N_49523,N_48279,N_48107);
nand U49524 (N_49524,N_48838,N_48087);
or U49525 (N_49525,N_48589,N_48531);
and U49526 (N_49526,N_48989,N_48317);
xnor U49527 (N_49527,N_48481,N_48137);
nor U49528 (N_49528,N_48265,N_48069);
and U49529 (N_49529,N_48070,N_48536);
nor U49530 (N_49530,N_48759,N_48654);
nor U49531 (N_49531,N_48238,N_48329);
nor U49532 (N_49532,N_48580,N_48925);
nor U49533 (N_49533,N_48669,N_48760);
nand U49534 (N_49534,N_48642,N_48842);
nand U49535 (N_49535,N_48436,N_48065);
nor U49536 (N_49536,N_48018,N_48038);
and U49537 (N_49537,N_48091,N_48735);
nand U49538 (N_49538,N_48853,N_48941);
nor U49539 (N_49539,N_48687,N_48518);
nor U49540 (N_49540,N_48723,N_48015);
and U49541 (N_49541,N_48572,N_48336);
nand U49542 (N_49542,N_48991,N_48236);
and U49543 (N_49543,N_48657,N_48939);
or U49544 (N_49544,N_48848,N_48447);
nand U49545 (N_49545,N_48535,N_48173);
xnor U49546 (N_49546,N_48646,N_48498);
and U49547 (N_49547,N_48703,N_48121);
nand U49548 (N_49548,N_48351,N_48440);
or U49549 (N_49549,N_48605,N_48046);
xnor U49550 (N_49550,N_48828,N_48155);
or U49551 (N_49551,N_48493,N_48423);
and U49552 (N_49552,N_48726,N_48952);
nor U49553 (N_49553,N_48743,N_48730);
nand U49554 (N_49554,N_48641,N_48594);
xor U49555 (N_49555,N_48000,N_48749);
nor U49556 (N_49556,N_48059,N_48861);
or U49557 (N_49557,N_48821,N_48125);
xor U49558 (N_49558,N_48206,N_48521);
and U49559 (N_49559,N_48490,N_48312);
nor U49560 (N_49560,N_48010,N_48308);
xnor U49561 (N_49561,N_48186,N_48716);
and U49562 (N_49562,N_48125,N_48390);
or U49563 (N_49563,N_48867,N_48577);
or U49564 (N_49564,N_48586,N_48019);
nor U49565 (N_49565,N_48323,N_48117);
nand U49566 (N_49566,N_48376,N_48718);
xnor U49567 (N_49567,N_48705,N_48432);
nor U49568 (N_49568,N_48327,N_48887);
nand U49569 (N_49569,N_48460,N_48737);
xor U49570 (N_49570,N_48948,N_48197);
and U49571 (N_49571,N_48279,N_48328);
xor U49572 (N_49572,N_48999,N_48767);
nand U49573 (N_49573,N_48297,N_48853);
xnor U49574 (N_49574,N_48646,N_48823);
or U49575 (N_49575,N_48968,N_48764);
xnor U49576 (N_49576,N_48820,N_48889);
nor U49577 (N_49577,N_48610,N_48619);
nor U49578 (N_49578,N_48038,N_48451);
nand U49579 (N_49579,N_48434,N_48077);
xor U49580 (N_49580,N_48253,N_48072);
nand U49581 (N_49581,N_48384,N_48021);
nand U49582 (N_49582,N_48826,N_48736);
nor U49583 (N_49583,N_48536,N_48473);
nor U49584 (N_49584,N_48543,N_48957);
or U49585 (N_49585,N_48301,N_48733);
nand U49586 (N_49586,N_48761,N_48183);
or U49587 (N_49587,N_48467,N_48061);
and U49588 (N_49588,N_48737,N_48358);
or U49589 (N_49589,N_48191,N_48246);
nand U49590 (N_49590,N_48856,N_48787);
or U49591 (N_49591,N_48777,N_48197);
and U49592 (N_49592,N_48206,N_48698);
nor U49593 (N_49593,N_48038,N_48101);
nor U49594 (N_49594,N_48935,N_48352);
and U49595 (N_49595,N_48496,N_48116);
xor U49596 (N_49596,N_48479,N_48609);
nand U49597 (N_49597,N_48218,N_48946);
nor U49598 (N_49598,N_48650,N_48945);
or U49599 (N_49599,N_48845,N_48254);
nand U49600 (N_49600,N_48136,N_48989);
and U49601 (N_49601,N_48735,N_48375);
nand U49602 (N_49602,N_48460,N_48516);
nor U49603 (N_49603,N_48793,N_48265);
and U49604 (N_49604,N_48446,N_48676);
nor U49605 (N_49605,N_48875,N_48830);
or U49606 (N_49606,N_48057,N_48608);
nor U49607 (N_49607,N_48519,N_48735);
xnor U49608 (N_49608,N_48971,N_48429);
nor U49609 (N_49609,N_48708,N_48225);
nor U49610 (N_49610,N_48427,N_48702);
and U49611 (N_49611,N_48638,N_48231);
and U49612 (N_49612,N_48744,N_48735);
xnor U49613 (N_49613,N_48659,N_48133);
xnor U49614 (N_49614,N_48465,N_48974);
and U49615 (N_49615,N_48721,N_48258);
nand U49616 (N_49616,N_48592,N_48244);
and U49617 (N_49617,N_48800,N_48327);
or U49618 (N_49618,N_48499,N_48395);
or U49619 (N_49619,N_48369,N_48930);
nand U49620 (N_49620,N_48813,N_48601);
xor U49621 (N_49621,N_48349,N_48987);
xor U49622 (N_49622,N_48647,N_48409);
xnor U49623 (N_49623,N_48328,N_48611);
nor U49624 (N_49624,N_48222,N_48491);
xor U49625 (N_49625,N_48003,N_48047);
or U49626 (N_49626,N_48930,N_48261);
and U49627 (N_49627,N_48564,N_48669);
and U49628 (N_49628,N_48465,N_48313);
nor U49629 (N_49629,N_48612,N_48404);
or U49630 (N_49630,N_48920,N_48126);
and U49631 (N_49631,N_48140,N_48025);
nor U49632 (N_49632,N_48720,N_48375);
or U49633 (N_49633,N_48718,N_48033);
xnor U49634 (N_49634,N_48264,N_48009);
nand U49635 (N_49635,N_48129,N_48389);
nor U49636 (N_49636,N_48055,N_48690);
nor U49637 (N_49637,N_48908,N_48137);
and U49638 (N_49638,N_48103,N_48354);
xor U49639 (N_49639,N_48139,N_48967);
or U49640 (N_49640,N_48757,N_48697);
nor U49641 (N_49641,N_48755,N_48870);
xnor U49642 (N_49642,N_48501,N_48871);
xnor U49643 (N_49643,N_48873,N_48702);
nor U49644 (N_49644,N_48028,N_48856);
or U49645 (N_49645,N_48621,N_48506);
xor U49646 (N_49646,N_48174,N_48674);
xor U49647 (N_49647,N_48165,N_48803);
and U49648 (N_49648,N_48356,N_48511);
and U49649 (N_49649,N_48946,N_48056);
nor U49650 (N_49650,N_48391,N_48774);
nor U49651 (N_49651,N_48284,N_48351);
and U49652 (N_49652,N_48659,N_48204);
or U49653 (N_49653,N_48680,N_48959);
xor U49654 (N_49654,N_48601,N_48432);
or U49655 (N_49655,N_48445,N_48476);
or U49656 (N_49656,N_48091,N_48968);
xor U49657 (N_49657,N_48444,N_48564);
nand U49658 (N_49658,N_48799,N_48294);
xnor U49659 (N_49659,N_48803,N_48991);
nand U49660 (N_49660,N_48245,N_48323);
nand U49661 (N_49661,N_48469,N_48500);
and U49662 (N_49662,N_48491,N_48828);
or U49663 (N_49663,N_48919,N_48553);
nor U49664 (N_49664,N_48268,N_48766);
nor U49665 (N_49665,N_48675,N_48714);
xnor U49666 (N_49666,N_48719,N_48417);
or U49667 (N_49667,N_48647,N_48562);
or U49668 (N_49668,N_48200,N_48679);
xor U49669 (N_49669,N_48721,N_48458);
and U49670 (N_49670,N_48654,N_48143);
nand U49671 (N_49671,N_48955,N_48154);
nand U49672 (N_49672,N_48685,N_48329);
xor U49673 (N_49673,N_48309,N_48364);
or U49674 (N_49674,N_48747,N_48412);
xor U49675 (N_49675,N_48195,N_48879);
and U49676 (N_49676,N_48230,N_48660);
xor U49677 (N_49677,N_48749,N_48753);
xor U49678 (N_49678,N_48244,N_48773);
or U49679 (N_49679,N_48051,N_48013);
and U49680 (N_49680,N_48147,N_48176);
xnor U49681 (N_49681,N_48497,N_48159);
or U49682 (N_49682,N_48341,N_48568);
nor U49683 (N_49683,N_48917,N_48292);
xnor U49684 (N_49684,N_48712,N_48043);
xor U49685 (N_49685,N_48608,N_48413);
nor U49686 (N_49686,N_48307,N_48407);
xnor U49687 (N_49687,N_48830,N_48685);
and U49688 (N_49688,N_48918,N_48674);
nor U49689 (N_49689,N_48362,N_48433);
and U49690 (N_49690,N_48288,N_48109);
and U49691 (N_49691,N_48749,N_48916);
nand U49692 (N_49692,N_48372,N_48195);
or U49693 (N_49693,N_48784,N_48797);
nor U49694 (N_49694,N_48021,N_48241);
nand U49695 (N_49695,N_48646,N_48288);
or U49696 (N_49696,N_48044,N_48316);
xor U49697 (N_49697,N_48174,N_48129);
or U49698 (N_49698,N_48896,N_48869);
nor U49699 (N_49699,N_48241,N_48533);
nor U49700 (N_49700,N_48081,N_48998);
nand U49701 (N_49701,N_48692,N_48399);
or U49702 (N_49702,N_48294,N_48325);
nor U49703 (N_49703,N_48445,N_48677);
nor U49704 (N_49704,N_48219,N_48760);
and U49705 (N_49705,N_48955,N_48587);
nor U49706 (N_49706,N_48989,N_48400);
xor U49707 (N_49707,N_48867,N_48503);
xor U49708 (N_49708,N_48309,N_48570);
nand U49709 (N_49709,N_48800,N_48995);
or U49710 (N_49710,N_48235,N_48363);
nand U49711 (N_49711,N_48295,N_48708);
or U49712 (N_49712,N_48186,N_48242);
nor U49713 (N_49713,N_48875,N_48327);
nand U49714 (N_49714,N_48304,N_48359);
nand U49715 (N_49715,N_48080,N_48286);
and U49716 (N_49716,N_48470,N_48207);
and U49717 (N_49717,N_48428,N_48870);
or U49718 (N_49718,N_48606,N_48228);
nor U49719 (N_49719,N_48173,N_48137);
nor U49720 (N_49720,N_48842,N_48415);
xor U49721 (N_49721,N_48466,N_48206);
nand U49722 (N_49722,N_48853,N_48716);
and U49723 (N_49723,N_48264,N_48455);
or U49724 (N_49724,N_48663,N_48429);
nor U49725 (N_49725,N_48076,N_48717);
or U49726 (N_49726,N_48452,N_48414);
or U49727 (N_49727,N_48386,N_48993);
nand U49728 (N_49728,N_48662,N_48031);
xor U49729 (N_49729,N_48206,N_48287);
or U49730 (N_49730,N_48178,N_48062);
and U49731 (N_49731,N_48452,N_48486);
nand U49732 (N_49732,N_48349,N_48388);
or U49733 (N_49733,N_48302,N_48542);
nor U49734 (N_49734,N_48068,N_48033);
nand U49735 (N_49735,N_48181,N_48706);
nor U49736 (N_49736,N_48628,N_48855);
and U49737 (N_49737,N_48654,N_48906);
xnor U49738 (N_49738,N_48600,N_48118);
xor U49739 (N_49739,N_48350,N_48901);
nor U49740 (N_49740,N_48734,N_48002);
and U49741 (N_49741,N_48642,N_48978);
nand U49742 (N_49742,N_48381,N_48176);
xor U49743 (N_49743,N_48744,N_48528);
and U49744 (N_49744,N_48838,N_48062);
and U49745 (N_49745,N_48291,N_48194);
nor U49746 (N_49746,N_48193,N_48514);
nand U49747 (N_49747,N_48138,N_48964);
nand U49748 (N_49748,N_48833,N_48414);
or U49749 (N_49749,N_48457,N_48173);
xnor U49750 (N_49750,N_48160,N_48800);
and U49751 (N_49751,N_48230,N_48728);
and U49752 (N_49752,N_48651,N_48576);
or U49753 (N_49753,N_48095,N_48656);
nand U49754 (N_49754,N_48823,N_48721);
nand U49755 (N_49755,N_48621,N_48537);
or U49756 (N_49756,N_48181,N_48077);
or U49757 (N_49757,N_48196,N_48412);
nand U49758 (N_49758,N_48828,N_48535);
nor U49759 (N_49759,N_48748,N_48259);
nor U49760 (N_49760,N_48508,N_48635);
or U49761 (N_49761,N_48590,N_48848);
or U49762 (N_49762,N_48281,N_48919);
xnor U49763 (N_49763,N_48191,N_48901);
or U49764 (N_49764,N_48601,N_48128);
nand U49765 (N_49765,N_48520,N_48502);
nand U49766 (N_49766,N_48965,N_48091);
or U49767 (N_49767,N_48673,N_48321);
and U49768 (N_49768,N_48679,N_48169);
or U49769 (N_49769,N_48922,N_48148);
nand U49770 (N_49770,N_48572,N_48945);
or U49771 (N_49771,N_48492,N_48226);
xor U49772 (N_49772,N_48658,N_48594);
and U49773 (N_49773,N_48040,N_48787);
nor U49774 (N_49774,N_48181,N_48862);
and U49775 (N_49775,N_48696,N_48262);
nand U49776 (N_49776,N_48913,N_48888);
or U49777 (N_49777,N_48356,N_48436);
or U49778 (N_49778,N_48905,N_48844);
xnor U49779 (N_49779,N_48072,N_48650);
nand U49780 (N_49780,N_48112,N_48109);
nand U49781 (N_49781,N_48429,N_48859);
nand U49782 (N_49782,N_48661,N_48558);
and U49783 (N_49783,N_48846,N_48275);
and U49784 (N_49784,N_48104,N_48265);
or U49785 (N_49785,N_48431,N_48745);
nor U49786 (N_49786,N_48497,N_48022);
nor U49787 (N_49787,N_48125,N_48870);
and U49788 (N_49788,N_48469,N_48888);
and U49789 (N_49789,N_48787,N_48706);
xor U49790 (N_49790,N_48115,N_48687);
and U49791 (N_49791,N_48261,N_48219);
and U49792 (N_49792,N_48957,N_48464);
xor U49793 (N_49793,N_48851,N_48766);
nand U49794 (N_49794,N_48847,N_48692);
xor U49795 (N_49795,N_48058,N_48813);
nor U49796 (N_49796,N_48930,N_48837);
or U49797 (N_49797,N_48919,N_48917);
xor U49798 (N_49798,N_48497,N_48101);
xnor U49799 (N_49799,N_48401,N_48829);
nor U49800 (N_49800,N_48713,N_48647);
or U49801 (N_49801,N_48516,N_48418);
and U49802 (N_49802,N_48491,N_48746);
and U49803 (N_49803,N_48216,N_48997);
nand U49804 (N_49804,N_48045,N_48466);
and U49805 (N_49805,N_48323,N_48803);
and U49806 (N_49806,N_48023,N_48265);
xor U49807 (N_49807,N_48151,N_48778);
nor U49808 (N_49808,N_48242,N_48166);
and U49809 (N_49809,N_48812,N_48446);
nand U49810 (N_49810,N_48856,N_48907);
nor U49811 (N_49811,N_48807,N_48496);
and U49812 (N_49812,N_48175,N_48296);
xnor U49813 (N_49813,N_48026,N_48543);
nor U49814 (N_49814,N_48955,N_48128);
and U49815 (N_49815,N_48107,N_48802);
or U49816 (N_49816,N_48826,N_48267);
xnor U49817 (N_49817,N_48403,N_48993);
nor U49818 (N_49818,N_48757,N_48799);
and U49819 (N_49819,N_48000,N_48178);
and U49820 (N_49820,N_48589,N_48323);
nand U49821 (N_49821,N_48288,N_48783);
xnor U49822 (N_49822,N_48989,N_48084);
and U49823 (N_49823,N_48469,N_48998);
and U49824 (N_49824,N_48578,N_48128);
and U49825 (N_49825,N_48171,N_48818);
nand U49826 (N_49826,N_48303,N_48275);
and U49827 (N_49827,N_48960,N_48240);
xor U49828 (N_49828,N_48412,N_48969);
or U49829 (N_49829,N_48922,N_48714);
xor U49830 (N_49830,N_48876,N_48186);
xnor U49831 (N_49831,N_48765,N_48599);
and U49832 (N_49832,N_48980,N_48656);
or U49833 (N_49833,N_48174,N_48832);
xor U49834 (N_49834,N_48311,N_48670);
nand U49835 (N_49835,N_48733,N_48807);
and U49836 (N_49836,N_48431,N_48947);
nand U49837 (N_49837,N_48384,N_48401);
nand U49838 (N_49838,N_48859,N_48535);
or U49839 (N_49839,N_48646,N_48873);
nor U49840 (N_49840,N_48242,N_48730);
and U49841 (N_49841,N_48362,N_48761);
nor U49842 (N_49842,N_48055,N_48346);
nand U49843 (N_49843,N_48003,N_48379);
or U49844 (N_49844,N_48674,N_48033);
nand U49845 (N_49845,N_48888,N_48083);
and U49846 (N_49846,N_48746,N_48026);
xnor U49847 (N_49847,N_48021,N_48945);
or U49848 (N_49848,N_48659,N_48481);
xnor U49849 (N_49849,N_48939,N_48807);
or U49850 (N_49850,N_48538,N_48616);
or U49851 (N_49851,N_48223,N_48630);
or U49852 (N_49852,N_48843,N_48717);
xnor U49853 (N_49853,N_48375,N_48954);
or U49854 (N_49854,N_48153,N_48589);
xnor U49855 (N_49855,N_48983,N_48169);
xnor U49856 (N_49856,N_48869,N_48619);
and U49857 (N_49857,N_48147,N_48817);
and U49858 (N_49858,N_48923,N_48286);
nor U49859 (N_49859,N_48454,N_48781);
and U49860 (N_49860,N_48360,N_48844);
nor U49861 (N_49861,N_48895,N_48770);
nand U49862 (N_49862,N_48556,N_48124);
nor U49863 (N_49863,N_48929,N_48642);
or U49864 (N_49864,N_48902,N_48975);
xor U49865 (N_49865,N_48826,N_48665);
nand U49866 (N_49866,N_48615,N_48188);
and U49867 (N_49867,N_48416,N_48616);
or U49868 (N_49868,N_48831,N_48418);
and U49869 (N_49869,N_48422,N_48264);
and U49870 (N_49870,N_48093,N_48893);
nand U49871 (N_49871,N_48490,N_48765);
nor U49872 (N_49872,N_48256,N_48273);
and U49873 (N_49873,N_48368,N_48564);
nor U49874 (N_49874,N_48293,N_48468);
and U49875 (N_49875,N_48924,N_48832);
nand U49876 (N_49876,N_48892,N_48692);
nor U49877 (N_49877,N_48000,N_48075);
nor U49878 (N_49878,N_48408,N_48784);
nand U49879 (N_49879,N_48241,N_48396);
and U49880 (N_49880,N_48609,N_48297);
nand U49881 (N_49881,N_48969,N_48596);
nand U49882 (N_49882,N_48858,N_48559);
and U49883 (N_49883,N_48493,N_48368);
and U49884 (N_49884,N_48144,N_48624);
nor U49885 (N_49885,N_48307,N_48270);
xor U49886 (N_49886,N_48262,N_48504);
and U49887 (N_49887,N_48936,N_48698);
xnor U49888 (N_49888,N_48710,N_48453);
xnor U49889 (N_49889,N_48428,N_48534);
and U49890 (N_49890,N_48149,N_48686);
or U49891 (N_49891,N_48497,N_48599);
and U49892 (N_49892,N_48197,N_48479);
or U49893 (N_49893,N_48807,N_48020);
nor U49894 (N_49894,N_48299,N_48778);
xor U49895 (N_49895,N_48858,N_48922);
xor U49896 (N_49896,N_48806,N_48562);
nor U49897 (N_49897,N_48480,N_48352);
xor U49898 (N_49898,N_48322,N_48821);
and U49899 (N_49899,N_48203,N_48735);
nand U49900 (N_49900,N_48732,N_48213);
nand U49901 (N_49901,N_48586,N_48542);
nand U49902 (N_49902,N_48352,N_48141);
or U49903 (N_49903,N_48541,N_48084);
nor U49904 (N_49904,N_48202,N_48314);
and U49905 (N_49905,N_48828,N_48223);
nand U49906 (N_49906,N_48866,N_48591);
nand U49907 (N_49907,N_48293,N_48797);
nand U49908 (N_49908,N_48801,N_48459);
nand U49909 (N_49909,N_48013,N_48097);
nor U49910 (N_49910,N_48867,N_48419);
nor U49911 (N_49911,N_48830,N_48485);
nand U49912 (N_49912,N_48932,N_48635);
xor U49913 (N_49913,N_48556,N_48402);
or U49914 (N_49914,N_48168,N_48530);
nor U49915 (N_49915,N_48112,N_48884);
xnor U49916 (N_49916,N_48973,N_48533);
nand U49917 (N_49917,N_48129,N_48743);
or U49918 (N_49918,N_48726,N_48286);
and U49919 (N_49919,N_48260,N_48417);
and U49920 (N_49920,N_48748,N_48867);
nor U49921 (N_49921,N_48856,N_48224);
xnor U49922 (N_49922,N_48484,N_48427);
xnor U49923 (N_49923,N_48869,N_48049);
and U49924 (N_49924,N_48806,N_48723);
and U49925 (N_49925,N_48815,N_48858);
and U49926 (N_49926,N_48185,N_48819);
nor U49927 (N_49927,N_48126,N_48684);
xnor U49928 (N_49928,N_48940,N_48513);
and U49929 (N_49929,N_48639,N_48926);
xnor U49930 (N_49930,N_48246,N_48594);
or U49931 (N_49931,N_48956,N_48826);
or U49932 (N_49932,N_48584,N_48673);
and U49933 (N_49933,N_48009,N_48107);
nand U49934 (N_49934,N_48440,N_48636);
nor U49935 (N_49935,N_48284,N_48326);
xor U49936 (N_49936,N_48113,N_48250);
or U49937 (N_49937,N_48257,N_48283);
xnor U49938 (N_49938,N_48840,N_48734);
or U49939 (N_49939,N_48710,N_48508);
or U49940 (N_49940,N_48980,N_48180);
and U49941 (N_49941,N_48484,N_48299);
nand U49942 (N_49942,N_48203,N_48861);
nand U49943 (N_49943,N_48931,N_48973);
xnor U49944 (N_49944,N_48307,N_48296);
and U49945 (N_49945,N_48657,N_48272);
xnor U49946 (N_49946,N_48800,N_48948);
xnor U49947 (N_49947,N_48878,N_48852);
nor U49948 (N_49948,N_48025,N_48884);
or U49949 (N_49949,N_48486,N_48328);
or U49950 (N_49950,N_48022,N_48014);
nor U49951 (N_49951,N_48415,N_48455);
nand U49952 (N_49952,N_48930,N_48789);
nor U49953 (N_49953,N_48694,N_48371);
or U49954 (N_49954,N_48923,N_48280);
xnor U49955 (N_49955,N_48580,N_48839);
nor U49956 (N_49956,N_48602,N_48451);
or U49957 (N_49957,N_48231,N_48322);
or U49958 (N_49958,N_48403,N_48440);
or U49959 (N_49959,N_48851,N_48300);
nand U49960 (N_49960,N_48139,N_48947);
or U49961 (N_49961,N_48218,N_48314);
or U49962 (N_49962,N_48755,N_48247);
and U49963 (N_49963,N_48152,N_48168);
nand U49964 (N_49964,N_48444,N_48436);
nand U49965 (N_49965,N_48151,N_48210);
xor U49966 (N_49966,N_48944,N_48134);
nor U49967 (N_49967,N_48545,N_48327);
or U49968 (N_49968,N_48566,N_48135);
and U49969 (N_49969,N_48937,N_48053);
xnor U49970 (N_49970,N_48247,N_48535);
and U49971 (N_49971,N_48588,N_48409);
nand U49972 (N_49972,N_48658,N_48049);
nand U49973 (N_49973,N_48804,N_48602);
or U49974 (N_49974,N_48402,N_48658);
nor U49975 (N_49975,N_48529,N_48757);
nand U49976 (N_49976,N_48209,N_48109);
nor U49977 (N_49977,N_48299,N_48259);
or U49978 (N_49978,N_48301,N_48024);
and U49979 (N_49979,N_48987,N_48243);
xor U49980 (N_49980,N_48903,N_48901);
xnor U49981 (N_49981,N_48917,N_48104);
nor U49982 (N_49982,N_48212,N_48096);
and U49983 (N_49983,N_48087,N_48573);
nor U49984 (N_49984,N_48998,N_48797);
nand U49985 (N_49985,N_48366,N_48815);
nor U49986 (N_49986,N_48331,N_48440);
nand U49987 (N_49987,N_48399,N_48335);
nand U49988 (N_49988,N_48165,N_48643);
and U49989 (N_49989,N_48029,N_48916);
xnor U49990 (N_49990,N_48641,N_48954);
xor U49991 (N_49991,N_48068,N_48788);
xnor U49992 (N_49992,N_48751,N_48127);
nand U49993 (N_49993,N_48505,N_48292);
nor U49994 (N_49994,N_48629,N_48812);
or U49995 (N_49995,N_48022,N_48253);
xnor U49996 (N_49996,N_48672,N_48210);
and U49997 (N_49997,N_48671,N_48246);
nand U49998 (N_49998,N_48981,N_48087);
xor U49999 (N_49999,N_48573,N_48878);
and UO_0 (O_0,N_49898,N_49716);
xor UO_1 (O_1,N_49867,N_49086);
or UO_2 (O_2,N_49620,N_49386);
nor UO_3 (O_3,N_49397,N_49407);
nor UO_4 (O_4,N_49769,N_49477);
or UO_5 (O_5,N_49402,N_49980);
and UO_6 (O_6,N_49515,N_49457);
nand UO_7 (O_7,N_49495,N_49277);
or UO_8 (O_8,N_49168,N_49066);
or UO_9 (O_9,N_49332,N_49344);
nand UO_10 (O_10,N_49036,N_49767);
and UO_11 (O_11,N_49764,N_49852);
and UO_12 (O_12,N_49736,N_49831);
xor UO_13 (O_13,N_49482,N_49935);
nand UO_14 (O_14,N_49917,N_49132);
xnor UO_15 (O_15,N_49448,N_49760);
or UO_16 (O_16,N_49556,N_49635);
nand UO_17 (O_17,N_49062,N_49173);
nand UO_18 (O_18,N_49626,N_49869);
or UO_19 (O_19,N_49941,N_49416);
or UO_20 (O_20,N_49424,N_49269);
or UO_21 (O_21,N_49456,N_49149);
nand UO_22 (O_22,N_49591,N_49485);
or UO_23 (O_23,N_49383,N_49193);
nand UO_24 (O_24,N_49678,N_49236);
or UO_25 (O_25,N_49589,N_49296);
nand UO_26 (O_26,N_49988,N_49458);
and UO_27 (O_27,N_49816,N_49195);
xnor UO_28 (O_28,N_49379,N_49549);
and UO_29 (O_29,N_49220,N_49048);
or UO_30 (O_30,N_49654,N_49046);
and UO_31 (O_31,N_49404,N_49892);
and UO_32 (O_32,N_49563,N_49721);
or UO_33 (O_33,N_49599,N_49704);
and UO_34 (O_34,N_49466,N_49776);
nand UO_35 (O_35,N_49749,N_49502);
and UO_36 (O_36,N_49717,N_49580);
and UO_37 (O_37,N_49042,N_49666);
xnor UO_38 (O_38,N_49178,N_49469);
or UO_39 (O_39,N_49262,N_49226);
and UO_40 (O_40,N_49737,N_49326);
xnor UO_41 (O_41,N_49634,N_49096);
xor UO_42 (O_42,N_49569,N_49774);
nand UO_43 (O_43,N_49371,N_49238);
nand UO_44 (O_44,N_49542,N_49446);
nand UO_45 (O_45,N_49090,N_49274);
nor UO_46 (O_46,N_49380,N_49423);
and UO_47 (O_47,N_49786,N_49224);
xor UO_48 (O_48,N_49143,N_49934);
nand UO_49 (O_49,N_49460,N_49147);
and UO_50 (O_50,N_49870,N_49798);
nor UO_51 (O_51,N_49433,N_49302);
nand UO_52 (O_52,N_49865,N_49612);
xor UO_53 (O_53,N_49328,N_49087);
nand UO_54 (O_54,N_49929,N_49291);
xnor UO_55 (O_55,N_49963,N_49520);
nand UO_56 (O_56,N_49053,N_49642);
nand UO_57 (O_57,N_49740,N_49413);
and UO_58 (O_58,N_49576,N_49398);
nor UO_59 (O_59,N_49507,N_49427);
nand UO_60 (O_60,N_49393,N_49058);
or UO_61 (O_61,N_49629,N_49572);
xor UO_62 (O_62,N_49151,N_49996);
and UO_63 (O_63,N_49573,N_49561);
or UO_64 (O_64,N_49000,N_49558);
or UO_65 (O_65,N_49304,N_49973);
and UO_66 (O_66,N_49616,N_49675);
nor UO_67 (O_67,N_49953,N_49182);
nor UO_68 (O_68,N_49258,N_49688);
or UO_69 (O_69,N_49944,N_49043);
or UO_70 (O_70,N_49719,N_49534);
and UO_71 (O_71,N_49985,N_49649);
or UO_72 (O_72,N_49602,N_49134);
and UO_73 (O_73,N_49400,N_49316);
or UO_74 (O_74,N_49505,N_49924);
nor UO_75 (O_75,N_49445,N_49512);
xnor UO_76 (O_76,N_49863,N_49664);
and UO_77 (O_77,N_49327,N_49733);
nor UO_78 (O_78,N_49860,N_49050);
and UO_79 (O_79,N_49028,N_49837);
xor UO_80 (O_80,N_49073,N_49029);
nor UO_81 (O_81,N_49686,N_49611);
or UO_82 (O_82,N_49876,N_49148);
and UO_83 (O_83,N_49116,N_49245);
nor UO_84 (O_84,N_49021,N_49844);
and UO_85 (O_85,N_49905,N_49851);
or UO_86 (O_86,N_49055,N_49259);
nor UO_87 (O_87,N_49590,N_49103);
nand UO_88 (O_88,N_49130,N_49685);
nand UO_89 (O_89,N_49074,N_49481);
or UO_90 (O_90,N_49916,N_49850);
xor UO_91 (O_91,N_49911,N_49637);
xnor UO_92 (O_92,N_49024,N_49191);
or UO_93 (O_93,N_49179,N_49155);
or UO_94 (O_94,N_49289,N_49297);
nand UO_95 (O_95,N_49984,N_49019);
nor UO_96 (O_96,N_49645,N_49468);
or UO_97 (O_97,N_49763,N_49287);
nor UO_98 (O_98,N_49990,N_49146);
or UO_99 (O_99,N_49160,N_49120);
nor UO_100 (O_100,N_49548,N_49267);
nand UO_101 (O_101,N_49777,N_49951);
nand UO_102 (O_102,N_49952,N_49720);
xnor UO_103 (O_103,N_49056,N_49683);
or UO_104 (O_104,N_49336,N_49578);
or UO_105 (O_105,N_49124,N_49701);
and UO_106 (O_106,N_49857,N_49026);
xor UO_107 (O_107,N_49330,N_49199);
xnor UO_108 (O_108,N_49295,N_49473);
nor UO_109 (O_109,N_49110,N_49937);
xnor UO_110 (O_110,N_49757,N_49268);
nor UO_111 (O_111,N_49276,N_49832);
nor UO_112 (O_112,N_49320,N_49765);
nand UO_113 (O_113,N_49725,N_49076);
nor UO_114 (O_114,N_49564,N_49894);
xor UO_115 (O_115,N_49491,N_49756);
and UO_116 (O_116,N_49047,N_49676);
xnor UO_117 (O_117,N_49483,N_49939);
nand UO_118 (O_118,N_49205,N_49444);
nor UO_119 (O_119,N_49750,N_49331);
and UO_120 (O_120,N_49356,N_49521);
or UO_121 (O_121,N_49766,N_49039);
or UO_122 (O_122,N_49970,N_49949);
nor UO_123 (O_123,N_49644,N_49023);
xnor UO_124 (O_124,N_49746,N_49387);
or UO_125 (O_125,N_49464,N_49997);
xnor UO_126 (O_126,N_49809,N_49214);
and UO_127 (O_127,N_49303,N_49715);
or UO_128 (O_128,N_49641,N_49974);
and UO_129 (O_129,N_49097,N_49421);
xnor UO_130 (O_130,N_49022,N_49847);
nand UO_131 (O_131,N_49885,N_49467);
xor UO_132 (O_132,N_49697,N_49801);
or UO_133 (O_133,N_49175,N_49270);
or UO_134 (O_134,N_49030,N_49680);
xnor UO_135 (O_135,N_49946,N_49689);
xnor UO_136 (O_136,N_49229,N_49382);
nand UO_137 (O_137,N_49968,N_49484);
nor UO_138 (O_138,N_49394,N_49188);
nand UO_139 (O_139,N_49511,N_49211);
nor UO_140 (O_140,N_49256,N_49450);
or UO_141 (O_141,N_49595,N_49643);
and UO_142 (O_142,N_49027,N_49044);
nor UO_143 (O_143,N_49806,N_49425);
or UO_144 (O_144,N_49319,N_49235);
and UO_145 (O_145,N_49417,N_49443);
or UO_146 (O_146,N_49560,N_49083);
and UO_147 (O_147,N_49105,N_49557);
and UO_148 (O_148,N_49334,N_49410);
nand UO_149 (O_149,N_49514,N_49159);
and UO_150 (O_150,N_49722,N_49550);
nand UO_151 (O_151,N_49035,N_49691);
nor UO_152 (O_152,N_49693,N_49998);
or UO_153 (O_153,N_49040,N_49755);
and UO_154 (O_154,N_49528,N_49845);
nor UO_155 (O_155,N_49509,N_49977);
nand UO_156 (O_156,N_49575,N_49987);
nor UO_157 (O_157,N_49438,N_49472);
xor UO_158 (O_158,N_49377,N_49165);
or UO_159 (O_159,N_49137,N_49227);
or UO_160 (O_160,N_49032,N_49075);
nor UO_161 (O_161,N_49525,N_49820);
or UO_162 (O_162,N_49903,N_49288);
and UO_163 (O_163,N_49114,N_49785);
and UO_164 (O_164,N_49566,N_49136);
xnor UO_165 (O_165,N_49360,N_49471);
or UO_166 (O_166,N_49872,N_49364);
or UO_167 (O_167,N_49210,N_49372);
xnor UO_168 (O_168,N_49099,N_49699);
nand UO_169 (O_169,N_49093,N_49357);
or UO_170 (O_170,N_49190,N_49546);
nor UO_171 (O_171,N_49418,N_49731);
nand UO_172 (O_172,N_49490,N_49315);
nand UO_173 (O_173,N_49373,N_49221);
and UO_174 (O_174,N_49758,N_49462);
xnor UO_175 (O_175,N_49249,N_49436);
and UO_176 (O_176,N_49636,N_49966);
xnor UO_177 (O_177,N_49228,N_49687);
and UO_178 (O_178,N_49014,N_49431);
and UO_179 (O_179,N_49011,N_49955);
and UO_180 (O_180,N_49871,N_49234);
or UO_181 (O_181,N_49950,N_49796);
or UO_182 (O_182,N_49582,N_49351);
nand UO_183 (O_183,N_49705,N_49031);
nand UO_184 (O_184,N_49792,N_49419);
and UO_185 (O_185,N_49913,N_49257);
and UO_186 (O_186,N_49299,N_49936);
xnor UO_187 (O_187,N_49598,N_49972);
or UO_188 (O_188,N_49638,N_49895);
or UO_189 (O_189,N_49735,N_49025);
nor UO_190 (O_190,N_49005,N_49426);
nor UO_191 (O_191,N_49565,N_49310);
xor UO_192 (O_192,N_49271,N_49216);
xnor UO_193 (O_193,N_49501,N_49335);
nor UO_194 (O_194,N_49745,N_49633);
nand UO_195 (O_195,N_49324,N_49923);
or UO_196 (O_196,N_49215,N_49140);
xor UO_197 (O_197,N_49298,N_49663);
nor UO_198 (O_198,N_49807,N_49054);
xor UO_199 (O_199,N_49711,N_49907);
nor UO_200 (O_200,N_49102,N_49539);
nand UO_201 (O_201,N_49399,N_49157);
or UO_202 (O_202,N_49442,N_49695);
or UO_203 (O_203,N_49346,N_49975);
xnor UO_204 (O_204,N_49339,N_49051);
and UO_205 (O_205,N_49883,N_49192);
nor UO_206 (O_206,N_49703,N_49574);
nor UO_207 (O_207,N_49170,N_49470);
xnor UO_208 (O_208,N_49150,N_49690);
and UO_209 (O_209,N_49367,N_49497);
nand UO_210 (O_210,N_49833,N_49194);
nor UO_211 (O_211,N_49583,N_49206);
and UO_212 (O_212,N_49932,N_49815);
or UO_213 (O_213,N_49655,N_49016);
nor UO_214 (O_214,N_49474,N_49899);
nand UO_215 (O_215,N_49255,N_49873);
nor UO_216 (O_216,N_49494,N_49240);
and UO_217 (O_217,N_49840,N_49180);
xor UO_218 (O_218,N_49762,N_49181);
and UO_219 (O_219,N_49734,N_49784);
nor UO_220 (O_220,N_49909,N_49329);
and UO_221 (O_221,N_49125,N_49706);
and UO_222 (O_222,N_49712,N_49825);
nand UO_223 (O_223,N_49788,N_49089);
xor UO_224 (O_224,N_49604,N_49354);
or UO_225 (O_225,N_49415,N_49392);
and UO_226 (O_226,N_49782,N_49004);
or UO_227 (O_227,N_49928,N_49012);
and UO_228 (O_228,N_49001,N_49080);
nand UO_229 (O_229,N_49547,N_49698);
nor UO_230 (O_230,N_49529,N_49463);
xnor UO_231 (O_231,N_49488,N_49059);
xnor UO_232 (O_232,N_49803,N_49586);
nor UO_233 (O_233,N_49897,N_49954);
xor UO_234 (O_234,N_49524,N_49239);
xor UO_235 (O_235,N_49640,N_49724);
and UO_236 (O_236,N_49684,N_49006);
xor UO_237 (O_237,N_49628,N_49605);
xnor UO_238 (O_238,N_49535,N_49945);
nand UO_239 (O_239,N_49829,N_49665);
or UO_240 (O_240,N_49652,N_49835);
or UO_241 (O_241,N_49246,N_49805);
nor UO_242 (O_242,N_49625,N_49587);
xnor UO_243 (O_243,N_49958,N_49186);
nand UO_244 (O_244,N_49848,N_49127);
nor UO_245 (O_245,N_49217,N_49250);
and UO_246 (O_246,N_49201,N_49748);
nor UO_247 (O_247,N_49993,N_49381);
or UO_248 (O_248,N_49893,N_49122);
nor UO_249 (O_249,N_49253,N_49992);
or UO_250 (O_250,N_49275,N_49668);
nor UO_251 (O_251,N_49614,N_49311);
nor UO_252 (O_252,N_49995,N_49409);
nand UO_253 (O_253,N_49607,N_49117);
nand UO_254 (O_254,N_49422,N_49077);
nor UO_255 (O_255,N_49478,N_49588);
or UO_256 (O_256,N_49121,N_49260);
or UO_257 (O_257,N_49523,N_49538);
nor UO_258 (O_258,N_49592,N_49522);
and UO_259 (O_259,N_49541,N_49811);
or UO_260 (O_260,N_49670,N_49709);
or UO_261 (O_261,N_49967,N_49317);
nand UO_262 (O_262,N_49553,N_49323);
nor UO_263 (O_263,N_49849,N_49779);
nor UO_264 (O_264,N_49904,N_49730);
nor UO_265 (O_265,N_49453,N_49577);
nand UO_266 (O_266,N_49884,N_49183);
nand UO_267 (O_267,N_49933,N_49219);
nor UO_268 (O_268,N_49536,N_49931);
nor UO_269 (O_269,N_49049,N_49771);
xor UO_270 (O_270,N_49139,N_49804);
xor UO_271 (O_271,N_49601,N_49808);
nand UO_272 (O_272,N_49751,N_49406);
xnor UO_273 (O_273,N_49496,N_49348);
nor UO_274 (O_274,N_49773,N_49994);
nor UO_275 (O_275,N_49233,N_49981);
nor UO_276 (O_276,N_49581,N_49651);
nor UO_277 (O_277,N_49864,N_49321);
nand UO_278 (O_278,N_49340,N_49437);
nor UO_279 (O_279,N_49648,N_49091);
xor UO_280 (O_280,N_49184,N_49278);
nor UO_281 (O_281,N_49878,N_49540);
and UO_282 (O_282,N_49414,N_49843);
and UO_283 (O_283,N_49113,N_49622);
and UO_284 (O_284,N_49358,N_49639);
or UO_285 (O_285,N_49119,N_49202);
or UO_286 (O_286,N_49133,N_49070);
or UO_287 (O_287,N_49013,N_49567);
nand UO_288 (O_288,N_49307,N_49244);
and UO_289 (O_289,N_49284,N_49243);
or UO_290 (O_290,N_49700,N_49728);
nand UO_291 (O_291,N_49208,N_49498);
and UO_292 (O_292,N_49608,N_49585);
nand UO_293 (O_293,N_49082,N_49964);
xnor UO_294 (O_294,N_49681,N_49999);
nand UO_295 (O_295,N_49842,N_49938);
nor UO_296 (O_296,N_49669,N_49508);
nand UO_297 (O_297,N_49617,N_49609);
and UO_298 (O_298,N_49353,N_49754);
nor UO_299 (O_299,N_49866,N_49230);
nor UO_300 (O_300,N_49362,N_49799);
and UO_301 (O_301,N_49504,N_49017);
or UO_302 (O_302,N_49085,N_49570);
and UO_303 (O_303,N_49991,N_49252);
and UO_304 (O_304,N_49828,N_49197);
nand UO_305 (O_305,N_49493,N_49887);
and UO_306 (O_306,N_49795,N_49727);
xor UO_307 (O_307,N_49962,N_49225);
or UO_308 (O_308,N_49374,N_49069);
xor UO_309 (O_309,N_49821,N_49266);
nor UO_310 (O_310,N_49823,N_49610);
or UO_311 (O_311,N_49623,N_49290);
nand UO_312 (O_312,N_49824,N_49812);
or UO_313 (O_313,N_49264,N_49817);
or UO_314 (O_314,N_49826,N_49794);
nor UO_315 (O_315,N_49942,N_49403);
xnor UO_316 (O_316,N_49562,N_49067);
nand UO_317 (O_317,N_49752,N_49888);
xnor UO_318 (O_318,N_49877,N_49692);
or UO_319 (O_319,N_49355,N_49956);
or UO_320 (O_320,N_49465,N_49673);
or UO_321 (O_321,N_49499,N_49231);
nand UO_322 (O_322,N_49447,N_49101);
or UO_323 (O_323,N_49510,N_49915);
nor UO_324 (O_324,N_49107,N_49247);
xor UO_325 (O_325,N_49218,N_49710);
or UO_326 (O_326,N_49279,N_49187);
or UO_327 (O_327,N_49272,N_49947);
nand UO_328 (O_328,N_49242,N_49532);
or UO_329 (O_329,N_49606,N_49982);
nand UO_330 (O_330,N_49880,N_49232);
nor UO_331 (O_331,N_49891,N_49775);
nand UO_332 (O_332,N_49209,N_49830);
nor UO_333 (O_333,N_49619,N_49677);
or UO_334 (O_334,N_49631,N_49144);
xnor UO_335 (O_335,N_49081,N_49434);
nand UO_336 (O_336,N_49002,N_49827);
and UO_337 (O_337,N_49435,N_49660);
xnor UO_338 (O_338,N_49385,N_49222);
or UO_339 (O_339,N_49248,N_49350);
nor UO_340 (O_340,N_49624,N_49411);
and UO_341 (O_341,N_49060,N_49797);
nand UO_342 (O_342,N_49312,N_49095);
nor UO_343 (O_343,N_49533,N_49976);
xnor UO_344 (O_344,N_49034,N_49742);
nor UO_345 (O_345,N_49322,N_49822);
or UO_346 (O_346,N_49943,N_49918);
and UO_347 (O_347,N_49818,N_49841);
and UO_348 (O_348,N_49780,N_49768);
or UO_349 (O_349,N_49875,N_49650);
or UO_350 (O_350,N_49037,N_49111);
xnor UO_351 (O_351,N_49166,N_49896);
nor UO_352 (O_352,N_49961,N_49571);
xnor UO_353 (O_353,N_49632,N_49855);
nand UO_354 (O_354,N_49858,N_49429);
and UO_355 (O_355,N_49057,N_49161);
nand UO_356 (O_356,N_49959,N_49738);
xnor UO_357 (O_357,N_49500,N_49045);
nor UO_358 (O_358,N_49084,N_49342);
and UO_359 (O_359,N_49171,N_49544);
xnor UO_360 (O_360,N_49531,N_49551);
nor UO_361 (O_361,N_49859,N_49273);
nand UO_362 (O_362,N_49106,N_49554);
and UO_363 (O_363,N_49714,N_49781);
and UO_364 (O_364,N_49789,N_49753);
nor UO_365 (O_365,N_49241,N_49621);
nand UO_366 (O_366,N_49378,N_49071);
and UO_367 (O_367,N_49886,N_49401);
nor UO_368 (O_368,N_49702,N_49128);
xnor UO_369 (O_369,N_49600,N_49008);
nand UO_370 (O_370,N_49492,N_49223);
nand UO_371 (O_371,N_49627,N_49881);
nor UO_372 (O_372,N_49741,N_49072);
nand UO_373 (O_373,N_49015,N_49674);
or UO_374 (O_374,N_49363,N_49459);
nor UO_375 (O_375,N_49603,N_49196);
or UO_376 (O_376,N_49527,N_49517);
xor UO_377 (O_377,N_49694,N_49889);
xor UO_378 (O_378,N_49552,N_49778);
nand UO_379 (O_379,N_49940,N_49439);
nand UO_380 (O_380,N_49347,N_49141);
or UO_381 (O_381,N_49518,N_49530);
nand UO_382 (O_382,N_49519,N_49819);
or UO_383 (O_383,N_49732,N_49454);
xor UO_384 (O_384,N_49584,N_49318);
and UO_385 (O_385,N_49169,N_49018);
nor UO_386 (O_386,N_49365,N_49543);
xor UO_387 (O_387,N_49920,N_49744);
and UO_388 (O_388,N_49203,N_49559);
nor UO_389 (O_389,N_49516,N_49679);
xnor UO_390 (O_390,N_49325,N_49428);
nor UO_391 (O_391,N_49957,N_49914);
xor UO_392 (O_392,N_49513,N_49979);
or UO_393 (O_393,N_49912,N_49667);
xnor UO_394 (O_394,N_49882,N_49910);
and UO_395 (O_395,N_49921,N_49930);
nor UO_396 (O_396,N_49747,N_49713);
nor UO_397 (O_397,N_49696,N_49254);
or UO_398 (O_398,N_49739,N_49900);
or UO_399 (O_399,N_49761,N_49856);
and UO_400 (O_400,N_49879,N_49009);
or UO_401 (O_401,N_49432,N_49671);
nor UO_402 (O_402,N_49594,N_49682);
nor UO_403 (O_403,N_49396,N_49568);
or UO_404 (O_404,N_49294,N_49853);
nor UO_405 (O_405,N_49185,N_49449);
or UO_406 (O_406,N_49301,N_49007);
nand UO_407 (O_407,N_49145,N_49306);
and UO_408 (O_408,N_49176,N_49345);
or UO_409 (O_409,N_49659,N_49265);
and UO_410 (O_410,N_49545,N_49376);
xnor UO_411 (O_411,N_49341,N_49476);
or UO_412 (O_412,N_49177,N_49813);
or UO_413 (O_413,N_49333,N_49451);
nor UO_414 (O_414,N_49292,N_49172);
nor UO_415 (O_415,N_49908,N_49926);
xor UO_416 (O_416,N_49109,N_49251);
xor UO_417 (O_417,N_49647,N_49352);
and UO_418 (O_418,N_49375,N_49906);
and UO_419 (O_419,N_49868,N_49068);
or UO_420 (O_420,N_49661,N_49092);
nor UO_421 (O_421,N_49033,N_49153);
or UO_422 (O_422,N_49237,N_49293);
nand UO_423 (O_423,N_49480,N_49486);
and UO_424 (O_424,N_49135,N_49919);
and UO_425 (O_425,N_49391,N_49041);
nand UO_426 (O_426,N_49922,N_49593);
nand UO_427 (O_427,N_49003,N_49479);
and UO_428 (O_428,N_49138,N_49729);
xnor UO_429 (O_429,N_49846,N_49198);
and UO_430 (O_430,N_49597,N_49280);
and UO_431 (O_431,N_49408,N_49978);
xnor UO_432 (O_432,N_49395,N_49369);
nor UO_433 (O_433,N_49154,N_49613);
or UO_434 (O_434,N_49174,N_49388);
xnor UO_435 (O_435,N_49723,N_49020);
nor UO_436 (O_436,N_49094,N_49207);
nor UO_437 (O_437,N_49506,N_49286);
and UO_438 (O_438,N_49118,N_49213);
or UO_439 (O_439,N_49098,N_49052);
and UO_440 (O_440,N_49800,N_49791);
nand UO_441 (O_441,N_49361,N_49440);
nand UO_442 (O_442,N_49455,N_49489);
or UO_443 (O_443,N_49285,N_49983);
nor UO_444 (O_444,N_49389,N_49309);
nor UO_445 (O_445,N_49142,N_49874);
xor UO_446 (O_446,N_49263,N_49167);
nor UO_447 (O_447,N_49861,N_49461);
nand UO_448 (O_448,N_49162,N_49010);
or UO_449 (O_449,N_49366,N_49989);
xor UO_450 (O_450,N_49038,N_49129);
or UO_451 (O_451,N_49960,N_49793);
nand UO_452 (O_452,N_49115,N_49718);
xor UO_453 (O_453,N_49305,N_49969);
and UO_454 (O_454,N_49579,N_49079);
nand UO_455 (O_455,N_49927,N_49338);
or UO_456 (O_456,N_49596,N_49064);
nor UO_457 (O_457,N_49475,N_49487);
xnor UO_458 (O_458,N_49646,N_49707);
nand UO_459 (O_459,N_49783,N_49152);
or UO_460 (O_460,N_49787,N_49759);
nand UO_461 (O_461,N_49065,N_49405);
and UO_462 (O_462,N_49063,N_49200);
and UO_463 (O_463,N_49313,N_49283);
or UO_464 (O_464,N_49810,N_49123);
xnor UO_465 (O_465,N_49163,N_49281);
nand UO_466 (O_466,N_49615,N_49537);
xnor UO_467 (O_467,N_49672,N_49503);
nand UO_468 (O_468,N_49158,N_49349);
nor UO_469 (O_469,N_49901,N_49986);
or UO_470 (O_470,N_49662,N_49839);
nor UO_471 (O_471,N_49854,N_49526);
and UO_472 (O_472,N_49390,N_49555);
xor UO_473 (O_473,N_49862,N_49925);
xor UO_474 (O_474,N_49261,N_49359);
nand UO_475 (O_475,N_49802,N_49420);
xor UO_476 (O_476,N_49314,N_49656);
nor UO_477 (O_477,N_49441,N_49061);
xor UO_478 (O_478,N_49189,N_49834);
xnor UO_479 (O_479,N_49630,N_49088);
nor UO_480 (O_480,N_49112,N_49836);
xor UO_481 (O_481,N_49343,N_49104);
or UO_482 (O_482,N_49948,N_49653);
nand UO_483 (O_483,N_49131,N_49838);
nor UO_484 (O_484,N_49204,N_49078);
and UO_485 (O_485,N_49708,N_49814);
or UO_486 (O_486,N_49156,N_49618);
and UO_487 (O_487,N_49212,N_49772);
or UO_488 (O_488,N_49726,N_49965);
xnor UO_489 (O_489,N_49971,N_49100);
nor UO_490 (O_490,N_49770,N_49308);
xor UO_491 (O_491,N_49430,N_49126);
nand UO_492 (O_492,N_49164,N_49368);
nand UO_493 (O_493,N_49890,N_49658);
nand UO_494 (O_494,N_49300,N_49282);
and UO_495 (O_495,N_49370,N_49902);
nand UO_496 (O_496,N_49412,N_49384);
and UO_497 (O_497,N_49452,N_49108);
nand UO_498 (O_498,N_49790,N_49743);
nand UO_499 (O_499,N_49337,N_49657);
xor UO_500 (O_500,N_49333,N_49112);
xnor UO_501 (O_501,N_49428,N_49523);
nand UO_502 (O_502,N_49759,N_49404);
nand UO_503 (O_503,N_49484,N_49147);
and UO_504 (O_504,N_49536,N_49363);
nor UO_505 (O_505,N_49229,N_49575);
or UO_506 (O_506,N_49930,N_49159);
and UO_507 (O_507,N_49995,N_49777);
nand UO_508 (O_508,N_49859,N_49245);
xnor UO_509 (O_509,N_49272,N_49913);
nand UO_510 (O_510,N_49961,N_49257);
nor UO_511 (O_511,N_49412,N_49852);
nand UO_512 (O_512,N_49298,N_49216);
xor UO_513 (O_513,N_49962,N_49312);
xor UO_514 (O_514,N_49253,N_49956);
or UO_515 (O_515,N_49904,N_49080);
and UO_516 (O_516,N_49549,N_49728);
nand UO_517 (O_517,N_49218,N_49367);
nand UO_518 (O_518,N_49862,N_49091);
or UO_519 (O_519,N_49719,N_49148);
nand UO_520 (O_520,N_49736,N_49554);
nand UO_521 (O_521,N_49665,N_49115);
nor UO_522 (O_522,N_49378,N_49972);
and UO_523 (O_523,N_49250,N_49282);
nand UO_524 (O_524,N_49866,N_49153);
nor UO_525 (O_525,N_49920,N_49226);
nand UO_526 (O_526,N_49950,N_49549);
nor UO_527 (O_527,N_49266,N_49614);
and UO_528 (O_528,N_49110,N_49261);
and UO_529 (O_529,N_49027,N_49430);
and UO_530 (O_530,N_49391,N_49614);
xor UO_531 (O_531,N_49644,N_49533);
xor UO_532 (O_532,N_49517,N_49365);
or UO_533 (O_533,N_49716,N_49947);
and UO_534 (O_534,N_49304,N_49279);
nand UO_535 (O_535,N_49241,N_49538);
nor UO_536 (O_536,N_49065,N_49675);
or UO_537 (O_537,N_49699,N_49910);
xor UO_538 (O_538,N_49614,N_49702);
nor UO_539 (O_539,N_49821,N_49646);
and UO_540 (O_540,N_49218,N_49435);
nand UO_541 (O_541,N_49239,N_49955);
nor UO_542 (O_542,N_49206,N_49892);
nand UO_543 (O_543,N_49175,N_49685);
nor UO_544 (O_544,N_49865,N_49979);
xor UO_545 (O_545,N_49507,N_49384);
xnor UO_546 (O_546,N_49041,N_49333);
nor UO_547 (O_547,N_49967,N_49581);
nor UO_548 (O_548,N_49313,N_49534);
nand UO_549 (O_549,N_49047,N_49013);
or UO_550 (O_550,N_49715,N_49644);
nor UO_551 (O_551,N_49198,N_49058);
nor UO_552 (O_552,N_49776,N_49931);
and UO_553 (O_553,N_49781,N_49851);
or UO_554 (O_554,N_49578,N_49125);
nand UO_555 (O_555,N_49958,N_49120);
and UO_556 (O_556,N_49793,N_49123);
xor UO_557 (O_557,N_49948,N_49511);
or UO_558 (O_558,N_49166,N_49130);
nand UO_559 (O_559,N_49011,N_49163);
or UO_560 (O_560,N_49873,N_49583);
or UO_561 (O_561,N_49650,N_49395);
or UO_562 (O_562,N_49306,N_49392);
and UO_563 (O_563,N_49506,N_49707);
nand UO_564 (O_564,N_49401,N_49443);
and UO_565 (O_565,N_49659,N_49518);
or UO_566 (O_566,N_49802,N_49540);
or UO_567 (O_567,N_49655,N_49273);
nand UO_568 (O_568,N_49449,N_49553);
and UO_569 (O_569,N_49582,N_49973);
nand UO_570 (O_570,N_49682,N_49653);
and UO_571 (O_571,N_49342,N_49968);
or UO_572 (O_572,N_49360,N_49877);
nor UO_573 (O_573,N_49302,N_49879);
or UO_574 (O_574,N_49285,N_49142);
xor UO_575 (O_575,N_49674,N_49053);
nor UO_576 (O_576,N_49561,N_49574);
and UO_577 (O_577,N_49955,N_49903);
or UO_578 (O_578,N_49670,N_49301);
or UO_579 (O_579,N_49484,N_49362);
or UO_580 (O_580,N_49673,N_49310);
nor UO_581 (O_581,N_49350,N_49232);
nor UO_582 (O_582,N_49020,N_49888);
nor UO_583 (O_583,N_49640,N_49948);
or UO_584 (O_584,N_49076,N_49003);
and UO_585 (O_585,N_49620,N_49052);
nand UO_586 (O_586,N_49989,N_49470);
nor UO_587 (O_587,N_49229,N_49293);
and UO_588 (O_588,N_49751,N_49098);
nor UO_589 (O_589,N_49692,N_49636);
nand UO_590 (O_590,N_49794,N_49937);
nand UO_591 (O_591,N_49129,N_49818);
and UO_592 (O_592,N_49101,N_49557);
nand UO_593 (O_593,N_49408,N_49884);
nand UO_594 (O_594,N_49643,N_49832);
xnor UO_595 (O_595,N_49676,N_49289);
and UO_596 (O_596,N_49649,N_49534);
nor UO_597 (O_597,N_49295,N_49703);
or UO_598 (O_598,N_49836,N_49361);
nand UO_599 (O_599,N_49089,N_49097);
nor UO_600 (O_600,N_49391,N_49445);
and UO_601 (O_601,N_49446,N_49273);
nor UO_602 (O_602,N_49802,N_49180);
nor UO_603 (O_603,N_49896,N_49135);
nand UO_604 (O_604,N_49765,N_49932);
nor UO_605 (O_605,N_49872,N_49874);
nor UO_606 (O_606,N_49715,N_49541);
nand UO_607 (O_607,N_49051,N_49458);
xnor UO_608 (O_608,N_49137,N_49218);
or UO_609 (O_609,N_49811,N_49144);
nor UO_610 (O_610,N_49777,N_49550);
xnor UO_611 (O_611,N_49799,N_49958);
or UO_612 (O_612,N_49315,N_49726);
or UO_613 (O_613,N_49038,N_49754);
or UO_614 (O_614,N_49123,N_49574);
xor UO_615 (O_615,N_49428,N_49128);
nand UO_616 (O_616,N_49410,N_49364);
xnor UO_617 (O_617,N_49128,N_49874);
and UO_618 (O_618,N_49306,N_49113);
or UO_619 (O_619,N_49204,N_49631);
or UO_620 (O_620,N_49702,N_49885);
or UO_621 (O_621,N_49669,N_49096);
nand UO_622 (O_622,N_49459,N_49997);
or UO_623 (O_623,N_49442,N_49544);
nand UO_624 (O_624,N_49912,N_49523);
xnor UO_625 (O_625,N_49424,N_49958);
xnor UO_626 (O_626,N_49100,N_49755);
or UO_627 (O_627,N_49461,N_49142);
nor UO_628 (O_628,N_49141,N_49503);
or UO_629 (O_629,N_49190,N_49415);
and UO_630 (O_630,N_49930,N_49933);
nor UO_631 (O_631,N_49116,N_49528);
and UO_632 (O_632,N_49975,N_49818);
and UO_633 (O_633,N_49455,N_49950);
nand UO_634 (O_634,N_49216,N_49929);
and UO_635 (O_635,N_49341,N_49766);
nand UO_636 (O_636,N_49300,N_49520);
and UO_637 (O_637,N_49163,N_49550);
nand UO_638 (O_638,N_49327,N_49061);
and UO_639 (O_639,N_49475,N_49323);
and UO_640 (O_640,N_49805,N_49893);
nand UO_641 (O_641,N_49847,N_49016);
xnor UO_642 (O_642,N_49873,N_49249);
nor UO_643 (O_643,N_49172,N_49589);
or UO_644 (O_644,N_49374,N_49370);
xor UO_645 (O_645,N_49461,N_49561);
nor UO_646 (O_646,N_49656,N_49537);
nor UO_647 (O_647,N_49329,N_49097);
or UO_648 (O_648,N_49357,N_49109);
or UO_649 (O_649,N_49462,N_49784);
or UO_650 (O_650,N_49167,N_49183);
nand UO_651 (O_651,N_49991,N_49344);
nor UO_652 (O_652,N_49017,N_49122);
or UO_653 (O_653,N_49793,N_49712);
and UO_654 (O_654,N_49735,N_49752);
nand UO_655 (O_655,N_49624,N_49676);
xor UO_656 (O_656,N_49925,N_49600);
or UO_657 (O_657,N_49936,N_49711);
or UO_658 (O_658,N_49074,N_49030);
xor UO_659 (O_659,N_49217,N_49037);
xnor UO_660 (O_660,N_49224,N_49655);
nor UO_661 (O_661,N_49764,N_49748);
xor UO_662 (O_662,N_49413,N_49857);
or UO_663 (O_663,N_49107,N_49427);
and UO_664 (O_664,N_49241,N_49602);
and UO_665 (O_665,N_49909,N_49254);
and UO_666 (O_666,N_49337,N_49153);
nor UO_667 (O_667,N_49048,N_49464);
and UO_668 (O_668,N_49508,N_49795);
or UO_669 (O_669,N_49894,N_49941);
and UO_670 (O_670,N_49791,N_49741);
nor UO_671 (O_671,N_49449,N_49082);
and UO_672 (O_672,N_49012,N_49497);
or UO_673 (O_673,N_49488,N_49945);
or UO_674 (O_674,N_49537,N_49751);
and UO_675 (O_675,N_49000,N_49810);
or UO_676 (O_676,N_49601,N_49760);
and UO_677 (O_677,N_49712,N_49741);
nand UO_678 (O_678,N_49559,N_49344);
and UO_679 (O_679,N_49370,N_49388);
and UO_680 (O_680,N_49782,N_49275);
nand UO_681 (O_681,N_49199,N_49288);
nor UO_682 (O_682,N_49840,N_49494);
or UO_683 (O_683,N_49969,N_49233);
or UO_684 (O_684,N_49880,N_49231);
nand UO_685 (O_685,N_49602,N_49550);
xor UO_686 (O_686,N_49389,N_49444);
nand UO_687 (O_687,N_49947,N_49051);
or UO_688 (O_688,N_49225,N_49427);
and UO_689 (O_689,N_49910,N_49362);
and UO_690 (O_690,N_49546,N_49375);
or UO_691 (O_691,N_49085,N_49691);
or UO_692 (O_692,N_49262,N_49394);
xor UO_693 (O_693,N_49283,N_49228);
nor UO_694 (O_694,N_49627,N_49451);
and UO_695 (O_695,N_49529,N_49507);
and UO_696 (O_696,N_49411,N_49676);
and UO_697 (O_697,N_49625,N_49357);
and UO_698 (O_698,N_49947,N_49871);
xnor UO_699 (O_699,N_49497,N_49979);
nor UO_700 (O_700,N_49256,N_49824);
nor UO_701 (O_701,N_49430,N_49593);
nor UO_702 (O_702,N_49739,N_49154);
xnor UO_703 (O_703,N_49282,N_49377);
or UO_704 (O_704,N_49684,N_49861);
xor UO_705 (O_705,N_49320,N_49038);
xor UO_706 (O_706,N_49077,N_49162);
nand UO_707 (O_707,N_49445,N_49493);
nand UO_708 (O_708,N_49337,N_49760);
or UO_709 (O_709,N_49963,N_49176);
or UO_710 (O_710,N_49293,N_49573);
nor UO_711 (O_711,N_49946,N_49823);
or UO_712 (O_712,N_49254,N_49772);
xnor UO_713 (O_713,N_49959,N_49932);
or UO_714 (O_714,N_49054,N_49713);
xnor UO_715 (O_715,N_49128,N_49912);
or UO_716 (O_716,N_49129,N_49513);
or UO_717 (O_717,N_49890,N_49452);
nand UO_718 (O_718,N_49220,N_49569);
xor UO_719 (O_719,N_49252,N_49977);
or UO_720 (O_720,N_49171,N_49555);
or UO_721 (O_721,N_49763,N_49045);
or UO_722 (O_722,N_49642,N_49393);
and UO_723 (O_723,N_49122,N_49422);
xnor UO_724 (O_724,N_49812,N_49610);
nor UO_725 (O_725,N_49788,N_49696);
xor UO_726 (O_726,N_49310,N_49136);
or UO_727 (O_727,N_49288,N_49781);
nand UO_728 (O_728,N_49055,N_49131);
or UO_729 (O_729,N_49070,N_49806);
nand UO_730 (O_730,N_49871,N_49894);
or UO_731 (O_731,N_49469,N_49291);
nand UO_732 (O_732,N_49599,N_49790);
nor UO_733 (O_733,N_49552,N_49395);
nand UO_734 (O_734,N_49984,N_49820);
and UO_735 (O_735,N_49326,N_49359);
nand UO_736 (O_736,N_49198,N_49131);
or UO_737 (O_737,N_49216,N_49715);
nand UO_738 (O_738,N_49587,N_49764);
xnor UO_739 (O_739,N_49046,N_49740);
or UO_740 (O_740,N_49241,N_49853);
or UO_741 (O_741,N_49710,N_49909);
xor UO_742 (O_742,N_49356,N_49409);
or UO_743 (O_743,N_49911,N_49638);
and UO_744 (O_744,N_49675,N_49491);
or UO_745 (O_745,N_49348,N_49424);
xnor UO_746 (O_746,N_49256,N_49107);
or UO_747 (O_747,N_49555,N_49047);
or UO_748 (O_748,N_49385,N_49930);
nand UO_749 (O_749,N_49921,N_49671);
xnor UO_750 (O_750,N_49495,N_49442);
or UO_751 (O_751,N_49857,N_49578);
nand UO_752 (O_752,N_49138,N_49801);
nand UO_753 (O_753,N_49322,N_49649);
xnor UO_754 (O_754,N_49130,N_49858);
or UO_755 (O_755,N_49532,N_49270);
nor UO_756 (O_756,N_49782,N_49276);
nor UO_757 (O_757,N_49021,N_49149);
nand UO_758 (O_758,N_49352,N_49200);
and UO_759 (O_759,N_49785,N_49205);
nand UO_760 (O_760,N_49978,N_49614);
nor UO_761 (O_761,N_49278,N_49964);
and UO_762 (O_762,N_49865,N_49986);
or UO_763 (O_763,N_49202,N_49905);
and UO_764 (O_764,N_49082,N_49791);
nor UO_765 (O_765,N_49451,N_49391);
nor UO_766 (O_766,N_49117,N_49154);
or UO_767 (O_767,N_49744,N_49636);
or UO_768 (O_768,N_49014,N_49889);
or UO_769 (O_769,N_49652,N_49072);
xnor UO_770 (O_770,N_49165,N_49907);
and UO_771 (O_771,N_49571,N_49306);
nand UO_772 (O_772,N_49785,N_49715);
nor UO_773 (O_773,N_49537,N_49077);
nor UO_774 (O_774,N_49455,N_49401);
xnor UO_775 (O_775,N_49412,N_49629);
and UO_776 (O_776,N_49724,N_49476);
and UO_777 (O_777,N_49471,N_49864);
xor UO_778 (O_778,N_49993,N_49828);
and UO_779 (O_779,N_49706,N_49107);
nor UO_780 (O_780,N_49817,N_49131);
nor UO_781 (O_781,N_49986,N_49075);
xnor UO_782 (O_782,N_49170,N_49845);
and UO_783 (O_783,N_49670,N_49193);
or UO_784 (O_784,N_49267,N_49956);
nand UO_785 (O_785,N_49828,N_49984);
nor UO_786 (O_786,N_49223,N_49210);
nor UO_787 (O_787,N_49398,N_49584);
xor UO_788 (O_788,N_49298,N_49882);
and UO_789 (O_789,N_49885,N_49983);
or UO_790 (O_790,N_49860,N_49598);
xnor UO_791 (O_791,N_49581,N_49677);
or UO_792 (O_792,N_49462,N_49610);
nand UO_793 (O_793,N_49525,N_49308);
or UO_794 (O_794,N_49275,N_49911);
or UO_795 (O_795,N_49214,N_49769);
xnor UO_796 (O_796,N_49058,N_49474);
nand UO_797 (O_797,N_49483,N_49672);
xnor UO_798 (O_798,N_49396,N_49921);
nor UO_799 (O_799,N_49161,N_49327);
nand UO_800 (O_800,N_49177,N_49857);
nand UO_801 (O_801,N_49848,N_49103);
xor UO_802 (O_802,N_49751,N_49850);
nand UO_803 (O_803,N_49858,N_49956);
nor UO_804 (O_804,N_49164,N_49023);
and UO_805 (O_805,N_49878,N_49089);
xnor UO_806 (O_806,N_49650,N_49880);
xor UO_807 (O_807,N_49791,N_49754);
and UO_808 (O_808,N_49104,N_49518);
xnor UO_809 (O_809,N_49376,N_49985);
nor UO_810 (O_810,N_49193,N_49388);
nor UO_811 (O_811,N_49716,N_49314);
xor UO_812 (O_812,N_49932,N_49509);
nand UO_813 (O_813,N_49875,N_49684);
xnor UO_814 (O_814,N_49742,N_49335);
xnor UO_815 (O_815,N_49095,N_49669);
or UO_816 (O_816,N_49799,N_49876);
or UO_817 (O_817,N_49426,N_49538);
or UO_818 (O_818,N_49019,N_49475);
or UO_819 (O_819,N_49222,N_49969);
nor UO_820 (O_820,N_49040,N_49484);
nor UO_821 (O_821,N_49643,N_49762);
or UO_822 (O_822,N_49196,N_49630);
xor UO_823 (O_823,N_49436,N_49097);
nor UO_824 (O_824,N_49344,N_49210);
or UO_825 (O_825,N_49284,N_49021);
nand UO_826 (O_826,N_49873,N_49932);
or UO_827 (O_827,N_49676,N_49970);
nand UO_828 (O_828,N_49191,N_49992);
or UO_829 (O_829,N_49557,N_49359);
xnor UO_830 (O_830,N_49126,N_49909);
or UO_831 (O_831,N_49431,N_49236);
xor UO_832 (O_832,N_49797,N_49942);
xor UO_833 (O_833,N_49332,N_49725);
or UO_834 (O_834,N_49730,N_49960);
xnor UO_835 (O_835,N_49460,N_49816);
or UO_836 (O_836,N_49859,N_49342);
xor UO_837 (O_837,N_49176,N_49272);
or UO_838 (O_838,N_49990,N_49433);
or UO_839 (O_839,N_49597,N_49331);
nor UO_840 (O_840,N_49358,N_49467);
and UO_841 (O_841,N_49144,N_49133);
and UO_842 (O_842,N_49963,N_49549);
and UO_843 (O_843,N_49405,N_49051);
and UO_844 (O_844,N_49884,N_49340);
xnor UO_845 (O_845,N_49792,N_49035);
and UO_846 (O_846,N_49154,N_49291);
nor UO_847 (O_847,N_49643,N_49901);
nor UO_848 (O_848,N_49991,N_49854);
xor UO_849 (O_849,N_49578,N_49959);
nor UO_850 (O_850,N_49183,N_49675);
nand UO_851 (O_851,N_49677,N_49244);
and UO_852 (O_852,N_49182,N_49392);
or UO_853 (O_853,N_49714,N_49302);
xor UO_854 (O_854,N_49067,N_49344);
nand UO_855 (O_855,N_49182,N_49661);
or UO_856 (O_856,N_49674,N_49805);
nor UO_857 (O_857,N_49114,N_49349);
and UO_858 (O_858,N_49642,N_49566);
xor UO_859 (O_859,N_49016,N_49680);
and UO_860 (O_860,N_49981,N_49148);
nand UO_861 (O_861,N_49535,N_49935);
nand UO_862 (O_862,N_49989,N_49455);
xor UO_863 (O_863,N_49948,N_49426);
nand UO_864 (O_864,N_49969,N_49061);
or UO_865 (O_865,N_49818,N_49639);
xor UO_866 (O_866,N_49312,N_49344);
xnor UO_867 (O_867,N_49181,N_49135);
nor UO_868 (O_868,N_49212,N_49601);
nor UO_869 (O_869,N_49222,N_49880);
nor UO_870 (O_870,N_49532,N_49795);
or UO_871 (O_871,N_49444,N_49824);
nor UO_872 (O_872,N_49297,N_49810);
nor UO_873 (O_873,N_49912,N_49465);
nand UO_874 (O_874,N_49759,N_49666);
or UO_875 (O_875,N_49348,N_49242);
and UO_876 (O_876,N_49590,N_49101);
nor UO_877 (O_877,N_49818,N_49117);
nor UO_878 (O_878,N_49248,N_49511);
or UO_879 (O_879,N_49954,N_49242);
nor UO_880 (O_880,N_49609,N_49598);
nor UO_881 (O_881,N_49872,N_49828);
and UO_882 (O_882,N_49709,N_49817);
nor UO_883 (O_883,N_49536,N_49103);
nand UO_884 (O_884,N_49135,N_49165);
or UO_885 (O_885,N_49982,N_49602);
and UO_886 (O_886,N_49282,N_49432);
xor UO_887 (O_887,N_49090,N_49126);
or UO_888 (O_888,N_49733,N_49101);
nor UO_889 (O_889,N_49639,N_49162);
and UO_890 (O_890,N_49285,N_49371);
nand UO_891 (O_891,N_49513,N_49279);
or UO_892 (O_892,N_49200,N_49673);
nand UO_893 (O_893,N_49722,N_49119);
and UO_894 (O_894,N_49845,N_49032);
and UO_895 (O_895,N_49034,N_49684);
xor UO_896 (O_896,N_49379,N_49947);
xnor UO_897 (O_897,N_49565,N_49073);
xnor UO_898 (O_898,N_49645,N_49707);
and UO_899 (O_899,N_49003,N_49276);
or UO_900 (O_900,N_49649,N_49995);
nand UO_901 (O_901,N_49342,N_49282);
and UO_902 (O_902,N_49845,N_49556);
and UO_903 (O_903,N_49065,N_49331);
nor UO_904 (O_904,N_49430,N_49381);
and UO_905 (O_905,N_49914,N_49093);
nand UO_906 (O_906,N_49742,N_49201);
nor UO_907 (O_907,N_49413,N_49321);
nor UO_908 (O_908,N_49740,N_49257);
or UO_909 (O_909,N_49737,N_49919);
nand UO_910 (O_910,N_49509,N_49448);
nand UO_911 (O_911,N_49040,N_49779);
nor UO_912 (O_912,N_49398,N_49191);
nand UO_913 (O_913,N_49505,N_49216);
and UO_914 (O_914,N_49061,N_49429);
xor UO_915 (O_915,N_49243,N_49943);
xnor UO_916 (O_916,N_49828,N_49673);
and UO_917 (O_917,N_49420,N_49101);
nor UO_918 (O_918,N_49562,N_49953);
xor UO_919 (O_919,N_49586,N_49730);
nor UO_920 (O_920,N_49594,N_49214);
or UO_921 (O_921,N_49440,N_49818);
and UO_922 (O_922,N_49172,N_49012);
nand UO_923 (O_923,N_49762,N_49132);
and UO_924 (O_924,N_49424,N_49174);
nand UO_925 (O_925,N_49224,N_49778);
nor UO_926 (O_926,N_49636,N_49078);
nand UO_927 (O_927,N_49009,N_49016);
nand UO_928 (O_928,N_49259,N_49324);
xnor UO_929 (O_929,N_49374,N_49083);
nor UO_930 (O_930,N_49727,N_49630);
and UO_931 (O_931,N_49863,N_49442);
nor UO_932 (O_932,N_49595,N_49132);
nor UO_933 (O_933,N_49771,N_49320);
and UO_934 (O_934,N_49533,N_49107);
or UO_935 (O_935,N_49085,N_49895);
or UO_936 (O_936,N_49480,N_49481);
xor UO_937 (O_937,N_49460,N_49070);
and UO_938 (O_938,N_49843,N_49879);
xnor UO_939 (O_939,N_49308,N_49194);
and UO_940 (O_940,N_49572,N_49952);
nor UO_941 (O_941,N_49883,N_49138);
xor UO_942 (O_942,N_49991,N_49310);
xnor UO_943 (O_943,N_49909,N_49502);
nor UO_944 (O_944,N_49455,N_49063);
nand UO_945 (O_945,N_49669,N_49106);
or UO_946 (O_946,N_49253,N_49842);
nand UO_947 (O_947,N_49716,N_49601);
xor UO_948 (O_948,N_49538,N_49888);
xnor UO_949 (O_949,N_49211,N_49164);
or UO_950 (O_950,N_49894,N_49509);
or UO_951 (O_951,N_49707,N_49499);
nor UO_952 (O_952,N_49119,N_49384);
or UO_953 (O_953,N_49852,N_49031);
nand UO_954 (O_954,N_49440,N_49999);
nand UO_955 (O_955,N_49443,N_49047);
nor UO_956 (O_956,N_49653,N_49403);
xor UO_957 (O_957,N_49148,N_49791);
nor UO_958 (O_958,N_49764,N_49743);
xor UO_959 (O_959,N_49462,N_49174);
nand UO_960 (O_960,N_49267,N_49924);
nand UO_961 (O_961,N_49031,N_49650);
nor UO_962 (O_962,N_49673,N_49589);
or UO_963 (O_963,N_49854,N_49105);
nor UO_964 (O_964,N_49492,N_49920);
nand UO_965 (O_965,N_49730,N_49258);
xnor UO_966 (O_966,N_49596,N_49209);
xor UO_967 (O_967,N_49348,N_49873);
xor UO_968 (O_968,N_49008,N_49713);
or UO_969 (O_969,N_49323,N_49706);
or UO_970 (O_970,N_49014,N_49463);
and UO_971 (O_971,N_49557,N_49516);
xnor UO_972 (O_972,N_49802,N_49586);
or UO_973 (O_973,N_49247,N_49733);
or UO_974 (O_974,N_49508,N_49480);
and UO_975 (O_975,N_49195,N_49846);
xor UO_976 (O_976,N_49404,N_49545);
nor UO_977 (O_977,N_49723,N_49228);
and UO_978 (O_978,N_49725,N_49442);
nor UO_979 (O_979,N_49181,N_49359);
or UO_980 (O_980,N_49225,N_49006);
nor UO_981 (O_981,N_49416,N_49876);
nand UO_982 (O_982,N_49883,N_49170);
and UO_983 (O_983,N_49795,N_49252);
xnor UO_984 (O_984,N_49861,N_49862);
and UO_985 (O_985,N_49735,N_49254);
nor UO_986 (O_986,N_49755,N_49266);
or UO_987 (O_987,N_49420,N_49428);
or UO_988 (O_988,N_49356,N_49610);
nor UO_989 (O_989,N_49271,N_49144);
nor UO_990 (O_990,N_49112,N_49957);
xnor UO_991 (O_991,N_49000,N_49050);
xor UO_992 (O_992,N_49297,N_49273);
nor UO_993 (O_993,N_49815,N_49204);
and UO_994 (O_994,N_49519,N_49844);
and UO_995 (O_995,N_49009,N_49152);
nor UO_996 (O_996,N_49293,N_49698);
or UO_997 (O_997,N_49814,N_49550);
and UO_998 (O_998,N_49065,N_49214);
nand UO_999 (O_999,N_49889,N_49452);
nand UO_1000 (O_1000,N_49229,N_49636);
or UO_1001 (O_1001,N_49395,N_49999);
and UO_1002 (O_1002,N_49265,N_49203);
xnor UO_1003 (O_1003,N_49633,N_49238);
nor UO_1004 (O_1004,N_49737,N_49325);
and UO_1005 (O_1005,N_49339,N_49199);
or UO_1006 (O_1006,N_49536,N_49070);
xnor UO_1007 (O_1007,N_49234,N_49059);
or UO_1008 (O_1008,N_49580,N_49044);
or UO_1009 (O_1009,N_49496,N_49709);
xnor UO_1010 (O_1010,N_49336,N_49704);
or UO_1011 (O_1011,N_49737,N_49814);
nand UO_1012 (O_1012,N_49364,N_49528);
or UO_1013 (O_1013,N_49068,N_49693);
nand UO_1014 (O_1014,N_49218,N_49990);
or UO_1015 (O_1015,N_49558,N_49938);
nand UO_1016 (O_1016,N_49576,N_49463);
xor UO_1017 (O_1017,N_49788,N_49563);
xnor UO_1018 (O_1018,N_49949,N_49861);
or UO_1019 (O_1019,N_49124,N_49472);
nand UO_1020 (O_1020,N_49623,N_49640);
nor UO_1021 (O_1021,N_49446,N_49598);
xor UO_1022 (O_1022,N_49275,N_49828);
nand UO_1023 (O_1023,N_49049,N_49323);
and UO_1024 (O_1024,N_49336,N_49920);
and UO_1025 (O_1025,N_49624,N_49487);
nand UO_1026 (O_1026,N_49020,N_49300);
and UO_1027 (O_1027,N_49620,N_49923);
and UO_1028 (O_1028,N_49992,N_49587);
or UO_1029 (O_1029,N_49711,N_49386);
nand UO_1030 (O_1030,N_49033,N_49694);
nand UO_1031 (O_1031,N_49697,N_49872);
or UO_1032 (O_1032,N_49315,N_49264);
and UO_1033 (O_1033,N_49877,N_49201);
xor UO_1034 (O_1034,N_49005,N_49559);
xor UO_1035 (O_1035,N_49959,N_49852);
nor UO_1036 (O_1036,N_49093,N_49720);
nand UO_1037 (O_1037,N_49191,N_49763);
xnor UO_1038 (O_1038,N_49402,N_49889);
nand UO_1039 (O_1039,N_49641,N_49925);
and UO_1040 (O_1040,N_49811,N_49075);
xnor UO_1041 (O_1041,N_49231,N_49841);
and UO_1042 (O_1042,N_49869,N_49918);
or UO_1043 (O_1043,N_49349,N_49948);
or UO_1044 (O_1044,N_49028,N_49612);
nand UO_1045 (O_1045,N_49920,N_49382);
xor UO_1046 (O_1046,N_49396,N_49755);
nand UO_1047 (O_1047,N_49813,N_49664);
nor UO_1048 (O_1048,N_49671,N_49223);
and UO_1049 (O_1049,N_49241,N_49452);
and UO_1050 (O_1050,N_49698,N_49450);
xnor UO_1051 (O_1051,N_49637,N_49203);
or UO_1052 (O_1052,N_49013,N_49569);
or UO_1053 (O_1053,N_49245,N_49050);
and UO_1054 (O_1054,N_49382,N_49518);
and UO_1055 (O_1055,N_49753,N_49213);
nor UO_1056 (O_1056,N_49686,N_49343);
nand UO_1057 (O_1057,N_49027,N_49571);
xnor UO_1058 (O_1058,N_49436,N_49651);
or UO_1059 (O_1059,N_49793,N_49877);
xnor UO_1060 (O_1060,N_49293,N_49525);
or UO_1061 (O_1061,N_49626,N_49638);
nand UO_1062 (O_1062,N_49859,N_49210);
and UO_1063 (O_1063,N_49241,N_49974);
xor UO_1064 (O_1064,N_49477,N_49547);
and UO_1065 (O_1065,N_49084,N_49700);
xnor UO_1066 (O_1066,N_49626,N_49778);
xnor UO_1067 (O_1067,N_49060,N_49294);
or UO_1068 (O_1068,N_49441,N_49806);
nor UO_1069 (O_1069,N_49820,N_49627);
and UO_1070 (O_1070,N_49903,N_49755);
xor UO_1071 (O_1071,N_49578,N_49912);
xnor UO_1072 (O_1072,N_49258,N_49731);
xor UO_1073 (O_1073,N_49515,N_49238);
nor UO_1074 (O_1074,N_49182,N_49147);
or UO_1075 (O_1075,N_49530,N_49637);
and UO_1076 (O_1076,N_49536,N_49852);
nand UO_1077 (O_1077,N_49376,N_49335);
nand UO_1078 (O_1078,N_49640,N_49531);
or UO_1079 (O_1079,N_49006,N_49775);
nand UO_1080 (O_1080,N_49349,N_49077);
or UO_1081 (O_1081,N_49289,N_49947);
nor UO_1082 (O_1082,N_49926,N_49947);
or UO_1083 (O_1083,N_49691,N_49278);
nor UO_1084 (O_1084,N_49967,N_49013);
and UO_1085 (O_1085,N_49954,N_49277);
nand UO_1086 (O_1086,N_49138,N_49390);
or UO_1087 (O_1087,N_49564,N_49363);
and UO_1088 (O_1088,N_49068,N_49154);
and UO_1089 (O_1089,N_49508,N_49288);
nor UO_1090 (O_1090,N_49079,N_49678);
and UO_1091 (O_1091,N_49162,N_49373);
or UO_1092 (O_1092,N_49573,N_49435);
nand UO_1093 (O_1093,N_49177,N_49420);
nand UO_1094 (O_1094,N_49639,N_49902);
nand UO_1095 (O_1095,N_49088,N_49145);
nor UO_1096 (O_1096,N_49790,N_49725);
nor UO_1097 (O_1097,N_49183,N_49118);
or UO_1098 (O_1098,N_49218,N_49266);
or UO_1099 (O_1099,N_49650,N_49575);
xor UO_1100 (O_1100,N_49675,N_49148);
nand UO_1101 (O_1101,N_49927,N_49552);
nand UO_1102 (O_1102,N_49394,N_49782);
nand UO_1103 (O_1103,N_49734,N_49847);
xor UO_1104 (O_1104,N_49746,N_49271);
nor UO_1105 (O_1105,N_49055,N_49548);
xor UO_1106 (O_1106,N_49700,N_49755);
nor UO_1107 (O_1107,N_49510,N_49095);
nor UO_1108 (O_1108,N_49727,N_49607);
nor UO_1109 (O_1109,N_49637,N_49385);
nand UO_1110 (O_1110,N_49826,N_49505);
nand UO_1111 (O_1111,N_49051,N_49856);
or UO_1112 (O_1112,N_49326,N_49244);
or UO_1113 (O_1113,N_49526,N_49286);
xor UO_1114 (O_1114,N_49931,N_49153);
nor UO_1115 (O_1115,N_49825,N_49287);
nand UO_1116 (O_1116,N_49939,N_49221);
xnor UO_1117 (O_1117,N_49793,N_49633);
or UO_1118 (O_1118,N_49473,N_49963);
nor UO_1119 (O_1119,N_49579,N_49490);
xnor UO_1120 (O_1120,N_49832,N_49171);
xor UO_1121 (O_1121,N_49851,N_49380);
nand UO_1122 (O_1122,N_49613,N_49727);
or UO_1123 (O_1123,N_49026,N_49985);
or UO_1124 (O_1124,N_49538,N_49368);
and UO_1125 (O_1125,N_49985,N_49021);
or UO_1126 (O_1126,N_49240,N_49729);
or UO_1127 (O_1127,N_49511,N_49807);
or UO_1128 (O_1128,N_49082,N_49387);
nor UO_1129 (O_1129,N_49425,N_49766);
nand UO_1130 (O_1130,N_49856,N_49643);
and UO_1131 (O_1131,N_49810,N_49606);
nor UO_1132 (O_1132,N_49418,N_49858);
nand UO_1133 (O_1133,N_49653,N_49396);
nor UO_1134 (O_1134,N_49210,N_49173);
nand UO_1135 (O_1135,N_49051,N_49940);
nand UO_1136 (O_1136,N_49957,N_49016);
nand UO_1137 (O_1137,N_49461,N_49063);
xor UO_1138 (O_1138,N_49877,N_49433);
nand UO_1139 (O_1139,N_49219,N_49740);
nor UO_1140 (O_1140,N_49502,N_49833);
or UO_1141 (O_1141,N_49043,N_49706);
and UO_1142 (O_1142,N_49027,N_49058);
nand UO_1143 (O_1143,N_49712,N_49111);
and UO_1144 (O_1144,N_49692,N_49960);
nand UO_1145 (O_1145,N_49133,N_49074);
or UO_1146 (O_1146,N_49661,N_49278);
or UO_1147 (O_1147,N_49910,N_49965);
xnor UO_1148 (O_1148,N_49853,N_49800);
and UO_1149 (O_1149,N_49960,N_49257);
xor UO_1150 (O_1150,N_49948,N_49097);
nand UO_1151 (O_1151,N_49589,N_49999);
and UO_1152 (O_1152,N_49949,N_49856);
and UO_1153 (O_1153,N_49794,N_49241);
nand UO_1154 (O_1154,N_49955,N_49995);
and UO_1155 (O_1155,N_49860,N_49045);
nor UO_1156 (O_1156,N_49887,N_49842);
nor UO_1157 (O_1157,N_49472,N_49338);
xnor UO_1158 (O_1158,N_49312,N_49122);
nand UO_1159 (O_1159,N_49085,N_49797);
or UO_1160 (O_1160,N_49204,N_49037);
and UO_1161 (O_1161,N_49428,N_49905);
xor UO_1162 (O_1162,N_49021,N_49794);
nor UO_1163 (O_1163,N_49625,N_49958);
and UO_1164 (O_1164,N_49978,N_49567);
or UO_1165 (O_1165,N_49265,N_49929);
and UO_1166 (O_1166,N_49644,N_49157);
and UO_1167 (O_1167,N_49351,N_49989);
and UO_1168 (O_1168,N_49364,N_49618);
xor UO_1169 (O_1169,N_49630,N_49195);
and UO_1170 (O_1170,N_49128,N_49954);
and UO_1171 (O_1171,N_49394,N_49894);
nor UO_1172 (O_1172,N_49964,N_49452);
or UO_1173 (O_1173,N_49095,N_49793);
nor UO_1174 (O_1174,N_49585,N_49411);
xor UO_1175 (O_1175,N_49555,N_49433);
nand UO_1176 (O_1176,N_49304,N_49025);
xor UO_1177 (O_1177,N_49950,N_49965);
nor UO_1178 (O_1178,N_49079,N_49129);
nand UO_1179 (O_1179,N_49315,N_49558);
nand UO_1180 (O_1180,N_49147,N_49511);
nor UO_1181 (O_1181,N_49560,N_49769);
nand UO_1182 (O_1182,N_49535,N_49247);
xor UO_1183 (O_1183,N_49521,N_49607);
nor UO_1184 (O_1184,N_49277,N_49153);
and UO_1185 (O_1185,N_49076,N_49810);
or UO_1186 (O_1186,N_49670,N_49977);
nor UO_1187 (O_1187,N_49059,N_49080);
nor UO_1188 (O_1188,N_49551,N_49071);
and UO_1189 (O_1189,N_49316,N_49500);
xnor UO_1190 (O_1190,N_49017,N_49411);
and UO_1191 (O_1191,N_49890,N_49560);
or UO_1192 (O_1192,N_49324,N_49160);
or UO_1193 (O_1193,N_49934,N_49920);
xnor UO_1194 (O_1194,N_49722,N_49384);
xnor UO_1195 (O_1195,N_49246,N_49643);
xor UO_1196 (O_1196,N_49736,N_49340);
or UO_1197 (O_1197,N_49259,N_49148);
xnor UO_1198 (O_1198,N_49591,N_49161);
and UO_1199 (O_1199,N_49006,N_49033);
and UO_1200 (O_1200,N_49335,N_49437);
nand UO_1201 (O_1201,N_49516,N_49682);
and UO_1202 (O_1202,N_49428,N_49340);
nor UO_1203 (O_1203,N_49024,N_49246);
nand UO_1204 (O_1204,N_49348,N_49594);
or UO_1205 (O_1205,N_49192,N_49629);
nor UO_1206 (O_1206,N_49807,N_49516);
or UO_1207 (O_1207,N_49446,N_49558);
or UO_1208 (O_1208,N_49866,N_49506);
xnor UO_1209 (O_1209,N_49106,N_49308);
or UO_1210 (O_1210,N_49782,N_49303);
nor UO_1211 (O_1211,N_49828,N_49849);
or UO_1212 (O_1212,N_49515,N_49226);
xnor UO_1213 (O_1213,N_49346,N_49154);
nand UO_1214 (O_1214,N_49931,N_49796);
nand UO_1215 (O_1215,N_49854,N_49615);
and UO_1216 (O_1216,N_49639,N_49343);
nor UO_1217 (O_1217,N_49142,N_49511);
or UO_1218 (O_1218,N_49359,N_49146);
xnor UO_1219 (O_1219,N_49935,N_49537);
xor UO_1220 (O_1220,N_49421,N_49839);
xnor UO_1221 (O_1221,N_49972,N_49487);
and UO_1222 (O_1222,N_49683,N_49161);
xor UO_1223 (O_1223,N_49529,N_49979);
nand UO_1224 (O_1224,N_49929,N_49270);
and UO_1225 (O_1225,N_49544,N_49665);
xor UO_1226 (O_1226,N_49752,N_49948);
and UO_1227 (O_1227,N_49042,N_49737);
and UO_1228 (O_1228,N_49057,N_49370);
nor UO_1229 (O_1229,N_49799,N_49734);
and UO_1230 (O_1230,N_49508,N_49583);
nor UO_1231 (O_1231,N_49690,N_49645);
and UO_1232 (O_1232,N_49568,N_49113);
xnor UO_1233 (O_1233,N_49295,N_49613);
xor UO_1234 (O_1234,N_49407,N_49177);
xor UO_1235 (O_1235,N_49153,N_49168);
and UO_1236 (O_1236,N_49055,N_49693);
nor UO_1237 (O_1237,N_49218,N_49510);
xnor UO_1238 (O_1238,N_49277,N_49473);
nor UO_1239 (O_1239,N_49095,N_49568);
or UO_1240 (O_1240,N_49204,N_49467);
and UO_1241 (O_1241,N_49040,N_49434);
nand UO_1242 (O_1242,N_49320,N_49967);
or UO_1243 (O_1243,N_49594,N_49756);
nor UO_1244 (O_1244,N_49130,N_49021);
nor UO_1245 (O_1245,N_49719,N_49079);
nand UO_1246 (O_1246,N_49207,N_49861);
or UO_1247 (O_1247,N_49073,N_49659);
xnor UO_1248 (O_1248,N_49398,N_49439);
nor UO_1249 (O_1249,N_49556,N_49411);
nand UO_1250 (O_1250,N_49998,N_49810);
xnor UO_1251 (O_1251,N_49751,N_49919);
or UO_1252 (O_1252,N_49835,N_49961);
xnor UO_1253 (O_1253,N_49132,N_49663);
nor UO_1254 (O_1254,N_49586,N_49527);
and UO_1255 (O_1255,N_49508,N_49352);
or UO_1256 (O_1256,N_49613,N_49222);
xnor UO_1257 (O_1257,N_49922,N_49504);
and UO_1258 (O_1258,N_49280,N_49037);
nor UO_1259 (O_1259,N_49016,N_49248);
nor UO_1260 (O_1260,N_49683,N_49343);
xor UO_1261 (O_1261,N_49941,N_49468);
nand UO_1262 (O_1262,N_49601,N_49790);
and UO_1263 (O_1263,N_49274,N_49146);
or UO_1264 (O_1264,N_49146,N_49880);
nand UO_1265 (O_1265,N_49887,N_49140);
or UO_1266 (O_1266,N_49401,N_49630);
nand UO_1267 (O_1267,N_49937,N_49518);
xnor UO_1268 (O_1268,N_49917,N_49399);
nand UO_1269 (O_1269,N_49905,N_49330);
nor UO_1270 (O_1270,N_49131,N_49708);
and UO_1271 (O_1271,N_49952,N_49595);
and UO_1272 (O_1272,N_49645,N_49593);
nand UO_1273 (O_1273,N_49009,N_49865);
and UO_1274 (O_1274,N_49169,N_49282);
and UO_1275 (O_1275,N_49622,N_49371);
xor UO_1276 (O_1276,N_49312,N_49667);
nand UO_1277 (O_1277,N_49257,N_49947);
or UO_1278 (O_1278,N_49877,N_49410);
and UO_1279 (O_1279,N_49308,N_49686);
nor UO_1280 (O_1280,N_49559,N_49713);
nor UO_1281 (O_1281,N_49377,N_49856);
and UO_1282 (O_1282,N_49547,N_49458);
xor UO_1283 (O_1283,N_49433,N_49223);
and UO_1284 (O_1284,N_49211,N_49136);
xor UO_1285 (O_1285,N_49321,N_49627);
nand UO_1286 (O_1286,N_49780,N_49754);
or UO_1287 (O_1287,N_49821,N_49043);
and UO_1288 (O_1288,N_49947,N_49596);
or UO_1289 (O_1289,N_49370,N_49893);
or UO_1290 (O_1290,N_49161,N_49991);
or UO_1291 (O_1291,N_49747,N_49698);
nand UO_1292 (O_1292,N_49418,N_49785);
or UO_1293 (O_1293,N_49530,N_49976);
nand UO_1294 (O_1294,N_49401,N_49224);
nor UO_1295 (O_1295,N_49128,N_49682);
or UO_1296 (O_1296,N_49951,N_49688);
and UO_1297 (O_1297,N_49549,N_49739);
nand UO_1298 (O_1298,N_49787,N_49795);
nand UO_1299 (O_1299,N_49031,N_49373);
nor UO_1300 (O_1300,N_49492,N_49628);
or UO_1301 (O_1301,N_49712,N_49754);
nor UO_1302 (O_1302,N_49121,N_49817);
and UO_1303 (O_1303,N_49792,N_49972);
nand UO_1304 (O_1304,N_49593,N_49919);
or UO_1305 (O_1305,N_49999,N_49718);
nor UO_1306 (O_1306,N_49942,N_49281);
nand UO_1307 (O_1307,N_49307,N_49577);
nand UO_1308 (O_1308,N_49149,N_49322);
and UO_1309 (O_1309,N_49463,N_49309);
or UO_1310 (O_1310,N_49395,N_49438);
and UO_1311 (O_1311,N_49015,N_49130);
and UO_1312 (O_1312,N_49190,N_49895);
nand UO_1313 (O_1313,N_49146,N_49314);
nand UO_1314 (O_1314,N_49655,N_49661);
xnor UO_1315 (O_1315,N_49103,N_49107);
or UO_1316 (O_1316,N_49768,N_49920);
xnor UO_1317 (O_1317,N_49226,N_49310);
or UO_1318 (O_1318,N_49944,N_49913);
or UO_1319 (O_1319,N_49005,N_49476);
or UO_1320 (O_1320,N_49772,N_49927);
xor UO_1321 (O_1321,N_49874,N_49727);
xnor UO_1322 (O_1322,N_49758,N_49769);
nor UO_1323 (O_1323,N_49525,N_49978);
and UO_1324 (O_1324,N_49838,N_49506);
and UO_1325 (O_1325,N_49221,N_49177);
nand UO_1326 (O_1326,N_49375,N_49139);
or UO_1327 (O_1327,N_49808,N_49964);
nand UO_1328 (O_1328,N_49980,N_49412);
and UO_1329 (O_1329,N_49439,N_49498);
xor UO_1330 (O_1330,N_49578,N_49371);
or UO_1331 (O_1331,N_49067,N_49782);
nor UO_1332 (O_1332,N_49665,N_49894);
or UO_1333 (O_1333,N_49041,N_49981);
nand UO_1334 (O_1334,N_49185,N_49848);
nand UO_1335 (O_1335,N_49881,N_49530);
or UO_1336 (O_1336,N_49564,N_49763);
xor UO_1337 (O_1337,N_49171,N_49813);
xnor UO_1338 (O_1338,N_49835,N_49663);
or UO_1339 (O_1339,N_49259,N_49323);
or UO_1340 (O_1340,N_49629,N_49390);
nor UO_1341 (O_1341,N_49651,N_49663);
nor UO_1342 (O_1342,N_49447,N_49668);
nor UO_1343 (O_1343,N_49996,N_49327);
and UO_1344 (O_1344,N_49884,N_49560);
nand UO_1345 (O_1345,N_49787,N_49710);
or UO_1346 (O_1346,N_49585,N_49710);
or UO_1347 (O_1347,N_49215,N_49172);
nor UO_1348 (O_1348,N_49435,N_49554);
nand UO_1349 (O_1349,N_49391,N_49747);
xor UO_1350 (O_1350,N_49489,N_49430);
and UO_1351 (O_1351,N_49615,N_49933);
xor UO_1352 (O_1352,N_49199,N_49738);
xor UO_1353 (O_1353,N_49083,N_49890);
nor UO_1354 (O_1354,N_49025,N_49356);
nand UO_1355 (O_1355,N_49919,N_49249);
nor UO_1356 (O_1356,N_49902,N_49439);
or UO_1357 (O_1357,N_49937,N_49642);
nor UO_1358 (O_1358,N_49074,N_49248);
or UO_1359 (O_1359,N_49778,N_49693);
nand UO_1360 (O_1360,N_49614,N_49590);
xnor UO_1361 (O_1361,N_49014,N_49286);
or UO_1362 (O_1362,N_49483,N_49811);
and UO_1363 (O_1363,N_49731,N_49855);
nor UO_1364 (O_1364,N_49426,N_49838);
and UO_1365 (O_1365,N_49878,N_49023);
and UO_1366 (O_1366,N_49919,N_49145);
xnor UO_1367 (O_1367,N_49571,N_49509);
xnor UO_1368 (O_1368,N_49151,N_49610);
and UO_1369 (O_1369,N_49164,N_49751);
and UO_1370 (O_1370,N_49332,N_49705);
nor UO_1371 (O_1371,N_49539,N_49736);
and UO_1372 (O_1372,N_49694,N_49906);
and UO_1373 (O_1373,N_49392,N_49473);
xor UO_1374 (O_1374,N_49596,N_49671);
nor UO_1375 (O_1375,N_49297,N_49153);
or UO_1376 (O_1376,N_49367,N_49225);
nor UO_1377 (O_1377,N_49178,N_49012);
nand UO_1378 (O_1378,N_49700,N_49608);
nand UO_1379 (O_1379,N_49108,N_49774);
nor UO_1380 (O_1380,N_49705,N_49310);
nand UO_1381 (O_1381,N_49849,N_49210);
or UO_1382 (O_1382,N_49745,N_49281);
and UO_1383 (O_1383,N_49455,N_49101);
nand UO_1384 (O_1384,N_49145,N_49713);
nand UO_1385 (O_1385,N_49639,N_49424);
or UO_1386 (O_1386,N_49524,N_49954);
and UO_1387 (O_1387,N_49531,N_49589);
and UO_1388 (O_1388,N_49092,N_49367);
and UO_1389 (O_1389,N_49805,N_49559);
and UO_1390 (O_1390,N_49679,N_49482);
nand UO_1391 (O_1391,N_49864,N_49138);
nor UO_1392 (O_1392,N_49753,N_49405);
nor UO_1393 (O_1393,N_49290,N_49031);
xnor UO_1394 (O_1394,N_49959,N_49246);
nor UO_1395 (O_1395,N_49236,N_49701);
and UO_1396 (O_1396,N_49778,N_49868);
and UO_1397 (O_1397,N_49004,N_49785);
or UO_1398 (O_1398,N_49982,N_49320);
nand UO_1399 (O_1399,N_49030,N_49510);
nand UO_1400 (O_1400,N_49467,N_49935);
and UO_1401 (O_1401,N_49767,N_49841);
and UO_1402 (O_1402,N_49256,N_49514);
or UO_1403 (O_1403,N_49744,N_49763);
nand UO_1404 (O_1404,N_49027,N_49043);
or UO_1405 (O_1405,N_49211,N_49370);
xor UO_1406 (O_1406,N_49884,N_49896);
xnor UO_1407 (O_1407,N_49546,N_49637);
and UO_1408 (O_1408,N_49905,N_49628);
xor UO_1409 (O_1409,N_49866,N_49334);
xnor UO_1410 (O_1410,N_49893,N_49082);
xor UO_1411 (O_1411,N_49858,N_49016);
xnor UO_1412 (O_1412,N_49997,N_49736);
or UO_1413 (O_1413,N_49243,N_49904);
nand UO_1414 (O_1414,N_49757,N_49861);
nand UO_1415 (O_1415,N_49501,N_49975);
or UO_1416 (O_1416,N_49744,N_49488);
or UO_1417 (O_1417,N_49886,N_49996);
nor UO_1418 (O_1418,N_49245,N_49942);
and UO_1419 (O_1419,N_49799,N_49546);
nor UO_1420 (O_1420,N_49535,N_49845);
or UO_1421 (O_1421,N_49177,N_49687);
and UO_1422 (O_1422,N_49638,N_49755);
and UO_1423 (O_1423,N_49424,N_49745);
xnor UO_1424 (O_1424,N_49084,N_49738);
or UO_1425 (O_1425,N_49948,N_49135);
nor UO_1426 (O_1426,N_49116,N_49331);
nor UO_1427 (O_1427,N_49812,N_49539);
nand UO_1428 (O_1428,N_49587,N_49229);
or UO_1429 (O_1429,N_49752,N_49743);
nor UO_1430 (O_1430,N_49199,N_49321);
nand UO_1431 (O_1431,N_49652,N_49622);
and UO_1432 (O_1432,N_49646,N_49051);
or UO_1433 (O_1433,N_49462,N_49742);
nor UO_1434 (O_1434,N_49565,N_49263);
or UO_1435 (O_1435,N_49618,N_49490);
xnor UO_1436 (O_1436,N_49240,N_49740);
nand UO_1437 (O_1437,N_49850,N_49975);
and UO_1438 (O_1438,N_49834,N_49581);
nor UO_1439 (O_1439,N_49889,N_49176);
and UO_1440 (O_1440,N_49886,N_49729);
or UO_1441 (O_1441,N_49609,N_49800);
or UO_1442 (O_1442,N_49553,N_49280);
and UO_1443 (O_1443,N_49055,N_49509);
xnor UO_1444 (O_1444,N_49603,N_49883);
and UO_1445 (O_1445,N_49835,N_49268);
or UO_1446 (O_1446,N_49935,N_49143);
nand UO_1447 (O_1447,N_49126,N_49952);
nor UO_1448 (O_1448,N_49724,N_49360);
and UO_1449 (O_1449,N_49394,N_49485);
nand UO_1450 (O_1450,N_49615,N_49164);
or UO_1451 (O_1451,N_49885,N_49246);
nand UO_1452 (O_1452,N_49634,N_49118);
nor UO_1453 (O_1453,N_49427,N_49308);
and UO_1454 (O_1454,N_49647,N_49531);
and UO_1455 (O_1455,N_49773,N_49327);
and UO_1456 (O_1456,N_49137,N_49756);
nand UO_1457 (O_1457,N_49003,N_49261);
nand UO_1458 (O_1458,N_49026,N_49680);
and UO_1459 (O_1459,N_49013,N_49902);
and UO_1460 (O_1460,N_49617,N_49215);
nand UO_1461 (O_1461,N_49410,N_49226);
nor UO_1462 (O_1462,N_49236,N_49984);
xnor UO_1463 (O_1463,N_49282,N_49024);
xor UO_1464 (O_1464,N_49128,N_49079);
xor UO_1465 (O_1465,N_49239,N_49412);
and UO_1466 (O_1466,N_49887,N_49029);
and UO_1467 (O_1467,N_49990,N_49892);
nand UO_1468 (O_1468,N_49622,N_49327);
xor UO_1469 (O_1469,N_49513,N_49272);
xor UO_1470 (O_1470,N_49887,N_49847);
or UO_1471 (O_1471,N_49120,N_49818);
and UO_1472 (O_1472,N_49529,N_49074);
and UO_1473 (O_1473,N_49394,N_49292);
nand UO_1474 (O_1474,N_49856,N_49801);
and UO_1475 (O_1475,N_49119,N_49332);
or UO_1476 (O_1476,N_49779,N_49096);
xnor UO_1477 (O_1477,N_49353,N_49542);
and UO_1478 (O_1478,N_49759,N_49343);
xnor UO_1479 (O_1479,N_49676,N_49195);
or UO_1480 (O_1480,N_49114,N_49000);
and UO_1481 (O_1481,N_49021,N_49568);
nand UO_1482 (O_1482,N_49299,N_49252);
or UO_1483 (O_1483,N_49713,N_49973);
xnor UO_1484 (O_1484,N_49864,N_49408);
xnor UO_1485 (O_1485,N_49397,N_49425);
xnor UO_1486 (O_1486,N_49618,N_49571);
xor UO_1487 (O_1487,N_49663,N_49197);
nand UO_1488 (O_1488,N_49114,N_49506);
and UO_1489 (O_1489,N_49413,N_49846);
and UO_1490 (O_1490,N_49194,N_49553);
and UO_1491 (O_1491,N_49535,N_49212);
or UO_1492 (O_1492,N_49931,N_49290);
and UO_1493 (O_1493,N_49367,N_49593);
nand UO_1494 (O_1494,N_49407,N_49052);
nor UO_1495 (O_1495,N_49863,N_49424);
or UO_1496 (O_1496,N_49122,N_49796);
or UO_1497 (O_1497,N_49015,N_49694);
nor UO_1498 (O_1498,N_49392,N_49303);
nor UO_1499 (O_1499,N_49181,N_49416);
xor UO_1500 (O_1500,N_49019,N_49451);
nand UO_1501 (O_1501,N_49078,N_49895);
xor UO_1502 (O_1502,N_49848,N_49548);
or UO_1503 (O_1503,N_49174,N_49560);
and UO_1504 (O_1504,N_49562,N_49445);
or UO_1505 (O_1505,N_49124,N_49482);
xnor UO_1506 (O_1506,N_49702,N_49534);
and UO_1507 (O_1507,N_49652,N_49132);
and UO_1508 (O_1508,N_49943,N_49245);
nor UO_1509 (O_1509,N_49648,N_49556);
xnor UO_1510 (O_1510,N_49974,N_49485);
or UO_1511 (O_1511,N_49026,N_49307);
nor UO_1512 (O_1512,N_49018,N_49745);
and UO_1513 (O_1513,N_49188,N_49532);
xor UO_1514 (O_1514,N_49922,N_49825);
nand UO_1515 (O_1515,N_49359,N_49262);
nor UO_1516 (O_1516,N_49367,N_49028);
nor UO_1517 (O_1517,N_49694,N_49459);
and UO_1518 (O_1518,N_49710,N_49503);
xnor UO_1519 (O_1519,N_49063,N_49326);
or UO_1520 (O_1520,N_49631,N_49930);
or UO_1521 (O_1521,N_49005,N_49946);
xnor UO_1522 (O_1522,N_49831,N_49365);
xnor UO_1523 (O_1523,N_49879,N_49802);
xor UO_1524 (O_1524,N_49098,N_49975);
or UO_1525 (O_1525,N_49604,N_49553);
or UO_1526 (O_1526,N_49005,N_49588);
nand UO_1527 (O_1527,N_49005,N_49312);
and UO_1528 (O_1528,N_49798,N_49955);
nand UO_1529 (O_1529,N_49101,N_49125);
nand UO_1530 (O_1530,N_49915,N_49675);
xor UO_1531 (O_1531,N_49082,N_49430);
nand UO_1532 (O_1532,N_49633,N_49237);
nand UO_1533 (O_1533,N_49620,N_49694);
or UO_1534 (O_1534,N_49815,N_49629);
nor UO_1535 (O_1535,N_49166,N_49563);
nor UO_1536 (O_1536,N_49060,N_49559);
xnor UO_1537 (O_1537,N_49881,N_49085);
or UO_1538 (O_1538,N_49007,N_49129);
and UO_1539 (O_1539,N_49643,N_49275);
or UO_1540 (O_1540,N_49660,N_49697);
or UO_1541 (O_1541,N_49956,N_49840);
nor UO_1542 (O_1542,N_49955,N_49423);
nor UO_1543 (O_1543,N_49765,N_49241);
nor UO_1544 (O_1544,N_49096,N_49158);
nand UO_1545 (O_1545,N_49696,N_49550);
xor UO_1546 (O_1546,N_49333,N_49357);
xnor UO_1547 (O_1547,N_49343,N_49381);
nand UO_1548 (O_1548,N_49099,N_49228);
xor UO_1549 (O_1549,N_49617,N_49485);
nor UO_1550 (O_1550,N_49216,N_49011);
and UO_1551 (O_1551,N_49522,N_49484);
nor UO_1552 (O_1552,N_49450,N_49400);
nor UO_1553 (O_1553,N_49837,N_49926);
nor UO_1554 (O_1554,N_49397,N_49231);
xnor UO_1555 (O_1555,N_49451,N_49067);
and UO_1556 (O_1556,N_49826,N_49388);
xnor UO_1557 (O_1557,N_49892,N_49009);
xnor UO_1558 (O_1558,N_49151,N_49713);
and UO_1559 (O_1559,N_49044,N_49490);
or UO_1560 (O_1560,N_49524,N_49557);
and UO_1561 (O_1561,N_49260,N_49937);
nand UO_1562 (O_1562,N_49066,N_49617);
xnor UO_1563 (O_1563,N_49262,N_49444);
and UO_1564 (O_1564,N_49636,N_49186);
or UO_1565 (O_1565,N_49965,N_49886);
nor UO_1566 (O_1566,N_49308,N_49147);
or UO_1567 (O_1567,N_49008,N_49280);
xor UO_1568 (O_1568,N_49642,N_49402);
nor UO_1569 (O_1569,N_49795,N_49290);
xnor UO_1570 (O_1570,N_49557,N_49038);
and UO_1571 (O_1571,N_49953,N_49651);
nor UO_1572 (O_1572,N_49068,N_49403);
xor UO_1573 (O_1573,N_49974,N_49687);
or UO_1574 (O_1574,N_49248,N_49387);
and UO_1575 (O_1575,N_49316,N_49280);
nor UO_1576 (O_1576,N_49959,N_49298);
xnor UO_1577 (O_1577,N_49753,N_49612);
xor UO_1578 (O_1578,N_49873,N_49463);
nor UO_1579 (O_1579,N_49339,N_49002);
nand UO_1580 (O_1580,N_49020,N_49988);
nor UO_1581 (O_1581,N_49607,N_49145);
nand UO_1582 (O_1582,N_49071,N_49224);
nand UO_1583 (O_1583,N_49185,N_49774);
nand UO_1584 (O_1584,N_49828,N_49472);
nand UO_1585 (O_1585,N_49093,N_49778);
or UO_1586 (O_1586,N_49508,N_49874);
nand UO_1587 (O_1587,N_49119,N_49334);
and UO_1588 (O_1588,N_49873,N_49990);
nor UO_1589 (O_1589,N_49332,N_49963);
or UO_1590 (O_1590,N_49221,N_49807);
xnor UO_1591 (O_1591,N_49655,N_49833);
nor UO_1592 (O_1592,N_49578,N_49434);
nand UO_1593 (O_1593,N_49579,N_49987);
or UO_1594 (O_1594,N_49946,N_49482);
and UO_1595 (O_1595,N_49040,N_49408);
nand UO_1596 (O_1596,N_49026,N_49378);
and UO_1597 (O_1597,N_49495,N_49028);
or UO_1598 (O_1598,N_49939,N_49546);
xor UO_1599 (O_1599,N_49532,N_49292);
nor UO_1600 (O_1600,N_49205,N_49174);
xnor UO_1601 (O_1601,N_49643,N_49677);
or UO_1602 (O_1602,N_49578,N_49436);
nand UO_1603 (O_1603,N_49640,N_49391);
nor UO_1604 (O_1604,N_49233,N_49691);
xnor UO_1605 (O_1605,N_49147,N_49338);
nand UO_1606 (O_1606,N_49024,N_49002);
xnor UO_1607 (O_1607,N_49264,N_49545);
xnor UO_1608 (O_1608,N_49911,N_49948);
nor UO_1609 (O_1609,N_49105,N_49772);
and UO_1610 (O_1610,N_49693,N_49502);
and UO_1611 (O_1611,N_49776,N_49693);
or UO_1612 (O_1612,N_49935,N_49082);
nor UO_1613 (O_1613,N_49566,N_49375);
or UO_1614 (O_1614,N_49740,N_49000);
and UO_1615 (O_1615,N_49491,N_49926);
nand UO_1616 (O_1616,N_49756,N_49009);
nor UO_1617 (O_1617,N_49574,N_49750);
nand UO_1618 (O_1618,N_49255,N_49729);
nor UO_1619 (O_1619,N_49355,N_49374);
nor UO_1620 (O_1620,N_49813,N_49033);
xnor UO_1621 (O_1621,N_49819,N_49586);
and UO_1622 (O_1622,N_49528,N_49275);
and UO_1623 (O_1623,N_49358,N_49443);
nand UO_1624 (O_1624,N_49328,N_49115);
nand UO_1625 (O_1625,N_49144,N_49710);
nand UO_1626 (O_1626,N_49174,N_49048);
nand UO_1627 (O_1627,N_49246,N_49200);
nor UO_1628 (O_1628,N_49597,N_49101);
and UO_1629 (O_1629,N_49811,N_49413);
nor UO_1630 (O_1630,N_49882,N_49255);
xor UO_1631 (O_1631,N_49901,N_49297);
nand UO_1632 (O_1632,N_49436,N_49085);
nor UO_1633 (O_1633,N_49480,N_49562);
or UO_1634 (O_1634,N_49947,N_49311);
nand UO_1635 (O_1635,N_49168,N_49682);
xnor UO_1636 (O_1636,N_49163,N_49141);
nor UO_1637 (O_1637,N_49502,N_49888);
xor UO_1638 (O_1638,N_49155,N_49232);
or UO_1639 (O_1639,N_49459,N_49966);
nor UO_1640 (O_1640,N_49378,N_49196);
or UO_1641 (O_1641,N_49735,N_49623);
nand UO_1642 (O_1642,N_49807,N_49647);
nor UO_1643 (O_1643,N_49511,N_49689);
nand UO_1644 (O_1644,N_49584,N_49855);
nor UO_1645 (O_1645,N_49838,N_49398);
and UO_1646 (O_1646,N_49085,N_49940);
and UO_1647 (O_1647,N_49332,N_49759);
nand UO_1648 (O_1648,N_49893,N_49183);
nand UO_1649 (O_1649,N_49149,N_49662);
nor UO_1650 (O_1650,N_49785,N_49933);
nand UO_1651 (O_1651,N_49555,N_49935);
nor UO_1652 (O_1652,N_49182,N_49932);
nand UO_1653 (O_1653,N_49256,N_49393);
nand UO_1654 (O_1654,N_49497,N_49376);
nand UO_1655 (O_1655,N_49867,N_49375);
nand UO_1656 (O_1656,N_49069,N_49572);
and UO_1657 (O_1657,N_49740,N_49442);
xnor UO_1658 (O_1658,N_49992,N_49934);
nor UO_1659 (O_1659,N_49790,N_49058);
and UO_1660 (O_1660,N_49863,N_49411);
nor UO_1661 (O_1661,N_49174,N_49539);
xor UO_1662 (O_1662,N_49074,N_49473);
or UO_1663 (O_1663,N_49445,N_49310);
nand UO_1664 (O_1664,N_49269,N_49915);
nand UO_1665 (O_1665,N_49700,N_49001);
xnor UO_1666 (O_1666,N_49614,N_49666);
nand UO_1667 (O_1667,N_49349,N_49611);
and UO_1668 (O_1668,N_49851,N_49200);
nor UO_1669 (O_1669,N_49828,N_49032);
or UO_1670 (O_1670,N_49469,N_49411);
and UO_1671 (O_1671,N_49943,N_49949);
and UO_1672 (O_1672,N_49006,N_49270);
nor UO_1673 (O_1673,N_49553,N_49347);
nand UO_1674 (O_1674,N_49137,N_49288);
nand UO_1675 (O_1675,N_49788,N_49383);
nand UO_1676 (O_1676,N_49320,N_49729);
nand UO_1677 (O_1677,N_49592,N_49124);
nor UO_1678 (O_1678,N_49271,N_49555);
nor UO_1679 (O_1679,N_49615,N_49260);
nand UO_1680 (O_1680,N_49416,N_49738);
nand UO_1681 (O_1681,N_49651,N_49185);
and UO_1682 (O_1682,N_49613,N_49591);
or UO_1683 (O_1683,N_49077,N_49713);
nand UO_1684 (O_1684,N_49322,N_49974);
and UO_1685 (O_1685,N_49610,N_49955);
and UO_1686 (O_1686,N_49625,N_49900);
and UO_1687 (O_1687,N_49902,N_49383);
and UO_1688 (O_1688,N_49181,N_49454);
nand UO_1689 (O_1689,N_49722,N_49502);
or UO_1690 (O_1690,N_49423,N_49840);
and UO_1691 (O_1691,N_49737,N_49609);
xor UO_1692 (O_1692,N_49911,N_49392);
or UO_1693 (O_1693,N_49730,N_49204);
or UO_1694 (O_1694,N_49636,N_49919);
or UO_1695 (O_1695,N_49565,N_49924);
xnor UO_1696 (O_1696,N_49195,N_49087);
and UO_1697 (O_1697,N_49871,N_49078);
and UO_1698 (O_1698,N_49398,N_49471);
xor UO_1699 (O_1699,N_49856,N_49518);
and UO_1700 (O_1700,N_49463,N_49358);
nor UO_1701 (O_1701,N_49354,N_49274);
nor UO_1702 (O_1702,N_49712,N_49239);
or UO_1703 (O_1703,N_49528,N_49115);
xor UO_1704 (O_1704,N_49282,N_49298);
or UO_1705 (O_1705,N_49907,N_49716);
nand UO_1706 (O_1706,N_49220,N_49257);
xor UO_1707 (O_1707,N_49693,N_49270);
and UO_1708 (O_1708,N_49212,N_49673);
nand UO_1709 (O_1709,N_49914,N_49091);
nor UO_1710 (O_1710,N_49216,N_49955);
or UO_1711 (O_1711,N_49645,N_49515);
nand UO_1712 (O_1712,N_49388,N_49479);
xnor UO_1713 (O_1713,N_49561,N_49953);
nand UO_1714 (O_1714,N_49484,N_49280);
xnor UO_1715 (O_1715,N_49350,N_49339);
nand UO_1716 (O_1716,N_49659,N_49310);
nand UO_1717 (O_1717,N_49913,N_49940);
xor UO_1718 (O_1718,N_49960,N_49871);
xor UO_1719 (O_1719,N_49754,N_49000);
nor UO_1720 (O_1720,N_49176,N_49875);
or UO_1721 (O_1721,N_49560,N_49998);
nor UO_1722 (O_1722,N_49634,N_49379);
or UO_1723 (O_1723,N_49059,N_49924);
and UO_1724 (O_1724,N_49491,N_49300);
or UO_1725 (O_1725,N_49873,N_49328);
and UO_1726 (O_1726,N_49932,N_49089);
or UO_1727 (O_1727,N_49786,N_49616);
nor UO_1728 (O_1728,N_49846,N_49316);
or UO_1729 (O_1729,N_49490,N_49939);
and UO_1730 (O_1730,N_49645,N_49273);
nor UO_1731 (O_1731,N_49100,N_49495);
xnor UO_1732 (O_1732,N_49118,N_49023);
xnor UO_1733 (O_1733,N_49458,N_49992);
or UO_1734 (O_1734,N_49579,N_49709);
xnor UO_1735 (O_1735,N_49109,N_49271);
xnor UO_1736 (O_1736,N_49229,N_49463);
nor UO_1737 (O_1737,N_49513,N_49353);
and UO_1738 (O_1738,N_49391,N_49420);
and UO_1739 (O_1739,N_49861,N_49855);
or UO_1740 (O_1740,N_49075,N_49055);
nand UO_1741 (O_1741,N_49493,N_49288);
nor UO_1742 (O_1742,N_49124,N_49983);
xnor UO_1743 (O_1743,N_49156,N_49497);
or UO_1744 (O_1744,N_49086,N_49565);
xor UO_1745 (O_1745,N_49904,N_49017);
nand UO_1746 (O_1746,N_49684,N_49245);
or UO_1747 (O_1747,N_49635,N_49331);
or UO_1748 (O_1748,N_49321,N_49115);
nand UO_1749 (O_1749,N_49809,N_49956);
and UO_1750 (O_1750,N_49621,N_49982);
or UO_1751 (O_1751,N_49962,N_49546);
or UO_1752 (O_1752,N_49401,N_49542);
nand UO_1753 (O_1753,N_49501,N_49642);
and UO_1754 (O_1754,N_49514,N_49401);
or UO_1755 (O_1755,N_49777,N_49590);
nor UO_1756 (O_1756,N_49863,N_49385);
nor UO_1757 (O_1757,N_49813,N_49267);
nand UO_1758 (O_1758,N_49021,N_49303);
nor UO_1759 (O_1759,N_49003,N_49001);
and UO_1760 (O_1760,N_49446,N_49801);
or UO_1761 (O_1761,N_49312,N_49800);
nor UO_1762 (O_1762,N_49908,N_49287);
or UO_1763 (O_1763,N_49952,N_49475);
nor UO_1764 (O_1764,N_49324,N_49218);
xnor UO_1765 (O_1765,N_49690,N_49932);
nand UO_1766 (O_1766,N_49942,N_49368);
nor UO_1767 (O_1767,N_49746,N_49440);
or UO_1768 (O_1768,N_49957,N_49705);
and UO_1769 (O_1769,N_49448,N_49067);
nor UO_1770 (O_1770,N_49999,N_49900);
nand UO_1771 (O_1771,N_49597,N_49542);
nand UO_1772 (O_1772,N_49196,N_49731);
nand UO_1773 (O_1773,N_49178,N_49584);
nor UO_1774 (O_1774,N_49308,N_49210);
nand UO_1775 (O_1775,N_49246,N_49044);
xor UO_1776 (O_1776,N_49314,N_49903);
and UO_1777 (O_1777,N_49807,N_49916);
nor UO_1778 (O_1778,N_49314,N_49391);
nor UO_1779 (O_1779,N_49575,N_49542);
nand UO_1780 (O_1780,N_49968,N_49130);
nand UO_1781 (O_1781,N_49841,N_49795);
nand UO_1782 (O_1782,N_49372,N_49264);
or UO_1783 (O_1783,N_49587,N_49267);
xor UO_1784 (O_1784,N_49242,N_49333);
and UO_1785 (O_1785,N_49521,N_49944);
xor UO_1786 (O_1786,N_49435,N_49572);
xnor UO_1787 (O_1787,N_49084,N_49686);
nand UO_1788 (O_1788,N_49564,N_49120);
nand UO_1789 (O_1789,N_49659,N_49567);
nand UO_1790 (O_1790,N_49514,N_49199);
and UO_1791 (O_1791,N_49676,N_49585);
xor UO_1792 (O_1792,N_49476,N_49061);
nor UO_1793 (O_1793,N_49863,N_49441);
nand UO_1794 (O_1794,N_49325,N_49349);
or UO_1795 (O_1795,N_49077,N_49775);
xnor UO_1796 (O_1796,N_49350,N_49814);
or UO_1797 (O_1797,N_49195,N_49298);
and UO_1798 (O_1798,N_49297,N_49859);
nor UO_1799 (O_1799,N_49773,N_49448);
or UO_1800 (O_1800,N_49210,N_49126);
nor UO_1801 (O_1801,N_49624,N_49045);
nor UO_1802 (O_1802,N_49403,N_49029);
nor UO_1803 (O_1803,N_49339,N_49730);
xor UO_1804 (O_1804,N_49168,N_49624);
or UO_1805 (O_1805,N_49441,N_49028);
nand UO_1806 (O_1806,N_49160,N_49316);
nor UO_1807 (O_1807,N_49291,N_49867);
or UO_1808 (O_1808,N_49284,N_49806);
nor UO_1809 (O_1809,N_49424,N_49036);
and UO_1810 (O_1810,N_49684,N_49049);
nor UO_1811 (O_1811,N_49193,N_49542);
or UO_1812 (O_1812,N_49203,N_49734);
or UO_1813 (O_1813,N_49166,N_49971);
xnor UO_1814 (O_1814,N_49030,N_49744);
nor UO_1815 (O_1815,N_49807,N_49177);
and UO_1816 (O_1816,N_49314,N_49398);
nand UO_1817 (O_1817,N_49561,N_49065);
nor UO_1818 (O_1818,N_49357,N_49977);
or UO_1819 (O_1819,N_49216,N_49866);
and UO_1820 (O_1820,N_49205,N_49070);
and UO_1821 (O_1821,N_49034,N_49889);
and UO_1822 (O_1822,N_49959,N_49556);
or UO_1823 (O_1823,N_49133,N_49729);
and UO_1824 (O_1824,N_49192,N_49064);
and UO_1825 (O_1825,N_49685,N_49308);
nand UO_1826 (O_1826,N_49460,N_49588);
nand UO_1827 (O_1827,N_49834,N_49462);
nor UO_1828 (O_1828,N_49686,N_49402);
nand UO_1829 (O_1829,N_49034,N_49301);
nand UO_1830 (O_1830,N_49775,N_49698);
or UO_1831 (O_1831,N_49864,N_49490);
and UO_1832 (O_1832,N_49213,N_49732);
nor UO_1833 (O_1833,N_49345,N_49682);
xor UO_1834 (O_1834,N_49987,N_49475);
nand UO_1835 (O_1835,N_49451,N_49018);
xnor UO_1836 (O_1836,N_49048,N_49778);
nor UO_1837 (O_1837,N_49797,N_49975);
or UO_1838 (O_1838,N_49862,N_49324);
nand UO_1839 (O_1839,N_49600,N_49927);
and UO_1840 (O_1840,N_49750,N_49326);
nor UO_1841 (O_1841,N_49752,N_49167);
nand UO_1842 (O_1842,N_49839,N_49046);
or UO_1843 (O_1843,N_49305,N_49288);
or UO_1844 (O_1844,N_49239,N_49806);
nor UO_1845 (O_1845,N_49661,N_49180);
and UO_1846 (O_1846,N_49891,N_49435);
nor UO_1847 (O_1847,N_49141,N_49533);
nor UO_1848 (O_1848,N_49850,N_49245);
nand UO_1849 (O_1849,N_49012,N_49799);
or UO_1850 (O_1850,N_49087,N_49610);
nand UO_1851 (O_1851,N_49650,N_49678);
nor UO_1852 (O_1852,N_49660,N_49583);
xor UO_1853 (O_1853,N_49240,N_49746);
nor UO_1854 (O_1854,N_49256,N_49224);
or UO_1855 (O_1855,N_49697,N_49296);
nor UO_1856 (O_1856,N_49578,N_49605);
nor UO_1857 (O_1857,N_49989,N_49465);
xor UO_1858 (O_1858,N_49417,N_49622);
nand UO_1859 (O_1859,N_49735,N_49937);
nor UO_1860 (O_1860,N_49837,N_49279);
nor UO_1861 (O_1861,N_49697,N_49239);
or UO_1862 (O_1862,N_49155,N_49512);
or UO_1863 (O_1863,N_49253,N_49283);
or UO_1864 (O_1864,N_49623,N_49307);
or UO_1865 (O_1865,N_49260,N_49701);
xor UO_1866 (O_1866,N_49242,N_49463);
or UO_1867 (O_1867,N_49679,N_49237);
xor UO_1868 (O_1868,N_49902,N_49742);
nand UO_1869 (O_1869,N_49169,N_49272);
xor UO_1870 (O_1870,N_49016,N_49356);
and UO_1871 (O_1871,N_49103,N_49053);
nand UO_1872 (O_1872,N_49159,N_49111);
nor UO_1873 (O_1873,N_49246,N_49075);
nand UO_1874 (O_1874,N_49961,N_49538);
and UO_1875 (O_1875,N_49312,N_49933);
and UO_1876 (O_1876,N_49339,N_49938);
nor UO_1877 (O_1877,N_49121,N_49395);
nand UO_1878 (O_1878,N_49833,N_49096);
nor UO_1879 (O_1879,N_49475,N_49388);
xor UO_1880 (O_1880,N_49286,N_49355);
nand UO_1881 (O_1881,N_49007,N_49016);
xor UO_1882 (O_1882,N_49913,N_49773);
nor UO_1883 (O_1883,N_49985,N_49174);
nor UO_1884 (O_1884,N_49207,N_49172);
nand UO_1885 (O_1885,N_49451,N_49619);
nor UO_1886 (O_1886,N_49483,N_49408);
nor UO_1887 (O_1887,N_49337,N_49762);
xor UO_1888 (O_1888,N_49293,N_49411);
nand UO_1889 (O_1889,N_49987,N_49935);
xor UO_1890 (O_1890,N_49025,N_49114);
nand UO_1891 (O_1891,N_49354,N_49195);
nand UO_1892 (O_1892,N_49266,N_49088);
nor UO_1893 (O_1893,N_49862,N_49706);
and UO_1894 (O_1894,N_49227,N_49459);
nand UO_1895 (O_1895,N_49789,N_49819);
and UO_1896 (O_1896,N_49465,N_49940);
nor UO_1897 (O_1897,N_49475,N_49854);
xnor UO_1898 (O_1898,N_49168,N_49515);
xnor UO_1899 (O_1899,N_49350,N_49674);
nand UO_1900 (O_1900,N_49632,N_49795);
xnor UO_1901 (O_1901,N_49501,N_49643);
nand UO_1902 (O_1902,N_49950,N_49776);
and UO_1903 (O_1903,N_49527,N_49902);
xor UO_1904 (O_1904,N_49644,N_49910);
nand UO_1905 (O_1905,N_49100,N_49877);
and UO_1906 (O_1906,N_49225,N_49798);
and UO_1907 (O_1907,N_49486,N_49907);
nor UO_1908 (O_1908,N_49460,N_49666);
nor UO_1909 (O_1909,N_49411,N_49942);
xnor UO_1910 (O_1910,N_49649,N_49746);
and UO_1911 (O_1911,N_49652,N_49857);
or UO_1912 (O_1912,N_49768,N_49720);
xnor UO_1913 (O_1913,N_49139,N_49532);
xnor UO_1914 (O_1914,N_49474,N_49866);
xor UO_1915 (O_1915,N_49657,N_49801);
nor UO_1916 (O_1916,N_49493,N_49634);
or UO_1917 (O_1917,N_49280,N_49726);
and UO_1918 (O_1918,N_49905,N_49318);
xor UO_1919 (O_1919,N_49661,N_49672);
and UO_1920 (O_1920,N_49098,N_49594);
or UO_1921 (O_1921,N_49717,N_49115);
nand UO_1922 (O_1922,N_49659,N_49048);
nand UO_1923 (O_1923,N_49817,N_49858);
nor UO_1924 (O_1924,N_49030,N_49956);
xnor UO_1925 (O_1925,N_49736,N_49885);
or UO_1926 (O_1926,N_49837,N_49125);
nand UO_1927 (O_1927,N_49117,N_49448);
nand UO_1928 (O_1928,N_49356,N_49922);
or UO_1929 (O_1929,N_49652,N_49728);
or UO_1930 (O_1930,N_49784,N_49094);
xnor UO_1931 (O_1931,N_49456,N_49060);
xnor UO_1932 (O_1932,N_49367,N_49885);
and UO_1933 (O_1933,N_49836,N_49289);
and UO_1934 (O_1934,N_49484,N_49720);
xor UO_1935 (O_1935,N_49543,N_49886);
xnor UO_1936 (O_1936,N_49265,N_49449);
or UO_1937 (O_1937,N_49276,N_49828);
nand UO_1938 (O_1938,N_49217,N_49162);
xor UO_1939 (O_1939,N_49496,N_49727);
and UO_1940 (O_1940,N_49341,N_49404);
and UO_1941 (O_1941,N_49621,N_49437);
or UO_1942 (O_1942,N_49823,N_49004);
or UO_1943 (O_1943,N_49801,N_49279);
nor UO_1944 (O_1944,N_49764,N_49032);
nor UO_1945 (O_1945,N_49432,N_49096);
or UO_1946 (O_1946,N_49184,N_49231);
nand UO_1947 (O_1947,N_49578,N_49666);
or UO_1948 (O_1948,N_49210,N_49242);
nand UO_1949 (O_1949,N_49691,N_49210);
nor UO_1950 (O_1950,N_49825,N_49584);
or UO_1951 (O_1951,N_49292,N_49422);
nor UO_1952 (O_1952,N_49366,N_49357);
nand UO_1953 (O_1953,N_49079,N_49119);
nand UO_1954 (O_1954,N_49635,N_49916);
nand UO_1955 (O_1955,N_49035,N_49381);
nor UO_1956 (O_1956,N_49878,N_49742);
xor UO_1957 (O_1957,N_49622,N_49791);
and UO_1958 (O_1958,N_49895,N_49097);
and UO_1959 (O_1959,N_49136,N_49073);
or UO_1960 (O_1960,N_49350,N_49734);
nor UO_1961 (O_1961,N_49148,N_49553);
nor UO_1962 (O_1962,N_49533,N_49219);
nand UO_1963 (O_1963,N_49170,N_49770);
nor UO_1964 (O_1964,N_49875,N_49028);
and UO_1965 (O_1965,N_49741,N_49073);
or UO_1966 (O_1966,N_49358,N_49246);
or UO_1967 (O_1967,N_49495,N_49614);
nand UO_1968 (O_1968,N_49878,N_49852);
nor UO_1969 (O_1969,N_49139,N_49650);
or UO_1970 (O_1970,N_49403,N_49363);
and UO_1971 (O_1971,N_49587,N_49208);
and UO_1972 (O_1972,N_49151,N_49694);
xnor UO_1973 (O_1973,N_49082,N_49943);
xnor UO_1974 (O_1974,N_49093,N_49489);
or UO_1975 (O_1975,N_49160,N_49610);
or UO_1976 (O_1976,N_49455,N_49674);
nand UO_1977 (O_1977,N_49910,N_49752);
nor UO_1978 (O_1978,N_49677,N_49408);
nor UO_1979 (O_1979,N_49503,N_49902);
xor UO_1980 (O_1980,N_49628,N_49504);
nand UO_1981 (O_1981,N_49122,N_49850);
nor UO_1982 (O_1982,N_49213,N_49549);
nor UO_1983 (O_1983,N_49425,N_49545);
nand UO_1984 (O_1984,N_49470,N_49368);
nand UO_1985 (O_1985,N_49806,N_49043);
nor UO_1986 (O_1986,N_49181,N_49063);
nor UO_1987 (O_1987,N_49737,N_49089);
nor UO_1988 (O_1988,N_49165,N_49591);
xnor UO_1989 (O_1989,N_49139,N_49214);
xor UO_1990 (O_1990,N_49221,N_49014);
or UO_1991 (O_1991,N_49226,N_49643);
nand UO_1992 (O_1992,N_49255,N_49716);
and UO_1993 (O_1993,N_49850,N_49030);
nor UO_1994 (O_1994,N_49087,N_49466);
xnor UO_1995 (O_1995,N_49735,N_49915);
and UO_1996 (O_1996,N_49903,N_49336);
nor UO_1997 (O_1997,N_49422,N_49262);
nand UO_1998 (O_1998,N_49606,N_49883);
xnor UO_1999 (O_1999,N_49044,N_49747);
or UO_2000 (O_2000,N_49946,N_49419);
nor UO_2001 (O_2001,N_49682,N_49998);
nand UO_2002 (O_2002,N_49124,N_49591);
nand UO_2003 (O_2003,N_49914,N_49320);
and UO_2004 (O_2004,N_49805,N_49966);
nor UO_2005 (O_2005,N_49493,N_49798);
and UO_2006 (O_2006,N_49357,N_49567);
nand UO_2007 (O_2007,N_49646,N_49656);
nor UO_2008 (O_2008,N_49961,N_49401);
xnor UO_2009 (O_2009,N_49936,N_49075);
or UO_2010 (O_2010,N_49968,N_49584);
xnor UO_2011 (O_2011,N_49273,N_49052);
nand UO_2012 (O_2012,N_49383,N_49067);
or UO_2013 (O_2013,N_49756,N_49011);
nand UO_2014 (O_2014,N_49322,N_49979);
xor UO_2015 (O_2015,N_49183,N_49233);
nor UO_2016 (O_2016,N_49495,N_49687);
or UO_2017 (O_2017,N_49804,N_49033);
nor UO_2018 (O_2018,N_49991,N_49822);
or UO_2019 (O_2019,N_49282,N_49715);
nor UO_2020 (O_2020,N_49617,N_49991);
nand UO_2021 (O_2021,N_49754,N_49386);
and UO_2022 (O_2022,N_49141,N_49026);
and UO_2023 (O_2023,N_49626,N_49906);
nand UO_2024 (O_2024,N_49466,N_49801);
nor UO_2025 (O_2025,N_49375,N_49459);
xor UO_2026 (O_2026,N_49336,N_49327);
and UO_2027 (O_2027,N_49867,N_49141);
and UO_2028 (O_2028,N_49143,N_49204);
xnor UO_2029 (O_2029,N_49736,N_49673);
and UO_2030 (O_2030,N_49899,N_49045);
nor UO_2031 (O_2031,N_49991,N_49329);
nor UO_2032 (O_2032,N_49886,N_49619);
nor UO_2033 (O_2033,N_49623,N_49982);
xnor UO_2034 (O_2034,N_49268,N_49338);
or UO_2035 (O_2035,N_49724,N_49187);
and UO_2036 (O_2036,N_49011,N_49526);
nor UO_2037 (O_2037,N_49480,N_49424);
nand UO_2038 (O_2038,N_49846,N_49328);
nor UO_2039 (O_2039,N_49600,N_49479);
or UO_2040 (O_2040,N_49890,N_49456);
and UO_2041 (O_2041,N_49591,N_49182);
or UO_2042 (O_2042,N_49475,N_49007);
nor UO_2043 (O_2043,N_49565,N_49666);
and UO_2044 (O_2044,N_49256,N_49149);
xnor UO_2045 (O_2045,N_49698,N_49080);
nand UO_2046 (O_2046,N_49180,N_49203);
nor UO_2047 (O_2047,N_49232,N_49391);
or UO_2048 (O_2048,N_49386,N_49539);
or UO_2049 (O_2049,N_49164,N_49898);
and UO_2050 (O_2050,N_49412,N_49783);
nor UO_2051 (O_2051,N_49474,N_49705);
nor UO_2052 (O_2052,N_49966,N_49310);
xor UO_2053 (O_2053,N_49928,N_49376);
nand UO_2054 (O_2054,N_49687,N_49352);
xnor UO_2055 (O_2055,N_49292,N_49055);
or UO_2056 (O_2056,N_49511,N_49501);
xor UO_2057 (O_2057,N_49345,N_49564);
and UO_2058 (O_2058,N_49783,N_49891);
or UO_2059 (O_2059,N_49137,N_49959);
nor UO_2060 (O_2060,N_49519,N_49155);
or UO_2061 (O_2061,N_49657,N_49048);
and UO_2062 (O_2062,N_49478,N_49550);
nand UO_2063 (O_2063,N_49826,N_49465);
nor UO_2064 (O_2064,N_49483,N_49025);
nor UO_2065 (O_2065,N_49453,N_49118);
xnor UO_2066 (O_2066,N_49624,N_49591);
nor UO_2067 (O_2067,N_49154,N_49314);
and UO_2068 (O_2068,N_49779,N_49282);
or UO_2069 (O_2069,N_49980,N_49009);
or UO_2070 (O_2070,N_49713,N_49764);
xor UO_2071 (O_2071,N_49881,N_49271);
or UO_2072 (O_2072,N_49038,N_49435);
or UO_2073 (O_2073,N_49961,N_49586);
nand UO_2074 (O_2074,N_49342,N_49205);
nand UO_2075 (O_2075,N_49481,N_49483);
or UO_2076 (O_2076,N_49539,N_49230);
nand UO_2077 (O_2077,N_49518,N_49750);
nand UO_2078 (O_2078,N_49386,N_49380);
nand UO_2079 (O_2079,N_49499,N_49001);
nor UO_2080 (O_2080,N_49166,N_49991);
nand UO_2081 (O_2081,N_49961,N_49589);
and UO_2082 (O_2082,N_49315,N_49227);
xor UO_2083 (O_2083,N_49087,N_49277);
or UO_2084 (O_2084,N_49078,N_49123);
xnor UO_2085 (O_2085,N_49366,N_49421);
nand UO_2086 (O_2086,N_49133,N_49387);
or UO_2087 (O_2087,N_49591,N_49928);
and UO_2088 (O_2088,N_49314,N_49265);
nor UO_2089 (O_2089,N_49072,N_49016);
xnor UO_2090 (O_2090,N_49094,N_49292);
nor UO_2091 (O_2091,N_49593,N_49030);
xor UO_2092 (O_2092,N_49167,N_49046);
or UO_2093 (O_2093,N_49169,N_49820);
nor UO_2094 (O_2094,N_49878,N_49400);
xnor UO_2095 (O_2095,N_49283,N_49185);
xnor UO_2096 (O_2096,N_49429,N_49189);
or UO_2097 (O_2097,N_49125,N_49992);
xor UO_2098 (O_2098,N_49400,N_49571);
nor UO_2099 (O_2099,N_49369,N_49949);
nand UO_2100 (O_2100,N_49491,N_49499);
or UO_2101 (O_2101,N_49440,N_49472);
nand UO_2102 (O_2102,N_49519,N_49356);
nor UO_2103 (O_2103,N_49084,N_49238);
nor UO_2104 (O_2104,N_49405,N_49643);
xor UO_2105 (O_2105,N_49619,N_49177);
nand UO_2106 (O_2106,N_49660,N_49780);
nor UO_2107 (O_2107,N_49150,N_49637);
nand UO_2108 (O_2108,N_49961,N_49510);
xnor UO_2109 (O_2109,N_49459,N_49441);
xor UO_2110 (O_2110,N_49838,N_49997);
nor UO_2111 (O_2111,N_49812,N_49486);
or UO_2112 (O_2112,N_49311,N_49341);
nand UO_2113 (O_2113,N_49030,N_49187);
and UO_2114 (O_2114,N_49677,N_49656);
and UO_2115 (O_2115,N_49647,N_49099);
xnor UO_2116 (O_2116,N_49601,N_49961);
xor UO_2117 (O_2117,N_49604,N_49107);
or UO_2118 (O_2118,N_49945,N_49309);
nor UO_2119 (O_2119,N_49330,N_49880);
nor UO_2120 (O_2120,N_49329,N_49613);
or UO_2121 (O_2121,N_49577,N_49031);
or UO_2122 (O_2122,N_49871,N_49083);
nand UO_2123 (O_2123,N_49288,N_49850);
nand UO_2124 (O_2124,N_49170,N_49897);
or UO_2125 (O_2125,N_49886,N_49169);
and UO_2126 (O_2126,N_49406,N_49972);
or UO_2127 (O_2127,N_49627,N_49890);
xnor UO_2128 (O_2128,N_49774,N_49431);
or UO_2129 (O_2129,N_49865,N_49592);
nor UO_2130 (O_2130,N_49298,N_49436);
nand UO_2131 (O_2131,N_49443,N_49101);
nor UO_2132 (O_2132,N_49576,N_49891);
or UO_2133 (O_2133,N_49772,N_49864);
nand UO_2134 (O_2134,N_49806,N_49850);
nand UO_2135 (O_2135,N_49047,N_49450);
nand UO_2136 (O_2136,N_49978,N_49554);
or UO_2137 (O_2137,N_49336,N_49937);
nand UO_2138 (O_2138,N_49067,N_49149);
nand UO_2139 (O_2139,N_49755,N_49918);
nor UO_2140 (O_2140,N_49306,N_49057);
xnor UO_2141 (O_2141,N_49788,N_49731);
and UO_2142 (O_2142,N_49919,N_49190);
nand UO_2143 (O_2143,N_49800,N_49747);
nor UO_2144 (O_2144,N_49105,N_49584);
nor UO_2145 (O_2145,N_49959,N_49186);
xnor UO_2146 (O_2146,N_49035,N_49996);
or UO_2147 (O_2147,N_49580,N_49997);
or UO_2148 (O_2148,N_49790,N_49551);
and UO_2149 (O_2149,N_49459,N_49286);
or UO_2150 (O_2150,N_49750,N_49050);
nor UO_2151 (O_2151,N_49703,N_49168);
nand UO_2152 (O_2152,N_49616,N_49596);
and UO_2153 (O_2153,N_49327,N_49053);
nand UO_2154 (O_2154,N_49564,N_49314);
and UO_2155 (O_2155,N_49818,N_49732);
xor UO_2156 (O_2156,N_49710,N_49212);
nor UO_2157 (O_2157,N_49449,N_49214);
and UO_2158 (O_2158,N_49003,N_49153);
or UO_2159 (O_2159,N_49453,N_49153);
nor UO_2160 (O_2160,N_49699,N_49217);
and UO_2161 (O_2161,N_49909,N_49778);
nor UO_2162 (O_2162,N_49469,N_49724);
or UO_2163 (O_2163,N_49594,N_49186);
or UO_2164 (O_2164,N_49698,N_49301);
and UO_2165 (O_2165,N_49678,N_49850);
nor UO_2166 (O_2166,N_49088,N_49021);
xnor UO_2167 (O_2167,N_49997,N_49276);
or UO_2168 (O_2168,N_49167,N_49818);
xnor UO_2169 (O_2169,N_49866,N_49670);
nor UO_2170 (O_2170,N_49325,N_49775);
xnor UO_2171 (O_2171,N_49010,N_49940);
nand UO_2172 (O_2172,N_49974,N_49102);
xnor UO_2173 (O_2173,N_49428,N_49911);
nand UO_2174 (O_2174,N_49412,N_49713);
nand UO_2175 (O_2175,N_49853,N_49874);
xor UO_2176 (O_2176,N_49773,N_49386);
xnor UO_2177 (O_2177,N_49520,N_49413);
nand UO_2178 (O_2178,N_49028,N_49100);
or UO_2179 (O_2179,N_49025,N_49974);
nor UO_2180 (O_2180,N_49932,N_49440);
nor UO_2181 (O_2181,N_49202,N_49901);
nor UO_2182 (O_2182,N_49727,N_49265);
xnor UO_2183 (O_2183,N_49397,N_49272);
and UO_2184 (O_2184,N_49175,N_49264);
nand UO_2185 (O_2185,N_49641,N_49130);
or UO_2186 (O_2186,N_49371,N_49049);
nor UO_2187 (O_2187,N_49405,N_49089);
nand UO_2188 (O_2188,N_49318,N_49313);
and UO_2189 (O_2189,N_49400,N_49240);
or UO_2190 (O_2190,N_49544,N_49356);
nor UO_2191 (O_2191,N_49016,N_49831);
nand UO_2192 (O_2192,N_49113,N_49871);
xor UO_2193 (O_2193,N_49350,N_49907);
or UO_2194 (O_2194,N_49983,N_49588);
or UO_2195 (O_2195,N_49144,N_49596);
or UO_2196 (O_2196,N_49061,N_49819);
nor UO_2197 (O_2197,N_49796,N_49142);
xor UO_2198 (O_2198,N_49094,N_49107);
xor UO_2199 (O_2199,N_49975,N_49996);
xor UO_2200 (O_2200,N_49867,N_49592);
nand UO_2201 (O_2201,N_49818,N_49359);
or UO_2202 (O_2202,N_49639,N_49797);
xnor UO_2203 (O_2203,N_49403,N_49303);
nand UO_2204 (O_2204,N_49691,N_49340);
or UO_2205 (O_2205,N_49583,N_49973);
and UO_2206 (O_2206,N_49423,N_49666);
and UO_2207 (O_2207,N_49406,N_49101);
or UO_2208 (O_2208,N_49270,N_49659);
or UO_2209 (O_2209,N_49608,N_49760);
nor UO_2210 (O_2210,N_49922,N_49579);
and UO_2211 (O_2211,N_49005,N_49393);
xnor UO_2212 (O_2212,N_49170,N_49246);
nand UO_2213 (O_2213,N_49938,N_49083);
and UO_2214 (O_2214,N_49268,N_49879);
and UO_2215 (O_2215,N_49213,N_49448);
or UO_2216 (O_2216,N_49258,N_49250);
nor UO_2217 (O_2217,N_49433,N_49207);
nand UO_2218 (O_2218,N_49116,N_49305);
or UO_2219 (O_2219,N_49233,N_49388);
nor UO_2220 (O_2220,N_49070,N_49642);
nor UO_2221 (O_2221,N_49649,N_49013);
nor UO_2222 (O_2222,N_49691,N_49930);
nand UO_2223 (O_2223,N_49549,N_49410);
and UO_2224 (O_2224,N_49154,N_49002);
xnor UO_2225 (O_2225,N_49782,N_49069);
nor UO_2226 (O_2226,N_49338,N_49630);
xnor UO_2227 (O_2227,N_49196,N_49907);
nand UO_2228 (O_2228,N_49865,N_49781);
xor UO_2229 (O_2229,N_49361,N_49927);
xnor UO_2230 (O_2230,N_49448,N_49573);
xor UO_2231 (O_2231,N_49152,N_49021);
nor UO_2232 (O_2232,N_49761,N_49862);
nand UO_2233 (O_2233,N_49486,N_49588);
xnor UO_2234 (O_2234,N_49434,N_49754);
nor UO_2235 (O_2235,N_49658,N_49920);
xor UO_2236 (O_2236,N_49917,N_49983);
nand UO_2237 (O_2237,N_49598,N_49659);
nor UO_2238 (O_2238,N_49055,N_49038);
and UO_2239 (O_2239,N_49231,N_49429);
nor UO_2240 (O_2240,N_49117,N_49602);
and UO_2241 (O_2241,N_49108,N_49512);
xnor UO_2242 (O_2242,N_49705,N_49521);
and UO_2243 (O_2243,N_49023,N_49871);
nand UO_2244 (O_2244,N_49564,N_49587);
and UO_2245 (O_2245,N_49563,N_49451);
nand UO_2246 (O_2246,N_49966,N_49372);
nor UO_2247 (O_2247,N_49330,N_49611);
xor UO_2248 (O_2248,N_49699,N_49278);
nand UO_2249 (O_2249,N_49007,N_49644);
nor UO_2250 (O_2250,N_49476,N_49166);
and UO_2251 (O_2251,N_49163,N_49940);
nand UO_2252 (O_2252,N_49476,N_49588);
or UO_2253 (O_2253,N_49465,N_49412);
and UO_2254 (O_2254,N_49598,N_49187);
xor UO_2255 (O_2255,N_49067,N_49225);
nand UO_2256 (O_2256,N_49818,N_49548);
nand UO_2257 (O_2257,N_49849,N_49116);
xnor UO_2258 (O_2258,N_49760,N_49294);
nand UO_2259 (O_2259,N_49670,N_49189);
nand UO_2260 (O_2260,N_49814,N_49137);
xnor UO_2261 (O_2261,N_49432,N_49659);
and UO_2262 (O_2262,N_49553,N_49959);
nor UO_2263 (O_2263,N_49895,N_49327);
xnor UO_2264 (O_2264,N_49410,N_49165);
xor UO_2265 (O_2265,N_49827,N_49619);
nor UO_2266 (O_2266,N_49225,N_49535);
xnor UO_2267 (O_2267,N_49891,N_49396);
or UO_2268 (O_2268,N_49386,N_49365);
and UO_2269 (O_2269,N_49212,N_49916);
nand UO_2270 (O_2270,N_49938,N_49585);
nand UO_2271 (O_2271,N_49517,N_49857);
nor UO_2272 (O_2272,N_49060,N_49403);
nor UO_2273 (O_2273,N_49948,N_49732);
and UO_2274 (O_2274,N_49824,N_49629);
and UO_2275 (O_2275,N_49103,N_49347);
nor UO_2276 (O_2276,N_49264,N_49240);
xnor UO_2277 (O_2277,N_49350,N_49426);
xor UO_2278 (O_2278,N_49754,N_49567);
and UO_2279 (O_2279,N_49796,N_49386);
nand UO_2280 (O_2280,N_49566,N_49897);
xor UO_2281 (O_2281,N_49054,N_49171);
nand UO_2282 (O_2282,N_49377,N_49740);
nor UO_2283 (O_2283,N_49094,N_49240);
or UO_2284 (O_2284,N_49996,N_49491);
and UO_2285 (O_2285,N_49300,N_49435);
and UO_2286 (O_2286,N_49654,N_49527);
nand UO_2287 (O_2287,N_49081,N_49014);
or UO_2288 (O_2288,N_49203,N_49105);
or UO_2289 (O_2289,N_49108,N_49164);
and UO_2290 (O_2290,N_49465,N_49043);
or UO_2291 (O_2291,N_49884,N_49373);
nor UO_2292 (O_2292,N_49443,N_49399);
nand UO_2293 (O_2293,N_49722,N_49979);
or UO_2294 (O_2294,N_49134,N_49078);
and UO_2295 (O_2295,N_49041,N_49792);
xor UO_2296 (O_2296,N_49322,N_49046);
xnor UO_2297 (O_2297,N_49335,N_49477);
and UO_2298 (O_2298,N_49573,N_49874);
and UO_2299 (O_2299,N_49535,N_49790);
nor UO_2300 (O_2300,N_49142,N_49295);
and UO_2301 (O_2301,N_49268,N_49667);
nand UO_2302 (O_2302,N_49467,N_49806);
nand UO_2303 (O_2303,N_49170,N_49282);
nand UO_2304 (O_2304,N_49714,N_49122);
nor UO_2305 (O_2305,N_49073,N_49841);
and UO_2306 (O_2306,N_49401,N_49684);
nor UO_2307 (O_2307,N_49654,N_49669);
nor UO_2308 (O_2308,N_49433,N_49954);
nand UO_2309 (O_2309,N_49484,N_49001);
nand UO_2310 (O_2310,N_49757,N_49891);
or UO_2311 (O_2311,N_49616,N_49630);
xnor UO_2312 (O_2312,N_49226,N_49686);
xor UO_2313 (O_2313,N_49630,N_49169);
or UO_2314 (O_2314,N_49415,N_49523);
and UO_2315 (O_2315,N_49251,N_49012);
or UO_2316 (O_2316,N_49371,N_49311);
xor UO_2317 (O_2317,N_49898,N_49045);
and UO_2318 (O_2318,N_49596,N_49282);
xnor UO_2319 (O_2319,N_49157,N_49225);
nand UO_2320 (O_2320,N_49715,N_49884);
nor UO_2321 (O_2321,N_49056,N_49168);
nor UO_2322 (O_2322,N_49198,N_49140);
nor UO_2323 (O_2323,N_49522,N_49101);
nor UO_2324 (O_2324,N_49536,N_49730);
or UO_2325 (O_2325,N_49305,N_49963);
nor UO_2326 (O_2326,N_49186,N_49334);
xor UO_2327 (O_2327,N_49589,N_49088);
nand UO_2328 (O_2328,N_49577,N_49979);
or UO_2329 (O_2329,N_49459,N_49697);
and UO_2330 (O_2330,N_49448,N_49010);
xnor UO_2331 (O_2331,N_49251,N_49657);
or UO_2332 (O_2332,N_49246,N_49397);
nand UO_2333 (O_2333,N_49822,N_49956);
nor UO_2334 (O_2334,N_49240,N_49689);
xnor UO_2335 (O_2335,N_49249,N_49941);
nand UO_2336 (O_2336,N_49211,N_49781);
xnor UO_2337 (O_2337,N_49977,N_49885);
nor UO_2338 (O_2338,N_49655,N_49191);
nand UO_2339 (O_2339,N_49531,N_49572);
nand UO_2340 (O_2340,N_49006,N_49741);
and UO_2341 (O_2341,N_49026,N_49995);
xor UO_2342 (O_2342,N_49062,N_49049);
or UO_2343 (O_2343,N_49319,N_49141);
nand UO_2344 (O_2344,N_49144,N_49272);
nor UO_2345 (O_2345,N_49609,N_49339);
xor UO_2346 (O_2346,N_49196,N_49195);
and UO_2347 (O_2347,N_49092,N_49435);
nor UO_2348 (O_2348,N_49669,N_49230);
xor UO_2349 (O_2349,N_49550,N_49133);
nand UO_2350 (O_2350,N_49108,N_49205);
or UO_2351 (O_2351,N_49278,N_49819);
nor UO_2352 (O_2352,N_49586,N_49116);
or UO_2353 (O_2353,N_49504,N_49182);
xor UO_2354 (O_2354,N_49408,N_49416);
xnor UO_2355 (O_2355,N_49983,N_49570);
nand UO_2356 (O_2356,N_49802,N_49133);
and UO_2357 (O_2357,N_49573,N_49539);
nand UO_2358 (O_2358,N_49752,N_49582);
nand UO_2359 (O_2359,N_49039,N_49685);
nor UO_2360 (O_2360,N_49282,N_49260);
or UO_2361 (O_2361,N_49015,N_49292);
nand UO_2362 (O_2362,N_49959,N_49034);
xor UO_2363 (O_2363,N_49320,N_49920);
and UO_2364 (O_2364,N_49887,N_49670);
or UO_2365 (O_2365,N_49344,N_49501);
nand UO_2366 (O_2366,N_49026,N_49198);
or UO_2367 (O_2367,N_49137,N_49849);
or UO_2368 (O_2368,N_49537,N_49091);
and UO_2369 (O_2369,N_49953,N_49782);
nand UO_2370 (O_2370,N_49159,N_49903);
or UO_2371 (O_2371,N_49842,N_49434);
or UO_2372 (O_2372,N_49525,N_49651);
and UO_2373 (O_2373,N_49852,N_49335);
nand UO_2374 (O_2374,N_49423,N_49846);
and UO_2375 (O_2375,N_49458,N_49263);
nor UO_2376 (O_2376,N_49841,N_49900);
or UO_2377 (O_2377,N_49228,N_49702);
or UO_2378 (O_2378,N_49902,N_49959);
or UO_2379 (O_2379,N_49277,N_49368);
and UO_2380 (O_2380,N_49394,N_49410);
nand UO_2381 (O_2381,N_49136,N_49937);
nor UO_2382 (O_2382,N_49887,N_49451);
or UO_2383 (O_2383,N_49686,N_49838);
nand UO_2384 (O_2384,N_49039,N_49435);
xnor UO_2385 (O_2385,N_49588,N_49569);
and UO_2386 (O_2386,N_49313,N_49202);
or UO_2387 (O_2387,N_49971,N_49363);
and UO_2388 (O_2388,N_49420,N_49834);
and UO_2389 (O_2389,N_49555,N_49559);
xor UO_2390 (O_2390,N_49748,N_49239);
nand UO_2391 (O_2391,N_49149,N_49515);
and UO_2392 (O_2392,N_49055,N_49245);
nor UO_2393 (O_2393,N_49183,N_49536);
xor UO_2394 (O_2394,N_49682,N_49922);
nor UO_2395 (O_2395,N_49490,N_49231);
nand UO_2396 (O_2396,N_49391,N_49478);
nor UO_2397 (O_2397,N_49752,N_49678);
or UO_2398 (O_2398,N_49762,N_49426);
and UO_2399 (O_2399,N_49756,N_49356);
and UO_2400 (O_2400,N_49418,N_49588);
or UO_2401 (O_2401,N_49769,N_49430);
xor UO_2402 (O_2402,N_49315,N_49195);
xnor UO_2403 (O_2403,N_49750,N_49134);
and UO_2404 (O_2404,N_49304,N_49992);
and UO_2405 (O_2405,N_49874,N_49801);
and UO_2406 (O_2406,N_49612,N_49447);
nand UO_2407 (O_2407,N_49989,N_49277);
and UO_2408 (O_2408,N_49198,N_49110);
nor UO_2409 (O_2409,N_49524,N_49522);
xnor UO_2410 (O_2410,N_49934,N_49269);
nor UO_2411 (O_2411,N_49803,N_49321);
xnor UO_2412 (O_2412,N_49569,N_49271);
xnor UO_2413 (O_2413,N_49404,N_49616);
or UO_2414 (O_2414,N_49879,N_49361);
nor UO_2415 (O_2415,N_49946,N_49909);
nor UO_2416 (O_2416,N_49420,N_49333);
and UO_2417 (O_2417,N_49105,N_49927);
and UO_2418 (O_2418,N_49298,N_49142);
xnor UO_2419 (O_2419,N_49942,N_49972);
and UO_2420 (O_2420,N_49993,N_49589);
nand UO_2421 (O_2421,N_49596,N_49450);
nor UO_2422 (O_2422,N_49374,N_49874);
or UO_2423 (O_2423,N_49235,N_49316);
or UO_2424 (O_2424,N_49900,N_49007);
nor UO_2425 (O_2425,N_49602,N_49983);
nand UO_2426 (O_2426,N_49581,N_49847);
xnor UO_2427 (O_2427,N_49544,N_49490);
nor UO_2428 (O_2428,N_49252,N_49926);
nor UO_2429 (O_2429,N_49184,N_49925);
and UO_2430 (O_2430,N_49715,N_49740);
nor UO_2431 (O_2431,N_49956,N_49155);
or UO_2432 (O_2432,N_49497,N_49611);
nor UO_2433 (O_2433,N_49716,N_49932);
nand UO_2434 (O_2434,N_49106,N_49592);
nand UO_2435 (O_2435,N_49462,N_49666);
or UO_2436 (O_2436,N_49049,N_49265);
or UO_2437 (O_2437,N_49267,N_49200);
nor UO_2438 (O_2438,N_49772,N_49112);
and UO_2439 (O_2439,N_49808,N_49100);
or UO_2440 (O_2440,N_49772,N_49220);
xor UO_2441 (O_2441,N_49492,N_49788);
nor UO_2442 (O_2442,N_49582,N_49066);
and UO_2443 (O_2443,N_49056,N_49726);
and UO_2444 (O_2444,N_49677,N_49905);
xor UO_2445 (O_2445,N_49679,N_49693);
nand UO_2446 (O_2446,N_49944,N_49229);
xor UO_2447 (O_2447,N_49560,N_49090);
and UO_2448 (O_2448,N_49600,N_49615);
or UO_2449 (O_2449,N_49192,N_49610);
nand UO_2450 (O_2450,N_49785,N_49452);
or UO_2451 (O_2451,N_49817,N_49280);
and UO_2452 (O_2452,N_49054,N_49880);
xor UO_2453 (O_2453,N_49827,N_49313);
nand UO_2454 (O_2454,N_49573,N_49699);
nor UO_2455 (O_2455,N_49533,N_49280);
xnor UO_2456 (O_2456,N_49863,N_49210);
nor UO_2457 (O_2457,N_49179,N_49900);
or UO_2458 (O_2458,N_49292,N_49542);
nand UO_2459 (O_2459,N_49990,N_49173);
and UO_2460 (O_2460,N_49100,N_49938);
and UO_2461 (O_2461,N_49300,N_49011);
nand UO_2462 (O_2462,N_49205,N_49237);
or UO_2463 (O_2463,N_49618,N_49105);
xor UO_2464 (O_2464,N_49078,N_49045);
nand UO_2465 (O_2465,N_49689,N_49149);
or UO_2466 (O_2466,N_49268,N_49304);
xnor UO_2467 (O_2467,N_49483,N_49745);
nand UO_2468 (O_2468,N_49988,N_49967);
nor UO_2469 (O_2469,N_49328,N_49705);
xor UO_2470 (O_2470,N_49546,N_49475);
and UO_2471 (O_2471,N_49842,N_49199);
nand UO_2472 (O_2472,N_49957,N_49819);
xnor UO_2473 (O_2473,N_49831,N_49806);
nand UO_2474 (O_2474,N_49589,N_49186);
xnor UO_2475 (O_2475,N_49981,N_49515);
or UO_2476 (O_2476,N_49283,N_49169);
or UO_2477 (O_2477,N_49553,N_49575);
nor UO_2478 (O_2478,N_49464,N_49388);
nand UO_2479 (O_2479,N_49527,N_49298);
xnor UO_2480 (O_2480,N_49300,N_49361);
nor UO_2481 (O_2481,N_49097,N_49013);
nor UO_2482 (O_2482,N_49428,N_49057);
nand UO_2483 (O_2483,N_49786,N_49451);
nor UO_2484 (O_2484,N_49042,N_49935);
or UO_2485 (O_2485,N_49715,N_49406);
and UO_2486 (O_2486,N_49838,N_49918);
nand UO_2487 (O_2487,N_49186,N_49537);
or UO_2488 (O_2488,N_49842,N_49594);
xnor UO_2489 (O_2489,N_49053,N_49665);
and UO_2490 (O_2490,N_49718,N_49349);
and UO_2491 (O_2491,N_49103,N_49557);
or UO_2492 (O_2492,N_49426,N_49957);
nor UO_2493 (O_2493,N_49212,N_49364);
nor UO_2494 (O_2494,N_49662,N_49943);
and UO_2495 (O_2495,N_49470,N_49779);
and UO_2496 (O_2496,N_49434,N_49998);
xor UO_2497 (O_2497,N_49629,N_49440);
nor UO_2498 (O_2498,N_49051,N_49622);
nor UO_2499 (O_2499,N_49829,N_49165);
and UO_2500 (O_2500,N_49888,N_49623);
and UO_2501 (O_2501,N_49066,N_49764);
and UO_2502 (O_2502,N_49247,N_49824);
nand UO_2503 (O_2503,N_49719,N_49118);
nor UO_2504 (O_2504,N_49978,N_49957);
and UO_2505 (O_2505,N_49876,N_49718);
and UO_2506 (O_2506,N_49143,N_49885);
nor UO_2507 (O_2507,N_49708,N_49731);
nand UO_2508 (O_2508,N_49873,N_49757);
nand UO_2509 (O_2509,N_49094,N_49560);
nor UO_2510 (O_2510,N_49890,N_49739);
or UO_2511 (O_2511,N_49809,N_49895);
nor UO_2512 (O_2512,N_49868,N_49200);
and UO_2513 (O_2513,N_49186,N_49885);
nand UO_2514 (O_2514,N_49956,N_49939);
xnor UO_2515 (O_2515,N_49857,N_49805);
and UO_2516 (O_2516,N_49712,N_49711);
xnor UO_2517 (O_2517,N_49875,N_49296);
nor UO_2518 (O_2518,N_49493,N_49047);
nand UO_2519 (O_2519,N_49645,N_49854);
or UO_2520 (O_2520,N_49206,N_49032);
nand UO_2521 (O_2521,N_49716,N_49562);
or UO_2522 (O_2522,N_49442,N_49678);
nor UO_2523 (O_2523,N_49423,N_49279);
nand UO_2524 (O_2524,N_49294,N_49245);
or UO_2525 (O_2525,N_49014,N_49701);
and UO_2526 (O_2526,N_49310,N_49035);
xor UO_2527 (O_2527,N_49405,N_49172);
nor UO_2528 (O_2528,N_49228,N_49218);
nor UO_2529 (O_2529,N_49537,N_49323);
nor UO_2530 (O_2530,N_49882,N_49998);
or UO_2531 (O_2531,N_49563,N_49436);
nand UO_2532 (O_2532,N_49301,N_49527);
nand UO_2533 (O_2533,N_49349,N_49677);
nor UO_2534 (O_2534,N_49254,N_49193);
or UO_2535 (O_2535,N_49104,N_49132);
nand UO_2536 (O_2536,N_49324,N_49938);
nor UO_2537 (O_2537,N_49484,N_49837);
or UO_2538 (O_2538,N_49691,N_49738);
nand UO_2539 (O_2539,N_49600,N_49709);
and UO_2540 (O_2540,N_49191,N_49650);
and UO_2541 (O_2541,N_49140,N_49732);
xor UO_2542 (O_2542,N_49157,N_49532);
and UO_2543 (O_2543,N_49388,N_49297);
nand UO_2544 (O_2544,N_49450,N_49541);
nor UO_2545 (O_2545,N_49898,N_49241);
xor UO_2546 (O_2546,N_49705,N_49488);
xor UO_2547 (O_2547,N_49065,N_49164);
or UO_2548 (O_2548,N_49462,N_49918);
nor UO_2549 (O_2549,N_49543,N_49961);
or UO_2550 (O_2550,N_49037,N_49032);
nand UO_2551 (O_2551,N_49205,N_49633);
xnor UO_2552 (O_2552,N_49544,N_49998);
xnor UO_2553 (O_2553,N_49687,N_49285);
and UO_2554 (O_2554,N_49620,N_49083);
and UO_2555 (O_2555,N_49318,N_49060);
or UO_2556 (O_2556,N_49109,N_49852);
nor UO_2557 (O_2557,N_49226,N_49006);
nand UO_2558 (O_2558,N_49614,N_49467);
nor UO_2559 (O_2559,N_49383,N_49724);
nand UO_2560 (O_2560,N_49180,N_49625);
nor UO_2561 (O_2561,N_49093,N_49042);
nand UO_2562 (O_2562,N_49294,N_49150);
xnor UO_2563 (O_2563,N_49796,N_49228);
and UO_2564 (O_2564,N_49136,N_49423);
xor UO_2565 (O_2565,N_49749,N_49590);
and UO_2566 (O_2566,N_49277,N_49711);
nor UO_2567 (O_2567,N_49638,N_49367);
nand UO_2568 (O_2568,N_49322,N_49536);
and UO_2569 (O_2569,N_49194,N_49169);
xor UO_2570 (O_2570,N_49260,N_49583);
and UO_2571 (O_2571,N_49545,N_49135);
or UO_2572 (O_2572,N_49765,N_49534);
or UO_2573 (O_2573,N_49273,N_49015);
or UO_2574 (O_2574,N_49238,N_49994);
and UO_2575 (O_2575,N_49889,N_49581);
and UO_2576 (O_2576,N_49074,N_49062);
nand UO_2577 (O_2577,N_49761,N_49085);
xnor UO_2578 (O_2578,N_49922,N_49088);
nor UO_2579 (O_2579,N_49578,N_49088);
nand UO_2580 (O_2580,N_49303,N_49156);
or UO_2581 (O_2581,N_49187,N_49179);
xor UO_2582 (O_2582,N_49012,N_49899);
xnor UO_2583 (O_2583,N_49334,N_49230);
nand UO_2584 (O_2584,N_49288,N_49896);
or UO_2585 (O_2585,N_49443,N_49197);
nor UO_2586 (O_2586,N_49527,N_49581);
xor UO_2587 (O_2587,N_49365,N_49702);
nor UO_2588 (O_2588,N_49340,N_49256);
and UO_2589 (O_2589,N_49381,N_49281);
or UO_2590 (O_2590,N_49928,N_49733);
and UO_2591 (O_2591,N_49992,N_49741);
or UO_2592 (O_2592,N_49221,N_49279);
nand UO_2593 (O_2593,N_49097,N_49083);
and UO_2594 (O_2594,N_49256,N_49147);
xnor UO_2595 (O_2595,N_49953,N_49817);
or UO_2596 (O_2596,N_49566,N_49787);
nor UO_2597 (O_2597,N_49606,N_49919);
xor UO_2598 (O_2598,N_49610,N_49983);
xor UO_2599 (O_2599,N_49255,N_49908);
and UO_2600 (O_2600,N_49788,N_49137);
nor UO_2601 (O_2601,N_49811,N_49815);
and UO_2602 (O_2602,N_49572,N_49077);
nor UO_2603 (O_2603,N_49922,N_49350);
or UO_2604 (O_2604,N_49866,N_49555);
nand UO_2605 (O_2605,N_49515,N_49754);
xor UO_2606 (O_2606,N_49267,N_49354);
and UO_2607 (O_2607,N_49232,N_49210);
or UO_2608 (O_2608,N_49500,N_49065);
xnor UO_2609 (O_2609,N_49485,N_49702);
nor UO_2610 (O_2610,N_49687,N_49460);
or UO_2611 (O_2611,N_49850,N_49048);
and UO_2612 (O_2612,N_49730,N_49870);
nand UO_2613 (O_2613,N_49781,N_49961);
or UO_2614 (O_2614,N_49046,N_49688);
and UO_2615 (O_2615,N_49403,N_49964);
or UO_2616 (O_2616,N_49139,N_49600);
nor UO_2617 (O_2617,N_49795,N_49867);
and UO_2618 (O_2618,N_49836,N_49863);
and UO_2619 (O_2619,N_49100,N_49888);
and UO_2620 (O_2620,N_49731,N_49491);
or UO_2621 (O_2621,N_49490,N_49495);
nand UO_2622 (O_2622,N_49534,N_49058);
nor UO_2623 (O_2623,N_49795,N_49381);
or UO_2624 (O_2624,N_49471,N_49252);
and UO_2625 (O_2625,N_49294,N_49773);
nand UO_2626 (O_2626,N_49170,N_49114);
nand UO_2627 (O_2627,N_49862,N_49756);
and UO_2628 (O_2628,N_49398,N_49301);
xor UO_2629 (O_2629,N_49032,N_49344);
nor UO_2630 (O_2630,N_49143,N_49790);
nor UO_2631 (O_2631,N_49228,N_49034);
nor UO_2632 (O_2632,N_49749,N_49704);
nand UO_2633 (O_2633,N_49879,N_49274);
xor UO_2634 (O_2634,N_49434,N_49313);
or UO_2635 (O_2635,N_49464,N_49963);
nand UO_2636 (O_2636,N_49081,N_49416);
and UO_2637 (O_2637,N_49662,N_49377);
nor UO_2638 (O_2638,N_49408,N_49943);
or UO_2639 (O_2639,N_49105,N_49262);
nand UO_2640 (O_2640,N_49270,N_49384);
nor UO_2641 (O_2641,N_49116,N_49814);
and UO_2642 (O_2642,N_49417,N_49682);
and UO_2643 (O_2643,N_49717,N_49027);
or UO_2644 (O_2644,N_49549,N_49373);
and UO_2645 (O_2645,N_49154,N_49012);
and UO_2646 (O_2646,N_49301,N_49712);
nand UO_2647 (O_2647,N_49972,N_49519);
and UO_2648 (O_2648,N_49259,N_49016);
nor UO_2649 (O_2649,N_49668,N_49136);
nor UO_2650 (O_2650,N_49708,N_49019);
xnor UO_2651 (O_2651,N_49140,N_49390);
xnor UO_2652 (O_2652,N_49604,N_49571);
and UO_2653 (O_2653,N_49498,N_49462);
xnor UO_2654 (O_2654,N_49166,N_49656);
xnor UO_2655 (O_2655,N_49732,N_49861);
nor UO_2656 (O_2656,N_49224,N_49330);
nand UO_2657 (O_2657,N_49870,N_49492);
nor UO_2658 (O_2658,N_49460,N_49941);
nor UO_2659 (O_2659,N_49597,N_49943);
nor UO_2660 (O_2660,N_49451,N_49490);
nor UO_2661 (O_2661,N_49759,N_49028);
xnor UO_2662 (O_2662,N_49402,N_49873);
or UO_2663 (O_2663,N_49446,N_49281);
nor UO_2664 (O_2664,N_49064,N_49850);
and UO_2665 (O_2665,N_49915,N_49396);
xor UO_2666 (O_2666,N_49270,N_49990);
or UO_2667 (O_2667,N_49575,N_49230);
nand UO_2668 (O_2668,N_49612,N_49389);
nand UO_2669 (O_2669,N_49800,N_49588);
xor UO_2670 (O_2670,N_49941,N_49345);
or UO_2671 (O_2671,N_49776,N_49602);
nor UO_2672 (O_2672,N_49045,N_49066);
xnor UO_2673 (O_2673,N_49050,N_49592);
and UO_2674 (O_2674,N_49465,N_49200);
and UO_2675 (O_2675,N_49965,N_49692);
nand UO_2676 (O_2676,N_49545,N_49197);
and UO_2677 (O_2677,N_49197,N_49810);
nand UO_2678 (O_2678,N_49002,N_49425);
or UO_2679 (O_2679,N_49761,N_49304);
xnor UO_2680 (O_2680,N_49739,N_49108);
or UO_2681 (O_2681,N_49238,N_49198);
nor UO_2682 (O_2682,N_49065,N_49236);
nand UO_2683 (O_2683,N_49106,N_49890);
or UO_2684 (O_2684,N_49601,N_49983);
nand UO_2685 (O_2685,N_49796,N_49729);
nor UO_2686 (O_2686,N_49535,N_49659);
or UO_2687 (O_2687,N_49793,N_49708);
and UO_2688 (O_2688,N_49348,N_49217);
and UO_2689 (O_2689,N_49018,N_49860);
or UO_2690 (O_2690,N_49333,N_49770);
or UO_2691 (O_2691,N_49618,N_49423);
nor UO_2692 (O_2692,N_49549,N_49846);
xnor UO_2693 (O_2693,N_49826,N_49966);
or UO_2694 (O_2694,N_49542,N_49678);
nand UO_2695 (O_2695,N_49591,N_49111);
xor UO_2696 (O_2696,N_49591,N_49090);
nor UO_2697 (O_2697,N_49122,N_49831);
nor UO_2698 (O_2698,N_49047,N_49842);
xor UO_2699 (O_2699,N_49322,N_49953);
nor UO_2700 (O_2700,N_49845,N_49140);
nand UO_2701 (O_2701,N_49194,N_49624);
and UO_2702 (O_2702,N_49264,N_49910);
and UO_2703 (O_2703,N_49465,N_49455);
nand UO_2704 (O_2704,N_49123,N_49995);
nand UO_2705 (O_2705,N_49288,N_49614);
or UO_2706 (O_2706,N_49501,N_49666);
nand UO_2707 (O_2707,N_49054,N_49677);
or UO_2708 (O_2708,N_49818,N_49503);
xor UO_2709 (O_2709,N_49016,N_49773);
and UO_2710 (O_2710,N_49686,N_49901);
or UO_2711 (O_2711,N_49790,N_49519);
xor UO_2712 (O_2712,N_49371,N_49866);
nand UO_2713 (O_2713,N_49255,N_49055);
xor UO_2714 (O_2714,N_49882,N_49008);
nor UO_2715 (O_2715,N_49619,N_49499);
nand UO_2716 (O_2716,N_49604,N_49597);
nor UO_2717 (O_2717,N_49403,N_49461);
xor UO_2718 (O_2718,N_49914,N_49154);
or UO_2719 (O_2719,N_49525,N_49673);
nand UO_2720 (O_2720,N_49597,N_49488);
xnor UO_2721 (O_2721,N_49259,N_49998);
or UO_2722 (O_2722,N_49764,N_49815);
or UO_2723 (O_2723,N_49547,N_49511);
nand UO_2724 (O_2724,N_49170,N_49808);
nand UO_2725 (O_2725,N_49599,N_49583);
or UO_2726 (O_2726,N_49695,N_49349);
or UO_2727 (O_2727,N_49911,N_49984);
nor UO_2728 (O_2728,N_49186,N_49743);
xnor UO_2729 (O_2729,N_49098,N_49923);
and UO_2730 (O_2730,N_49092,N_49939);
xor UO_2731 (O_2731,N_49359,N_49816);
or UO_2732 (O_2732,N_49338,N_49194);
xnor UO_2733 (O_2733,N_49488,N_49073);
nand UO_2734 (O_2734,N_49250,N_49605);
nand UO_2735 (O_2735,N_49823,N_49604);
and UO_2736 (O_2736,N_49740,N_49559);
and UO_2737 (O_2737,N_49669,N_49597);
xor UO_2738 (O_2738,N_49296,N_49433);
nor UO_2739 (O_2739,N_49869,N_49533);
nand UO_2740 (O_2740,N_49257,N_49602);
or UO_2741 (O_2741,N_49785,N_49624);
xnor UO_2742 (O_2742,N_49638,N_49327);
and UO_2743 (O_2743,N_49526,N_49044);
xnor UO_2744 (O_2744,N_49467,N_49742);
nand UO_2745 (O_2745,N_49920,N_49187);
or UO_2746 (O_2746,N_49179,N_49928);
nor UO_2747 (O_2747,N_49500,N_49590);
xnor UO_2748 (O_2748,N_49571,N_49464);
nor UO_2749 (O_2749,N_49993,N_49178);
and UO_2750 (O_2750,N_49613,N_49603);
and UO_2751 (O_2751,N_49513,N_49396);
xor UO_2752 (O_2752,N_49699,N_49478);
xor UO_2753 (O_2753,N_49863,N_49267);
nand UO_2754 (O_2754,N_49219,N_49778);
or UO_2755 (O_2755,N_49508,N_49775);
and UO_2756 (O_2756,N_49461,N_49658);
and UO_2757 (O_2757,N_49036,N_49095);
xor UO_2758 (O_2758,N_49559,N_49605);
nand UO_2759 (O_2759,N_49717,N_49784);
nor UO_2760 (O_2760,N_49266,N_49216);
and UO_2761 (O_2761,N_49425,N_49409);
nand UO_2762 (O_2762,N_49262,N_49865);
or UO_2763 (O_2763,N_49616,N_49277);
xor UO_2764 (O_2764,N_49735,N_49065);
nor UO_2765 (O_2765,N_49451,N_49312);
xnor UO_2766 (O_2766,N_49956,N_49940);
nand UO_2767 (O_2767,N_49462,N_49303);
nor UO_2768 (O_2768,N_49694,N_49097);
and UO_2769 (O_2769,N_49616,N_49204);
or UO_2770 (O_2770,N_49581,N_49444);
nor UO_2771 (O_2771,N_49588,N_49799);
nand UO_2772 (O_2772,N_49778,N_49009);
or UO_2773 (O_2773,N_49193,N_49716);
nor UO_2774 (O_2774,N_49567,N_49566);
nor UO_2775 (O_2775,N_49471,N_49443);
nand UO_2776 (O_2776,N_49109,N_49436);
xor UO_2777 (O_2777,N_49475,N_49789);
or UO_2778 (O_2778,N_49024,N_49303);
nand UO_2779 (O_2779,N_49746,N_49968);
and UO_2780 (O_2780,N_49569,N_49070);
xnor UO_2781 (O_2781,N_49461,N_49581);
xnor UO_2782 (O_2782,N_49823,N_49493);
xor UO_2783 (O_2783,N_49868,N_49338);
nor UO_2784 (O_2784,N_49319,N_49596);
nand UO_2785 (O_2785,N_49280,N_49958);
nor UO_2786 (O_2786,N_49775,N_49198);
and UO_2787 (O_2787,N_49617,N_49942);
nand UO_2788 (O_2788,N_49567,N_49176);
nand UO_2789 (O_2789,N_49351,N_49839);
nand UO_2790 (O_2790,N_49847,N_49704);
or UO_2791 (O_2791,N_49291,N_49509);
nand UO_2792 (O_2792,N_49614,N_49922);
xor UO_2793 (O_2793,N_49214,N_49945);
or UO_2794 (O_2794,N_49194,N_49905);
or UO_2795 (O_2795,N_49247,N_49597);
and UO_2796 (O_2796,N_49205,N_49757);
or UO_2797 (O_2797,N_49386,N_49510);
or UO_2798 (O_2798,N_49530,N_49818);
nor UO_2799 (O_2799,N_49528,N_49974);
xor UO_2800 (O_2800,N_49641,N_49646);
xnor UO_2801 (O_2801,N_49167,N_49015);
and UO_2802 (O_2802,N_49255,N_49582);
nand UO_2803 (O_2803,N_49468,N_49495);
nand UO_2804 (O_2804,N_49994,N_49930);
or UO_2805 (O_2805,N_49704,N_49629);
and UO_2806 (O_2806,N_49830,N_49154);
nor UO_2807 (O_2807,N_49718,N_49884);
nand UO_2808 (O_2808,N_49709,N_49259);
or UO_2809 (O_2809,N_49798,N_49241);
or UO_2810 (O_2810,N_49989,N_49294);
nor UO_2811 (O_2811,N_49615,N_49941);
xnor UO_2812 (O_2812,N_49895,N_49428);
xor UO_2813 (O_2813,N_49384,N_49074);
nand UO_2814 (O_2814,N_49250,N_49394);
and UO_2815 (O_2815,N_49799,N_49071);
and UO_2816 (O_2816,N_49216,N_49816);
or UO_2817 (O_2817,N_49612,N_49508);
nand UO_2818 (O_2818,N_49476,N_49041);
and UO_2819 (O_2819,N_49017,N_49453);
and UO_2820 (O_2820,N_49461,N_49640);
xor UO_2821 (O_2821,N_49515,N_49143);
nand UO_2822 (O_2822,N_49411,N_49522);
nor UO_2823 (O_2823,N_49072,N_49380);
nand UO_2824 (O_2824,N_49538,N_49421);
xnor UO_2825 (O_2825,N_49864,N_49765);
or UO_2826 (O_2826,N_49323,N_49349);
nor UO_2827 (O_2827,N_49045,N_49163);
nor UO_2828 (O_2828,N_49121,N_49862);
and UO_2829 (O_2829,N_49169,N_49250);
nand UO_2830 (O_2830,N_49954,N_49977);
nand UO_2831 (O_2831,N_49943,N_49807);
and UO_2832 (O_2832,N_49707,N_49487);
xnor UO_2833 (O_2833,N_49117,N_49897);
and UO_2834 (O_2834,N_49667,N_49089);
or UO_2835 (O_2835,N_49231,N_49543);
nor UO_2836 (O_2836,N_49967,N_49599);
nor UO_2837 (O_2837,N_49845,N_49750);
and UO_2838 (O_2838,N_49820,N_49326);
nand UO_2839 (O_2839,N_49689,N_49102);
and UO_2840 (O_2840,N_49462,N_49967);
and UO_2841 (O_2841,N_49160,N_49738);
and UO_2842 (O_2842,N_49149,N_49168);
xor UO_2843 (O_2843,N_49664,N_49316);
nor UO_2844 (O_2844,N_49723,N_49773);
xnor UO_2845 (O_2845,N_49998,N_49418);
xnor UO_2846 (O_2846,N_49315,N_49761);
and UO_2847 (O_2847,N_49073,N_49863);
and UO_2848 (O_2848,N_49423,N_49647);
nand UO_2849 (O_2849,N_49138,N_49803);
xnor UO_2850 (O_2850,N_49706,N_49703);
or UO_2851 (O_2851,N_49311,N_49361);
or UO_2852 (O_2852,N_49620,N_49817);
xor UO_2853 (O_2853,N_49617,N_49152);
nor UO_2854 (O_2854,N_49378,N_49992);
xnor UO_2855 (O_2855,N_49548,N_49317);
nand UO_2856 (O_2856,N_49213,N_49311);
xor UO_2857 (O_2857,N_49149,N_49223);
xor UO_2858 (O_2858,N_49167,N_49887);
xor UO_2859 (O_2859,N_49963,N_49036);
nor UO_2860 (O_2860,N_49513,N_49377);
and UO_2861 (O_2861,N_49150,N_49588);
xnor UO_2862 (O_2862,N_49220,N_49899);
nor UO_2863 (O_2863,N_49051,N_49245);
xnor UO_2864 (O_2864,N_49056,N_49594);
or UO_2865 (O_2865,N_49045,N_49555);
nand UO_2866 (O_2866,N_49609,N_49640);
nand UO_2867 (O_2867,N_49953,N_49673);
nor UO_2868 (O_2868,N_49197,N_49107);
and UO_2869 (O_2869,N_49629,N_49226);
and UO_2870 (O_2870,N_49516,N_49701);
or UO_2871 (O_2871,N_49290,N_49634);
xor UO_2872 (O_2872,N_49811,N_49585);
or UO_2873 (O_2873,N_49927,N_49128);
nand UO_2874 (O_2874,N_49270,N_49887);
xnor UO_2875 (O_2875,N_49052,N_49060);
and UO_2876 (O_2876,N_49016,N_49547);
and UO_2877 (O_2877,N_49913,N_49017);
and UO_2878 (O_2878,N_49325,N_49154);
nor UO_2879 (O_2879,N_49803,N_49292);
and UO_2880 (O_2880,N_49304,N_49334);
nand UO_2881 (O_2881,N_49336,N_49637);
nor UO_2882 (O_2882,N_49801,N_49504);
xnor UO_2883 (O_2883,N_49470,N_49604);
or UO_2884 (O_2884,N_49353,N_49718);
xnor UO_2885 (O_2885,N_49933,N_49128);
or UO_2886 (O_2886,N_49974,N_49787);
nand UO_2887 (O_2887,N_49379,N_49401);
nor UO_2888 (O_2888,N_49913,N_49260);
and UO_2889 (O_2889,N_49186,N_49941);
nor UO_2890 (O_2890,N_49745,N_49594);
nor UO_2891 (O_2891,N_49789,N_49275);
nand UO_2892 (O_2892,N_49980,N_49997);
or UO_2893 (O_2893,N_49611,N_49857);
or UO_2894 (O_2894,N_49190,N_49430);
xnor UO_2895 (O_2895,N_49367,N_49238);
and UO_2896 (O_2896,N_49809,N_49254);
xor UO_2897 (O_2897,N_49233,N_49780);
or UO_2898 (O_2898,N_49006,N_49645);
or UO_2899 (O_2899,N_49369,N_49662);
or UO_2900 (O_2900,N_49722,N_49988);
xor UO_2901 (O_2901,N_49647,N_49480);
and UO_2902 (O_2902,N_49120,N_49355);
nor UO_2903 (O_2903,N_49666,N_49592);
nor UO_2904 (O_2904,N_49816,N_49889);
xnor UO_2905 (O_2905,N_49294,N_49679);
nand UO_2906 (O_2906,N_49591,N_49706);
and UO_2907 (O_2907,N_49267,N_49818);
xnor UO_2908 (O_2908,N_49769,N_49874);
or UO_2909 (O_2909,N_49708,N_49357);
xnor UO_2910 (O_2910,N_49900,N_49898);
nand UO_2911 (O_2911,N_49209,N_49081);
nand UO_2912 (O_2912,N_49423,N_49216);
and UO_2913 (O_2913,N_49807,N_49247);
and UO_2914 (O_2914,N_49016,N_49115);
or UO_2915 (O_2915,N_49027,N_49868);
or UO_2916 (O_2916,N_49147,N_49214);
or UO_2917 (O_2917,N_49917,N_49706);
nand UO_2918 (O_2918,N_49767,N_49925);
nand UO_2919 (O_2919,N_49488,N_49689);
xnor UO_2920 (O_2920,N_49324,N_49073);
nand UO_2921 (O_2921,N_49389,N_49529);
nand UO_2922 (O_2922,N_49191,N_49677);
xnor UO_2923 (O_2923,N_49780,N_49190);
and UO_2924 (O_2924,N_49409,N_49159);
nand UO_2925 (O_2925,N_49772,N_49147);
and UO_2926 (O_2926,N_49724,N_49405);
or UO_2927 (O_2927,N_49216,N_49915);
nand UO_2928 (O_2928,N_49266,N_49597);
or UO_2929 (O_2929,N_49964,N_49416);
xor UO_2930 (O_2930,N_49340,N_49490);
or UO_2931 (O_2931,N_49867,N_49256);
or UO_2932 (O_2932,N_49861,N_49853);
nor UO_2933 (O_2933,N_49712,N_49423);
nor UO_2934 (O_2934,N_49325,N_49163);
xor UO_2935 (O_2935,N_49019,N_49236);
xor UO_2936 (O_2936,N_49439,N_49905);
nand UO_2937 (O_2937,N_49841,N_49844);
or UO_2938 (O_2938,N_49022,N_49597);
and UO_2939 (O_2939,N_49866,N_49679);
or UO_2940 (O_2940,N_49728,N_49621);
and UO_2941 (O_2941,N_49536,N_49792);
nor UO_2942 (O_2942,N_49557,N_49131);
nand UO_2943 (O_2943,N_49524,N_49640);
xnor UO_2944 (O_2944,N_49910,N_49680);
xnor UO_2945 (O_2945,N_49478,N_49740);
or UO_2946 (O_2946,N_49477,N_49342);
nand UO_2947 (O_2947,N_49583,N_49989);
and UO_2948 (O_2948,N_49171,N_49522);
and UO_2949 (O_2949,N_49377,N_49607);
nand UO_2950 (O_2950,N_49593,N_49280);
or UO_2951 (O_2951,N_49339,N_49261);
nor UO_2952 (O_2952,N_49152,N_49933);
xor UO_2953 (O_2953,N_49398,N_49893);
nor UO_2954 (O_2954,N_49348,N_49112);
or UO_2955 (O_2955,N_49738,N_49094);
and UO_2956 (O_2956,N_49369,N_49852);
or UO_2957 (O_2957,N_49644,N_49174);
xnor UO_2958 (O_2958,N_49911,N_49167);
and UO_2959 (O_2959,N_49600,N_49623);
or UO_2960 (O_2960,N_49835,N_49340);
nor UO_2961 (O_2961,N_49220,N_49673);
and UO_2962 (O_2962,N_49342,N_49446);
nor UO_2963 (O_2963,N_49090,N_49450);
and UO_2964 (O_2964,N_49148,N_49661);
xnor UO_2965 (O_2965,N_49385,N_49967);
nand UO_2966 (O_2966,N_49912,N_49032);
or UO_2967 (O_2967,N_49079,N_49169);
nor UO_2968 (O_2968,N_49515,N_49148);
or UO_2969 (O_2969,N_49522,N_49220);
nor UO_2970 (O_2970,N_49831,N_49915);
and UO_2971 (O_2971,N_49913,N_49969);
nand UO_2972 (O_2972,N_49258,N_49763);
xnor UO_2973 (O_2973,N_49429,N_49518);
xnor UO_2974 (O_2974,N_49368,N_49651);
or UO_2975 (O_2975,N_49016,N_49207);
or UO_2976 (O_2976,N_49843,N_49502);
nor UO_2977 (O_2977,N_49848,N_49755);
nor UO_2978 (O_2978,N_49421,N_49748);
nor UO_2979 (O_2979,N_49466,N_49165);
xnor UO_2980 (O_2980,N_49870,N_49410);
xnor UO_2981 (O_2981,N_49179,N_49487);
xor UO_2982 (O_2982,N_49502,N_49531);
or UO_2983 (O_2983,N_49185,N_49807);
and UO_2984 (O_2984,N_49418,N_49173);
nor UO_2985 (O_2985,N_49258,N_49917);
or UO_2986 (O_2986,N_49603,N_49852);
nor UO_2987 (O_2987,N_49138,N_49357);
nor UO_2988 (O_2988,N_49768,N_49239);
nand UO_2989 (O_2989,N_49766,N_49708);
or UO_2990 (O_2990,N_49797,N_49989);
nand UO_2991 (O_2991,N_49976,N_49653);
xor UO_2992 (O_2992,N_49616,N_49614);
nor UO_2993 (O_2993,N_49188,N_49256);
nor UO_2994 (O_2994,N_49123,N_49139);
and UO_2995 (O_2995,N_49635,N_49607);
or UO_2996 (O_2996,N_49051,N_49420);
nor UO_2997 (O_2997,N_49828,N_49087);
and UO_2998 (O_2998,N_49071,N_49168);
xnor UO_2999 (O_2999,N_49509,N_49158);
and UO_3000 (O_3000,N_49458,N_49864);
xor UO_3001 (O_3001,N_49998,N_49758);
nand UO_3002 (O_3002,N_49532,N_49729);
xor UO_3003 (O_3003,N_49443,N_49030);
nor UO_3004 (O_3004,N_49212,N_49422);
or UO_3005 (O_3005,N_49891,N_49470);
xor UO_3006 (O_3006,N_49632,N_49298);
or UO_3007 (O_3007,N_49111,N_49670);
xor UO_3008 (O_3008,N_49250,N_49144);
and UO_3009 (O_3009,N_49496,N_49113);
nor UO_3010 (O_3010,N_49361,N_49092);
nand UO_3011 (O_3011,N_49406,N_49610);
or UO_3012 (O_3012,N_49324,N_49794);
nor UO_3013 (O_3013,N_49735,N_49987);
xnor UO_3014 (O_3014,N_49718,N_49348);
xor UO_3015 (O_3015,N_49126,N_49307);
nor UO_3016 (O_3016,N_49829,N_49920);
nand UO_3017 (O_3017,N_49136,N_49989);
nor UO_3018 (O_3018,N_49075,N_49117);
nor UO_3019 (O_3019,N_49702,N_49432);
and UO_3020 (O_3020,N_49344,N_49065);
or UO_3021 (O_3021,N_49400,N_49668);
and UO_3022 (O_3022,N_49095,N_49864);
nor UO_3023 (O_3023,N_49163,N_49604);
nor UO_3024 (O_3024,N_49777,N_49340);
nand UO_3025 (O_3025,N_49164,N_49831);
and UO_3026 (O_3026,N_49941,N_49161);
xor UO_3027 (O_3027,N_49874,N_49286);
xor UO_3028 (O_3028,N_49028,N_49514);
nor UO_3029 (O_3029,N_49596,N_49905);
or UO_3030 (O_3030,N_49950,N_49937);
or UO_3031 (O_3031,N_49884,N_49894);
nor UO_3032 (O_3032,N_49325,N_49788);
and UO_3033 (O_3033,N_49042,N_49444);
and UO_3034 (O_3034,N_49671,N_49828);
xnor UO_3035 (O_3035,N_49367,N_49171);
nand UO_3036 (O_3036,N_49365,N_49950);
nand UO_3037 (O_3037,N_49758,N_49790);
and UO_3038 (O_3038,N_49663,N_49185);
and UO_3039 (O_3039,N_49219,N_49796);
nand UO_3040 (O_3040,N_49649,N_49840);
or UO_3041 (O_3041,N_49550,N_49852);
nand UO_3042 (O_3042,N_49211,N_49298);
nand UO_3043 (O_3043,N_49439,N_49341);
nor UO_3044 (O_3044,N_49057,N_49445);
or UO_3045 (O_3045,N_49338,N_49116);
or UO_3046 (O_3046,N_49431,N_49310);
xor UO_3047 (O_3047,N_49317,N_49112);
nor UO_3048 (O_3048,N_49082,N_49108);
nand UO_3049 (O_3049,N_49970,N_49413);
xor UO_3050 (O_3050,N_49252,N_49736);
nor UO_3051 (O_3051,N_49879,N_49442);
nand UO_3052 (O_3052,N_49262,N_49020);
xnor UO_3053 (O_3053,N_49983,N_49026);
or UO_3054 (O_3054,N_49445,N_49392);
nor UO_3055 (O_3055,N_49012,N_49203);
xnor UO_3056 (O_3056,N_49798,N_49731);
nand UO_3057 (O_3057,N_49511,N_49214);
and UO_3058 (O_3058,N_49189,N_49382);
and UO_3059 (O_3059,N_49398,N_49603);
or UO_3060 (O_3060,N_49324,N_49205);
xor UO_3061 (O_3061,N_49451,N_49938);
or UO_3062 (O_3062,N_49154,N_49145);
nand UO_3063 (O_3063,N_49077,N_49604);
and UO_3064 (O_3064,N_49112,N_49163);
or UO_3065 (O_3065,N_49665,N_49821);
nand UO_3066 (O_3066,N_49629,N_49571);
or UO_3067 (O_3067,N_49529,N_49586);
nand UO_3068 (O_3068,N_49301,N_49254);
xnor UO_3069 (O_3069,N_49251,N_49418);
xor UO_3070 (O_3070,N_49133,N_49170);
or UO_3071 (O_3071,N_49103,N_49296);
nor UO_3072 (O_3072,N_49264,N_49321);
nor UO_3073 (O_3073,N_49841,N_49012);
xor UO_3074 (O_3074,N_49570,N_49796);
nand UO_3075 (O_3075,N_49481,N_49190);
xor UO_3076 (O_3076,N_49363,N_49594);
or UO_3077 (O_3077,N_49583,N_49474);
xor UO_3078 (O_3078,N_49335,N_49084);
and UO_3079 (O_3079,N_49320,N_49584);
and UO_3080 (O_3080,N_49333,N_49514);
and UO_3081 (O_3081,N_49583,N_49598);
nand UO_3082 (O_3082,N_49749,N_49977);
xnor UO_3083 (O_3083,N_49452,N_49962);
and UO_3084 (O_3084,N_49233,N_49164);
nand UO_3085 (O_3085,N_49158,N_49375);
xnor UO_3086 (O_3086,N_49676,N_49134);
or UO_3087 (O_3087,N_49025,N_49575);
nor UO_3088 (O_3088,N_49026,N_49683);
nand UO_3089 (O_3089,N_49884,N_49259);
nor UO_3090 (O_3090,N_49996,N_49445);
nand UO_3091 (O_3091,N_49102,N_49196);
nand UO_3092 (O_3092,N_49294,N_49993);
xnor UO_3093 (O_3093,N_49432,N_49132);
and UO_3094 (O_3094,N_49503,N_49790);
and UO_3095 (O_3095,N_49789,N_49727);
xnor UO_3096 (O_3096,N_49108,N_49064);
nand UO_3097 (O_3097,N_49946,N_49295);
nand UO_3098 (O_3098,N_49071,N_49843);
nand UO_3099 (O_3099,N_49811,N_49118);
xor UO_3100 (O_3100,N_49054,N_49213);
or UO_3101 (O_3101,N_49106,N_49352);
or UO_3102 (O_3102,N_49425,N_49099);
or UO_3103 (O_3103,N_49297,N_49990);
xor UO_3104 (O_3104,N_49524,N_49476);
and UO_3105 (O_3105,N_49497,N_49338);
and UO_3106 (O_3106,N_49166,N_49985);
and UO_3107 (O_3107,N_49259,N_49624);
xnor UO_3108 (O_3108,N_49505,N_49113);
xnor UO_3109 (O_3109,N_49465,N_49012);
or UO_3110 (O_3110,N_49680,N_49876);
nand UO_3111 (O_3111,N_49286,N_49339);
or UO_3112 (O_3112,N_49151,N_49593);
or UO_3113 (O_3113,N_49581,N_49341);
nor UO_3114 (O_3114,N_49278,N_49990);
xnor UO_3115 (O_3115,N_49617,N_49537);
nor UO_3116 (O_3116,N_49069,N_49729);
xnor UO_3117 (O_3117,N_49473,N_49906);
or UO_3118 (O_3118,N_49208,N_49773);
and UO_3119 (O_3119,N_49523,N_49708);
or UO_3120 (O_3120,N_49753,N_49961);
or UO_3121 (O_3121,N_49916,N_49856);
or UO_3122 (O_3122,N_49876,N_49216);
nand UO_3123 (O_3123,N_49834,N_49574);
xor UO_3124 (O_3124,N_49029,N_49835);
nand UO_3125 (O_3125,N_49466,N_49579);
xnor UO_3126 (O_3126,N_49992,N_49062);
xnor UO_3127 (O_3127,N_49891,N_49184);
xor UO_3128 (O_3128,N_49465,N_49235);
nand UO_3129 (O_3129,N_49576,N_49058);
and UO_3130 (O_3130,N_49653,N_49464);
and UO_3131 (O_3131,N_49584,N_49692);
nor UO_3132 (O_3132,N_49987,N_49807);
nor UO_3133 (O_3133,N_49574,N_49689);
xnor UO_3134 (O_3134,N_49108,N_49198);
or UO_3135 (O_3135,N_49960,N_49399);
or UO_3136 (O_3136,N_49965,N_49960);
xnor UO_3137 (O_3137,N_49532,N_49075);
xnor UO_3138 (O_3138,N_49529,N_49267);
nand UO_3139 (O_3139,N_49034,N_49700);
or UO_3140 (O_3140,N_49781,N_49654);
or UO_3141 (O_3141,N_49695,N_49140);
nor UO_3142 (O_3142,N_49923,N_49374);
nand UO_3143 (O_3143,N_49527,N_49165);
xor UO_3144 (O_3144,N_49541,N_49834);
nand UO_3145 (O_3145,N_49170,N_49331);
nand UO_3146 (O_3146,N_49155,N_49949);
nand UO_3147 (O_3147,N_49598,N_49775);
and UO_3148 (O_3148,N_49067,N_49532);
xnor UO_3149 (O_3149,N_49619,N_49638);
and UO_3150 (O_3150,N_49563,N_49691);
xor UO_3151 (O_3151,N_49648,N_49469);
xor UO_3152 (O_3152,N_49373,N_49165);
nor UO_3153 (O_3153,N_49409,N_49160);
xor UO_3154 (O_3154,N_49648,N_49894);
xnor UO_3155 (O_3155,N_49161,N_49141);
and UO_3156 (O_3156,N_49923,N_49815);
nor UO_3157 (O_3157,N_49702,N_49570);
nor UO_3158 (O_3158,N_49042,N_49289);
or UO_3159 (O_3159,N_49733,N_49250);
or UO_3160 (O_3160,N_49032,N_49314);
nand UO_3161 (O_3161,N_49346,N_49097);
nor UO_3162 (O_3162,N_49213,N_49877);
nor UO_3163 (O_3163,N_49361,N_49380);
and UO_3164 (O_3164,N_49143,N_49608);
nand UO_3165 (O_3165,N_49833,N_49692);
or UO_3166 (O_3166,N_49230,N_49905);
nor UO_3167 (O_3167,N_49327,N_49943);
or UO_3168 (O_3168,N_49730,N_49009);
and UO_3169 (O_3169,N_49754,N_49559);
xor UO_3170 (O_3170,N_49853,N_49715);
xor UO_3171 (O_3171,N_49947,N_49425);
and UO_3172 (O_3172,N_49619,N_49709);
nor UO_3173 (O_3173,N_49018,N_49491);
xor UO_3174 (O_3174,N_49056,N_49526);
and UO_3175 (O_3175,N_49608,N_49139);
nor UO_3176 (O_3176,N_49728,N_49405);
nor UO_3177 (O_3177,N_49447,N_49530);
or UO_3178 (O_3178,N_49975,N_49730);
or UO_3179 (O_3179,N_49582,N_49681);
and UO_3180 (O_3180,N_49704,N_49341);
nand UO_3181 (O_3181,N_49380,N_49559);
xnor UO_3182 (O_3182,N_49836,N_49507);
or UO_3183 (O_3183,N_49230,N_49185);
nand UO_3184 (O_3184,N_49633,N_49125);
nor UO_3185 (O_3185,N_49681,N_49876);
and UO_3186 (O_3186,N_49287,N_49726);
nor UO_3187 (O_3187,N_49819,N_49717);
xor UO_3188 (O_3188,N_49810,N_49129);
or UO_3189 (O_3189,N_49788,N_49081);
nand UO_3190 (O_3190,N_49231,N_49441);
nor UO_3191 (O_3191,N_49771,N_49585);
and UO_3192 (O_3192,N_49919,N_49768);
nor UO_3193 (O_3193,N_49479,N_49098);
nand UO_3194 (O_3194,N_49568,N_49411);
nand UO_3195 (O_3195,N_49887,N_49978);
nor UO_3196 (O_3196,N_49041,N_49525);
nand UO_3197 (O_3197,N_49288,N_49430);
xor UO_3198 (O_3198,N_49860,N_49321);
or UO_3199 (O_3199,N_49501,N_49154);
or UO_3200 (O_3200,N_49737,N_49948);
xor UO_3201 (O_3201,N_49318,N_49816);
or UO_3202 (O_3202,N_49416,N_49716);
nor UO_3203 (O_3203,N_49110,N_49361);
and UO_3204 (O_3204,N_49727,N_49987);
nor UO_3205 (O_3205,N_49702,N_49427);
and UO_3206 (O_3206,N_49767,N_49931);
nand UO_3207 (O_3207,N_49407,N_49887);
or UO_3208 (O_3208,N_49619,N_49626);
and UO_3209 (O_3209,N_49403,N_49570);
and UO_3210 (O_3210,N_49680,N_49499);
nand UO_3211 (O_3211,N_49555,N_49048);
nand UO_3212 (O_3212,N_49631,N_49459);
or UO_3213 (O_3213,N_49202,N_49739);
and UO_3214 (O_3214,N_49374,N_49178);
and UO_3215 (O_3215,N_49974,N_49487);
nand UO_3216 (O_3216,N_49651,N_49327);
or UO_3217 (O_3217,N_49806,N_49610);
and UO_3218 (O_3218,N_49414,N_49502);
xnor UO_3219 (O_3219,N_49890,N_49226);
or UO_3220 (O_3220,N_49148,N_49161);
nand UO_3221 (O_3221,N_49714,N_49442);
and UO_3222 (O_3222,N_49284,N_49635);
or UO_3223 (O_3223,N_49455,N_49214);
or UO_3224 (O_3224,N_49862,N_49380);
nand UO_3225 (O_3225,N_49194,N_49720);
or UO_3226 (O_3226,N_49212,N_49370);
xor UO_3227 (O_3227,N_49640,N_49213);
nor UO_3228 (O_3228,N_49456,N_49674);
xor UO_3229 (O_3229,N_49511,N_49041);
and UO_3230 (O_3230,N_49745,N_49721);
xnor UO_3231 (O_3231,N_49325,N_49782);
nand UO_3232 (O_3232,N_49449,N_49616);
nand UO_3233 (O_3233,N_49169,N_49600);
nor UO_3234 (O_3234,N_49272,N_49902);
or UO_3235 (O_3235,N_49643,N_49364);
nand UO_3236 (O_3236,N_49386,N_49453);
nor UO_3237 (O_3237,N_49561,N_49430);
and UO_3238 (O_3238,N_49550,N_49673);
xor UO_3239 (O_3239,N_49355,N_49669);
or UO_3240 (O_3240,N_49578,N_49917);
nand UO_3241 (O_3241,N_49340,N_49301);
nor UO_3242 (O_3242,N_49289,N_49703);
nand UO_3243 (O_3243,N_49497,N_49843);
nor UO_3244 (O_3244,N_49396,N_49771);
xor UO_3245 (O_3245,N_49932,N_49522);
or UO_3246 (O_3246,N_49341,N_49880);
and UO_3247 (O_3247,N_49807,N_49914);
xor UO_3248 (O_3248,N_49757,N_49449);
nor UO_3249 (O_3249,N_49148,N_49871);
nor UO_3250 (O_3250,N_49047,N_49425);
nor UO_3251 (O_3251,N_49745,N_49776);
nor UO_3252 (O_3252,N_49112,N_49198);
nand UO_3253 (O_3253,N_49687,N_49115);
nor UO_3254 (O_3254,N_49507,N_49645);
xnor UO_3255 (O_3255,N_49816,N_49671);
xnor UO_3256 (O_3256,N_49751,N_49408);
or UO_3257 (O_3257,N_49845,N_49585);
and UO_3258 (O_3258,N_49743,N_49231);
nand UO_3259 (O_3259,N_49862,N_49244);
or UO_3260 (O_3260,N_49548,N_49148);
nor UO_3261 (O_3261,N_49907,N_49545);
nand UO_3262 (O_3262,N_49523,N_49855);
xnor UO_3263 (O_3263,N_49007,N_49748);
nor UO_3264 (O_3264,N_49802,N_49276);
nor UO_3265 (O_3265,N_49802,N_49497);
xnor UO_3266 (O_3266,N_49918,N_49408);
and UO_3267 (O_3267,N_49103,N_49683);
and UO_3268 (O_3268,N_49246,N_49770);
or UO_3269 (O_3269,N_49289,N_49049);
and UO_3270 (O_3270,N_49363,N_49723);
xnor UO_3271 (O_3271,N_49526,N_49720);
and UO_3272 (O_3272,N_49291,N_49620);
xor UO_3273 (O_3273,N_49284,N_49329);
nand UO_3274 (O_3274,N_49275,N_49217);
nor UO_3275 (O_3275,N_49632,N_49228);
nor UO_3276 (O_3276,N_49922,N_49924);
nand UO_3277 (O_3277,N_49588,N_49722);
xnor UO_3278 (O_3278,N_49275,N_49819);
nand UO_3279 (O_3279,N_49603,N_49770);
or UO_3280 (O_3280,N_49928,N_49949);
or UO_3281 (O_3281,N_49219,N_49390);
xor UO_3282 (O_3282,N_49295,N_49144);
xnor UO_3283 (O_3283,N_49211,N_49674);
nor UO_3284 (O_3284,N_49484,N_49656);
nand UO_3285 (O_3285,N_49458,N_49365);
nor UO_3286 (O_3286,N_49935,N_49799);
and UO_3287 (O_3287,N_49351,N_49495);
nor UO_3288 (O_3288,N_49446,N_49096);
or UO_3289 (O_3289,N_49173,N_49252);
and UO_3290 (O_3290,N_49066,N_49975);
nor UO_3291 (O_3291,N_49122,N_49351);
or UO_3292 (O_3292,N_49297,N_49750);
or UO_3293 (O_3293,N_49245,N_49020);
or UO_3294 (O_3294,N_49114,N_49447);
xor UO_3295 (O_3295,N_49492,N_49433);
nand UO_3296 (O_3296,N_49249,N_49459);
or UO_3297 (O_3297,N_49527,N_49248);
and UO_3298 (O_3298,N_49683,N_49285);
nand UO_3299 (O_3299,N_49646,N_49512);
xor UO_3300 (O_3300,N_49171,N_49853);
nand UO_3301 (O_3301,N_49420,N_49863);
nand UO_3302 (O_3302,N_49540,N_49975);
nor UO_3303 (O_3303,N_49299,N_49845);
xnor UO_3304 (O_3304,N_49832,N_49933);
or UO_3305 (O_3305,N_49011,N_49707);
nand UO_3306 (O_3306,N_49903,N_49975);
xnor UO_3307 (O_3307,N_49723,N_49583);
or UO_3308 (O_3308,N_49213,N_49804);
nor UO_3309 (O_3309,N_49820,N_49856);
nand UO_3310 (O_3310,N_49854,N_49943);
xor UO_3311 (O_3311,N_49441,N_49162);
xor UO_3312 (O_3312,N_49991,N_49296);
nand UO_3313 (O_3313,N_49914,N_49939);
xnor UO_3314 (O_3314,N_49548,N_49123);
or UO_3315 (O_3315,N_49585,N_49013);
or UO_3316 (O_3316,N_49118,N_49574);
xor UO_3317 (O_3317,N_49301,N_49347);
and UO_3318 (O_3318,N_49369,N_49786);
or UO_3319 (O_3319,N_49617,N_49705);
nand UO_3320 (O_3320,N_49171,N_49378);
and UO_3321 (O_3321,N_49066,N_49083);
and UO_3322 (O_3322,N_49934,N_49067);
xor UO_3323 (O_3323,N_49360,N_49751);
nand UO_3324 (O_3324,N_49677,N_49617);
xnor UO_3325 (O_3325,N_49410,N_49969);
nor UO_3326 (O_3326,N_49999,N_49333);
or UO_3327 (O_3327,N_49567,N_49047);
nor UO_3328 (O_3328,N_49218,N_49389);
xor UO_3329 (O_3329,N_49286,N_49046);
nand UO_3330 (O_3330,N_49399,N_49102);
nand UO_3331 (O_3331,N_49645,N_49673);
and UO_3332 (O_3332,N_49112,N_49012);
or UO_3333 (O_3333,N_49892,N_49836);
or UO_3334 (O_3334,N_49226,N_49503);
nor UO_3335 (O_3335,N_49948,N_49650);
xor UO_3336 (O_3336,N_49011,N_49212);
and UO_3337 (O_3337,N_49771,N_49223);
xnor UO_3338 (O_3338,N_49955,N_49133);
xor UO_3339 (O_3339,N_49636,N_49399);
nand UO_3340 (O_3340,N_49780,N_49331);
and UO_3341 (O_3341,N_49686,N_49369);
xor UO_3342 (O_3342,N_49552,N_49639);
nor UO_3343 (O_3343,N_49003,N_49140);
xor UO_3344 (O_3344,N_49232,N_49908);
nor UO_3345 (O_3345,N_49266,N_49381);
and UO_3346 (O_3346,N_49386,N_49177);
and UO_3347 (O_3347,N_49391,N_49549);
and UO_3348 (O_3348,N_49881,N_49878);
nand UO_3349 (O_3349,N_49501,N_49981);
nor UO_3350 (O_3350,N_49833,N_49142);
or UO_3351 (O_3351,N_49360,N_49136);
nand UO_3352 (O_3352,N_49337,N_49057);
nand UO_3353 (O_3353,N_49497,N_49288);
or UO_3354 (O_3354,N_49774,N_49882);
nand UO_3355 (O_3355,N_49230,N_49741);
and UO_3356 (O_3356,N_49148,N_49162);
xnor UO_3357 (O_3357,N_49990,N_49685);
nor UO_3358 (O_3358,N_49937,N_49729);
or UO_3359 (O_3359,N_49150,N_49470);
xor UO_3360 (O_3360,N_49361,N_49068);
nand UO_3361 (O_3361,N_49461,N_49407);
or UO_3362 (O_3362,N_49826,N_49699);
or UO_3363 (O_3363,N_49297,N_49768);
or UO_3364 (O_3364,N_49410,N_49727);
nor UO_3365 (O_3365,N_49264,N_49436);
and UO_3366 (O_3366,N_49833,N_49504);
xor UO_3367 (O_3367,N_49134,N_49138);
or UO_3368 (O_3368,N_49702,N_49343);
xnor UO_3369 (O_3369,N_49154,N_49663);
xnor UO_3370 (O_3370,N_49887,N_49939);
xor UO_3371 (O_3371,N_49462,N_49808);
and UO_3372 (O_3372,N_49245,N_49686);
and UO_3373 (O_3373,N_49088,N_49800);
and UO_3374 (O_3374,N_49807,N_49867);
or UO_3375 (O_3375,N_49800,N_49807);
xor UO_3376 (O_3376,N_49422,N_49145);
nand UO_3377 (O_3377,N_49451,N_49795);
nand UO_3378 (O_3378,N_49452,N_49186);
or UO_3379 (O_3379,N_49394,N_49908);
xnor UO_3380 (O_3380,N_49039,N_49032);
nand UO_3381 (O_3381,N_49543,N_49571);
nor UO_3382 (O_3382,N_49997,N_49977);
nor UO_3383 (O_3383,N_49950,N_49224);
and UO_3384 (O_3384,N_49785,N_49269);
xnor UO_3385 (O_3385,N_49462,N_49021);
nand UO_3386 (O_3386,N_49473,N_49323);
nand UO_3387 (O_3387,N_49718,N_49225);
or UO_3388 (O_3388,N_49073,N_49888);
and UO_3389 (O_3389,N_49952,N_49762);
nor UO_3390 (O_3390,N_49695,N_49434);
xor UO_3391 (O_3391,N_49451,N_49716);
xor UO_3392 (O_3392,N_49907,N_49899);
nand UO_3393 (O_3393,N_49061,N_49127);
nor UO_3394 (O_3394,N_49841,N_49606);
or UO_3395 (O_3395,N_49151,N_49174);
nor UO_3396 (O_3396,N_49073,N_49396);
or UO_3397 (O_3397,N_49304,N_49199);
nand UO_3398 (O_3398,N_49983,N_49593);
nand UO_3399 (O_3399,N_49797,N_49082);
xor UO_3400 (O_3400,N_49513,N_49634);
nand UO_3401 (O_3401,N_49533,N_49262);
nand UO_3402 (O_3402,N_49717,N_49829);
nor UO_3403 (O_3403,N_49495,N_49048);
nor UO_3404 (O_3404,N_49883,N_49840);
or UO_3405 (O_3405,N_49860,N_49429);
and UO_3406 (O_3406,N_49635,N_49883);
xnor UO_3407 (O_3407,N_49566,N_49158);
xnor UO_3408 (O_3408,N_49663,N_49800);
and UO_3409 (O_3409,N_49003,N_49409);
xor UO_3410 (O_3410,N_49272,N_49508);
and UO_3411 (O_3411,N_49272,N_49911);
nor UO_3412 (O_3412,N_49591,N_49132);
nor UO_3413 (O_3413,N_49074,N_49009);
xnor UO_3414 (O_3414,N_49892,N_49042);
nor UO_3415 (O_3415,N_49424,N_49179);
xnor UO_3416 (O_3416,N_49423,N_49726);
and UO_3417 (O_3417,N_49568,N_49808);
and UO_3418 (O_3418,N_49548,N_49149);
nand UO_3419 (O_3419,N_49169,N_49501);
nand UO_3420 (O_3420,N_49640,N_49608);
nor UO_3421 (O_3421,N_49674,N_49128);
or UO_3422 (O_3422,N_49052,N_49794);
and UO_3423 (O_3423,N_49170,N_49343);
nand UO_3424 (O_3424,N_49741,N_49526);
or UO_3425 (O_3425,N_49811,N_49036);
and UO_3426 (O_3426,N_49762,N_49668);
nand UO_3427 (O_3427,N_49871,N_49669);
or UO_3428 (O_3428,N_49025,N_49527);
nand UO_3429 (O_3429,N_49532,N_49786);
nand UO_3430 (O_3430,N_49763,N_49574);
nand UO_3431 (O_3431,N_49919,N_49101);
and UO_3432 (O_3432,N_49131,N_49658);
xnor UO_3433 (O_3433,N_49937,N_49815);
nand UO_3434 (O_3434,N_49619,N_49191);
nand UO_3435 (O_3435,N_49004,N_49558);
nand UO_3436 (O_3436,N_49182,N_49014);
xor UO_3437 (O_3437,N_49645,N_49040);
nor UO_3438 (O_3438,N_49095,N_49297);
xor UO_3439 (O_3439,N_49331,N_49149);
nand UO_3440 (O_3440,N_49794,N_49185);
xnor UO_3441 (O_3441,N_49647,N_49198);
or UO_3442 (O_3442,N_49733,N_49631);
and UO_3443 (O_3443,N_49199,N_49279);
or UO_3444 (O_3444,N_49381,N_49396);
xnor UO_3445 (O_3445,N_49024,N_49488);
or UO_3446 (O_3446,N_49763,N_49908);
and UO_3447 (O_3447,N_49648,N_49492);
nand UO_3448 (O_3448,N_49005,N_49650);
nor UO_3449 (O_3449,N_49248,N_49714);
and UO_3450 (O_3450,N_49385,N_49994);
and UO_3451 (O_3451,N_49729,N_49561);
and UO_3452 (O_3452,N_49768,N_49190);
nor UO_3453 (O_3453,N_49748,N_49759);
or UO_3454 (O_3454,N_49170,N_49269);
nor UO_3455 (O_3455,N_49594,N_49974);
xnor UO_3456 (O_3456,N_49679,N_49771);
nor UO_3457 (O_3457,N_49321,N_49587);
nor UO_3458 (O_3458,N_49561,N_49030);
xnor UO_3459 (O_3459,N_49940,N_49561);
nand UO_3460 (O_3460,N_49178,N_49929);
nor UO_3461 (O_3461,N_49262,N_49135);
nand UO_3462 (O_3462,N_49646,N_49950);
and UO_3463 (O_3463,N_49781,N_49752);
xor UO_3464 (O_3464,N_49137,N_49843);
nor UO_3465 (O_3465,N_49298,N_49380);
nand UO_3466 (O_3466,N_49000,N_49057);
nand UO_3467 (O_3467,N_49358,N_49025);
or UO_3468 (O_3468,N_49281,N_49947);
nor UO_3469 (O_3469,N_49684,N_49775);
nor UO_3470 (O_3470,N_49209,N_49650);
nor UO_3471 (O_3471,N_49370,N_49356);
and UO_3472 (O_3472,N_49593,N_49253);
nand UO_3473 (O_3473,N_49480,N_49428);
nor UO_3474 (O_3474,N_49428,N_49376);
or UO_3475 (O_3475,N_49811,N_49573);
nor UO_3476 (O_3476,N_49513,N_49102);
nand UO_3477 (O_3477,N_49283,N_49837);
xnor UO_3478 (O_3478,N_49575,N_49599);
or UO_3479 (O_3479,N_49369,N_49214);
and UO_3480 (O_3480,N_49739,N_49420);
and UO_3481 (O_3481,N_49395,N_49864);
nand UO_3482 (O_3482,N_49510,N_49586);
nand UO_3483 (O_3483,N_49282,N_49640);
xnor UO_3484 (O_3484,N_49249,N_49764);
xnor UO_3485 (O_3485,N_49873,N_49751);
and UO_3486 (O_3486,N_49845,N_49551);
or UO_3487 (O_3487,N_49078,N_49759);
and UO_3488 (O_3488,N_49791,N_49885);
and UO_3489 (O_3489,N_49704,N_49755);
xnor UO_3490 (O_3490,N_49549,N_49942);
and UO_3491 (O_3491,N_49023,N_49287);
xor UO_3492 (O_3492,N_49373,N_49843);
nand UO_3493 (O_3493,N_49894,N_49834);
xnor UO_3494 (O_3494,N_49104,N_49178);
and UO_3495 (O_3495,N_49817,N_49889);
nand UO_3496 (O_3496,N_49060,N_49770);
or UO_3497 (O_3497,N_49989,N_49228);
and UO_3498 (O_3498,N_49682,N_49691);
nand UO_3499 (O_3499,N_49522,N_49714);
nand UO_3500 (O_3500,N_49238,N_49141);
or UO_3501 (O_3501,N_49921,N_49872);
xnor UO_3502 (O_3502,N_49634,N_49631);
and UO_3503 (O_3503,N_49788,N_49823);
xor UO_3504 (O_3504,N_49285,N_49796);
and UO_3505 (O_3505,N_49064,N_49859);
or UO_3506 (O_3506,N_49531,N_49710);
or UO_3507 (O_3507,N_49432,N_49806);
or UO_3508 (O_3508,N_49536,N_49517);
and UO_3509 (O_3509,N_49690,N_49166);
and UO_3510 (O_3510,N_49170,N_49175);
and UO_3511 (O_3511,N_49554,N_49534);
nand UO_3512 (O_3512,N_49345,N_49520);
xnor UO_3513 (O_3513,N_49023,N_49971);
and UO_3514 (O_3514,N_49485,N_49431);
and UO_3515 (O_3515,N_49930,N_49107);
xnor UO_3516 (O_3516,N_49679,N_49692);
nor UO_3517 (O_3517,N_49426,N_49008);
nand UO_3518 (O_3518,N_49906,N_49566);
nor UO_3519 (O_3519,N_49938,N_49566);
nor UO_3520 (O_3520,N_49532,N_49999);
nand UO_3521 (O_3521,N_49461,N_49723);
and UO_3522 (O_3522,N_49209,N_49352);
and UO_3523 (O_3523,N_49014,N_49187);
nor UO_3524 (O_3524,N_49663,N_49474);
and UO_3525 (O_3525,N_49096,N_49128);
or UO_3526 (O_3526,N_49847,N_49679);
and UO_3527 (O_3527,N_49253,N_49854);
xor UO_3528 (O_3528,N_49271,N_49575);
nand UO_3529 (O_3529,N_49987,N_49863);
or UO_3530 (O_3530,N_49788,N_49663);
xnor UO_3531 (O_3531,N_49023,N_49751);
nand UO_3532 (O_3532,N_49121,N_49788);
nand UO_3533 (O_3533,N_49178,N_49031);
xor UO_3534 (O_3534,N_49845,N_49614);
nor UO_3535 (O_3535,N_49709,N_49395);
xnor UO_3536 (O_3536,N_49847,N_49218);
or UO_3537 (O_3537,N_49965,N_49349);
nand UO_3538 (O_3538,N_49950,N_49374);
nand UO_3539 (O_3539,N_49717,N_49431);
nand UO_3540 (O_3540,N_49018,N_49484);
nor UO_3541 (O_3541,N_49790,N_49080);
nor UO_3542 (O_3542,N_49585,N_49245);
nand UO_3543 (O_3543,N_49120,N_49941);
or UO_3544 (O_3544,N_49116,N_49057);
nor UO_3545 (O_3545,N_49602,N_49095);
and UO_3546 (O_3546,N_49284,N_49668);
or UO_3547 (O_3547,N_49864,N_49810);
nand UO_3548 (O_3548,N_49622,N_49145);
and UO_3549 (O_3549,N_49677,N_49250);
and UO_3550 (O_3550,N_49150,N_49362);
nor UO_3551 (O_3551,N_49193,N_49409);
nand UO_3552 (O_3552,N_49793,N_49442);
xor UO_3553 (O_3553,N_49976,N_49610);
or UO_3554 (O_3554,N_49501,N_49804);
xor UO_3555 (O_3555,N_49731,N_49445);
and UO_3556 (O_3556,N_49315,N_49642);
nand UO_3557 (O_3557,N_49562,N_49852);
nand UO_3558 (O_3558,N_49886,N_49943);
and UO_3559 (O_3559,N_49234,N_49801);
xnor UO_3560 (O_3560,N_49264,N_49169);
nand UO_3561 (O_3561,N_49953,N_49587);
or UO_3562 (O_3562,N_49466,N_49559);
and UO_3563 (O_3563,N_49567,N_49097);
and UO_3564 (O_3564,N_49575,N_49070);
and UO_3565 (O_3565,N_49796,N_49271);
and UO_3566 (O_3566,N_49168,N_49046);
nor UO_3567 (O_3567,N_49037,N_49545);
xor UO_3568 (O_3568,N_49393,N_49276);
or UO_3569 (O_3569,N_49577,N_49146);
or UO_3570 (O_3570,N_49299,N_49452);
or UO_3571 (O_3571,N_49835,N_49131);
xnor UO_3572 (O_3572,N_49557,N_49770);
and UO_3573 (O_3573,N_49259,N_49879);
nor UO_3574 (O_3574,N_49408,N_49967);
and UO_3575 (O_3575,N_49402,N_49724);
nor UO_3576 (O_3576,N_49251,N_49145);
nand UO_3577 (O_3577,N_49647,N_49863);
nand UO_3578 (O_3578,N_49526,N_49908);
nor UO_3579 (O_3579,N_49629,N_49698);
or UO_3580 (O_3580,N_49422,N_49898);
xor UO_3581 (O_3581,N_49438,N_49233);
xnor UO_3582 (O_3582,N_49076,N_49180);
nand UO_3583 (O_3583,N_49649,N_49607);
nand UO_3584 (O_3584,N_49392,N_49450);
and UO_3585 (O_3585,N_49702,N_49953);
xor UO_3586 (O_3586,N_49658,N_49298);
and UO_3587 (O_3587,N_49542,N_49105);
nand UO_3588 (O_3588,N_49362,N_49837);
and UO_3589 (O_3589,N_49059,N_49470);
or UO_3590 (O_3590,N_49634,N_49183);
nand UO_3591 (O_3591,N_49748,N_49069);
xor UO_3592 (O_3592,N_49288,N_49975);
nand UO_3593 (O_3593,N_49190,N_49320);
nand UO_3594 (O_3594,N_49253,N_49298);
and UO_3595 (O_3595,N_49003,N_49781);
xor UO_3596 (O_3596,N_49850,N_49019);
nor UO_3597 (O_3597,N_49887,N_49873);
nand UO_3598 (O_3598,N_49913,N_49349);
or UO_3599 (O_3599,N_49948,N_49693);
nor UO_3600 (O_3600,N_49476,N_49954);
or UO_3601 (O_3601,N_49681,N_49812);
or UO_3602 (O_3602,N_49122,N_49833);
nor UO_3603 (O_3603,N_49885,N_49270);
xor UO_3604 (O_3604,N_49906,N_49363);
nor UO_3605 (O_3605,N_49957,N_49265);
and UO_3606 (O_3606,N_49832,N_49757);
xnor UO_3607 (O_3607,N_49515,N_49724);
xnor UO_3608 (O_3608,N_49415,N_49984);
and UO_3609 (O_3609,N_49618,N_49260);
nand UO_3610 (O_3610,N_49687,N_49697);
and UO_3611 (O_3611,N_49481,N_49395);
or UO_3612 (O_3612,N_49718,N_49390);
or UO_3613 (O_3613,N_49725,N_49532);
nor UO_3614 (O_3614,N_49044,N_49225);
or UO_3615 (O_3615,N_49022,N_49986);
and UO_3616 (O_3616,N_49738,N_49505);
and UO_3617 (O_3617,N_49035,N_49275);
and UO_3618 (O_3618,N_49970,N_49179);
xnor UO_3619 (O_3619,N_49200,N_49115);
nor UO_3620 (O_3620,N_49194,N_49449);
and UO_3621 (O_3621,N_49353,N_49411);
and UO_3622 (O_3622,N_49105,N_49856);
nor UO_3623 (O_3623,N_49457,N_49715);
xnor UO_3624 (O_3624,N_49114,N_49754);
and UO_3625 (O_3625,N_49019,N_49902);
xor UO_3626 (O_3626,N_49445,N_49345);
or UO_3627 (O_3627,N_49405,N_49167);
or UO_3628 (O_3628,N_49287,N_49365);
or UO_3629 (O_3629,N_49494,N_49636);
xor UO_3630 (O_3630,N_49723,N_49285);
nand UO_3631 (O_3631,N_49077,N_49486);
nand UO_3632 (O_3632,N_49821,N_49811);
nand UO_3633 (O_3633,N_49389,N_49773);
nand UO_3634 (O_3634,N_49225,N_49467);
or UO_3635 (O_3635,N_49606,N_49584);
nor UO_3636 (O_3636,N_49497,N_49056);
and UO_3637 (O_3637,N_49111,N_49675);
and UO_3638 (O_3638,N_49604,N_49928);
xor UO_3639 (O_3639,N_49074,N_49407);
and UO_3640 (O_3640,N_49924,N_49630);
and UO_3641 (O_3641,N_49732,N_49598);
xnor UO_3642 (O_3642,N_49483,N_49769);
and UO_3643 (O_3643,N_49963,N_49193);
xor UO_3644 (O_3644,N_49800,N_49287);
xor UO_3645 (O_3645,N_49422,N_49774);
and UO_3646 (O_3646,N_49819,N_49097);
nor UO_3647 (O_3647,N_49977,N_49390);
xor UO_3648 (O_3648,N_49552,N_49587);
xnor UO_3649 (O_3649,N_49174,N_49574);
xor UO_3650 (O_3650,N_49913,N_49229);
or UO_3651 (O_3651,N_49156,N_49550);
or UO_3652 (O_3652,N_49601,N_49607);
xnor UO_3653 (O_3653,N_49399,N_49577);
or UO_3654 (O_3654,N_49362,N_49185);
and UO_3655 (O_3655,N_49294,N_49158);
or UO_3656 (O_3656,N_49259,N_49153);
xnor UO_3657 (O_3657,N_49073,N_49879);
xnor UO_3658 (O_3658,N_49745,N_49242);
xor UO_3659 (O_3659,N_49185,N_49461);
xor UO_3660 (O_3660,N_49743,N_49530);
or UO_3661 (O_3661,N_49373,N_49685);
nor UO_3662 (O_3662,N_49556,N_49073);
nand UO_3663 (O_3663,N_49245,N_49185);
or UO_3664 (O_3664,N_49362,N_49633);
nor UO_3665 (O_3665,N_49026,N_49770);
or UO_3666 (O_3666,N_49883,N_49767);
nor UO_3667 (O_3667,N_49431,N_49622);
xnor UO_3668 (O_3668,N_49173,N_49226);
and UO_3669 (O_3669,N_49837,N_49479);
nor UO_3670 (O_3670,N_49116,N_49627);
nand UO_3671 (O_3671,N_49426,N_49969);
xor UO_3672 (O_3672,N_49491,N_49726);
nor UO_3673 (O_3673,N_49323,N_49810);
nor UO_3674 (O_3674,N_49324,N_49698);
or UO_3675 (O_3675,N_49321,N_49298);
nand UO_3676 (O_3676,N_49146,N_49583);
nor UO_3677 (O_3677,N_49184,N_49616);
nor UO_3678 (O_3678,N_49559,N_49551);
and UO_3679 (O_3679,N_49864,N_49429);
nor UO_3680 (O_3680,N_49638,N_49173);
nor UO_3681 (O_3681,N_49058,N_49892);
nand UO_3682 (O_3682,N_49098,N_49253);
xnor UO_3683 (O_3683,N_49603,N_49469);
nor UO_3684 (O_3684,N_49979,N_49702);
xor UO_3685 (O_3685,N_49319,N_49261);
nand UO_3686 (O_3686,N_49989,N_49265);
nor UO_3687 (O_3687,N_49896,N_49312);
nand UO_3688 (O_3688,N_49208,N_49592);
and UO_3689 (O_3689,N_49221,N_49322);
or UO_3690 (O_3690,N_49505,N_49474);
or UO_3691 (O_3691,N_49208,N_49145);
and UO_3692 (O_3692,N_49593,N_49226);
nor UO_3693 (O_3693,N_49757,N_49167);
xor UO_3694 (O_3694,N_49129,N_49277);
or UO_3695 (O_3695,N_49984,N_49077);
or UO_3696 (O_3696,N_49697,N_49763);
nand UO_3697 (O_3697,N_49831,N_49050);
nand UO_3698 (O_3698,N_49846,N_49966);
xnor UO_3699 (O_3699,N_49621,N_49270);
and UO_3700 (O_3700,N_49576,N_49744);
nor UO_3701 (O_3701,N_49810,N_49185);
nand UO_3702 (O_3702,N_49647,N_49499);
and UO_3703 (O_3703,N_49997,N_49370);
or UO_3704 (O_3704,N_49580,N_49039);
or UO_3705 (O_3705,N_49511,N_49612);
nand UO_3706 (O_3706,N_49334,N_49086);
or UO_3707 (O_3707,N_49733,N_49232);
nor UO_3708 (O_3708,N_49092,N_49866);
or UO_3709 (O_3709,N_49927,N_49693);
nor UO_3710 (O_3710,N_49556,N_49736);
and UO_3711 (O_3711,N_49046,N_49049);
xnor UO_3712 (O_3712,N_49188,N_49647);
or UO_3713 (O_3713,N_49111,N_49203);
and UO_3714 (O_3714,N_49097,N_49613);
or UO_3715 (O_3715,N_49383,N_49600);
and UO_3716 (O_3716,N_49018,N_49687);
nor UO_3717 (O_3717,N_49203,N_49335);
xor UO_3718 (O_3718,N_49402,N_49107);
and UO_3719 (O_3719,N_49799,N_49140);
nor UO_3720 (O_3720,N_49819,N_49753);
or UO_3721 (O_3721,N_49970,N_49939);
nor UO_3722 (O_3722,N_49565,N_49042);
xor UO_3723 (O_3723,N_49085,N_49703);
nand UO_3724 (O_3724,N_49894,N_49720);
and UO_3725 (O_3725,N_49844,N_49296);
xnor UO_3726 (O_3726,N_49952,N_49220);
nor UO_3727 (O_3727,N_49548,N_49974);
and UO_3728 (O_3728,N_49588,N_49318);
nor UO_3729 (O_3729,N_49210,N_49814);
xnor UO_3730 (O_3730,N_49645,N_49573);
or UO_3731 (O_3731,N_49239,N_49245);
and UO_3732 (O_3732,N_49962,N_49848);
nand UO_3733 (O_3733,N_49740,N_49631);
xor UO_3734 (O_3734,N_49818,N_49261);
or UO_3735 (O_3735,N_49449,N_49526);
nor UO_3736 (O_3736,N_49338,N_49019);
xor UO_3737 (O_3737,N_49048,N_49210);
nand UO_3738 (O_3738,N_49024,N_49253);
nand UO_3739 (O_3739,N_49472,N_49014);
and UO_3740 (O_3740,N_49286,N_49094);
nand UO_3741 (O_3741,N_49678,N_49425);
or UO_3742 (O_3742,N_49979,N_49494);
or UO_3743 (O_3743,N_49690,N_49322);
or UO_3744 (O_3744,N_49394,N_49924);
nand UO_3745 (O_3745,N_49173,N_49234);
xor UO_3746 (O_3746,N_49105,N_49137);
or UO_3747 (O_3747,N_49022,N_49545);
and UO_3748 (O_3748,N_49846,N_49224);
xnor UO_3749 (O_3749,N_49166,N_49562);
xor UO_3750 (O_3750,N_49069,N_49711);
or UO_3751 (O_3751,N_49205,N_49528);
or UO_3752 (O_3752,N_49783,N_49759);
nand UO_3753 (O_3753,N_49997,N_49725);
and UO_3754 (O_3754,N_49303,N_49807);
and UO_3755 (O_3755,N_49816,N_49288);
nand UO_3756 (O_3756,N_49361,N_49589);
xor UO_3757 (O_3757,N_49437,N_49498);
or UO_3758 (O_3758,N_49293,N_49911);
nor UO_3759 (O_3759,N_49463,N_49590);
or UO_3760 (O_3760,N_49613,N_49911);
xnor UO_3761 (O_3761,N_49855,N_49643);
and UO_3762 (O_3762,N_49282,N_49048);
or UO_3763 (O_3763,N_49747,N_49732);
nor UO_3764 (O_3764,N_49359,N_49194);
and UO_3765 (O_3765,N_49188,N_49666);
nor UO_3766 (O_3766,N_49665,N_49406);
xnor UO_3767 (O_3767,N_49299,N_49338);
or UO_3768 (O_3768,N_49165,N_49521);
nand UO_3769 (O_3769,N_49761,N_49955);
or UO_3770 (O_3770,N_49727,N_49027);
nand UO_3771 (O_3771,N_49797,N_49841);
nor UO_3772 (O_3772,N_49389,N_49417);
xor UO_3773 (O_3773,N_49099,N_49416);
xnor UO_3774 (O_3774,N_49326,N_49720);
xnor UO_3775 (O_3775,N_49935,N_49224);
xnor UO_3776 (O_3776,N_49132,N_49872);
xnor UO_3777 (O_3777,N_49759,N_49417);
and UO_3778 (O_3778,N_49070,N_49483);
xnor UO_3779 (O_3779,N_49439,N_49897);
nand UO_3780 (O_3780,N_49821,N_49261);
or UO_3781 (O_3781,N_49303,N_49437);
nand UO_3782 (O_3782,N_49873,N_49729);
xnor UO_3783 (O_3783,N_49289,N_49772);
nor UO_3784 (O_3784,N_49079,N_49533);
xnor UO_3785 (O_3785,N_49932,N_49042);
and UO_3786 (O_3786,N_49832,N_49684);
nor UO_3787 (O_3787,N_49548,N_49676);
xor UO_3788 (O_3788,N_49029,N_49523);
xor UO_3789 (O_3789,N_49597,N_49978);
or UO_3790 (O_3790,N_49047,N_49031);
xor UO_3791 (O_3791,N_49845,N_49554);
and UO_3792 (O_3792,N_49041,N_49167);
and UO_3793 (O_3793,N_49627,N_49364);
or UO_3794 (O_3794,N_49460,N_49510);
and UO_3795 (O_3795,N_49416,N_49922);
or UO_3796 (O_3796,N_49914,N_49968);
nor UO_3797 (O_3797,N_49359,N_49797);
or UO_3798 (O_3798,N_49500,N_49439);
nand UO_3799 (O_3799,N_49091,N_49877);
and UO_3800 (O_3800,N_49093,N_49450);
nor UO_3801 (O_3801,N_49641,N_49376);
or UO_3802 (O_3802,N_49699,N_49658);
and UO_3803 (O_3803,N_49901,N_49352);
xnor UO_3804 (O_3804,N_49277,N_49784);
xnor UO_3805 (O_3805,N_49168,N_49464);
and UO_3806 (O_3806,N_49074,N_49088);
xnor UO_3807 (O_3807,N_49098,N_49979);
or UO_3808 (O_3808,N_49232,N_49100);
and UO_3809 (O_3809,N_49490,N_49257);
nor UO_3810 (O_3810,N_49200,N_49211);
nor UO_3811 (O_3811,N_49105,N_49670);
xor UO_3812 (O_3812,N_49281,N_49516);
or UO_3813 (O_3813,N_49152,N_49544);
xor UO_3814 (O_3814,N_49606,N_49168);
or UO_3815 (O_3815,N_49439,N_49375);
and UO_3816 (O_3816,N_49641,N_49521);
nand UO_3817 (O_3817,N_49384,N_49188);
nor UO_3818 (O_3818,N_49692,N_49925);
nor UO_3819 (O_3819,N_49096,N_49744);
and UO_3820 (O_3820,N_49113,N_49476);
xnor UO_3821 (O_3821,N_49247,N_49748);
xor UO_3822 (O_3822,N_49612,N_49761);
nand UO_3823 (O_3823,N_49510,N_49088);
nor UO_3824 (O_3824,N_49337,N_49986);
xnor UO_3825 (O_3825,N_49840,N_49163);
nor UO_3826 (O_3826,N_49630,N_49636);
nand UO_3827 (O_3827,N_49016,N_49551);
or UO_3828 (O_3828,N_49222,N_49551);
xnor UO_3829 (O_3829,N_49531,N_49174);
xor UO_3830 (O_3830,N_49578,N_49010);
nor UO_3831 (O_3831,N_49468,N_49976);
or UO_3832 (O_3832,N_49791,N_49054);
or UO_3833 (O_3833,N_49101,N_49958);
and UO_3834 (O_3834,N_49036,N_49904);
and UO_3835 (O_3835,N_49918,N_49062);
nor UO_3836 (O_3836,N_49621,N_49535);
xor UO_3837 (O_3837,N_49536,N_49353);
and UO_3838 (O_3838,N_49773,N_49978);
and UO_3839 (O_3839,N_49542,N_49019);
and UO_3840 (O_3840,N_49531,N_49273);
or UO_3841 (O_3841,N_49799,N_49213);
or UO_3842 (O_3842,N_49118,N_49620);
nor UO_3843 (O_3843,N_49253,N_49532);
nand UO_3844 (O_3844,N_49703,N_49162);
or UO_3845 (O_3845,N_49027,N_49107);
nand UO_3846 (O_3846,N_49198,N_49565);
and UO_3847 (O_3847,N_49770,N_49450);
xnor UO_3848 (O_3848,N_49231,N_49310);
and UO_3849 (O_3849,N_49809,N_49080);
and UO_3850 (O_3850,N_49079,N_49832);
or UO_3851 (O_3851,N_49710,N_49757);
nor UO_3852 (O_3852,N_49681,N_49675);
and UO_3853 (O_3853,N_49621,N_49813);
and UO_3854 (O_3854,N_49669,N_49279);
or UO_3855 (O_3855,N_49302,N_49449);
and UO_3856 (O_3856,N_49942,N_49561);
nor UO_3857 (O_3857,N_49175,N_49758);
xor UO_3858 (O_3858,N_49186,N_49627);
nor UO_3859 (O_3859,N_49130,N_49050);
nand UO_3860 (O_3860,N_49457,N_49294);
nand UO_3861 (O_3861,N_49723,N_49134);
nor UO_3862 (O_3862,N_49806,N_49606);
and UO_3863 (O_3863,N_49825,N_49417);
or UO_3864 (O_3864,N_49841,N_49413);
and UO_3865 (O_3865,N_49102,N_49304);
nand UO_3866 (O_3866,N_49371,N_49539);
or UO_3867 (O_3867,N_49472,N_49484);
xor UO_3868 (O_3868,N_49191,N_49084);
nor UO_3869 (O_3869,N_49067,N_49836);
or UO_3870 (O_3870,N_49494,N_49139);
and UO_3871 (O_3871,N_49968,N_49102);
xor UO_3872 (O_3872,N_49183,N_49629);
and UO_3873 (O_3873,N_49589,N_49434);
xnor UO_3874 (O_3874,N_49548,N_49823);
nand UO_3875 (O_3875,N_49060,N_49268);
and UO_3876 (O_3876,N_49308,N_49412);
or UO_3877 (O_3877,N_49201,N_49200);
or UO_3878 (O_3878,N_49160,N_49633);
and UO_3879 (O_3879,N_49340,N_49883);
and UO_3880 (O_3880,N_49665,N_49023);
nand UO_3881 (O_3881,N_49568,N_49586);
and UO_3882 (O_3882,N_49184,N_49351);
nand UO_3883 (O_3883,N_49623,N_49512);
or UO_3884 (O_3884,N_49568,N_49450);
or UO_3885 (O_3885,N_49833,N_49679);
nor UO_3886 (O_3886,N_49764,N_49426);
or UO_3887 (O_3887,N_49146,N_49376);
and UO_3888 (O_3888,N_49581,N_49085);
nor UO_3889 (O_3889,N_49084,N_49662);
nand UO_3890 (O_3890,N_49789,N_49551);
or UO_3891 (O_3891,N_49399,N_49260);
nand UO_3892 (O_3892,N_49394,N_49015);
or UO_3893 (O_3893,N_49680,N_49427);
and UO_3894 (O_3894,N_49858,N_49793);
and UO_3895 (O_3895,N_49909,N_49031);
or UO_3896 (O_3896,N_49317,N_49751);
and UO_3897 (O_3897,N_49751,N_49729);
nand UO_3898 (O_3898,N_49315,N_49037);
xor UO_3899 (O_3899,N_49069,N_49763);
or UO_3900 (O_3900,N_49430,N_49366);
and UO_3901 (O_3901,N_49411,N_49177);
or UO_3902 (O_3902,N_49592,N_49443);
nand UO_3903 (O_3903,N_49741,N_49800);
xnor UO_3904 (O_3904,N_49701,N_49450);
nand UO_3905 (O_3905,N_49267,N_49082);
xnor UO_3906 (O_3906,N_49597,N_49737);
nand UO_3907 (O_3907,N_49014,N_49998);
nand UO_3908 (O_3908,N_49427,N_49774);
nand UO_3909 (O_3909,N_49405,N_49325);
nand UO_3910 (O_3910,N_49220,N_49484);
xnor UO_3911 (O_3911,N_49709,N_49603);
and UO_3912 (O_3912,N_49386,N_49696);
nand UO_3913 (O_3913,N_49694,N_49363);
xnor UO_3914 (O_3914,N_49271,N_49802);
and UO_3915 (O_3915,N_49751,N_49241);
and UO_3916 (O_3916,N_49659,N_49384);
xnor UO_3917 (O_3917,N_49408,N_49338);
and UO_3918 (O_3918,N_49892,N_49335);
nand UO_3919 (O_3919,N_49908,N_49848);
or UO_3920 (O_3920,N_49387,N_49678);
nor UO_3921 (O_3921,N_49346,N_49608);
and UO_3922 (O_3922,N_49679,N_49162);
and UO_3923 (O_3923,N_49033,N_49506);
and UO_3924 (O_3924,N_49530,N_49927);
nor UO_3925 (O_3925,N_49491,N_49588);
xnor UO_3926 (O_3926,N_49160,N_49749);
nor UO_3927 (O_3927,N_49097,N_49374);
nor UO_3928 (O_3928,N_49255,N_49323);
nor UO_3929 (O_3929,N_49781,N_49396);
and UO_3930 (O_3930,N_49602,N_49541);
and UO_3931 (O_3931,N_49610,N_49764);
xnor UO_3932 (O_3932,N_49123,N_49973);
xor UO_3933 (O_3933,N_49115,N_49489);
nand UO_3934 (O_3934,N_49941,N_49184);
nand UO_3935 (O_3935,N_49085,N_49905);
xnor UO_3936 (O_3936,N_49217,N_49683);
nand UO_3937 (O_3937,N_49116,N_49220);
or UO_3938 (O_3938,N_49653,N_49788);
or UO_3939 (O_3939,N_49739,N_49402);
xnor UO_3940 (O_3940,N_49215,N_49549);
nand UO_3941 (O_3941,N_49924,N_49923);
and UO_3942 (O_3942,N_49778,N_49730);
nor UO_3943 (O_3943,N_49987,N_49503);
xor UO_3944 (O_3944,N_49561,N_49827);
and UO_3945 (O_3945,N_49266,N_49047);
or UO_3946 (O_3946,N_49966,N_49625);
or UO_3947 (O_3947,N_49922,N_49746);
or UO_3948 (O_3948,N_49677,N_49401);
nor UO_3949 (O_3949,N_49179,N_49241);
nand UO_3950 (O_3950,N_49556,N_49528);
and UO_3951 (O_3951,N_49247,N_49212);
nor UO_3952 (O_3952,N_49706,N_49218);
nor UO_3953 (O_3953,N_49511,N_49311);
xnor UO_3954 (O_3954,N_49833,N_49600);
and UO_3955 (O_3955,N_49307,N_49271);
and UO_3956 (O_3956,N_49672,N_49952);
or UO_3957 (O_3957,N_49814,N_49466);
or UO_3958 (O_3958,N_49146,N_49871);
or UO_3959 (O_3959,N_49803,N_49452);
nand UO_3960 (O_3960,N_49333,N_49055);
or UO_3961 (O_3961,N_49678,N_49179);
and UO_3962 (O_3962,N_49203,N_49460);
xor UO_3963 (O_3963,N_49861,N_49993);
nor UO_3964 (O_3964,N_49220,N_49259);
and UO_3965 (O_3965,N_49450,N_49839);
and UO_3966 (O_3966,N_49671,N_49249);
and UO_3967 (O_3967,N_49630,N_49103);
xnor UO_3968 (O_3968,N_49364,N_49623);
nand UO_3969 (O_3969,N_49210,N_49602);
xor UO_3970 (O_3970,N_49524,N_49495);
nor UO_3971 (O_3971,N_49237,N_49778);
or UO_3972 (O_3972,N_49177,N_49449);
or UO_3973 (O_3973,N_49345,N_49706);
and UO_3974 (O_3974,N_49255,N_49375);
nor UO_3975 (O_3975,N_49739,N_49729);
xnor UO_3976 (O_3976,N_49031,N_49669);
and UO_3977 (O_3977,N_49222,N_49411);
xnor UO_3978 (O_3978,N_49686,N_49872);
and UO_3979 (O_3979,N_49055,N_49783);
and UO_3980 (O_3980,N_49833,N_49947);
nor UO_3981 (O_3981,N_49146,N_49427);
or UO_3982 (O_3982,N_49117,N_49690);
or UO_3983 (O_3983,N_49011,N_49306);
xnor UO_3984 (O_3984,N_49753,N_49597);
nor UO_3985 (O_3985,N_49881,N_49759);
nor UO_3986 (O_3986,N_49452,N_49778);
xnor UO_3987 (O_3987,N_49623,N_49980);
or UO_3988 (O_3988,N_49902,N_49661);
nor UO_3989 (O_3989,N_49424,N_49868);
xor UO_3990 (O_3990,N_49418,N_49704);
xnor UO_3991 (O_3991,N_49759,N_49815);
or UO_3992 (O_3992,N_49831,N_49018);
or UO_3993 (O_3993,N_49096,N_49857);
nand UO_3994 (O_3994,N_49182,N_49767);
nor UO_3995 (O_3995,N_49566,N_49820);
or UO_3996 (O_3996,N_49470,N_49383);
nand UO_3997 (O_3997,N_49624,N_49270);
or UO_3998 (O_3998,N_49177,N_49763);
and UO_3999 (O_3999,N_49689,N_49453);
nand UO_4000 (O_4000,N_49654,N_49370);
nor UO_4001 (O_4001,N_49786,N_49023);
nand UO_4002 (O_4002,N_49930,N_49477);
or UO_4003 (O_4003,N_49198,N_49260);
and UO_4004 (O_4004,N_49890,N_49580);
and UO_4005 (O_4005,N_49421,N_49414);
nand UO_4006 (O_4006,N_49444,N_49363);
nand UO_4007 (O_4007,N_49899,N_49598);
nor UO_4008 (O_4008,N_49221,N_49449);
or UO_4009 (O_4009,N_49468,N_49071);
nor UO_4010 (O_4010,N_49727,N_49596);
nand UO_4011 (O_4011,N_49200,N_49068);
nor UO_4012 (O_4012,N_49866,N_49181);
xor UO_4013 (O_4013,N_49700,N_49976);
nor UO_4014 (O_4014,N_49484,N_49876);
nand UO_4015 (O_4015,N_49392,N_49860);
nor UO_4016 (O_4016,N_49439,N_49577);
and UO_4017 (O_4017,N_49060,N_49552);
and UO_4018 (O_4018,N_49458,N_49824);
nand UO_4019 (O_4019,N_49511,N_49241);
nor UO_4020 (O_4020,N_49212,N_49899);
and UO_4021 (O_4021,N_49168,N_49560);
and UO_4022 (O_4022,N_49547,N_49345);
xor UO_4023 (O_4023,N_49742,N_49820);
xor UO_4024 (O_4024,N_49952,N_49512);
or UO_4025 (O_4025,N_49895,N_49016);
or UO_4026 (O_4026,N_49032,N_49584);
or UO_4027 (O_4027,N_49935,N_49149);
nand UO_4028 (O_4028,N_49617,N_49980);
and UO_4029 (O_4029,N_49208,N_49784);
nand UO_4030 (O_4030,N_49159,N_49163);
nand UO_4031 (O_4031,N_49293,N_49130);
and UO_4032 (O_4032,N_49075,N_49394);
xor UO_4033 (O_4033,N_49762,N_49913);
nor UO_4034 (O_4034,N_49238,N_49413);
and UO_4035 (O_4035,N_49765,N_49163);
nand UO_4036 (O_4036,N_49014,N_49383);
xor UO_4037 (O_4037,N_49223,N_49297);
xnor UO_4038 (O_4038,N_49780,N_49817);
nor UO_4039 (O_4039,N_49774,N_49353);
or UO_4040 (O_4040,N_49503,N_49161);
xor UO_4041 (O_4041,N_49360,N_49723);
or UO_4042 (O_4042,N_49613,N_49875);
nand UO_4043 (O_4043,N_49798,N_49684);
nand UO_4044 (O_4044,N_49436,N_49670);
or UO_4045 (O_4045,N_49685,N_49392);
nor UO_4046 (O_4046,N_49235,N_49287);
and UO_4047 (O_4047,N_49296,N_49700);
xor UO_4048 (O_4048,N_49127,N_49271);
nand UO_4049 (O_4049,N_49942,N_49184);
or UO_4050 (O_4050,N_49723,N_49398);
or UO_4051 (O_4051,N_49472,N_49138);
nor UO_4052 (O_4052,N_49130,N_49351);
or UO_4053 (O_4053,N_49568,N_49298);
xor UO_4054 (O_4054,N_49257,N_49988);
or UO_4055 (O_4055,N_49272,N_49054);
nor UO_4056 (O_4056,N_49675,N_49100);
xnor UO_4057 (O_4057,N_49836,N_49406);
and UO_4058 (O_4058,N_49942,N_49341);
nor UO_4059 (O_4059,N_49159,N_49238);
and UO_4060 (O_4060,N_49173,N_49602);
and UO_4061 (O_4061,N_49071,N_49469);
or UO_4062 (O_4062,N_49449,N_49977);
nor UO_4063 (O_4063,N_49452,N_49194);
nor UO_4064 (O_4064,N_49041,N_49520);
nor UO_4065 (O_4065,N_49168,N_49627);
nor UO_4066 (O_4066,N_49848,N_49874);
or UO_4067 (O_4067,N_49966,N_49650);
xor UO_4068 (O_4068,N_49784,N_49061);
nand UO_4069 (O_4069,N_49074,N_49938);
nand UO_4070 (O_4070,N_49046,N_49037);
nor UO_4071 (O_4071,N_49229,N_49103);
nor UO_4072 (O_4072,N_49851,N_49978);
xor UO_4073 (O_4073,N_49834,N_49932);
xor UO_4074 (O_4074,N_49932,N_49762);
xor UO_4075 (O_4075,N_49820,N_49718);
nor UO_4076 (O_4076,N_49514,N_49752);
or UO_4077 (O_4077,N_49273,N_49414);
xor UO_4078 (O_4078,N_49998,N_49694);
xor UO_4079 (O_4079,N_49020,N_49394);
or UO_4080 (O_4080,N_49496,N_49968);
or UO_4081 (O_4081,N_49785,N_49200);
nand UO_4082 (O_4082,N_49011,N_49710);
xor UO_4083 (O_4083,N_49471,N_49223);
and UO_4084 (O_4084,N_49472,N_49511);
xor UO_4085 (O_4085,N_49575,N_49268);
and UO_4086 (O_4086,N_49127,N_49294);
or UO_4087 (O_4087,N_49603,N_49505);
xor UO_4088 (O_4088,N_49954,N_49206);
or UO_4089 (O_4089,N_49403,N_49550);
xor UO_4090 (O_4090,N_49021,N_49709);
xor UO_4091 (O_4091,N_49596,N_49114);
nor UO_4092 (O_4092,N_49992,N_49066);
and UO_4093 (O_4093,N_49363,N_49254);
xor UO_4094 (O_4094,N_49272,N_49690);
and UO_4095 (O_4095,N_49514,N_49584);
and UO_4096 (O_4096,N_49902,N_49330);
nand UO_4097 (O_4097,N_49672,N_49993);
xor UO_4098 (O_4098,N_49143,N_49574);
nand UO_4099 (O_4099,N_49174,N_49964);
nor UO_4100 (O_4100,N_49498,N_49802);
nor UO_4101 (O_4101,N_49469,N_49857);
and UO_4102 (O_4102,N_49907,N_49507);
or UO_4103 (O_4103,N_49086,N_49576);
or UO_4104 (O_4104,N_49205,N_49192);
xnor UO_4105 (O_4105,N_49633,N_49417);
nand UO_4106 (O_4106,N_49331,N_49876);
xor UO_4107 (O_4107,N_49705,N_49085);
nor UO_4108 (O_4108,N_49965,N_49366);
and UO_4109 (O_4109,N_49462,N_49941);
xnor UO_4110 (O_4110,N_49134,N_49277);
and UO_4111 (O_4111,N_49054,N_49781);
nor UO_4112 (O_4112,N_49147,N_49014);
nand UO_4113 (O_4113,N_49653,N_49701);
nor UO_4114 (O_4114,N_49754,N_49148);
nor UO_4115 (O_4115,N_49441,N_49151);
or UO_4116 (O_4116,N_49241,N_49170);
or UO_4117 (O_4117,N_49020,N_49793);
nand UO_4118 (O_4118,N_49450,N_49792);
or UO_4119 (O_4119,N_49740,N_49585);
nor UO_4120 (O_4120,N_49120,N_49580);
xnor UO_4121 (O_4121,N_49571,N_49898);
nor UO_4122 (O_4122,N_49615,N_49296);
nor UO_4123 (O_4123,N_49948,N_49044);
or UO_4124 (O_4124,N_49229,N_49097);
or UO_4125 (O_4125,N_49638,N_49132);
and UO_4126 (O_4126,N_49192,N_49087);
and UO_4127 (O_4127,N_49610,N_49359);
and UO_4128 (O_4128,N_49413,N_49980);
xnor UO_4129 (O_4129,N_49097,N_49987);
or UO_4130 (O_4130,N_49246,N_49181);
nand UO_4131 (O_4131,N_49509,N_49391);
or UO_4132 (O_4132,N_49416,N_49113);
nand UO_4133 (O_4133,N_49884,N_49323);
nor UO_4134 (O_4134,N_49539,N_49722);
nand UO_4135 (O_4135,N_49087,N_49395);
nand UO_4136 (O_4136,N_49559,N_49680);
xnor UO_4137 (O_4137,N_49752,N_49929);
nand UO_4138 (O_4138,N_49596,N_49376);
xor UO_4139 (O_4139,N_49653,N_49282);
and UO_4140 (O_4140,N_49020,N_49056);
nor UO_4141 (O_4141,N_49458,N_49621);
and UO_4142 (O_4142,N_49229,N_49117);
nor UO_4143 (O_4143,N_49028,N_49949);
or UO_4144 (O_4144,N_49157,N_49147);
or UO_4145 (O_4145,N_49094,N_49541);
nand UO_4146 (O_4146,N_49639,N_49308);
xnor UO_4147 (O_4147,N_49118,N_49857);
and UO_4148 (O_4148,N_49610,N_49870);
nand UO_4149 (O_4149,N_49729,N_49117);
xnor UO_4150 (O_4150,N_49959,N_49988);
xor UO_4151 (O_4151,N_49652,N_49038);
or UO_4152 (O_4152,N_49856,N_49321);
nor UO_4153 (O_4153,N_49589,N_49981);
nor UO_4154 (O_4154,N_49327,N_49528);
nor UO_4155 (O_4155,N_49397,N_49149);
or UO_4156 (O_4156,N_49595,N_49679);
or UO_4157 (O_4157,N_49705,N_49661);
and UO_4158 (O_4158,N_49578,N_49215);
nor UO_4159 (O_4159,N_49363,N_49043);
xnor UO_4160 (O_4160,N_49439,N_49392);
xnor UO_4161 (O_4161,N_49435,N_49681);
nor UO_4162 (O_4162,N_49936,N_49202);
nor UO_4163 (O_4163,N_49682,N_49529);
nand UO_4164 (O_4164,N_49464,N_49875);
nand UO_4165 (O_4165,N_49516,N_49165);
or UO_4166 (O_4166,N_49556,N_49405);
nor UO_4167 (O_4167,N_49693,N_49244);
and UO_4168 (O_4168,N_49770,N_49132);
nor UO_4169 (O_4169,N_49839,N_49225);
or UO_4170 (O_4170,N_49824,N_49576);
xnor UO_4171 (O_4171,N_49904,N_49801);
xor UO_4172 (O_4172,N_49172,N_49805);
or UO_4173 (O_4173,N_49237,N_49036);
xor UO_4174 (O_4174,N_49990,N_49729);
nand UO_4175 (O_4175,N_49691,N_49510);
xnor UO_4176 (O_4176,N_49815,N_49259);
xnor UO_4177 (O_4177,N_49361,N_49705);
nand UO_4178 (O_4178,N_49156,N_49059);
nand UO_4179 (O_4179,N_49071,N_49055);
nand UO_4180 (O_4180,N_49755,N_49627);
and UO_4181 (O_4181,N_49114,N_49652);
xor UO_4182 (O_4182,N_49944,N_49479);
and UO_4183 (O_4183,N_49224,N_49289);
nor UO_4184 (O_4184,N_49099,N_49147);
nand UO_4185 (O_4185,N_49285,N_49893);
and UO_4186 (O_4186,N_49041,N_49088);
nor UO_4187 (O_4187,N_49885,N_49223);
xnor UO_4188 (O_4188,N_49237,N_49002);
xor UO_4189 (O_4189,N_49042,N_49132);
xnor UO_4190 (O_4190,N_49848,N_49423);
nor UO_4191 (O_4191,N_49641,N_49402);
nor UO_4192 (O_4192,N_49976,N_49677);
and UO_4193 (O_4193,N_49197,N_49135);
nor UO_4194 (O_4194,N_49249,N_49587);
and UO_4195 (O_4195,N_49384,N_49593);
and UO_4196 (O_4196,N_49222,N_49168);
or UO_4197 (O_4197,N_49565,N_49776);
nand UO_4198 (O_4198,N_49653,N_49545);
nor UO_4199 (O_4199,N_49916,N_49882);
and UO_4200 (O_4200,N_49855,N_49357);
and UO_4201 (O_4201,N_49213,N_49842);
and UO_4202 (O_4202,N_49813,N_49902);
and UO_4203 (O_4203,N_49459,N_49282);
or UO_4204 (O_4204,N_49464,N_49085);
xor UO_4205 (O_4205,N_49656,N_49468);
and UO_4206 (O_4206,N_49333,N_49096);
and UO_4207 (O_4207,N_49694,N_49908);
and UO_4208 (O_4208,N_49855,N_49271);
xnor UO_4209 (O_4209,N_49259,N_49329);
or UO_4210 (O_4210,N_49125,N_49306);
and UO_4211 (O_4211,N_49891,N_49558);
nor UO_4212 (O_4212,N_49770,N_49045);
or UO_4213 (O_4213,N_49123,N_49597);
nand UO_4214 (O_4214,N_49367,N_49735);
xnor UO_4215 (O_4215,N_49349,N_49867);
nor UO_4216 (O_4216,N_49673,N_49086);
nand UO_4217 (O_4217,N_49741,N_49748);
xor UO_4218 (O_4218,N_49546,N_49422);
nand UO_4219 (O_4219,N_49670,N_49550);
and UO_4220 (O_4220,N_49852,N_49441);
and UO_4221 (O_4221,N_49357,N_49622);
nor UO_4222 (O_4222,N_49147,N_49178);
nor UO_4223 (O_4223,N_49528,N_49271);
nand UO_4224 (O_4224,N_49792,N_49279);
and UO_4225 (O_4225,N_49441,N_49742);
nand UO_4226 (O_4226,N_49310,N_49961);
and UO_4227 (O_4227,N_49729,N_49820);
or UO_4228 (O_4228,N_49699,N_49424);
or UO_4229 (O_4229,N_49762,N_49276);
and UO_4230 (O_4230,N_49292,N_49964);
xor UO_4231 (O_4231,N_49389,N_49953);
nand UO_4232 (O_4232,N_49602,N_49791);
xor UO_4233 (O_4233,N_49221,N_49890);
or UO_4234 (O_4234,N_49152,N_49372);
or UO_4235 (O_4235,N_49567,N_49436);
and UO_4236 (O_4236,N_49723,N_49432);
nor UO_4237 (O_4237,N_49686,N_49455);
and UO_4238 (O_4238,N_49168,N_49873);
nand UO_4239 (O_4239,N_49837,N_49439);
nor UO_4240 (O_4240,N_49044,N_49257);
xnor UO_4241 (O_4241,N_49482,N_49424);
nand UO_4242 (O_4242,N_49117,N_49147);
nor UO_4243 (O_4243,N_49980,N_49539);
or UO_4244 (O_4244,N_49974,N_49449);
and UO_4245 (O_4245,N_49484,N_49343);
nand UO_4246 (O_4246,N_49928,N_49685);
or UO_4247 (O_4247,N_49821,N_49810);
nor UO_4248 (O_4248,N_49482,N_49541);
and UO_4249 (O_4249,N_49071,N_49174);
xor UO_4250 (O_4250,N_49118,N_49564);
or UO_4251 (O_4251,N_49950,N_49295);
nor UO_4252 (O_4252,N_49563,N_49750);
xor UO_4253 (O_4253,N_49019,N_49805);
and UO_4254 (O_4254,N_49071,N_49795);
and UO_4255 (O_4255,N_49354,N_49232);
nand UO_4256 (O_4256,N_49673,N_49396);
nand UO_4257 (O_4257,N_49800,N_49921);
xnor UO_4258 (O_4258,N_49326,N_49403);
xor UO_4259 (O_4259,N_49384,N_49675);
and UO_4260 (O_4260,N_49511,N_49663);
xnor UO_4261 (O_4261,N_49309,N_49115);
and UO_4262 (O_4262,N_49184,N_49125);
nor UO_4263 (O_4263,N_49759,N_49696);
and UO_4264 (O_4264,N_49004,N_49831);
and UO_4265 (O_4265,N_49104,N_49220);
and UO_4266 (O_4266,N_49603,N_49548);
and UO_4267 (O_4267,N_49590,N_49192);
nor UO_4268 (O_4268,N_49599,N_49171);
nand UO_4269 (O_4269,N_49666,N_49837);
or UO_4270 (O_4270,N_49877,N_49767);
and UO_4271 (O_4271,N_49738,N_49059);
and UO_4272 (O_4272,N_49223,N_49157);
or UO_4273 (O_4273,N_49306,N_49834);
nor UO_4274 (O_4274,N_49083,N_49766);
or UO_4275 (O_4275,N_49471,N_49286);
or UO_4276 (O_4276,N_49469,N_49428);
xnor UO_4277 (O_4277,N_49797,N_49535);
nor UO_4278 (O_4278,N_49148,N_49163);
nor UO_4279 (O_4279,N_49336,N_49613);
xnor UO_4280 (O_4280,N_49223,N_49845);
xnor UO_4281 (O_4281,N_49229,N_49817);
nand UO_4282 (O_4282,N_49204,N_49858);
nand UO_4283 (O_4283,N_49030,N_49161);
and UO_4284 (O_4284,N_49331,N_49027);
nand UO_4285 (O_4285,N_49943,N_49964);
nand UO_4286 (O_4286,N_49822,N_49843);
nor UO_4287 (O_4287,N_49587,N_49562);
xor UO_4288 (O_4288,N_49781,N_49452);
or UO_4289 (O_4289,N_49342,N_49170);
nor UO_4290 (O_4290,N_49888,N_49852);
nand UO_4291 (O_4291,N_49372,N_49545);
xor UO_4292 (O_4292,N_49477,N_49243);
and UO_4293 (O_4293,N_49580,N_49170);
nand UO_4294 (O_4294,N_49657,N_49184);
and UO_4295 (O_4295,N_49513,N_49038);
and UO_4296 (O_4296,N_49040,N_49920);
or UO_4297 (O_4297,N_49784,N_49526);
or UO_4298 (O_4298,N_49884,N_49343);
nand UO_4299 (O_4299,N_49067,N_49850);
and UO_4300 (O_4300,N_49419,N_49146);
nand UO_4301 (O_4301,N_49075,N_49553);
xor UO_4302 (O_4302,N_49085,N_49417);
or UO_4303 (O_4303,N_49848,N_49693);
nand UO_4304 (O_4304,N_49865,N_49335);
or UO_4305 (O_4305,N_49587,N_49627);
nor UO_4306 (O_4306,N_49411,N_49330);
and UO_4307 (O_4307,N_49413,N_49313);
nor UO_4308 (O_4308,N_49958,N_49957);
and UO_4309 (O_4309,N_49343,N_49406);
or UO_4310 (O_4310,N_49176,N_49440);
xnor UO_4311 (O_4311,N_49641,N_49320);
nor UO_4312 (O_4312,N_49139,N_49779);
xor UO_4313 (O_4313,N_49591,N_49184);
and UO_4314 (O_4314,N_49463,N_49490);
nor UO_4315 (O_4315,N_49058,N_49623);
or UO_4316 (O_4316,N_49571,N_49454);
xor UO_4317 (O_4317,N_49053,N_49146);
nand UO_4318 (O_4318,N_49810,N_49334);
nor UO_4319 (O_4319,N_49268,N_49945);
or UO_4320 (O_4320,N_49251,N_49827);
and UO_4321 (O_4321,N_49131,N_49070);
and UO_4322 (O_4322,N_49508,N_49075);
nor UO_4323 (O_4323,N_49058,N_49225);
or UO_4324 (O_4324,N_49878,N_49687);
or UO_4325 (O_4325,N_49930,N_49755);
nor UO_4326 (O_4326,N_49738,N_49973);
and UO_4327 (O_4327,N_49877,N_49594);
nor UO_4328 (O_4328,N_49714,N_49870);
nor UO_4329 (O_4329,N_49649,N_49779);
nand UO_4330 (O_4330,N_49739,N_49026);
nand UO_4331 (O_4331,N_49173,N_49814);
nand UO_4332 (O_4332,N_49469,N_49172);
xor UO_4333 (O_4333,N_49621,N_49623);
and UO_4334 (O_4334,N_49203,N_49631);
and UO_4335 (O_4335,N_49739,N_49916);
or UO_4336 (O_4336,N_49239,N_49442);
xor UO_4337 (O_4337,N_49761,N_49741);
and UO_4338 (O_4338,N_49843,N_49749);
xnor UO_4339 (O_4339,N_49722,N_49728);
and UO_4340 (O_4340,N_49777,N_49802);
xor UO_4341 (O_4341,N_49299,N_49463);
nand UO_4342 (O_4342,N_49173,N_49302);
xor UO_4343 (O_4343,N_49712,N_49284);
nand UO_4344 (O_4344,N_49579,N_49308);
nand UO_4345 (O_4345,N_49148,N_49923);
and UO_4346 (O_4346,N_49074,N_49750);
or UO_4347 (O_4347,N_49533,N_49525);
nand UO_4348 (O_4348,N_49320,N_49950);
nor UO_4349 (O_4349,N_49802,N_49698);
or UO_4350 (O_4350,N_49174,N_49528);
nor UO_4351 (O_4351,N_49274,N_49774);
and UO_4352 (O_4352,N_49851,N_49303);
xor UO_4353 (O_4353,N_49751,N_49833);
nand UO_4354 (O_4354,N_49229,N_49483);
nand UO_4355 (O_4355,N_49761,N_49717);
and UO_4356 (O_4356,N_49241,N_49614);
nor UO_4357 (O_4357,N_49470,N_49952);
and UO_4358 (O_4358,N_49161,N_49931);
and UO_4359 (O_4359,N_49341,N_49739);
nand UO_4360 (O_4360,N_49861,N_49396);
nor UO_4361 (O_4361,N_49683,N_49058);
and UO_4362 (O_4362,N_49229,N_49957);
nand UO_4363 (O_4363,N_49127,N_49781);
and UO_4364 (O_4364,N_49895,N_49284);
nand UO_4365 (O_4365,N_49146,N_49035);
nor UO_4366 (O_4366,N_49674,N_49584);
xor UO_4367 (O_4367,N_49179,N_49557);
xor UO_4368 (O_4368,N_49201,N_49633);
nor UO_4369 (O_4369,N_49771,N_49233);
nand UO_4370 (O_4370,N_49051,N_49434);
nand UO_4371 (O_4371,N_49197,N_49382);
or UO_4372 (O_4372,N_49555,N_49072);
or UO_4373 (O_4373,N_49471,N_49450);
or UO_4374 (O_4374,N_49653,N_49923);
nor UO_4375 (O_4375,N_49965,N_49238);
or UO_4376 (O_4376,N_49264,N_49735);
xor UO_4377 (O_4377,N_49197,N_49075);
nor UO_4378 (O_4378,N_49747,N_49733);
nand UO_4379 (O_4379,N_49078,N_49577);
nor UO_4380 (O_4380,N_49385,N_49859);
or UO_4381 (O_4381,N_49505,N_49793);
xnor UO_4382 (O_4382,N_49835,N_49219);
xor UO_4383 (O_4383,N_49431,N_49163);
nor UO_4384 (O_4384,N_49985,N_49802);
xnor UO_4385 (O_4385,N_49483,N_49052);
xnor UO_4386 (O_4386,N_49512,N_49524);
nand UO_4387 (O_4387,N_49995,N_49272);
nand UO_4388 (O_4388,N_49238,N_49697);
nand UO_4389 (O_4389,N_49403,N_49128);
and UO_4390 (O_4390,N_49050,N_49571);
and UO_4391 (O_4391,N_49142,N_49033);
nor UO_4392 (O_4392,N_49124,N_49189);
or UO_4393 (O_4393,N_49030,N_49874);
and UO_4394 (O_4394,N_49067,N_49191);
or UO_4395 (O_4395,N_49975,N_49345);
nand UO_4396 (O_4396,N_49311,N_49596);
and UO_4397 (O_4397,N_49999,N_49872);
or UO_4398 (O_4398,N_49356,N_49094);
and UO_4399 (O_4399,N_49829,N_49428);
nor UO_4400 (O_4400,N_49055,N_49296);
nor UO_4401 (O_4401,N_49152,N_49326);
and UO_4402 (O_4402,N_49255,N_49581);
nand UO_4403 (O_4403,N_49026,N_49347);
or UO_4404 (O_4404,N_49449,N_49338);
and UO_4405 (O_4405,N_49884,N_49761);
xnor UO_4406 (O_4406,N_49184,N_49220);
and UO_4407 (O_4407,N_49550,N_49991);
or UO_4408 (O_4408,N_49741,N_49927);
or UO_4409 (O_4409,N_49194,N_49563);
xor UO_4410 (O_4410,N_49947,N_49015);
and UO_4411 (O_4411,N_49367,N_49620);
nand UO_4412 (O_4412,N_49486,N_49366);
xor UO_4413 (O_4413,N_49547,N_49772);
nand UO_4414 (O_4414,N_49844,N_49268);
nand UO_4415 (O_4415,N_49916,N_49098);
nand UO_4416 (O_4416,N_49671,N_49107);
xnor UO_4417 (O_4417,N_49741,N_49150);
xor UO_4418 (O_4418,N_49571,N_49515);
nand UO_4419 (O_4419,N_49305,N_49212);
nor UO_4420 (O_4420,N_49535,N_49455);
or UO_4421 (O_4421,N_49421,N_49372);
and UO_4422 (O_4422,N_49768,N_49074);
or UO_4423 (O_4423,N_49201,N_49493);
nor UO_4424 (O_4424,N_49587,N_49772);
xor UO_4425 (O_4425,N_49597,N_49479);
or UO_4426 (O_4426,N_49788,N_49235);
xor UO_4427 (O_4427,N_49949,N_49578);
or UO_4428 (O_4428,N_49191,N_49617);
nand UO_4429 (O_4429,N_49214,N_49478);
xor UO_4430 (O_4430,N_49429,N_49407);
xnor UO_4431 (O_4431,N_49431,N_49148);
xnor UO_4432 (O_4432,N_49473,N_49748);
xnor UO_4433 (O_4433,N_49130,N_49951);
or UO_4434 (O_4434,N_49812,N_49821);
nor UO_4435 (O_4435,N_49618,N_49393);
xnor UO_4436 (O_4436,N_49700,N_49094);
or UO_4437 (O_4437,N_49911,N_49317);
xnor UO_4438 (O_4438,N_49131,N_49080);
xnor UO_4439 (O_4439,N_49345,N_49035);
nor UO_4440 (O_4440,N_49668,N_49622);
nor UO_4441 (O_4441,N_49057,N_49132);
xor UO_4442 (O_4442,N_49926,N_49629);
or UO_4443 (O_4443,N_49303,N_49153);
or UO_4444 (O_4444,N_49096,N_49843);
nand UO_4445 (O_4445,N_49057,N_49855);
or UO_4446 (O_4446,N_49986,N_49425);
xor UO_4447 (O_4447,N_49328,N_49860);
or UO_4448 (O_4448,N_49321,N_49400);
xnor UO_4449 (O_4449,N_49479,N_49860);
nand UO_4450 (O_4450,N_49716,N_49247);
or UO_4451 (O_4451,N_49501,N_49826);
nand UO_4452 (O_4452,N_49852,N_49480);
nor UO_4453 (O_4453,N_49768,N_49306);
and UO_4454 (O_4454,N_49995,N_49933);
and UO_4455 (O_4455,N_49119,N_49636);
nand UO_4456 (O_4456,N_49029,N_49155);
nor UO_4457 (O_4457,N_49858,N_49075);
nand UO_4458 (O_4458,N_49126,N_49050);
or UO_4459 (O_4459,N_49353,N_49140);
and UO_4460 (O_4460,N_49124,N_49977);
or UO_4461 (O_4461,N_49861,N_49171);
nor UO_4462 (O_4462,N_49777,N_49898);
and UO_4463 (O_4463,N_49843,N_49541);
nor UO_4464 (O_4464,N_49540,N_49020);
xnor UO_4465 (O_4465,N_49228,N_49993);
nor UO_4466 (O_4466,N_49517,N_49019);
xnor UO_4467 (O_4467,N_49031,N_49819);
nor UO_4468 (O_4468,N_49647,N_49319);
or UO_4469 (O_4469,N_49682,N_49769);
and UO_4470 (O_4470,N_49096,N_49047);
and UO_4471 (O_4471,N_49176,N_49354);
xnor UO_4472 (O_4472,N_49071,N_49689);
or UO_4473 (O_4473,N_49608,N_49034);
or UO_4474 (O_4474,N_49983,N_49985);
nand UO_4475 (O_4475,N_49819,N_49702);
nor UO_4476 (O_4476,N_49320,N_49763);
xor UO_4477 (O_4477,N_49633,N_49257);
and UO_4478 (O_4478,N_49191,N_49815);
or UO_4479 (O_4479,N_49983,N_49448);
nor UO_4480 (O_4480,N_49526,N_49690);
nor UO_4481 (O_4481,N_49367,N_49129);
and UO_4482 (O_4482,N_49156,N_49107);
nor UO_4483 (O_4483,N_49655,N_49517);
nor UO_4484 (O_4484,N_49257,N_49254);
nor UO_4485 (O_4485,N_49614,N_49603);
nand UO_4486 (O_4486,N_49089,N_49726);
or UO_4487 (O_4487,N_49039,N_49869);
nor UO_4488 (O_4488,N_49048,N_49684);
xor UO_4489 (O_4489,N_49249,N_49434);
and UO_4490 (O_4490,N_49148,N_49953);
nand UO_4491 (O_4491,N_49789,N_49579);
or UO_4492 (O_4492,N_49120,N_49852);
nand UO_4493 (O_4493,N_49452,N_49527);
and UO_4494 (O_4494,N_49828,N_49154);
xor UO_4495 (O_4495,N_49513,N_49459);
and UO_4496 (O_4496,N_49024,N_49675);
and UO_4497 (O_4497,N_49749,N_49829);
nor UO_4498 (O_4498,N_49055,N_49142);
and UO_4499 (O_4499,N_49717,N_49697);
nand UO_4500 (O_4500,N_49189,N_49733);
or UO_4501 (O_4501,N_49459,N_49872);
nor UO_4502 (O_4502,N_49875,N_49501);
nand UO_4503 (O_4503,N_49450,N_49361);
and UO_4504 (O_4504,N_49145,N_49639);
xnor UO_4505 (O_4505,N_49999,N_49342);
nand UO_4506 (O_4506,N_49150,N_49656);
nand UO_4507 (O_4507,N_49846,N_49672);
or UO_4508 (O_4508,N_49861,N_49990);
nor UO_4509 (O_4509,N_49114,N_49535);
and UO_4510 (O_4510,N_49082,N_49419);
and UO_4511 (O_4511,N_49519,N_49087);
nand UO_4512 (O_4512,N_49982,N_49886);
and UO_4513 (O_4513,N_49962,N_49545);
nand UO_4514 (O_4514,N_49785,N_49527);
or UO_4515 (O_4515,N_49814,N_49122);
nand UO_4516 (O_4516,N_49783,N_49182);
nand UO_4517 (O_4517,N_49448,N_49530);
nand UO_4518 (O_4518,N_49566,N_49992);
nor UO_4519 (O_4519,N_49849,N_49537);
and UO_4520 (O_4520,N_49327,N_49471);
nand UO_4521 (O_4521,N_49163,N_49967);
nand UO_4522 (O_4522,N_49265,N_49821);
xnor UO_4523 (O_4523,N_49432,N_49297);
xnor UO_4524 (O_4524,N_49444,N_49108);
nand UO_4525 (O_4525,N_49276,N_49325);
or UO_4526 (O_4526,N_49096,N_49390);
or UO_4527 (O_4527,N_49906,N_49523);
or UO_4528 (O_4528,N_49101,N_49321);
and UO_4529 (O_4529,N_49352,N_49313);
or UO_4530 (O_4530,N_49228,N_49675);
or UO_4531 (O_4531,N_49829,N_49971);
nand UO_4532 (O_4532,N_49186,N_49225);
nor UO_4533 (O_4533,N_49315,N_49421);
or UO_4534 (O_4534,N_49179,N_49837);
or UO_4535 (O_4535,N_49563,N_49466);
nand UO_4536 (O_4536,N_49932,N_49590);
nand UO_4537 (O_4537,N_49842,N_49665);
nor UO_4538 (O_4538,N_49083,N_49941);
nor UO_4539 (O_4539,N_49987,N_49082);
nand UO_4540 (O_4540,N_49083,N_49661);
or UO_4541 (O_4541,N_49777,N_49497);
xor UO_4542 (O_4542,N_49349,N_49497);
nor UO_4543 (O_4543,N_49637,N_49194);
xor UO_4544 (O_4544,N_49170,N_49538);
xnor UO_4545 (O_4545,N_49448,N_49516);
nor UO_4546 (O_4546,N_49136,N_49512);
xnor UO_4547 (O_4547,N_49948,N_49962);
or UO_4548 (O_4548,N_49001,N_49636);
and UO_4549 (O_4549,N_49366,N_49420);
or UO_4550 (O_4550,N_49488,N_49581);
or UO_4551 (O_4551,N_49898,N_49653);
xnor UO_4552 (O_4552,N_49385,N_49426);
nor UO_4553 (O_4553,N_49055,N_49380);
xor UO_4554 (O_4554,N_49963,N_49111);
xor UO_4555 (O_4555,N_49153,N_49217);
and UO_4556 (O_4556,N_49214,N_49589);
or UO_4557 (O_4557,N_49969,N_49582);
nor UO_4558 (O_4558,N_49078,N_49703);
nand UO_4559 (O_4559,N_49361,N_49706);
xor UO_4560 (O_4560,N_49615,N_49848);
nor UO_4561 (O_4561,N_49581,N_49022);
or UO_4562 (O_4562,N_49792,N_49043);
xor UO_4563 (O_4563,N_49481,N_49956);
or UO_4564 (O_4564,N_49638,N_49936);
or UO_4565 (O_4565,N_49031,N_49744);
xor UO_4566 (O_4566,N_49589,N_49072);
or UO_4567 (O_4567,N_49777,N_49465);
or UO_4568 (O_4568,N_49246,N_49595);
nor UO_4569 (O_4569,N_49056,N_49602);
nor UO_4570 (O_4570,N_49565,N_49619);
nor UO_4571 (O_4571,N_49327,N_49397);
xnor UO_4572 (O_4572,N_49913,N_49549);
or UO_4573 (O_4573,N_49899,N_49414);
and UO_4574 (O_4574,N_49317,N_49618);
nor UO_4575 (O_4575,N_49506,N_49839);
nand UO_4576 (O_4576,N_49661,N_49358);
nand UO_4577 (O_4577,N_49740,N_49788);
or UO_4578 (O_4578,N_49009,N_49605);
xnor UO_4579 (O_4579,N_49922,N_49607);
xnor UO_4580 (O_4580,N_49444,N_49981);
nand UO_4581 (O_4581,N_49658,N_49468);
xor UO_4582 (O_4582,N_49237,N_49887);
or UO_4583 (O_4583,N_49056,N_49846);
nor UO_4584 (O_4584,N_49948,N_49433);
nor UO_4585 (O_4585,N_49409,N_49951);
or UO_4586 (O_4586,N_49374,N_49266);
nor UO_4587 (O_4587,N_49329,N_49384);
xnor UO_4588 (O_4588,N_49360,N_49102);
or UO_4589 (O_4589,N_49548,N_49577);
xnor UO_4590 (O_4590,N_49904,N_49083);
and UO_4591 (O_4591,N_49050,N_49950);
and UO_4592 (O_4592,N_49797,N_49468);
xor UO_4593 (O_4593,N_49049,N_49988);
xor UO_4594 (O_4594,N_49745,N_49907);
xnor UO_4595 (O_4595,N_49154,N_49970);
or UO_4596 (O_4596,N_49249,N_49103);
and UO_4597 (O_4597,N_49232,N_49665);
nor UO_4598 (O_4598,N_49022,N_49188);
and UO_4599 (O_4599,N_49869,N_49029);
and UO_4600 (O_4600,N_49896,N_49060);
nor UO_4601 (O_4601,N_49146,N_49831);
xor UO_4602 (O_4602,N_49248,N_49445);
or UO_4603 (O_4603,N_49051,N_49406);
nor UO_4604 (O_4604,N_49860,N_49486);
and UO_4605 (O_4605,N_49326,N_49622);
nor UO_4606 (O_4606,N_49682,N_49814);
or UO_4607 (O_4607,N_49968,N_49105);
and UO_4608 (O_4608,N_49638,N_49521);
xnor UO_4609 (O_4609,N_49030,N_49933);
nor UO_4610 (O_4610,N_49150,N_49234);
nand UO_4611 (O_4611,N_49489,N_49908);
nor UO_4612 (O_4612,N_49580,N_49117);
xnor UO_4613 (O_4613,N_49277,N_49990);
xor UO_4614 (O_4614,N_49247,N_49000);
and UO_4615 (O_4615,N_49503,N_49130);
and UO_4616 (O_4616,N_49705,N_49301);
xnor UO_4617 (O_4617,N_49074,N_49691);
nor UO_4618 (O_4618,N_49478,N_49332);
or UO_4619 (O_4619,N_49624,N_49611);
nor UO_4620 (O_4620,N_49028,N_49340);
nor UO_4621 (O_4621,N_49482,N_49528);
or UO_4622 (O_4622,N_49447,N_49275);
nor UO_4623 (O_4623,N_49843,N_49369);
nor UO_4624 (O_4624,N_49652,N_49763);
nor UO_4625 (O_4625,N_49681,N_49208);
and UO_4626 (O_4626,N_49916,N_49738);
or UO_4627 (O_4627,N_49060,N_49037);
xnor UO_4628 (O_4628,N_49883,N_49391);
xnor UO_4629 (O_4629,N_49799,N_49820);
xor UO_4630 (O_4630,N_49558,N_49128);
and UO_4631 (O_4631,N_49633,N_49349);
or UO_4632 (O_4632,N_49416,N_49993);
and UO_4633 (O_4633,N_49034,N_49857);
and UO_4634 (O_4634,N_49055,N_49672);
or UO_4635 (O_4635,N_49687,N_49428);
or UO_4636 (O_4636,N_49991,N_49313);
nor UO_4637 (O_4637,N_49145,N_49282);
nand UO_4638 (O_4638,N_49155,N_49645);
nor UO_4639 (O_4639,N_49931,N_49232);
nand UO_4640 (O_4640,N_49693,N_49490);
nor UO_4641 (O_4641,N_49984,N_49411);
or UO_4642 (O_4642,N_49504,N_49613);
and UO_4643 (O_4643,N_49104,N_49779);
or UO_4644 (O_4644,N_49957,N_49681);
and UO_4645 (O_4645,N_49719,N_49368);
or UO_4646 (O_4646,N_49715,N_49095);
nand UO_4647 (O_4647,N_49177,N_49240);
nor UO_4648 (O_4648,N_49103,N_49624);
and UO_4649 (O_4649,N_49256,N_49937);
and UO_4650 (O_4650,N_49418,N_49736);
or UO_4651 (O_4651,N_49899,N_49099);
and UO_4652 (O_4652,N_49418,N_49152);
xor UO_4653 (O_4653,N_49040,N_49383);
and UO_4654 (O_4654,N_49394,N_49995);
or UO_4655 (O_4655,N_49094,N_49126);
nor UO_4656 (O_4656,N_49107,N_49905);
and UO_4657 (O_4657,N_49071,N_49431);
and UO_4658 (O_4658,N_49218,N_49382);
nor UO_4659 (O_4659,N_49823,N_49333);
or UO_4660 (O_4660,N_49379,N_49341);
and UO_4661 (O_4661,N_49670,N_49459);
and UO_4662 (O_4662,N_49991,N_49626);
nor UO_4663 (O_4663,N_49221,N_49513);
or UO_4664 (O_4664,N_49872,N_49750);
nor UO_4665 (O_4665,N_49760,N_49532);
xor UO_4666 (O_4666,N_49553,N_49286);
nand UO_4667 (O_4667,N_49469,N_49230);
nor UO_4668 (O_4668,N_49907,N_49927);
nor UO_4669 (O_4669,N_49066,N_49540);
or UO_4670 (O_4670,N_49844,N_49180);
nand UO_4671 (O_4671,N_49577,N_49115);
nor UO_4672 (O_4672,N_49735,N_49216);
nor UO_4673 (O_4673,N_49074,N_49265);
and UO_4674 (O_4674,N_49559,N_49240);
nor UO_4675 (O_4675,N_49089,N_49163);
nand UO_4676 (O_4676,N_49402,N_49658);
nand UO_4677 (O_4677,N_49676,N_49612);
nor UO_4678 (O_4678,N_49523,N_49429);
or UO_4679 (O_4679,N_49487,N_49603);
and UO_4680 (O_4680,N_49921,N_49430);
and UO_4681 (O_4681,N_49055,N_49747);
nand UO_4682 (O_4682,N_49276,N_49769);
nand UO_4683 (O_4683,N_49999,N_49072);
nand UO_4684 (O_4684,N_49026,N_49835);
or UO_4685 (O_4685,N_49984,N_49789);
nor UO_4686 (O_4686,N_49822,N_49452);
nor UO_4687 (O_4687,N_49883,N_49084);
xor UO_4688 (O_4688,N_49961,N_49018);
xor UO_4689 (O_4689,N_49228,N_49516);
nand UO_4690 (O_4690,N_49246,N_49514);
xnor UO_4691 (O_4691,N_49617,N_49471);
nor UO_4692 (O_4692,N_49370,N_49462);
nor UO_4693 (O_4693,N_49244,N_49864);
or UO_4694 (O_4694,N_49043,N_49196);
nor UO_4695 (O_4695,N_49521,N_49477);
xor UO_4696 (O_4696,N_49725,N_49756);
nor UO_4697 (O_4697,N_49048,N_49166);
xnor UO_4698 (O_4698,N_49522,N_49239);
nor UO_4699 (O_4699,N_49489,N_49631);
xor UO_4700 (O_4700,N_49925,N_49981);
xnor UO_4701 (O_4701,N_49626,N_49518);
xnor UO_4702 (O_4702,N_49869,N_49438);
nand UO_4703 (O_4703,N_49206,N_49005);
xnor UO_4704 (O_4704,N_49324,N_49696);
and UO_4705 (O_4705,N_49928,N_49814);
and UO_4706 (O_4706,N_49931,N_49969);
or UO_4707 (O_4707,N_49232,N_49199);
or UO_4708 (O_4708,N_49112,N_49051);
nand UO_4709 (O_4709,N_49359,N_49426);
and UO_4710 (O_4710,N_49017,N_49934);
and UO_4711 (O_4711,N_49257,N_49884);
and UO_4712 (O_4712,N_49438,N_49256);
nor UO_4713 (O_4713,N_49316,N_49660);
nor UO_4714 (O_4714,N_49248,N_49754);
nor UO_4715 (O_4715,N_49053,N_49813);
nor UO_4716 (O_4716,N_49726,N_49422);
and UO_4717 (O_4717,N_49139,N_49897);
nand UO_4718 (O_4718,N_49216,N_49267);
xnor UO_4719 (O_4719,N_49037,N_49313);
xor UO_4720 (O_4720,N_49298,N_49190);
and UO_4721 (O_4721,N_49656,N_49248);
and UO_4722 (O_4722,N_49918,N_49003);
xnor UO_4723 (O_4723,N_49384,N_49342);
and UO_4724 (O_4724,N_49796,N_49898);
nor UO_4725 (O_4725,N_49961,N_49221);
and UO_4726 (O_4726,N_49092,N_49659);
and UO_4727 (O_4727,N_49003,N_49019);
nor UO_4728 (O_4728,N_49409,N_49037);
and UO_4729 (O_4729,N_49402,N_49557);
nor UO_4730 (O_4730,N_49659,N_49930);
nor UO_4731 (O_4731,N_49639,N_49420);
and UO_4732 (O_4732,N_49162,N_49172);
nand UO_4733 (O_4733,N_49640,N_49652);
nor UO_4734 (O_4734,N_49744,N_49551);
and UO_4735 (O_4735,N_49924,N_49123);
nand UO_4736 (O_4736,N_49241,N_49247);
and UO_4737 (O_4737,N_49825,N_49962);
xor UO_4738 (O_4738,N_49949,N_49014);
nor UO_4739 (O_4739,N_49892,N_49593);
and UO_4740 (O_4740,N_49936,N_49952);
nand UO_4741 (O_4741,N_49094,N_49527);
and UO_4742 (O_4742,N_49724,N_49637);
and UO_4743 (O_4743,N_49884,N_49776);
and UO_4744 (O_4744,N_49678,N_49336);
nand UO_4745 (O_4745,N_49172,N_49267);
nand UO_4746 (O_4746,N_49344,N_49608);
and UO_4747 (O_4747,N_49060,N_49972);
nor UO_4748 (O_4748,N_49623,N_49859);
or UO_4749 (O_4749,N_49747,N_49107);
nor UO_4750 (O_4750,N_49867,N_49834);
xor UO_4751 (O_4751,N_49138,N_49019);
nor UO_4752 (O_4752,N_49010,N_49243);
nand UO_4753 (O_4753,N_49608,N_49633);
nor UO_4754 (O_4754,N_49082,N_49639);
nand UO_4755 (O_4755,N_49441,N_49262);
nand UO_4756 (O_4756,N_49509,N_49094);
xnor UO_4757 (O_4757,N_49962,N_49790);
nand UO_4758 (O_4758,N_49998,N_49156);
nor UO_4759 (O_4759,N_49839,N_49150);
nand UO_4760 (O_4760,N_49795,N_49285);
nor UO_4761 (O_4761,N_49520,N_49234);
nand UO_4762 (O_4762,N_49667,N_49195);
xor UO_4763 (O_4763,N_49427,N_49037);
and UO_4764 (O_4764,N_49563,N_49695);
nor UO_4765 (O_4765,N_49366,N_49287);
xnor UO_4766 (O_4766,N_49245,N_49604);
or UO_4767 (O_4767,N_49229,N_49946);
nand UO_4768 (O_4768,N_49273,N_49497);
nor UO_4769 (O_4769,N_49803,N_49212);
nor UO_4770 (O_4770,N_49707,N_49108);
and UO_4771 (O_4771,N_49813,N_49499);
xnor UO_4772 (O_4772,N_49428,N_49576);
or UO_4773 (O_4773,N_49167,N_49007);
and UO_4774 (O_4774,N_49135,N_49766);
nor UO_4775 (O_4775,N_49306,N_49133);
nand UO_4776 (O_4776,N_49931,N_49506);
or UO_4777 (O_4777,N_49023,N_49463);
nand UO_4778 (O_4778,N_49777,N_49711);
and UO_4779 (O_4779,N_49973,N_49960);
xnor UO_4780 (O_4780,N_49682,N_49545);
or UO_4781 (O_4781,N_49659,N_49837);
xor UO_4782 (O_4782,N_49638,N_49332);
and UO_4783 (O_4783,N_49238,N_49676);
nor UO_4784 (O_4784,N_49054,N_49006);
nor UO_4785 (O_4785,N_49169,N_49350);
xor UO_4786 (O_4786,N_49004,N_49720);
nor UO_4787 (O_4787,N_49759,N_49170);
and UO_4788 (O_4788,N_49179,N_49411);
and UO_4789 (O_4789,N_49827,N_49820);
xnor UO_4790 (O_4790,N_49693,N_49328);
xor UO_4791 (O_4791,N_49008,N_49699);
xor UO_4792 (O_4792,N_49826,N_49567);
nor UO_4793 (O_4793,N_49328,N_49563);
nand UO_4794 (O_4794,N_49865,N_49411);
nand UO_4795 (O_4795,N_49518,N_49404);
or UO_4796 (O_4796,N_49165,N_49644);
and UO_4797 (O_4797,N_49622,N_49338);
nand UO_4798 (O_4798,N_49014,N_49248);
or UO_4799 (O_4799,N_49270,N_49960);
nor UO_4800 (O_4800,N_49165,N_49778);
and UO_4801 (O_4801,N_49427,N_49800);
nor UO_4802 (O_4802,N_49565,N_49762);
nand UO_4803 (O_4803,N_49482,N_49960);
nor UO_4804 (O_4804,N_49279,N_49953);
nor UO_4805 (O_4805,N_49447,N_49955);
nor UO_4806 (O_4806,N_49611,N_49464);
nor UO_4807 (O_4807,N_49281,N_49065);
nand UO_4808 (O_4808,N_49284,N_49401);
xor UO_4809 (O_4809,N_49945,N_49397);
or UO_4810 (O_4810,N_49197,N_49704);
and UO_4811 (O_4811,N_49387,N_49254);
or UO_4812 (O_4812,N_49048,N_49756);
nor UO_4813 (O_4813,N_49579,N_49235);
or UO_4814 (O_4814,N_49239,N_49823);
or UO_4815 (O_4815,N_49920,N_49263);
or UO_4816 (O_4816,N_49339,N_49854);
nor UO_4817 (O_4817,N_49179,N_49861);
and UO_4818 (O_4818,N_49670,N_49547);
nand UO_4819 (O_4819,N_49450,N_49342);
xor UO_4820 (O_4820,N_49799,N_49577);
or UO_4821 (O_4821,N_49327,N_49734);
or UO_4822 (O_4822,N_49001,N_49353);
nand UO_4823 (O_4823,N_49758,N_49359);
and UO_4824 (O_4824,N_49504,N_49948);
xnor UO_4825 (O_4825,N_49940,N_49608);
nand UO_4826 (O_4826,N_49210,N_49810);
nor UO_4827 (O_4827,N_49284,N_49085);
nand UO_4828 (O_4828,N_49205,N_49319);
or UO_4829 (O_4829,N_49080,N_49270);
or UO_4830 (O_4830,N_49170,N_49679);
nor UO_4831 (O_4831,N_49364,N_49838);
xor UO_4832 (O_4832,N_49885,N_49363);
and UO_4833 (O_4833,N_49004,N_49540);
xnor UO_4834 (O_4834,N_49266,N_49570);
xor UO_4835 (O_4835,N_49670,N_49426);
nor UO_4836 (O_4836,N_49727,N_49764);
nor UO_4837 (O_4837,N_49950,N_49524);
nor UO_4838 (O_4838,N_49629,N_49599);
nor UO_4839 (O_4839,N_49189,N_49728);
nand UO_4840 (O_4840,N_49336,N_49324);
and UO_4841 (O_4841,N_49350,N_49340);
xnor UO_4842 (O_4842,N_49773,N_49710);
or UO_4843 (O_4843,N_49524,N_49077);
or UO_4844 (O_4844,N_49027,N_49496);
nor UO_4845 (O_4845,N_49704,N_49861);
nor UO_4846 (O_4846,N_49633,N_49896);
or UO_4847 (O_4847,N_49820,N_49065);
nand UO_4848 (O_4848,N_49601,N_49236);
and UO_4849 (O_4849,N_49328,N_49949);
nand UO_4850 (O_4850,N_49731,N_49192);
and UO_4851 (O_4851,N_49938,N_49731);
or UO_4852 (O_4852,N_49601,N_49813);
nand UO_4853 (O_4853,N_49033,N_49448);
nor UO_4854 (O_4854,N_49741,N_49456);
xnor UO_4855 (O_4855,N_49337,N_49523);
nor UO_4856 (O_4856,N_49526,N_49066);
nand UO_4857 (O_4857,N_49471,N_49460);
nor UO_4858 (O_4858,N_49432,N_49652);
xnor UO_4859 (O_4859,N_49753,N_49174);
nand UO_4860 (O_4860,N_49373,N_49547);
nand UO_4861 (O_4861,N_49951,N_49346);
or UO_4862 (O_4862,N_49361,N_49895);
or UO_4863 (O_4863,N_49917,N_49885);
nand UO_4864 (O_4864,N_49831,N_49641);
and UO_4865 (O_4865,N_49895,N_49977);
nor UO_4866 (O_4866,N_49080,N_49941);
nor UO_4867 (O_4867,N_49558,N_49475);
and UO_4868 (O_4868,N_49055,N_49660);
xnor UO_4869 (O_4869,N_49277,N_49316);
nand UO_4870 (O_4870,N_49052,N_49333);
nor UO_4871 (O_4871,N_49615,N_49225);
nor UO_4872 (O_4872,N_49919,N_49687);
nor UO_4873 (O_4873,N_49434,N_49215);
and UO_4874 (O_4874,N_49593,N_49536);
nand UO_4875 (O_4875,N_49705,N_49442);
nor UO_4876 (O_4876,N_49526,N_49437);
and UO_4877 (O_4877,N_49788,N_49514);
nor UO_4878 (O_4878,N_49923,N_49959);
and UO_4879 (O_4879,N_49970,N_49654);
xnor UO_4880 (O_4880,N_49444,N_49360);
nand UO_4881 (O_4881,N_49612,N_49492);
xor UO_4882 (O_4882,N_49579,N_49853);
xnor UO_4883 (O_4883,N_49175,N_49149);
nor UO_4884 (O_4884,N_49368,N_49574);
or UO_4885 (O_4885,N_49868,N_49237);
nand UO_4886 (O_4886,N_49295,N_49970);
nor UO_4887 (O_4887,N_49819,N_49162);
nand UO_4888 (O_4888,N_49885,N_49722);
or UO_4889 (O_4889,N_49290,N_49140);
xnor UO_4890 (O_4890,N_49509,N_49862);
nand UO_4891 (O_4891,N_49291,N_49882);
or UO_4892 (O_4892,N_49444,N_49447);
nand UO_4893 (O_4893,N_49938,N_49745);
xor UO_4894 (O_4894,N_49199,N_49188);
or UO_4895 (O_4895,N_49988,N_49905);
nor UO_4896 (O_4896,N_49718,N_49758);
nor UO_4897 (O_4897,N_49965,N_49496);
and UO_4898 (O_4898,N_49493,N_49302);
nand UO_4899 (O_4899,N_49479,N_49402);
and UO_4900 (O_4900,N_49022,N_49470);
and UO_4901 (O_4901,N_49424,N_49202);
and UO_4902 (O_4902,N_49977,N_49811);
nor UO_4903 (O_4903,N_49086,N_49406);
nor UO_4904 (O_4904,N_49094,N_49066);
or UO_4905 (O_4905,N_49370,N_49660);
and UO_4906 (O_4906,N_49053,N_49719);
and UO_4907 (O_4907,N_49299,N_49913);
and UO_4908 (O_4908,N_49483,N_49105);
and UO_4909 (O_4909,N_49786,N_49870);
nand UO_4910 (O_4910,N_49228,N_49594);
xor UO_4911 (O_4911,N_49843,N_49295);
nand UO_4912 (O_4912,N_49964,N_49918);
nor UO_4913 (O_4913,N_49708,N_49062);
nor UO_4914 (O_4914,N_49428,N_49678);
or UO_4915 (O_4915,N_49557,N_49985);
xnor UO_4916 (O_4916,N_49375,N_49503);
nand UO_4917 (O_4917,N_49841,N_49913);
nand UO_4918 (O_4918,N_49723,N_49906);
and UO_4919 (O_4919,N_49014,N_49520);
nor UO_4920 (O_4920,N_49118,N_49366);
or UO_4921 (O_4921,N_49305,N_49188);
nor UO_4922 (O_4922,N_49749,N_49857);
nand UO_4923 (O_4923,N_49143,N_49016);
and UO_4924 (O_4924,N_49819,N_49429);
xor UO_4925 (O_4925,N_49550,N_49333);
xor UO_4926 (O_4926,N_49392,N_49276);
nand UO_4927 (O_4927,N_49813,N_49668);
xor UO_4928 (O_4928,N_49329,N_49990);
nand UO_4929 (O_4929,N_49877,N_49264);
nor UO_4930 (O_4930,N_49978,N_49332);
or UO_4931 (O_4931,N_49595,N_49579);
and UO_4932 (O_4932,N_49393,N_49814);
nor UO_4933 (O_4933,N_49216,N_49792);
nand UO_4934 (O_4934,N_49312,N_49825);
xnor UO_4935 (O_4935,N_49313,N_49244);
or UO_4936 (O_4936,N_49298,N_49581);
xnor UO_4937 (O_4937,N_49518,N_49683);
xnor UO_4938 (O_4938,N_49856,N_49639);
nand UO_4939 (O_4939,N_49038,N_49611);
and UO_4940 (O_4940,N_49780,N_49733);
nor UO_4941 (O_4941,N_49323,N_49790);
and UO_4942 (O_4942,N_49676,N_49461);
xor UO_4943 (O_4943,N_49950,N_49169);
xnor UO_4944 (O_4944,N_49622,N_49062);
xnor UO_4945 (O_4945,N_49873,N_49764);
and UO_4946 (O_4946,N_49311,N_49725);
nand UO_4947 (O_4947,N_49650,N_49118);
and UO_4948 (O_4948,N_49797,N_49439);
nor UO_4949 (O_4949,N_49908,N_49676);
and UO_4950 (O_4950,N_49400,N_49040);
nor UO_4951 (O_4951,N_49527,N_49119);
and UO_4952 (O_4952,N_49709,N_49771);
nor UO_4953 (O_4953,N_49136,N_49284);
and UO_4954 (O_4954,N_49293,N_49285);
nand UO_4955 (O_4955,N_49939,N_49481);
nand UO_4956 (O_4956,N_49255,N_49352);
nor UO_4957 (O_4957,N_49064,N_49437);
nor UO_4958 (O_4958,N_49529,N_49036);
xor UO_4959 (O_4959,N_49328,N_49046);
nand UO_4960 (O_4960,N_49865,N_49421);
and UO_4961 (O_4961,N_49773,N_49163);
xor UO_4962 (O_4962,N_49492,N_49571);
and UO_4963 (O_4963,N_49017,N_49084);
or UO_4964 (O_4964,N_49046,N_49561);
and UO_4965 (O_4965,N_49378,N_49833);
and UO_4966 (O_4966,N_49593,N_49758);
or UO_4967 (O_4967,N_49178,N_49530);
nor UO_4968 (O_4968,N_49610,N_49662);
nand UO_4969 (O_4969,N_49646,N_49637);
nor UO_4970 (O_4970,N_49064,N_49442);
xor UO_4971 (O_4971,N_49543,N_49207);
or UO_4972 (O_4972,N_49572,N_49881);
nor UO_4973 (O_4973,N_49660,N_49948);
xnor UO_4974 (O_4974,N_49090,N_49929);
nand UO_4975 (O_4975,N_49848,N_49635);
or UO_4976 (O_4976,N_49801,N_49545);
nor UO_4977 (O_4977,N_49099,N_49240);
xor UO_4978 (O_4978,N_49907,N_49491);
nor UO_4979 (O_4979,N_49880,N_49371);
xnor UO_4980 (O_4980,N_49991,N_49600);
nand UO_4981 (O_4981,N_49299,N_49313);
nor UO_4982 (O_4982,N_49618,N_49462);
nand UO_4983 (O_4983,N_49899,N_49833);
xor UO_4984 (O_4984,N_49232,N_49625);
nor UO_4985 (O_4985,N_49712,N_49766);
and UO_4986 (O_4986,N_49640,N_49087);
nor UO_4987 (O_4987,N_49071,N_49009);
and UO_4988 (O_4988,N_49345,N_49199);
nor UO_4989 (O_4989,N_49480,N_49534);
xnor UO_4990 (O_4990,N_49862,N_49811);
xor UO_4991 (O_4991,N_49027,N_49883);
xor UO_4992 (O_4992,N_49916,N_49442);
xor UO_4993 (O_4993,N_49447,N_49973);
xnor UO_4994 (O_4994,N_49052,N_49652);
and UO_4995 (O_4995,N_49864,N_49744);
xnor UO_4996 (O_4996,N_49897,N_49772);
and UO_4997 (O_4997,N_49230,N_49779);
and UO_4998 (O_4998,N_49585,N_49112);
nand UO_4999 (O_4999,N_49557,N_49635);
endmodule