module basic_1000_10000_1500_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_944,In_862);
xnor U1 (N_1,In_252,In_710);
xnor U2 (N_2,In_453,In_0);
nand U3 (N_3,In_620,In_288);
and U4 (N_4,In_557,In_977);
or U5 (N_5,In_326,In_256);
nor U6 (N_6,In_970,In_383);
nor U7 (N_7,In_184,In_425);
nor U8 (N_8,In_522,In_817);
or U9 (N_9,In_518,In_692);
nor U10 (N_10,In_319,In_8);
xnor U11 (N_11,In_180,In_437);
and U12 (N_12,In_962,In_896);
or U13 (N_13,In_119,In_534);
or U14 (N_14,In_146,In_483);
nand U15 (N_15,In_279,In_237);
xnor U16 (N_16,In_428,In_596);
or U17 (N_17,In_148,In_354);
nor U18 (N_18,In_983,In_638);
or U19 (N_19,In_418,In_512);
nand U20 (N_20,In_276,In_766);
nand U21 (N_21,In_703,In_650);
xnor U22 (N_22,In_565,In_982);
nand U23 (N_23,In_786,In_932);
nand U24 (N_24,In_948,In_574);
xor U25 (N_25,In_716,In_702);
xor U26 (N_26,In_395,In_517);
xnor U27 (N_27,In_992,In_116);
nand U28 (N_28,In_743,In_617);
nor U29 (N_29,In_22,In_471);
or U30 (N_30,In_888,In_622);
xnor U31 (N_31,In_836,In_723);
or U32 (N_32,In_771,In_975);
nor U33 (N_33,In_467,In_449);
xor U34 (N_34,In_285,In_464);
nor U35 (N_35,In_774,In_839);
and U36 (N_36,In_752,In_226);
nand U37 (N_37,In_735,In_876);
nor U38 (N_38,In_451,In_742);
nand U39 (N_39,In_287,In_871);
xnor U40 (N_40,In_583,In_782);
or U41 (N_41,In_657,In_588);
nor U42 (N_42,In_481,In_36);
or U43 (N_43,In_582,In_34);
nand U44 (N_44,In_893,In_753);
or U45 (N_45,In_155,In_928);
and U46 (N_46,In_333,In_814);
nand U47 (N_47,In_535,In_648);
and U48 (N_48,In_589,In_159);
xor U49 (N_49,In_682,In_853);
or U50 (N_50,In_821,In_442);
nand U51 (N_51,In_974,In_934);
nor U52 (N_52,In_851,In_731);
nand U53 (N_53,In_502,In_441);
xnor U54 (N_54,In_128,In_688);
xor U55 (N_55,In_619,In_967);
nand U56 (N_56,In_640,In_216);
and U57 (N_57,In_706,In_564);
and U58 (N_58,In_163,In_651);
xor U59 (N_59,In_533,In_584);
xor U60 (N_60,In_199,In_487);
nand U61 (N_61,In_40,In_403);
nand U62 (N_62,In_310,In_980);
xor U63 (N_63,In_892,In_624);
nand U64 (N_64,In_318,In_173);
nand U65 (N_65,In_505,In_834);
xnor U66 (N_66,In_768,In_811);
xor U67 (N_67,In_592,In_496);
nor U68 (N_68,In_99,In_431);
or U69 (N_69,In_791,In_795);
or U70 (N_70,In_719,In_833);
nor U71 (N_71,In_936,In_515);
xor U72 (N_72,In_826,In_749);
nor U73 (N_73,In_604,In_446);
and U74 (N_74,In_764,In_633);
xnor U75 (N_75,In_520,In_423);
nand U76 (N_76,In_745,In_664);
nor U77 (N_77,In_578,In_13);
and U78 (N_78,In_73,In_626);
nor U79 (N_79,In_772,In_837);
nand U80 (N_80,In_72,In_410);
nor U81 (N_81,In_486,In_259);
nor U82 (N_82,In_990,In_891);
or U83 (N_83,In_438,In_755);
nand U84 (N_84,In_57,In_910);
or U85 (N_85,In_981,In_819);
nand U86 (N_86,In_636,In_142);
nor U87 (N_87,In_368,In_358);
and U88 (N_88,In_705,In_976);
nand U89 (N_89,In_166,In_314);
or U90 (N_90,In_445,In_639);
and U91 (N_91,In_218,In_929);
nor U92 (N_92,In_879,In_661);
xnor U93 (N_93,In_615,In_769);
nor U94 (N_94,In_24,In_290);
nand U95 (N_95,In_689,In_874);
or U96 (N_96,In_351,In_201);
xor U97 (N_97,In_634,In_525);
and U98 (N_98,In_586,In_371);
and U99 (N_99,In_240,In_920);
and U100 (N_100,In_452,In_537);
nand U101 (N_101,In_60,In_5);
and U102 (N_102,In_642,In_379);
and U103 (N_103,In_775,In_221);
and U104 (N_104,In_317,In_440);
nand U105 (N_105,In_687,In_31);
xnor U106 (N_106,In_92,In_516);
nand U107 (N_107,In_540,In_866);
nand U108 (N_108,In_567,In_978);
or U109 (N_109,In_720,In_124);
nand U110 (N_110,In_426,In_511);
xor U111 (N_111,In_998,In_391);
nand U112 (N_112,In_649,In_385);
nor U113 (N_113,In_543,In_121);
xnor U114 (N_114,In_239,In_448);
xor U115 (N_115,In_396,In_204);
or U116 (N_116,In_341,In_925);
or U117 (N_117,In_222,In_591);
nand U118 (N_118,In_647,In_541);
xor U119 (N_119,In_299,In_562);
or U120 (N_120,In_644,In_889);
nor U121 (N_121,In_363,In_744);
nor U122 (N_122,In_253,In_832);
and U123 (N_123,In_727,In_169);
and U124 (N_124,In_924,In_508);
xor U125 (N_125,In_114,In_472);
and U126 (N_126,In_713,In_190);
and U127 (N_127,In_968,In_227);
and U128 (N_128,In_304,In_10);
or U129 (N_129,In_219,In_401);
and U130 (N_130,In_278,In_918);
nor U131 (N_131,In_74,In_366);
and U132 (N_132,In_105,In_233);
nand U133 (N_133,In_316,In_556);
nand U134 (N_134,In_264,In_329);
xnor U135 (N_135,In_570,In_77);
nand U136 (N_136,In_873,In_645);
nand U137 (N_137,In_608,In_656);
nand U138 (N_138,In_677,In_504);
nor U139 (N_139,In_193,In_544);
nand U140 (N_140,In_51,In_254);
and U141 (N_141,In_457,In_497);
xor U142 (N_142,In_229,In_64);
and U143 (N_143,In_463,In_308);
and U144 (N_144,In_359,In_773);
xnor U145 (N_145,In_777,In_84);
and U146 (N_146,In_156,In_653);
xor U147 (N_147,In_182,In_849);
or U148 (N_148,In_154,In_600);
and U149 (N_149,In_272,In_914);
nor U150 (N_150,In_262,In_711);
xor U151 (N_151,In_337,In_215);
nor U152 (N_152,In_20,In_922);
nand U153 (N_153,In_965,In_784);
nand U154 (N_154,In_126,In_315);
and U155 (N_155,In_205,In_323);
or U156 (N_156,In_546,In_59);
and U157 (N_157,In_946,In_112);
or U158 (N_158,In_738,In_629);
nand U159 (N_159,In_271,In_460);
nand U160 (N_160,In_655,In_740);
nand U161 (N_161,In_248,In_593);
and U162 (N_162,In_579,In_123);
xor U163 (N_163,In_381,In_898);
nand U164 (N_164,In_686,In_700);
and U165 (N_165,In_200,In_654);
or U166 (N_166,In_151,In_364);
or U167 (N_167,In_869,In_999);
nand U168 (N_168,In_170,In_513);
nor U169 (N_169,In_660,In_760);
and U170 (N_170,In_214,In_375);
or U171 (N_171,In_963,In_959);
nand U172 (N_172,In_954,In_841);
or U173 (N_173,In_859,In_850);
nor U174 (N_174,In_38,In_98);
nand U175 (N_175,In_815,In_294);
and U176 (N_176,In_408,In_186);
nand U177 (N_177,In_61,In_307);
nor U178 (N_178,In_397,In_41);
xnor U179 (N_179,In_812,In_28);
nor U180 (N_180,In_996,In_236);
xnor U181 (N_181,In_960,In_985);
nor U182 (N_182,In_547,In_790);
xnor U183 (N_183,In_691,In_210);
nor U184 (N_184,In_606,In_127);
nor U185 (N_185,In_906,In_627);
nor U186 (N_186,In_11,In_417);
nor U187 (N_187,In_4,In_113);
nor U188 (N_188,In_348,In_658);
and U189 (N_189,In_66,In_320);
or U190 (N_190,In_412,In_150);
or U191 (N_191,In_132,In_915);
nand U192 (N_192,In_637,In_115);
xnor U193 (N_193,In_555,In_454);
and U194 (N_194,In_803,In_257);
and U195 (N_195,In_529,In_781);
nand U196 (N_196,In_730,In_697);
and U197 (N_197,In_350,In_389);
and U198 (N_198,In_701,In_185);
nand U199 (N_199,In_572,In_88);
nand U200 (N_200,In_599,In_663);
nand U201 (N_201,In_933,In_545);
and U202 (N_202,In_286,In_455);
or U203 (N_203,In_824,In_554);
xnor U204 (N_204,In_714,In_799);
xor U205 (N_205,In_942,In_949);
or U206 (N_206,In_133,In_797);
and U207 (N_207,In_900,In_693);
nor U208 (N_208,In_217,In_461);
and U209 (N_209,In_712,In_208);
nand U210 (N_210,In_748,In_103);
and U211 (N_211,In_152,In_203);
nand U212 (N_212,In_552,In_695);
and U213 (N_213,In_856,In_979);
and U214 (N_214,In_957,In_779);
or U215 (N_215,In_756,In_507);
nor U216 (N_216,In_872,In_561);
or U217 (N_217,In_206,In_668);
xor U218 (N_218,In_414,In_804);
and U219 (N_219,In_830,In_725);
nand U220 (N_220,In_322,In_147);
and U221 (N_221,In_984,In_228);
and U222 (N_222,In_298,In_842);
or U223 (N_223,In_794,In_598);
nor U224 (N_224,In_607,In_458);
or U225 (N_225,In_39,In_443);
or U226 (N_226,In_400,In_573);
and U227 (N_227,In_757,In_831);
xor U228 (N_228,In_82,In_388);
nand U229 (N_229,In_83,In_117);
or U230 (N_230,In_491,In_519);
nand U231 (N_231,In_882,In_739);
or U232 (N_232,In_699,In_243);
or U233 (N_233,In_476,In_536);
nor U234 (N_234,In_490,In_413);
nor U235 (N_235,In_224,In_136);
nand U236 (N_236,In_630,In_747);
xnor U237 (N_237,In_498,In_857);
xor U238 (N_238,In_93,In_244);
or U239 (N_239,In_56,In_897);
or U240 (N_240,In_792,In_746);
xor U241 (N_241,In_347,In_800);
or U242 (N_242,In_602,In_346);
or U243 (N_243,In_376,In_96);
nand U244 (N_244,In_75,In_390);
and U245 (N_245,In_62,In_432);
nor U246 (N_246,In_296,In_673);
xnor U247 (N_247,In_838,In_282);
xor U248 (N_248,In_269,In_191);
and U249 (N_249,In_104,In_265);
nor U250 (N_250,In_85,In_274);
nand U251 (N_251,In_895,In_16);
nand U252 (N_252,In_450,In_762);
xor U253 (N_253,In_931,In_338);
and U254 (N_254,In_494,In_58);
xnor U255 (N_255,In_245,In_676);
nor U256 (N_256,In_958,In_503);
nor U257 (N_257,In_17,In_788);
nand U258 (N_258,In_377,In_662);
and U259 (N_259,In_621,In_171);
nand U260 (N_260,In_175,In_548);
xnor U261 (N_261,In_281,In_101);
xnor U262 (N_262,In_109,In_7);
nand U263 (N_263,In_560,In_46);
xor U264 (N_264,In_987,In_192);
and U265 (N_265,In_421,In_801);
nor U266 (N_266,In_181,In_538);
xor U267 (N_267,In_2,In_724);
or U268 (N_268,In_683,In_30);
nand U269 (N_269,In_671,In_902);
nand U270 (N_270,In_230,In_696);
nor U271 (N_271,In_751,In_631);
nor U272 (N_272,In_776,In_580);
nor U273 (N_273,In_409,In_309);
xor U274 (N_274,In_118,In_386);
nand U275 (N_275,In_829,In_986);
and U276 (N_276,In_167,In_581);
nor U277 (N_277,In_488,In_867);
and U278 (N_278,In_447,In_48);
nor U279 (N_279,In_94,In_275);
nor U280 (N_280,In_300,In_336);
and U281 (N_281,In_793,In_852);
and U282 (N_282,In_251,In_726);
or U283 (N_283,In_153,In_531);
and U284 (N_284,In_951,In_27);
nand U285 (N_285,In_137,In_950);
or U286 (N_286,In_258,In_340);
or U287 (N_287,In_179,In_997);
xor U288 (N_288,In_667,In_177);
nand U289 (N_289,In_162,In_249);
and U290 (N_290,In_209,In_884);
nor U291 (N_291,In_378,In_71);
and U292 (N_292,In_477,In_609);
and U293 (N_293,In_325,In_816);
nor U294 (N_294,In_405,In_553);
or U295 (N_295,In_903,In_911);
nand U296 (N_296,In_614,In_969);
or U297 (N_297,In_909,In_825);
xnor U298 (N_298,In_270,In_131);
and U299 (N_299,In_666,In_835);
nor U300 (N_300,In_549,In_674);
or U301 (N_301,In_35,In_44);
and U302 (N_302,In_69,In_569);
nor U303 (N_303,In_344,In_904);
and U304 (N_304,In_384,In_875);
nor U305 (N_305,In_189,In_12);
xnor U306 (N_306,In_301,In_550);
and U307 (N_307,In_780,In_164);
or U308 (N_308,In_349,In_1);
xnor U309 (N_309,In_763,In_860);
and U310 (N_310,In_945,In_19);
nand U311 (N_311,In_357,In_809);
nor U312 (N_312,In_321,In_612);
and U313 (N_313,In_665,In_844);
and U314 (N_314,In_362,In_42);
xnor U315 (N_315,In_704,In_225);
nor U316 (N_316,In_961,In_439);
nor U317 (N_317,In_989,In_174);
xnor U318 (N_318,In_994,In_901);
or U319 (N_319,In_15,In_563);
and U320 (N_320,In_802,In_292);
nor U321 (N_321,In_459,In_652);
xor U322 (N_322,In_427,In_480);
xnor U323 (N_323,In_886,In_238);
nand U324 (N_324,In_670,In_474);
nor U325 (N_325,In_865,In_473);
and U326 (N_326,In_778,In_495);
or U327 (N_327,In_890,In_313);
or U328 (N_328,In_411,In_345);
nand U329 (N_329,In_528,In_947);
nand U330 (N_330,In_685,In_469);
xor U331 (N_331,In_334,In_161);
nor U332 (N_332,In_9,In_930);
nor U333 (N_333,In_927,In_404);
nor U334 (N_334,In_659,In_143);
nand U335 (N_335,In_732,In_370);
or U336 (N_336,In_47,In_361);
or U337 (N_337,In_302,In_595);
nor U338 (N_338,In_953,In_241);
xnor U339 (N_339,In_770,In_880);
nor U340 (N_340,In_32,In_107);
and U341 (N_341,In_721,In_235);
nand U342 (N_342,In_306,In_263);
or U343 (N_343,In_289,In_372);
xor U344 (N_344,In_616,In_500);
nand U345 (N_345,In_509,In_168);
nor U346 (N_346,In_941,In_149);
xnor U347 (N_347,In_669,In_679);
and U348 (N_348,In_466,In_144);
xor U349 (N_349,In_356,In_178);
or U350 (N_350,In_387,In_157);
xnor U351 (N_351,In_273,In_202);
nand U352 (N_352,In_160,In_327);
nand U353 (N_353,In_808,In_926);
xnor U354 (N_354,In_484,In_135);
xnor U355 (N_355,In_172,In_328);
or U356 (N_356,In_861,In_758);
nor U357 (N_357,In_729,In_767);
and U358 (N_358,In_183,In_165);
nor U359 (N_359,In_232,In_848);
nor U360 (N_360,In_37,In_899);
and U361 (N_361,In_995,In_76);
and U362 (N_362,In_955,In_733);
or U363 (N_363,In_759,In_303);
nor U364 (N_364,In_736,In_722);
xor U365 (N_365,In_125,In_416);
and U366 (N_366,In_475,In_806);
xor U367 (N_367,In_120,In_470);
and U368 (N_368,In_810,In_43);
nand U369 (N_369,In_331,In_65);
nand U370 (N_370,In_694,In_293);
nand U371 (N_371,In_524,In_80);
or U372 (N_372,In_330,In_242);
nor U373 (N_373,In_87,In_95);
and U374 (N_374,In_559,In_90);
nor U375 (N_375,In_89,In_324);
and U376 (N_376,In_130,In_988);
nor U377 (N_377,In_392,In_485);
and U378 (N_378,In_420,In_878);
nand U379 (N_379,In_680,In_158);
and U380 (N_380,In_6,In_684);
nor U381 (N_381,In_335,In_29);
xnor U382 (N_382,In_715,In_122);
nand U383 (N_383,In_250,In_374);
nor U384 (N_384,In_50,In_939);
xnor U385 (N_385,In_81,In_912);
xnor U386 (N_386,In_501,In_741);
xor U387 (N_387,In_868,In_21);
xor U388 (N_388,In_971,In_261);
xnor U389 (N_389,In_681,In_526);
nor U390 (N_390,In_785,In_643);
or U391 (N_391,In_108,In_863);
xnor U392 (N_392,In_68,In_618);
xnor U393 (N_393,In_576,In_641);
and U394 (N_394,In_141,In_295);
xnor U395 (N_395,In_212,In_594);
nor U396 (N_396,In_291,In_787);
xnor U397 (N_397,In_601,In_921);
nor U398 (N_398,In_415,In_539);
nand U399 (N_399,In_367,In_196);
nand U400 (N_400,In_365,In_25);
xnor U401 (N_401,In_91,In_422);
and U402 (N_402,In_530,In_840);
nor U403 (N_403,In_943,In_129);
and U404 (N_404,In_690,In_194);
and U405 (N_405,In_737,In_623);
nor U406 (N_406,In_429,In_462);
or U407 (N_407,In_937,In_783);
nor U408 (N_408,In_398,In_499);
xnor U409 (N_409,In_907,In_393);
xnor U410 (N_410,In_964,In_352);
nor U411 (N_411,In_635,In_268);
and U412 (N_412,In_106,In_585);
nor U413 (N_413,In_284,In_870);
nor U414 (N_414,In_603,In_198);
nand U415 (N_415,In_728,In_956);
or U416 (N_416,In_577,In_283);
nor U417 (N_417,In_188,In_54);
xnor U418 (N_418,In_465,In_332);
nor U419 (N_419,In_993,In_718);
xnor U420 (N_420,In_482,In_887);
and U421 (N_421,In_138,In_207);
nor U422 (N_422,In_672,In_823);
nand U423 (N_423,In_197,In_223);
and U424 (N_424,In_33,In_613);
and U425 (N_425,In_708,In_877);
or U426 (N_426,In_605,In_843);
nor U427 (N_427,In_807,In_813);
and U428 (N_428,In_456,In_312);
xor U429 (N_429,In_492,In_646);
nand U430 (N_430,In_858,In_246);
xnor U431 (N_431,In_435,In_267);
xor U432 (N_432,In_514,In_430);
or U433 (N_433,In_632,In_266);
or U434 (N_434,In_940,In_220);
nand U435 (N_435,In_991,In_966);
xor U436 (N_436,In_493,In_847);
and U437 (N_437,In_894,In_628);
xor U438 (N_438,In_145,In_213);
nor U439 (N_439,In_542,In_3);
and U440 (N_440,In_527,In_734);
and U441 (N_441,In_311,In_952);
or U442 (N_442,In_489,In_187);
and U443 (N_443,In_297,In_818);
nor U444 (N_444,In_63,In_369);
or U445 (N_445,In_881,In_305);
or U446 (N_446,In_339,In_855);
nand U447 (N_447,In_709,In_231);
nor U448 (N_448,In_765,In_255);
nand U449 (N_449,In_78,In_406);
or U450 (N_450,In_67,In_399);
nor U451 (N_451,In_551,In_247);
nand U452 (N_452,In_566,In_407);
or U453 (N_453,In_343,In_805);
or U454 (N_454,In_18,In_134);
nor U455 (N_455,In_611,In_521);
and U456 (N_456,In_49,In_45);
xor U457 (N_457,In_761,In_822);
xnor U458 (N_458,In_575,In_913);
xnor U459 (N_459,In_26,In_14);
nand U460 (N_460,In_885,In_789);
and U461 (N_461,In_798,In_360);
xor U462 (N_462,In_590,In_973);
nor U463 (N_463,In_625,In_854);
xnor U464 (N_464,In_434,In_111);
and U465 (N_465,In_917,In_678);
xnor U466 (N_466,In_923,In_234);
or U467 (N_467,In_707,In_610);
xor U468 (N_468,In_820,In_479);
nand U469 (N_469,In_23,In_510);
or U470 (N_470,In_382,In_717);
or U471 (N_471,In_828,In_597);
or U472 (N_472,In_587,In_845);
and U473 (N_473,In_433,In_100);
or U474 (N_474,In_280,In_478);
and U475 (N_475,In_698,In_139);
or U476 (N_476,In_86,In_52);
or U477 (N_477,In_277,In_846);
nand U478 (N_478,In_55,In_506);
nor U479 (N_479,In_394,In_140);
nand U480 (N_480,In_97,In_79);
nor U481 (N_481,In_675,In_373);
xor U482 (N_482,In_468,In_905);
nor U483 (N_483,In_796,In_754);
xor U484 (N_484,In_353,In_195);
and U485 (N_485,In_935,In_750);
nand U486 (N_486,In_355,In_419);
nor U487 (N_487,In_919,In_916);
nand U488 (N_488,In_402,In_424);
or U489 (N_489,In_176,In_444);
or U490 (N_490,In_260,In_938);
or U491 (N_491,In_827,In_70);
or U492 (N_492,In_342,In_436);
nand U493 (N_493,In_102,In_523);
nor U494 (N_494,In_568,In_532);
xnor U495 (N_495,In_883,In_864);
nor U496 (N_496,In_211,In_53);
and U497 (N_497,In_380,In_571);
nor U498 (N_498,In_972,In_110);
or U499 (N_499,In_558,In_908);
nand U500 (N_500,In_157,In_491);
nand U501 (N_501,In_485,In_923);
xor U502 (N_502,In_977,In_884);
xor U503 (N_503,In_676,In_622);
xnor U504 (N_504,In_560,In_302);
nor U505 (N_505,In_867,In_894);
or U506 (N_506,In_778,In_928);
and U507 (N_507,In_626,In_718);
or U508 (N_508,In_610,In_173);
and U509 (N_509,In_540,In_877);
nor U510 (N_510,In_371,In_540);
nor U511 (N_511,In_312,In_378);
and U512 (N_512,In_980,In_117);
xnor U513 (N_513,In_377,In_721);
or U514 (N_514,In_975,In_998);
nand U515 (N_515,In_29,In_131);
or U516 (N_516,In_536,In_876);
and U517 (N_517,In_451,In_409);
xnor U518 (N_518,In_907,In_712);
or U519 (N_519,In_778,In_782);
nor U520 (N_520,In_953,In_539);
and U521 (N_521,In_781,In_589);
and U522 (N_522,In_51,In_858);
and U523 (N_523,In_431,In_376);
xor U524 (N_524,In_267,In_88);
nor U525 (N_525,In_3,In_271);
nor U526 (N_526,In_369,In_880);
or U527 (N_527,In_876,In_216);
or U528 (N_528,In_760,In_351);
nor U529 (N_529,In_221,In_631);
and U530 (N_530,In_843,In_989);
or U531 (N_531,In_587,In_778);
or U532 (N_532,In_28,In_757);
and U533 (N_533,In_791,In_752);
nand U534 (N_534,In_601,In_657);
nand U535 (N_535,In_289,In_406);
and U536 (N_536,In_64,In_298);
or U537 (N_537,In_716,In_875);
and U538 (N_538,In_421,In_215);
nor U539 (N_539,In_649,In_745);
nand U540 (N_540,In_339,In_638);
or U541 (N_541,In_78,In_73);
nor U542 (N_542,In_618,In_300);
or U543 (N_543,In_837,In_914);
nor U544 (N_544,In_9,In_938);
xor U545 (N_545,In_449,In_977);
xor U546 (N_546,In_514,In_769);
xnor U547 (N_547,In_442,In_260);
nand U548 (N_548,In_359,In_695);
nor U549 (N_549,In_366,In_848);
nor U550 (N_550,In_161,In_831);
nor U551 (N_551,In_633,In_935);
xor U552 (N_552,In_429,In_866);
nand U553 (N_553,In_177,In_373);
xor U554 (N_554,In_508,In_986);
or U555 (N_555,In_812,In_294);
and U556 (N_556,In_965,In_694);
nand U557 (N_557,In_947,In_358);
and U558 (N_558,In_138,In_813);
or U559 (N_559,In_891,In_468);
nor U560 (N_560,In_777,In_338);
nor U561 (N_561,In_699,In_322);
xor U562 (N_562,In_395,In_956);
nor U563 (N_563,In_124,In_757);
nor U564 (N_564,In_817,In_414);
and U565 (N_565,In_857,In_213);
nand U566 (N_566,In_907,In_546);
and U567 (N_567,In_880,In_722);
or U568 (N_568,In_201,In_71);
xnor U569 (N_569,In_195,In_79);
nor U570 (N_570,In_803,In_474);
nand U571 (N_571,In_11,In_378);
or U572 (N_572,In_491,In_516);
and U573 (N_573,In_756,In_522);
xnor U574 (N_574,In_364,In_377);
xnor U575 (N_575,In_727,In_486);
xor U576 (N_576,In_151,In_36);
and U577 (N_577,In_491,In_645);
xor U578 (N_578,In_824,In_961);
nand U579 (N_579,In_320,In_148);
xnor U580 (N_580,In_352,In_436);
or U581 (N_581,In_177,In_767);
and U582 (N_582,In_717,In_769);
xnor U583 (N_583,In_121,In_621);
nand U584 (N_584,In_488,In_911);
and U585 (N_585,In_788,In_555);
xor U586 (N_586,In_641,In_740);
or U587 (N_587,In_549,In_425);
and U588 (N_588,In_911,In_285);
nor U589 (N_589,In_281,In_191);
nand U590 (N_590,In_438,In_946);
and U591 (N_591,In_922,In_685);
xnor U592 (N_592,In_854,In_642);
or U593 (N_593,In_876,In_994);
nor U594 (N_594,In_677,In_934);
or U595 (N_595,In_545,In_446);
or U596 (N_596,In_688,In_638);
or U597 (N_597,In_467,In_102);
xor U598 (N_598,In_209,In_190);
and U599 (N_599,In_242,In_603);
and U600 (N_600,In_208,In_479);
and U601 (N_601,In_964,In_297);
or U602 (N_602,In_115,In_486);
nand U603 (N_603,In_857,In_649);
and U604 (N_604,In_160,In_417);
and U605 (N_605,In_119,In_53);
nor U606 (N_606,In_985,In_370);
and U607 (N_607,In_107,In_949);
xor U608 (N_608,In_830,In_329);
xnor U609 (N_609,In_232,In_420);
nand U610 (N_610,In_657,In_797);
or U611 (N_611,In_916,In_411);
xnor U612 (N_612,In_906,In_304);
or U613 (N_613,In_664,In_951);
xnor U614 (N_614,In_851,In_468);
or U615 (N_615,In_391,In_833);
xnor U616 (N_616,In_463,In_812);
and U617 (N_617,In_113,In_88);
and U618 (N_618,In_185,In_366);
or U619 (N_619,In_860,In_335);
xnor U620 (N_620,In_359,In_549);
nand U621 (N_621,In_574,In_879);
xnor U622 (N_622,In_419,In_267);
or U623 (N_623,In_399,In_783);
nand U624 (N_624,In_601,In_965);
or U625 (N_625,In_494,In_227);
and U626 (N_626,In_538,In_278);
or U627 (N_627,In_523,In_206);
xor U628 (N_628,In_500,In_783);
nand U629 (N_629,In_426,In_649);
nand U630 (N_630,In_580,In_854);
nor U631 (N_631,In_43,In_360);
xor U632 (N_632,In_656,In_117);
nor U633 (N_633,In_8,In_467);
xor U634 (N_634,In_712,In_732);
or U635 (N_635,In_919,In_630);
nor U636 (N_636,In_46,In_148);
and U637 (N_637,In_64,In_23);
xnor U638 (N_638,In_959,In_583);
nor U639 (N_639,In_868,In_540);
nor U640 (N_640,In_874,In_796);
nor U641 (N_641,In_737,In_590);
and U642 (N_642,In_906,In_440);
and U643 (N_643,In_473,In_509);
or U644 (N_644,In_267,In_196);
xnor U645 (N_645,In_588,In_900);
xor U646 (N_646,In_494,In_318);
xor U647 (N_647,In_298,In_130);
xnor U648 (N_648,In_968,In_159);
nor U649 (N_649,In_331,In_481);
xnor U650 (N_650,In_949,In_672);
nor U651 (N_651,In_857,In_953);
or U652 (N_652,In_966,In_699);
nor U653 (N_653,In_661,In_147);
nor U654 (N_654,In_811,In_272);
and U655 (N_655,In_738,In_219);
xor U656 (N_656,In_235,In_676);
or U657 (N_657,In_460,In_654);
nor U658 (N_658,In_148,In_584);
xor U659 (N_659,In_512,In_947);
xnor U660 (N_660,In_204,In_570);
xor U661 (N_661,In_823,In_650);
nand U662 (N_662,In_312,In_734);
xor U663 (N_663,In_952,In_982);
nor U664 (N_664,In_166,In_588);
xor U665 (N_665,In_684,In_576);
or U666 (N_666,In_308,In_93);
nand U667 (N_667,In_82,In_752);
and U668 (N_668,In_346,In_818);
or U669 (N_669,In_766,In_809);
or U670 (N_670,In_446,In_613);
or U671 (N_671,In_46,In_593);
nand U672 (N_672,In_695,In_127);
and U673 (N_673,In_14,In_64);
and U674 (N_674,In_974,In_76);
nand U675 (N_675,In_923,In_955);
or U676 (N_676,In_812,In_445);
nand U677 (N_677,In_205,In_407);
nor U678 (N_678,In_843,In_907);
or U679 (N_679,In_390,In_588);
nand U680 (N_680,In_438,In_384);
nand U681 (N_681,In_108,In_703);
nand U682 (N_682,In_995,In_973);
or U683 (N_683,In_352,In_781);
and U684 (N_684,In_131,In_246);
xnor U685 (N_685,In_455,In_525);
xor U686 (N_686,In_18,In_837);
and U687 (N_687,In_92,In_491);
nor U688 (N_688,In_605,In_67);
xor U689 (N_689,In_428,In_366);
or U690 (N_690,In_828,In_163);
or U691 (N_691,In_254,In_850);
xor U692 (N_692,In_112,In_234);
xnor U693 (N_693,In_221,In_145);
and U694 (N_694,In_377,In_380);
or U695 (N_695,In_626,In_96);
and U696 (N_696,In_939,In_952);
xor U697 (N_697,In_808,In_123);
nor U698 (N_698,In_841,In_942);
or U699 (N_699,In_922,In_609);
xnor U700 (N_700,In_264,In_987);
and U701 (N_701,In_167,In_548);
and U702 (N_702,In_319,In_203);
xor U703 (N_703,In_129,In_216);
and U704 (N_704,In_958,In_337);
nand U705 (N_705,In_543,In_12);
nand U706 (N_706,In_441,In_212);
nand U707 (N_707,In_999,In_385);
nor U708 (N_708,In_449,In_677);
and U709 (N_709,In_450,In_514);
nand U710 (N_710,In_153,In_49);
nor U711 (N_711,In_318,In_909);
nand U712 (N_712,In_457,In_108);
nor U713 (N_713,In_745,In_114);
nand U714 (N_714,In_13,In_972);
nor U715 (N_715,In_970,In_378);
xor U716 (N_716,In_807,In_856);
and U717 (N_717,In_447,In_856);
or U718 (N_718,In_900,In_893);
nor U719 (N_719,In_300,In_974);
nand U720 (N_720,In_991,In_807);
xor U721 (N_721,In_812,In_572);
and U722 (N_722,In_477,In_980);
nand U723 (N_723,In_427,In_694);
nand U724 (N_724,In_547,In_818);
or U725 (N_725,In_573,In_224);
or U726 (N_726,In_551,In_129);
nor U727 (N_727,In_841,In_91);
nand U728 (N_728,In_750,In_578);
or U729 (N_729,In_153,In_924);
xor U730 (N_730,In_196,In_11);
and U731 (N_731,In_586,In_319);
nor U732 (N_732,In_726,In_401);
or U733 (N_733,In_776,In_570);
nor U734 (N_734,In_970,In_846);
and U735 (N_735,In_316,In_676);
nor U736 (N_736,In_669,In_759);
nand U737 (N_737,In_526,In_370);
and U738 (N_738,In_678,In_204);
or U739 (N_739,In_292,In_974);
nand U740 (N_740,In_307,In_352);
nand U741 (N_741,In_511,In_246);
nor U742 (N_742,In_413,In_149);
nor U743 (N_743,In_893,In_998);
or U744 (N_744,In_615,In_338);
or U745 (N_745,In_306,In_387);
or U746 (N_746,In_967,In_562);
and U747 (N_747,In_439,In_238);
nand U748 (N_748,In_353,In_677);
xor U749 (N_749,In_745,In_396);
nor U750 (N_750,In_81,In_378);
or U751 (N_751,In_428,In_502);
xor U752 (N_752,In_319,In_615);
nand U753 (N_753,In_463,In_323);
xnor U754 (N_754,In_400,In_901);
nor U755 (N_755,In_578,In_265);
and U756 (N_756,In_792,In_16);
and U757 (N_757,In_787,In_564);
and U758 (N_758,In_356,In_273);
nand U759 (N_759,In_157,In_949);
nor U760 (N_760,In_69,In_541);
nor U761 (N_761,In_940,In_879);
nand U762 (N_762,In_104,In_777);
nand U763 (N_763,In_223,In_42);
nor U764 (N_764,In_756,In_136);
or U765 (N_765,In_565,In_701);
and U766 (N_766,In_323,In_837);
or U767 (N_767,In_450,In_527);
nor U768 (N_768,In_15,In_341);
xnor U769 (N_769,In_970,In_142);
xor U770 (N_770,In_664,In_843);
nand U771 (N_771,In_618,In_775);
xor U772 (N_772,In_505,In_808);
or U773 (N_773,In_226,In_671);
and U774 (N_774,In_495,In_592);
xor U775 (N_775,In_644,In_286);
or U776 (N_776,In_576,In_663);
xor U777 (N_777,In_407,In_623);
and U778 (N_778,In_312,In_554);
nor U779 (N_779,In_252,In_277);
nand U780 (N_780,In_617,In_869);
nand U781 (N_781,In_528,In_686);
or U782 (N_782,In_320,In_484);
nor U783 (N_783,In_297,In_201);
xor U784 (N_784,In_878,In_678);
nor U785 (N_785,In_469,In_605);
or U786 (N_786,In_50,In_96);
or U787 (N_787,In_973,In_166);
or U788 (N_788,In_153,In_98);
nor U789 (N_789,In_153,In_296);
nand U790 (N_790,In_771,In_589);
or U791 (N_791,In_576,In_474);
nand U792 (N_792,In_645,In_223);
nor U793 (N_793,In_833,In_86);
and U794 (N_794,In_872,In_981);
xor U795 (N_795,In_174,In_127);
nor U796 (N_796,In_198,In_15);
xnor U797 (N_797,In_465,In_354);
and U798 (N_798,In_445,In_481);
xor U799 (N_799,In_553,In_974);
and U800 (N_800,In_248,In_779);
and U801 (N_801,In_560,In_137);
and U802 (N_802,In_927,In_117);
nor U803 (N_803,In_595,In_347);
and U804 (N_804,In_836,In_220);
nand U805 (N_805,In_288,In_424);
xnor U806 (N_806,In_57,In_830);
nor U807 (N_807,In_736,In_586);
nand U808 (N_808,In_990,In_48);
or U809 (N_809,In_536,In_970);
and U810 (N_810,In_474,In_932);
or U811 (N_811,In_584,In_942);
or U812 (N_812,In_852,In_173);
and U813 (N_813,In_67,In_773);
nor U814 (N_814,In_664,In_37);
nand U815 (N_815,In_349,In_664);
or U816 (N_816,In_191,In_164);
xnor U817 (N_817,In_723,In_680);
nand U818 (N_818,In_89,In_944);
nor U819 (N_819,In_422,In_787);
nor U820 (N_820,In_455,In_369);
nor U821 (N_821,In_861,In_309);
and U822 (N_822,In_336,In_845);
or U823 (N_823,In_8,In_409);
and U824 (N_824,In_844,In_162);
or U825 (N_825,In_197,In_201);
nor U826 (N_826,In_976,In_919);
or U827 (N_827,In_288,In_382);
xnor U828 (N_828,In_74,In_466);
xor U829 (N_829,In_587,In_747);
nor U830 (N_830,In_922,In_810);
nand U831 (N_831,In_651,In_978);
nor U832 (N_832,In_289,In_532);
nand U833 (N_833,In_723,In_780);
or U834 (N_834,In_916,In_92);
xnor U835 (N_835,In_963,In_340);
and U836 (N_836,In_475,In_883);
nand U837 (N_837,In_6,In_958);
nand U838 (N_838,In_958,In_787);
xor U839 (N_839,In_536,In_73);
nor U840 (N_840,In_459,In_679);
xnor U841 (N_841,In_882,In_961);
xor U842 (N_842,In_81,In_753);
and U843 (N_843,In_655,In_573);
or U844 (N_844,In_723,In_75);
nand U845 (N_845,In_995,In_833);
or U846 (N_846,In_66,In_737);
nor U847 (N_847,In_243,In_469);
xor U848 (N_848,In_528,In_478);
nor U849 (N_849,In_857,In_190);
nand U850 (N_850,In_43,In_205);
nand U851 (N_851,In_457,In_202);
nor U852 (N_852,In_250,In_768);
nor U853 (N_853,In_240,In_273);
nor U854 (N_854,In_60,In_382);
nor U855 (N_855,In_342,In_488);
nor U856 (N_856,In_95,In_672);
xor U857 (N_857,In_825,In_926);
nand U858 (N_858,In_847,In_403);
or U859 (N_859,In_279,In_346);
and U860 (N_860,In_788,In_766);
and U861 (N_861,In_406,In_405);
and U862 (N_862,In_775,In_751);
and U863 (N_863,In_766,In_624);
nor U864 (N_864,In_418,In_238);
or U865 (N_865,In_580,In_997);
nand U866 (N_866,In_299,In_161);
xnor U867 (N_867,In_680,In_182);
xor U868 (N_868,In_213,In_493);
and U869 (N_869,In_165,In_636);
nand U870 (N_870,In_378,In_786);
xor U871 (N_871,In_31,In_135);
and U872 (N_872,In_267,In_359);
nand U873 (N_873,In_535,In_927);
or U874 (N_874,In_456,In_217);
and U875 (N_875,In_46,In_618);
or U876 (N_876,In_72,In_832);
or U877 (N_877,In_149,In_137);
xor U878 (N_878,In_829,In_828);
xor U879 (N_879,In_380,In_457);
nor U880 (N_880,In_289,In_469);
nor U881 (N_881,In_390,In_764);
nor U882 (N_882,In_844,In_980);
xor U883 (N_883,In_70,In_652);
or U884 (N_884,In_161,In_673);
xor U885 (N_885,In_897,In_387);
nor U886 (N_886,In_368,In_684);
xor U887 (N_887,In_838,In_199);
nor U888 (N_888,In_215,In_663);
nor U889 (N_889,In_290,In_475);
and U890 (N_890,In_60,In_949);
and U891 (N_891,In_911,In_969);
nor U892 (N_892,In_561,In_370);
or U893 (N_893,In_782,In_762);
and U894 (N_894,In_34,In_672);
nor U895 (N_895,In_186,In_933);
nand U896 (N_896,In_158,In_542);
nor U897 (N_897,In_919,In_588);
nand U898 (N_898,In_980,In_755);
or U899 (N_899,In_303,In_849);
or U900 (N_900,In_222,In_478);
xnor U901 (N_901,In_330,In_961);
nand U902 (N_902,In_826,In_821);
nand U903 (N_903,In_983,In_729);
nand U904 (N_904,In_98,In_309);
xnor U905 (N_905,In_527,In_66);
xnor U906 (N_906,In_900,In_548);
nand U907 (N_907,In_291,In_807);
and U908 (N_908,In_469,In_344);
nand U909 (N_909,In_944,In_627);
nor U910 (N_910,In_911,In_282);
and U911 (N_911,In_444,In_255);
nand U912 (N_912,In_322,In_612);
xor U913 (N_913,In_144,In_952);
and U914 (N_914,In_593,In_762);
xnor U915 (N_915,In_616,In_142);
and U916 (N_916,In_81,In_343);
xnor U917 (N_917,In_917,In_700);
or U918 (N_918,In_698,In_760);
xnor U919 (N_919,In_775,In_188);
xor U920 (N_920,In_745,In_922);
xnor U921 (N_921,In_497,In_563);
or U922 (N_922,In_539,In_671);
and U923 (N_923,In_988,In_853);
nor U924 (N_924,In_181,In_141);
nand U925 (N_925,In_860,In_970);
and U926 (N_926,In_238,In_685);
nand U927 (N_927,In_154,In_247);
or U928 (N_928,In_669,In_342);
nor U929 (N_929,In_803,In_959);
nand U930 (N_930,In_828,In_865);
nor U931 (N_931,In_512,In_874);
and U932 (N_932,In_167,In_833);
nand U933 (N_933,In_706,In_919);
nand U934 (N_934,In_967,In_640);
xnor U935 (N_935,In_619,In_442);
nand U936 (N_936,In_679,In_286);
xor U937 (N_937,In_249,In_727);
nor U938 (N_938,In_343,In_953);
nor U939 (N_939,In_425,In_415);
or U940 (N_940,In_87,In_371);
xnor U941 (N_941,In_714,In_959);
nand U942 (N_942,In_448,In_137);
nand U943 (N_943,In_157,In_363);
and U944 (N_944,In_287,In_317);
or U945 (N_945,In_98,In_182);
nor U946 (N_946,In_161,In_43);
or U947 (N_947,In_416,In_763);
nand U948 (N_948,In_503,In_514);
nand U949 (N_949,In_371,In_25);
nor U950 (N_950,In_53,In_696);
and U951 (N_951,In_995,In_808);
nand U952 (N_952,In_479,In_297);
and U953 (N_953,In_549,In_690);
and U954 (N_954,In_171,In_590);
and U955 (N_955,In_418,In_549);
nand U956 (N_956,In_440,In_376);
nand U957 (N_957,In_753,In_882);
nand U958 (N_958,In_737,In_147);
nor U959 (N_959,In_65,In_312);
or U960 (N_960,In_596,In_69);
and U961 (N_961,In_293,In_886);
and U962 (N_962,In_938,In_697);
or U963 (N_963,In_25,In_250);
or U964 (N_964,In_800,In_152);
and U965 (N_965,In_624,In_791);
or U966 (N_966,In_580,In_455);
nor U967 (N_967,In_437,In_833);
nor U968 (N_968,In_637,In_63);
nor U969 (N_969,In_200,In_304);
nand U970 (N_970,In_212,In_576);
nor U971 (N_971,In_405,In_283);
nand U972 (N_972,In_133,In_538);
xnor U973 (N_973,In_989,In_490);
or U974 (N_974,In_834,In_164);
xor U975 (N_975,In_772,In_909);
nor U976 (N_976,In_554,In_313);
and U977 (N_977,In_354,In_134);
xnor U978 (N_978,In_867,In_358);
and U979 (N_979,In_61,In_565);
nor U980 (N_980,In_841,In_344);
or U981 (N_981,In_406,In_34);
or U982 (N_982,In_385,In_773);
nand U983 (N_983,In_369,In_414);
xnor U984 (N_984,In_545,In_160);
and U985 (N_985,In_940,In_0);
and U986 (N_986,In_737,In_367);
nand U987 (N_987,In_492,In_158);
xor U988 (N_988,In_648,In_92);
nand U989 (N_989,In_885,In_339);
nor U990 (N_990,In_691,In_507);
nand U991 (N_991,In_768,In_741);
nand U992 (N_992,In_873,In_559);
or U993 (N_993,In_920,In_683);
or U994 (N_994,In_67,In_685);
and U995 (N_995,In_866,In_411);
nor U996 (N_996,In_576,In_795);
xor U997 (N_997,In_991,In_916);
nand U998 (N_998,In_784,In_444);
or U999 (N_999,In_205,In_972);
or U1000 (N_1000,In_357,In_650);
or U1001 (N_1001,In_883,In_648);
and U1002 (N_1002,In_606,In_367);
xnor U1003 (N_1003,In_95,In_41);
nor U1004 (N_1004,In_920,In_562);
or U1005 (N_1005,In_492,In_682);
xor U1006 (N_1006,In_623,In_651);
nand U1007 (N_1007,In_762,In_868);
xnor U1008 (N_1008,In_396,In_267);
nor U1009 (N_1009,In_473,In_422);
or U1010 (N_1010,In_120,In_766);
xor U1011 (N_1011,In_935,In_379);
nor U1012 (N_1012,In_672,In_362);
nor U1013 (N_1013,In_716,In_776);
nand U1014 (N_1014,In_930,In_722);
or U1015 (N_1015,In_440,In_445);
nor U1016 (N_1016,In_623,In_422);
nand U1017 (N_1017,In_320,In_85);
nor U1018 (N_1018,In_309,In_253);
xnor U1019 (N_1019,In_978,In_529);
xor U1020 (N_1020,In_691,In_127);
nor U1021 (N_1021,In_180,In_966);
or U1022 (N_1022,In_538,In_161);
nand U1023 (N_1023,In_859,In_547);
nor U1024 (N_1024,In_778,In_375);
or U1025 (N_1025,In_345,In_747);
and U1026 (N_1026,In_705,In_457);
nor U1027 (N_1027,In_89,In_901);
nor U1028 (N_1028,In_483,In_257);
nor U1029 (N_1029,In_230,In_585);
nand U1030 (N_1030,In_727,In_962);
xnor U1031 (N_1031,In_394,In_432);
nand U1032 (N_1032,In_881,In_735);
nor U1033 (N_1033,In_174,In_777);
and U1034 (N_1034,In_632,In_514);
nand U1035 (N_1035,In_161,In_25);
nand U1036 (N_1036,In_963,In_840);
nand U1037 (N_1037,In_840,In_260);
xnor U1038 (N_1038,In_308,In_973);
nand U1039 (N_1039,In_281,In_584);
xor U1040 (N_1040,In_714,In_94);
or U1041 (N_1041,In_477,In_529);
or U1042 (N_1042,In_414,In_862);
nor U1043 (N_1043,In_378,In_248);
xnor U1044 (N_1044,In_620,In_372);
nand U1045 (N_1045,In_420,In_113);
or U1046 (N_1046,In_154,In_639);
or U1047 (N_1047,In_877,In_322);
nor U1048 (N_1048,In_475,In_964);
or U1049 (N_1049,In_895,In_592);
and U1050 (N_1050,In_666,In_234);
and U1051 (N_1051,In_475,In_816);
nor U1052 (N_1052,In_630,In_898);
nor U1053 (N_1053,In_10,In_897);
or U1054 (N_1054,In_411,In_236);
nand U1055 (N_1055,In_46,In_393);
nand U1056 (N_1056,In_866,In_50);
nor U1057 (N_1057,In_609,In_565);
or U1058 (N_1058,In_606,In_967);
xor U1059 (N_1059,In_291,In_653);
and U1060 (N_1060,In_808,In_690);
nor U1061 (N_1061,In_372,In_87);
nor U1062 (N_1062,In_455,In_994);
nand U1063 (N_1063,In_998,In_560);
nand U1064 (N_1064,In_605,In_147);
and U1065 (N_1065,In_894,In_961);
nor U1066 (N_1066,In_178,In_808);
nand U1067 (N_1067,In_638,In_457);
or U1068 (N_1068,In_975,In_848);
nor U1069 (N_1069,In_677,In_523);
nand U1070 (N_1070,In_308,In_268);
and U1071 (N_1071,In_140,In_528);
xnor U1072 (N_1072,In_796,In_363);
xnor U1073 (N_1073,In_667,In_597);
and U1074 (N_1074,In_266,In_18);
and U1075 (N_1075,In_978,In_889);
nand U1076 (N_1076,In_832,In_980);
nand U1077 (N_1077,In_706,In_456);
or U1078 (N_1078,In_798,In_728);
xor U1079 (N_1079,In_912,In_423);
nand U1080 (N_1080,In_784,In_788);
or U1081 (N_1081,In_753,In_707);
xor U1082 (N_1082,In_54,In_296);
nand U1083 (N_1083,In_982,In_522);
nand U1084 (N_1084,In_984,In_342);
nor U1085 (N_1085,In_237,In_813);
xor U1086 (N_1086,In_488,In_797);
or U1087 (N_1087,In_768,In_682);
or U1088 (N_1088,In_214,In_85);
or U1089 (N_1089,In_972,In_291);
nand U1090 (N_1090,In_97,In_506);
and U1091 (N_1091,In_843,In_717);
nand U1092 (N_1092,In_774,In_180);
nor U1093 (N_1093,In_322,In_633);
or U1094 (N_1094,In_287,In_240);
xnor U1095 (N_1095,In_72,In_266);
nor U1096 (N_1096,In_261,In_325);
nand U1097 (N_1097,In_206,In_984);
xor U1098 (N_1098,In_163,In_958);
nor U1099 (N_1099,In_708,In_229);
or U1100 (N_1100,In_48,In_43);
or U1101 (N_1101,In_86,In_94);
nor U1102 (N_1102,In_101,In_392);
and U1103 (N_1103,In_856,In_838);
nor U1104 (N_1104,In_805,In_734);
and U1105 (N_1105,In_312,In_901);
nor U1106 (N_1106,In_920,In_311);
and U1107 (N_1107,In_536,In_680);
nand U1108 (N_1108,In_415,In_658);
or U1109 (N_1109,In_441,In_796);
or U1110 (N_1110,In_246,In_300);
nor U1111 (N_1111,In_99,In_495);
and U1112 (N_1112,In_956,In_994);
and U1113 (N_1113,In_486,In_337);
xor U1114 (N_1114,In_878,In_362);
and U1115 (N_1115,In_578,In_587);
or U1116 (N_1116,In_390,In_572);
nand U1117 (N_1117,In_383,In_477);
nor U1118 (N_1118,In_746,In_613);
xnor U1119 (N_1119,In_736,In_756);
nor U1120 (N_1120,In_214,In_287);
and U1121 (N_1121,In_305,In_246);
and U1122 (N_1122,In_213,In_653);
or U1123 (N_1123,In_931,In_50);
and U1124 (N_1124,In_530,In_171);
nand U1125 (N_1125,In_308,In_853);
or U1126 (N_1126,In_607,In_620);
or U1127 (N_1127,In_261,In_641);
or U1128 (N_1128,In_66,In_685);
nor U1129 (N_1129,In_206,In_903);
nor U1130 (N_1130,In_378,In_355);
xnor U1131 (N_1131,In_154,In_665);
and U1132 (N_1132,In_152,In_162);
and U1133 (N_1133,In_678,In_603);
xor U1134 (N_1134,In_382,In_232);
and U1135 (N_1135,In_954,In_823);
xnor U1136 (N_1136,In_945,In_76);
xor U1137 (N_1137,In_600,In_687);
nor U1138 (N_1138,In_689,In_124);
or U1139 (N_1139,In_89,In_665);
xor U1140 (N_1140,In_604,In_988);
nand U1141 (N_1141,In_48,In_657);
and U1142 (N_1142,In_909,In_69);
or U1143 (N_1143,In_293,In_635);
xor U1144 (N_1144,In_460,In_453);
nor U1145 (N_1145,In_302,In_384);
and U1146 (N_1146,In_627,In_208);
xor U1147 (N_1147,In_536,In_167);
nand U1148 (N_1148,In_410,In_967);
nor U1149 (N_1149,In_309,In_687);
or U1150 (N_1150,In_682,In_844);
nand U1151 (N_1151,In_611,In_639);
or U1152 (N_1152,In_534,In_732);
nand U1153 (N_1153,In_203,In_15);
nor U1154 (N_1154,In_644,In_749);
xnor U1155 (N_1155,In_101,In_343);
xnor U1156 (N_1156,In_415,In_489);
nand U1157 (N_1157,In_440,In_611);
or U1158 (N_1158,In_619,In_280);
and U1159 (N_1159,In_718,In_483);
nor U1160 (N_1160,In_556,In_340);
nand U1161 (N_1161,In_873,In_333);
or U1162 (N_1162,In_526,In_794);
nor U1163 (N_1163,In_178,In_208);
and U1164 (N_1164,In_937,In_166);
and U1165 (N_1165,In_47,In_698);
or U1166 (N_1166,In_928,In_353);
nor U1167 (N_1167,In_952,In_665);
and U1168 (N_1168,In_827,In_309);
nor U1169 (N_1169,In_990,In_92);
nand U1170 (N_1170,In_281,In_796);
xor U1171 (N_1171,In_432,In_756);
nor U1172 (N_1172,In_987,In_829);
xnor U1173 (N_1173,In_181,In_584);
nand U1174 (N_1174,In_597,In_982);
and U1175 (N_1175,In_461,In_15);
xor U1176 (N_1176,In_53,In_471);
xor U1177 (N_1177,In_291,In_957);
and U1178 (N_1178,In_906,In_716);
nand U1179 (N_1179,In_364,In_529);
and U1180 (N_1180,In_57,In_370);
or U1181 (N_1181,In_487,In_370);
nor U1182 (N_1182,In_779,In_378);
xor U1183 (N_1183,In_464,In_217);
and U1184 (N_1184,In_561,In_684);
nor U1185 (N_1185,In_294,In_609);
nor U1186 (N_1186,In_371,In_211);
nand U1187 (N_1187,In_857,In_527);
nor U1188 (N_1188,In_784,In_225);
xnor U1189 (N_1189,In_446,In_477);
and U1190 (N_1190,In_543,In_769);
and U1191 (N_1191,In_335,In_165);
or U1192 (N_1192,In_566,In_213);
and U1193 (N_1193,In_806,In_427);
or U1194 (N_1194,In_16,In_13);
nor U1195 (N_1195,In_140,In_531);
nand U1196 (N_1196,In_193,In_620);
xnor U1197 (N_1197,In_309,In_998);
and U1198 (N_1198,In_54,In_811);
nand U1199 (N_1199,In_910,In_102);
xnor U1200 (N_1200,In_692,In_298);
nand U1201 (N_1201,In_434,In_983);
nand U1202 (N_1202,In_384,In_43);
xor U1203 (N_1203,In_681,In_932);
and U1204 (N_1204,In_858,In_298);
or U1205 (N_1205,In_170,In_210);
or U1206 (N_1206,In_776,In_780);
nand U1207 (N_1207,In_20,In_605);
and U1208 (N_1208,In_863,In_122);
xor U1209 (N_1209,In_102,In_538);
nand U1210 (N_1210,In_269,In_75);
nor U1211 (N_1211,In_523,In_572);
or U1212 (N_1212,In_797,In_729);
nor U1213 (N_1213,In_22,In_931);
and U1214 (N_1214,In_394,In_202);
and U1215 (N_1215,In_134,In_661);
xnor U1216 (N_1216,In_68,In_295);
xor U1217 (N_1217,In_731,In_908);
nand U1218 (N_1218,In_225,In_496);
nor U1219 (N_1219,In_571,In_18);
and U1220 (N_1220,In_57,In_532);
or U1221 (N_1221,In_782,In_847);
and U1222 (N_1222,In_41,In_994);
or U1223 (N_1223,In_484,In_630);
or U1224 (N_1224,In_552,In_99);
or U1225 (N_1225,In_467,In_153);
nand U1226 (N_1226,In_806,In_492);
nand U1227 (N_1227,In_882,In_38);
or U1228 (N_1228,In_320,In_87);
nand U1229 (N_1229,In_676,In_800);
nand U1230 (N_1230,In_612,In_68);
nor U1231 (N_1231,In_254,In_161);
nor U1232 (N_1232,In_882,In_461);
xor U1233 (N_1233,In_947,In_705);
or U1234 (N_1234,In_607,In_755);
nand U1235 (N_1235,In_861,In_449);
and U1236 (N_1236,In_803,In_392);
and U1237 (N_1237,In_817,In_435);
and U1238 (N_1238,In_246,In_345);
or U1239 (N_1239,In_574,In_244);
xnor U1240 (N_1240,In_273,In_290);
nand U1241 (N_1241,In_101,In_869);
or U1242 (N_1242,In_423,In_845);
or U1243 (N_1243,In_870,In_935);
or U1244 (N_1244,In_735,In_861);
nand U1245 (N_1245,In_218,In_386);
nand U1246 (N_1246,In_490,In_301);
xnor U1247 (N_1247,In_596,In_463);
nor U1248 (N_1248,In_928,In_623);
nand U1249 (N_1249,In_457,In_146);
xnor U1250 (N_1250,In_933,In_645);
xnor U1251 (N_1251,In_51,In_76);
and U1252 (N_1252,In_793,In_559);
nand U1253 (N_1253,In_517,In_634);
xnor U1254 (N_1254,In_170,In_270);
and U1255 (N_1255,In_183,In_933);
or U1256 (N_1256,In_588,In_334);
xor U1257 (N_1257,In_70,In_867);
or U1258 (N_1258,In_717,In_418);
or U1259 (N_1259,In_650,In_400);
and U1260 (N_1260,In_35,In_681);
xor U1261 (N_1261,In_931,In_584);
xor U1262 (N_1262,In_612,In_984);
nor U1263 (N_1263,In_882,In_769);
nand U1264 (N_1264,In_279,In_759);
xnor U1265 (N_1265,In_669,In_847);
nand U1266 (N_1266,In_0,In_716);
and U1267 (N_1267,In_87,In_272);
nand U1268 (N_1268,In_294,In_219);
or U1269 (N_1269,In_951,In_835);
nor U1270 (N_1270,In_544,In_679);
nand U1271 (N_1271,In_929,In_870);
and U1272 (N_1272,In_318,In_320);
nor U1273 (N_1273,In_130,In_291);
xnor U1274 (N_1274,In_690,In_774);
and U1275 (N_1275,In_830,In_944);
nor U1276 (N_1276,In_350,In_944);
and U1277 (N_1277,In_553,In_318);
nand U1278 (N_1278,In_199,In_787);
xor U1279 (N_1279,In_821,In_449);
nand U1280 (N_1280,In_257,In_865);
and U1281 (N_1281,In_941,In_690);
and U1282 (N_1282,In_66,In_419);
and U1283 (N_1283,In_536,In_714);
nor U1284 (N_1284,In_336,In_130);
or U1285 (N_1285,In_319,In_72);
or U1286 (N_1286,In_948,In_918);
xor U1287 (N_1287,In_800,In_623);
and U1288 (N_1288,In_902,In_11);
or U1289 (N_1289,In_731,In_644);
nor U1290 (N_1290,In_307,In_847);
or U1291 (N_1291,In_600,In_438);
xor U1292 (N_1292,In_505,In_400);
or U1293 (N_1293,In_50,In_469);
xor U1294 (N_1294,In_604,In_529);
or U1295 (N_1295,In_204,In_879);
nor U1296 (N_1296,In_205,In_571);
and U1297 (N_1297,In_423,In_273);
or U1298 (N_1298,In_520,In_941);
and U1299 (N_1299,In_151,In_738);
and U1300 (N_1300,In_801,In_529);
and U1301 (N_1301,In_977,In_708);
or U1302 (N_1302,In_354,In_983);
or U1303 (N_1303,In_998,In_677);
xor U1304 (N_1304,In_778,In_556);
and U1305 (N_1305,In_909,In_467);
nand U1306 (N_1306,In_470,In_290);
nand U1307 (N_1307,In_931,In_646);
nand U1308 (N_1308,In_45,In_761);
and U1309 (N_1309,In_967,In_704);
nand U1310 (N_1310,In_741,In_349);
or U1311 (N_1311,In_40,In_891);
or U1312 (N_1312,In_427,In_234);
or U1313 (N_1313,In_963,In_438);
nor U1314 (N_1314,In_777,In_962);
xnor U1315 (N_1315,In_83,In_371);
and U1316 (N_1316,In_393,In_5);
nand U1317 (N_1317,In_174,In_169);
nand U1318 (N_1318,In_939,In_290);
nor U1319 (N_1319,In_638,In_190);
and U1320 (N_1320,In_617,In_196);
xnor U1321 (N_1321,In_458,In_203);
or U1322 (N_1322,In_731,In_720);
xor U1323 (N_1323,In_291,In_91);
nand U1324 (N_1324,In_46,In_501);
and U1325 (N_1325,In_716,In_653);
or U1326 (N_1326,In_83,In_226);
and U1327 (N_1327,In_288,In_21);
nor U1328 (N_1328,In_942,In_610);
nor U1329 (N_1329,In_1,In_545);
or U1330 (N_1330,In_345,In_972);
xor U1331 (N_1331,In_340,In_111);
xor U1332 (N_1332,In_705,In_658);
xor U1333 (N_1333,In_400,In_718);
and U1334 (N_1334,In_788,In_133);
nand U1335 (N_1335,In_958,In_769);
or U1336 (N_1336,In_662,In_74);
xnor U1337 (N_1337,In_843,In_267);
nand U1338 (N_1338,In_495,In_339);
or U1339 (N_1339,In_4,In_191);
xor U1340 (N_1340,In_368,In_118);
nor U1341 (N_1341,In_709,In_587);
nand U1342 (N_1342,In_856,In_691);
or U1343 (N_1343,In_409,In_988);
nand U1344 (N_1344,In_266,In_368);
xor U1345 (N_1345,In_21,In_159);
xnor U1346 (N_1346,In_852,In_355);
xnor U1347 (N_1347,In_184,In_791);
or U1348 (N_1348,In_214,In_258);
or U1349 (N_1349,In_582,In_47);
nand U1350 (N_1350,In_738,In_163);
and U1351 (N_1351,In_75,In_961);
or U1352 (N_1352,In_522,In_805);
and U1353 (N_1353,In_792,In_237);
or U1354 (N_1354,In_272,In_542);
nand U1355 (N_1355,In_19,In_310);
and U1356 (N_1356,In_911,In_995);
xor U1357 (N_1357,In_357,In_252);
or U1358 (N_1358,In_47,In_955);
and U1359 (N_1359,In_60,In_450);
and U1360 (N_1360,In_892,In_575);
xnor U1361 (N_1361,In_498,In_346);
nor U1362 (N_1362,In_189,In_628);
xnor U1363 (N_1363,In_816,In_926);
nand U1364 (N_1364,In_180,In_612);
or U1365 (N_1365,In_67,In_751);
and U1366 (N_1366,In_656,In_710);
nor U1367 (N_1367,In_545,In_113);
or U1368 (N_1368,In_609,In_985);
nand U1369 (N_1369,In_626,In_427);
xor U1370 (N_1370,In_513,In_359);
and U1371 (N_1371,In_315,In_247);
and U1372 (N_1372,In_242,In_817);
or U1373 (N_1373,In_812,In_976);
nand U1374 (N_1374,In_551,In_577);
or U1375 (N_1375,In_631,In_446);
nand U1376 (N_1376,In_901,In_94);
xor U1377 (N_1377,In_858,In_287);
nor U1378 (N_1378,In_318,In_613);
or U1379 (N_1379,In_111,In_636);
xor U1380 (N_1380,In_605,In_679);
and U1381 (N_1381,In_291,In_297);
nor U1382 (N_1382,In_23,In_946);
nor U1383 (N_1383,In_450,In_773);
nand U1384 (N_1384,In_735,In_319);
nand U1385 (N_1385,In_668,In_712);
or U1386 (N_1386,In_774,In_175);
and U1387 (N_1387,In_208,In_147);
and U1388 (N_1388,In_248,In_730);
or U1389 (N_1389,In_603,In_595);
xnor U1390 (N_1390,In_422,In_284);
and U1391 (N_1391,In_411,In_418);
or U1392 (N_1392,In_664,In_337);
nor U1393 (N_1393,In_453,In_689);
nand U1394 (N_1394,In_962,In_143);
or U1395 (N_1395,In_819,In_273);
or U1396 (N_1396,In_221,In_545);
and U1397 (N_1397,In_594,In_491);
xnor U1398 (N_1398,In_210,In_587);
and U1399 (N_1399,In_878,In_786);
xor U1400 (N_1400,In_227,In_538);
or U1401 (N_1401,In_736,In_944);
and U1402 (N_1402,In_386,In_224);
or U1403 (N_1403,In_849,In_363);
or U1404 (N_1404,In_744,In_809);
or U1405 (N_1405,In_242,In_64);
xor U1406 (N_1406,In_539,In_723);
and U1407 (N_1407,In_937,In_439);
and U1408 (N_1408,In_16,In_786);
xnor U1409 (N_1409,In_381,In_556);
nand U1410 (N_1410,In_719,In_484);
and U1411 (N_1411,In_656,In_536);
nand U1412 (N_1412,In_165,In_138);
or U1413 (N_1413,In_808,In_38);
or U1414 (N_1414,In_386,In_873);
nand U1415 (N_1415,In_843,In_17);
nand U1416 (N_1416,In_366,In_465);
nand U1417 (N_1417,In_114,In_190);
and U1418 (N_1418,In_627,In_399);
or U1419 (N_1419,In_169,In_585);
nand U1420 (N_1420,In_458,In_740);
nor U1421 (N_1421,In_979,In_179);
nor U1422 (N_1422,In_728,In_749);
nor U1423 (N_1423,In_314,In_98);
nand U1424 (N_1424,In_457,In_674);
nand U1425 (N_1425,In_710,In_102);
xor U1426 (N_1426,In_902,In_908);
and U1427 (N_1427,In_332,In_262);
nand U1428 (N_1428,In_292,In_945);
or U1429 (N_1429,In_699,In_909);
xnor U1430 (N_1430,In_800,In_969);
or U1431 (N_1431,In_259,In_664);
nor U1432 (N_1432,In_323,In_78);
nand U1433 (N_1433,In_64,In_810);
or U1434 (N_1434,In_283,In_13);
nor U1435 (N_1435,In_468,In_79);
or U1436 (N_1436,In_600,In_737);
or U1437 (N_1437,In_827,In_412);
nor U1438 (N_1438,In_614,In_192);
xnor U1439 (N_1439,In_25,In_413);
nor U1440 (N_1440,In_103,In_283);
nor U1441 (N_1441,In_360,In_204);
and U1442 (N_1442,In_367,In_346);
nor U1443 (N_1443,In_208,In_720);
nor U1444 (N_1444,In_501,In_632);
or U1445 (N_1445,In_554,In_128);
xor U1446 (N_1446,In_342,In_180);
or U1447 (N_1447,In_966,In_337);
nand U1448 (N_1448,In_503,In_64);
nand U1449 (N_1449,In_655,In_731);
and U1450 (N_1450,In_535,In_717);
or U1451 (N_1451,In_362,In_674);
nand U1452 (N_1452,In_418,In_435);
xor U1453 (N_1453,In_905,In_374);
and U1454 (N_1454,In_818,In_340);
xor U1455 (N_1455,In_597,In_914);
and U1456 (N_1456,In_921,In_937);
xor U1457 (N_1457,In_586,In_13);
xor U1458 (N_1458,In_682,In_872);
nand U1459 (N_1459,In_166,In_760);
and U1460 (N_1460,In_236,In_896);
or U1461 (N_1461,In_469,In_486);
xnor U1462 (N_1462,In_652,In_398);
xor U1463 (N_1463,In_168,In_420);
nand U1464 (N_1464,In_157,In_806);
xor U1465 (N_1465,In_665,In_392);
xor U1466 (N_1466,In_520,In_213);
xnor U1467 (N_1467,In_570,In_972);
nand U1468 (N_1468,In_224,In_586);
or U1469 (N_1469,In_377,In_713);
or U1470 (N_1470,In_694,In_941);
nor U1471 (N_1471,In_525,In_370);
nand U1472 (N_1472,In_70,In_793);
nand U1473 (N_1473,In_886,In_429);
and U1474 (N_1474,In_139,In_875);
xnor U1475 (N_1475,In_952,In_138);
or U1476 (N_1476,In_747,In_471);
and U1477 (N_1477,In_491,In_331);
xor U1478 (N_1478,In_559,In_652);
nor U1479 (N_1479,In_358,In_844);
and U1480 (N_1480,In_38,In_684);
and U1481 (N_1481,In_108,In_213);
nor U1482 (N_1482,In_778,In_381);
and U1483 (N_1483,In_768,In_200);
or U1484 (N_1484,In_257,In_924);
or U1485 (N_1485,In_939,In_659);
and U1486 (N_1486,In_270,In_107);
or U1487 (N_1487,In_527,In_716);
nand U1488 (N_1488,In_363,In_791);
or U1489 (N_1489,In_56,In_779);
or U1490 (N_1490,In_936,In_123);
or U1491 (N_1491,In_846,In_374);
and U1492 (N_1492,In_785,In_929);
nor U1493 (N_1493,In_138,In_241);
or U1494 (N_1494,In_470,In_802);
or U1495 (N_1495,In_93,In_478);
nor U1496 (N_1496,In_457,In_511);
nand U1497 (N_1497,In_244,In_635);
or U1498 (N_1498,In_886,In_583);
nor U1499 (N_1499,In_746,In_342);
xnor U1500 (N_1500,In_449,In_675);
nor U1501 (N_1501,In_783,In_931);
nand U1502 (N_1502,In_29,In_304);
or U1503 (N_1503,In_964,In_147);
xnor U1504 (N_1504,In_656,In_693);
nor U1505 (N_1505,In_977,In_671);
or U1506 (N_1506,In_390,In_775);
xnor U1507 (N_1507,In_79,In_193);
nand U1508 (N_1508,In_784,In_800);
nand U1509 (N_1509,In_398,In_32);
and U1510 (N_1510,In_780,In_619);
nand U1511 (N_1511,In_95,In_586);
nand U1512 (N_1512,In_835,In_899);
nor U1513 (N_1513,In_9,In_901);
or U1514 (N_1514,In_450,In_516);
nand U1515 (N_1515,In_633,In_924);
xor U1516 (N_1516,In_850,In_641);
and U1517 (N_1517,In_141,In_916);
or U1518 (N_1518,In_680,In_177);
or U1519 (N_1519,In_287,In_636);
nand U1520 (N_1520,In_774,In_833);
nand U1521 (N_1521,In_17,In_478);
and U1522 (N_1522,In_321,In_277);
xnor U1523 (N_1523,In_126,In_454);
nand U1524 (N_1524,In_470,In_601);
and U1525 (N_1525,In_232,In_357);
xor U1526 (N_1526,In_495,In_733);
xor U1527 (N_1527,In_530,In_124);
or U1528 (N_1528,In_468,In_954);
or U1529 (N_1529,In_317,In_417);
nor U1530 (N_1530,In_37,In_711);
or U1531 (N_1531,In_59,In_907);
and U1532 (N_1532,In_489,In_661);
and U1533 (N_1533,In_21,In_738);
nand U1534 (N_1534,In_116,In_866);
or U1535 (N_1535,In_963,In_390);
nand U1536 (N_1536,In_261,In_905);
and U1537 (N_1537,In_5,In_130);
nor U1538 (N_1538,In_411,In_406);
and U1539 (N_1539,In_215,In_916);
nor U1540 (N_1540,In_115,In_574);
xor U1541 (N_1541,In_165,In_815);
nor U1542 (N_1542,In_595,In_752);
nor U1543 (N_1543,In_336,In_972);
nor U1544 (N_1544,In_506,In_844);
or U1545 (N_1545,In_787,In_284);
nand U1546 (N_1546,In_31,In_633);
nand U1547 (N_1547,In_311,In_150);
nor U1548 (N_1548,In_788,In_364);
nand U1549 (N_1549,In_413,In_304);
nor U1550 (N_1550,In_423,In_121);
or U1551 (N_1551,In_867,In_239);
nand U1552 (N_1552,In_271,In_221);
nor U1553 (N_1553,In_312,In_946);
or U1554 (N_1554,In_631,In_692);
xnor U1555 (N_1555,In_997,In_25);
and U1556 (N_1556,In_961,In_499);
nand U1557 (N_1557,In_69,In_964);
or U1558 (N_1558,In_960,In_736);
nor U1559 (N_1559,In_379,In_127);
or U1560 (N_1560,In_781,In_43);
and U1561 (N_1561,In_802,In_655);
nor U1562 (N_1562,In_972,In_896);
nand U1563 (N_1563,In_475,In_623);
nand U1564 (N_1564,In_582,In_636);
nor U1565 (N_1565,In_951,In_686);
or U1566 (N_1566,In_175,In_856);
or U1567 (N_1567,In_731,In_537);
and U1568 (N_1568,In_901,In_799);
nor U1569 (N_1569,In_629,In_459);
xor U1570 (N_1570,In_264,In_523);
nand U1571 (N_1571,In_114,In_830);
xor U1572 (N_1572,In_872,In_71);
nand U1573 (N_1573,In_687,In_487);
or U1574 (N_1574,In_505,In_204);
nor U1575 (N_1575,In_724,In_345);
or U1576 (N_1576,In_927,In_519);
and U1577 (N_1577,In_515,In_644);
nand U1578 (N_1578,In_77,In_686);
xnor U1579 (N_1579,In_839,In_208);
or U1580 (N_1580,In_429,In_507);
nor U1581 (N_1581,In_413,In_0);
nor U1582 (N_1582,In_202,In_288);
and U1583 (N_1583,In_782,In_285);
or U1584 (N_1584,In_759,In_737);
nand U1585 (N_1585,In_415,In_794);
xor U1586 (N_1586,In_201,In_365);
or U1587 (N_1587,In_797,In_1);
xnor U1588 (N_1588,In_313,In_928);
nor U1589 (N_1589,In_846,In_155);
nand U1590 (N_1590,In_982,In_149);
and U1591 (N_1591,In_679,In_379);
or U1592 (N_1592,In_530,In_616);
or U1593 (N_1593,In_861,In_218);
nand U1594 (N_1594,In_834,In_436);
xor U1595 (N_1595,In_449,In_44);
and U1596 (N_1596,In_523,In_985);
and U1597 (N_1597,In_191,In_66);
nand U1598 (N_1598,In_83,In_623);
or U1599 (N_1599,In_170,In_540);
and U1600 (N_1600,In_527,In_783);
and U1601 (N_1601,In_144,In_275);
and U1602 (N_1602,In_799,In_793);
and U1603 (N_1603,In_722,In_740);
nor U1604 (N_1604,In_306,In_934);
nand U1605 (N_1605,In_251,In_20);
xor U1606 (N_1606,In_800,In_616);
and U1607 (N_1607,In_735,In_843);
xnor U1608 (N_1608,In_835,In_319);
and U1609 (N_1609,In_621,In_140);
nor U1610 (N_1610,In_845,In_227);
and U1611 (N_1611,In_189,In_650);
nand U1612 (N_1612,In_23,In_155);
and U1613 (N_1613,In_226,In_316);
nand U1614 (N_1614,In_493,In_706);
nand U1615 (N_1615,In_806,In_724);
nand U1616 (N_1616,In_465,In_5);
nor U1617 (N_1617,In_438,In_437);
xor U1618 (N_1618,In_957,In_371);
xor U1619 (N_1619,In_487,In_442);
xor U1620 (N_1620,In_550,In_873);
xor U1621 (N_1621,In_538,In_843);
xor U1622 (N_1622,In_972,In_993);
and U1623 (N_1623,In_231,In_534);
or U1624 (N_1624,In_673,In_698);
and U1625 (N_1625,In_387,In_490);
or U1626 (N_1626,In_991,In_49);
nand U1627 (N_1627,In_999,In_525);
or U1628 (N_1628,In_351,In_464);
or U1629 (N_1629,In_275,In_850);
and U1630 (N_1630,In_230,In_688);
and U1631 (N_1631,In_644,In_541);
or U1632 (N_1632,In_871,In_651);
and U1633 (N_1633,In_731,In_981);
or U1634 (N_1634,In_642,In_197);
or U1635 (N_1635,In_412,In_582);
xor U1636 (N_1636,In_148,In_290);
nand U1637 (N_1637,In_249,In_126);
xnor U1638 (N_1638,In_724,In_404);
and U1639 (N_1639,In_877,In_718);
nand U1640 (N_1640,In_431,In_718);
or U1641 (N_1641,In_546,In_991);
nand U1642 (N_1642,In_530,In_10);
xor U1643 (N_1643,In_926,In_461);
or U1644 (N_1644,In_760,In_399);
nand U1645 (N_1645,In_693,In_608);
nor U1646 (N_1646,In_105,In_760);
nor U1647 (N_1647,In_217,In_768);
nand U1648 (N_1648,In_497,In_58);
xor U1649 (N_1649,In_851,In_212);
nand U1650 (N_1650,In_973,In_545);
xor U1651 (N_1651,In_388,In_401);
nor U1652 (N_1652,In_87,In_427);
xnor U1653 (N_1653,In_542,In_181);
nand U1654 (N_1654,In_149,In_638);
nor U1655 (N_1655,In_357,In_598);
or U1656 (N_1656,In_28,In_546);
xor U1657 (N_1657,In_369,In_96);
or U1658 (N_1658,In_600,In_211);
nand U1659 (N_1659,In_177,In_374);
and U1660 (N_1660,In_76,In_767);
nand U1661 (N_1661,In_666,In_907);
and U1662 (N_1662,In_72,In_815);
and U1663 (N_1663,In_333,In_426);
xnor U1664 (N_1664,In_1,In_225);
nor U1665 (N_1665,In_557,In_857);
or U1666 (N_1666,In_519,In_537);
or U1667 (N_1667,In_357,In_953);
or U1668 (N_1668,In_428,In_295);
nand U1669 (N_1669,In_569,In_634);
xnor U1670 (N_1670,In_603,In_786);
nand U1671 (N_1671,In_249,In_600);
or U1672 (N_1672,In_588,In_974);
or U1673 (N_1673,In_680,In_693);
or U1674 (N_1674,In_194,In_829);
and U1675 (N_1675,In_500,In_409);
xor U1676 (N_1676,In_505,In_161);
nand U1677 (N_1677,In_421,In_756);
nor U1678 (N_1678,In_641,In_776);
nand U1679 (N_1679,In_318,In_924);
nor U1680 (N_1680,In_291,In_9);
and U1681 (N_1681,In_611,In_523);
or U1682 (N_1682,In_538,In_497);
xnor U1683 (N_1683,In_460,In_482);
nor U1684 (N_1684,In_879,In_964);
nand U1685 (N_1685,In_976,In_935);
xnor U1686 (N_1686,In_265,In_422);
nor U1687 (N_1687,In_257,In_743);
and U1688 (N_1688,In_479,In_187);
xor U1689 (N_1689,In_155,In_696);
nor U1690 (N_1690,In_832,In_492);
nor U1691 (N_1691,In_929,In_766);
nor U1692 (N_1692,In_165,In_997);
and U1693 (N_1693,In_445,In_854);
or U1694 (N_1694,In_31,In_441);
or U1695 (N_1695,In_913,In_169);
and U1696 (N_1696,In_378,In_412);
nand U1697 (N_1697,In_852,In_142);
nor U1698 (N_1698,In_750,In_716);
xnor U1699 (N_1699,In_93,In_45);
and U1700 (N_1700,In_25,In_618);
nor U1701 (N_1701,In_711,In_80);
xor U1702 (N_1702,In_45,In_506);
nor U1703 (N_1703,In_626,In_447);
nand U1704 (N_1704,In_978,In_25);
nor U1705 (N_1705,In_170,In_357);
or U1706 (N_1706,In_998,In_699);
or U1707 (N_1707,In_782,In_219);
nand U1708 (N_1708,In_138,In_663);
nor U1709 (N_1709,In_525,In_857);
or U1710 (N_1710,In_206,In_777);
nand U1711 (N_1711,In_662,In_979);
and U1712 (N_1712,In_118,In_379);
or U1713 (N_1713,In_288,In_321);
or U1714 (N_1714,In_169,In_602);
xor U1715 (N_1715,In_873,In_468);
nor U1716 (N_1716,In_418,In_180);
xor U1717 (N_1717,In_972,In_940);
nand U1718 (N_1718,In_586,In_26);
xor U1719 (N_1719,In_42,In_744);
or U1720 (N_1720,In_337,In_216);
and U1721 (N_1721,In_698,In_467);
nand U1722 (N_1722,In_39,In_638);
or U1723 (N_1723,In_665,In_902);
or U1724 (N_1724,In_987,In_10);
and U1725 (N_1725,In_852,In_941);
xor U1726 (N_1726,In_823,In_223);
and U1727 (N_1727,In_614,In_823);
nor U1728 (N_1728,In_962,In_838);
nor U1729 (N_1729,In_192,In_832);
or U1730 (N_1730,In_543,In_922);
nor U1731 (N_1731,In_47,In_383);
nor U1732 (N_1732,In_921,In_137);
xnor U1733 (N_1733,In_319,In_538);
and U1734 (N_1734,In_787,In_36);
nor U1735 (N_1735,In_73,In_25);
and U1736 (N_1736,In_638,In_283);
xnor U1737 (N_1737,In_759,In_848);
xor U1738 (N_1738,In_766,In_34);
nand U1739 (N_1739,In_69,In_846);
nand U1740 (N_1740,In_456,In_976);
or U1741 (N_1741,In_528,In_414);
nand U1742 (N_1742,In_513,In_552);
nand U1743 (N_1743,In_476,In_10);
xor U1744 (N_1744,In_333,In_95);
nor U1745 (N_1745,In_93,In_647);
and U1746 (N_1746,In_880,In_403);
xnor U1747 (N_1747,In_460,In_671);
nand U1748 (N_1748,In_884,In_671);
and U1749 (N_1749,In_284,In_625);
nand U1750 (N_1750,In_945,In_371);
or U1751 (N_1751,In_594,In_776);
nand U1752 (N_1752,In_114,In_571);
and U1753 (N_1753,In_702,In_553);
or U1754 (N_1754,In_714,In_519);
xor U1755 (N_1755,In_104,In_117);
xnor U1756 (N_1756,In_108,In_857);
xor U1757 (N_1757,In_778,In_524);
nor U1758 (N_1758,In_445,In_996);
nor U1759 (N_1759,In_788,In_83);
nor U1760 (N_1760,In_479,In_803);
and U1761 (N_1761,In_219,In_691);
nor U1762 (N_1762,In_234,In_15);
nand U1763 (N_1763,In_180,In_843);
or U1764 (N_1764,In_694,In_56);
xnor U1765 (N_1765,In_239,In_544);
or U1766 (N_1766,In_789,In_891);
nand U1767 (N_1767,In_351,In_769);
and U1768 (N_1768,In_152,In_852);
and U1769 (N_1769,In_464,In_297);
xnor U1770 (N_1770,In_535,In_864);
nor U1771 (N_1771,In_494,In_72);
nand U1772 (N_1772,In_729,In_207);
xor U1773 (N_1773,In_999,In_821);
nand U1774 (N_1774,In_347,In_263);
and U1775 (N_1775,In_269,In_339);
xor U1776 (N_1776,In_447,In_121);
nor U1777 (N_1777,In_134,In_903);
nand U1778 (N_1778,In_941,In_440);
and U1779 (N_1779,In_771,In_763);
nand U1780 (N_1780,In_512,In_104);
nor U1781 (N_1781,In_783,In_471);
xnor U1782 (N_1782,In_151,In_880);
nand U1783 (N_1783,In_609,In_453);
and U1784 (N_1784,In_343,In_453);
nand U1785 (N_1785,In_118,In_538);
and U1786 (N_1786,In_793,In_271);
xor U1787 (N_1787,In_352,In_743);
nand U1788 (N_1788,In_415,In_25);
xor U1789 (N_1789,In_641,In_789);
and U1790 (N_1790,In_566,In_637);
nand U1791 (N_1791,In_117,In_979);
nor U1792 (N_1792,In_319,In_151);
and U1793 (N_1793,In_81,In_758);
nor U1794 (N_1794,In_76,In_649);
xor U1795 (N_1795,In_358,In_363);
nand U1796 (N_1796,In_210,In_24);
and U1797 (N_1797,In_182,In_846);
nand U1798 (N_1798,In_17,In_171);
nor U1799 (N_1799,In_515,In_698);
and U1800 (N_1800,In_284,In_85);
and U1801 (N_1801,In_477,In_848);
or U1802 (N_1802,In_436,In_403);
or U1803 (N_1803,In_346,In_351);
nor U1804 (N_1804,In_758,In_39);
and U1805 (N_1805,In_814,In_736);
nor U1806 (N_1806,In_836,In_138);
xnor U1807 (N_1807,In_439,In_690);
or U1808 (N_1808,In_816,In_733);
nor U1809 (N_1809,In_57,In_268);
and U1810 (N_1810,In_975,In_67);
or U1811 (N_1811,In_483,In_207);
or U1812 (N_1812,In_22,In_240);
xor U1813 (N_1813,In_225,In_890);
xnor U1814 (N_1814,In_829,In_977);
nor U1815 (N_1815,In_641,In_90);
xor U1816 (N_1816,In_434,In_147);
and U1817 (N_1817,In_482,In_347);
nand U1818 (N_1818,In_145,In_629);
xnor U1819 (N_1819,In_533,In_466);
nor U1820 (N_1820,In_10,In_106);
xor U1821 (N_1821,In_908,In_278);
nor U1822 (N_1822,In_837,In_317);
and U1823 (N_1823,In_126,In_803);
and U1824 (N_1824,In_202,In_333);
nand U1825 (N_1825,In_887,In_881);
nor U1826 (N_1826,In_483,In_10);
or U1827 (N_1827,In_621,In_886);
and U1828 (N_1828,In_421,In_138);
nand U1829 (N_1829,In_811,In_140);
xnor U1830 (N_1830,In_528,In_117);
nor U1831 (N_1831,In_386,In_120);
or U1832 (N_1832,In_356,In_832);
and U1833 (N_1833,In_714,In_756);
and U1834 (N_1834,In_397,In_169);
nand U1835 (N_1835,In_562,In_305);
and U1836 (N_1836,In_704,In_900);
or U1837 (N_1837,In_558,In_397);
nor U1838 (N_1838,In_225,In_462);
nand U1839 (N_1839,In_764,In_287);
nor U1840 (N_1840,In_428,In_595);
nand U1841 (N_1841,In_272,In_941);
nor U1842 (N_1842,In_556,In_787);
xnor U1843 (N_1843,In_687,In_870);
or U1844 (N_1844,In_71,In_851);
and U1845 (N_1845,In_804,In_415);
or U1846 (N_1846,In_698,In_49);
or U1847 (N_1847,In_403,In_348);
or U1848 (N_1848,In_937,In_202);
xor U1849 (N_1849,In_645,In_78);
and U1850 (N_1850,In_301,In_331);
xnor U1851 (N_1851,In_688,In_96);
and U1852 (N_1852,In_424,In_239);
nand U1853 (N_1853,In_507,In_127);
nand U1854 (N_1854,In_700,In_463);
or U1855 (N_1855,In_863,In_906);
xor U1856 (N_1856,In_850,In_168);
and U1857 (N_1857,In_335,In_551);
nor U1858 (N_1858,In_658,In_830);
nor U1859 (N_1859,In_71,In_149);
and U1860 (N_1860,In_255,In_923);
nand U1861 (N_1861,In_697,In_979);
and U1862 (N_1862,In_458,In_739);
or U1863 (N_1863,In_698,In_73);
nand U1864 (N_1864,In_521,In_865);
and U1865 (N_1865,In_176,In_848);
nand U1866 (N_1866,In_279,In_74);
nand U1867 (N_1867,In_885,In_234);
nor U1868 (N_1868,In_894,In_833);
xnor U1869 (N_1869,In_904,In_908);
nor U1870 (N_1870,In_161,In_264);
and U1871 (N_1871,In_590,In_235);
xnor U1872 (N_1872,In_503,In_224);
or U1873 (N_1873,In_842,In_505);
and U1874 (N_1874,In_54,In_677);
nor U1875 (N_1875,In_790,In_919);
or U1876 (N_1876,In_172,In_488);
or U1877 (N_1877,In_343,In_437);
or U1878 (N_1878,In_895,In_508);
or U1879 (N_1879,In_148,In_435);
nand U1880 (N_1880,In_815,In_293);
nand U1881 (N_1881,In_570,In_876);
nor U1882 (N_1882,In_294,In_62);
xnor U1883 (N_1883,In_133,In_647);
xor U1884 (N_1884,In_990,In_498);
nand U1885 (N_1885,In_615,In_987);
nand U1886 (N_1886,In_948,In_621);
nand U1887 (N_1887,In_105,In_526);
and U1888 (N_1888,In_996,In_760);
and U1889 (N_1889,In_859,In_917);
or U1890 (N_1890,In_634,In_250);
or U1891 (N_1891,In_203,In_409);
and U1892 (N_1892,In_191,In_595);
or U1893 (N_1893,In_67,In_710);
xor U1894 (N_1894,In_92,In_215);
and U1895 (N_1895,In_95,In_622);
nor U1896 (N_1896,In_557,In_979);
nor U1897 (N_1897,In_853,In_468);
or U1898 (N_1898,In_377,In_236);
xnor U1899 (N_1899,In_750,In_547);
xor U1900 (N_1900,In_896,In_339);
or U1901 (N_1901,In_975,In_431);
xnor U1902 (N_1902,In_597,In_615);
and U1903 (N_1903,In_587,In_630);
nand U1904 (N_1904,In_479,In_986);
xor U1905 (N_1905,In_822,In_146);
nor U1906 (N_1906,In_353,In_825);
xnor U1907 (N_1907,In_787,In_807);
nor U1908 (N_1908,In_244,In_540);
xor U1909 (N_1909,In_922,In_962);
xor U1910 (N_1910,In_276,In_561);
nand U1911 (N_1911,In_34,In_647);
nor U1912 (N_1912,In_523,In_58);
or U1913 (N_1913,In_309,In_734);
nand U1914 (N_1914,In_502,In_899);
nand U1915 (N_1915,In_454,In_479);
or U1916 (N_1916,In_937,In_119);
or U1917 (N_1917,In_324,In_331);
xnor U1918 (N_1918,In_927,In_686);
xnor U1919 (N_1919,In_64,In_891);
nand U1920 (N_1920,In_211,In_275);
nor U1921 (N_1921,In_934,In_826);
nand U1922 (N_1922,In_203,In_840);
nor U1923 (N_1923,In_940,In_310);
nor U1924 (N_1924,In_463,In_727);
xor U1925 (N_1925,In_662,In_840);
or U1926 (N_1926,In_652,In_893);
nand U1927 (N_1927,In_716,In_94);
and U1928 (N_1928,In_432,In_3);
xnor U1929 (N_1929,In_636,In_705);
nand U1930 (N_1930,In_893,In_777);
xor U1931 (N_1931,In_365,In_403);
nand U1932 (N_1932,In_124,In_310);
and U1933 (N_1933,In_117,In_655);
xor U1934 (N_1934,In_969,In_802);
xor U1935 (N_1935,In_471,In_139);
nand U1936 (N_1936,In_263,In_729);
or U1937 (N_1937,In_76,In_189);
xor U1938 (N_1938,In_397,In_639);
nand U1939 (N_1939,In_802,In_604);
and U1940 (N_1940,In_621,In_235);
and U1941 (N_1941,In_80,In_200);
or U1942 (N_1942,In_934,In_636);
xor U1943 (N_1943,In_786,In_695);
nor U1944 (N_1944,In_61,In_396);
nand U1945 (N_1945,In_760,In_103);
nand U1946 (N_1946,In_185,In_459);
or U1947 (N_1947,In_483,In_199);
xor U1948 (N_1948,In_686,In_489);
nor U1949 (N_1949,In_257,In_382);
and U1950 (N_1950,In_554,In_58);
nor U1951 (N_1951,In_513,In_374);
xnor U1952 (N_1952,In_60,In_62);
nand U1953 (N_1953,In_703,In_887);
nand U1954 (N_1954,In_752,In_825);
nand U1955 (N_1955,In_826,In_135);
nor U1956 (N_1956,In_254,In_141);
nor U1957 (N_1957,In_142,In_199);
nor U1958 (N_1958,In_716,In_460);
nand U1959 (N_1959,In_424,In_624);
and U1960 (N_1960,In_665,In_612);
nor U1961 (N_1961,In_990,In_688);
and U1962 (N_1962,In_627,In_35);
nor U1963 (N_1963,In_435,In_293);
nor U1964 (N_1964,In_93,In_548);
and U1965 (N_1965,In_576,In_929);
nor U1966 (N_1966,In_51,In_419);
or U1967 (N_1967,In_599,In_473);
and U1968 (N_1968,In_982,In_148);
nand U1969 (N_1969,In_842,In_277);
nand U1970 (N_1970,In_807,In_867);
or U1971 (N_1971,In_413,In_960);
xnor U1972 (N_1972,In_347,In_202);
or U1973 (N_1973,In_34,In_875);
xnor U1974 (N_1974,In_872,In_215);
xnor U1975 (N_1975,In_930,In_355);
and U1976 (N_1976,In_713,In_964);
and U1977 (N_1977,In_765,In_806);
or U1978 (N_1978,In_380,In_308);
nand U1979 (N_1979,In_67,In_153);
xnor U1980 (N_1980,In_202,In_120);
xnor U1981 (N_1981,In_456,In_985);
nor U1982 (N_1982,In_580,In_730);
nor U1983 (N_1983,In_64,In_406);
and U1984 (N_1984,In_359,In_19);
and U1985 (N_1985,In_189,In_230);
nor U1986 (N_1986,In_509,In_844);
xnor U1987 (N_1987,In_5,In_967);
nand U1988 (N_1988,In_894,In_708);
xor U1989 (N_1989,In_849,In_499);
or U1990 (N_1990,In_914,In_416);
nand U1991 (N_1991,In_200,In_494);
nor U1992 (N_1992,In_706,In_46);
nand U1993 (N_1993,In_28,In_623);
xnor U1994 (N_1994,In_339,In_330);
and U1995 (N_1995,In_745,In_417);
nand U1996 (N_1996,In_991,In_205);
or U1997 (N_1997,In_766,In_264);
nor U1998 (N_1998,In_758,In_883);
or U1999 (N_1999,In_976,In_270);
or U2000 (N_2000,N_1666,N_517);
xor U2001 (N_2001,N_506,N_775);
xnor U2002 (N_2002,N_588,N_779);
xor U2003 (N_2003,N_1344,N_397);
nor U2004 (N_2004,N_1038,N_1581);
xnor U2005 (N_2005,N_669,N_185);
nand U2006 (N_2006,N_784,N_1016);
nand U2007 (N_2007,N_974,N_1373);
or U2008 (N_2008,N_194,N_1821);
xor U2009 (N_2009,N_165,N_1175);
nand U2010 (N_2010,N_842,N_412);
nor U2011 (N_2011,N_308,N_1777);
xor U2012 (N_2012,N_248,N_1906);
nor U2013 (N_2013,N_1416,N_660);
and U2014 (N_2014,N_523,N_1300);
or U2015 (N_2015,N_755,N_1315);
or U2016 (N_2016,N_1636,N_664);
nand U2017 (N_2017,N_605,N_613);
nand U2018 (N_2018,N_965,N_1524);
nand U2019 (N_2019,N_320,N_1455);
or U2020 (N_2020,N_35,N_373);
nand U2021 (N_2021,N_1469,N_1705);
xor U2022 (N_2022,N_977,N_57);
or U2023 (N_2023,N_744,N_935);
nor U2024 (N_2024,N_1905,N_887);
or U2025 (N_2025,N_601,N_541);
and U2026 (N_2026,N_1685,N_529);
xnor U2027 (N_2027,N_95,N_1638);
and U2028 (N_2028,N_573,N_1425);
nand U2029 (N_2029,N_1111,N_370);
nand U2030 (N_2030,N_807,N_1348);
xnor U2031 (N_2031,N_1378,N_1163);
xor U2032 (N_2032,N_1372,N_279);
or U2033 (N_2033,N_737,N_69);
or U2034 (N_2034,N_661,N_836);
nor U2035 (N_2035,N_136,N_681);
or U2036 (N_2036,N_1494,N_1883);
and U2037 (N_2037,N_415,N_1311);
nand U2038 (N_2038,N_1971,N_83);
xnor U2039 (N_2039,N_521,N_1245);
xor U2040 (N_2040,N_897,N_1676);
nand U2041 (N_2041,N_983,N_310);
xor U2042 (N_2042,N_1166,N_558);
nor U2043 (N_2043,N_1305,N_98);
and U2044 (N_2044,N_799,N_1789);
xor U2045 (N_2045,N_1030,N_1023);
nor U2046 (N_2046,N_577,N_1648);
xor U2047 (N_2047,N_76,N_111);
xnor U2048 (N_2048,N_1034,N_19);
xor U2049 (N_2049,N_1398,N_1428);
nor U2050 (N_2050,N_1154,N_1626);
nand U2051 (N_2051,N_1439,N_1321);
xor U2052 (N_2052,N_1691,N_543);
and U2053 (N_2053,N_422,N_1800);
xor U2054 (N_2054,N_1095,N_1483);
nor U2055 (N_2055,N_1830,N_1674);
and U2056 (N_2056,N_198,N_774);
and U2057 (N_2057,N_958,N_877);
xor U2058 (N_2058,N_1476,N_1675);
nor U2059 (N_2059,N_137,N_1934);
and U2060 (N_2060,N_270,N_876);
or U2061 (N_2061,N_666,N_1731);
or U2062 (N_2062,N_170,N_611);
nor U2063 (N_2063,N_479,N_1482);
or U2064 (N_2064,N_335,N_466);
and U2065 (N_2065,N_1096,N_742);
nor U2066 (N_2066,N_1249,N_1422);
and U2067 (N_2067,N_74,N_552);
xnor U2068 (N_2068,N_495,N_702);
and U2069 (N_2069,N_1002,N_122);
nor U2070 (N_2070,N_1670,N_222);
nand U2071 (N_2071,N_546,N_731);
nand U2072 (N_2072,N_1955,N_1790);
xor U2073 (N_2073,N_1324,N_1260);
nor U2074 (N_2074,N_336,N_570);
xor U2075 (N_2075,N_1099,N_1639);
and U2076 (N_2076,N_572,N_845);
nand U2077 (N_2077,N_1486,N_1962);
or U2078 (N_2078,N_239,N_369);
nor U2079 (N_2079,N_1823,N_431);
and U2080 (N_2080,N_1155,N_1271);
and U2081 (N_2081,N_579,N_372);
xnor U2082 (N_2082,N_1668,N_1704);
or U2083 (N_2083,N_338,N_690);
nand U2084 (N_2084,N_938,N_1501);
xnor U2085 (N_2085,N_1829,N_1472);
nor U2086 (N_2086,N_113,N_1762);
xnor U2087 (N_2087,N_1263,N_1911);
nor U2088 (N_2088,N_1555,N_1873);
xor U2089 (N_2089,N_1082,N_339);
nand U2090 (N_2090,N_707,N_1185);
xnor U2091 (N_2091,N_1813,N_399);
and U2092 (N_2092,N_578,N_1242);
nand U2093 (N_2093,N_484,N_1902);
nand U2094 (N_2094,N_1990,N_1525);
nand U2095 (N_2095,N_378,N_1778);
and U2096 (N_2096,N_286,N_1839);
and U2097 (N_2097,N_1499,N_853);
nand U2098 (N_2098,N_1760,N_1448);
and U2099 (N_2099,N_1584,N_1203);
or U2100 (N_2100,N_70,N_1144);
and U2101 (N_2101,N_182,N_926);
xor U2102 (N_2102,N_1410,N_1818);
nor U2103 (N_2103,N_1449,N_1815);
nor U2104 (N_2104,N_438,N_251);
xnor U2105 (N_2105,N_49,N_1152);
and U2106 (N_2106,N_1097,N_1963);
xnor U2107 (N_2107,N_655,N_1307);
nor U2108 (N_2108,N_161,N_627);
nand U2109 (N_2109,N_1606,N_1750);
xor U2110 (N_2110,N_1006,N_107);
nor U2111 (N_2111,N_567,N_538);
nor U2112 (N_2112,N_211,N_1037);
nand U2113 (N_2113,N_536,N_991);
or U2114 (N_2114,N_491,N_1631);
nor U2115 (N_2115,N_1115,N_1585);
or U2116 (N_2116,N_1660,N_387);
xor U2117 (N_2117,N_1328,N_1600);
and U2118 (N_2118,N_1804,N_1877);
or U2119 (N_2119,N_1663,N_1366);
or U2120 (N_2120,N_1898,N_1220);
and U2121 (N_2121,N_266,N_409);
or U2122 (N_2122,N_1699,N_1383);
nand U2123 (N_2123,N_1081,N_1050);
nand U2124 (N_2124,N_1914,N_1210);
and U2125 (N_2125,N_777,N_1954);
or U2126 (N_2126,N_1080,N_835);
and U2127 (N_2127,N_1586,N_238);
and U2128 (N_2128,N_1722,N_1644);
xor U2129 (N_2129,N_1947,N_989);
or U2130 (N_2130,N_1618,N_947);
nand U2131 (N_2131,N_1635,N_511);
nand U2132 (N_2132,N_86,N_1332);
xor U2133 (N_2133,N_64,N_1749);
and U2134 (N_2134,N_1664,N_1709);
or U2135 (N_2135,N_944,N_52);
and U2136 (N_2136,N_846,N_647);
xor U2137 (N_2137,N_769,N_1143);
nand U2138 (N_2138,N_1292,N_867);
and U2139 (N_2139,N_1826,N_1733);
or U2140 (N_2140,N_949,N_396);
xnor U2141 (N_2141,N_493,N_1172);
xnor U2142 (N_2142,N_982,N_1506);
or U2143 (N_2143,N_90,N_1884);
xor U2144 (N_2144,N_604,N_250);
or U2145 (N_2145,N_1860,N_130);
xor U2146 (N_2146,N_514,N_528);
and U2147 (N_2147,N_649,N_1473);
and U2148 (N_2148,N_1736,N_1255);
xor U2149 (N_2149,N_1960,N_223);
nor U2150 (N_2150,N_527,N_416);
and U2151 (N_2151,N_1201,N_1682);
and U2152 (N_2152,N_1021,N_740);
nand U2153 (N_2153,N_1768,N_1545);
nor U2154 (N_2154,N_1151,N_89);
nand U2155 (N_2155,N_599,N_448);
nor U2156 (N_2156,N_208,N_1984);
nand U2157 (N_2157,N_104,N_1688);
and U2158 (N_2158,N_946,N_1949);
xnor U2159 (N_2159,N_1858,N_241);
nand U2160 (N_2160,N_1452,N_1417);
and U2161 (N_2161,N_1576,N_395);
or U2162 (N_2162,N_1803,N_856);
nand U2163 (N_2163,N_1619,N_71);
and U2164 (N_2164,N_460,N_614);
or U2165 (N_2165,N_1078,N_1089);
nand U2166 (N_2166,N_1930,N_1248);
or U2167 (N_2167,N_571,N_1156);
or U2168 (N_2168,N_1624,N_1407);
and U2169 (N_2169,N_1544,N_48);
and U2170 (N_2170,N_637,N_39);
nand U2171 (N_2171,N_1693,N_88);
nand U2172 (N_2172,N_1017,N_376);
xor U2173 (N_2173,N_823,N_1230);
nor U2174 (N_2174,N_189,N_1488);
xor U2175 (N_2175,N_1857,N_1132);
xnor U2176 (N_2176,N_621,N_103);
nor U2177 (N_2177,N_1182,N_1217);
or U2178 (N_2178,N_1518,N_1414);
nand U2179 (N_2179,N_942,N_1924);
and U2180 (N_2180,N_47,N_631);
and U2181 (N_2181,N_1293,N_1523);
xnor U2182 (N_2182,N_1267,N_1098);
or U2183 (N_2183,N_1885,N_1401);
xor U2184 (N_2184,N_507,N_1521);
and U2185 (N_2185,N_1411,N_966);
or U2186 (N_2186,N_245,N_1807);
xor U2187 (N_2187,N_406,N_1872);
nand U2188 (N_2188,N_1084,N_252);
nand U2189 (N_2189,N_1827,N_1350);
or U2190 (N_2190,N_1751,N_910);
nor U2191 (N_2191,N_1596,N_1254);
nor U2192 (N_2192,N_157,N_1478);
nor U2193 (N_2193,N_1667,N_948);
and U2194 (N_2194,N_1289,N_765);
nor U2195 (N_2195,N_1967,N_524);
and U2196 (N_2196,N_153,N_1958);
and U2197 (N_2197,N_990,N_228);
xor U2198 (N_2198,N_1948,N_826);
or U2199 (N_2199,N_37,N_886);
or U2200 (N_2200,N_1765,N_1649);
nand U2201 (N_2201,N_334,N_883);
nand U2202 (N_2202,N_287,N_1176);
nand U2203 (N_2203,N_726,N_1568);
nand U2204 (N_2204,N_1920,N_782);
or U2205 (N_2205,N_1308,N_679);
and U2206 (N_2206,N_816,N_1338);
nor U2207 (N_2207,N_4,N_1429);
nand U2208 (N_2208,N_1892,N_1679);
nand U2209 (N_2209,N_1604,N_269);
or U2210 (N_2210,N_1643,N_778);
xor U2211 (N_2211,N_1171,N_1077);
and U2212 (N_2212,N_829,N_1916);
xor U2213 (N_2213,N_1725,N_560);
xor U2214 (N_2214,N_1552,N_1118);
nand U2215 (N_2215,N_872,N_616);
nand U2216 (N_2216,N_12,N_1970);
nand U2217 (N_2217,N_1394,N_1141);
or U2218 (N_2218,N_328,N_1375);
and U2219 (N_2219,N_467,N_358);
and U2220 (N_2220,N_303,N_1784);
nor U2221 (N_2221,N_476,N_1773);
or U2222 (N_2222,N_1150,N_1577);
xnor U2223 (N_2223,N_1240,N_1758);
nor U2224 (N_2224,N_1766,N_20);
nand U2225 (N_2225,N_1167,N_636);
and U2226 (N_2226,N_869,N_1265);
and U2227 (N_2227,N_160,N_317);
and U2228 (N_2228,N_1866,N_1629);
xnor U2229 (N_2229,N_213,N_1579);
xor U2230 (N_2230,N_1500,N_9);
or U2231 (N_2231,N_1899,N_973);
xnor U2232 (N_2232,N_318,N_704);
xor U2233 (N_2233,N_224,N_1162);
nor U2234 (N_2234,N_1381,N_1367);
and U2235 (N_2235,N_1388,N_686);
and U2236 (N_2236,N_367,N_689);
xnor U2237 (N_2237,N_331,N_1262);
or U2238 (N_2238,N_533,N_825);
or U2239 (N_2239,N_327,N_1409);
or U2240 (N_2240,N_821,N_1405);
nor U2241 (N_2241,N_634,N_1437);
or U2242 (N_2242,N_1646,N_246);
and U2243 (N_2243,N_1431,N_321);
nor U2244 (N_2244,N_1932,N_1863);
nor U2245 (N_2245,N_1741,N_968);
xnor U2246 (N_2246,N_1752,N_635);
nand U2247 (N_2247,N_1280,N_1997);
nand U2248 (N_2248,N_184,N_899);
or U2249 (N_2249,N_1622,N_486);
and U2250 (N_2250,N_1029,N_1513);
nor U2251 (N_2251,N_1468,N_1546);
xor U2252 (N_2252,N_473,N_1404);
or U2253 (N_2253,N_173,N_1194);
or U2254 (N_2254,N_53,N_500);
nand U2255 (N_2255,N_805,N_1893);
and U2256 (N_2256,N_1197,N_445);
nand U2257 (N_2257,N_1453,N_1020);
or U2258 (N_2258,N_734,N_554);
and U2259 (N_2259,N_875,N_801);
nand U2260 (N_2260,N_994,N_863);
and U2261 (N_2261,N_1191,N_1218);
or U2262 (N_2262,N_1000,N_1073);
or U2263 (N_2263,N_1047,N_767);
xnor U2264 (N_2264,N_589,N_1811);
nand U2265 (N_2265,N_315,N_404);
and U2266 (N_2266,N_201,N_485);
nor U2267 (N_2267,N_1542,N_1923);
or U2268 (N_2268,N_1462,N_56);
or U2269 (N_2269,N_1767,N_1538);
xor U2270 (N_2270,N_1612,N_437);
xnor U2271 (N_2271,N_293,N_809);
or U2272 (N_2272,N_1052,N_1785);
xor U2273 (N_2273,N_566,N_1320);
nor U2274 (N_2274,N_1285,N_1754);
and U2275 (N_2275,N_1879,N_607);
nor U2276 (N_2276,N_1092,N_1269);
and U2277 (N_2277,N_191,N_216);
xor U2278 (N_2278,N_447,N_1341);
or U2279 (N_2279,N_1213,N_1522);
or U2280 (N_2280,N_1371,N_143);
xnor U2281 (N_2281,N_1620,N_1548);
and U2282 (N_2282,N_261,N_960);
xnor U2283 (N_2283,N_770,N_914);
nor U2284 (N_2284,N_124,N_1816);
nor U2285 (N_2285,N_1198,N_141);
or U2286 (N_2286,N_1805,N_710);
or U2287 (N_2287,N_1445,N_1969);
nand U2288 (N_2288,N_247,N_633);
nand U2289 (N_2289,N_1671,N_1356);
nand U2290 (N_2290,N_1244,N_81);
and U2291 (N_2291,N_1850,N_1972);
or U2292 (N_2292,N_230,N_1756);
xor U2293 (N_2293,N_1687,N_295);
and U2294 (N_2294,N_932,N_706);
xnor U2295 (N_2295,N_1258,N_903);
or U2296 (N_2296,N_954,N_1862);
and U2297 (N_2297,N_1694,N_314);
nand U2298 (N_2298,N_1157,N_1894);
xnor U2299 (N_2299,N_17,N_884);
or U2300 (N_2300,N_892,N_1842);
nand U2301 (N_2301,N_1102,N_42);
and U2302 (N_2302,N_181,N_1537);
nand U2303 (N_2303,N_764,N_144);
and U2304 (N_2304,N_1661,N_273);
nor U2305 (N_2305,N_1284,N_840);
nor U2306 (N_2306,N_1423,N_357);
xnor U2307 (N_2307,N_446,N_351);
xnor U2308 (N_2308,N_909,N_786);
nor U2309 (N_2309,N_243,N_174);
xor U2310 (N_2310,N_1216,N_1008);
xnor U2311 (N_2311,N_981,N_953);
nor U2312 (N_2312,N_67,N_741);
nand U2313 (N_2313,N_596,N_1168);
nand U2314 (N_2314,N_1653,N_597);
nand U2315 (N_2315,N_1065,N_1992);
xor U2316 (N_2316,N_561,N_1946);
and U2317 (N_2317,N_371,N_1540);
nand U2318 (N_2318,N_168,N_544);
or U2319 (N_2319,N_1505,N_898);
nand U2320 (N_2320,N_1226,N_488);
xor U2321 (N_2321,N_377,N_1441);
and U2322 (N_2322,N_508,N_8);
xnor U2323 (N_2323,N_1470,N_1632);
xor U2324 (N_2324,N_407,N_502);
xor U2325 (N_2325,N_1178,N_1359);
or U2326 (N_2326,N_1788,N_615);
or U2327 (N_2327,N_1817,N_691);
nor U2328 (N_2328,N_565,N_30);
nand U2329 (N_2329,N_855,N_1515);
and U2330 (N_2330,N_662,N_400);
nor U2331 (N_2331,N_699,N_1282);
nand U2332 (N_2332,N_641,N_1330);
and U2333 (N_2333,N_383,N_1655);
nor U2334 (N_2334,N_419,N_365);
nand U2335 (N_2335,N_868,N_815);
or U2336 (N_2336,N_975,N_1748);
xnor U2337 (N_2337,N_1945,N_1491);
nand U2338 (N_2338,N_319,N_1786);
nor U2339 (N_2339,N_852,N_232);
nand U2340 (N_2340,N_1306,N_1325);
xnor U2341 (N_2341,N_659,N_1880);
and U2342 (N_2342,N_687,N_1974);
and U2343 (N_2343,N_119,N_648);
and U2344 (N_2344,N_329,N_392);
or U2345 (N_2345,N_811,N_1588);
or U2346 (N_2346,N_393,N_1046);
nand U2347 (N_2347,N_585,N_939);
nor U2348 (N_2348,N_1147,N_1146);
nor U2349 (N_2349,N_894,N_459);
nand U2350 (N_2350,N_715,N_348);
xor U2351 (N_2351,N_1814,N_539);
nor U2352 (N_2352,N_1004,N_1775);
nand U2353 (N_2353,N_429,N_1665);
xnor U2354 (N_2354,N_259,N_1108);
or U2355 (N_2355,N_1454,N_1318);
or U2356 (N_2356,N_1953,N_1937);
xnor U2357 (N_2357,N_275,N_1808);
or U2358 (N_2358,N_1312,N_7);
xor U2359 (N_2359,N_212,N_498);
nor U2360 (N_2360,N_257,N_575);
nor U2361 (N_2361,N_1125,N_758);
and U2362 (N_2362,N_1068,N_941);
nand U2363 (N_2363,N_490,N_792);
nor U2364 (N_2364,N_470,N_1);
or U2365 (N_2365,N_908,N_1412);
or U2366 (N_2366,N_1011,N_1792);
and U2367 (N_2367,N_414,N_234);
or U2368 (N_2368,N_717,N_444);
and U2369 (N_2369,N_1799,N_1519);
nand U2370 (N_2370,N_5,N_644);
or U2371 (N_2371,N_757,N_1497);
nor U2372 (N_2372,N_296,N_23);
and U2373 (N_2373,N_221,N_1735);
xor U2374 (N_2374,N_1692,N_857);
xnor U2375 (N_2375,N_1045,N_432);
or U2376 (N_2376,N_1276,N_425);
or U2377 (N_2377,N_1492,N_1935);
nor U2378 (N_2378,N_1994,N_66);
or U2379 (N_2379,N_1313,N_709);
or U2380 (N_2380,N_1810,N_1559);
xnor U2381 (N_2381,N_878,N_1868);
xor U2382 (N_2382,N_1702,N_1189);
xnor U2383 (N_2383,N_1802,N_763);
and U2384 (N_2384,N_754,N_426);
nand U2385 (N_2385,N_1295,N_749);
nand U2386 (N_2386,N_603,N_209);
and U2387 (N_2387,N_1364,N_766);
xnor U2388 (N_2388,N_1594,N_197);
and U2389 (N_2389,N_1233,N_997);
xor U2390 (N_2390,N_1053,N_790);
nand U2391 (N_2391,N_1901,N_525);
or U2392 (N_2392,N_716,N_1223);
xnor U2393 (N_2393,N_417,N_780);
nor U2394 (N_2394,N_555,N_1076);
nor U2395 (N_2395,N_1243,N_1033);
xnor U2396 (N_2396,N_987,N_1275);
nor U2397 (N_2397,N_984,N_540);
or U2398 (N_2398,N_106,N_683);
and U2399 (N_2399,N_1235,N_1986);
and U2400 (N_2400,N_695,N_772);
or U2401 (N_2401,N_176,N_1496);
nand U2402 (N_2402,N_82,N_1541);
and U2403 (N_2403,N_46,N_1349);
nand U2404 (N_2404,N_1134,N_1067);
nor U2405 (N_2405,N_1798,N_988);
xnor U2406 (N_2406,N_1103,N_326);
or U2407 (N_2407,N_1133,N_537);
or U2408 (N_2408,N_1039,N_360);
nand U2409 (N_2409,N_1058,N_350);
or U2410 (N_2410,N_1959,N_32);
or U2411 (N_2411,N_54,N_1094);
nor U2412 (N_2412,N_421,N_1764);
nor U2413 (N_2413,N_465,N_1621);
and U2414 (N_2414,N_265,N_187);
nand U2415 (N_2415,N_1869,N_1028);
xnor U2416 (N_2416,N_553,N_494);
or U2417 (N_2417,N_264,N_483);
nor U2418 (N_2418,N_1870,N_1979);
xor U2419 (N_2419,N_827,N_2);
or U2420 (N_2420,N_1290,N_1239);
nand U2421 (N_2421,N_557,N_274);
xnor U2422 (N_2422,N_309,N_118);
nor U2423 (N_2423,N_630,N_1031);
and U2424 (N_2424,N_1838,N_674);
nor U2425 (N_2425,N_618,N_1957);
xor U2426 (N_2426,N_1995,N_186);
and U2427 (N_2427,N_1279,N_1086);
or U2428 (N_2428,N_945,N_27);
nor U2429 (N_2429,N_199,N_1981);
xor U2430 (N_2430,N_1467,N_15);
nand U2431 (N_2431,N_458,N_1950);
or U2432 (N_2432,N_1940,N_1927);
nor U2433 (N_2433,N_1801,N_1534);
nand U2434 (N_2434,N_628,N_1461);
and U2435 (N_2435,N_164,N_653);
or U2436 (N_2436,N_1656,N_1149);
nor U2437 (N_2437,N_1558,N_135);
nand U2438 (N_2438,N_1874,N_1630);
and U2439 (N_2439,N_562,N_87);
nor U2440 (N_2440,N_481,N_298);
and U2441 (N_2441,N_1022,N_833);
nand U2442 (N_2442,N_1598,N_272);
nor U2443 (N_2443,N_456,N_1382);
nand U2444 (N_2444,N_405,N_684);
nor U2445 (N_2445,N_1806,N_549);
or U2446 (N_2446,N_1164,N_1343);
nand U2447 (N_2447,N_356,N_1434);
or U2448 (N_2448,N_817,N_1861);
and U2449 (N_2449,N_1673,N_1380);
xnor U2450 (N_2450,N_1983,N_1442);
or U2451 (N_2451,N_240,N_343);
xor U2452 (N_2452,N_1177,N_115);
or U2453 (N_2453,N_1003,N_1420);
or U2454 (N_2454,N_880,N_1895);
and U2455 (N_2455,N_10,N_1651);
nand U2456 (N_2456,N_1836,N_797);
xnor U2457 (N_2457,N_888,N_617);
nand U2458 (N_2458,N_1936,N_885);
and U2459 (N_2459,N_1783,N_860);
xor U2460 (N_2460,N_673,N_955);
nor U2461 (N_2461,N_1683,N_583);
and U2462 (N_2462,N_866,N_1697);
xor U2463 (N_2463,N_1296,N_1456);
nand U2464 (N_2464,N_692,N_1379);
nor U2465 (N_2465,N_1726,N_824);
or U2466 (N_2466,N_1173,N_1993);
or U2467 (N_2467,N_969,N_1977);
nand U2468 (N_2468,N_1591,N_1738);
xor U2469 (N_2469,N_102,N_1319);
or U2470 (N_2470,N_101,N_1221);
xor U2471 (N_2471,N_1677,N_284);
xor U2472 (N_2472,N_505,N_1719);
xor U2473 (N_2473,N_1358,N_1302);
nand U2474 (N_2474,N_548,N_1933);
and U2475 (N_2475,N_1460,N_902);
xnor U2476 (N_2476,N_117,N_1389);
xor U2477 (N_2477,N_1566,N_218);
and U2478 (N_2478,N_1159,N_890);
and U2479 (N_2479,N_463,N_1896);
or U2480 (N_2480,N_1854,N_1557);
xor U2481 (N_2481,N_998,N_891);
nor U2482 (N_2482,N_155,N_455);
nand U2483 (N_2483,N_762,N_688);
xor U2484 (N_2484,N_776,N_1781);
and U2485 (N_2485,N_451,N_1973);
xor U2486 (N_2486,N_671,N_718);
nand U2487 (N_2487,N_1406,N_225);
nand U2488 (N_2488,N_229,N_1527);
nand U2489 (N_2489,N_564,N_25);
nand U2490 (N_2490,N_812,N_970);
xnor U2491 (N_2491,N_912,N_1988);
xnor U2492 (N_2492,N_530,N_1310);
nand U2493 (N_2493,N_236,N_895);
nand U2494 (N_2494,N_1113,N_150);
and U2495 (N_2495,N_1294,N_729);
nand U2496 (N_2496,N_980,N_1878);
nand U2497 (N_2497,N_1931,N_93);
nand U2498 (N_2498,N_1480,N_1309);
nand U2499 (N_2499,N_347,N_1238);
xor U2500 (N_2500,N_676,N_748);
xor U2501 (N_2501,N_1508,N_177);
nor U2502 (N_2502,N_62,N_714);
nand U2503 (N_2503,N_206,N_1304);
nand U2504 (N_2504,N_640,N_1763);
nand U2505 (N_2505,N_1484,N_1794);
xnor U2506 (N_2506,N_169,N_1026);
nor U2507 (N_2507,N_453,N_1384);
nor U2508 (N_2508,N_1721,N_1291);
nor U2509 (N_2509,N_1051,N_1772);
or U2510 (N_2510,N_1186,N_1362);
nor U2511 (N_2511,N_1712,N_1966);
or U2512 (N_2512,N_1912,N_1225);
xor U2513 (N_2513,N_242,N_837);
xnor U2514 (N_2514,N_889,N_1903);
and U2515 (N_2515,N_1317,N_1640);
nand U2516 (N_2516,N_1729,N_1464);
and U2517 (N_2517,N_1528,N_950);
nor U2518 (N_2518,N_323,N_590);
nor U2519 (N_2519,N_482,N_1613);
nand U2520 (N_2520,N_911,N_768);
nand U2521 (N_2521,N_1057,N_962);
xor U2522 (N_2522,N_1710,N_480);
nand U2523 (N_2523,N_1138,N_1261);
and U2524 (N_2524,N_13,N_793);
nand U2525 (N_2525,N_1840,N_645);
nand U2526 (N_2526,N_154,N_1421);
or U2527 (N_2527,N_1129,N_1917);
xnor U2528 (N_2528,N_1283,N_1834);
or U2529 (N_2529,N_1517,N_1723);
xor U2530 (N_2530,N_1530,N_800);
nand U2531 (N_2531,N_1408,N_1014);
xnor U2532 (N_2532,N_1662,N_834);
nand U2533 (N_2533,N_1753,N_1193);
or U2534 (N_2534,N_593,N_1264);
nand U2535 (N_2535,N_1770,N_773);
and U2536 (N_2536,N_667,N_1761);
or U2537 (N_2537,N_297,N_598);
nor U2538 (N_2538,N_1563,N_11);
or U2539 (N_2539,N_1048,N_1871);
nor U2540 (N_2540,N_1553,N_1529);
nor U2541 (N_2541,N_1828,N_475);
or U2542 (N_2542,N_313,N_1510);
xor U2543 (N_2543,N_1451,N_442);
nand U2544 (N_2544,N_1109,N_267);
or U2545 (N_2545,N_307,N_428);
xor U2546 (N_2546,N_1444,N_77);
nand U2547 (N_2547,N_956,N_1659);
or U2548 (N_2548,N_99,N_1700);
or U2549 (N_2549,N_424,N_971);
nand U2550 (N_2550,N_934,N_423);
or U2551 (N_2551,N_788,N_1145);
nor U2552 (N_2552,N_925,N_1180);
nor U2553 (N_2553,N_1610,N_159);
or U2554 (N_2554,N_680,N_283);
xnor U2555 (N_2555,N_848,N_1774);
xor U2556 (N_2556,N_1387,N_854);
nand U2557 (N_2557,N_1390,N_276);
xnor U2558 (N_2558,N_814,N_1299);
xnor U2559 (N_2559,N_1864,N_1686);
nor U2560 (N_2560,N_1650,N_1286);
and U2561 (N_2561,N_1090,N_986);
or U2562 (N_2562,N_1377,N_1246);
xor U2563 (N_2563,N_1287,N_1658);
xor U2564 (N_2564,N_1281,N_1116);
xor U2565 (N_2565,N_720,N_3);
or U2566 (N_2566,N_504,N_31);
and U2567 (N_2567,N_1996,N_1493);
nand U2568 (N_2568,N_292,N_759);
nand U2569 (N_2569,N_411,N_1270);
nor U2570 (N_2570,N_1843,N_1256);
nor U2571 (N_2571,N_1718,N_1695);
and U2572 (N_2572,N_398,N_355);
or U2573 (N_2573,N_1504,N_1139);
nor U2574 (N_2574,N_1915,N_1329);
and U2575 (N_2575,N_859,N_830);
or U2576 (N_2576,N_18,N_97);
xor U2577 (N_2577,N_450,N_1465);
nand U2578 (N_2578,N_1288,N_332);
or U2579 (N_2579,N_1645,N_1855);
or U2580 (N_2580,N_436,N_464);
nor U2581 (N_2581,N_919,N_487);
nand U2582 (N_2582,N_1479,N_736);
and U2583 (N_2583,N_384,N_282);
nand U2584 (N_2584,N_166,N_364);
and U2585 (N_2585,N_606,N_915);
nand U2586 (N_2586,N_864,N_713);
or U2587 (N_2587,N_220,N_324);
nand U2588 (N_2588,N_501,N_1782);
nor U2589 (N_2589,N_1689,N_1049);
and U2590 (N_2590,N_260,N_721);
nor U2591 (N_2591,N_1054,N_359);
nand U2592 (N_2592,N_803,N_497);
or U2593 (N_2593,N_403,N_1849);
nor U2594 (N_2594,N_1567,N_893);
xor U2595 (N_2595,N_1713,N_922);
nand U2596 (N_2596,N_959,N_569);
nand U2597 (N_2597,N_140,N_280);
xnor U2598 (N_2598,N_1104,N_1919);
nand U2599 (N_2599,N_1490,N_874);
and U2600 (N_2600,N_712,N_114);
nand U2601 (N_2601,N_1797,N_1569);
nand U2602 (N_2602,N_1363,N_1212);
nor U2603 (N_2603,N_1474,N_1060);
and U2604 (N_2604,N_291,N_496);
nand U2605 (N_2605,N_531,N_738);
xor U2606 (N_2606,N_1056,N_1812);
nand U2607 (N_2607,N_937,N_810);
xor U2608 (N_2608,N_516,N_1376);
and U2609 (N_2609,N_747,N_1314);
xor U2610 (N_2610,N_1698,N_1922);
or U2611 (N_2611,N_843,N_304);
xnor U2612 (N_2612,N_1183,N_492);
nor U2613 (N_2613,N_1040,N_787);
and U2614 (N_2614,N_1148,N_263);
nand U2615 (N_2615,N_179,N_1273);
or U2616 (N_2616,N_1865,N_1222);
and U2617 (N_2617,N_1897,N_1153);
and U2618 (N_2618,N_26,N_587);
xor U2619 (N_2619,N_513,N_1925);
nand U2620 (N_2620,N_91,N_656);
nand U2621 (N_2621,N_1085,N_1447);
and U2622 (N_2622,N_957,N_1079);
or U2623 (N_2623,N_443,N_1430);
nor U2624 (N_2624,N_936,N_510);
xnor U2625 (N_2625,N_45,N_930);
xnor U2626 (N_2626,N_1392,N_1578);
nand U2627 (N_2627,N_389,N_1368);
or U2628 (N_2628,N_694,N_126);
or U2629 (N_2629,N_563,N_1044);
and U2630 (N_2630,N_1316,N_921);
and U2631 (N_2631,N_1117,N_258);
nand U2632 (N_2632,N_1779,N_535);
xor U2633 (N_2633,N_390,N_591);
nand U2634 (N_2634,N_281,N_1908);
xnor U2635 (N_2635,N_873,N_1214);
nor U2636 (N_2636,N_870,N_379);
nand U2637 (N_2637,N_643,N_1205);
xnor U2638 (N_2638,N_639,N_1195);
or U2639 (N_2639,N_226,N_200);
xnor U2640 (N_2640,N_1202,N_700);
nand U2641 (N_2641,N_518,N_195);
nor U2642 (N_2642,N_80,N_1609);
nand U2643 (N_2643,N_333,N_1965);
and U2644 (N_2644,N_1961,N_586);
and U2645 (N_2645,N_375,N_1204);
nand U2646 (N_2646,N_1776,N_1565);
nand U2647 (N_2647,N_1337,N_24);
or U2648 (N_2648,N_325,N_78);
and U2649 (N_2649,N_730,N_626);
or U2650 (N_2650,N_1386,N_1793);
xor U2651 (N_2651,N_1744,N_1882);
nor U2652 (N_2652,N_1251,N_1824);
nor U2653 (N_2653,N_1019,N_1769);
xnor U2654 (N_2654,N_1066,N_1137);
or U2655 (N_2655,N_1122,N_916);
or U2656 (N_2656,N_1841,N_1607);
nor U2657 (N_2657,N_1696,N_1140);
xnor U2658 (N_2658,N_1791,N_1743);
and U2659 (N_2659,N_1991,N_1601);
nor U2660 (N_2660,N_996,N_205);
and U2661 (N_2661,N_1707,N_1413);
xor U2662 (N_2662,N_1352,N_1061);
and U2663 (N_2663,N_1323,N_839);
xnor U2664 (N_2664,N_871,N_1900);
or U2665 (N_2665,N_132,N_147);
xnor U2666 (N_2666,N_158,N_1757);
xor U2667 (N_2667,N_1796,N_1457);
nor U2668 (N_2668,N_1876,N_1706);
xor U2669 (N_2669,N_924,N_722);
xor U2670 (N_2670,N_896,N_1070);
xnor U2671 (N_2671,N_632,N_1547);
or U2672 (N_2672,N_745,N_1746);
and U2673 (N_2673,N_440,N_701);
nand U2674 (N_2674,N_861,N_1353);
or U2675 (N_2675,N_1859,N_1603);
nand U2676 (N_2676,N_1432,N_723);
nand U2677 (N_2677,N_756,N_380);
or U2678 (N_2678,N_532,N_262);
or U2679 (N_2679,N_288,N_1370);
nand U2680 (N_2680,N_850,N_1013);
xor U2681 (N_2681,N_1005,N_1711);
and U2682 (N_2682,N_1593,N_985);
and U2683 (N_2683,N_1064,N_1728);
or U2684 (N_2684,N_1227,N_63);
nand U2685 (N_2685,N_256,N_299);
nor U2686 (N_2686,N_1485,N_675);
or U2687 (N_2687,N_820,N_940);
nor U2688 (N_2688,N_1001,N_1351);
or U2689 (N_2689,N_519,N_931);
nor U2690 (N_2690,N_51,N_366);
nor U2691 (N_2691,N_1742,N_1327);
nand U2692 (N_2692,N_844,N_719);
nor U2693 (N_2693,N_305,N_1503);
nand U2694 (N_2694,N_1819,N_1322);
nand U2695 (N_2695,N_1599,N_1554);
nor U2696 (N_2696,N_1142,N_219);
xnor U2697 (N_2697,N_413,N_992);
or U2698 (N_2698,N_1259,N_85);
xor U2699 (N_2699,N_929,N_1495);
and U2700 (N_2700,N_1551,N_512);
nor U2701 (N_2701,N_1374,N_1207);
or U2702 (N_2702,N_1027,N_210);
nor U2703 (N_2703,N_255,N_1652);
and U2704 (N_2704,N_1978,N_798);
nor U2705 (N_2705,N_584,N_1628);
or U2706 (N_2706,N_1130,N_434);
or U2707 (N_2707,N_271,N_1739);
nor U2708 (N_2708,N_1678,N_808);
and U2709 (N_2709,N_472,N_1574);
nand U2710 (N_2710,N_1331,N_1889);
xnor U2711 (N_2711,N_1043,N_391);
xnor U2712 (N_2712,N_1015,N_1944);
and U2713 (N_2713,N_1419,N_1904);
and U2714 (N_2714,N_522,N_1681);
xnor U2715 (N_2715,N_629,N_1120);
and U2716 (N_2716,N_1397,N_1272);
nand U2717 (N_2717,N_612,N_1393);
nor U2718 (N_2718,N_771,N_668);
nand U2719 (N_2719,N_441,N_60);
nand U2720 (N_2720,N_1268,N_125);
and U2721 (N_2721,N_1184,N_340);
nand U2722 (N_2722,N_1121,N_882);
or U2723 (N_2723,N_193,N_469);
or U2724 (N_2724,N_1266,N_901);
or U2725 (N_2725,N_1999,N_595);
or U2726 (N_2726,N_1277,N_881);
xor U2727 (N_2727,N_907,N_1887);
nor U2728 (N_2728,N_36,N_1589);
or U2729 (N_2729,N_253,N_1642);
and U2730 (N_2730,N_344,N_386);
xnor U2731 (N_2731,N_1234,N_217);
nor U2732 (N_2732,N_374,N_1128);
nor U2733 (N_2733,N_1334,N_1229);
nand U2734 (N_2734,N_698,N_1161);
or U2735 (N_2735,N_685,N_979);
nand U2736 (N_2736,N_1072,N_337);
and U2737 (N_2737,N_1342,N_382);
nand U2738 (N_2738,N_112,N_294);
or U2739 (N_2739,N_733,N_146);
nor U2740 (N_2740,N_94,N_1025);
nor U2741 (N_2741,N_724,N_120);
xor U2742 (N_2742,N_1627,N_277);
or U2743 (N_2743,N_545,N_862);
xor U2744 (N_2744,N_1088,N_568);
nand U2745 (N_2745,N_1907,N_116);
xor U2746 (N_2746,N_1740,N_917);
xor U2747 (N_2747,N_430,N_1787);
xor U2748 (N_2748,N_672,N_1572);
xnor U2749 (N_2749,N_622,N_1055);
nor U2750 (N_2750,N_1009,N_138);
xor U2751 (N_2751,N_1403,N_832);
nand U2752 (N_2752,N_1976,N_1929);
xor U2753 (N_2753,N_818,N_148);
or U2754 (N_2754,N_1365,N_1252);
xor U2755 (N_2755,N_418,N_534);
and U2756 (N_2756,N_1536,N_1165);
or U2757 (N_2757,N_638,N_1637);
or U2758 (N_2758,N_1395,N_1708);
or U2759 (N_2759,N_600,N_1190);
xnor U2760 (N_2760,N_665,N_703);
or U2761 (N_2761,N_993,N_1208);
and U2762 (N_2762,N_1985,N_795);
xor U2763 (N_2763,N_906,N_1587);
xor U2764 (N_2764,N_50,N_1361);
xor U2765 (N_2765,N_1440,N_693);
or U2766 (N_2766,N_1845,N_1507);
xor U2767 (N_2767,N_139,N_1402);
or U2768 (N_2768,N_1059,N_732);
and U2769 (N_2769,N_1759,N_963);
or U2770 (N_2770,N_1035,N_1623);
nor U2771 (N_2771,N_1415,N_41);
nor U2772 (N_2772,N_28,N_1867);
nand U2773 (N_2773,N_1354,N_1975);
nand U2774 (N_2774,N_752,N_828);
nor U2775 (N_2775,N_1580,N_1980);
and U2776 (N_2776,N_1590,N_1888);
nor U2777 (N_2777,N_582,N_1124);
xnor U2778 (N_2778,N_156,N_385);
nor U2779 (N_2779,N_1160,N_789);
or U2780 (N_2780,N_515,N_38);
or U2781 (N_2781,N_967,N_1418);
nor U2782 (N_2782,N_1335,N_708);
nand U2783 (N_2783,N_1093,N_559);
nand U2784 (N_2784,N_1968,N_904);
nand U2785 (N_2785,N_1301,N_1573);
or U2786 (N_2786,N_1583,N_978);
nor U2787 (N_2787,N_1206,N_1041);
xor U2788 (N_2788,N_1570,N_1672);
and U2789 (N_2789,N_1087,N_1347);
xor U2790 (N_2790,N_1123,N_933);
and U2791 (N_2791,N_22,N_918);
and U2792 (N_2792,N_109,N_1875);
xor U2793 (N_2793,N_1012,N_1481);
or U2794 (N_2794,N_1657,N_620);
nor U2795 (N_2795,N_1105,N_300);
nand U2796 (N_2796,N_1851,N_244);
nor U2797 (N_2797,N_452,N_1926);
or U2798 (N_2798,N_1616,N_0);
xnor U2799 (N_2799,N_349,N_1669);
or U2800 (N_2800,N_1236,N_581);
and U2801 (N_2801,N_1755,N_1998);
nor U2802 (N_2802,N_1703,N_1357);
and U2803 (N_2803,N_1237,N_1369);
and U2804 (N_2804,N_410,N_920);
nand U2805 (N_2805,N_152,N_468);
nor U2806 (N_2806,N_1730,N_342);
xor U2807 (N_2807,N_489,N_188);
nand U2808 (N_2808,N_751,N_1188);
nand U2809 (N_2809,N_1556,N_92);
or U2810 (N_2810,N_976,N_237);
xnor U2811 (N_2811,N_625,N_471);
nand U2812 (N_2812,N_905,N_1512);
nand U2813 (N_2813,N_551,N_654);
nor U2814 (N_2814,N_129,N_1114);
nor U2815 (N_2815,N_1532,N_1846);
nand U2816 (N_2816,N_1466,N_73);
xor U2817 (N_2817,N_1170,N_477);
and U2818 (N_2818,N_1427,N_207);
or U2819 (N_2819,N_753,N_1734);
nor U2820 (N_2820,N_1745,N_576);
nand U2821 (N_2821,N_322,N_952);
xor U2822 (N_2822,N_167,N_1918);
or U2823 (N_2823,N_1435,N_227);
or U2824 (N_2824,N_363,N_330);
xor U2825 (N_2825,N_1771,N_1820);
and U2826 (N_2826,N_1340,N_1471);
or U2827 (N_2827,N_806,N_791);
nor U2828 (N_2828,N_362,N_943);
nand U2829 (N_2829,N_1690,N_290);
nor U2830 (N_2830,N_1886,N_1535);
nor U2831 (N_2831,N_100,N_841);
and U2832 (N_2832,N_1475,N_402);
or U2833 (N_2833,N_1582,N_1219);
nand U2834 (N_2834,N_145,N_1100);
xor U2835 (N_2835,N_1450,N_761);
or U2836 (N_2836,N_1253,N_995);
or U2837 (N_2837,N_1634,N_449);
or U2838 (N_2838,N_1119,N_658);
nor U2839 (N_2839,N_1297,N_1433);
or U2840 (N_2840,N_1943,N_1680);
xnor U2841 (N_2841,N_1127,N_204);
nor U2842 (N_2842,N_728,N_1247);
nand U2843 (N_2843,N_1571,N_21);
and U2844 (N_2844,N_1400,N_1516);
xnor U2845 (N_2845,N_1187,N_847);
or U2846 (N_2846,N_1560,N_746);
xor U2847 (N_2847,N_1561,N_1333);
and U2848 (N_2848,N_59,N_1112);
or U2849 (N_2849,N_1071,N_1355);
and U2850 (N_2850,N_196,N_1611);
xnor U2851 (N_2851,N_183,N_1241);
and U2852 (N_2852,N_1032,N_354);
nand U2853 (N_2853,N_478,N_33);
and U2854 (N_2854,N_796,N_1179);
xnor U2855 (N_2855,N_1391,N_1250);
or U2856 (N_2856,N_1641,N_203);
or U2857 (N_2857,N_727,N_394);
and U2858 (N_2858,N_1533,N_1833);
nand U2859 (N_2859,N_785,N_381);
nor U2860 (N_2860,N_79,N_171);
nor U2861 (N_2861,N_1091,N_838);
nor U2862 (N_2862,N_1526,N_1952);
and U2863 (N_2863,N_401,N_1158);
or U2864 (N_2864,N_40,N_289);
nand U2865 (N_2865,N_302,N_1075);
nand U2866 (N_2866,N_163,N_1825);
and U2867 (N_2867,N_61,N_951);
nor U2868 (N_2868,N_108,N_1910);
nand U2869 (N_2869,N_1199,N_192);
xor U2870 (N_2870,N_121,N_110);
nand U2871 (N_2871,N_1617,N_1715);
nor U2872 (N_2872,N_1716,N_439);
nand U2873 (N_2873,N_162,N_1385);
and U2874 (N_2874,N_427,N_306);
nor U2875 (N_2875,N_1549,N_1007);
nor U2876 (N_2876,N_1438,N_663);
nand U2877 (N_2877,N_624,N_1720);
and U2878 (N_2878,N_1531,N_1520);
and U2879 (N_2879,N_1360,N_1326);
or U2880 (N_2880,N_1951,N_913);
xor U2881 (N_2881,N_849,N_678);
nor U2882 (N_2882,N_133,N_231);
nor U2883 (N_2883,N_1831,N_999);
nor U2884 (N_2884,N_652,N_1209);
nor U2885 (N_2885,N_368,N_499);
and U2886 (N_2886,N_1856,N_646);
nand U2887 (N_2887,N_1196,N_341);
nor U2888 (N_2888,N_1228,N_550);
and U2889 (N_2889,N_1200,N_388);
and U2890 (N_2890,N_1832,N_1633);
nand U2891 (N_2891,N_1780,N_190);
xnor U2892 (N_2892,N_1564,N_865);
or U2893 (N_2893,N_642,N_697);
or U2894 (N_2894,N_964,N_750);
nor U2895 (N_2895,N_68,N_1498);
nor U2896 (N_2896,N_149,N_254);
nor U2897 (N_2897,N_1024,N_1837);
nor U2898 (N_2898,N_739,N_1399);
or U2899 (N_2899,N_1336,N_461);
nor U2900 (N_2900,N_1169,N_72);
nor U2901 (N_2901,N_705,N_822);
xor U2902 (N_2902,N_1502,N_1847);
and U2903 (N_2903,N_1224,N_175);
nand U2904 (N_2904,N_1443,N_1458);
or U2905 (N_2905,N_361,N_1110);
and U2906 (N_2906,N_34,N_609);
xnor U2907 (N_2907,N_65,N_285);
xor U2908 (N_2908,N_1608,N_346);
xnor U2909 (N_2909,N_131,N_435);
nand U2910 (N_2910,N_1822,N_84);
or U2911 (N_2911,N_1717,N_711);
or U2912 (N_2912,N_735,N_520);
nand U2913 (N_2913,N_1543,N_1174);
nand U2914 (N_2914,N_58,N_1890);
or U2915 (N_2915,N_1036,N_1956);
xor U2916 (N_2916,N_1181,N_1848);
and U2917 (N_2917,N_1913,N_214);
nand U2918 (N_2918,N_202,N_1562);
xnor U2919 (N_2919,N_819,N_1597);
xor U2920 (N_2920,N_1101,N_1477);
nand U2921 (N_2921,N_1274,N_783);
or U2922 (N_2922,N_900,N_556);
or U2923 (N_2923,N_1852,N_657);
nand U2924 (N_2924,N_928,N_542);
xnor U2925 (N_2925,N_1303,N_1795);
or U2926 (N_2926,N_1921,N_16);
nor U2927 (N_2927,N_127,N_1135);
or U2928 (N_2928,N_420,N_233);
xnor U2929 (N_2929,N_1844,N_1231);
and U2930 (N_2930,N_353,N_1909);
nor U2931 (N_2931,N_1625,N_128);
nand U2932 (N_2932,N_1511,N_608);
nand U2933 (N_2933,N_682,N_1459);
nor U2934 (N_2934,N_1215,N_879);
xnor U2935 (N_2935,N_574,N_1928);
and U2936 (N_2936,N_6,N_1727);
and U2937 (N_2937,N_134,N_1339);
or U2938 (N_2938,N_43,N_142);
xnor U2939 (N_2939,N_96,N_1345);
nor U2940 (N_2940,N_1987,N_1550);
xnor U2941 (N_2941,N_923,N_1592);
nor U2942 (N_2942,N_1069,N_1136);
and U2943 (N_2943,N_312,N_1809);
nor U2944 (N_2944,N_1714,N_1982);
and U2945 (N_2945,N_1942,N_105);
and U2946 (N_2946,N_547,N_592);
nand U2947 (N_2947,N_851,N_1489);
or U2948 (N_2948,N_14,N_151);
nand U2949 (N_2949,N_696,N_1232);
xnor U2950 (N_2950,N_1436,N_602);
nor U2951 (N_2951,N_1446,N_345);
nand U2952 (N_2952,N_454,N_1424);
and U2953 (N_2953,N_1684,N_1881);
nand U2954 (N_2954,N_804,N_1747);
or U2955 (N_2955,N_215,N_610);
or U2956 (N_2956,N_1939,N_813);
or U2957 (N_2957,N_1211,N_457);
nand U2958 (N_2958,N_961,N_1724);
xor U2959 (N_2959,N_619,N_650);
and U2960 (N_2960,N_268,N_760);
nor U2961 (N_2961,N_509,N_1487);
or U2962 (N_2962,N_55,N_858);
nand U2963 (N_2963,N_1396,N_1257);
nand U2964 (N_2964,N_1514,N_1615);
or U2965 (N_2965,N_1509,N_1853);
xor U2966 (N_2966,N_172,N_831);
xor U2967 (N_2967,N_1131,N_1614);
xor U2968 (N_2968,N_1938,N_311);
nand U2969 (N_2969,N_352,N_1192);
nor U2970 (N_2970,N_474,N_249);
nor U2971 (N_2971,N_123,N_1732);
and U2972 (N_2972,N_1605,N_1010);
nor U2973 (N_2973,N_301,N_1426);
or U2974 (N_2974,N_651,N_1989);
or U2975 (N_2975,N_180,N_1835);
xnor U2976 (N_2976,N_433,N_1042);
xnor U2977 (N_2977,N_1298,N_743);
and U2978 (N_2978,N_781,N_1654);
xnor U2979 (N_2979,N_1346,N_1602);
xnor U2980 (N_2980,N_526,N_972);
and U2981 (N_2981,N_1647,N_1964);
and U2982 (N_2982,N_670,N_1074);
nand U2983 (N_2983,N_316,N_235);
or U2984 (N_2984,N_1083,N_794);
and U2985 (N_2985,N_503,N_1126);
or U2986 (N_2986,N_677,N_1278);
and U2987 (N_2987,N_802,N_29);
and U2988 (N_2988,N_1062,N_580);
or U2989 (N_2989,N_1595,N_462);
or U2990 (N_2990,N_1941,N_927);
nand U2991 (N_2991,N_623,N_1701);
xnor U2992 (N_2992,N_408,N_44);
or U2993 (N_2993,N_1107,N_1063);
and U2994 (N_2994,N_278,N_178);
xnor U2995 (N_2995,N_1737,N_1891);
nor U2996 (N_2996,N_1575,N_1539);
xnor U2997 (N_2997,N_1463,N_75);
or U2998 (N_2998,N_1106,N_1018);
nor U2999 (N_2999,N_725,N_594);
and U3000 (N_3000,N_1840,N_1424);
nor U3001 (N_3001,N_1132,N_178);
or U3002 (N_3002,N_1262,N_436);
xnor U3003 (N_3003,N_46,N_1128);
nor U3004 (N_3004,N_1774,N_1383);
or U3005 (N_3005,N_878,N_1264);
and U3006 (N_3006,N_103,N_1275);
nor U3007 (N_3007,N_990,N_1289);
xor U3008 (N_3008,N_643,N_664);
xor U3009 (N_3009,N_1179,N_1333);
nand U3010 (N_3010,N_912,N_1066);
or U3011 (N_3011,N_388,N_200);
and U3012 (N_3012,N_451,N_6);
nand U3013 (N_3013,N_1356,N_1078);
nand U3014 (N_3014,N_1256,N_176);
and U3015 (N_3015,N_1694,N_716);
or U3016 (N_3016,N_1352,N_1997);
nor U3017 (N_3017,N_1793,N_718);
nor U3018 (N_3018,N_1706,N_168);
or U3019 (N_3019,N_1701,N_631);
and U3020 (N_3020,N_1572,N_1884);
and U3021 (N_3021,N_1636,N_1679);
and U3022 (N_3022,N_1354,N_647);
and U3023 (N_3023,N_1612,N_946);
nand U3024 (N_3024,N_397,N_450);
xnor U3025 (N_3025,N_1312,N_1146);
nand U3026 (N_3026,N_1420,N_792);
and U3027 (N_3027,N_1426,N_577);
and U3028 (N_3028,N_1866,N_1491);
xnor U3029 (N_3029,N_1589,N_953);
and U3030 (N_3030,N_1645,N_510);
and U3031 (N_3031,N_457,N_84);
nand U3032 (N_3032,N_893,N_1261);
and U3033 (N_3033,N_1664,N_1276);
nor U3034 (N_3034,N_1618,N_59);
nor U3035 (N_3035,N_113,N_1549);
or U3036 (N_3036,N_1545,N_1536);
nor U3037 (N_3037,N_1675,N_550);
nand U3038 (N_3038,N_394,N_148);
xnor U3039 (N_3039,N_944,N_891);
and U3040 (N_3040,N_132,N_1411);
and U3041 (N_3041,N_1815,N_1349);
nor U3042 (N_3042,N_1697,N_1665);
nor U3043 (N_3043,N_1798,N_1843);
nand U3044 (N_3044,N_1462,N_1956);
or U3045 (N_3045,N_400,N_1063);
and U3046 (N_3046,N_1464,N_183);
and U3047 (N_3047,N_445,N_1272);
xnor U3048 (N_3048,N_590,N_473);
xor U3049 (N_3049,N_709,N_1867);
xnor U3050 (N_3050,N_615,N_123);
xnor U3051 (N_3051,N_1829,N_908);
and U3052 (N_3052,N_1562,N_1997);
and U3053 (N_3053,N_499,N_1572);
xor U3054 (N_3054,N_229,N_1728);
and U3055 (N_3055,N_581,N_1576);
nor U3056 (N_3056,N_1356,N_1299);
nor U3057 (N_3057,N_8,N_539);
and U3058 (N_3058,N_1416,N_937);
or U3059 (N_3059,N_1663,N_737);
xor U3060 (N_3060,N_1328,N_282);
and U3061 (N_3061,N_1058,N_94);
or U3062 (N_3062,N_679,N_543);
xor U3063 (N_3063,N_111,N_337);
and U3064 (N_3064,N_842,N_1317);
nand U3065 (N_3065,N_759,N_493);
nand U3066 (N_3066,N_708,N_1115);
or U3067 (N_3067,N_1575,N_862);
or U3068 (N_3068,N_1596,N_1539);
or U3069 (N_3069,N_1590,N_1794);
nor U3070 (N_3070,N_1502,N_739);
nor U3071 (N_3071,N_1831,N_416);
or U3072 (N_3072,N_685,N_367);
and U3073 (N_3073,N_491,N_660);
nor U3074 (N_3074,N_77,N_1917);
nand U3075 (N_3075,N_775,N_1161);
or U3076 (N_3076,N_145,N_149);
and U3077 (N_3077,N_1911,N_1027);
nand U3078 (N_3078,N_1654,N_1683);
nor U3079 (N_3079,N_1227,N_1818);
xnor U3080 (N_3080,N_993,N_669);
xor U3081 (N_3081,N_799,N_1153);
nand U3082 (N_3082,N_1458,N_713);
or U3083 (N_3083,N_1756,N_267);
nor U3084 (N_3084,N_333,N_681);
xnor U3085 (N_3085,N_1514,N_166);
or U3086 (N_3086,N_1985,N_1484);
or U3087 (N_3087,N_1679,N_1397);
nor U3088 (N_3088,N_911,N_1412);
nor U3089 (N_3089,N_1973,N_147);
or U3090 (N_3090,N_1628,N_1781);
nand U3091 (N_3091,N_1598,N_1047);
nand U3092 (N_3092,N_714,N_1003);
nand U3093 (N_3093,N_1483,N_1925);
nor U3094 (N_3094,N_877,N_1586);
nand U3095 (N_3095,N_67,N_360);
xor U3096 (N_3096,N_501,N_1763);
nor U3097 (N_3097,N_684,N_1461);
nor U3098 (N_3098,N_221,N_782);
nor U3099 (N_3099,N_176,N_350);
or U3100 (N_3100,N_291,N_1168);
xor U3101 (N_3101,N_20,N_1598);
and U3102 (N_3102,N_1053,N_1762);
and U3103 (N_3103,N_374,N_1910);
nor U3104 (N_3104,N_72,N_457);
and U3105 (N_3105,N_1031,N_692);
nor U3106 (N_3106,N_1397,N_758);
nand U3107 (N_3107,N_1894,N_378);
nor U3108 (N_3108,N_1974,N_847);
nor U3109 (N_3109,N_72,N_1852);
or U3110 (N_3110,N_1255,N_332);
xnor U3111 (N_3111,N_1376,N_439);
and U3112 (N_3112,N_1985,N_114);
xnor U3113 (N_3113,N_1760,N_649);
and U3114 (N_3114,N_41,N_1949);
and U3115 (N_3115,N_1013,N_1037);
nor U3116 (N_3116,N_1677,N_1718);
or U3117 (N_3117,N_1145,N_1974);
nand U3118 (N_3118,N_1994,N_1674);
xor U3119 (N_3119,N_259,N_61);
xor U3120 (N_3120,N_204,N_229);
or U3121 (N_3121,N_297,N_1548);
nand U3122 (N_3122,N_272,N_1901);
nand U3123 (N_3123,N_306,N_975);
and U3124 (N_3124,N_410,N_1129);
xnor U3125 (N_3125,N_711,N_121);
and U3126 (N_3126,N_1433,N_1026);
nand U3127 (N_3127,N_1359,N_535);
nor U3128 (N_3128,N_1290,N_514);
nor U3129 (N_3129,N_265,N_1457);
nand U3130 (N_3130,N_592,N_240);
nand U3131 (N_3131,N_99,N_1728);
or U3132 (N_3132,N_135,N_1498);
or U3133 (N_3133,N_609,N_717);
nor U3134 (N_3134,N_32,N_663);
xor U3135 (N_3135,N_61,N_1263);
xor U3136 (N_3136,N_1380,N_1511);
and U3137 (N_3137,N_1183,N_1428);
nand U3138 (N_3138,N_1469,N_1204);
xnor U3139 (N_3139,N_873,N_812);
xnor U3140 (N_3140,N_1258,N_1237);
xor U3141 (N_3141,N_1196,N_925);
and U3142 (N_3142,N_793,N_1751);
xnor U3143 (N_3143,N_1598,N_1972);
nand U3144 (N_3144,N_677,N_955);
or U3145 (N_3145,N_1320,N_154);
and U3146 (N_3146,N_1263,N_564);
nor U3147 (N_3147,N_1258,N_486);
or U3148 (N_3148,N_473,N_349);
nand U3149 (N_3149,N_426,N_1429);
nor U3150 (N_3150,N_1949,N_406);
nand U3151 (N_3151,N_1656,N_991);
or U3152 (N_3152,N_76,N_541);
and U3153 (N_3153,N_1675,N_1058);
nand U3154 (N_3154,N_1789,N_868);
xnor U3155 (N_3155,N_846,N_576);
xor U3156 (N_3156,N_1749,N_201);
nor U3157 (N_3157,N_191,N_450);
nand U3158 (N_3158,N_1359,N_518);
nand U3159 (N_3159,N_564,N_5);
and U3160 (N_3160,N_1930,N_1488);
or U3161 (N_3161,N_1388,N_269);
or U3162 (N_3162,N_41,N_1618);
and U3163 (N_3163,N_158,N_322);
nand U3164 (N_3164,N_705,N_30);
and U3165 (N_3165,N_176,N_487);
nand U3166 (N_3166,N_1627,N_1454);
xnor U3167 (N_3167,N_1225,N_1280);
and U3168 (N_3168,N_651,N_1450);
or U3169 (N_3169,N_1503,N_1720);
and U3170 (N_3170,N_586,N_83);
xor U3171 (N_3171,N_1099,N_907);
and U3172 (N_3172,N_1915,N_1394);
and U3173 (N_3173,N_730,N_1740);
nor U3174 (N_3174,N_1045,N_1095);
and U3175 (N_3175,N_1746,N_652);
and U3176 (N_3176,N_512,N_979);
or U3177 (N_3177,N_662,N_1566);
nand U3178 (N_3178,N_1595,N_1955);
nor U3179 (N_3179,N_445,N_115);
or U3180 (N_3180,N_1251,N_1167);
and U3181 (N_3181,N_1913,N_1127);
and U3182 (N_3182,N_988,N_1791);
xor U3183 (N_3183,N_120,N_698);
nor U3184 (N_3184,N_1508,N_760);
nand U3185 (N_3185,N_1804,N_1651);
nor U3186 (N_3186,N_908,N_1129);
nand U3187 (N_3187,N_341,N_266);
nor U3188 (N_3188,N_1064,N_189);
or U3189 (N_3189,N_51,N_151);
or U3190 (N_3190,N_649,N_157);
or U3191 (N_3191,N_960,N_292);
and U3192 (N_3192,N_1310,N_883);
nand U3193 (N_3193,N_116,N_1428);
nor U3194 (N_3194,N_1960,N_558);
or U3195 (N_3195,N_502,N_1140);
or U3196 (N_3196,N_1195,N_988);
xor U3197 (N_3197,N_1648,N_854);
nor U3198 (N_3198,N_1664,N_1262);
and U3199 (N_3199,N_959,N_1365);
nand U3200 (N_3200,N_774,N_523);
or U3201 (N_3201,N_1228,N_1082);
nand U3202 (N_3202,N_1308,N_972);
or U3203 (N_3203,N_1196,N_1379);
and U3204 (N_3204,N_1002,N_1308);
nor U3205 (N_3205,N_56,N_740);
or U3206 (N_3206,N_71,N_515);
and U3207 (N_3207,N_1262,N_852);
xor U3208 (N_3208,N_134,N_1555);
or U3209 (N_3209,N_1989,N_1362);
and U3210 (N_3210,N_1378,N_1438);
and U3211 (N_3211,N_372,N_297);
xnor U3212 (N_3212,N_1012,N_1071);
nor U3213 (N_3213,N_727,N_288);
nor U3214 (N_3214,N_1329,N_1945);
xor U3215 (N_3215,N_1814,N_1037);
nand U3216 (N_3216,N_1169,N_1905);
nand U3217 (N_3217,N_1202,N_169);
and U3218 (N_3218,N_674,N_220);
and U3219 (N_3219,N_569,N_176);
or U3220 (N_3220,N_1045,N_287);
nand U3221 (N_3221,N_1369,N_247);
xnor U3222 (N_3222,N_1466,N_94);
or U3223 (N_3223,N_122,N_89);
xor U3224 (N_3224,N_756,N_1665);
xnor U3225 (N_3225,N_1098,N_421);
nor U3226 (N_3226,N_227,N_1913);
nand U3227 (N_3227,N_414,N_1481);
xor U3228 (N_3228,N_1913,N_1669);
or U3229 (N_3229,N_1084,N_348);
or U3230 (N_3230,N_1922,N_282);
nand U3231 (N_3231,N_63,N_34);
nor U3232 (N_3232,N_920,N_407);
and U3233 (N_3233,N_705,N_1412);
nand U3234 (N_3234,N_334,N_771);
nand U3235 (N_3235,N_1562,N_71);
nor U3236 (N_3236,N_22,N_1974);
xnor U3237 (N_3237,N_470,N_1681);
nand U3238 (N_3238,N_661,N_133);
nand U3239 (N_3239,N_593,N_98);
and U3240 (N_3240,N_1137,N_991);
nand U3241 (N_3241,N_1999,N_1641);
xor U3242 (N_3242,N_1428,N_1666);
nor U3243 (N_3243,N_616,N_823);
nor U3244 (N_3244,N_1875,N_668);
and U3245 (N_3245,N_138,N_487);
nor U3246 (N_3246,N_829,N_1691);
or U3247 (N_3247,N_1259,N_768);
nand U3248 (N_3248,N_631,N_1082);
xor U3249 (N_3249,N_1206,N_761);
nor U3250 (N_3250,N_904,N_307);
nor U3251 (N_3251,N_8,N_417);
xor U3252 (N_3252,N_921,N_722);
and U3253 (N_3253,N_645,N_1711);
nor U3254 (N_3254,N_2,N_1065);
nand U3255 (N_3255,N_442,N_599);
nor U3256 (N_3256,N_192,N_196);
and U3257 (N_3257,N_498,N_1531);
and U3258 (N_3258,N_783,N_1626);
nor U3259 (N_3259,N_606,N_447);
nand U3260 (N_3260,N_81,N_904);
xor U3261 (N_3261,N_1557,N_905);
nand U3262 (N_3262,N_375,N_743);
nor U3263 (N_3263,N_972,N_1432);
nor U3264 (N_3264,N_1400,N_954);
and U3265 (N_3265,N_997,N_1000);
and U3266 (N_3266,N_792,N_1755);
or U3267 (N_3267,N_856,N_849);
or U3268 (N_3268,N_89,N_182);
nor U3269 (N_3269,N_1902,N_663);
nor U3270 (N_3270,N_318,N_661);
nor U3271 (N_3271,N_24,N_57);
xnor U3272 (N_3272,N_560,N_1849);
nand U3273 (N_3273,N_558,N_1780);
and U3274 (N_3274,N_1610,N_1385);
and U3275 (N_3275,N_889,N_1854);
nor U3276 (N_3276,N_216,N_943);
and U3277 (N_3277,N_1146,N_786);
nand U3278 (N_3278,N_821,N_508);
nor U3279 (N_3279,N_607,N_436);
xnor U3280 (N_3280,N_490,N_33);
nor U3281 (N_3281,N_1247,N_170);
and U3282 (N_3282,N_13,N_1195);
xnor U3283 (N_3283,N_1914,N_853);
and U3284 (N_3284,N_1201,N_270);
or U3285 (N_3285,N_1055,N_761);
and U3286 (N_3286,N_1825,N_1082);
or U3287 (N_3287,N_1919,N_1416);
nand U3288 (N_3288,N_693,N_1913);
nand U3289 (N_3289,N_1112,N_52);
nor U3290 (N_3290,N_757,N_756);
or U3291 (N_3291,N_223,N_977);
and U3292 (N_3292,N_1025,N_40);
xor U3293 (N_3293,N_1782,N_1485);
xnor U3294 (N_3294,N_362,N_998);
and U3295 (N_3295,N_1594,N_590);
or U3296 (N_3296,N_1435,N_1320);
and U3297 (N_3297,N_140,N_1535);
and U3298 (N_3298,N_699,N_977);
xnor U3299 (N_3299,N_34,N_611);
and U3300 (N_3300,N_922,N_333);
and U3301 (N_3301,N_99,N_895);
or U3302 (N_3302,N_1351,N_361);
and U3303 (N_3303,N_1237,N_438);
nor U3304 (N_3304,N_1663,N_1757);
and U3305 (N_3305,N_932,N_1757);
or U3306 (N_3306,N_1398,N_1589);
or U3307 (N_3307,N_166,N_895);
nor U3308 (N_3308,N_1693,N_1074);
nor U3309 (N_3309,N_475,N_322);
and U3310 (N_3310,N_535,N_1242);
xor U3311 (N_3311,N_1941,N_1254);
and U3312 (N_3312,N_314,N_1662);
xor U3313 (N_3313,N_435,N_1233);
nand U3314 (N_3314,N_1857,N_1439);
nor U3315 (N_3315,N_587,N_175);
nor U3316 (N_3316,N_256,N_1037);
and U3317 (N_3317,N_64,N_1252);
nor U3318 (N_3318,N_859,N_1575);
and U3319 (N_3319,N_1913,N_171);
nor U3320 (N_3320,N_1986,N_681);
or U3321 (N_3321,N_211,N_1088);
xor U3322 (N_3322,N_0,N_1861);
nor U3323 (N_3323,N_309,N_1311);
or U3324 (N_3324,N_1977,N_837);
xnor U3325 (N_3325,N_1833,N_1655);
and U3326 (N_3326,N_1050,N_892);
xnor U3327 (N_3327,N_817,N_331);
nor U3328 (N_3328,N_207,N_595);
xor U3329 (N_3329,N_1369,N_1684);
or U3330 (N_3330,N_1343,N_203);
and U3331 (N_3331,N_1763,N_1044);
or U3332 (N_3332,N_931,N_1359);
nand U3333 (N_3333,N_1316,N_356);
and U3334 (N_3334,N_1898,N_132);
xor U3335 (N_3335,N_1200,N_120);
or U3336 (N_3336,N_1085,N_1772);
nor U3337 (N_3337,N_166,N_1047);
or U3338 (N_3338,N_1261,N_1789);
xor U3339 (N_3339,N_1770,N_735);
xnor U3340 (N_3340,N_995,N_143);
nor U3341 (N_3341,N_1727,N_1619);
and U3342 (N_3342,N_965,N_785);
or U3343 (N_3343,N_1550,N_394);
xor U3344 (N_3344,N_831,N_1743);
xnor U3345 (N_3345,N_637,N_398);
or U3346 (N_3346,N_853,N_1539);
and U3347 (N_3347,N_1573,N_1223);
and U3348 (N_3348,N_141,N_833);
nor U3349 (N_3349,N_1029,N_793);
or U3350 (N_3350,N_188,N_1224);
and U3351 (N_3351,N_1879,N_580);
nand U3352 (N_3352,N_472,N_1985);
or U3353 (N_3353,N_132,N_977);
nand U3354 (N_3354,N_354,N_990);
or U3355 (N_3355,N_760,N_993);
nand U3356 (N_3356,N_401,N_1748);
and U3357 (N_3357,N_1515,N_700);
or U3358 (N_3358,N_559,N_482);
or U3359 (N_3359,N_1143,N_1496);
nand U3360 (N_3360,N_609,N_588);
xor U3361 (N_3361,N_1172,N_549);
and U3362 (N_3362,N_1658,N_415);
or U3363 (N_3363,N_1959,N_995);
and U3364 (N_3364,N_1913,N_1678);
nand U3365 (N_3365,N_1141,N_604);
nand U3366 (N_3366,N_1610,N_264);
nor U3367 (N_3367,N_1666,N_634);
and U3368 (N_3368,N_1194,N_243);
and U3369 (N_3369,N_1514,N_1333);
or U3370 (N_3370,N_58,N_1554);
nor U3371 (N_3371,N_26,N_1152);
xnor U3372 (N_3372,N_1790,N_489);
nand U3373 (N_3373,N_524,N_1942);
and U3374 (N_3374,N_139,N_1887);
nor U3375 (N_3375,N_1249,N_10);
nor U3376 (N_3376,N_924,N_632);
xnor U3377 (N_3377,N_371,N_77);
nor U3378 (N_3378,N_1020,N_147);
and U3379 (N_3379,N_865,N_839);
nor U3380 (N_3380,N_776,N_964);
nor U3381 (N_3381,N_1409,N_273);
nand U3382 (N_3382,N_349,N_1865);
and U3383 (N_3383,N_1831,N_452);
or U3384 (N_3384,N_975,N_518);
nor U3385 (N_3385,N_683,N_1908);
nand U3386 (N_3386,N_265,N_1036);
nor U3387 (N_3387,N_701,N_1089);
xor U3388 (N_3388,N_1312,N_1307);
or U3389 (N_3389,N_1259,N_354);
xor U3390 (N_3390,N_229,N_744);
nor U3391 (N_3391,N_1119,N_912);
and U3392 (N_3392,N_24,N_310);
xor U3393 (N_3393,N_814,N_430);
and U3394 (N_3394,N_1387,N_1194);
nand U3395 (N_3395,N_741,N_224);
xor U3396 (N_3396,N_1639,N_707);
xnor U3397 (N_3397,N_1429,N_213);
xor U3398 (N_3398,N_1878,N_1743);
nand U3399 (N_3399,N_1544,N_128);
or U3400 (N_3400,N_1102,N_1105);
xor U3401 (N_3401,N_1138,N_776);
xnor U3402 (N_3402,N_1636,N_1535);
xor U3403 (N_3403,N_1824,N_713);
and U3404 (N_3404,N_938,N_595);
or U3405 (N_3405,N_1126,N_60);
xor U3406 (N_3406,N_539,N_1845);
or U3407 (N_3407,N_567,N_949);
nor U3408 (N_3408,N_667,N_661);
and U3409 (N_3409,N_1889,N_1657);
or U3410 (N_3410,N_484,N_358);
xor U3411 (N_3411,N_952,N_662);
nor U3412 (N_3412,N_899,N_70);
nand U3413 (N_3413,N_1609,N_1312);
and U3414 (N_3414,N_1187,N_1441);
nand U3415 (N_3415,N_874,N_788);
and U3416 (N_3416,N_1242,N_255);
nor U3417 (N_3417,N_541,N_174);
and U3418 (N_3418,N_270,N_1202);
xnor U3419 (N_3419,N_280,N_1815);
or U3420 (N_3420,N_1673,N_1136);
nand U3421 (N_3421,N_1559,N_1460);
and U3422 (N_3422,N_1510,N_187);
nand U3423 (N_3423,N_494,N_1440);
xor U3424 (N_3424,N_203,N_587);
xor U3425 (N_3425,N_1433,N_833);
nand U3426 (N_3426,N_295,N_608);
nand U3427 (N_3427,N_85,N_316);
and U3428 (N_3428,N_1409,N_638);
and U3429 (N_3429,N_91,N_387);
or U3430 (N_3430,N_1571,N_445);
or U3431 (N_3431,N_681,N_804);
nand U3432 (N_3432,N_1860,N_895);
xnor U3433 (N_3433,N_1577,N_737);
or U3434 (N_3434,N_1455,N_718);
nor U3435 (N_3435,N_298,N_492);
or U3436 (N_3436,N_1916,N_1882);
nand U3437 (N_3437,N_776,N_1869);
nand U3438 (N_3438,N_462,N_1502);
or U3439 (N_3439,N_1647,N_172);
and U3440 (N_3440,N_761,N_1950);
nand U3441 (N_3441,N_1495,N_258);
xnor U3442 (N_3442,N_608,N_799);
or U3443 (N_3443,N_115,N_1748);
nor U3444 (N_3444,N_134,N_1968);
xnor U3445 (N_3445,N_1110,N_1843);
or U3446 (N_3446,N_1692,N_1043);
nor U3447 (N_3447,N_1502,N_365);
nor U3448 (N_3448,N_1233,N_709);
xor U3449 (N_3449,N_155,N_967);
and U3450 (N_3450,N_1051,N_1731);
or U3451 (N_3451,N_583,N_27);
nor U3452 (N_3452,N_1580,N_1332);
nand U3453 (N_3453,N_950,N_384);
nand U3454 (N_3454,N_1948,N_1241);
xor U3455 (N_3455,N_887,N_549);
nor U3456 (N_3456,N_1028,N_1683);
or U3457 (N_3457,N_1576,N_841);
or U3458 (N_3458,N_986,N_848);
and U3459 (N_3459,N_1721,N_906);
nor U3460 (N_3460,N_1774,N_1307);
and U3461 (N_3461,N_1807,N_247);
xnor U3462 (N_3462,N_290,N_1521);
xnor U3463 (N_3463,N_720,N_1215);
nor U3464 (N_3464,N_336,N_1647);
nor U3465 (N_3465,N_250,N_644);
nor U3466 (N_3466,N_1781,N_413);
xnor U3467 (N_3467,N_1662,N_1542);
nor U3468 (N_3468,N_485,N_1002);
nand U3469 (N_3469,N_141,N_113);
xor U3470 (N_3470,N_1524,N_762);
and U3471 (N_3471,N_648,N_985);
and U3472 (N_3472,N_880,N_0);
xnor U3473 (N_3473,N_606,N_590);
nand U3474 (N_3474,N_1225,N_1942);
nor U3475 (N_3475,N_175,N_544);
nor U3476 (N_3476,N_1384,N_1779);
or U3477 (N_3477,N_1506,N_555);
and U3478 (N_3478,N_614,N_1596);
and U3479 (N_3479,N_1405,N_1933);
or U3480 (N_3480,N_1612,N_694);
xnor U3481 (N_3481,N_229,N_1211);
nor U3482 (N_3482,N_1496,N_787);
and U3483 (N_3483,N_693,N_613);
nor U3484 (N_3484,N_28,N_1452);
and U3485 (N_3485,N_10,N_145);
and U3486 (N_3486,N_243,N_643);
xnor U3487 (N_3487,N_102,N_362);
or U3488 (N_3488,N_376,N_741);
nand U3489 (N_3489,N_1717,N_526);
nor U3490 (N_3490,N_1641,N_325);
xor U3491 (N_3491,N_658,N_1509);
nand U3492 (N_3492,N_466,N_688);
nor U3493 (N_3493,N_1176,N_1460);
nor U3494 (N_3494,N_1128,N_1927);
and U3495 (N_3495,N_881,N_1799);
xnor U3496 (N_3496,N_1304,N_967);
or U3497 (N_3497,N_643,N_1967);
nand U3498 (N_3498,N_1457,N_93);
xor U3499 (N_3499,N_1961,N_1593);
or U3500 (N_3500,N_785,N_350);
and U3501 (N_3501,N_198,N_1786);
nor U3502 (N_3502,N_609,N_1316);
or U3503 (N_3503,N_560,N_457);
xnor U3504 (N_3504,N_1694,N_410);
or U3505 (N_3505,N_791,N_1293);
xor U3506 (N_3506,N_1661,N_963);
or U3507 (N_3507,N_1427,N_1637);
xor U3508 (N_3508,N_773,N_670);
and U3509 (N_3509,N_502,N_331);
and U3510 (N_3510,N_1944,N_1040);
or U3511 (N_3511,N_1617,N_1883);
or U3512 (N_3512,N_815,N_1297);
and U3513 (N_3513,N_71,N_1060);
nand U3514 (N_3514,N_1791,N_200);
xor U3515 (N_3515,N_707,N_1582);
and U3516 (N_3516,N_1362,N_492);
and U3517 (N_3517,N_563,N_997);
xnor U3518 (N_3518,N_325,N_23);
xnor U3519 (N_3519,N_21,N_1427);
nor U3520 (N_3520,N_856,N_1683);
nor U3521 (N_3521,N_1644,N_1019);
xor U3522 (N_3522,N_1103,N_1363);
and U3523 (N_3523,N_384,N_1269);
xor U3524 (N_3524,N_1209,N_1208);
nand U3525 (N_3525,N_240,N_1193);
or U3526 (N_3526,N_508,N_1967);
or U3527 (N_3527,N_1317,N_1197);
or U3528 (N_3528,N_1216,N_964);
nor U3529 (N_3529,N_534,N_1048);
or U3530 (N_3530,N_380,N_610);
or U3531 (N_3531,N_1016,N_562);
xnor U3532 (N_3532,N_1346,N_1506);
nand U3533 (N_3533,N_476,N_321);
and U3534 (N_3534,N_520,N_484);
nor U3535 (N_3535,N_1422,N_1365);
xor U3536 (N_3536,N_28,N_406);
nand U3537 (N_3537,N_1433,N_1768);
and U3538 (N_3538,N_726,N_1573);
and U3539 (N_3539,N_1260,N_89);
xor U3540 (N_3540,N_1895,N_722);
nand U3541 (N_3541,N_1307,N_478);
xnor U3542 (N_3542,N_1709,N_432);
nand U3543 (N_3543,N_983,N_119);
xnor U3544 (N_3544,N_1541,N_1837);
nor U3545 (N_3545,N_1461,N_1326);
nor U3546 (N_3546,N_693,N_1044);
xnor U3547 (N_3547,N_311,N_965);
and U3548 (N_3548,N_1302,N_1362);
or U3549 (N_3549,N_1889,N_233);
nor U3550 (N_3550,N_507,N_1867);
and U3551 (N_3551,N_1231,N_1269);
nor U3552 (N_3552,N_29,N_657);
and U3553 (N_3553,N_1679,N_869);
xnor U3554 (N_3554,N_692,N_23);
and U3555 (N_3555,N_1242,N_1197);
and U3556 (N_3556,N_137,N_1626);
xor U3557 (N_3557,N_790,N_1378);
or U3558 (N_3558,N_1282,N_1576);
xnor U3559 (N_3559,N_1211,N_1104);
nor U3560 (N_3560,N_556,N_1131);
nand U3561 (N_3561,N_782,N_1207);
or U3562 (N_3562,N_1012,N_468);
nor U3563 (N_3563,N_1151,N_652);
or U3564 (N_3564,N_1051,N_192);
or U3565 (N_3565,N_1787,N_1729);
or U3566 (N_3566,N_490,N_1592);
nor U3567 (N_3567,N_925,N_1462);
xor U3568 (N_3568,N_1806,N_1278);
or U3569 (N_3569,N_812,N_1486);
nand U3570 (N_3570,N_226,N_899);
and U3571 (N_3571,N_731,N_1168);
nor U3572 (N_3572,N_493,N_1372);
and U3573 (N_3573,N_523,N_1458);
nor U3574 (N_3574,N_1388,N_1187);
and U3575 (N_3575,N_991,N_1647);
xnor U3576 (N_3576,N_1593,N_273);
nand U3577 (N_3577,N_851,N_946);
nand U3578 (N_3578,N_1055,N_1069);
or U3579 (N_3579,N_1119,N_990);
nor U3580 (N_3580,N_936,N_1946);
and U3581 (N_3581,N_1139,N_1286);
xor U3582 (N_3582,N_1209,N_761);
nor U3583 (N_3583,N_685,N_504);
nor U3584 (N_3584,N_108,N_1953);
nand U3585 (N_3585,N_735,N_1707);
xnor U3586 (N_3586,N_541,N_129);
and U3587 (N_3587,N_1242,N_10);
or U3588 (N_3588,N_1579,N_1657);
nand U3589 (N_3589,N_759,N_394);
or U3590 (N_3590,N_1015,N_1654);
xnor U3591 (N_3591,N_1959,N_1430);
or U3592 (N_3592,N_634,N_1661);
and U3593 (N_3593,N_1636,N_467);
nand U3594 (N_3594,N_1285,N_178);
or U3595 (N_3595,N_955,N_1574);
xnor U3596 (N_3596,N_1676,N_730);
nor U3597 (N_3597,N_732,N_1397);
xnor U3598 (N_3598,N_1590,N_1855);
nor U3599 (N_3599,N_667,N_1918);
nor U3600 (N_3600,N_295,N_1943);
xor U3601 (N_3601,N_170,N_474);
nor U3602 (N_3602,N_215,N_1944);
or U3603 (N_3603,N_757,N_1530);
and U3604 (N_3604,N_229,N_1086);
nand U3605 (N_3605,N_1485,N_337);
or U3606 (N_3606,N_1536,N_1105);
and U3607 (N_3607,N_458,N_946);
or U3608 (N_3608,N_748,N_1567);
nor U3609 (N_3609,N_556,N_898);
nor U3610 (N_3610,N_1729,N_574);
nor U3611 (N_3611,N_1927,N_1127);
nor U3612 (N_3612,N_1552,N_835);
nand U3613 (N_3613,N_1146,N_972);
or U3614 (N_3614,N_605,N_96);
xor U3615 (N_3615,N_1740,N_1138);
and U3616 (N_3616,N_229,N_1770);
nand U3617 (N_3617,N_90,N_407);
nor U3618 (N_3618,N_615,N_1120);
xor U3619 (N_3619,N_525,N_1485);
and U3620 (N_3620,N_1083,N_1043);
and U3621 (N_3621,N_526,N_134);
xor U3622 (N_3622,N_51,N_1572);
or U3623 (N_3623,N_853,N_192);
and U3624 (N_3624,N_277,N_1001);
nor U3625 (N_3625,N_324,N_126);
xor U3626 (N_3626,N_1531,N_800);
and U3627 (N_3627,N_1596,N_1597);
and U3628 (N_3628,N_169,N_301);
nor U3629 (N_3629,N_91,N_657);
xor U3630 (N_3630,N_469,N_1338);
nand U3631 (N_3631,N_57,N_1141);
nand U3632 (N_3632,N_701,N_226);
and U3633 (N_3633,N_1788,N_381);
and U3634 (N_3634,N_1208,N_1705);
xnor U3635 (N_3635,N_1972,N_984);
xor U3636 (N_3636,N_1744,N_471);
and U3637 (N_3637,N_1257,N_45);
nor U3638 (N_3638,N_810,N_1935);
or U3639 (N_3639,N_1038,N_477);
or U3640 (N_3640,N_432,N_1393);
and U3641 (N_3641,N_1363,N_953);
or U3642 (N_3642,N_1161,N_1229);
nor U3643 (N_3643,N_1518,N_540);
nor U3644 (N_3644,N_1447,N_19);
xnor U3645 (N_3645,N_1938,N_134);
or U3646 (N_3646,N_1326,N_72);
or U3647 (N_3647,N_683,N_1177);
and U3648 (N_3648,N_196,N_1394);
and U3649 (N_3649,N_335,N_444);
nor U3650 (N_3650,N_1537,N_1642);
nor U3651 (N_3651,N_512,N_225);
xnor U3652 (N_3652,N_1196,N_1927);
and U3653 (N_3653,N_1946,N_1839);
nand U3654 (N_3654,N_597,N_1973);
xor U3655 (N_3655,N_1877,N_312);
and U3656 (N_3656,N_1723,N_1100);
nand U3657 (N_3657,N_302,N_512);
or U3658 (N_3658,N_344,N_939);
or U3659 (N_3659,N_734,N_1515);
xnor U3660 (N_3660,N_619,N_20);
xor U3661 (N_3661,N_1445,N_202);
nor U3662 (N_3662,N_317,N_676);
and U3663 (N_3663,N_1471,N_1783);
and U3664 (N_3664,N_610,N_260);
and U3665 (N_3665,N_1807,N_1373);
and U3666 (N_3666,N_903,N_39);
or U3667 (N_3667,N_1995,N_1915);
nand U3668 (N_3668,N_479,N_1834);
or U3669 (N_3669,N_1056,N_456);
nand U3670 (N_3670,N_1626,N_315);
or U3671 (N_3671,N_1937,N_1962);
nor U3672 (N_3672,N_819,N_1115);
or U3673 (N_3673,N_945,N_273);
nand U3674 (N_3674,N_811,N_1839);
and U3675 (N_3675,N_275,N_1972);
nand U3676 (N_3676,N_1863,N_895);
nor U3677 (N_3677,N_1947,N_74);
and U3678 (N_3678,N_1656,N_1831);
or U3679 (N_3679,N_1191,N_179);
and U3680 (N_3680,N_114,N_1201);
or U3681 (N_3681,N_1736,N_858);
or U3682 (N_3682,N_1422,N_158);
nand U3683 (N_3683,N_1959,N_1950);
nor U3684 (N_3684,N_1790,N_973);
nand U3685 (N_3685,N_1997,N_281);
xnor U3686 (N_3686,N_1306,N_548);
nand U3687 (N_3687,N_922,N_1733);
xor U3688 (N_3688,N_954,N_349);
xor U3689 (N_3689,N_1542,N_1907);
or U3690 (N_3690,N_1327,N_1504);
nor U3691 (N_3691,N_1995,N_179);
xnor U3692 (N_3692,N_807,N_1996);
or U3693 (N_3693,N_804,N_840);
xnor U3694 (N_3694,N_1809,N_497);
and U3695 (N_3695,N_610,N_373);
nand U3696 (N_3696,N_1268,N_643);
and U3697 (N_3697,N_1267,N_1449);
nor U3698 (N_3698,N_866,N_1952);
and U3699 (N_3699,N_1750,N_1755);
nand U3700 (N_3700,N_1033,N_253);
nand U3701 (N_3701,N_1555,N_609);
nor U3702 (N_3702,N_1748,N_839);
nor U3703 (N_3703,N_1446,N_914);
xor U3704 (N_3704,N_1684,N_1689);
or U3705 (N_3705,N_1676,N_1403);
and U3706 (N_3706,N_163,N_1072);
and U3707 (N_3707,N_566,N_1077);
and U3708 (N_3708,N_1356,N_130);
xor U3709 (N_3709,N_630,N_1569);
xnor U3710 (N_3710,N_409,N_1233);
nor U3711 (N_3711,N_1273,N_1914);
nand U3712 (N_3712,N_425,N_1383);
or U3713 (N_3713,N_724,N_757);
nand U3714 (N_3714,N_884,N_1218);
and U3715 (N_3715,N_1206,N_394);
xor U3716 (N_3716,N_747,N_1169);
nand U3717 (N_3717,N_695,N_1030);
nand U3718 (N_3718,N_1682,N_315);
nand U3719 (N_3719,N_856,N_106);
nor U3720 (N_3720,N_1554,N_731);
and U3721 (N_3721,N_1550,N_843);
and U3722 (N_3722,N_881,N_1558);
and U3723 (N_3723,N_1442,N_1919);
nor U3724 (N_3724,N_1496,N_83);
xor U3725 (N_3725,N_263,N_1425);
nor U3726 (N_3726,N_1575,N_1211);
and U3727 (N_3727,N_852,N_4);
nor U3728 (N_3728,N_480,N_775);
and U3729 (N_3729,N_489,N_1638);
or U3730 (N_3730,N_921,N_187);
or U3731 (N_3731,N_622,N_1508);
nand U3732 (N_3732,N_325,N_707);
xnor U3733 (N_3733,N_710,N_1255);
and U3734 (N_3734,N_224,N_1616);
xnor U3735 (N_3735,N_38,N_1134);
nand U3736 (N_3736,N_933,N_524);
or U3737 (N_3737,N_1237,N_1382);
nand U3738 (N_3738,N_685,N_1701);
nor U3739 (N_3739,N_905,N_1589);
and U3740 (N_3740,N_149,N_377);
or U3741 (N_3741,N_363,N_173);
and U3742 (N_3742,N_1200,N_1663);
or U3743 (N_3743,N_543,N_1499);
nand U3744 (N_3744,N_1361,N_1820);
nand U3745 (N_3745,N_1832,N_1068);
or U3746 (N_3746,N_479,N_188);
nor U3747 (N_3747,N_978,N_120);
xor U3748 (N_3748,N_991,N_1132);
and U3749 (N_3749,N_1433,N_358);
nor U3750 (N_3750,N_880,N_1144);
nor U3751 (N_3751,N_1061,N_929);
and U3752 (N_3752,N_1715,N_15);
nor U3753 (N_3753,N_414,N_450);
nand U3754 (N_3754,N_476,N_1817);
nand U3755 (N_3755,N_1782,N_1186);
xnor U3756 (N_3756,N_264,N_563);
nor U3757 (N_3757,N_1765,N_1513);
nor U3758 (N_3758,N_1360,N_844);
and U3759 (N_3759,N_882,N_1350);
nand U3760 (N_3760,N_590,N_589);
nand U3761 (N_3761,N_994,N_120);
xnor U3762 (N_3762,N_1427,N_466);
nor U3763 (N_3763,N_336,N_474);
or U3764 (N_3764,N_375,N_1013);
nand U3765 (N_3765,N_870,N_484);
xor U3766 (N_3766,N_807,N_1192);
nor U3767 (N_3767,N_1525,N_1582);
or U3768 (N_3768,N_1022,N_963);
or U3769 (N_3769,N_1010,N_1092);
nor U3770 (N_3770,N_389,N_215);
or U3771 (N_3771,N_558,N_641);
nand U3772 (N_3772,N_1635,N_673);
xor U3773 (N_3773,N_594,N_1399);
or U3774 (N_3774,N_1778,N_1403);
or U3775 (N_3775,N_1795,N_970);
and U3776 (N_3776,N_1301,N_761);
or U3777 (N_3777,N_1588,N_786);
xnor U3778 (N_3778,N_761,N_1212);
nand U3779 (N_3779,N_717,N_1152);
xor U3780 (N_3780,N_1685,N_894);
nand U3781 (N_3781,N_668,N_1315);
or U3782 (N_3782,N_1471,N_603);
xor U3783 (N_3783,N_163,N_1680);
nand U3784 (N_3784,N_1164,N_1739);
nor U3785 (N_3785,N_999,N_489);
nand U3786 (N_3786,N_1600,N_300);
nor U3787 (N_3787,N_468,N_354);
xor U3788 (N_3788,N_1060,N_197);
and U3789 (N_3789,N_653,N_150);
nor U3790 (N_3790,N_981,N_791);
or U3791 (N_3791,N_896,N_92);
nor U3792 (N_3792,N_952,N_776);
and U3793 (N_3793,N_1699,N_985);
xnor U3794 (N_3794,N_619,N_330);
xor U3795 (N_3795,N_541,N_1979);
nand U3796 (N_3796,N_1959,N_1362);
nor U3797 (N_3797,N_1808,N_1072);
nor U3798 (N_3798,N_328,N_80);
and U3799 (N_3799,N_1319,N_1298);
or U3800 (N_3800,N_126,N_89);
xnor U3801 (N_3801,N_1656,N_912);
or U3802 (N_3802,N_1564,N_1343);
or U3803 (N_3803,N_403,N_733);
and U3804 (N_3804,N_1886,N_1599);
nor U3805 (N_3805,N_399,N_1662);
nor U3806 (N_3806,N_1885,N_423);
nand U3807 (N_3807,N_1593,N_571);
xnor U3808 (N_3808,N_1923,N_1456);
xnor U3809 (N_3809,N_113,N_1233);
nor U3810 (N_3810,N_1254,N_72);
nor U3811 (N_3811,N_1371,N_1706);
and U3812 (N_3812,N_1036,N_1396);
nor U3813 (N_3813,N_1168,N_710);
nor U3814 (N_3814,N_1514,N_1507);
nor U3815 (N_3815,N_610,N_362);
xnor U3816 (N_3816,N_173,N_777);
nor U3817 (N_3817,N_399,N_249);
or U3818 (N_3818,N_961,N_805);
or U3819 (N_3819,N_1875,N_44);
nand U3820 (N_3820,N_371,N_89);
nor U3821 (N_3821,N_328,N_466);
or U3822 (N_3822,N_957,N_363);
and U3823 (N_3823,N_944,N_1594);
or U3824 (N_3824,N_1279,N_1322);
nand U3825 (N_3825,N_1359,N_681);
or U3826 (N_3826,N_1291,N_1381);
and U3827 (N_3827,N_773,N_606);
xor U3828 (N_3828,N_1230,N_1441);
nor U3829 (N_3829,N_1871,N_418);
nor U3830 (N_3830,N_818,N_705);
nand U3831 (N_3831,N_1124,N_136);
nand U3832 (N_3832,N_900,N_1576);
nor U3833 (N_3833,N_1995,N_78);
xnor U3834 (N_3834,N_46,N_1896);
xor U3835 (N_3835,N_1392,N_597);
and U3836 (N_3836,N_1585,N_131);
and U3837 (N_3837,N_326,N_705);
and U3838 (N_3838,N_1130,N_1690);
xnor U3839 (N_3839,N_1386,N_1927);
nand U3840 (N_3840,N_1146,N_780);
or U3841 (N_3841,N_1072,N_313);
or U3842 (N_3842,N_759,N_834);
nand U3843 (N_3843,N_843,N_1960);
and U3844 (N_3844,N_383,N_1436);
and U3845 (N_3845,N_849,N_338);
nor U3846 (N_3846,N_620,N_1925);
nor U3847 (N_3847,N_1782,N_1561);
nor U3848 (N_3848,N_512,N_508);
xor U3849 (N_3849,N_1129,N_1340);
nor U3850 (N_3850,N_1104,N_772);
nand U3851 (N_3851,N_1603,N_665);
nand U3852 (N_3852,N_480,N_647);
xnor U3853 (N_3853,N_253,N_1553);
xor U3854 (N_3854,N_1423,N_812);
and U3855 (N_3855,N_1119,N_1434);
or U3856 (N_3856,N_1293,N_1536);
or U3857 (N_3857,N_155,N_491);
and U3858 (N_3858,N_1109,N_1531);
and U3859 (N_3859,N_1188,N_649);
nand U3860 (N_3860,N_847,N_575);
xnor U3861 (N_3861,N_1464,N_1386);
or U3862 (N_3862,N_183,N_675);
or U3863 (N_3863,N_122,N_840);
xnor U3864 (N_3864,N_263,N_1070);
nor U3865 (N_3865,N_35,N_927);
or U3866 (N_3866,N_1623,N_651);
and U3867 (N_3867,N_1164,N_694);
and U3868 (N_3868,N_1705,N_1595);
nand U3869 (N_3869,N_1987,N_194);
xor U3870 (N_3870,N_1345,N_1901);
nor U3871 (N_3871,N_648,N_706);
nand U3872 (N_3872,N_968,N_452);
nor U3873 (N_3873,N_683,N_1447);
or U3874 (N_3874,N_1991,N_154);
and U3875 (N_3875,N_705,N_784);
and U3876 (N_3876,N_1932,N_1346);
or U3877 (N_3877,N_1499,N_433);
xor U3878 (N_3878,N_1774,N_1366);
xor U3879 (N_3879,N_540,N_1279);
xor U3880 (N_3880,N_189,N_1366);
or U3881 (N_3881,N_1746,N_1273);
nor U3882 (N_3882,N_1089,N_1218);
and U3883 (N_3883,N_1012,N_110);
or U3884 (N_3884,N_1286,N_946);
nand U3885 (N_3885,N_1214,N_835);
or U3886 (N_3886,N_979,N_1731);
nor U3887 (N_3887,N_57,N_1352);
nor U3888 (N_3888,N_1273,N_261);
nor U3889 (N_3889,N_1030,N_519);
nand U3890 (N_3890,N_1279,N_230);
nand U3891 (N_3891,N_1814,N_1381);
and U3892 (N_3892,N_1920,N_53);
nor U3893 (N_3893,N_139,N_337);
and U3894 (N_3894,N_6,N_1093);
nand U3895 (N_3895,N_83,N_1528);
nor U3896 (N_3896,N_429,N_508);
or U3897 (N_3897,N_608,N_281);
or U3898 (N_3898,N_336,N_377);
or U3899 (N_3899,N_1576,N_1194);
and U3900 (N_3900,N_420,N_700);
xnor U3901 (N_3901,N_280,N_1959);
nor U3902 (N_3902,N_53,N_411);
nand U3903 (N_3903,N_1987,N_1838);
xor U3904 (N_3904,N_217,N_451);
nand U3905 (N_3905,N_337,N_268);
xnor U3906 (N_3906,N_474,N_123);
and U3907 (N_3907,N_1917,N_154);
xor U3908 (N_3908,N_579,N_899);
or U3909 (N_3909,N_1682,N_540);
xor U3910 (N_3910,N_105,N_610);
or U3911 (N_3911,N_587,N_1055);
and U3912 (N_3912,N_1956,N_1782);
nor U3913 (N_3913,N_1573,N_1658);
and U3914 (N_3914,N_1840,N_1113);
nor U3915 (N_3915,N_293,N_939);
and U3916 (N_3916,N_608,N_1772);
and U3917 (N_3917,N_1177,N_602);
xor U3918 (N_3918,N_1704,N_1200);
nand U3919 (N_3919,N_484,N_1825);
nand U3920 (N_3920,N_319,N_129);
nand U3921 (N_3921,N_1399,N_190);
nor U3922 (N_3922,N_1358,N_1450);
nor U3923 (N_3923,N_1752,N_346);
nand U3924 (N_3924,N_678,N_257);
and U3925 (N_3925,N_1157,N_194);
nor U3926 (N_3926,N_1988,N_32);
or U3927 (N_3927,N_1788,N_39);
or U3928 (N_3928,N_882,N_1095);
or U3929 (N_3929,N_1228,N_1373);
nand U3930 (N_3930,N_1767,N_370);
xor U3931 (N_3931,N_131,N_990);
nand U3932 (N_3932,N_1095,N_1028);
and U3933 (N_3933,N_1335,N_1247);
and U3934 (N_3934,N_1811,N_787);
or U3935 (N_3935,N_38,N_1012);
or U3936 (N_3936,N_1878,N_1586);
xor U3937 (N_3937,N_1984,N_10);
or U3938 (N_3938,N_465,N_327);
nand U3939 (N_3939,N_1951,N_940);
nand U3940 (N_3940,N_1468,N_1274);
nand U3941 (N_3941,N_100,N_264);
or U3942 (N_3942,N_1734,N_1221);
nand U3943 (N_3943,N_909,N_1578);
nor U3944 (N_3944,N_163,N_1625);
nor U3945 (N_3945,N_989,N_484);
or U3946 (N_3946,N_649,N_1322);
or U3947 (N_3947,N_1232,N_1500);
xnor U3948 (N_3948,N_447,N_949);
or U3949 (N_3949,N_1884,N_386);
nand U3950 (N_3950,N_1109,N_4);
and U3951 (N_3951,N_11,N_1820);
nor U3952 (N_3952,N_1475,N_367);
nor U3953 (N_3953,N_1046,N_735);
nor U3954 (N_3954,N_1959,N_1913);
or U3955 (N_3955,N_1906,N_739);
or U3956 (N_3956,N_473,N_1515);
and U3957 (N_3957,N_1876,N_750);
or U3958 (N_3958,N_1962,N_844);
and U3959 (N_3959,N_203,N_670);
or U3960 (N_3960,N_1219,N_1642);
or U3961 (N_3961,N_574,N_1602);
nor U3962 (N_3962,N_769,N_512);
and U3963 (N_3963,N_2,N_1976);
and U3964 (N_3964,N_908,N_767);
xnor U3965 (N_3965,N_1595,N_1805);
nand U3966 (N_3966,N_689,N_1890);
nor U3967 (N_3967,N_735,N_915);
nand U3968 (N_3968,N_528,N_905);
and U3969 (N_3969,N_1684,N_1749);
or U3970 (N_3970,N_1790,N_356);
nor U3971 (N_3971,N_1243,N_427);
nor U3972 (N_3972,N_1053,N_975);
nand U3973 (N_3973,N_1815,N_1962);
or U3974 (N_3974,N_119,N_1951);
xnor U3975 (N_3975,N_558,N_84);
and U3976 (N_3976,N_1143,N_1370);
or U3977 (N_3977,N_378,N_1597);
nand U3978 (N_3978,N_450,N_840);
and U3979 (N_3979,N_393,N_512);
and U3980 (N_3980,N_1570,N_1025);
nor U3981 (N_3981,N_1409,N_110);
or U3982 (N_3982,N_416,N_1651);
xnor U3983 (N_3983,N_950,N_1489);
xor U3984 (N_3984,N_1988,N_762);
nor U3985 (N_3985,N_1741,N_528);
xnor U3986 (N_3986,N_1607,N_1844);
xnor U3987 (N_3987,N_939,N_198);
xor U3988 (N_3988,N_302,N_28);
and U3989 (N_3989,N_1669,N_847);
or U3990 (N_3990,N_121,N_1466);
and U3991 (N_3991,N_1507,N_490);
or U3992 (N_3992,N_6,N_1457);
nand U3993 (N_3993,N_495,N_1041);
nor U3994 (N_3994,N_1148,N_1434);
or U3995 (N_3995,N_684,N_121);
or U3996 (N_3996,N_997,N_1431);
xor U3997 (N_3997,N_1569,N_928);
nor U3998 (N_3998,N_591,N_1019);
and U3999 (N_3999,N_986,N_676);
and U4000 (N_4000,N_3135,N_2759);
xnor U4001 (N_4001,N_3472,N_3981);
xor U4002 (N_4002,N_2585,N_2122);
or U4003 (N_4003,N_3658,N_2256);
or U4004 (N_4004,N_2506,N_3361);
nand U4005 (N_4005,N_2396,N_2682);
nand U4006 (N_4006,N_3807,N_3786);
or U4007 (N_4007,N_3196,N_3469);
nor U4008 (N_4008,N_2721,N_3443);
xor U4009 (N_4009,N_3206,N_3440);
and U4010 (N_4010,N_2061,N_3181);
or U4011 (N_4011,N_3987,N_3737);
nor U4012 (N_4012,N_2041,N_3360);
nand U4013 (N_4013,N_2444,N_3405);
nand U4014 (N_4014,N_2312,N_2640);
nand U4015 (N_4015,N_2090,N_2969);
xor U4016 (N_4016,N_2279,N_3757);
and U4017 (N_4017,N_3130,N_3780);
and U4018 (N_4018,N_3003,N_3725);
nor U4019 (N_4019,N_2622,N_2539);
nor U4020 (N_4020,N_3313,N_3842);
xor U4021 (N_4021,N_2915,N_2820);
and U4022 (N_4022,N_3754,N_2810);
nor U4023 (N_4023,N_3393,N_3805);
or U4024 (N_4024,N_3076,N_2386);
nand U4025 (N_4025,N_3178,N_2275);
and U4026 (N_4026,N_2778,N_3494);
nor U4027 (N_4027,N_3389,N_3948);
nor U4028 (N_4028,N_3518,N_3704);
or U4029 (N_4029,N_3403,N_2616);
nand U4030 (N_4030,N_3101,N_2450);
xor U4031 (N_4031,N_2557,N_2966);
or U4032 (N_4032,N_2562,N_3061);
or U4033 (N_4033,N_3237,N_3363);
or U4034 (N_4034,N_2590,N_3722);
or U4035 (N_4035,N_3572,N_3610);
and U4036 (N_4036,N_2814,N_2344);
nor U4037 (N_4037,N_3983,N_2528);
xnor U4038 (N_4038,N_2319,N_3249);
xor U4039 (N_4039,N_2037,N_3154);
or U4040 (N_4040,N_2132,N_2025);
xnor U4041 (N_4041,N_2161,N_3930);
or U4042 (N_4042,N_3335,N_3123);
nor U4043 (N_4043,N_2001,N_3497);
nor U4044 (N_4044,N_2210,N_3604);
xor U4045 (N_4045,N_2375,N_3296);
nand U4046 (N_4046,N_2179,N_2443);
xor U4047 (N_4047,N_3671,N_2304);
nand U4048 (N_4048,N_2584,N_3120);
xnor U4049 (N_4049,N_3751,N_2599);
nand U4050 (N_4050,N_2978,N_3906);
xnor U4051 (N_4051,N_2068,N_2149);
or U4052 (N_4052,N_3759,N_2769);
nand U4053 (N_4053,N_2441,N_2994);
nor U4054 (N_4054,N_2937,N_3862);
nand U4055 (N_4055,N_3039,N_2614);
nor U4056 (N_4056,N_3687,N_2070);
nor U4057 (N_4057,N_3733,N_3090);
or U4058 (N_4058,N_2799,N_3033);
or U4059 (N_4059,N_3150,N_2148);
nor U4060 (N_4060,N_2415,N_2788);
nor U4061 (N_4061,N_3867,N_3750);
or U4062 (N_4062,N_3266,N_3878);
or U4063 (N_4063,N_3345,N_2139);
xnor U4064 (N_4064,N_3125,N_3846);
and U4065 (N_4065,N_3517,N_2589);
and U4066 (N_4066,N_3634,N_3096);
and U4067 (N_4067,N_3635,N_3895);
nand U4068 (N_4068,N_3719,N_3121);
or U4069 (N_4069,N_3740,N_3914);
nor U4070 (N_4070,N_2125,N_2498);
nand U4071 (N_4071,N_3617,N_2992);
and U4072 (N_4072,N_2389,N_3378);
or U4073 (N_4073,N_2427,N_2483);
nand U4074 (N_4074,N_2845,N_3225);
and U4075 (N_4075,N_3590,N_2475);
and U4076 (N_4076,N_2896,N_3253);
nand U4077 (N_4077,N_2348,N_3723);
and U4078 (N_4078,N_3556,N_3925);
nand U4079 (N_4079,N_2251,N_3007);
nor U4080 (N_4080,N_2807,N_3713);
nand U4081 (N_4081,N_3770,N_3765);
nor U4082 (N_4082,N_2363,N_3029);
and U4083 (N_4083,N_2581,N_2648);
or U4084 (N_4084,N_2397,N_2071);
nand U4085 (N_4085,N_2979,N_3038);
xor U4086 (N_4086,N_3674,N_3201);
xor U4087 (N_4087,N_2487,N_3295);
nor U4088 (N_4088,N_3383,N_2752);
nand U4089 (N_4089,N_2980,N_3407);
nor U4090 (N_4090,N_3025,N_2123);
or U4091 (N_4091,N_2257,N_2138);
or U4092 (N_4092,N_3756,N_2631);
xnor U4093 (N_4093,N_3338,N_2731);
xor U4094 (N_4094,N_2954,N_2129);
xor U4095 (N_4095,N_3406,N_2091);
nand U4096 (N_4096,N_3220,N_3709);
nor U4097 (N_4097,N_3479,N_2962);
or U4098 (N_4098,N_3174,N_3002);
nor U4099 (N_4099,N_2824,N_2703);
nor U4100 (N_4100,N_2701,N_2904);
and U4101 (N_4101,N_3422,N_3144);
nand U4102 (N_4102,N_2783,N_3790);
nand U4103 (N_4103,N_3591,N_3132);
nand U4104 (N_4104,N_2505,N_2827);
nand U4105 (N_4105,N_2474,N_3369);
nor U4106 (N_4106,N_3398,N_2288);
nand U4107 (N_4107,N_2033,N_2185);
xor U4108 (N_4108,N_2740,N_2838);
and U4109 (N_4109,N_3385,N_2228);
and U4110 (N_4110,N_2677,N_3021);
nor U4111 (N_4111,N_3928,N_2434);
and U4112 (N_4112,N_3062,N_2993);
or U4113 (N_4113,N_3368,N_3362);
nand U4114 (N_4114,N_2891,N_3173);
xor U4115 (N_4115,N_3341,N_2008);
xnor U4116 (N_4116,N_2758,N_3379);
nor U4117 (N_4117,N_3030,N_3921);
nor U4118 (N_4118,N_3277,N_3834);
and U4119 (N_4119,N_3016,N_2446);
nand U4120 (N_4120,N_3408,N_2399);
nand U4121 (N_4121,N_2750,N_3886);
nand U4122 (N_4122,N_3190,N_3084);
nand U4123 (N_4123,N_2354,N_3170);
or U4124 (N_4124,N_2239,N_2739);
nand U4125 (N_4125,N_2930,N_3923);
nand U4126 (N_4126,N_3143,N_2565);
nor U4127 (N_4127,N_3718,N_3911);
nor U4128 (N_4128,N_3072,N_2559);
nand U4129 (N_4129,N_2236,N_2801);
nor U4130 (N_4130,N_2112,N_2477);
nand U4131 (N_4131,N_3108,N_2267);
xnor U4132 (N_4132,N_3186,N_2658);
or U4133 (N_4133,N_3373,N_2080);
xor U4134 (N_4134,N_2381,N_2699);
nor U4135 (N_4135,N_3870,N_3013);
xor U4136 (N_4136,N_3187,N_3789);
nor U4137 (N_4137,N_2202,N_2400);
or U4138 (N_4138,N_3328,N_2489);
xor U4139 (N_4139,N_3285,N_2544);
xnor U4140 (N_4140,N_2253,N_2413);
nand U4141 (N_4141,N_2373,N_2651);
nand U4142 (N_4142,N_3419,N_2482);
and U4143 (N_4143,N_2774,N_3648);
and U4144 (N_4144,N_2812,N_3997);
or U4145 (N_4145,N_3926,N_3668);
nand U4146 (N_4146,N_2481,N_2555);
xnor U4147 (N_4147,N_3031,N_2021);
or U4148 (N_4148,N_2195,N_2337);
nor U4149 (N_4149,N_2765,N_2999);
nand U4150 (N_4150,N_3066,N_3631);
and U4151 (N_4151,N_2895,N_3017);
xnor U4152 (N_4152,N_2905,N_2645);
or U4153 (N_4153,N_2164,N_3176);
and U4154 (N_4154,N_3166,N_2696);
or U4155 (N_4155,N_3149,N_2833);
nor U4156 (N_4156,N_2692,N_2115);
nand U4157 (N_4157,N_3571,N_3113);
nor U4158 (N_4158,N_2851,N_2763);
nor U4159 (N_4159,N_2791,N_3649);
nor U4160 (N_4160,N_3514,N_2742);
and U4161 (N_4161,N_2675,N_3755);
or U4162 (N_4162,N_3357,N_3473);
and U4163 (N_4163,N_3601,N_3550);
and U4164 (N_4164,N_3816,N_2917);
and U4165 (N_4165,N_2366,N_2294);
or U4166 (N_4166,N_2554,N_3441);
and U4167 (N_4167,N_2307,N_2280);
and U4168 (N_4168,N_3814,N_3138);
nor U4169 (N_4169,N_3808,N_2828);
nand U4170 (N_4170,N_3425,N_2802);
or U4171 (N_4171,N_3124,N_3359);
xnor U4172 (N_4172,N_3258,N_2031);
or U4173 (N_4173,N_2469,N_2748);
nor U4174 (N_4174,N_2015,N_2159);
xor U4175 (N_4175,N_2087,N_3436);
nor U4176 (N_4176,N_2078,N_2325);
or U4177 (N_4177,N_3105,N_3574);
or U4178 (N_4178,N_3792,N_2367);
and U4179 (N_4179,N_3223,N_2704);
or U4180 (N_4180,N_3411,N_2852);
nor U4181 (N_4181,N_3724,N_2391);
nor U4182 (N_4182,N_2884,N_3071);
nand U4183 (N_4183,N_2153,N_2277);
or U4184 (N_4184,N_3698,N_3730);
nand U4185 (N_4185,N_3250,N_2881);
nand U4186 (N_4186,N_2231,N_2949);
nand U4187 (N_4187,N_2611,N_3483);
or U4188 (N_4188,N_2732,N_2005);
or U4189 (N_4189,N_3712,N_3855);
xnor U4190 (N_4190,N_2020,N_2735);
nand U4191 (N_4191,N_2471,N_3191);
nor U4192 (N_4192,N_3578,N_2686);
and U4193 (N_4193,N_2500,N_2951);
and U4194 (N_4194,N_2203,N_2309);
and U4195 (N_4195,N_3133,N_3804);
nor U4196 (N_4196,N_3056,N_2835);
or U4197 (N_4197,N_3640,N_2933);
nand U4198 (N_4198,N_3330,N_2550);
xnor U4199 (N_4199,N_3800,N_2250);
nor U4200 (N_4200,N_2330,N_3563);
xnor U4201 (N_4201,N_3868,N_3859);
or U4202 (N_4202,N_2369,N_2627);
or U4203 (N_4203,N_2998,N_3717);
or U4204 (N_4204,N_3207,N_3197);
and U4205 (N_4205,N_2743,N_3284);
and U4206 (N_4206,N_3972,N_3613);
or U4207 (N_4207,N_2160,N_2026);
and U4208 (N_4208,N_3307,N_2177);
xnor U4209 (N_4209,N_2972,N_2119);
or U4210 (N_4210,N_3272,N_3795);
or U4211 (N_4211,N_3290,N_2313);
nor U4212 (N_4212,N_2927,N_3561);
nand U4213 (N_4213,N_2379,N_2150);
or U4214 (N_4214,N_2853,N_3882);
nand U4215 (N_4215,N_2105,N_2570);
xor U4216 (N_4216,N_3965,N_3141);
nand U4217 (N_4217,N_3232,N_3305);
or U4218 (N_4218,N_2051,N_3306);
or U4219 (N_4219,N_3465,N_2734);
xor U4220 (N_4220,N_3890,N_3597);
nor U4221 (N_4221,N_3727,N_2308);
xor U4222 (N_4222,N_3519,N_2270);
nand U4223 (N_4223,N_2878,N_2720);
nor U4224 (N_4224,N_2662,N_3492);
nor U4225 (N_4225,N_3278,N_3034);
nand U4226 (N_4226,N_3523,N_2568);
and U4227 (N_4227,N_2871,N_2310);
and U4228 (N_4228,N_3689,N_2221);
xnor U4229 (N_4229,N_2002,N_3311);
and U4230 (N_4230,N_2754,N_2401);
xnor U4231 (N_4231,N_2155,N_2198);
nor U4232 (N_4232,N_3421,N_2587);
xor U4233 (N_4233,N_2844,N_2715);
and U4234 (N_4234,N_3380,N_3998);
nor U4235 (N_4235,N_2054,N_2111);
nand U4236 (N_4236,N_3785,N_2421);
nor U4237 (N_4237,N_3666,N_2047);
xnor U4238 (N_4238,N_2772,N_2695);
nor U4239 (N_4239,N_3264,N_3970);
or U4240 (N_4240,N_3280,N_2208);
xnor U4241 (N_4241,N_2350,N_3018);
xor U4242 (N_4242,N_2594,N_2245);
or U4243 (N_4243,N_2121,N_2151);
and U4244 (N_4244,N_3244,N_2171);
nand U4245 (N_4245,N_2635,N_2916);
xnor U4246 (N_4246,N_3619,N_2621);
nand U4247 (N_4247,N_3701,N_3739);
nand U4248 (N_4248,N_2362,N_3760);
nand U4249 (N_4249,N_2235,N_2628);
or U4250 (N_4250,N_3657,N_2227);
nor U4251 (N_4251,N_2777,N_3035);
or U4252 (N_4252,N_3200,N_2689);
nor U4253 (N_4253,N_2560,N_2900);
nand U4254 (N_4254,N_3447,N_2861);
xnor U4255 (N_4255,N_3866,N_3324);
nor U4256 (N_4256,N_2664,N_3820);
nand U4257 (N_4257,N_2302,N_3188);
nor U4258 (N_4258,N_2580,N_3884);
xor U4259 (N_4259,N_2947,N_2417);
or U4260 (N_4260,N_2893,N_3944);
xnor U4261 (N_4261,N_3799,N_2744);
xor U4262 (N_4262,N_2394,N_3559);
or U4263 (N_4263,N_3894,N_3158);
xnor U4264 (N_4264,N_3932,N_2839);
and U4265 (N_4265,N_3773,N_2960);
nor U4266 (N_4266,N_3252,N_3055);
nor U4267 (N_4267,N_2175,N_2058);
xor U4268 (N_4268,N_3539,N_2452);
or U4269 (N_4269,N_3516,N_2096);
and U4270 (N_4270,N_3414,N_2242);
xor U4271 (N_4271,N_3122,N_3481);
nor U4272 (N_4272,N_2234,N_3747);
nand U4273 (N_4273,N_3630,N_3708);
nor U4274 (N_4274,N_2535,N_3929);
nand U4275 (N_4275,N_3140,N_2079);
nor U4276 (N_4276,N_2049,N_3475);
and U4277 (N_4277,N_3391,N_3297);
xnor U4278 (N_4278,N_2502,N_3491);
or U4279 (N_4279,N_2120,N_3938);
nand U4280 (N_4280,N_2848,N_2532);
xnor U4281 (N_4281,N_3169,N_2263);
and U4282 (N_4282,N_2605,N_3962);
or U4283 (N_4283,N_2693,N_3893);
nand U4284 (N_4284,N_2097,N_3697);
and U4285 (N_4285,N_2448,N_3386);
or U4286 (N_4286,N_2118,N_2901);
nand U4287 (N_4287,N_2856,N_2521);
and U4288 (N_4288,N_2062,N_3008);
and U4289 (N_4289,N_2886,N_2538);
xor U4290 (N_4290,N_2874,N_3524);
nand U4291 (N_4291,N_2178,N_2547);
or U4292 (N_4292,N_2322,N_3194);
nand U4293 (N_4293,N_2305,N_2066);
or U4294 (N_4294,N_3675,N_2619);
and U4295 (N_4295,N_2016,N_2811);
or U4296 (N_4296,N_3470,N_3001);
and U4297 (N_4297,N_3788,N_2166);
or U4298 (N_4298,N_2790,N_2552);
nor U4299 (N_4299,N_2238,N_2470);
or U4300 (N_4300,N_3986,N_3706);
or U4301 (N_4301,N_3486,N_3390);
and U4302 (N_4302,N_3507,N_3288);
and U4303 (N_4303,N_2958,N_3243);
or U4304 (N_4304,N_2387,N_2600);
and U4305 (N_4305,N_3241,N_2566);
nand U4306 (N_4306,N_2287,N_2467);
nand U4307 (N_4307,N_2113,N_2406);
nand U4308 (N_4308,N_3769,N_2233);
nand U4309 (N_4309,N_3199,N_2085);
or U4310 (N_4310,N_3683,N_3294);
nor U4311 (N_4311,N_3364,N_2081);
or U4312 (N_4312,N_2717,N_2840);
or U4313 (N_4313,N_2768,N_2215);
or U4314 (N_4314,N_3980,N_3248);
or U4315 (N_4315,N_2723,N_2045);
or U4316 (N_4316,N_2558,N_3899);
nor U4317 (N_4317,N_3323,N_2593);
nand U4318 (N_4318,N_2244,N_3404);
nor U4319 (N_4319,N_3812,N_3234);
nor U4320 (N_4320,N_2847,N_3106);
and U4321 (N_4321,N_2213,N_3839);
and U4322 (N_4322,N_2346,N_2914);
nor U4323 (N_4323,N_3114,N_3829);
xnor U4324 (N_4324,N_3728,N_3694);
xnor U4325 (N_4325,N_2464,N_3978);
and U4326 (N_4326,N_3869,N_3427);
and U4327 (N_4327,N_3749,N_2518);
nor U4328 (N_4328,N_2286,N_2935);
and U4329 (N_4329,N_3794,N_2869);
and U4330 (N_4330,N_3267,N_3119);
and U4331 (N_4331,N_2412,N_2542);
xor U4332 (N_4332,N_2347,N_3576);
nand U4333 (N_4333,N_3742,N_2385);
nand U4334 (N_4334,N_2495,N_3355);
or U4335 (N_4335,N_3209,N_2598);
nand U4336 (N_4336,N_2331,N_2109);
xnor U4337 (N_4337,N_3005,N_2410);
or U4338 (N_4338,N_3976,N_2629);
nor U4339 (N_4339,N_2486,N_2702);
xnor U4340 (N_4340,N_3195,N_2977);
xor U4341 (N_4341,N_3402,N_2345);
xor U4342 (N_4342,N_2249,N_2336);
nand U4343 (N_4343,N_3953,N_2255);
nand U4344 (N_4344,N_3115,N_2268);
xnor U4345 (N_4345,N_3919,N_2083);
nand U4346 (N_4346,N_3908,N_2667);
or U4347 (N_4347,N_3924,N_3089);
nor U4348 (N_4348,N_2468,N_2318);
and U4349 (N_4349,N_2541,N_2719);
xnor U4350 (N_4350,N_2700,N_2529);
xor U4351 (N_4351,N_3684,N_3830);
nor U4352 (N_4352,N_2816,N_3283);
or U4353 (N_4353,N_3850,N_2760);
nand U4354 (N_4354,N_3471,N_3058);
or U4355 (N_4355,N_2128,N_3399);
and U4356 (N_4356,N_2491,N_2747);
or U4357 (N_4357,N_3575,N_3877);
or U4358 (N_4358,N_3889,N_3450);
and U4359 (N_4359,N_3989,N_3845);
xor U4360 (N_4360,N_2826,N_3735);
xnor U4361 (N_4361,N_3676,N_2613);
nor U4362 (N_4362,N_3536,N_3961);
nor U4363 (N_4363,N_2197,N_2194);
and U4364 (N_4364,N_3641,N_2984);
nand U4365 (N_4365,N_3616,N_3875);
or U4366 (N_4366,N_3024,N_3336);
nor U4367 (N_4367,N_3478,N_2862);
and U4368 (N_4368,N_3065,N_3269);
and U4369 (N_4369,N_3831,N_3111);
xnor U4370 (N_4370,N_3711,N_3358);
nand U4371 (N_4371,N_3192,N_3552);
xor U4372 (N_4372,N_3157,N_3618);
xnor U4373 (N_4373,N_2261,N_2134);
and U4374 (N_4374,N_2618,N_3857);
and U4375 (N_4375,N_3520,N_3088);
and U4376 (N_4376,N_3412,N_3973);
or U4377 (N_4377,N_3851,N_3340);
and U4378 (N_4378,N_2019,N_3185);
nor U4379 (N_4379,N_2656,N_3710);
and U4380 (N_4380,N_3881,N_3963);
xor U4381 (N_4381,N_2059,N_2334);
nand U4382 (N_4382,N_2205,N_2642);
nand U4383 (N_4383,N_3876,N_3535);
and U4384 (N_4384,N_3334,N_3605);
and U4385 (N_4385,N_3049,N_3462);
and U4386 (N_4386,N_3325,N_2918);
and U4387 (N_4387,N_2782,N_3651);
or U4388 (N_4388,N_3164,N_2865);
nor U4389 (N_4389,N_3463,N_3621);
xnor U4390 (N_4390,N_3104,N_3037);
or U4391 (N_4391,N_3318,N_3594);
nor U4392 (N_4392,N_3655,N_3316);
nand U4393 (N_4393,N_3918,N_2643);
xor U4394 (N_4394,N_2990,N_3162);
nand U4395 (N_4395,N_2463,N_3303);
xnor U4396 (N_4396,N_3409,N_3160);
nor U4397 (N_4397,N_2982,N_3118);
and U4398 (N_4398,N_2104,N_3901);
nor U4399 (N_4399,N_3545,N_2110);
nand U4400 (N_4400,N_2262,N_3585);
xnor U4401 (N_4401,N_2784,N_2252);
xnor U4402 (N_4402,N_3579,N_2316);
xor U4403 (N_4403,N_2923,N_2329);
nand U4404 (N_4404,N_2357,N_2407);
and U4405 (N_4405,N_3082,N_3534);
nand U4406 (N_4406,N_3951,N_2511);
nand U4407 (N_4407,N_3716,N_2892);
xnor U4408 (N_4408,N_3246,N_2564);
nor U4409 (N_4409,N_3047,N_2516);
nor U4410 (N_4410,N_2416,N_3686);
xnor U4411 (N_4411,N_3080,N_3966);
xnor U4412 (N_4412,N_3569,N_2145);
nand U4413 (N_4413,N_2805,N_3646);
xor U4414 (N_4414,N_2187,N_2950);
nor U4415 (N_4415,N_3401,N_3499);
xor U4416 (N_4416,N_2147,N_2738);
and U4417 (N_4417,N_3078,N_2439);
and U4418 (N_4418,N_3212,N_2885);
or U4419 (N_4419,N_2575,N_2430);
nand U4420 (N_4420,N_2665,N_3954);
nor U4421 (N_4421,N_2237,N_2536);
nand U4422 (N_4422,N_2991,N_2243);
xnor U4423 (N_4423,N_2165,N_3809);
xor U4424 (N_4424,N_2246,N_2649);
nor U4425 (N_4425,N_2934,N_2995);
nor U4426 (N_4426,N_3073,N_2158);
xnor U4427 (N_4427,N_2447,N_2609);
xor U4428 (N_4428,N_2124,N_3521);
nand U4429 (N_4429,N_3134,N_3537);
or U4430 (N_4430,N_2741,N_3947);
xor U4431 (N_4431,N_3079,N_3087);
nand U4432 (N_4432,N_3028,N_3660);
nor U4433 (N_4433,N_2968,N_2157);
or U4434 (N_4434,N_2435,N_3202);
nor U4435 (N_4435,N_3484,N_3665);
nand U4436 (N_4436,N_2390,N_2606);
and U4437 (N_4437,N_2659,N_3275);
nor U4438 (N_4438,N_2548,N_3456);
or U4439 (N_4439,N_2297,N_2259);
or U4440 (N_4440,N_3815,N_3544);
or U4441 (N_4441,N_2060,N_2180);
or U4442 (N_4442,N_3172,N_2780);
nor U4443 (N_4443,N_2282,N_3247);
nand U4444 (N_4444,N_2545,N_3934);
and U4445 (N_4445,N_3229,N_2269);
nor U4446 (N_4446,N_3356,N_2911);
nor U4447 (N_4447,N_3221,N_3418);
nand U4448 (N_4448,N_3179,N_3300);
nand U4449 (N_4449,N_2776,N_3764);
nor U4450 (N_4450,N_3580,N_2501);
and U4451 (N_4451,N_3350,N_3848);
xnor U4452 (N_4452,N_3500,N_3548);
or U4453 (N_4453,N_2663,N_2479);
nand U4454 (N_4454,N_2797,N_2207);
nor U4455 (N_4455,N_3153,N_2515);
or U4456 (N_4456,N_2569,N_2056);
and U4457 (N_4457,N_3731,N_3326);
nand U4458 (N_4458,N_2680,N_2372);
xor U4459 (N_4459,N_3679,N_3053);
and U4460 (N_4460,N_2519,N_2284);
or U4461 (N_4461,N_3045,N_3622);
nand U4462 (N_4462,N_2290,N_2781);
nand U4463 (N_4463,N_3653,N_2945);
and U4464 (N_4464,N_2292,N_3161);
and U4465 (N_4465,N_3353,N_2556);
nor U4466 (N_4466,N_3596,N_3540);
or U4467 (N_4467,N_3533,N_3265);
or U4468 (N_4468,N_2661,N_3589);
nor U4469 (N_4469,N_3695,N_2929);
and U4470 (N_4470,N_2384,N_2494);
or U4471 (N_4471,N_2582,N_3817);
or U4472 (N_4472,N_3331,N_3688);
and U4473 (N_4473,N_3245,N_2258);
and U4474 (N_4474,N_2364,N_3026);
or U4475 (N_4475,N_3841,N_3063);
and U4476 (N_4476,N_3032,N_3803);
or U4477 (N_4477,N_2108,N_2484);
xor U4478 (N_4478,N_2460,N_2457);
nor U4479 (N_4479,N_3768,N_3074);
nor U4480 (N_4480,N_2424,N_2496);
nand U4481 (N_4481,N_3703,N_2254);
or U4482 (N_4482,N_3060,N_3573);
nor U4483 (N_4483,N_3453,N_3661);
or U4484 (N_4484,N_2089,N_2745);
nor U4485 (N_4485,N_3667,N_2967);
or U4486 (N_4486,N_2355,N_3217);
xor U4487 (N_4487,N_2959,N_3847);
xnor U4488 (N_4488,N_3871,N_2981);
nor U4489 (N_4489,N_3798,N_3228);
or U4490 (N_4490,N_3147,N_3319);
nand U4491 (N_4491,N_3603,N_2340);
or U4492 (N_4492,N_3910,N_3933);
and U4493 (N_4493,N_2462,N_3915);
nand U4494 (N_4494,N_3515,N_2652);
xnor U4495 (N_4495,N_3198,N_3916);
and U4496 (N_4496,N_3818,N_2785);
xnor U4497 (N_4497,N_3957,N_3913);
nand U4498 (N_4498,N_2508,N_3644);
xor U4499 (N_4499,N_3289,N_2011);
nor U4500 (N_4500,N_2866,N_3046);
and U4501 (N_4501,N_2919,N_2010);
nand U4502 (N_4502,N_3083,N_3638);
or U4503 (N_4503,N_3672,N_2674);
nor U4504 (N_4504,N_2746,N_2879);
and U4505 (N_4505,N_3586,N_2889);
xnor U4506 (N_4506,N_2809,N_3485);
and U4507 (N_4507,N_2755,N_3214);
xnor U4508 (N_4508,N_2039,N_2034);
or U4509 (N_4509,N_2480,N_2006);
nor U4510 (N_4510,N_2300,N_2055);
and U4511 (N_4511,N_3287,N_3779);
xor U4512 (N_4512,N_3394,N_2492);
nand U4513 (N_4513,N_2574,N_3057);
nand U4514 (N_4514,N_3493,N_3222);
nor U4515 (N_4515,N_2193,N_3782);
xor U4516 (N_4516,N_2209,N_2647);
nor U4517 (N_4517,N_3967,N_2473);
or U4518 (N_4518,N_3752,N_3896);
nand U4519 (N_4519,N_3117,N_3673);
and U4520 (N_4520,N_3943,N_2099);
and U4521 (N_4521,N_3367,N_2004);
nand U4522 (N_4522,N_3595,N_3006);
nor U4523 (N_4523,N_3587,N_3797);
or U4524 (N_4524,N_3270,N_2817);
xnor U4525 (N_4525,N_3064,N_2795);
nand U4526 (N_4526,N_3778,N_2425);
nor U4527 (N_4527,N_2098,N_3165);
nor U4528 (N_4528,N_2436,N_2708);
nor U4529 (N_4529,N_3027,N_2442);
nand U4530 (N_4530,N_2311,N_3844);
nand U4531 (N_4531,N_2453,N_2383);
or U4532 (N_4532,N_2749,N_2465);
or U4533 (N_4533,N_2940,N_2398);
nor U4534 (N_4534,N_2632,N_2888);
xor U4535 (N_4535,N_2855,N_3744);
nor U4536 (N_4536,N_2315,N_2638);
nor U4537 (N_4537,N_2729,N_2023);
and U4538 (N_4538,N_2846,N_2504);
or U4539 (N_4539,N_3235,N_3175);
and U4540 (N_4540,N_3417,N_2077);
and U4541 (N_4541,N_2012,N_3819);
xnor U4542 (N_4542,N_2349,N_3459);
nor U4543 (N_4543,N_2974,N_2009);
nor U4544 (N_4544,N_3433,N_2567);
or U4545 (N_4545,N_3041,N_3909);
xor U4546 (N_4546,N_2830,N_3467);
and U4547 (N_4547,N_3009,N_3067);
xor U4548 (N_4548,N_2872,N_3282);
xor U4549 (N_4549,N_3628,N_2859);
xnor U4550 (N_4550,N_3240,N_2028);
or U4551 (N_4551,N_2660,N_2192);
nand U4552 (N_4552,N_2762,N_2211);
nand U4553 (N_4553,N_2378,N_2718);
nor U4554 (N_4554,N_3570,N_3670);
nand U4555 (N_4555,N_2377,N_2408);
nand U4556 (N_4556,N_3663,N_3236);
nand U4557 (N_4557,N_2324,N_3446);
nand U4558 (N_4558,N_2342,N_3992);
or U4559 (N_4559,N_2189,N_3690);
and U4560 (N_4560,N_2142,N_3042);
or U4561 (N_4561,N_3262,N_3366);
or U4562 (N_4562,N_3156,N_2524);
nand U4563 (N_4563,N_3513,N_3825);
or U4564 (N_4564,N_2633,N_3969);
or U4565 (N_4565,N_2201,N_3151);
nor U4566 (N_4566,N_2490,N_2730);
xor U4567 (N_4567,N_3642,N_2514);
nor U4568 (N_4568,N_3381,N_3416);
and U4569 (N_4569,N_2437,N_2141);
or U4570 (N_4570,N_2775,N_2043);
xor U4571 (N_4571,N_3127,N_3508);
nand U4572 (N_4572,N_3736,N_2285);
nor U4573 (N_4573,N_3310,N_2069);
nor U4574 (N_4574,N_2172,N_2100);
and U4575 (N_4575,N_3023,N_2102);
xnor U4576 (N_4576,N_2230,N_2067);
and U4577 (N_4577,N_2405,N_2973);
xnor U4578 (N_4578,N_2458,N_2733);
xnor U4579 (N_4579,N_3950,N_2678);
nor U4580 (N_4580,N_2832,N_3955);
and U4581 (N_4581,N_2092,N_3321);
or U4582 (N_4582,N_2503,N_2032);
and U4583 (N_4583,N_3208,N_3551);
or U4584 (N_4584,N_2291,N_3854);
or U4585 (N_4585,N_2987,N_3354);
and U4586 (N_4586,N_3971,N_3216);
xor U4587 (N_4587,N_2353,N_2610);
xnor U4588 (N_4588,N_3685,N_2976);
nand U4589 (N_4589,N_2154,N_3112);
nand U4590 (N_4590,N_3614,N_2169);
nand U4591 (N_4591,N_3952,N_2368);
and U4592 (N_4592,N_3883,N_2298);
or U4593 (N_4593,N_2668,N_3822);
and U4594 (N_4594,N_3256,N_2295);
nor U4595 (N_4595,N_2624,N_2823);
xnor U4596 (N_4596,N_2654,N_3542);
and U4597 (N_4597,N_2724,N_2328);
nor U4598 (N_4598,N_2975,N_2922);
nand U4599 (N_4599,N_3371,N_3912);
xor U4600 (N_4600,N_2455,N_3714);
nand U4601 (N_4601,N_3802,N_2939);
or U4602 (N_4602,N_3146,N_3168);
xor U4603 (N_4603,N_2697,N_2137);
xnor U4604 (N_4604,N_3011,N_2577);
nor U4605 (N_4605,N_2792,N_2323);
nor U4606 (N_4606,N_3048,N_2320);
nor U4607 (N_4607,N_3810,N_2116);
and U4608 (N_4608,N_3939,N_3054);
xor U4609 (N_4609,N_3015,N_2726);
xor U4610 (N_4610,N_3531,N_3873);
and U4611 (N_4611,N_2093,N_3092);
or U4612 (N_4612,N_2418,N_3439);
xnor U4613 (N_4613,N_3776,N_3238);
xor U4614 (N_4614,N_2870,N_2860);
and U4615 (N_4615,N_2672,N_2793);
and U4616 (N_4616,N_2880,N_3643);
xor U4617 (N_4617,N_3274,N_3979);
or U4618 (N_4618,N_3721,N_3692);
nand U4619 (N_4619,N_2030,N_3273);
nor U4620 (N_4620,N_3949,N_3044);
or U4621 (N_4621,N_2957,N_3213);
nand U4622 (N_4622,N_2920,N_2800);
or U4623 (N_4623,N_2586,N_2265);
and U4624 (N_4624,N_3647,N_2216);
or U4625 (N_4625,N_2226,N_3532);
or U4626 (N_4626,N_2965,N_2694);
nand U4627 (N_4627,N_2140,N_3423);
xnor U4628 (N_4628,N_2666,N_2725);
nand U4629 (N_4629,N_3488,N_2409);
nor U4630 (N_4630,N_2932,N_3856);
and U4631 (N_4631,N_2796,N_2167);
and U4632 (N_4632,N_3329,N_2561);
or U4633 (N_4633,N_3777,N_2411);
and U4634 (N_4634,N_3598,N_2513);
nand U4635 (N_4635,N_2200,N_2520);
xor U4636 (N_4636,N_3577,N_2710);
and U4637 (N_4637,N_3512,N_3593);
or U4638 (N_4638,N_3257,N_2493);
xnor U4639 (N_4639,N_2822,N_2065);
nor U4640 (N_4640,N_3958,N_2358);
and U4641 (N_4641,N_3696,N_3155);
and U4642 (N_4642,N_2630,N_3171);
nor U4643 (N_4643,N_3339,N_3592);
nand U4644 (N_4644,N_3180,N_3458);
nor U4645 (N_4645,N_3620,N_3504);
nor U4646 (N_4646,N_3292,N_2537);
and U4647 (N_4647,N_2076,N_3254);
nand U4648 (N_4648,N_3299,N_2898);
or U4649 (N_4649,N_2509,N_2639);
or U4650 (N_4650,N_3824,N_3239);
and U4651 (N_4651,N_3014,N_2637);
or U4652 (N_4652,N_2683,N_3681);
or U4653 (N_4653,N_3506,N_2897);
or U4654 (N_4654,N_3775,N_3602);
nor U4655 (N_4655,N_2591,N_3343);
and U4656 (N_4656,N_3960,N_3650);
nand U4657 (N_4657,N_3445,N_3000);
nor U4658 (N_4658,N_2705,N_2359);
nand U4659 (N_4659,N_2517,N_2926);
nand U4660 (N_4660,N_3931,N_3995);
nor U4661 (N_4661,N_2553,N_2266);
nor U4662 (N_4662,N_2224,N_2716);
and U4663 (N_4663,N_3784,N_3342);
nor U4664 (N_4664,N_3332,N_2419);
and U4665 (N_4665,N_2332,N_2264);
xnor U4666 (N_4666,N_2608,N_2212);
and U4667 (N_4667,N_3702,N_2422);
nand U4668 (N_4668,N_3286,N_3993);
and U4669 (N_4669,N_3503,N_3940);
nor U4670 (N_4670,N_3496,N_2000);
nor U4671 (N_4671,N_3434,N_3557);
and U4672 (N_4672,N_3541,N_3495);
nor U4673 (N_4673,N_2525,N_2064);
nand U4674 (N_4674,N_3774,N_2634);
nor U4675 (N_4675,N_2299,N_3193);
xnor U4676 (N_4676,N_2451,N_2825);
xnor U4677 (N_4677,N_2691,N_3858);
xor U4678 (N_4678,N_3599,N_3036);
and U4679 (N_4679,N_2174,N_2670);
or U4680 (N_4680,N_3093,N_2022);
nand U4681 (N_4681,N_3397,N_3761);
or U4682 (N_4682,N_2512,N_2924);
and U4683 (N_4683,N_3298,N_3828);
xor U4684 (N_4684,N_3167,N_3936);
and U4685 (N_4685,N_3203,N_2806);
nor U4686 (N_4686,N_3271,N_2423);
and U4687 (N_4687,N_2858,N_2523);
xnor U4688 (N_4688,N_2612,N_3384);
and U4689 (N_4689,N_2943,N_3043);
nor U4690 (N_4690,N_3293,N_3231);
nand U4691 (N_4691,N_2615,N_2751);
or U4692 (N_4692,N_2868,N_2072);
or U4693 (N_4693,N_2834,N_2402);
nand U4694 (N_4694,N_3806,N_2601);
xnor U4695 (N_4695,N_2038,N_3430);
nand U4696 (N_4696,N_2260,N_2414);
or U4697 (N_4697,N_2184,N_3796);
nor U4698 (N_4698,N_3075,N_3466);
or U4699 (N_4699,N_2841,N_2908);
and U4700 (N_4700,N_2563,N_2497);
xor U4701 (N_4701,N_2190,N_3526);
and U4702 (N_4702,N_2127,N_2374);
and U4703 (N_4703,N_2936,N_3490);
nor U4704 (N_4704,N_2433,N_2983);
nand U4705 (N_4705,N_3314,N_2478);
nor U4706 (N_4706,N_2223,N_3142);
and U4707 (N_4707,N_3555,N_2094);
and U4708 (N_4708,N_3344,N_2476);
nand U4709 (N_4709,N_2626,N_2048);
or U4710 (N_4710,N_2527,N_2843);
and U4711 (N_4711,N_3437,N_3327);
nor U4712 (N_4712,N_3699,N_2617);
xnor U4713 (N_4713,N_2819,N_2727);
nand U4714 (N_4714,N_2728,N_3543);
nand U4715 (N_4715,N_3793,N_3086);
nor U4716 (N_4716,N_2887,N_2676);
or U4717 (N_4717,N_2219,N_3069);
xnor U4718 (N_4718,N_3177,N_2404);
and U4719 (N_4719,N_2876,N_2229);
or U4720 (N_4720,N_3852,N_3975);
nor U4721 (N_4721,N_2222,N_3553);
nor U4722 (N_4722,N_2773,N_2510);
nand U4723 (N_4723,N_3315,N_2798);
xnor U4724 (N_4724,N_3268,N_3633);
nand U4725 (N_4725,N_3460,N_3392);
nand U4726 (N_4726,N_2985,N_2296);
nand U4727 (N_4727,N_2327,N_3413);
xnor U4728 (N_4728,N_2107,N_3251);
nor U4729 (N_4729,N_3732,N_2829);
or U4730 (N_4730,N_3629,N_2821);
and U4731 (N_4731,N_3639,N_3428);
nor U4732 (N_4732,N_2456,N_3291);
nor U4733 (N_4733,N_3626,N_2445);
xnor U4734 (N_4734,N_2913,N_3522);
or U4735 (N_4735,N_3837,N_3182);
and U4736 (N_4736,N_2803,N_3455);
xor U4737 (N_4737,N_3230,N_2956);
nor U4738 (N_4738,N_3126,N_3637);
nor U4739 (N_4739,N_2952,N_2813);
nand U4740 (N_4740,N_3410,N_3729);
and U4741 (N_4741,N_3659,N_3865);
and U4742 (N_4742,N_3811,N_2472);
or U4743 (N_4743,N_2588,N_3509);
and U4744 (N_4744,N_2218,N_2592);
xnor U4745 (N_4745,N_2018,N_2894);
and U4746 (N_4746,N_3263,N_3110);
nand U4747 (N_4747,N_3489,N_2135);
and U4748 (N_4748,N_3477,N_2281);
or U4749 (N_4749,N_2247,N_3861);
or U4750 (N_4750,N_3449,N_3012);
nand U4751 (N_4751,N_2131,N_2953);
xor U4752 (N_4752,N_3564,N_3020);
nor U4753 (N_4753,N_3680,N_3052);
and U4754 (N_4754,N_3549,N_3741);
or U4755 (N_4755,N_3838,N_3420);
nand U4756 (N_4756,N_3128,N_3615);
or U4757 (N_4757,N_2428,N_3623);
nor U4758 (N_4758,N_3652,N_2168);
xnor U4759 (N_4759,N_3625,N_3107);
or U4760 (N_4760,N_2392,N_2756);
nand U4761 (N_4761,N_2641,N_2204);
nor U4762 (N_4762,N_3498,N_2931);
nand U4763 (N_4763,N_2278,N_2289);
nor U4764 (N_4764,N_2024,N_2961);
xnor U4765 (N_4765,N_3678,N_2925);
or U4766 (N_4766,N_2583,N_2075);
xnor U4767 (N_4767,N_3438,N_2214);
nand U4768 (N_4768,N_3554,N_3461);
xor U4769 (N_4769,N_3547,N_3276);
nor U4770 (N_4770,N_3457,N_3656);
and U4771 (N_4771,N_2596,N_2017);
and U4772 (N_4772,N_2650,N_3094);
or U4773 (N_4773,N_3607,N_2143);
nand U4774 (N_4774,N_3511,N_3051);
and U4775 (N_4775,N_2403,N_2955);
nand U4776 (N_4776,N_2183,N_3738);
or U4777 (N_4777,N_3219,N_3991);
nand U4778 (N_4778,N_3977,N_3415);
nor U4779 (N_4779,N_3382,N_2910);
nor U4780 (N_4780,N_2057,N_2604);
nor U4781 (N_4781,N_3823,N_2948);
and U4782 (N_4782,N_3726,N_3964);
nand U4783 (N_4783,N_3843,N_2095);
or U4784 (N_4784,N_3609,N_2191);
nand U4785 (N_4785,N_2432,N_2857);
nand U4786 (N_4786,N_2485,N_2273);
or U4787 (N_4787,N_3211,N_3102);
and U4788 (N_4788,N_2867,N_2707);
xor U4789 (N_4789,N_2546,N_3707);
nand U4790 (N_4790,N_3984,N_3163);
or U4791 (N_4791,N_2380,N_3974);
xnor U4792 (N_4792,N_3309,N_2787);
or U4793 (N_4793,N_3885,N_2522);
and U4794 (N_4794,N_3566,N_2333);
or U4795 (N_4795,N_2293,N_2551);
nor U4796 (N_4796,N_2186,N_3654);
or U4797 (N_4797,N_2176,N_2971);
xnor U4798 (N_4798,N_3581,N_2042);
nor U4799 (N_4799,N_3771,N_2794);
nor U4800 (N_4800,N_2303,N_2343);
nand U4801 (N_4801,N_3396,N_3864);
or U4802 (N_4802,N_3567,N_2620);
nor U4803 (N_4803,N_2335,N_2679);
xor U4804 (N_4804,N_2766,N_2655);
and U4805 (N_4805,N_3582,N_2388);
nor U4806 (N_4806,N_3426,N_3474);
nand U4807 (N_4807,N_2274,N_3432);
nand U4808 (N_4808,N_2206,N_2877);
or U4809 (N_4809,N_2365,N_3996);
nand U4810 (N_4810,N_2106,N_2044);
nor U4811 (N_4811,N_2602,N_3827);
xor U4812 (N_4812,N_2549,N_2152);
xnor U4813 (N_4813,N_2646,N_2540);
or U4814 (N_4814,N_2241,N_3791);
and U4815 (N_4815,N_3322,N_3636);
or U4816 (N_4816,N_3255,N_2162);
or U4817 (N_4817,N_3260,N_2942);
nor U4818 (N_4818,N_3183,N_2126);
nor U4819 (N_4819,N_2101,N_3903);
nor U4820 (N_4820,N_3982,N_2903);
and U4821 (N_4821,N_3152,N_2103);
and U4822 (N_4822,N_2534,N_3905);
or U4823 (N_4823,N_2317,N_3279);
nor U4824 (N_4824,N_3131,N_2382);
nand U4825 (N_4825,N_2301,N_2376);
xnor U4826 (N_4826,N_3662,N_3900);
nand U4827 (N_4827,N_3040,N_2182);
xor U4828 (N_4828,N_2786,N_2007);
nand U4829 (N_4829,N_2082,N_2709);
or U4830 (N_4830,N_3347,N_3853);
and U4831 (N_4831,N_2863,N_3624);
nand U4832 (N_4832,N_2909,N_3068);
nor U4833 (N_4833,N_2837,N_2393);
and U4834 (N_4834,N_3312,N_3558);
or U4835 (N_4835,N_2063,N_2181);
or U4836 (N_4836,N_2804,N_2314);
or U4837 (N_4837,N_3959,N_3880);
or U4838 (N_4838,N_2272,N_3081);
xnor U4839 (N_4839,N_2849,N_3677);
xnor U4840 (N_4840,N_2963,N_2644);
xnor U4841 (N_4841,N_2603,N_3351);
xor U4842 (N_4842,N_3091,N_3070);
nand U4843 (N_4843,N_3985,N_3528);
nand U4844 (N_4844,N_3233,N_3442);
or U4845 (N_4845,N_3787,N_2271);
nand U4846 (N_4846,N_3205,N_3874);
nand U4847 (N_4847,N_3400,N_3424);
or U4848 (N_4848,N_3826,N_3753);
nand U4849 (N_4849,N_3700,N_3451);
and U4850 (N_4850,N_2970,N_3376);
nand U4851 (N_4851,N_3387,N_2928);
nand U4852 (N_4852,N_2117,N_2815);
or U4853 (N_4853,N_2466,N_3444);
and U4854 (N_4854,N_2706,N_3099);
xor U4855 (N_4855,N_3372,N_2040);
nor U4856 (N_4856,N_3525,N_2906);
nand U4857 (N_4857,N_2921,N_2964);
nand U4858 (N_4858,N_2767,N_2899);
nand U4859 (N_4859,N_2890,N_2499);
xor U4860 (N_4860,N_2687,N_3346);
xnor U4861 (N_4861,N_3898,N_2370);
or U4862 (N_4862,N_2912,N_2461);
or U4863 (N_4863,N_2531,N_3781);
nand U4864 (N_4864,N_2688,N_3664);
xnor U4865 (N_4865,N_2027,N_2426);
or U4866 (N_4866,N_2144,N_3529);
xor U4867 (N_4867,N_2321,N_2836);
and U4868 (N_4868,N_2597,N_3337);
and U4869 (N_4869,N_3762,N_3468);
nand U4870 (N_4870,N_3204,N_2217);
nand U4871 (N_4871,N_3600,N_2146);
or U4872 (N_4872,N_3546,N_2579);
or U4873 (N_4873,N_3946,N_2156);
and U4874 (N_4874,N_3860,N_3887);
xor U4875 (N_4875,N_3431,N_3464);
and U4876 (N_4876,N_2351,N_2248);
and U4877 (N_4877,N_2713,N_2882);
nor U4878 (N_4878,N_3320,N_2053);
xor U4879 (N_4879,N_3693,N_3059);
nand U4880 (N_4880,N_2737,N_2013);
xnor U4881 (N_4881,N_3999,N_2420);
or U4882 (N_4882,N_2873,N_2029);
and U4883 (N_4883,N_2996,N_2225);
nor U4884 (N_4884,N_3748,N_2173);
xnor U4885 (N_4885,N_2220,N_3669);
xnor U4886 (N_4886,N_3085,N_2088);
and U4887 (N_4887,N_3502,N_3994);
and U4888 (N_4888,N_3224,N_3302);
nor U4889 (N_4889,N_3100,N_2779);
xor U4890 (N_4890,N_2673,N_2997);
or U4891 (N_4891,N_3836,N_3821);
nor U4892 (N_4892,N_2395,N_2712);
nand U4893 (N_4893,N_3922,N_3888);
and U4894 (N_4894,N_2938,N_2685);
or U4895 (N_4895,N_3527,N_3941);
or U4896 (N_4896,N_3103,N_3429);
or U4897 (N_4897,N_2276,N_2232);
nand U4898 (N_4898,N_3281,N_3897);
nand U4899 (N_4899,N_2761,N_3184);
xnor U4900 (N_4900,N_3583,N_3763);
nand U4901 (N_4901,N_3482,N_2530);
nor U4902 (N_4902,N_2625,N_3945);
and U4903 (N_4903,N_3022,N_2526);
nor U4904 (N_4904,N_3879,N_2854);
xnor U4905 (N_4905,N_2572,N_3374);
nand U4906 (N_4906,N_2533,N_3333);
xnor U4907 (N_4907,N_2488,N_2818);
and U4908 (N_4908,N_2684,N_2576);
or U4909 (N_4909,N_2074,N_3766);
nand U4910 (N_4910,N_3375,N_2941);
xor U4911 (N_4911,N_3767,N_3632);
nand U4912 (N_4912,N_3377,N_2864);
nand U4913 (N_4913,N_3927,N_2808);
nand U4914 (N_4914,N_3019,N_3352);
or U4915 (N_4915,N_3988,N_2753);
or U4916 (N_4916,N_2757,N_3487);
and U4917 (N_4917,N_3956,N_3095);
and U4918 (N_4918,N_2657,N_3645);
nor U4919 (N_4919,N_2306,N_3783);
nor U4920 (N_4920,N_3813,N_2636);
xor U4921 (N_4921,N_3148,N_3937);
xor U4922 (N_4922,N_3116,N_2698);
xor U4923 (N_4923,N_2371,N_2690);
nor U4924 (N_4924,N_3606,N_3452);
and U4925 (N_4925,N_3109,N_2133);
or U4926 (N_4926,N_3840,N_2986);
xor U4927 (N_4927,N_3608,N_3902);
xnor U4928 (N_4928,N_3833,N_2669);
nor U4929 (N_4929,N_2449,N_2035);
or U4930 (N_4930,N_3308,N_3261);
nand U4931 (N_4931,N_3530,N_2341);
nand U4932 (N_4932,N_2607,N_2431);
xnor U4933 (N_4933,N_2086,N_3010);
or U4934 (N_4934,N_3935,N_3301);
or U4935 (N_4935,N_3218,N_2338);
nand U4936 (N_4936,N_3720,N_2946);
nand U4937 (N_4937,N_3772,N_2429);
and U4938 (N_4938,N_2352,N_3242);
nand U4939 (N_4939,N_2771,N_2883);
nor U4940 (N_4940,N_3743,N_2736);
or U4941 (N_4941,N_3304,N_2573);
xor U4942 (N_4942,N_3568,N_2283);
nor U4943 (N_4943,N_3227,N_3145);
xor U4944 (N_4944,N_2361,N_2163);
and U4945 (N_4945,N_3691,N_3611);
xnor U4946 (N_4946,N_2578,N_3137);
nor U4947 (N_4947,N_2356,N_3189);
nand U4948 (N_4948,N_3004,N_3476);
nor U4949 (N_4949,N_3907,N_2360);
and U4950 (N_4950,N_3758,N_3835);
nand U4951 (N_4951,N_2770,N_2084);
or U4952 (N_4952,N_2459,N_2989);
or U4953 (N_4953,N_3215,N_2199);
nand U4954 (N_4954,N_2046,N_2789);
xor U4955 (N_4955,N_3917,N_3968);
or U4956 (N_4956,N_3682,N_3349);
xnor U4957 (N_4957,N_3734,N_3538);
xnor U4958 (N_4958,N_3077,N_2507);
or U4959 (N_4959,N_2339,N_3565);
and U4960 (N_4960,N_3863,N_3715);
and U4961 (N_4961,N_3584,N_2902);
nor U4962 (N_4962,N_3501,N_3050);
nand U4963 (N_4963,N_2326,N_3801);
and U4964 (N_4964,N_3370,N_3317);
nor U4965 (N_4965,N_2454,N_3098);
nor U4966 (N_4966,N_2136,N_3159);
and U4967 (N_4967,N_3892,N_3348);
nand U4968 (N_4968,N_3745,N_2050);
xor U4969 (N_4969,N_2988,N_2188);
or U4970 (N_4970,N_2073,N_2196);
xor U4971 (N_4971,N_3872,N_2438);
or U4972 (N_4972,N_2170,N_3588);
or U4973 (N_4973,N_3139,N_2842);
and U4974 (N_4974,N_3990,N_3226);
nand U4975 (N_4975,N_3612,N_2875);
xor U4976 (N_4976,N_2240,N_2907);
and U4977 (N_4977,N_3259,N_2052);
or U4978 (N_4978,N_3560,N_2831);
or U4979 (N_4979,N_3388,N_2850);
xnor U4980 (N_4980,N_3832,N_2671);
nor U4981 (N_4981,N_2440,N_2130);
or U4982 (N_4982,N_3891,N_3435);
nand U4983 (N_4983,N_2114,N_2764);
nand U4984 (N_4984,N_3920,N_2014);
or U4985 (N_4985,N_2003,N_2543);
nor U4986 (N_4986,N_3129,N_3210);
and U4987 (N_4987,N_3454,N_3849);
or U4988 (N_4988,N_3746,N_3136);
nand U4989 (N_4989,N_2722,N_3480);
nor U4990 (N_4990,N_3097,N_3904);
or U4991 (N_4991,N_2653,N_3505);
and U4992 (N_4992,N_3395,N_2595);
and U4993 (N_4993,N_3365,N_2711);
nor U4994 (N_4994,N_2944,N_3705);
nand U4995 (N_4995,N_2714,N_3448);
xnor U4996 (N_4996,N_3562,N_2623);
xnor U4997 (N_4997,N_2571,N_3942);
nor U4998 (N_4998,N_2036,N_3627);
or U4999 (N_4999,N_3510,N_2681);
and U5000 (N_5000,N_3949,N_3711);
xor U5001 (N_5001,N_2666,N_3283);
nand U5002 (N_5002,N_2425,N_2867);
and U5003 (N_5003,N_2186,N_2944);
nor U5004 (N_5004,N_2865,N_3864);
xor U5005 (N_5005,N_2847,N_3095);
or U5006 (N_5006,N_2360,N_2487);
nor U5007 (N_5007,N_2614,N_2665);
nor U5008 (N_5008,N_3940,N_2090);
and U5009 (N_5009,N_3798,N_2011);
or U5010 (N_5010,N_2323,N_3826);
or U5011 (N_5011,N_2869,N_2605);
xor U5012 (N_5012,N_2932,N_3974);
nand U5013 (N_5013,N_3905,N_3017);
or U5014 (N_5014,N_3192,N_2876);
xnor U5015 (N_5015,N_2770,N_3030);
and U5016 (N_5016,N_3916,N_3523);
nand U5017 (N_5017,N_3102,N_2887);
nand U5018 (N_5018,N_2377,N_3188);
and U5019 (N_5019,N_2355,N_2482);
nand U5020 (N_5020,N_3513,N_3132);
nand U5021 (N_5021,N_2411,N_2034);
and U5022 (N_5022,N_3923,N_3719);
xnor U5023 (N_5023,N_2157,N_2082);
xnor U5024 (N_5024,N_3823,N_2426);
nor U5025 (N_5025,N_3077,N_3799);
and U5026 (N_5026,N_2452,N_3937);
nor U5027 (N_5027,N_2362,N_2925);
or U5028 (N_5028,N_2288,N_3344);
or U5029 (N_5029,N_2184,N_2628);
or U5030 (N_5030,N_3646,N_2452);
nand U5031 (N_5031,N_2445,N_3087);
nand U5032 (N_5032,N_3213,N_2717);
nor U5033 (N_5033,N_3903,N_2935);
nor U5034 (N_5034,N_3576,N_2925);
nor U5035 (N_5035,N_2791,N_2752);
and U5036 (N_5036,N_3193,N_3966);
or U5037 (N_5037,N_2474,N_2007);
and U5038 (N_5038,N_2661,N_2785);
nor U5039 (N_5039,N_3622,N_3946);
or U5040 (N_5040,N_2638,N_2903);
or U5041 (N_5041,N_3408,N_3353);
nor U5042 (N_5042,N_3981,N_3364);
nand U5043 (N_5043,N_3834,N_3205);
nand U5044 (N_5044,N_2019,N_2755);
and U5045 (N_5045,N_2895,N_2251);
nand U5046 (N_5046,N_3227,N_3255);
or U5047 (N_5047,N_3698,N_2125);
nor U5048 (N_5048,N_2838,N_2857);
nor U5049 (N_5049,N_2881,N_2035);
or U5050 (N_5050,N_3656,N_3840);
xor U5051 (N_5051,N_2172,N_3777);
nor U5052 (N_5052,N_2190,N_3273);
nor U5053 (N_5053,N_3029,N_3172);
nand U5054 (N_5054,N_2286,N_3695);
nor U5055 (N_5055,N_2604,N_2971);
or U5056 (N_5056,N_3111,N_3398);
or U5057 (N_5057,N_2512,N_3209);
nor U5058 (N_5058,N_3557,N_3715);
xor U5059 (N_5059,N_3184,N_2250);
or U5060 (N_5060,N_3311,N_2575);
nand U5061 (N_5061,N_3411,N_2288);
or U5062 (N_5062,N_2372,N_3808);
nand U5063 (N_5063,N_3270,N_3141);
or U5064 (N_5064,N_2063,N_3878);
nor U5065 (N_5065,N_2385,N_3663);
nor U5066 (N_5066,N_3148,N_3400);
nor U5067 (N_5067,N_3544,N_3127);
and U5068 (N_5068,N_2303,N_2933);
nor U5069 (N_5069,N_2157,N_3195);
xor U5070 (N_5070,N_3968,N_2503);
and U5071 (N_5071,N_2525,N_2360);
or U5072 (N_5072,N_3683,N_3166);
or U5073 (N_5073,N_2449,N_2913);
or U5074 (N_5074,N_2458,N_3969);
or U5075 (N_5075,N_3135,N_3137);
nor U5076 (N_5076,N_2678,N_2033);
nor U5077 (N_5077,N_2947,N_3533);
nor U5078 (N_5078,N_2770,N_2101);
or U5079 (N_5079,N_3600,N_2182);
xor U5080 (N_5080,N_3014,N_3572);
xnor U5081 (N_5081,N_2650,N_3899);
nor U5082 (N_5082,N_2183,N_3783);
and U5083 (N_5083,N_3632,N_2774);
xor U5084 (N_5084,N_3745,N_2620);
nand U5085 (N_5085,N_3697,N_2761);
nand U5086 (N_5086,N_3210,N_3168);
nor U5087 (N_5087,N_3846,N_3152);
and U5088 (N_5088,N_2870,N_2482);
nand U5089 (N_5089,N_2282,N_2462);
nand U5090 (N_5090,N_2678,N_3587);
nand U5091 (N_5091,N_3451,N_2781);
nor U5092 (N_5092,N_3382,N_2633);
or U5093 (N_5093,N_2372,N_3707);
xnor U5094 (N_5094,N_3057,N_3989);
nor U5095 (N_5095,N_2261,N_2940);
nand U5096 (N_5096,N_3835,N_3714);
or U5097 (N_5097,N_2578,N_3482);
nor U5098 (N_5098,N_3251,N_2891);
xor U5099 (N_5099,N_2773,N_2363);
nor U5100 (N_5100,N_2925,N_3321);
nor U5101 (N_5101,N_3761,N_3814);
nand U5102 (N_5102,N_2487,N_2402);
and U5103 (N_5103,N_2849,N_2002);
nand U5104 (N_5104,N_2392,N_3767);
xor U5105 (N_5105,N_3886,N_3333);
nor U5106 (N_5106,N_2892,N_3619);
xor U5107 (N_5107,N_2066,N_3842);
nor U5108 (N_5108,N_3559,N_3523);
and U5109 (N_5109,N_3201,N_3347);
nor U5110 (N_5110,N_2222,N_3297);
and U5111 (N_5111,N_2139,N_3844);
and U5112 (N_5112,N_3261,N_3511);
nand U5113 (N_5113,N_3234,N_2578);
nand U5114 (N_5114,N_3794,N_3142);
nor U5115 (N_5115,N_3558,N_3716);
nor U5116 (N_5116,N_3551,N_3763);
nor U5117 (N_5117,N_2297,N_2910);
or U5118 (N_5118,N_3704,N_3803);
or U5119 (N_5119,N_2741,N_2525);
nor U5120 (N_5120,N_2538,N_2725);
nor U5121 (N_5121,N_3365,N_3034);
or U5122 (N_5122,N_2154,N_2852);
or U5123 (N_5123,N_2353,N_2703);
or U5124 (N_5124,N_2024,N_2590);
xor U5125 (N_5125,N_3229,N_2303);
or U5126 (N_5126,N_3057,N_2524);
or U5127 (N_5127,N_2767,N_3133);
xor U5128 (N_5128,N_2131,N_3308);
or U5129 (N_5129,N_3258,N_3004);
nor U5130 (N_5130,N_3283,N_3633);
and U5131 (N_5131,N_3401,N_3793);
nor U5132 (N_5132,N_3977,N_2140);
and U5133 (N_5133,N_2513,N_2160);
xnor U5134 (N_5134,N_3565,N_2676);
or U5135 (N_5135,N_2693,N_2191);
xnor U5136 (N_5136,N_2029,N_3316);
nand U5137 (N_5137,N_3857,N_3395);
nor U5138 (N_5138,N_3614,N_2147);
nor U5139 (N_5139,N_3578,N_3501);
nand U5140 (N_5140,N_3628,N_3486);
xnor U5141 (N_5141,N_2418,N_2478);
nor U5142 (N_5142,N_3613,N_3713);
or U5143 (N_5143,N_3699,N_2377);
xnor U5144 (N_5144,N_3380,N_3598);
or U5145 (N_5145,N_3032,N_3636);
nand U5146 (N_5146,N_3895,N_2046);
or U5147 (N_5147,N_3141,N_2077);
and U5148 (N_5148,N_3967,N_2191);
or U5149 (N_5149,N_3470,N_2898);
or U5150 (N_5150,N_2293,N_2974);
nand U5151 (N_5151,N_3216,N_2805);
nor U5152 (N_5152,N_2453,N_3152);
xor U5153 (N_5153,N_2145,N_3160);
nand U5154 (N_5154,N_2200,N_2789);
nor U5155 (N_5155,N_2618,N_2984);
nand U5156 (N_5156,N_3985,N_2244);
nand U5157 (N_5157,N_2916,N_2433);
nor U5158 (N_5158,N_3515,N_2528);
nand U5159 (N_5159,N_2489,N_2834);
or U5160 (N_5160,N_2665,N_2071);
xor U5161 (N_5161,N_3328,N_3590);
nor U5162 (N_5162,N_2661,N_3533);
nand U5163 (N_5163,N_2660,N_3539);
xor U5164 (N_5164,N_2067,N_3260);
nor U5165 (N_5165,N_2318,N_2986);
nand U5166 (N_5166,N_2538,N_2636);
and U5167 (N_5167,N_3086,N_3448);
and U5168 (N_5168,N_3402,N_2185);
nand U5169 (N_5169,N_2825,N_2689);
and U5170 (N_5170,N_2277,N_3829);
nand U5171 (N_5171,N_3130,N_3110);
and U5172 (N_5172,N_2302,N_3887);
and U5173 (N_5173,N_3258,N_2203);
and U5174 (N_5174,N_2886,N_3586);
and U5175 (N_5175,N_2217,N_3246);
xor U5176 (N_5176,N_2722,N_2534);
and U5177 (N_5177,N_2114,N_3530);
and U5178 (N_5178,N_3761,N_3206);
and U5179 (N_5179,N_2782,N_3290);
or U5180 (N_5180,N_3383,N_2864);
nand U5181 (N_5181,N_3158,N_3784);
nor U5182 (N_5182,N_2664,N_3293);
or U5183 (N_5183,N_2114,N_3118);
xor U5184 (N_5184,N_2935,N_3526);
nand U5185 (N_5185,N_2323,N_2828);
xnor U5186 (N_5186,N_3180,N_2492);
nand U5187 (N_5187,N_3061,N_3992);
nor U5188 (N_5188,N_3978,N_2563);
nor U5189 (N_5189,N_2414,N_2301);
xor U5190 (N_5190,N_2092,N_3071);
and U5191 (N_5191,N_3178,N_3799);
nand U5192 (N_5192,N_3939,N_2597);
nor U5193 (N_5193,N_2111,N_3022);
xnor U5194 (N_5194,N_3763,N_3441);
xnor U5195 (N_5195,N_3912,N_2779);
xnor U5196 (N_5196,N_3697,N_2149);
and U5197 (N_5197,N_3338,N_3706);
and U5198 (N_5198,N_3069,N_2311);
or U5199 (N_5199,N_2648,N_3805);
nand U5200 (N_5200,N_3863,N_2710);
nand U5201 (N_5201,N_3981,N_2164);
nor U5202 (N_5202,N_2695,N_2948);
xnor U5203 (N_5203,N_2989,N_3902);
nand U5204 (N_5204,N_2864,N_3690);
or U5205 (N_5205,N_3385,N_2044);
xnor U5206 (N_5206,N_3542,N_3464);
nor U5207 (N_5207,N_3027,N_3954);
nor U5208 (N_5208,N_3773,N_2221);
and U5209 (N_5209,N_3581,N_2483);
nor U5210 (N_5210,N_2372,N_2363);
nand U5211 (N_5211,N_3502,N_3934);
xor U5212 (N_5212,N_2745,N_3128);
and U5213 (N_5213,N_2970,N_2671);
nor U5214 (N_5214,N_3951,N_3111);
nor U5215 (N_5215,N_2111,N_2145);
or U5216 (N_5216,N_2719,N_3798);
or U5217 (N_5217,N_3518,N_3411);
nand U5218 (N_5218,N_3593,N_2885);
or U5219 (N_5219,N_2038,N_3891);
and U5220 (N_5220,N_3697,N_2337);
or U5221 (N_5221,N_3440,N_2153);
and U5222 (N_5222,N_3733,N_3920);
nand U5223 (N_5223,N_2487,N_3673);
xnor U5224 (N_5224,N_2318,N_3911);
or U5225 (N_5225,N_3935,N_3975);
xnor U5226 (N_5226,N_3314,N_2956);
and U5227 (N_5227,N_3866,N_3896);
or U5228 (N_5228,N_2415,N_2329);
or U5229 (N_5229,N_3557,N_2448);
xor U5230 (N_5230,N_2122,N_3016);
xnor U5231 (N_5231,N_2036,N_3113);
and U5232 (N_5232,N_3180,N_2468);
or U5233 (N_5233,N_3164,N_2146);
and U5234 (N_5234,N_3417,N_3546);
nor U5235 (N_5235,N_3779,N_2955);
and U5236 (N_5236,N_3997,N_2524);
xor U5237 (N_5237,N_3160,N_2124);
or U5238 (N_5238,N_3946,N_3584);
or U5239 (N_5239,N_3866,N_3084);
nand U5240 (N_5240,N_2072,N_2729);
xnor U5241 (N_5241,N_2731,N_3331);
and U5242 (N_5242,N_3624,N_2870);
and U5243 (N_5243,N_2557,N_3054);
and U5244 (N_5244,N_3013,N_2560);
xnor U5245 (N_5245,N_3170,N_3605);
nor U5246 (N_5246,N_3390,N_2068);
or U5247 (N_5247,N_3019,N_2839);
nor U5248 (N_5248,N_2238,N_2390);
nor U5249 (N_5249,N_2765,N_3518);
nor U5250 (N_5250,N_3467,N_2965);
nand U5251 (N_5251,N_2716,N_2008);
nand U5252 (N_5252,N_3973,N_2010);
and U5253 (N_5253,N_2851,N_3291);
nand U5254 (N_5254,N_2540,N_3970);
or U5255 (N_5255,N_3446,N_3641);
nand U5256 (N_5256,N_2912,N_3421);
xor U5257 (N_5257,N_2637,N_2832);
xnor U5258 (N_5258,N_3540,N_2221);
or U5259 (N_5259,N_2186,N_3899);
nand U5260 (N_5260,N_3368,N_3311);
nor U5261 (N_5261,N_2087,N_3507);
xnor U5262 (N_5262,N_2756,N_2546);
and U5263 (N_5263,N_3284,N_2978);
and U5264 (N_5264,N_3107,N_2156);
and U5265 (N_5265,N_2902,N_2169);
or U5266 (N_5266,N_3182,N_3807);
xor U5267 (N_5267,N_2703,N_2741);
or U5268 (N_5268,N_3830,N_3760);
nand U5269 (N_5269,N_3056,N_2011);
nor U5270 (N_5270,N_3581,N_2517);
nor U5271 (N_5271,N_2150,N_3129);
or U5272 (N_5272,N_2538,N_2079);
nand U5273 (N_5273,N_2154,N_3259);
xor U5274 (N_5274,N_2978,N_2762);
xnor U5275 (N_5275,N_3355,N_2626);
nor U5276 (N_5276,N_3744,N_2052);
nand U5277 (N_5277,N_2002,N_2490);
nand U5278 (N_5278,N_2162,N_3179);
or U5279 (N_5279,N_3693,N_2892);
or U5280 (N_5280,N_3569,N_3171);
nor U5281 (N_5281,N_2119,N_3570);
and U5282 (N_5282,N_3757,N_3476);
and U5283 (N_5283,N_2609,N_3268);
xor U5284 (N_5284,N_3850,N_2528);
nand U5285 (N_5285,N_3168,N_3910);
or U5286 (N_5286,N_2175,N_3772);
or U5287 (N_5287,N_3493,N_2505);
nor U5288 (N_5288,N_2355,N_2233);
nor U5289 (N_5289,N_3286,N_2925);
xor U5290 (N_5290,N_2798,N_3821);
nor U5291 (N_5291,N_3884,N_3306);
or U5292 (N_5292,N_3949,N_2397);
or U5293 (N_5293,N_3506,N_2216);
or U5294 (N_5294,N_2460,N_2352);
or U5295 (N_5295,N_2327,N_2752);
nand U5296 (N_5296,N_2678,N_3779);
xor U5297 (N_5297,N_2303,N_3996);
nand U5298 (N_5298,N_2619,N_3579);
nor U5299 (N_5299,N_2269,N_2572);
or U5300 (N_5300,N_2840,N_2617);
nor U5301 (N_5301,N_2628,N_2787);
nand U5302 (N_5302,N_3496,N_2184);
nor U5303 (N_5303,N_2350,N_3840);
nor U5304 (N_5304,N_2968,N_2929);
nor U5305 (N_5305,N_3621,N_3244);
or U5306 (N_5306,N_2227,N_3791);
or U5307 (N_5307,N_3788,N_2371);
nor U5308 (N_5308,N_3723,N_2613);
xnor U5309 (N_5309,N_3237,N_3487);
or U5310 (N_5310,N_2345,N_3629);
and U5311 (N_5311,N_2867,N_2297);
or U5312 (N_5312,N_3053,N_3060);
nor U5313 (N_5313,N_2327,N_2002);
xor U5314 (N_5314,N_3157,N_3668);
or U5315 (N_5315,N_3627,N_2523);
xor U5316 (N_5316,N_2363,N_2949);
xnor U5317 (N_5317,N_3758,N_3981);
xnor U5318 (N_5318,N_3277,N_2935);
nor U5319 (N_5319,N_2410,N_3564);
nand U5320 (N_5320,N_2950,N_3350);
xor U5321 (N_5321,N_3035,N_3542);
xor U5322 (N_5322,N_3458,N_2420);
xor U5323 (N_5323,N_3949,N_3590);
nor U5324 (N_5324,N_2566,N_3482);
and U5325 (N_5325,N_3737,N_2805);
nor U5326 (N_5326,N_3696,N_2954);
nor U5327 (N_5327,N_2058,N_3761);
or U5328 (N_5328,N_3805,N_2338);
and U5329 (N_5329,N_3062,N_2234);
or U5330 (N_5330,N_2399,N_3466);
nand U5331 (N_5331,N_2914,N_2268);
xnor U5332 (N_5332,N_2955,N_3479);
xnor U5333 (N_5333,N_2054,N_2135);
and U5334 (N_5334,N_3979,N_3629);
or U5335 (N_5335,N_2224,N_3614);
or U5336 (N_5336,N_3384,N_3052);
and U5337 (N_5337,N_2328,N_3066);
or U5338 (N_5338,N_3191,N_2108);
or U5339 (N_5339,N_3540,N_3366);
xor U5340 (N_5340,N_2386,N_2751);
or U5341 (N_5341,N_2817,N_3105);
xor U5342 (N_5342,N_3240,N_2393);
xor U5343 (N_5343,N_2930,N_2158);
nand U5344 (N_5344,N_2316,N_2645);
nand U5345 (N_5345,N_2022,N_2173);
or U5346 (N_5346,N_2884,N_3666);
nor U5347 (N_5347,N_3126,N_3272);
nor U5348 (N_5348,N_2653,N_2113);
nor U5349 (N_5349,N_3271,N_2165);
nand U5350 (N_5350,N_2607,N_2798);
or U5351 (N_5351,N_2970,N_2418);
nor U5352 (N_5352,N_2150,N_3568);
nor U5353 (N_5353,N_2019,N_3652);
or U5354 (N_5354,N_2714,N_2204);
xor U5355 (N_5355,N_2313,N_2036);
xnor U5356 (N_5356,N_2005,N_2747);
and U5357 (N_5357,N_2063,N_2306);
xor U5358 (N_5358,N_3825,N_3493);
nand U5359 (N_5359,N_2648,N_2107);
nand U5360 (N_5360,N_2706,N_3850);
xor U5361 (N_5361,N_3322,N_2334);
xor U5362 (N_5362,N_2421,N_3864);
nor U5363 (N_5363,N_2618,N_2302);
nor U5364 (N_5364,N_3501,N_2047);
nand U5365 (N_5365,N_3451,N_3308);
nor U5366 (N_5366,N_2755,N_3183);
and U5367 (N_5367,N_3887,N_2521);
or U5368 (N_5368,N_3957,N_3113);
and U5369 (N_5369,N_2200,N_2618);
and U5370 (N_5370,N_2164,N_2597);
nor U5371 (N_5371,N_3134,N_3654);
or U5372 (N_5372,N_2333,N_3422);
nor U5373 (N_5373,N_3453,N_2401);
or U5374 (N_5374,N_3394,N_2058);
xor U5375 (N_5375,N_2492,N_3501);
or U5376 (N_5376,N_2031,N_3925);
and U5377 (N_5377,N_2541,N_3999);
nor U5378 (N_5378,N_2843,N_2668);
or U5379 (N_5379,N_2328,N_3872);
nand U5380 (N_5380,N_3858,N_3413);
nor U5381 (N_5381,N_2613,N_3492);
nor U5382 (N_5382,N_3059,N_2384);
or U5383 (N_5383,N_2182,N_2062);
nand U5384 (N_5384,N_3350,N_3110);
nand U5385 (N_5385,N_2857,N_2702);
nor U5386 (N_5386,N_2500,N_3418);
xor U5387 (N_5387,N_3171,N_3994);
and U5388 (N_5388,N_2271,N_2225);
xor U5389 (N_5389,N_3036,N_2941);
xor U5390 (N_5390,N_2237,N_2923);
nor U5391 (N_5391,N_3295,N_2857);
xor U5392 (N_5392,N_3552,N_3054);
or U5393 (N_5393,N_3950,N_2471);
nand U5394 (N_5394,N_3043,N_2269);
or U5395 (N_5395,N_2042,N_3679);
and U5396 (N_5396,N_3453,N_2257);
or U5397 (N_5397,N_2529,N_2393);
xor U5398 (N_5398,N_2918,N_3470);
nand U5399 (N_5399,N_2038,N_2308);
xnor U5400 (N_5400,N_2737,N_3257);
xor U5401 (N_5401,N_3697,N_2867);
or U5402 (N_5402,N_3229,N_3178);
nand U5403 (N_5403,N_3242,N_2528);
and U5404 (N_5404,N_3044,N_2605);
and U5405 (N_5405,N_3233,N_2355);
or U5406 (N_5406,N_2045,N_3734);
xor U5407 (N_5407,N_3633,N_3877);
nor U5408 (N_5408,N_3685,N_3784);
or U5409 (N_5409,N_2833,N_2991);
nand U5410 (N_5410,N_2506,N_2583);
nand U5411 (N_5411,N_3246,N_3979);
xor U5412 (N_5412,N_2853,N_3443);
and U5413 (N_5413,N_2195,N_3119);
nor U5414 (N_5414,N_2641,N_3434);
xor U5415 (N_5415,N_3527,N_2344);
or U5416 (N_5416,N_3828,N_3082);
xor U5417 (N_5417,N_2986,N_2836);
and U5418 (N_5418,N_2663,N_3903);
nand U5419 (N_5419,N_3141,N_3275);
nor U5420 (N_5420,N_2155,N_2469);
nand U5421 (N_5421,N_2848,N_3195);
nand U5422 (N_5422,N_2548,N_2761);
nand U5423 (N_5423,N_2479,N_2871);
or U5424 (N_5424,N_2224,N_3328);
xnor U5425 (N_5425,N_2080,N_2468);
nand U5426 (N_5426,N_3990,N_2995);
nand U5427 (N_5427,N_2962,N_3957);
nor U5428 (N_5428,N_2723,N_2404);
and U5429 (N_5429,N_2850,N_2064);
nor U5430 (N_5430,N_2005,N_2558);
nand U5431 (N_5431,N_3719,N_3119);
nand U5432 (N_5432,N_3364,N_2625);
and U5433 (N_5433,N_2196,N_3145);
xnor U5434 (N_5434,N_2920,N_2303);
nor U5435 (N_5435,N_3821,N_3144);
and U5436 (N_5436,N_2327,N_2786);
nor U5437 (N_5437,N_2612,N_3913);
or U5438 (N_5438,N_2912,N_3989);
nor U5439 (N_5439,N_2230,N_2934);
and U5440 (N_5440,N_3494,N_3078);
or U5441 (N_5441,N_3288,N_2147);
xor U5442 (N_5442,N_3678,N_2365);
and U5443 (N_5443,N_3767,N_2477);
xor U5444 (N_5444,N_3931,N_2600);
xnor U5445 (N_5445,N_3799,N_3327);
or U5446 (N_5446,N_2733,N_2340);
nand U5447 (N_5447,N_2518,N_2410);
xor U5448 (N_5448,N_2275,N_3088);
nor U5449 (N_5449,N_3516,N_2110);
or U5450 (N_5450,N_2274,N_3443);
nor U5451 (N_5451,N_3353,N_2794);
nor U5452 (N_5452,N_2227,N_2823);
and U5453 (N_5453,N_3716,N_3686);
nor U5454 (N_5454,N_3035,N_2519);
and U5455 (N_5455,N_2310,N_2824);
xnor U5456 (N_5456,N_3148,N_2906);
and U5457 (N_5457,N_3246,N_3658);
or U5458 (N_5458,N_2361,N_3310);
nand U5459 (N_5459,N_2619,N_3460);
nand U5460 (N_5460,N_2928,N_2213);
nor U5461 (N_5461,N_2853,N_3043);
nor U5462 (N_5462,N_3903,N_3807);
or U5463 (N_5463,N_3968,N_2771);
and U5464 (N_5464,N_2085,N_3907);
or U5465 (N_5465,N_3217,N_2101);
and U5466 (N_5466,N_3409,N_3948);
nor U5467 (N_5467,N_2493,N_2660);
and U5468 (N_5468,N_3713,N_3650);
nor U5469 (N_5469,N_2843,N_3248);
nand U5470 (N_5470,N_2633,N_2926);
and U5471 (N_5471,N_2906,N_3329);
or U5472 (N_5472,N_3003,N_2654);
or U5473 (N_5473,N_3591,N_2495);
or U5474 (N_5474,N_2286,N_2406);
nand U5475 (N_5475,N_3827,N_2685);
xnor U5476 (N_5476,N_3512,N_2847);
and U5477 (N_5477,N_3172,N_3666);
and U5478 (N_5478,N_3805,N_2993);
xor U5479 (N_5479,N_3614,N_3119);
or U5480 (N_5480,N_3781,N_2355);
xor U5481 (N_5481,N_3240,N_2879);
and U5482 (N_5482,N_2039,N_2529);
nor U5483 (N_5483,N_3918,N_3575);
or U5484 (N_5484,N_2560,N_3927);
nand U5485 (N_5485,N_2893,N_3784);
nand U5486 (N_5486,N_2956,N_2366);
and U5487 (N_5487,N_2378,N_3443);
nand U5488 (N_5488,N_3947,N_3559);
nand U5489 (N_5489,N_2722,N_2824);
nand U5490 (N_5490,N_2870,N_3821);
or U5491 (N_5491,N_3858,N_2084);
and U5492 (N_5492,N_3846,N_2074);
or U5493 (N_5493,N_2667,N_2951);
or U5494 (N_5494,N_2348,N_3312);
or U5495 (N_5495,N_3640,N_2431);
or U5496 (N_5496,N_2694,N_2961);
xnor U5497 (N_5497,N_3792,N_3481);
nor U5498 (N_5498,N_2003,N_3715);
xnor U5499 (N_5499,N_2258,N_2149);
xnor U5500 (N_5500,N_3289,N_2865);
or U5501 (N_5501,N_2538,N_2394);
nand U5502 (N_5502,N_3409,N_3189);
and U5503 (N_5503,N_3920,N_3825);
or U5504 (N_5504,N_2537,N_3901);
or U5505 (N_5505,N_2977,N_2736);
nand U5506 (N_5506,N_2190,N_3240);
and U5507 (N_5507,N_3014,N_2761);
and U5508 (N_5508,N_2562,N_2721);
or U5509 (N_5509,N_3843,N_3182);
xnor U5510 (N_5510,N_3341,N_3925);
or U5511 (N_5511,N_2006,N_3542);
nor U5512 (N_5512,N_2221,N_2554);
nor U5513 (N_5513,N_3824,N_2728);
and U5514 (N_5514,N_3146,N_3576);
nand U5515 (N_5515,N_3062,N_3915);
and U5516 (N_5516,N_3083,N_3946);
and U5517 (N_5517,N_3808,N_3995);
xor U5518 (N_5518,N_2731,N_3596);
nand U5519 (N_5519,N_2223,N_3264);
xnor U5520 (N_5520,N_3724,N_3109);
nand U5521 (N_5521,N_3265,N_2864);
xnor U5522 (N_5522,N_3298,N_3928);
nor U5523 (N_5523,N_2104,N_3103);
xor U5524 (N_5524,N_3467,N_3112);
nand U5525 (N_5525,N_3602,N_3917);
nand U5526 (N_5526,N_3608,N_2347);
xor U5527 (N_5527,N_2044,N_3303);
nand U5528 (N_5528,N_2107,N_2244);
and U5529 (N_5529,N_3210,N_3667);
or U5530 (N_5530,N_3996,N_2105);
nand U5531 (N_5531,N_3736,N_2815);
xor U5532 (N_5532,N_2388,N_2180);
xor U5533 (N_5533,N_3989,N_2613);
or U5534 (N_5534,N_2611,N_2231);
or U5535 (N_5535,N_2987,N_2477);
xor U5536 (N_5536,N_3457,N_2838);
nor U5537 (N_5537,N_2935,N_3425);
xnor U5538 (N_5538,N_3472,N_3284);
xnor U5539 (N_5539,N_3885,N_2958);
nand U5540 (N_5540,N_3045,N_3677);
and U5541 (N_5541,N_3314,N_2459);
nand U5542 (N_5542,N_3874,N_2421);
and U5543 (N_5543,N_2847,N_3368);
xnor U5544 (N_5544,N_2581,N_2820);
and U5545 (N_5545,N_3728,N_3592);
nor U5546 (N_5546,N_2316,N_3692);
xor U5547 (N_5547,N_3274,N_2321);
xnor U5548 (N_5548,N_3478,N_3549);
nor U5549 (N_5549,N_2668,N_2580);
xor U5550 (N_5550,N_2962,N_3144);
nand U5551 (N_5551,N_2466,N_2903);
xor U5552 (N_5552,N_3532,N_2652);
xnor U5553 (N_5553,N_2334,N_2818);
and U5554 (N_5554,N_2612,N_2015);
nand U5555 (N_5555,N_3182,N_3009);
nand U5556 (N_5556,N_2427,N_2137);
xnor U5557 (N_5557,N_2882,N_2273);
xnor U5558 (N_5558,N_3329,N_3737);
nand U5559 (N_5559,N_2622,N_2023);
xnor U5560 (N_5560,N_2441,N_3645);
and U5561 (N_5561,N_2172,N_3308);
or U5562 (N_5562,N_2196,N_2134);
and U5563 (N_5563,N_3886,N_3633);
xor U5564 (N_5564,N_2792,N_2076);
or U5565 (N_5565,N_2651,N_3168);
nand U5566 (N_5566,N_3304,N_2050);
or U5567 (N_5567,N_2932,N_2001);
nand U5568 (N_5568,N_2519,N_2714);
xnor U5569 (N_5569,N_3343,N_2758);
nand U5570 (N_5570,N_3456,N_2227);
nor U5571 (N_5571,N_3270,N_2520);
nor U5572 (N_5572,N_3318,N_3774);
or U5573 (N_5573,N_2471,N_2914);
nor U5574 (N_5574,N_2626,N_2660);
and U5575 (N_5575,N_3211,N_2774);
and U5576 (N_5576,N_2574,N_2063);
nor U5577 (N_5577,N_2691,N_3188);
nor U5578 (N_5578,N_3363,N_2318);
xnor U5579 (N_5579,N_3139,N_3483);
or U5580 (N_5580,N_3087,N_3658);
xor U5581 (N_5581,N_3723,N_2034);
and U5582 (N_5582,N_3247,N_3732);
nor U5583 (N_5583,N_2280,N_2825);
or U5584 (N_5584,N_2011,N_2292);
or U5585 (N_5585,N_3184,N_3567);
nand U5586 (N_5586,N_3291,N_3869);
nor U5587 (N_5587,N_3118,N_3554);
nand U5588 (N_5588,N_3398,N_3372);
nor U5589 (N_5589,N_2520,N_3782);
or U5590 (N_5590,N_3091,N_3014);
and U5591 (N_5591,N_2029,N_2798);
nor U5592 (N_5592,N_2771,N_2837);
or U5593 (N_5593,N_2201,N_2842);
and U5594 (N_5594,N_3930,N_3910);
or U5595 (N_5595,N_2818,N_3618);
and U5596 (N_5596,N_2338,N_3746);
or U5597 (N_5597,N_3011,N_2876);
nand U5598 (N_5598,N_2284,N_2238);
nand U5599 (N_5599,N_3153,N_2256);
nor U5600 (N_5600,N_3720,N_2494);
and U5601 (N_5601,N_3664,N_2983);
nand U5602 (N_5602,N_3801,N_3082);
xnor U5603 (N_5603,N_3048,N_3108);
and U5604 (N_5604,N_2842,N_3522);
nor U5605 (N_5605,N_2861,N_2466);
and U5606 (N_5606,N_3011,N_3028);
nor U5607 (N_5607,N_2662,N_2614);
xnor U5608 (N_5608,N_3331,N_3705);
and U5609 (N_5609,N_2840,N_2022);
or U5610 (N_5610,N_3920,N_3984);
xnor U5611 (N_5611,N_2037,N_2206);
nor U5612 (N_5612,N_3942,N_2063);
and U5613 (N_5613,N_3046,N_3367);
or U5614 (N_5614,N_3707,N_2861);
or U5615 (N_5615,N_3742,N_3452);
or U5616 (N_5616,N_2326,N_2645);
or U5617 (N_5617,N_2363,N_3246);
xor U5618 (N_5618,N_3735,N_2623);
and U5619 (N_5619,N_3308,N_2518);
and U5620 (N_5620,N_3146,N_3259);
or U5621 (N_5621,N_3543,N_3279);
xor U5622 (N_5622,N_2171,N_2116);
or U5623 (N_5623,N_2754,N_2252);
xor U5624 (N_5624,N_2702,N_2500);
xnor U5625 (N_5625,N_2493,N_3893);
nor U5626 (N_5626,N_3387,N_3099);
and U5627 (N_5627,N_3142,N_3813);
nand U5628 (N_5628,N_2526,N_2379);
xor U5629 (N_5629,N_3013,N_2268);
nand U5630 (N_5630,N_2534,N_2772);
nand U5631 (N_5631,N_2292,N_3321);
and U5632 (N_5632,N_2262,N_3721);
or U5633 (N_5633,N_3280,N_2571);
and U5634 (N_5634,N_2463,N_2925);
xnor U5635 (N_5635,N_3682,N_2035);
or U5636 (N_5636,N_2107,N_3846);
or U5637 (N_5637,N_2611,N_3866);
and U5638 (N_5638,N_2485,N_3350);
and U5639 (N_5639,N_3245,N_3919);
and U5640 (N_5640,N_3412,N_3354);
or U5641 (N_5641,N_2081,N_2025);
or U5642 (N_5642,N_3162,N_3248);
or U5643 (N_5643,N_2670,N_2207);
or U5644 (N_5644,N_2967,N_2813);
xor U5645 (N_5645,N_2295,N_3717);
xnor U5646 (N_5646,N_2880,N_2340);
xor U5647 (N_5647,N_3950,N_2250);
and U5648 (N_5648,N_3204,N_2734);
and U5649 (N_5649,N_2666,N_3738);
or U5650 (N_5650,N_3983,N_3320);
or U5651 (N_5651,N_2613,N_2756);
and U5652 (N_5652,N_2259,N_3101);
and U5653 (N_5653,N_2222,N_3418);
nand U5654 (N_5654,N_2042,N_2657);
xor U5655 (N_5655,N_3802,N_2541);
and U5656 (N_5656,N_3987,N_3917);
or U5657 (N_5657,N_3046,N_3837);
and U5658 (N_5658,N_2324,N_3431);
or U5659 (N_5659,N_3516,N_2326);
and U5660 (N_5660,N_2168,N_2292);
nand U5661 (N_5661,N_2241,N_3727);
or U5662 (N_5662,N_2674,N_3035);
and U5663 (N_5663,N_2959,N_3405);
nor U5664 (N_5664,N_2618,N_3822);
and U5665 (N_5665,N_3589,N_2378);
xor U5666 (N_5666,N_2720,N_3309);
nor U5667 (N_5667,N_2590,N_3921);
xor U5668 (N_5668,N_2127,N_2205);
nor U5669 (N_5669,N_3011,N_3668);
or U5670 (N_5670,N_3088,N_3255);
xnor U5671 (N_5671,N_3796,N_3768);
nor U5672 (N_5672,N_2254,N_3875);
or U5673 (N_5673,N_2944,N_2040);
and U5674 (N_5674,N_3704,N_2034);
and U5675 (N_5675,N_3195,N_2630);
or U5676 (N_5676,N_3383,N_2165);
and U5677 (N_5677,N_2373,N_3580);
or U5678 (N_5678,N_2870,N_2332);
and U5679 (N_5679,N_3470,N_2821);
nor U5680 (N_5680,N_3800,N_2131);
xnor U5681 (N_5681,N_3825,N_3502);
nor U5682 (N_5682,N_3064,N_2499);
nor U5683 (N_5683,N_3705,N_3190);
and U5684 (N_5684,N_2946,N_3484);
and U5685 (N_5685,N_3676,N_2106);
or U5686 (N_5686,N_3675,N_2329);
and U5687 (N_5687,N_2965,N_2461);
or U5688 (N_5688,N_2618,N_2587);
nor U5689 (N_5689,N_3502,N_3356);
or U5690 (N_5690,N_2291,N_3838);
or U5691 (N_5691,N_3517,N_3665);
nor U5692 (N_5692,N_2944,N_3574);
xor U5693 (N_5693,N_2184,N_3448);
and U5694 (N_5694,N_3711,N_2767);
or U5695 (N_5695,N_2552,N_3331);
and U5696 (N_5696,N_3824,N_3215);
and U5697 (N_5697,N_3137,N_3383);
xnor U5698 (N_5698,N_3715,N_3697);
nand U5699 (N_5699,N_2881,N_3422);
and U5700 (N_5700,N_2754,N_3342);
and U5701 (N_5701,N_3685,N_2810);
nand U5702 (N_5702,N_3607,N_3182);
and U5703 (N_5703,N_3784,N_2418);
nand U5704 (N_5704,N_3859,N_2870);
nand U5705 (N_5705,N_3637,N_3261);
and U5706 (N_5706,N_2734,N_2648);
xor U5707 (N_5707,N_2141,N_3576);
xnor U5708 (N_5708,N_2570,N_2276);
and U5709 (N_5709,N_2563,N_2446);
or U5710 (N_5710,N_2989,N_2111);
nor U5711 (N_5711,N_2176,N_2597);
nor U5712 (N_5712,N_3411,N_3728);
nand U5713 (N_5713,N_3542,N_2725);
and U5714 (N_5714,N_2221,N_2165);
and U5715 (N_5715,N_2651,N_3977);
nor U5716 (N_5716,N_2780,N_2372);
or U5717 (N_5717,N_2422,N_3738);
nor U5718 (N_5718,N_2060,N_3673);
nor U5719 (N_5719,N_3992,N_3046);
nor U5720 (N_5720,N_3558,N_3461);
nor U5721 (N_5721,N_3754,N_3163);
nand U5722 (N_5722,N_2031,N_2141);
xnor U5723 (N_5723,N_2929,N_2738);
nand U5724 (N_5724,N_3854,N_3832);
nand U5725 (N_5725,N_2390,N_3958);
or U5726 (N_5726,N_3128,N_2135);
and U5727 (N_5727,N_3572,N_2572);
xnor U5728 (N_5728,N_2571,N_2955);
nand U5729 (N_5729,N_3462,N_2671);
nor U5730 (N_5730,N_2932,N_3359);
nand U5731 (N_5731,N_2657,N_3936);
xnor U5732 (N_5732,N_3475,N_3973);
nand U5733 (N_5733,N_3375,N_2098);
xor U5734 (N_5734,N_3656,N_2380);
xnor U5735 (N_5735,N_2692,N_3309);
xor U5736 (N_5736,N_2567,N_3507);
nor U5737 (N_5737,N_3015,N_2482);
nor U5738 (N_5738,N_2345,N_3336);
nand U5739 (N_5739,N_2834,N_3341);
nor U5740 (N_5740,N_3621,N_2018);
or U5741 (N_5741,N_2684,N_2493);
xnor U5742 (N_5742,N_3870,N_2002);
nand U5743 (N_5743,N_3282,N_2610);
nor U5744 (N_5744,N_2904,N_2711);
xor U5745 (N_5745,N_3908,N_3774);
nor U5746 (N_5746,N_2136,N_2376);
or U5747 (N_5747,N_3135,N_2852);
nor U5748 (N_5748,N_2530,N_2409);
nand U5749 (N_5749,N_3682,N_2380);
nor U5750 (N_5750,N_2686,N_2796);
nor U5751 (N_5751,N_2040,N_2128);
xor U5752 (N_5752,N_3969,N_3743);
or U5753 (N_5753,N_3827,N_3960);
xor U5754 (N_5754,N_2347,N_2573);
nor U5755 (N_5755,N_3721,N_2497);
or U5756 (N_5756,N_3936,N_2274);
nor U5757 (N_5757,N_3362,N_2544);
nor U5758 (N_5758,N_3388,N_2804);
or U5759 (N_5759,N_3890,N_3628);
xnor U5760 (N_5760,N_3269,N_3816);
and U5761 (N_5761,N_3830,N_2239);
nor U5762 (N_5762,N_3024,N_3569);
nor U5763 (N_5763,N_2293,N_2084);
and U5764 (N_5764,N_3174,N_2634);
or U5765 (N_5765,N_3055,N_2327);
and U5766 (N_5766,N_2350,N_2071);
xnor U5767 (N_5767,N_3011,N_2244);
nand U5768 (N_5768,N_2940,N_2448);
nor U5769 (N_5769,N_3455,N_3795);
nand U5770 (N_5770,N_2531,N_3459);
nand U5771 (N_5771,N_2527,N_3657);
or U5772 (N_5772,N_2644,N_3444);
nand U5773 (N_5773,N_2701,N_3195);
nor U5774 (N_5774,N_2687,N_3860);
nor U5775 (N_5775,N_2152,N_3656);
nor U5776 (N_5776,N_2819,N_2348);
and U5777 (N_5777,N_3357,N_2787);
nand U5778 (N_5778,N_3801,N_2593);
nor U5779 (N_5779,N_3558,N_3160);
nor U5780 (N_5780,N_2415,N_3710);
xor U5781 (N_5781,N_2202,N_3723);
xnor U5782 (N_5782,N_2607,N_2918);
nand U5783 (N_5783,N_2468,N_2155);
xnor U5784 (N_5784,N_3441,N_3862);
nand U5785 (N_5785,N_3577,N_2788);
and U5786 (N_5786,N_3492,N_3688);
nor U5787 (N_5787,N_3503,N_2940);
or U5788 (N_5788,N_2878,N_3396);
nor U5789 (N_5789,N_2559,N_3063);
and U5790 (N_5790,N_2144,N_2569);
or U5791 (N_5791,N_3502,N_3842);
nand U5792 (N_5792,N_3621,N_2363);
nor U5793 (N_5793,N_3581,N_2865);
or U5794 (N_5794,N_2244,N_3860);
xnor U5795 (N_5795,N_3871,N_2943);
or U5796 (N_5796,N_2293,N_3877);
and U5797 (N_5797,N_3405,N_3198);
and U5798 (N_5798,N_2608,N_3269);
nor U5799 (N_5799,N_2907,N_2621);
nor U5800 (N_5800,N_2288,N_3472);
xnor U5801 (N_5801,N_3597,N_3569);
or U5802 (N_5802,N_3660,N_3662);
xnor U5803 (N_5803,N_2893,N_3434);
and U5804 (N_5804,N_2369,N_3507);
and U5805 (N_5805,N_2126,N_3267);
and U5806 (N_5806,N_2007,N_3206);
or U5807 (N_5807,N_3194,N_2812);
nand U5808 (N_5808,N_2949,N_2173);
or U5809 (N_5809,N_3935,N_2093);
xor U5810 (N_5810,N_3556,N_2149);
nor U5811 (N_5811,N_3349,N_3029);
nand U5812 (N_5812,N_2165,N_3485);
nand U5813 (N_5813,N_3070,N_2338);
xnor U5814 (N_5814,N_2040,N_2262);
and U5815 (N_5815,N_3069,N_3114);
nand U5816 (N_5816,N_2263,N_3674);
nor U5817 (N_5817,N_3894,N_2093);
or U5818 (N_5818,N_2686,N_3468);
nand U5819 (N_5819,N_3265,N_2777);
or U5820 (N_5820,N_2875,N_2418);
and U5821 (N_5821,N_2583,N_2274);
and U5822 (N_5822,N_3442,N_3644);
and U5823 (N_5823,N_2256,N_2224);
nor U5824 (N_5824,N_3252,N_2885);
nand U5825 (N_5825,N_2216,N_3591);
xnor U5826 (N_5826,N_3452,N_2861);
and U5827 (N_5827,N_3956,N_2458);
nor U5828 (N_5828,N_3830,N_2644);
nand U5829 (N_5829,N_3091,N_3505);
xnor U5830 (N_5830,N_2233,N_3670);
and U5831 (N_5831,N_3506,N_2496);
nor U5832 (N_5832,N_3178,N_2779);
or U5833 (N_5833,N_3137,N_3055);
nor U5834 (N_5834,N_3139,N_2968);
nand U5835 (N_5835,N_2381,N_3675);
or U5836 (N_5836,N_3580,N_3283);
nand U5837 (N_5837,N_3297,N_2097);
nand U5838 (N_5838,N_3991,N_3844);
nor U5839 (N_5839,N_3428,N_3062);
and U5840 (N_5840,N_3344,N_2754);
xnor U5841 (N_5841,N_3454,N_3134);
or U5842 (N_5842,N_3367,N_2370);
nand U5843 (N_5843,N_3122,N_2841);
nand U5844 (N_5844,N_3487,N_3583);
nor U5845 (N_5845,N_2327,N_2662);
and U5846 (N_5846,N_3419,N_2935);
xor U5847 (N_5847,N_2304,N_3569);
nor U5848 (N_5848,N_2983,N_3140);
or U5849 (N_5849,N_2966,N_2547);
nor U5850 (N_5850,N_3110,N_2266);
xnor U5851 (N_5851,N_2363,N_3175);
xor U5852 (N_5852,N_2300,N_3291);
nor U5853 (N_5853,N_2924,N_3156);
and U5854 (N_5854,N_2258,N_2523);
nor U5855 (N_5855,N_3769,N_3823);
or U5856 (N_5856,N_3429,N_3058);
nor U5857 (N_5857,N_2706,N_3103);
and U5858 (N_5858,N_2723,N_2858);
nand U5859 (N_5859,N_3496,N_3726);
and U5860 (N_5860,N_3568,N_3018);
nand U5861 (N_5861,N_2238,N_2767);
xnor U5862 (N_5862,N_3794,N_2246);
or U5863 (N_5863,N_2007,N_3717);
or U5864 (N_5864,N_3800,N_2377);
nand U5865 (N_5865,N_3328,N_3764);
nand U5866 (N_5866,N_2335,N_2452);
and U5867 (N_5867,N_2746,N_3611);
xnor U5868 (N_5868,N_2743,N_3994);
nor U5869 (N_5869,N_3370,N_3270);
or U5870 (N_5870,N_3199,N_2143);
xor U5871 (N_5871,N_2612,N_2639);
nand U5872 (N_5872,N_2478,N_3137);
nand U5873 (N_5873,N_2889,N_2645);
nand U5874 (N_5874,N_3073,N_3524);
nand U5875 (N_5875,N_2864,N_2592);
nand U5876 (N_5876,N_3865,N_3185);
or U5877 (N_5877,N_2804,N_3383);
nand U5878 (N_5878,N_3610,N_2652);
nand U5879 (N_5879,N_3109,N_2029);
xnor U5880 (N_5880,N_3811,N_2854);
nor U5881 (N_5881,N_3277,N_3723);
or U5882 (N_5882,N_3004,N_3049);
nor U5883 (N_5883,N_2285,N_3079);
or U5884 (N_5884,N_2088,N_2196);
nand U5885 (N_5885,N_3001,N_3368);
xor U5886 (N_5886,N_3358,N_2399);
nand U5887 (N_5887,N_2218,N_2872);
or U5888 (N_5888,N_2947,N_2645);
or U5889 (N_5889,N_3752,N_3751);
and U5890 (N_5890,N_2224,N_2673);
nor U5891 (N_5891,N_3152,N_2283);
and U5892 (N_5892,N_3708,N_3850);
and U5893 (N_5893,N_3107,N_3040);
and U5894 (N_5894,N_2338,N_3549);
xnor U5895 (N_5895,N_2483,N_2722);
xnor U5896 (N_5896,N_3826,N_2256);
nor U5897 (N_5897,N_3782,N_2379);
nor U5898 (N_5898,N_2214,N_2107);
or U5899 (N_5899,N_3026,N_3716);
nand U5900 (N_5900,N_3396,N_2809);
nor U5901 (N_5901,N_2280,N_2487);
nor U5902 (N_5902,N_2922,N_3039);
xor U5903 (N_5903,N_2318,N_2659);
xnor U5904 (N_5904,N_3364,N_2047);
nor U5905 (N_5905,N_2671,N_2702);
nand U5906 (N_5906,N_2883,N_2924);
and U5907 (N_5907,N_3288,N_3516);
xor U5908 (N_5908,N_2486,N_2370);
or U5909 (N_5909,N_3061,N_3979);
nand U5910 (N_5910,N_2351,N_2260);
nor U5911 (N_5911,N_3799,N_3746);
and U5912 (N_5912,N_2569,N_2859);
nand U5913 (N_5913,N_3395,N_2039);
nor U5914 (N_5914,N_2618,N_2414);
or U5915 (N_5915,N_3975,N_3175);
and U5916 (N_5916,N_2537,N_3653);
nor U5917 (N_5917,N_3678,N_3152);
xor U5918 (N_5918,N_3405,N_3785);
nand U5919 (N_5919,N_3837,N_3489);
xor U5920 (N_5920,N_3389,N_3555);
nand U5921 (N_5921,N_3379,N_3664);
nor U5922 (N_5922,N_3457,N_2977);
nor U5923 (N_5923,N_2325,N_2063);
or U5924 (N_5924,N_2440,N_3007);
nor U5925 (N_5925,N_3914,N_2661);
or U5926 (N_5926,N_3268,N_3923);
nor U5927 (N_5927,N_2595,N_3519);
nor U5928 (N_5928,N_3707,N_3098);
nand U5929 (N_5929,N_3645,N_2852);
and U5930 (N_5930,N_3842,N_3382);
nor U5931 (N_5931,N_2351,N_2084);
xor U5932 (N_5932,N_2540,N_3185);
xor U5933 (N_5933,N_3855,N_2927);
nor U5934 (N_5934,N_2743,N_3282);
and U5935 (N_5935,N_3840,N_3634);
or U5936 (N_5936,N_3458,N_2181);
xnor U5937 (N_5937,N_3453,N_2247);
or U5938 (N_5938,N_2515,N_3749);
xor U5939 (N_5939,N_2836,N_2369);
or U5940 (N_5940,N_3953,N_2262);
and U5941 (N_5941,N_3759,N_2246);
nand U5942 (N_5942,N_2014,N_3740);
or U5943 (N_5943,N_3897,N_3293);
nor U5944 (N_5944,N_2673,N_3791);
nand U5945 (N_5945,N_2081,N_2997);
or U5946 (N_5946,N_3638,N_3331);
and U5947 (N_5947,N_3883,N_3328);
nor U5948 (N_5948,N_3758,N_3497);
nor U5949 (N_5949,N_2445,N_3614);
and U5950 (N_5950,N_2813,N_3595);
nand U5951 (N_5951,N_2485,N_2248);
and U5952 (N_5952,N_3925,N_3805);
nand U5953 (N_5953,N_3500,N_2313);
xnor U5954 (N_5954,N_3582,N_3213);
nand U5955 (N_5955,N_3314,N_2106);
nand U5956 (N_5956,N_3932,N_3346);
nor U5957 (N_5957,N_3633,N_3964);
nor U5958 (N_5958,N_3605,N_2561);
nor U5959 (N_5959,N_3773,N_3939);
nor U5960 (N_5960,N_2905,N_2180);
and U5961 (N_5961,N_3909,N_2080);
nor U5962 (N_5962,N_3409,N_3484);
nor U5963 (N_5963,N_3420,N_2104);
nor U5964 (N_5964,N_2324,N_2969);
or U5965 (N_5965,N_2262,N_3095);
or U5966 (N_5966,N_2752,N_2867);
or U5967 (N_5967,N_3609,N_2921);
nor U5968 (N_5968,N_2247,N_3397);
nor U5969 (N_5969,N_3204,N_2421);
nand U5970 (N_5970,N_3229,N_2778);
and U5971 (N_5971,N_3995,N_3578);
or U5972 (N_5972,N_3070,N_2414);
or U5973 (N_5973,N_3920,N_3865);
nor U5974 (N_5974,N_2150,N_2123);
or U5975 (N_5975,N_2150,N_2439);
xnor U5976 (N_5976,N_2076,N_3283);
or U5977 (N_5977,N_3353,N_3515);
xor U5978 (N_5978,N_2885,N_3682);
xor U5979 (N_5979,N_3703,N_2952);
nor U5980 (N_5980,N_3950,N_2925);
nor U5981 (N_5981,N_2804,N_2171);
and U5982 (N_5982,N_2574,N_2281);
nor U5983 (N_5983,N_2546,N_2593);
nand U5984 (N_5984,N_2277,N_3549);
or U5985 (N_5985,N_2701,N_2435);
nand U5986 (N_5986,N_3390,N_3940);
nand U5987 (N_5987,N_2404,N_2108);
or U5988 (N_5988,N_2019,N_2501);
and U5989 (N_5989,N_2747,N_2562);
and U5990 (N_5990,N_2714,N_2439);
xor U5991 (N_5991,N_3854,N_2724);
xnor U5992 (N_5992,N_2471,N_3267);
and U5993 (N_5993,N_3066,N_3095);
or U5994 (N_5994,N_2557,N_2588);
nor U5995 (N_5995,N_3499,N_2622);
nand U5996 (N_5996,N_3443,N_2440);
nor U5997 (N_5997,N_2206,N_3961);
and U5998 (N_5998,N_2440,N_2754);
nor U5999 (N_5999,N_2120,N_3100);
nor U6000 (N_6000,N_4033,N_4450);
nand U6001 (N_6001,N_4041,N_4480);
xor U6002 (N_6002,N_5322,N_5471);
and U6003 (N_6003,N_5534,N_5447);
xor U6004 (N_6004,N_5090,N_4476);
nand U6005 (N_6005,N_4846,N_4562);
xnor U6006 (N_6006,N_5124,N_4704);
nor U6007 (N_6007,N_5335,N_4975);
nor U6008 (N_6008,N_5824,N_4171);
nand U6009 (N_6009,N_5413,N_5648);
or U6010 (N_6010,N_4003,N_5700);
nand U6011 (N_6011,N_4513,N_4848);
or U6012 (N_6012,N_4248,N_5876);
xor U6013 (N_6013,N_4817,N_4646);
xor U6014 (N_6014,N_4272,N_4954);
nor U6015 (N_6015,N_4967,N_4095);
and U6016 (N_6016,N_5160,N_4469);
nand U6017 (N_6017,N_5491,N_5671);
and U6018 (N_6018,N_5070,N_4166);
xnor U6019 (N_6019,N_4580,N_4705);
nor U6020 (N_6020,N_4579,N_4507);
or U6021 (N_6021,N_4374,N_5523);
or U6022 (N_6022,N_4853,N_4305);
nor U6023 (N_6023,N_4263,N_4155);
or U6024 (N_6024,N_4983,N_4608);
xor U6025 (N_6025,N_5507,N_5302);
or U6026 (N_6026,N_4677,N_4981);
nand U6027 (N_6027,N_4300,N_5309);
or U6028 (N_6028,N_5842,N_5767);
nor U6029 (N_6029,N_4539,N_5715);
nor U6030 (N_6030,N_5906,N_4837);
and U6031 (N_6031,N_4192,N_5011);
nor U6032 (N_6032,N_4721,N_5268);
xnor U6033 (N_6033,N_4093,N_4386);
or U6034 (N_6034,N_5755,N_5622);
xnor U6035 (N_6035,N_4423,N_5705);
nand U6036 (N_6036,N_4605,N_5836);
or U6037 (N_6037,N_5449,N_5199);
or U6038 (N_6038,N_5995,N_5644);
nor U6039 (N_6039,N_5345,N_4655);
xor U6040 (N_6040,N_5247,N_5544);
xnor U6041 (N_6041,N_5063,N_4997);
nand U6042 (N_6042,N_5240,N_4553);
or U6043 (N_6043,N_5058,N_5765);
nor U6044 (N_6044,N_4910,N_4360);
and U6045 (N_6045,N_4213,N_4780);
nand U6046 (N_6046,N_4663,N_4068);
nand U6047 (N_6047,N_4153,N_5900);
or U6048 (N_6048,N_5628,N_5559);
nor U6049 (N_6049,N_5381,N_4748);
or U6050 (N_6050,N_4031,N_5045);
or U6051 (N_6051,N_5225,N_5997);
nor U6052 (N_6052,N_4912,N_5457);
nand U6053 (N_6053,N_5952,N_4464);
xor U6054 (N_6054,N_4109,N_4479);
and U6055 (N_6055,N_5719,N_4428);
nand U6056 (N_6056,N_5157,N_5286);
xor U6057 (N_6057,N_5366,N_4180);
xor U6058 (N_6058,N_5870,N_4494);
xnor U6059 (N_6059,N_5795,N_5281);
or U6060 (N_6060,N_5394,N_5908);
and U6061 (N_6061,N_4368,N_5062);
xnor U6062 (N_6062,N_4738,N_4867);
nor U6063 (N_6063,N_5518,N_4509);
nand U6064 (N_6064,N_4208,N_5179);
nand U6065 (N_6065,N_5789,N_4085);
xnor U6066 (N_6066,N_4865,N_4994);
xor U6067 (N_6067,N_5557,N_5643);
xnor U6068 (N_6068,N_5667,N_5444);
xnor U6069 (N_6069,N_5243,N_4542);
xnor U6070 (N_6070,N_5142,N_5076);
nor U6071 (N_6071,N_4407,N_5012);
and U6072 (N_6072,N_5693,N_5419);
nand U6073 (N_6073,N_5771,N_4687);
nand U6074 (N_6074,N_4991,N_4445);
nor U6075 (N_6075,N_5373,N_4894);
and U6076 (N_6076,N_4736,N_4559);
nand U6077 (N_6077,N_5500,N_5331);
xor U6078 (N_6078,N_5440,N_4990);
nor U6079 (N_6079,N_5015,N_5552);
nand U6080 (N_6080,N_4413,N_4298);
nand U6081 (N_6081,N_5928,N_4652);
nand U6082 (N_6082,N_4661,N_5100);
or U6083 (N_6083,N_5053,N_4276);
or U6084 (N_6084,N_4301,N_4266);
or U6085 (N_6085,N_5535,N_5213);
nand U6086 (N_6086,N_5543,N_4287);
nor U6087 (N_6087,N_5528,N_5135);
nor U6088 (N_6088,N_4676,N_4518);
and U6089 (N_6089,N_4498,N_5730);
or U6090 (N_6090,N_5219,N_4066);
xnor U6091 (N_6091,N_5542,N_4366);
xor U6092 (N_6092,N_4819,N_4601);
xor U6093 (N_6093,N_4822,N_5792);
nor U6094 (N_6094,N_5947,N_5016);
and U6095 (N_6095,N_4129,N_4236);
nand U6096 (N_6096,N_5835,N_4890);
nand U6097 (N_6097,N_5333,N_4173);
xnor U6098 (N_6098,N_5129,N_4055);
nand U6099 (N_6099,N_4941,N_5781);
xor U6100 (N_6100,N_5403,N_4038);
and U6101 (N_6101,N_5714,N_5329);
and U6102 (N_6102,N_4984,N_4120);
and U6103 (N_6103,N_4678,N_5987);
xor U6104 (N_6104,N_5607,N_4483);
nand U6105 (N_6105,N_5769,N_5258);
nand U6106 (N_6106,N_4511,N_5530);
nor U6107 (N_6107,N_5059,N_4945);
and U6108 (N_6108,N_5085,N_4081);
xor U6109 (N_6109,N_5486,N_4787);
or U6110 (N_6110,N_4325,N_5960);
and U6111 (N_6111,N_5862,N_5039);
and U6112 (N_6112,N_4574,N_5222);
or U6113 (N_6113,N_4307,N_5490);
nand U6114 (N_6114,N_5128,N_4987);
nand U6115 (N_6115,N_5158,N_5364);
nor U6116 (N_6116,N_5326,N_4800);
xnor U6117 (N_6117,N_5577,N_5269);
nor U6118 (N_6118,N_4919,N_4348);
or U6119 (N_6119,N_5986,N_5169);
xor U6120 (N_6120,N_5999,N_4082);
or U6121 (N_6121,N_5985,N_5355);
or U6122 (N_6122,N_4660,N_4292);
nor U6123 (N_6123,N_5936,N_4179);
nor U6124 (N_6124,N_4274,N_4878);
and U6125 (N_6125,N_5031,N_4029);
nor U6126 (N_6126,N_4638,N_4004);
nand U6127 (N_6127,N_5476,N_4555);
xnor U6128 (N_6128,N_5297,N_5810);
and U6129 (N_6129,N_4098,N_4543);
or U6130 (N_6130,N_5586,N_5007);
xnor U6131 (N_6131,N_5119,N_5889);
or U6132 (N_6132,N_4146,N_5657);
and U6133 (N_6133,N_5910,N_4679);
nand U6134 (N_6134,N_5925,N_4026);
nor U6135 (N_6135,N_4231,N_4933);
and U6136 (N_6136,N_5159,N_5321);
nor U6137 (N_6137,N_5590,N_5598);
xor U6138 (N_6138,N_4462,N_4640);
nor U6139 (N_6139,N_5474,N_4770);
and U6140 (N_6140,N_4802,N_4895);
nor U6141 (N_6141,N_5887,N_5298);
nor U6142 (N_6142,N_4317,N_4874);
nor U6143 (N_6143,N_5939,N_5639);
or U6144 (N_6144,N_5699,N_4497);
xor U6145 (N_6145,N_5086,N_5097);
or U6146 (N_6146,N_4645,N_5660);
and U6147 (N_6147,N_5234,N_4730);
xor U6148 (N_6148,N_5470,N_5950);
xnor U6149 (N_6149,N_4299,N_4484);
xnor U6150 (N_6150,N_4091,N_4959);
and U6151 (N_6151,N_4045,N_5442);
and U6152 (N_6152,N_4914,N_5075);
nor U6153 (N_6153,N_4972,N_4644);
or U6154 (N_6154,N_5501,N_4383);
or U6155 (N_6155,N_4604,N_5718);
nor U6156 (N_6156,N_5456,N_4233);
and U6157 (N_6157,N_4815,N_4399);
nand U6158 (N_6158,N_4556,N_5791);
and U6159 (N_6159,N_4456,N_5953);
xor U6160 (N_6160,N_5230,N_5347);
or U6161 (N_6161,N_4499,N_5582);
xnor U6162 (N_6162,N_5207,N_4797);
nor U6163 (N_6163,N_4906,N_5111);
nand U6164 (N_6164,N_4779,N_5077);
or U6165 (N_6165,N_4000,N_5130);
xor U6166 (N_6166,N_4757,N_4680);
nand U6167 (N_6167,N_5959,N_5742);
or U6168 (N_6168,N_5416,N_5691);
xnor U6169 (N_6169,N_5662,N_5988);
or U6170 (N_6170,N_5175,N_5775);
nor U6171 (N_6171,N_4771,N_5481);
xor U6172 (N_6172,N_5658,N_4939);
nor U6173 (N_6173,N_4627,N_5010);
nor U6174 (N_6174,N_5702,N_4279);
nor U6175 (N_6175,N_4826,N_4632);
xor U6176 (N_6176,N_5924,N_4013);
or U6177 (N_6177,N_4212,N_4336);
nand U6178 (N_6178,N_5651,N_4930);
nand U6179 (N_6179,N_4648,N_5382);
xnor U6180 (N_6180,N_5632,N_4942);
nand U6181 (N_6181,N_4896,N_4578);
and U6182 (N_6182,N_5185,N_4978);
or U6183 (N_6183,N_5346,N_5935);
or U6184 (N_6184,N_5496,N_5738);
xor U6185 (N_6185,N_5663,N_5672);
xor U6186 (N_6186,N_5592,N_5433);
xnor U6187 (N_6187,N_4491,N_4143);
xnor U6188 (N_6188,N_4056,N_5441);
or U6189 (N_6189,N_5990,N_4949);
nor U6190 (N_6190,N_5880,N_4079);
and U6191 (N_6191,N_4753,N_5450);
nand U6192 (N_6192,N_4027,N_4183);
xnor U6193 (N_6193,N_5074,N_4566);
xnor U6194 (N_6194,N_4203,N_4228);
and U6195 (N_6195,N_4882,N_5479);
or U6196 (N_6196,N_5246,N_5517);
xor U6197 (N_6197,N_4102,N_4893);
nand U6198 (N_6198,N_5525,N_5674);
nor U6199 (N_6199,N_5037,N_4436);
and U6200 (N_6200,N_5375,N_4432);
nor U6201 (N_6201,N_4868,N_5429);
or U6202 (N_6202,N_4801,N_5018);
xor U6203 (N_6203,N_5430,N_4391);
nor U6204 (N_6204,N_5740,N_4007);
and U6205 (N_6205,N_4724,N_5872);
nand U6206 (N_6206,N_5844,N_4793);
nor U6207 (N_6207,N_4825,N_5485);
nand U6208 (N_6208,N_4546,N_5165);
and U6209 (N_6209,N_5197,N_5885);
or U6210 (N_6210,N_5890,N_5806);
and U6211 (N_6211,N_4623,N_5669);
or U6212 (N_6212,N_4370,N_4584);
and U6213 (N_6213,N_5732,N_5608);
nand U6214 (N_6214,N_4227,N_5772);
or U6215 (N_6215,N_5593,N_4599);
nand U6216 (N_6216,N_5808,N_5955);
nand U6217 (N_6217,N_4214,N_5370);
or U6218 (N_6218,N_4139,N_4977);
xnor U6219 (N_6219,N_5673,N_4851);
xnor U6220 (N_6220,N_5365,N_5584);
or U6221 (N_6221,N_5646,N_5984);
and U6222 (N_6222,N_4998,N_5073);
xnor U6223 (N_6223,N_5841,N_4995);
and U6224 (N_6224,N_5815,N_4658);
xnor U6225 (N_6225,N_4037,N_4406);
or U6226 (N_6226,N_4395,N_4060);
nand U6227 (N_6227,N_5531,N_4582);
or U6228 (N_6228,N_4267,N_5654);
xnor U6229 (N_6229,N_5864,N_5274);
or U6230 (N_6230,N_5541,N_5549);
and U6231 (N_6231,N_4812,N_4160);
or U6232 (N_6232,N_5484,N_4200);
xor U6233 (N_6233,N_4295,N_5304);
or U6234 (N_6234,N_5971,N_5261);
nand U6235 (N_6235,N_4782,N_5023);
nand U6236 (N_6236,N_5736,N_5478);
and U6237 (N_6237,N_4694,N_5563);
xor U6238 (N_6238,N_5524,N_4576);
or U6239 (N_6239,N_4936,N_5827);
and U6240 (N_6240,N_4962,N_5882);
and U6241 (N_6241,N_5993,N_4794);
nor U6242 (N_6242,N_5706,N_4829);
nand U6243 (N_6243,N_4653,N_4788);
or U6244 (N_6244,N_5907,N_5389);
nor U6245 (N_6245,N_5548,N_5316);
nor U6246 (N_6246,N_4455,N_4193);
xnor U6247 (N_6247,N_5652,N_5323);
or U6248 (N_6248,N_5601,N_4282);
xnor U6249 (N_6249,N_4525,N_4903);
xnor U6250 (N_6250,N_5623,N_4493);
nand U6251 (N_6251,N_4538,N_5339);
xnor U6252 (N_6252,N_5152,N_5773);
xor U6253 (N_6253,N_4289,N_5121);
nor U6254 (N_6254,N_4918,N_4877);
nand U6255 (N_6255,N_4734,N_5728);
or U6256 (N_6256,N_5104,N_5251);
nor U6257 (N_6257,N_5828,N_4232);
nand U6258 (N_6258,N_5380,N_5432);
or U6259 (N_6259,N_4859,N_5205);
nor U6260 (N_6260,N_5102,N_4008);
or U6261 (N_6261,N_5685,N_5176);
xor U6262 (N_6262,N_4732,N_5707);
or U6263 (N_6263,N_4698,N_4696);
nor U6264 (N_6264,N_4205,N_4626);
and U6265 (N_6265,N_4937,N_4879);
nor U6266 (N_6266,N_4306,N_5363);
xor U6267 (N_6267,N_4440,N_5797);
xnor U6268 (N_6268,N_5303,N_5932);
and U6269 (N_6269,N_5362,N_5218);
or U6270 (N_6270,N_4354,N_4598);
and U6271 (N_6271,N_5492,N_5711);
xnor U6272 (N_6272,N_5992,N_4375);
nor U6273 (N_6273,N_4904,N_5962);
xor U6274 (N_6274,N_4841,N_5570);
nand U6275 (N_6275,N_4531,N_4224);
xnor U6276 (N_6276,N_4950,N_5353);
nor U6277 (N_6277,N_4387,N_4527);
and U6278 (N_6278,N_5743,N_4594);
xor U6279 (N_6279,N_4537,N_4720);
nor U6280 (N_6280,N_4683,N_4958);
xor U6281 (N_6281,N_5150,N_4052);
xnor U6282 (N_6282,N_5242,N_4080);
or U6283 (N_6283,N_4589,N_4570);
xor U6284 (N_6284,N_5081,N_5799);
xnor U6285 (N_6285,N_5256,N_5678);
nor U6286 (N_6286,N_4659,N_4427);
nor U6287 (N_6287,N_5972,N_4350);
or U6288 (N_6288,N_4402,N_4377);
or U6289 (N_6289,N_5386,N_4367);
nand U6290 (N_6290,N_4144,N_4749);
nand U6291 (N_6291,N_5757,N_5241);
nand U6292 (N_6292,N_4051,N_5968);
or U6293 (N_6293,N_5676,N_4265);
or U6294 (N_6294,N_5725,N_5493);
and U6295 (N_6295,N_5227,N_4397);
or U6296 (N_6296,N_5894,N_5406);
xor U6297 (N_6297,N_4642,N_4197);
nor U6298 (N_6298,N_5560,N_5417);
or U6299 (N_6299,N_5438,N_5591);
or U6300 (N_6300,N_5259,N_4790);
or U6301 (N_6301,N_5066,N_5282);
xnor U6302 (N_6302,N_5589,N_4773);
nor U6303 (N_6303,N_5927,N_4884);
xor U6304 (N_6304,N_4152,N_4839);
or U6305 (N_6305,N_5578,N_5445);
xor U6306 (N_6306,N_5047,N_5522);
or U6307 (N_6307,N_5279,N_5290);
xnor U6308 (N_6308,N_4145,N_4250);
nand U6309 (N_6309,N_5454,N_4709);
and U6310 (N_6310,N_4832,N_4636);
or U6311 (N_6311,N_5125,N_4795);
xor U6312 (N_6312,N_5930,N_5777);
or U6313 (N_6313,N_5830,N_4989);
and U6314 (N_6314,N_5285,N_5392);
and U6315 (N_6315,N_5554,N_4765);
nor U6316 (N_6316,N_4575,N_5099);
nand U6317 (N_6317,N_4611,N_4988);
and U6318 (N_6318,N_4421,N_4714);
xnor U6319 (N_6319,N_5049,N_4411);
xnor U6320 (N_6320,N_4500,N_5991);
nor U6321 (N_6321,N_4073,N_4828);
nor U6322 (N_6322,N_5127,N_5854);
nand U6323 (N_6323,N_4666,N_4836);
nand U6324 (N_6324,N_5284,N_5720);
xor U6325 (N_6325,N_5878,N_5946);
xor U6326 (N_6326,N_4178,N_4293);
nor U6327 (N_6327,N_5000,N_4590);
nor U6328 (N_6328,N_5195,N_5891);
nand U6329 (N_6329,N_5605,N_4747);
and U6330 (N_6330,N_5372,N_4597);
xor U6331 (N_6331,N_5349,N_5087);
and U6332 (N_6332,N_4215,N_4861);
nand U6333 (N_6333,N_4487,N_4092);
and U6334 (N_6334,N_5458,N_4563);
xnor U6335 (N_6335,N_4799,N_5480);
nand U6336 (N_6336,N_4613,N_5027);
nand U6337 (N_6337,N_5411,N_4070);
nor U6338 (N_6338,N_4742,N_4380);
nand U6339 (N_6339,N_4186,N_4113);
xnor U6340 (N_6340,N_5790,N_5182);
nand U6341 (N_6341,N_5847,N_4225);
and U6342 (N_6342,N_4347,N_5938);
and U6343 (N_6343,N_5469,N_5237);
and U6344 (N_6344,N_5171,N_4125);
nand U6345 (N_6345,N_5788,N_4264);
xnor U6346 (N_6346,N_4755,N_5311);
nand U6347 (N_6347,N_5055,N_4296);
nand U6348 (N_6348,N_4544,N_4430);
nor U6349 (N_6349,N_4345,N_4137);
xor U6350 (N_6350,N_5191,N_5005);
nand U6351 (N_6351,N_5398,N_4302);
nor U6352 (N_6352,N_5856,N_5040);
and U6353 (N_6353,N_5922,N_4554);
nor U6354 (N_6354,N_5221,N_5970);
and U6355 (N_6355,N_5278,N_4743);
and U6356 (N_6356,N_4530,N_5001);
nor U6357 (N_6357,N_4651,N_4385);
and U6358 (N_6358,N_4047,N_5538);
xnor U6359 (N_6359,N_5168,N_5198);
and U6360 (N_6360,N_5606,N_4686);
and U6361 (N_6361,N_4774,N_4415);
xnor U6362 (N_6362,N_4681,N_5424);
and U6363 (N_6363,N_4217,N_5903);
xor U6364 (N_6364,N_4618,N_4591);
or U6365 (N_6365,N_4364,N_5271);
and U6366 (N_6366,N_4438,N_4833);
nor U6367 (N_6367,N_5201,N_4435);
nand U6368 (N_6368,N_5209,N_5495);
nor U6369 (N_6369,N_5164,N_4123);
and U6370 (N_6370,N_5314,N_4211);
xnor U6371 (N_6371,N_5499,N_5342);
or U6372 (N_6372,N_5146,N_4885);
nand U6373 (N_6373,N_4495,N_4581);
nand U6374 (N_6374,N_4077,N_4585);
or U6375 (N_6375,N_5181,N_4813);
and U6376 (N_6376,N_4784,N_4925);
or U6377 (N_6377,N_4634,N_5024);
and U6378 (N_6378,N_5327,N_4280);
or U6379 (N_6379,N_5112,N_4177);
and U6380 (N_6380,N_5871,N_4718);
nand U6381 (N_6381,N_5819,N_4012);
or U6382 (N_6382,N_5186,N_5371);
nor U6383 (N_6383,N_4496,N_4439);
and U6384 (N_6384,N_4195,N_4631);
or U6385 (N_6385,N_4806,N_4856);
and U6386 (N_6386,N_4058,N_5902);
and U6387 (N_6387,N_4913,N_5096);
nor U6388 (N_6388,N_5266,N_5734);
or U6389 (N_6389,N_4021,N_4053);
xor U6390 (N_6390,N_4275,N_4326);
or U6391 (N_6391,N_5294,N_4259);
and U6392 (N_6392,N_5579,N_4147);
or U6393 (N_6393,N_4323,N_4946);
xor U6394 (N_6394,N_5735,N_4961);
or U6395 (N_6395,N_5954,N_5211);
xnor U6396 (N_6396,N_4722,N_4405);
nand U6397 (N_6397,N_5410,N_5916);
xor U6398 (N_6398,N_4548,N_4169);
nor U6399 (N_6399,N_5395,N_4222);
nor U6400 (N_6400,N_5162,N_5798);
and U6401 (N_6401,N_5154,N_5802);
nand U6402 (N_6402,N_4750,N_5338);
nand U6403 (N_6403,N_5180,N_4786);
xor U6404 (N_6404,N_4332,N_5110);
xnor U6405 (N_6405,N_5974,N_5132);
nor U6406 (N_6406,N_5336,N_5141);
xnor U6407 (N_6407,N_5255,N_4478);
nor U6408 (N_6408,N_5566,N_4669);
xor U6409 (N_6409,N_5459,N_5768);
nor U6410 (N_6410,N_5793,N_5238);
nand U6411 (N_6411,N_4022,N_5034);
or U6412 (N_6412,N_4811,N_5519);
nand U6413 (N_6413,N_5510,N_5758);
or U6414 (N_6414,N_5123,N_5703);
nor U6415 (N_6415,N_4752,N_5875);
nand U6416 (N_6416,N_4595,N_5625);
or U6417 (N_6417,N_4711,N_4116);
or U6418 (N_6418,N_4286,N_4313);
nor U6419 (N_6419,N_5546,N_4444);
xor U6420 (N_6420,N_5686,N_5937);
nand U6421 (N_6421,N_4094,N_5727);
nor U6422 (N_6422,N_4522,N_5325);
nor U6423 (N_6423,N_5785,N_5020);
xor U6424 (N_6424,N_5067,N_5273);
and U6425 (N_6425,N_4372,N_4869);
or U6426 (N_6426,N_5229,N_4219);
nand U6427 (N_6427,N_4561,N_4664);
and U6428 (N_6428,N_4624,N_4573);
and U6429 (N_6429,N_4400,N_4515);
or U6430 (N_6430,N_4713,N_4100);
nor U6431 (N_6431,N_4514,N_4396);
and U6432 (N_6432,N_4019,N_5611);
nor U6433 (N_6433,N_5717,N_4737);
nor U6434 (N_6434,N_4754,N_4957);
nor U6435 (N_6435,N_4571,N_5301);
nand U6436 (N_6436,N_4426,N_5989);
xnor U6437 (N_6437,N_4524,N_5957);
xnor U6438 (N_6438,N_5803,N_5330);
nor U6439 (N_6439,N_5145,N_5929);
xor U6440 (N_6440,N_4229,N_5640);
xor U6441 (N_6441,N_4294,N_5551);
xor U6442 (N_6442,N_4410,N_4682);
xor U6443 (N_6443,N_4695,N_5427);
nand U6444 (N_6444,N_4670,N_4703);
nand U6445 (N_6445,N_5529,N_5387);
and U6446 (N_6446,N_4588,N_4729);
nor U6447 (N_6447,N_5504,N_5724);
nor U6448 (N_6448,N_5264,N_4206);
xnor U6449 (N_6449,N_4965,N_4097);
and U6450 (N_6450,N_4168,N_4980);
or U6451 (N_6451,N_5307,N_4603);
nor U6452 (N_6452,N_5713,N_4124);
nand U6453 (N_6453,N_5204,N_5783);
or U6454 (N_6454,N_5813,N_4459);
nand U6455 (N_6455,N_5254,N_4121);
or U6456 (N_6456,N_4532,N_4897);
or U6457 (N_6457,N_5943,N_4049);
xnor U6458 (N_6458,N_5376,N_4460);
or U6459 (N_6459,N_4069,N_5352);
nand U6460 (N_6460,N_5217,N_4550);
and U6461 (N_6461,N_5461,N_4629);
xor U6462 (N_6462,N_4412,N_5809);
nor U6463 (N_6463,N_4150,N_4772);
and U6464 (N_6464,N_4087,N_4569);
xor U6465 (N_6465,N_4111,N_5451);
xor U6466 (N_6466,N_4216,N_4334);
and U6467 (N_6467,N_5821,N_5681);
nand U6468 (N_6468,N_4766,N_4020);
xor U6469 (N_6469,N_4928,N_5439);
xor U6470 (N_6470,N_5776,N_5917);
xnor U6471 (N_6471,N_4242,N_5635);
or U6472 (N_6472,N_5656,N_4017);
nor U6473 (N_6473,N_5919,N_4916);
and U6474 (N_6474,N_4132,N_4615);
nor U6475 (N_6475,N_5751,N_5036);
or U6476 (N_6476,N_4014,N_4130);
xor U6477 (N_6477,N_5909,N_4767);
nand U6478 (N_6478,N_5423,N_4172);
nand U6479 (N_6479,N_5228,N_4324);
or U6480 (N_6480,N_5443,N_5782);
nand U6481 (N_6481,N_4157,N_4067);
xnor U6482 (N_6482,N_4947,N_5041);
nand U6483 (N_6483,N_5649,N_4838);
or U6484 (N_6484,N_4974,N_5624);
nand U6485 (N_6485,N_5196,N_4844);
nor U6486 (N_6486,N_4744,N_5536);
or U6487 (N_6487,N_5556,N_5565);
or U6488 (N_6488,N_5134,N_5633);
or U6489 (N_6489,N_5980,N_4520);
xor U6490 (N_6490,N_5745,N_5756);
or U6491 (N_6491,N_5636,N_5019);
nor U6492 (N_6492,N_5462,N_5621);
nand U6493 (N_6493,N_5638,N_5631);
nor U6494 (N_6494,N_4419,N_5194);
and U6495 (N_6495,N_4526,N_4740);
nor U6496 (N_6496,N_5283,N_4798);
or U6497 (N_6497,N_5540,N_5561);
or U6498 (N_6498,N_5028,N_4873);
nor U6499 (N_6499,N_4420,N_4447);
nor U6500 (N_6500,N_5641,N_4078);
and U6501 (N_6501,N_5661,N_4246);
nand U6502 (N_6502,N_5343,N_4359);
or U6503 (N_6503,N_4731,N_5167);
and U6504 (N_6504,N_4448,N_5422);
xor U6505 (N_6505,N_5739,N_5299);
xor U6506 (N_6506,N_4074,N_5401);
xnor U6507 (N_6507,N_5516,N_5083);
xnor U6508 (N_6508,N_5982,N_5328);
and U6509 (N_6509,N_5899,N_5337);
or U6510 (N_6510,N_4508,N_4471);
nand U6511 (N_6511,N_5095,N_5383);
nand U6512 (N_6512,N_4159,N_4751);
xor U6513 (N_6513,N_5192,N_4715);
and U6514 (N_6514,N_5208,N_5829);
nor U6515 (N_6515,N_5276,N_4039);
nand U6516 (N_6516,N_5428,N_5231);
nor U6517 (N_6517,N_5961,N_5613);
nand U6518 (N_6518,N_5103,N_4088);
nor U6519 (N_6519,N_5721,N_4938);
xor U6520 (N_6520,N_5203,N_5668);
nand U6521 (N_6521,N_4356,N_4639);
or U6522 (N_6522,N_4362,N_5701);
or U6523 (N_6523,N_4401,N_4908);
nand U6524 (N_6524,N_4956,N_4131);
and U6525 (N_6525,N_4127,N_5388);
or U6526 (N_6526,N_5588,N_5761);
nor U6527 (N_6527,N_4218,N_4437);
and U6528 (N_6528,N_5468,N_4256);
xnor U6529 (N_6529,N_4671,N_5915);
xnor U6530 (N_6530,N_4643,N_4327);
xnor U6531 (N_6531,N_5232,N_5147);
or U6532 (N_6532,N_4789,N_4245);
xor U6533 (N_6533,N_4905,N_4807);
and U6534 (N_6534,N_5022,N_5473);
nand U6535 (N_6535,N_4700,N_4441);
or U6536 (N_6536,N_5568,N_5619);
nor U6537 (N_6537,N_4072,N_5369);
and U6538 (N_6538,N_4727,N_4257);
nand U6539 (N_6539,N_5184,N_4917);
nand U6540 (N_6540,N_5116,N_4188);
or U6541 (N_6541,N_4547,N_4084);
nand U6542 (N_6542,N_4628,N_4076);
or U6543 (N_6543,N_4392,N_4971);
nand U6544 (N_6544,N_5637,N_5949);
nand U6545 (N_6545,N_4993,N_5295);
or U6546 (N_6546,N_5448,N_4973);
xor U6547 (N_6547,N_4115,N_4185);
nand U6548 (N_6548,N_4607,N_5697);
or U6549 (N_6549,N_5655,N_5825);
or U6550 (N_6550,N_4909,N_5926);
nand U6551 (N_6551,N_4376,N_5453);
xor U6552 (N_6552,N_5766,N_4048);
or U6553 (N_6553,N_4529,N_4226);
nor U6554 (N_6554,N_4136,N_5396);
or U6555 (N_6555,N_5215,N_5503);
or U6556 (N_6556,N_5630,N_5080);
and U6557 (N_6557,N_5004,N_4783);
nand U6558 (N_6558,N_5341,N_5571);
nand U6559 (N_6559,N_4625,N_5558);
nand U6560 (N_6560,N_5308,N_5187);
xor U6561 (N_6561,N_5839,N_5101);
nor U6562 (N_6562,N_4816,N_5144);
xnor U6563 (N_6563,N_5811,N_5051);
and U6564 (N_6564,N_5845,N_4835);
nand U6565 (N_6565,N_5688,N_5868);
nor U6566 (N_6566,N_5866,N_5078);
xnor U6567 (N_6567,N_4810,N_4650);
or U6568 (N_6568,N_4863,N_4018);
nand U6569 (N_6569,N_4057,N_4273);
xor U6570 (N_6570,N_4308,N_4234);
nor U6571 (N_6571,N_5515,N_5071);
nor U6572 (N_6572,N_5360,N_4330);
xor U6573 (N_6573,N_4823,N_4924);
nand U6574 (N_6574,N_5188,N_4099);
xnor U6575 (N_6575,N_4475,N_5117);
nor U6576 (N_6576,N_4845,N_5137);
nand U6577 (N_6577,N_5178,N_5537);
nand U6578 (N_6578,N_5778,N_4176);
or U6579 (N_6579,N_5057,N_4649);
xor U6580 (N_6580,N_4443,N_5467);
and U6581 (N_6581,N_4831,N_4010);
or U6582 (N_6582,N_5061,N_4764);
and U6583 (N_6583,N_4071,N_5506);
or U6584 (N_6584,N_5709,N_4353);
nor U6585 (N_6585,N_5514,N_4119);
and U6586 (N_6586,N_5645,N_5780);
or U6587 (N_6587,N_4244,N_4596);
xnor U6588 (N_6588,N_4059,N_4446);
or U6589 (N_6589,N_4042,N_5942);
and U6590 (N_6590,N_5072,N_5452);
xnor U6591 (N_6591,N_4281,N_4251);
nand U6592 (N_6592,N_5006,N_5886);
nor U6593 (N_6593,N_4175,N_4321);
and U6594 (N_6594,N_5400,N_5804);
or U6595 (N_6595,N_5604,N_4149);
and U6596 (N_6596,N_4196,N_4254);
nand U6597 (N_6597,N_5555,N_5287);
nand U6598 (N_6598,N_5620,N_5173);
xor U6599 (N_6599,N_4620,N_4763);
nand U6600 (N_6600,N_4898,N_4290);
nand U6601 (N_6601,N_4221,N_4723);
or U6602 (N_6602,N_4291,N_5694);
xnor U6603 (N_6603,N_5665,N_4174);
and U6604 (N_6604,N_4210,N_4468);
nand U6605 (N_6605,N_4866,N_4717);
nor U6606 (N_6606,N_5404,N_4966);
or U6607 (N_6607,N_4504,N_4050);
nor U6608 (N_6608,N_4202,N_4593);
nor U6609 (N_6609,N_5418,N_5934);
or U6610 (N_6610,N_5161,N_4619);
xnor U6611 (N_6611,N_5105,N_4331);
or U6612 (N_6612,N_5402,N_5350);
xnor U6613 (N_6613,N_5690,N_4382);
or U6614 (N_6614,N_5089,N_4269);
and U6615 (N_6615,N_5288,N_4818);
nor U6616 (N_6616,N_4424,N_5733);
xor U6617 (N_6617,N_4927,N_4025);
or U6618 (N_6618,N_4830,N_4960);
nand U6619 (N_6619,N_5650,N_5267);
nand U6620 (N_6620,N_5750,N_4034);
nor U6621 (N_6621,N_5659,N_5708);
nand U6622 (N_6622,N_5405,N_4996);
xnor U6623 (N_6623,N_4485,N_4114);
xnor U6624 (N_6624,N_4388,N_5465);
or U6625 (N_6625,N_4320,N_5497);
xnor U6626 (N_6626,N_4768,N_4122);
and U6627 (N_6627,N_5737,N_4931);
and U6628 (N_6628,N_5113,N_4249);
or U6629 (N_6629,N_5190,N_4090);
nand U6630 (N_6630,N_5567,N_5223);
and U6631 (N_6631,N_5716,N_5280);
or U6632 (N_6632,N_5312,N_5877);
xnor U6633 (N_6633,N_4466,N_5779);
nor U6634 (N_6634,N_4899,N_4541);
or U6635 (N_6635,N_4064,N_4028);
nor U6636 (N_6636,N_4148,N_4834);
nand U6637 (N_6637,N_5634,N_4338);
xor U6638 (N_6638,N_5069,N_5834);
xor U6639 (N_6639,N_5046,N_5319);
xnor U6640 (N_6640,N_5580,N_4690);
nand U6641 (N_6641,N_5026,N_4577);
and U6642 (N_6642,N_4481,N_5963);
or U6643 (N_6643,N_5747,N_4032);
and U6644 (N_6644,N_5973,N_4379);
nor U6645 (N_6645,N_4156,N_4344);
and U6646 (N_6646,N_5435,N_5446);
nor U6647 (N_6647,N_5177,N_5911);
xnor U6648 (N_6648,N_5807,N_5114);
and U6649 (N_6649,N_4463,N_5357);
xor U6650 (N_6650,N_4921,N_5865);
xor U6651 (N_6651,N_4283,N_5088);
xnor U6652 (N_6652,N_4449,N_4907);
nor U6653 (N_6653,N_4612,N_4852);
xnor U6654 (N_6654,N_5800,N_4434);
nand U6655 (N_6655,N_4668,N_4948);
nand U6656 (N_6656,N_4394,N_5214);
xnor U6657 (N_6657,N_4621,N_4785);
nand U6658 (N_6658,N_5933,N_5511);
nand U6659 (N_6659,N_4699,N_4689);
or U6660 (N_6660,N_4923,N_4587);
nand U6661 (N_6661,N_4549,N_4384);
xor U6662 (N_6662,N_4270,N_5260);
xor U6663 (N_6663,N_5367,N_4535);
and U6664 (N_6664,N_5901,N_4418);
and U6665 (N_6665,N_4103,N_4241);
nand U6666 (N_6666,N_5091,N_4209);
nor U6667 (N_6667,N_5126,N_5408);
or U6668 (N_6668,N_4633,N_4952);
and U6669 (N_6669,N_4862,N_4647);
or U6670 (N_6670,N_5155,N_5320);
xor U6671 (N_6671,N_4181,N_5754);
nand U6672 (N_6672,N_4610,N_5550);
xor U6673 (N_6673,N_4506,N_4329);
xnor U6674 (N_6674,N_4922,N_5434);
nand U6675 (N_6675,N_4381,N_4635);
or U6676 (N_6676,N_5385,N_5994);
xor U6677 (N_6677,N_4842,N_5617);
xnor U6678 (N_6678,N_5921,N_5873);
xor U6679 (N_6679,N_5817,N_5596);
nand U6680 (N_6680,N_4328,N_4458);
or U6681 (N_6681,N_5814,N_4207);
nand U6682 (N_6682,N_5996,N_4190);
xor U6683 (N_6683,N_5014,N_5391);
or U6684 (N_6684,N_4716,N_5863);
nor U6685 (N_6685,N_5426,N_4309);
nand U6686 (N_6686,N_4880,N_4756);
or U6687 (N_6687,N_5883,N_5210);
nand U6688 (N_6688,N_5292,N_4086);
nand U6689 (N_6689,N_5245,N_5595);
nand U6690 (N_6690,N_4775,N_4312);
nand U6691 (N_6691,N_4517,N_4617);
xor U6692 (N_6692,N_5043,N_4701);
nor U6693 (N_6693,N_4404,N_5532);
nor U6694 (N_6694,N_4986,N_4791);
or U6695 (N_6695,N_5272,N_4821);
nor U6696 (N_6696,N_5216,N_4706);
nand U6697 (N_6697,N_4255,N_5874);
or U6698 (N_6698,N_5220,N_5860);
or U6699 (N_6699,N_4151,N_4762);
or U6700 (N_6700,N_4142,N_5030);
nand U6701 (N_6701,N_5764,N_4429);
nor U6702 (N_6702,N_4141,N_5581);
or U6703 (N_6703,N_4335,N_4201);
and U6704 (N_6704,N_5969,N_4505);
and U6705 (N_6705,N_4015,N_5770);
nand U6706 (N_6706,N_5393,N_4776);
nor U6707 (N_6707,N_5892,N_4803);
nand U6708 (N_6708,N_5614,N_5494);
nand U6709 (N_6709,N_5033,N_5574);
and U6710 (N_6710,N_4488,N_4089);
or U6711 (N_6711,N_4252,N_5318);
nor U6712 (N_6712,N_4106,N_5675);
and U6713 (N_6713,N_4708,N_5784);
nor U6714 (N_6714,N_4920,N_5884);
nor U6715 (N_6715,N_4107,N_5533);
nand U6716 (N_6716,N_5120,N_4849);
xor U6717 (N_6717,N_4871,N_5421);
or U6718 (N_6718,N_5746,N_4016);
and U6719 (N_6719,N_4726,N_5502);
or U6720 (N_6720,N_5965,N_5626);
and U6721 (N_6721,N_5079,N_5850);
nand U6722 (N_6722,N_5140,N_4393);
or U6723 (N_6723,N_5615,N_4002);
nor U6724 (N_6724,N_5384,N_5460);
or U6725 (N_6725,N_5677,N_4858);
xnor U6726 (N_6726,N_5893,N_4943);
and U6727 (N_6727,N_5275,N_4482);
nor U6728 (N_6728,N_5851,N_5958);
and U6729 (N_6729,N_4191,N_5966);
nand U6730 (N_6730,N_4339,N_5390);
xnor U6731 (N_6731,N_5553,N_4284);
nor U6732 (N_6732,N_5763,N_5670);
and U6733 (N_6733,N_4416,N_5898);
nand U6734 (N_6734,N_4881,N_4902);
and U6735 (N_6735,N_4741,N_4240);
and U6736 (N_6736,N_4969,N_5163);
nor U6737 (N_6737,N_5931,N_4614);
nor U6738 (N_6738,N_5978,N_4940);
nor U6739 (N_6739,N_4352,N_5857);
xor U6740 (N_6740,N_5324,N_5148);
xor U6741 (N_6741,N_4691,N_4528);
and U6742 (N_6742,N_4194,N_4536);
and U6743 (N_6743,N_4061,N_5224);
xnor U6744 (N_6744,N_5545,N_5594);
nor U6745 (N_6745,N_5849,N_5576);
or U6746 (N_6746,N_5206,N_5358);
or U6747 (N_6747,N_4083,N_4616);
and U6748 (N_6748,N_5689,N_5975);
nor U6749 (N_6749,N_5683,N_4230);
nand U6750 (N_6750,N_5712,N_4477);
or U6751 (N_6751,N_4888,N_4953);
xnor U6752 (N_6752,N_5483,N_4271);
and U6753 (N_6753,N_4892,N_4390);
xnor U6754 (N_6754,N_4808,N_5153);
nor U6755 (N_6755,N_5977,N_4985);
or U6756 (N_6756,N_5084,N_4285);
or U6757 (N_6757,N_4365,N_4237);
or U6758 (N_6758,N_5945,N_5044);
nand U6759 (N_6759,N_5923,N_5008);
nor U6760 (N_6760,N_5744,N_5796);
nor U6761 (N_6761,N_5840,N_4043);
xnor U6762 (N_6762,N_5368,N_5054);
nand U6763 (N_6763,N_5981,N_4134);
nand U6764 (N_6764,N_4243,N_5603);
and U6765 (N_6765,N_4850,N_4030);
nand U6766 (N_6766,N_5263,N_4260);
nand U6767 (N_6767,N_4900,N_4009);
xor U6768 (N_6768,N_4674,N_5399);
and U6769 (N_6769,N_5489,N_5038);
or U6770 (N_6770,N_5156,N_4105);
xor U6771 (N_6771,N_5826,N_5569);
nand U6772 (N_6772,N_4847,N_4667);
or U6773 (N_6773,N_5172,N_4685);
or U6774 (N_6774,N_5032,N_5998);
nor U6775 (N_6775,N_5642,N_4707);
nor U6776 (N_6776,N_4804,N_4746);
and U6777 (N_6777,N_5139,N_4165);
nand U6778 (N_6778,N_5521,N_5235);
nor U6779 (N_6779,N_4697,N_4138);
and U6780 (N_6780,N_5853,N_5823);
and U6781 (N_6781,N_5455,N_5913);
nand U6782 (N_6782,N_5378,N_4371);
or U6783 (N_6783,N_5509,N_4944);
or U6784 (N_6784,N_4710,N_5305);
nor U6785 (N_6785,N_4461,N_5526);
and U6786 (N_6786,N_4693,N_5547);
nand U6787 (N_6787,N_4929,N_5976);
nand U6788 (N_6788,N_4164,N_5679);
nor U6789 (N_6789,N_5695,N_5202);
or U6790 (N_6790,N_4557,N_4820);
nor U6791 (N_6791,N_4792,N_4519);
xor U6792 (N_6792,N_5226,N_5236);
xor U6793 (N_6793,N_5682,N_4023);
nor U6794 (N_6794,N_5048,N_5354);
xnor U6795 (N_6795,N_5482,N_5361);
nor U6796 (N_6796,N_4545,N_4451);
nand U6797 (N_6797,N_4035,N_5956);
nor U6798 (N_6798,N_5239,N_4901);
nor U6799 (N_6799,N_4654,N_5520);
and U6800 (N_6800,N_4341,N_4108);
nand U6801 (N_6801,N_4662,N_4337);
and U6802 (N_6802,N_5106,N_4322);
xor U6803 (N_6803,N_4110,N_4005);
and U6804 (N_6804,N_4602,N_5816);
nand U6805 (N_6805,N_4870,N_5729);
or U6806 (N_6806,N_5002,N_4872);
and U6807 (N_6807,N_5664,N_5600);
xnor U6808 (N_6808,N_5914,N_4692);
and U6809 (N_6809,N_4075,N_5262);
nand U6810 (N_6810,N_4135,N_5377);
or U6811 (N_6811,N_4040,N_4968);
xor U6812 (N_6812,N_4316,N_5300);
nand U6813 (N_6813,N_4465,N_5951);
and U6814 (N_6814,N_4970,N_5359);
or U6815 (N_6815,N_5332,N_5912);
xor U6816 (N_6816,N_5291,N_5436);
or U6817 (N_6817,N_4128,N_4198);
xor U6818 (N_6818,N_5837,N_5244);
and U6819 (N_6819,N_4133,N_4304);
or U6820 (N_6820,N_4592,N_4247);
and U6821 (N_6821,N_5174,N_5115);
or U6822 (N_6822,N_5334,N_4104);
xnor U6823 (N_6823,N_4860,N_5881);
nor U6824 (N_6824,N_5498,N_4006);
nand U6825 (N_6825,N_4062,N_4657);
nand U6826 (N_6826,N_4735,N_5692);
xor U6827 (N_6827,N_4063,N_4358);
and U6828 (N_6828,N_4778,N_5944);
or U6829 (N_6829,N_4684,N_4964);
or U6830 (N_6830,N_4158,N_5068);
nor U6831 (N_6831,N_4702,N_4346);
nand U6832 (N_6832,N_5021,N_4760);
nor U6833 (N_6833,N_4915,N_4431);
and U6834 (N_6834,N_5602,N_4665);
nand U6835 (N_6835,N_4503,N_5093);
and U6836 (N_6836,N_5351,N_5488);
nand U6837 (N_6837,N_5415,N_4389);
nand U6838 (N_6838,N_5964,N_5249);
nor U6839 (N_6839,N_4982,N_5948);
xnor U6840 (N_6840,N_5722,N_4167);
nand U6841 (N_6841,N_5846,N_5609);
xnor U6842 (N_6842,N_5979,N_5472);
xnor U6843 (N_6843,N_4712,N_5253);
xnor U6844 (N_6844,N_5832,N_5527);
and U6845 (N_6845,N_4510,N_5879);
or U6846 (N_6846,N_5653,N_5296);
nand U6847 (N_6847,N_4759,N_4622);
nor U6848 (N_6848,N_4725,N_4963);
and U6849 (N_6849,N_5753,N_4126);
or U6850 (N_6850,N_5464,N_5306);
or U6851 (N_6851,N_5583,N_5833);
xor U6852 (N_6852,N_4992,N_5094);
or U6853 (N_6853,N_5466,N_5616);
nor U6854 (N_6854,N_5562,N_5508);
and U6855 (N_6855,N_5741,N_5629);
and U6856 (N_6856,N_4363,N_4452);
nor U6857 (N_6857,N_4277,N_5374);
and U6858 (N_6858,N_4238,N_4001);
nor U6859 (N_6859,N_5166,N_5151);
and U6860 (N_6860,N_5170,N_4777);
or U6861 (N_6861,N_4673,N_5861);
nor U6862 (N_6862,N_4926,N_5897);
nand U6863 (N_6863,N_5731,N_4220);
or U6864 (N_6864,N_5774,N_5138);
xor U6865 (N_6865,N_4999,N_4184);
xor U6866 (N_6866,N_5136,N_4540);
nand U6867 (N_6867,N_4855,N_4606);
and U6868 (N_6868,N_4911,N_4470);
or U6869 (N_6869,N_4398,N_5118);
and U6870 (N_6870,N_4521,N_5612);
nor U6871 (N_6871,N_5888,N_4036);
nand U6872 (N_6872,N_5293,N_4170);
xnor U6873 (N_6873,N_5257,N_4745);
nor U6874 (N_6874,N_4096,N_4189);
xor U6875 (N_6875,N_4814,N_4163);
or U6876 (N_6876,N_4501,N_5122);
xor U6877 (N_6877,N_4567,N_5505);
or U6878 (N_6878,N_5983,N_4425);
or U6879 (N_6879,N_4467,N_5277);
nor U6880 (N_6880,N_4568,N_4672);
and U6881 (N_6881,N_5941,N_4739);
nor U6882 (N_6882,N_5064,N_5822);
and U6883 (N_6883,N_4408,N_5794);
and U6884 (N_6884,N_5869,N_4630);
and U6885 (N_6885,N_4349,N_5017);
or U6886 (N_6886,N_4357,N_4840);
nor U6887 (N_6887,N_4351,N_4512);
nand U6888 (N_6888,N_4875,N_5183);
nand U6889 (N_6889,N_4932,N_5065);
xor U6890 (N_6890,N_4565,N_5787);
nor U6891 (N_6891,N_5585,N_4935);
xnor U6892 (N_6892,N_5564,N_4378);
and U6893 (N_6893,N_5696,N_4889);
nor U6894 (N_6894,N_4805,N_4857);
and U6895 (N_6895,N_5317,N_5042);
xor U6896 (N_6896,N_4600,N_4442);
nand U6897 (N_6897,N_5109,N_4311);
xor U6898 (N_6898,N_4319,N_4891);
and U6899 (N_6899,N_4572,N_5749);
xor U6900 (N_6900,N_4761,N_4262);
nor U6901 (N_6901,N_5092,N_5698);
nor U6902 (N_6902,N_4887,N_4489);
nand U6903 (N_6903,N_5726,N_5610);
xnor U6904 (N_6904,N_4046,N_5487);
or U6905 (N_6905,N_4318,N_4827);
and U6906 (N_6906,N_4199,N_4502);
or U6907 (N_6907,N_5060,N_5704);
xor U6908 (N_6908,N_4204,N_5618);
and U6909 (N_6909,N_4472,N_4490);
xor U6910 (N_6910,N_5248,N_4979);
or U6911 (N_6911,N_5573,N_5820);
xor U6912 (N_6912,N_4552,N_5539);
or U6913 (N_6913,N_4182,N_5867);
and U6914 (N_6914,N_4886,N_4883);
and U6915 (N_6915,N_5250,N_4934);
and U6916 (N_6916,N_4054,N_4656);
or U6917 (N_6917,N_4310,N_4101);
nand U6918 (N_6918,N_5760,N_4976);
xnor U6919 (N_6919,N_5340,N_4641);
xor U6920 (N_6920,N_5855,N_4355);
nor U6921 (N_6921,N_4409,N_5477);
and U6922 (N_6922,N_5805,N_4523);
xnor U6923 (N_6923,N_5940,N_5818);
nand U6924 (N_6924,N_4474,N_5407);
xor U6925 (N_6925,N_5356,N_4951);
nand U6926 (N_6926,N_4258,N_5918);
and U6927 (N_6927,N_5050,N_4024);
nand U6928 (N_6928,N_4809,N_4583);
nand U6929 (N_6929,N_5003,N_4162);
or U6930 (N_6930,N_4854,N_5896);
xor U6931 (N_6931,N_4268,N_4422);
nand U6932 (N_6932,N_4609,N_5098);
xor U6933 (N_6933,N_5149,N_5838);
nor U6934 (N_6934,N_5599,N_4457);
xnor U6935 (N_6935,N_4315,N_5475);
nor U6936 (N_6936,N_4876,N_5848);
xnor U6937 (N_6937,N_4781,N_5904);
or U6938 (N_6938,N_4564,N_5786);
and U6939 (N_6939,N_5315,N_5133);
xnor U6940 (N_6940,N_5052,N_4314);
and U6941 (N_6941,N_4369,N_5463);
or U6942 (N_6942,N_5313,N_4955);
nor U6943 (N_6943,N_4864,N_5752);
and U6944 (N_6944,N_5812,N_5409);
nand U6945 (N_6945,N_4235,N_5420);
and U6946 (N_6946,N_5762,N_5597);
nand U6947 (N_6947,N_4486,N_4403);
nor U6948 (N_6948,N_5265,N_5759);
or U6949 (N_6949,N_4533,N_5512);
nand U6950 (N_6950,N_5344,N_4288);
nand U6951 (N_6951,N_4333,N_5025);
nor U6952 (N_6952,N_5013,N_4140);
and U6953 (N_6953,N_4340,N_5270);
or U6954 (N_6954,N_5905,N_5108);
xnor U6955 (N_6955,N_4733,N_4011);
nand U6956 (N_6956,N_5437,N_5425);
or U6957 (N_6957,N_5852,N_4044);
or U6958 (N_6958,N_5189,N_5379);
nor U6959 (N_6959,N_4342,N_4253);
nand U6960 (N_6960,N_5575,N_5587);
xor U6961 (N_6961,N_4453,N_4843);
and U6962 (N_6962,N_5895,N_5687);
or U6963 (N_6963,N_5831,N_5200);
or U6964 (N_6964,N_5858,N_5082);
and U6965 (N_6965,N_4586,N_5131);
nor U6966 (N_6966,N_4769,N_4261);
and U6967 (N_6967,N_4187,N_5666);
and U6968 (N_6968,N_5252,N_4796);
nand U6969 (N_6969,N_5193,N_5572);
xnor U6970 (N_6970,N_4758,N_5029);
and U6971 (N_6971,N_5680,N_4492);
nand U6972 (N_6972,N_5967,N_5412);
xor U6973 (N_6973,N_5431,N_4297);
nor U6974 (N_6974,N_4637,N_5289);
and U6975 (N_6975,N_4675,N_5035);
or U6976 (N_6976,N_4161,N_5143);
nand U6977 (N_6977,N_5843,N_4373);
and U6978 (N_6978,N_4728,N_4558);
or U6979 (N_6979,N_5310,N_5723);
and U6980 (N_6980,N_4118,N_5627);
nor U6981 (N_6981,N_4688,N_4239);
nor U6982 (N_6982,N_4414,N_5212);
nor U6983 (N_6983,N_4065,N_5801);
and U6984 (N_6984,N_5414,N_4223);
nor U6985 (N_6985,N_5748,N_5056);
xnor U6986 (N_6986,N_4551,N_4473);
and U6987 (N_6987,N_5859,N_5233);
nor U6988 (N_6988,N_4117,N_5009);
and U6989 (N_6989,N_5647,N_5348);
or U6990 (N_6990,N_4278,N_4343);
or U6991 (N_6991,N_4454,N_4154);
and U6992 (N_6992,N_4433,N_4112);
and U6993 (N_6993,N_4361,N_4516);
or U6994 (N_6994,N_5684,N_5397);
and U6995 (N_6995,N_5513,N_5920);
or U6996 (N_6996,N_4719,N_4534);
or U6997 (N_6997,N_4417,N_5107);
and U6998 (N_6998,N_4303,N_4824);
nand U6999 (N_6999,N_5710,N_4560);
or U7000 (N_7000,N_5607,N_4892);
xnor U7001 (N_7001,N_5814,N_5242);
and U7002 (N_7002,N_4632,N_5723);
nor U7003 (N_7003,N_5827,N_4158);
nor U7004 (N_7004,N_4187,N_4913);
xnor U7005 (N_7005,N_4725,N_5364);
and U7006 (N_7006,N_5735,N_5608);
nor U7007 (N_7007,N_5443,N_5676);
nor U7008 (N_7008,N_5505,N_4019);
nor U7009 (N_7009,N_5215,N_4498);
xor U7010 (N_7010,N_4922,N_5728);
nand U7011 (N_7011,N_4057,N_5244);
or U7012 (N_7012,N_4657,N_4839);
nor U7013 (N_7013,N_4921,N_5687);
xor U7014 (N_7014,N_4569,N_5634);
nand U7015 (N_7015,N_4975,N_5739);
nor U7016 (N_7016,N_5294,N_4489);
nor U7017 (N_7017,N_4420,N_4243);
nor U7018 (N_7018,N_5539,N_4386);
nor U7019 (N_7019,N_4415,N_4981);
nand U7020 (N_7020,N_5856,N_5263);
nand U7021 (N_7021,N_4667,N_4823);
and U7022 (N_7022,N_5005,N_4054);
nor U7023 (N_7023,N_5483,N_4415);
xor U7024 (N_7024,N_4904,N_4093);
nand U7025 (N_7025,N_4213,N_4767);
and U7026 (N_7026,N_5967,N_4293);
and U7027 (N_7027,N_5113,N_4245);
xnor U7028 (N_7028,N_4354,N_4957);
xnor U7029 (N_7029,N_5034,N_5021);
nand U7030 (N_7030,N_5599,N_4192);
xnor U7031 (N_7031,N_4084,N_4807);
and U7032 (N_7032,N_5372,N_5066);
xor U7033 (N_7033,N_4107,N_4985);
and U7034 (N_7034,N_4827,N_4459);
nand U7035 (N_7035,N_5520,N_4068);
or U7036 (N_7036,N_5650,N_5302);
and U7037 (N_7037,N_5814,N_4057);
nor U7038 (N_7038,N_5912,N_5955);
and U7039 (N_7039,N_4617,N_5795);
nor U7040 (N_7040,N_5740,N_4462);
and U7041 (N_7041,N_4641,N_5143);
and U7042 (N_7042,N_4934,N_4346);
nor U7043 (N_7043,N_5842,N_5378);
xor U7044 (N_7044,N_4980,N_5311);
nor U7045 (N_7045,N_5391,N_5670);
nor U7046 (N_7046,N_5560,N_5694);
xor U7047 (N_7047,N_5831,N_5438);
xnor U7048 (N_7048,N_5176,N_4617);
or U7049 (N_7049,N_5022,N_4895);
nand U7050 (N_7050,N_5259,N_4466);
xor U7051 (N_7051,N_4115,N_5234);
or U7052 (N_7052,N_4846,N_5116);
xnor U7053 (N_7053,N_5560,N_5763);
xnor U7054 (N_7054,N_5013,N_5207);
and U7055 (N_7055,N_4713,N_4186);
xnor U7056 (N_7056,N_4209,N_5913);
and U7057 (N_7057,N_4190,N_4606);
nand U7058 (N_7058,N_5909,N_4332);
nand U7059 (N_7059,N_5590,N_5804);
nand U7060 (N_7060,N_5315,N_4867);
xnor U7061 (N_7061,N_5916,N_4834);
and U7062 (N_7062,N_5578,N_5200);
and U7063 (N_7063,N_4587,N_4418);
and U7064 (N_7064,N_5241,N_5857);
and U7065 (N_7065,N_4977,N_5494);
nor U7066 (N_7066,N_5743,N_4432);
or U7067 (N_7067,N_4366,N_5633);
and U7068 (N_7068,N_4626,N_5959);
nand U7069 (N_7069,N_4924,N_4673);
nor U7070 (N_7070,N_4711,N_5873);
or U7071 (N_7071,N_4772,N_4018);
xor U7072 (N_7072,N_4930,N_5370);
nand U7073 (N_7073,N_4008,N_5078);
nor U7074 (N_7074,N_5174,N_4734);
or U7075 (N_7075,N_4171,N_5343);
xnor U7076 (N_7076,N_5227,N_5023);
xor U7077 (N_7077,N_4698,N_4415);
xor U7078 (N_7078,N_4456,N_4502);
or U7079 (N_7079,N_5985,N_5069);
xnor U7080 (N_7080,N_5903,N_5172);
or U7081 (N_7081,N_5089,N_5000);
and U7082 (N_7082,N_4508,N_4932);
nor U7083 (N_7083,N_4212,N_5779);
xor U7084 (N_7084,N_4921,N_5512);
nand U7085 (N_7085,N_5953,N_5896);
nor U7086 (N_7086,N_4215,N_5512);
nand U7087 (N_7087,N_4291,N_4136);
and U7088 (N_7088,N_5961,N_5527);
or U7089 (N_7089,N_4543,N_5578);
nor U7090 (N_7090,N_5148,N_4318);
and U7091 (N_7091,N_5400,N_4252);
nand U7092 (N_7092,N_5236,N_5000);
and U7093 (N_7093,N_4358,N_5398);
and U7094 (N_7094,N_5463,N_4491);
xor U7095 (N_7095,N_4378,N_5236);
nand U7096 (N_7096,N_4548,N_5954);
nand U7097 (N_7097,N_5378,N_4501);
nand U7098 (N_7098,N_5098,N_4407);
and U7099 (N_7099,N_5750,N_4669);
nor U7100 (N_7100,N_4842,N_4281);
and U7101 (N_7101,N_5893,N_4290);
xnor U7102 (N_7102,N_5952,N_5210);
nand U7103 (N_7103,N_5748,N_5903);
nor U7104 (N_7104,N_5833,N_4262);
or U7105 (N_7105,N_5852,N_4769);
xnor U7106 (N_7106,N_4006,N_4534);
xnor U7107 (N_7107,N_5272,N_5684);
or U7108 (N_7108,N_5321,N_4937);
or U7109 (N_7109,N_5395,N_5141);
and U7110 (N_7110,N_5700,N_5926);
nand U7111 (N_7111,N_4323,N_4413);
and U7112 (N_7112,N_4893,N_4711);
nand U7113 (N_7113,N_5144,N_5305);
xor U7114 (N_7114,N_4509,N_5036);
and U7115 (N_7115,N_5329,N_5205);
or U7116 (N_7116,N_5871,N_5765);
or U7117 (N_7117,N_5944,N_4422);
nor U7118 (N_7118,N_4991,N_5731);
and U7119 (N_7119,N_4686,N_5774);
xnor U7120 (N_7120,N_4658,N_5402);
nor U7121 (N_7121,N_4838,N_5714);
and U7122 (N_7122,N_4391,N_4195);
xnor U7123 (N_7123,N_4570,N_4115);
nor U7124 (N_7124,N_5939,N_5074);
and U7125 (N_7125,N_5560,N_5839);
and U7126 (N_7126,N_5109,N_5344);
or U7127 (N_7127,N_5741,N_4324);
nand U7128 (N_7128,N_5743,N_4303);
xnor U7129 (N_7129,N_5333,N_4715);
xor U7130 (N_7130,N_5316,N_4677);
nor U7131 (N_7131,N_4185,N_5658);
nand U7132 (N_7132,N_5575,N_4918);
or U7133 (N_7133,N_4568,N_5723);
xnor U7134 (N_7134,N_4222,N_4426);
or U7135 (N_7135,N_4299,N_4050);
or U7136 (N_7136,N_5503,N_5733);
nor U7137 (N_7137,N_5405,N_5721);
nand U7138 (N_7138,N_4938,N_5378);
nor U7139 (N_7139,N_4854,N_4304);
xnor U7140 (N_7140,N_4099,N_4175);
nor U7141 (N_7141,N_5003,N_5449);
xor U7142 (N_7142,N_5631,N_5284);
xor U7143 (N_7143,N_4966,N_5695);
nand U7144 (N_7144,N_5108,N_5199);
nand U7145 (N_7145,N_5110,N_4571);
xor U7146 (N_7146,N_5121,N_5565);
or U7147 (N_7147,N_4955,N_5671);
nand U7148 (N_7148,N_4729,N_5610);
nor U7149 (N_7149,N_5738,N_4157);
xor U7150 (N_7150,N_4513,N_4389);
or U7151 (N_7151,N_5079,N_4324);
nor U7152 (N_7152,N_5157,N_5129);
or U7153 (N_7153,N_5768,N_4578);
or U7154 (N_7154,N_5148,N_5097);
or U7155 (N_7155,N_4098,N_4038);
and U7156 (N_7156,N_4048,N_4291);
nor U7157 (N_7157,N_4080,N_5418);
xor U7158 (N_7158,N_4634,N_5389);
nand U7159 (N_7159,N_5743,N_5102);
or U7160 (N_7160,N_4530,N_5410);
or U7161 (N_7161,N_5728,N_5892);
nor U7162 (N_7162,N_4295,N_5328);
nor U7163 (N_7163,N_5682,N_5155);
and U7164 (N_7164,N_4179,N_4438);
nand U7165 (N_7165,N_5894,N_5694);
or U7166 (N_7166,N_4393,N_5745);
nand U7167 (N_7167,N_4651,N_5063);
or U7168 (N_7168,N_4741,N_4658);
or U7169 (N_7169,N_4561,N_5686);
or U7170 (N_7170,N_4056,N_4689);
nor U7171 (N_7171,N_5811,N_5805);
and U7172 (N_7172,N_4600,N_5487);
nand U7173 (N_7173,N_5503,N_4128);
nor U7174 (N_7174,N_5058,N_5052);
or U7175 (N_7175,N_5820,N_5214);
and U7176 (N_7176,N_4241,N_5873);
nor U7177 (N_7177,N_5892,N_5859);
xor U7178 (N_7178,N_4322,N_5042);
xor U7179 (N_7179,N_5416,N_5934);
xnor U7180 (N_7180,N_5865,N_5475);
xor U7181 (N_7181,N_4306,N_5655);
xnor U7182 (N_7182,N_4383,N_4626);
or U7183 (N_7183,N_5170,N_5376);
nand U7184 (N_7184,N_4320,N_4236);
nand U7185 (N_7185,N_4876,N_4717);
xor U7186 (N_7186,N_4131,N_5258);
nand U7187 (N_7187,N_4523,N_5758);
nand U7188 (N_7188,N_5028,N_5642);
or U7189 (N_7189,N_5571,N_4043);
or U7190 (N_7190,N_4616,N_4953);
nor U7191 (N_7191,N_5744,N_5309);
xnor U7192 (N_7192,N_4972,N_4463);
xnor U7193 (N_7193,N_4547,N_5747);
and U7194 (N_7194,N_5291,N_5882);
xor U7195 (N_7195,N_5775,N_4840);
or U7196 (N_7196,N_4734,N_4005);
nand U7197 (N_7197,N_4495,N_5417);
nor U7198 (N_7198,N_5806,N_5042);
nor U7199 (N_7199,N_5775,N_5540);
xnor U7200 (N_7200,N_4163,N_5651);
nor U7201 (N_7201,N_5352,N_5416);
xor U7202 (N_7202,N_5718,N_5485);
or U7203 (N_7203,N_5063,N_4554);
or U7204 (N_7204,N_4481,N_4063);
nor U7205 (N_7205,N_4187,N_5679);
nand U7206 (N_7206,N_4152,N_4954);
xor U7207 (N_7207,N_4701,N_5662);
nor U7208 (N_7208,N_5470,N_4825);
and U7209 (N_7209,N_4033,N_5552);
nor U7210 (N_7210,N_4053,N_5494);
or U7211 (N_7211,N_5071,N_5079);
and U7212 (N_7212,N_4734,N_5613);
or U7213 (N_7213,N_4019,N_5945);
and U7214 (N_7214,N_4718,N_5214);
nand U7215 (N_7215,N_5605,N_4542);
nor U7216 (N_7216,N_4923,N_5394);
or U7217 (N_7217,N_4832,N_5917);
and U7218 (N_7218,N_5969,N_4166);
and U7219 (N_7219,N_4758,N_4224);
nand U7220 (N_7220,N_5724,N_4314);
nor U7221 (N_7221,N_5509,N_5958);
nor U7222 (N_7222,N_5263,N_4267);
nor U7223 (N_7223,N_5810,N_5135);
or U7224 (N_7224,N_4007,N_5881);
xnor U7225 (N_7225,N_4587,N_5598);
nand U7226 (N_7226,N_4062,N_5581);
xnor U7227 (N_7227,N_4397,N_4028);
nand U7228 (N_7228,N_4071,N_5694);
nand U7229 (N_7229,N_5085,N_4552);
xor U7230 (N_7230,N_4651,N_5801);
nor U7231 (N_7231,N_5026,N_5786);
and U7232 (N_7232,N_5004,N_5931);
or U7233 (N_7233,N_5994,N_4378);
nand U7234 (N_7234,N_5252,N_4170);
nor U7235 (N_7235,N_5755,N_5880);
xnor U7236 (N_7236,N_5530,N_4110);
or U7237 (N_7237,N_4647,N_4468);
xnor U7238 (N_7238,N_4870,N_5095);
nor U7239 (N_7239,N_4722,N_5403);
and U7240 (N_7240,N_4254,N_4651);
or U7241 (N_7241,N_4974,N_4041);
and U7242 (N_7242,N_5501,N_4637);
nor U7243 (N_7243,N_5139,N_5234);
nor U7244 (N_7244,N_4828,N_5349);
nor U7245 (N_7245,N_4155,N_5682);
nand U7246 (N_7246,N_4103,N_4923);
xor U7247 (N_7247,N_4058,N_5207);
nand U7248 (N_7248,N_4172,N_4058);
or U7249 (N_7249,N_4902,N_4452);
nor U7250 (N_7250,N_4000,N_5464);
nor U7251 (N_7251,N_4316,N_4754);
nor U7252 (N_7252,N_4674,N_5198);
and U7253 (N_7253,N_5456,N_5455);
nor U7254 (N_7254,N_5875,N_5365);
xnor U7255 (N_7255,N_5977,N_5101);
xnor U7256 (N_7256,N_5646,N_5395);
and U7257 (N_7257,N_4157,N_5526);
or U7258 (N_7258,N_4332,N_5090);
and U7259 (N_7259,N_5910,N_5750);
nor U7260 (N_7260,N_4036,N_5405);
and U7261 (N_7261,N_5119,N_5169);
nand U7262 (N_7262,N_4028,N_4002);
or U7263 (N_7263,N_4817,N_5427);
xor U7264 (N_7264,N_4029,N_5766);
and U7265 (N_7265,N_4854,N_4712);
xnor U7266 (N_7266,N_5836,N_5551);
nand U7267 (N_7267,N_4788,N_5368);
and U7268 (N_7268,N_5682,N_5902);
nor U7269 (N_7269,N_4732,N_5316);
nor U7270 (N_7270,N_5017,N_4718);
or U7271 (N_7271,N_5256,N_4775);
and U7272 (N_7272,N_4137,N_5300);
or U7273 (N_7273,N_5962,N_4102);
nand U7274 (N_7274,N_4279,N_5934);
nand U7275 (N_7275,N_4304,N_5508);
xor U7276 (N_7276,N_4850,N_5220);
or U7277 (N_7277,N_5735,N_5977);
nand U7278 (N_7278,N_4021,N_4426);
and U7279 (N_7279,N_4234,N_5640);
nand U7280 (N_7280,N_4487,N_5113);
nor U7281 (N_7281,N_4685,N_5874);
nor U7282 (N_7282,N_5163,N_5053);
and U7283 (N_7283,N_5196,N_5720);
and U7284 (N_7284,N_4863,N_4464);
nor U7285 (N_7285,N_5402,N_4790);
nor U7286 (N_7286,N_5006,N_5433);
xor U7287 (N_7287,N_5275,N_5424);
or U7288 (N_7288,N_5330,N_4120);
nand U7289 (N_7289,N_4942,N_4411);
xnor U7290 (N_7290,N_5725,N_5464);
nor U7291 (N_7291,N_5261,N_5631);
or U7292 (N_7292,N_5839,N_4387);
nand U7293 (N_7293,N_4714,N_4180);
or U7294 (N_7294,N_4223,N_5651);
nor U7295 (N_7295,N_4208,N_5575);
nor U7296 (N_7296,N_4266,N_4276);
xnor U7297 (N_7297,N_4487,N_4228);
or U7298 (N_7298,N_4260,N_4811);
or U7299 (N_7299,N_4845,N_5531);
and U7300 (N_7300,N_5667,N_5727);
xor U7301 (N_7301,N_5300,N_4163);
nor U7302 (N_7302,N_4118,N_5695);
or U7303 (N_7303,N_5095,N_5663);
nor U7304 (N_7304,N_5761,N_5561);
and U7305 (N_7305,N_5038,N_4305);
nand U7306 (N_7306,N_5146,N_4909);
nor U7307 (N_7307,N_4282,N_5172);
xnor U7308 (N_7308,N_4488,N_5577);
nor U7309 (N_7309,N_4279,N_4203);
nand U7310 (N_7310,N_4517,N_5899);
or U7311 (N_7311,N_5768,N_4345);
or U7312 (N_7312,N_4890,N_5115);
nor U7313 (N_7313,N_4348,N_5766);
xor U7314 (N_7314,N_4010,N_4833);
and U7315 (N_7315,N_5970,N_4993);
xnor U7316 (N_7316,N_5872,N_5307);
and U7317 (N_7317,N_4323,N_4117);
or U7318 (N_7318,N_5562,N_5771);
nand U7319 (N_7319,N_4322,N_4784);
nor U7320 (N_7320,N_5618,N_4769);
nand U7321 (N_7321,N_5298,N_4708);
nor U7322 (N_7322,N_5796,N_4088);
xor U7323 (N_7323,N_4349,N_5322);
or U7324 (N_7324,N_4207,N_4279);
nor U7325 (N_7325,N_4624,N_5441);
nand U7326 (N_7326,N_4538,N_5649);
xor U7327 (N_7327,N_4574,N_4107);
and U7328 (N_7328,N_4115,N_4425);
xnor U7329 (N_7329,N_4879,N_5390);
or U7330 (N_7330,N_4558,N_5668);
and U7331 (N_7331,N_4865,N_5564);
and U7332 (N_7332,N_5266,N_4715);
xor U7333 (N_7333,N_4701,N_5485);
xor U7334 (N_7334,N_5811,N_5907);
nand U7335 (N_7335,N_4863,N_4274);
nand U7336 (N_7336,N_4282,N_4170);
nand U7337 (N_7337,N_4930,N_4558);
and U7338 (N_7338,N_5911,N_5949);
nor U7339 (N_7339,N_4260,N_4902);
or U7340 (N_7340,N_4277,N_4815);
or U7341 (N_7341,N_4727,N_4075);
and U7342 (N_7342,N_4041,N_4527);
nor U7343 (N_7343,N_5338,N_4691);
nand U7344 (N_7344,N_4588,N_5261);
and U7345 (N_7345,N_5510,N_4509);
nor U7346 (N_7346,N_5918,N_4340);
xor U7347 (N_7347,N_5303,N_4797);
nand U7348 (N_7348,N_4070,N_5749);
xnor U7349 (N_7349,N_5915,N_5761);
nand U7350 (N_7350,N_5501,N_5942);
and U7351 (N_7351,N_5467,N_5965);
or U7352 (N_7352,N_4702,N_5113);
or U7353 (N_7353,N_4132,N_5942);
nand U7354 (N_7354,N_5063,N_4710);
and U7355 (N_7355,N_5288,N_5824);
nand U7356 (N_7356,N_5392,N_5577);
xor U7357 (N_7357,N_5185,N_5680);
and U7358 (N_7358,N_4933,N_5402);
nor U7359 (N_7359,N_4932,N_4762);
and U7360 (N_7360,N_5781,N_5131);
xnor U7361 (N_7361,N_5577,N_4357);
or U7362 (N_7362,N_4657,N_4545);
nor U7363 (N_7363,N_5972,N_5502);
or U7364 (N_7364,N_4603,N_4005);
xnor U7365 (N_7365,N_5642,N_5063);
xor U7366 (N_7366,N_4140,N_5864);
or U7367 (N_7367,N_5525,N_5815);
nor U7368 (N_7368,N_4080,N_4640);
nor U7369 (N_7369,N_4654,N_5341);
nor U7370 (N_7370,N_4032,N_5935);
nor U7371 (N_7371,N_5011,N_4032);
nand U7372 (N_7372,N_5263,N_5851);
and U7373 (N_7373,N_4438,N_4625);
or U7374 (N_7374,N_5634,N_5222);
xor U7375 (N_7375,N_4628,N_5704);
xor U7376 (N_7376,N_4336,N_5258);
nand U7377 (N_7377,N_4799,N_5320);
or U7378 (N_7378,N_4561,N_4267);
xnor U7379 (N_7379,N_5828,N_4558);
and U7380 (N_7380,N_4093,N_4209);
or U7381 (N_7381,N_4353,N_4709);
nand U7382 (N_7382,N_4568,N_4342);
nor U7383 (N_7383,N_5384,N_5663);
xnor U7384 (N_7384,N_4771,N_5132);
xnor U7385 (N_7385,N_5320,N_5247);
nand U7386 (N_7386,N_5574,N_5560);
nand U7387 (N_7387,N_4056,N_4944);
or U7388 (N_7388,N_5482,N_5736);
or U7389 (N_7389,N_4420,N_4204);
or U7390 (N_7390,N_5267,N_4358);
nor U7391 (N_7391,N_5883,N_5603);
and U7392 (N_7392,N_4499,N_5389);
or U7393 (N_7393,N_4570,N_5892);
nor U7394 (N_7394,N_5872,N_4054);
and U7395 (N_7395,N_4831,N_5244);
nand U7396 (N_7396,N_4826,N_4257);
and U7397 (N_7397,N_5045,N_5184);
and U7398 (N_7398,N_4086,N_4546);
or U7399 (N_7399,N_5037,N_4463);
and U7400 (N_7400,N_4812,N_4351);
or U7401 (N_7401,N_4586,N_5127);
and U7402 (N_7402,N_5162,N_4916);
or U7403 (N_7403,N_5685,N_5142);
or U7404 (N_7404,N_4964,N_4341);
or U7405 (N_7405,N_5453,N_5496);
or U7406 (N_7406,N_5424,N_5470);
and U7407 (N_7407,N_5280,N_5695);
nor U7408 (N_7408,N_5966,N_5793);
or U7409 (N_7409,N_4207,N_5142);
nor U7410 (N_7410,N_5784,N_4040);
or U7411 (N_7411,N_5965,N_5497);
xnor U7412 (N_7412,N_4093,N_5643);
nand U7413 (N_7413,N_4814,N_4890);
xor U7414 (N_7414,N_5250,N_4269);
and U7415 (N_7415,N_4407,N_4958);
nor U7416 (N_7416,N_5278,N_5437);
xnor U7417 (N_7417,N_4291,N_4514);
xnor U7418 (N_7418,N_4653,N_4313);
xor U7419 (N_7419,N_5695,N_5455);
or U7420 (N_7420,N_4945,N_4365);
or U7421 (N_7421,N_4278,N_4187);
or U7422 (N_7422,N_4290,N_5328);
and U7423 (N_7423,N_5814,N_5014);
xor U7424 (N_7424,N_4559,N_5071);
and U7425 (N_7425,N_5403,N_5517);
or U7426 (N_7426,N_4409,N_4251);
nor U7427 (N_7427,N_5415,N_4521);
nor U7428 (N_7428,N_4498,N_4104);
xnor U7429 (N_7429,N_5457,N_4584);
nor U7430 (N_7430,N_4613,N_4784);
nor U7431 (N_7431,N_4412,N_4129);
and U7432 (N_7432,N_5692,N_5630);
nor U7433 (N_7433,N_4992,N_5344);
xor U7434 (N_7434,N_4640,N_5725);
nor U7435 (N_7435,N_4587,N_4250);
nor U7436 (N_7436,N_5439,N_4059);
nand U7437 (N_7437,N_5366,N_5465);
and U7438 (N_7438,N_4762,N_5180);
and U7439 (N_7439,N_4258,N_4517);
xnor U7440 (N_7440,N_4101,N_4314);
xnor U7441 (N_7441,N_4137,N_4218);
nor U7442 (N_7442,N_5783,N_4281);
nor U7443 (N_7443,N_4922,N_5607);
nand U7444 (N_7444,N_5526,N_5794);
and U7445 (N_7445,N_5812,N_4944);
and U7446 (N_7446,N_5914,N_4262);
or U7447 (N_7447,N_5749,N_5778);
nor U7448 (N_7448,N_4261,N_4553);
or U7449 (N_7449,N_5462,N_4187);
xnor U7450 (N_7450,N_5145,N_5498);
or U7451 (N_7451,N_5725,N_5898);
xnor U7452 (N_7452,N_5312,N_4553);
xor U7453 (N_7453,N_5293,N_4789);
nor U7454 (N_7454,N_4608,N_4671);
nor U7455 (N_7455,N_4688,N_5680);
nor U7456 (N_7456,N_5122,N_5611);
or U7457 (N_7457,N_4423,N_5712);
xor U7458 (N_7458,N_5167,N_4228);
nor U7459 (N_7459,N_5827,N_4043);
nand U7460 (N_7460,N_5171,N_4468);
nand U7461 (N_7461,N_5425,N_4351);
nor U7462 (N_7462,N_4283,N_5724);
xor U7463 (N_7463,N_5971,N_5097);
nand U7464 (N_7464,N_5657,N_5524);
nand U7465 (N_7465,N_5309,N_5402);
nand U7466 (N_7466,N_4378,N_4561);
xor U7467 (N_7467,N_5986,N_5590);
nand U7468 (N_7468,N_5159,N_4976);
or U7469 (N_7469,N_4497,N_5646);
nor U7470 (N_7470,N_5631,N_5674);
or U7471 (N_7471,N_5696,N_5982);
nand U7472 (N_7472,N_4496,N_5033);
nand U7473 (N_7473,N_4023,N_5331);
and U7474 (N_7474,N_4931,N_5246);
nor U7475 (N_7475,N_5377,N_4233);
or U7476 (N_7476,N_4878,N_5783);
xor U7477 (N_7477,N_4136,N_4978);
nand U7478 (N_7478,N_5145,N_5806);
or U7479 (N_7479,N_4204,N_4323);
nand U7480 (N_7480,N_4140,N_5651);
nor U7481 (N_7481,N_5032,N_5150);
and U7482 (N_7482,N_4566,N_5480);
xor U7483 (N_7483,N_4422,N_5757);
or U7484 (N_7484,N_4931,N_4398);
nor U7485 (N_7485,N_4902,N_5356);
nor U7486 (N_7486,N_5009,N_5068);
nor U7487 (N_7487,N_4836,N_5799);
xnor U7488 (N_7488,N_4231,N_5324);
xor U7489 (N_7489,N_5955,N_5132);
xnor U7490 (N_7490,N_4470,N_5971);
nor U7491 (N_7491,N_5431,N_5939);
or U7492 (N_7492,N_4456,N_5398);
nor U7493 (N_7493,N_4267,N_4752);
xor U7494 (N_7494,N_4545,N_4366);
or U7495 (N_7495,N_5891,N_5319);
or U7496 (N_7496,N_5206,N_5893);
xnor U7497 (N_7497,N_5047,N_4725);
nand U7498 (N_7498,N_5247,N_4685);
nor U7499 (N_7499,N_4104,N_5523);
and U7500 (N_7500,N_5480,N_4252);
nand U7501 (N_7501,N_5031,N_5546);
xor U7502 (N_7502,N_5579,N_4612);
and U7503 (N_7503,N_4827,N_5423);
or U7504 (N_7504,N_5747,N_4155);
and U7505 (N_7505,N_4421,N_5707);
and U7506 (N_7506,N_5923,N_4509);
nor U7507 (N_7507,N_5960,N_5864);
xnor U7508 (N_7508,N_5590,N_4231);
nor U7509 (N_7509,N_4838,N_4982);
and U7510 (N_7510,N_5688,N_5331);
and U7511 (N_7511,N_5750,N_5290);
xor U7512 (N_7512,N_5665,N_5365);
nand U7513 (N_7513,N_4643,N_5781);
and U7514 (N_7514,N_4468,N_5662);
xnor U7515 (N_7515,N_4122,N_5325);
xor U7516 (N_7516,N_5088,N_4443);
or U7517 (N_7517,N_4035,N_4136);
nand U7518 (N_7518,N_5511,N_4044);
nor U7519 (N_7519,N_5676,N_5958);
and U7520 (N_7520,N_5399,N_5095);
and U7521 (N_7521,N_4648,N_4777);
nand U7522 (N_7522,N_5927,N_5000);
nor U7523 (N_7523,N_5190,N_5191);
or U7524 (N_7524,N_4954,N_4830);
xnor U7525 (N_7525,N_5141,N_5130);
nor U7526 (N_7526,N_5336,N_4031);
or U7527 (N_7527,N_4540,N_5889);
or U7528 (N_7528,N_4792,N_5366);
nor U7529 (N_7529,N_4188,N_5290);
xor U7530 (N_7530,N_4975,N_5932);
or U7531 (N_7531,N_4486,N_5667);
or U7532 (N_7532,N_4931,N_4731);
nand U7533 (N_7533,N_4935,N_5671);
nand U7534 (N_7534,N_5158,N_5787);
xnor U7535 (N_7535,N_5652,N_4527);
or U7536 (N_7536,N_4755,N_5646);
or U7537 (N_7537,N_5949,N_4949);
and U7538 (N_7538,N_5515,N_4151);
or U7539 (N_7539,N_5507,N_4420);
nor U7540 (N_7540,N_5082,N_5759);
xnor U7541 (N_7541,N_5009,N_4539);
xor U7542 (N_7542,N_4659,N_5932);
or U7543 (N_7543,N_4514,N_4861);
or U7544 (N_7544,N_4223,N_4248);
or U7545 (N_7545,N_5817,N_4393);
nand U7546 (N_7546,N_5079,N_5896);
nor U7547 (N_7547,N_5050,N_5455);
or U7548 (N_7548,N_4070,N_5665);
nand U7549 (N_7549,N_5714,N_5114);
and U7550 (N_7550,N_5260,N_4318);
xor U7551 (N_7551,N_5668,N_5490);
nor U7552 (N_7552,N_5175,N_5696);
nand U7553 (N_7553,N_4864,N_4498);
and U7554 (N_7554,N_4733,N_5254);
nor U7555 (N_7555,N_5624,N_4444);
xnor U7556 (N_7556,N_5694,N_5165);
nor U7557 (N_7557,N_4812,N_5393);
xor U7558 (N_7558,N_5303,N_4731);
or U7559 (N_7559,N_4068,N_4399);
nor U7560 (N_7560,N_4653,N_4318);
nor U7561 (N_7561,N_4362,N_5178);
and U7562 (N_7562,N_4875,N_5276);
nand U7563 (N_7563,N_5089,N_5428);
nand U7564 (N_7564,N_4587,N_5531);
or U7565 (N_7565,N_4188,N_5432);
and U7566 (N_7566,N_5704,N_5731);
or U7567 (N_7567,N_5824,N_5406);
nor U7568 (N_7568,N_5383,N_5840);
nand U7569 (N_7569,N_5339,N_5514);
xnor U7570 (N_7570,N_4599,N_5813);
and U7571 (N_7571,N_4915,N_5259);
nand U7572 (N_7572,N_4092,N_5880);
nor U7573 (N_7573,N_5055,N_5833);
xnor U7574 (N_7574,N_4330,N_4436);
or U7575 (N_7575,N_5961,N_4883);
nor U7576 (N_7576,N_5264,N_4557);
or U7577 (N_7577,N_4649,N_4079);
nand U7578 (N_7578,N_4707,N_4612);
nor U7579 (N_7579,N_5816,N_4597);
xor U7580 (N_7580,N_4602,N_4445);
and U7581 (N_7581,N_5439,N_5646);
and U7582 (N_7582,N_4297,N_5350);
nand U7583 (N_7583,N_4016,N_4483);
xnor U7584 (N_7584,N_5342,N_5246);
and U7585 (N_7585,N_4885,N_4491);
and U7586 (N_7586,N_5639,N_5900);
and U7587 (N_7587,N_5452,N_5885);
nor U7588 (N_7588,N_4862,N_4299);
and U7589 (N_7589,N_5428,N_5592);
and U7590 (N_7590,N_5528,N_4373);
nand U7591 (N_7591,N_4752,N_4190);
and U7592 (N_7592,N_4624,N_4278);
nand U7593 (N_7593,N_5868,N_5645);
nor U7594 (N_7594,N_5552,N_5898);
xnor U7595 (N_7595,N_4462,N_4704);
xor U7596 (N_7596,N_5243,N_5167);
xnor U7597 (N_7597,N_4314,N_4366);
nand U7598 (N_7598,N_5308,N_5163);
nor U7599 (N_7599,N_5899,N_5195);
nor U7600 (N_7600,N_5637,N_5490);
nand U7601 (N_7601,N_4864,N_5414);
and U7602 (N_7602,N_5783,N_5025);
or U7603 (N_7603,N_4395,N_5339);
or U7604 (N_7604,N_5485,N_4514);
and U7605 (N_7605,N_5572,N_4408);
or U7606 (N_7606,N_5583,N_5033);
or U7607 (N_7607,N_4607,N_4223);
and U7608 (N_7608,N_5740,N_5743);
or U7609 (N_7609,N_4266,N_5851);
and U7610 (N_7610,N_4047,N_5127);
nor U7611 (N_7611,N_5426,N_4112);
xnor U7612 (N_7612,N_4218,N_5957);
or U7613 (N_7613,N_4970,N_5489);
xnor U7614 (N_7614,N_5983,N_5735);
xnor U7615 (N_7615,N_4047,N_4356);
xnor U7616 (N_7616,N_5774,N_5147);
xor U7617 (N_7617,N_5140,N_5669);
nand U7618 (N_7618,N_4139,N_5633);
and U7619 (N_7619,N_5676,N_4421);
nand U7620 (N_7620,N_4293,N_5652);
and U7621 (N_7621,N_4518,N_4076);
nand U7622 (N_7622,N_4631,N_5267);
or U7623 (N_7623,N_5666,N_5100);
nor U7624 (N_7624,N_4611,N_5001);
nor U7625 (N_7625,N_5065,N_4633);
and U7626 (N_7626,N_5892,N_4076);
xor U7627 (N_7627,N_4287,N_5783);
or U7628 (N_7628,N_4131,N_4167);
nand U7629 (N_7629,N_5010,N_5124);
or U7630 (N_7630,N_5543,N_5477);
or U7631 (N_7631,N_4719,N_4641);
or U7632 (N_7632,N_5868,N_4415);
and U7633 (N_7633,N_4324,N_4002);
or U7634 (N_7634,N_4987,N_4586);
nor U7635 (N_7635,N_4614,N_5581);
nor U7636 (N_7636,N_4205,N_4151);
and U7637 (N_7637,N_5415,N_5771);
and U7638 (N_7638,N_4977,N_4786);
xor U7639 (N_7639,N_4131,N_5644);
xnor U7640 (N_7640,N_5508,N_4709);
or U7641 (N_7641,N_5262,N_5221);
nor U7642 (N_7642,N_4297,N_5045);
and U7643 (N_7643,N_5176,N_5075);
or U7644 (N_7644,N_5664,N_4654);
and U7645 (N_7645,N_4370,N_5734);
or U7646 (N_7646,N_4837,N_4944);
nand U7647 (N_7647,N_4749,N_4718);
or U7648 (N_7648,N_5767,N_5307);
xor U7649 (N_7649,N_4019,N_5707);
nand U7650 (N_7650,N_4341,N_5820);
xnor U7651 (N_7651,N_4684,N_4580);
nor U7652 (N_7652,N_4992,N_5553);
nand U7653 (N_7653,N_4771,N_4934);
or U7654 (N_7654,N_5347,N_4083);
or U7655 (N_7655,N_4483,N_5468);
nand U7656 (N_7656,N_4264,N_4326);
nand U7657 (N_7657,N_5639,N_4738);
or U7658 (N_7658,N_4545,N_4186);
or U7659 (N_7659,N_5164,N_4521);
or U7660 (N_7660,N_5490,N_4864);
nand U7661 (N_7661,N_5577,N_5497);
nand U7662 (N_7662,N_4052,N_5484);
and U7663 (N_7663,N_5438,N_4788);
nor U7664 (N_7664,N_5459,N_4565);
nand U7665 (N_7665,N_5678,N_4641);
and U7666 (N_7666,N_5375,N_4650);
or U7667 (N_7667,N_4484,N_5645);
nor U7668 (N_7668,N_4385,N_4572);
xor U7669 (N_7669,N_4411,N_4874);
nor U7670 (N_7670,N_5249,N_5107);
or U7671 (N_7671,N_5215,N_5179);
or U7672 (N_7672,N_4729,N_4745);
or U7673 (N_7673,N_4212,N_4203);
nor U7674 (N_7674,N_5435,N_5693);
or U7675 (N_7675,N_4334,N_5765);
xor U7676 (N_7676,N_5899,N_5093);
nor U7677 (N_7677,N_4349,N_4093);
nand U7678 (N_7678,N_4210,N_5723);
and U7679 (N_7679,N_5956,N_5972);
nand U7680 (N_7680,N_5467,N_4200);
xnor U7681 (N_7681,N_5298,N_5572);
nor U7682 (N_7682,N_5327,N_4505);
and U7683 (N_7683,N_5349,N_4374);
xor U7684 (N_7684,N_5038,N_5166);
nor U7685 (N_7685,N_4205,N_5961);
xnor U7686 (N_7686,N_4613,N_5065);
or U7687 (N_7687,N_5363,N_5580);
or U7688 (N_7688,N_4686,N_5214);
and U7689 (N_7689,N_4960,N_5780);
nor U7690 (N_7690,N_4826,N_4192);
nand U7691 (N_7691,N_4538,N_4241);
xnor U7692 (N_7692,N_4274,N_5862);
and U7693 (N_7693,N_4600,N_4859);
and U7694 (N_7694,N_5139,N_5148);
and U7695 (N_7695,N_4696,N_4371);
nor U7696 (N_7696,N_5376,N_4801);
nor U7697 (N_7697,N_5898,N_4862);
and U7698 (N_7698,N_4984,N_4725);
and U7699 (N_7699,N_5485,N_5576);
xnor U7700 (N_7700,N_4451,N_4504);
or U7701 (N_7701,N_4587,N_5017);
or U7702 (N_7702,N_4399,N_5001);
xor U7703 (N_7703,N_4401,N_4477);
or U7704 (N_7704,N_5314,N_4515);
nand U7705 (N_7705,N_4905,N_4504);
nand U7706 (N_7706,N_4849,N_4615);
or U7707 (N_7707,N_5439,N_5210);
xnor U7708 (N_7708,N_5114,N_5824);
xnor U7709 (N_7709,N_4980,N_5737);
xor U7710 (N_7710,N_5380,N_5554);
nor U7711 (N_7711,N_5784,N_5002);
or U7712 (N_7712,N_5923,N_5656);
xnor U7713 (N_7713,N_5324,N_4941);
nand U7714 (N_7714,N_4288,N_5041);
xor U7715 (N_7715,N_4259,N_5532);
or U7716 (N_7716,N_4486,N_4302);
nor U7717 (N_7717,N_4334,N_5537);
xor U7718 (N_7718,N_4802,N_4027);
nor U7719 (N_7719,N_4086,N_5550);
nand U7720 (N_7720,N_5080,N_4363);
and U7721 (N_7721,N_5524,N_4181);
xor U7722 (N_7722,N_5912,N_4651);
xor U7723 (N_7723,N_5613,N_5042);
nor U7724 (N_7724,N_4826,N_5661);
and U7725 (N_7725,N_4121,N_5536);
xnor U7726 (N_7726,N_4680,N_5713);
nor U7727 (N_7727,N_5306,N_5012);
nand U7728 (N_7728,N_5499,N_5932);
and U7729 (N_7729,N_4443,N_4923);
nand U7730 (N_7730,N_4147,N_5937);
xnor U7731 (N_7731,N_4226,N_4012);
or U7732 (N_7732,N_5669,N_4670);
and U7733 (N_7733,N_4246,N_5333);
xnor U7734 (N_7734,N_4390,N_5333);
nor U7735 (N_7735,N_4307,N_4357);
nor U7736 (N_7736,N_4991,N_4511);
nand U7737 (N_7737,N_5987,N_5699);
or U7738 (N_7738,N_5193,N_5795);
and U7739 (N_7739,N_4337,N_5623);
or U7740 (N_7740,N_5320,N_5656);
xor U7741 (N_7741,N_5566,N_4718);
nor U7742 (N_7742,N_4912,N_5225);
or U7743 (N_7743,N_5518,N_5876);
nor U7744 (N_7744,N_5736,N_5648);
xor U7745 (N_7745,N_4925,N_4402);
or U7746 (N_7746,N_4965,N_5938);
nand U7747 (N_7747,N_5212,N_4605);
nand U7748 (N_7748,N_4194,N_5647);
xor U7749 (N_7749,N_4037,N_4838);
or U7750 (N_7750,N_4293,N_5158);
and U7751 (N_7751,N_4646,N_5240);
nand U7752 (N_7752,N_5490,N_4652);
xnor U7753 (N_7753,N_5762,N_4781);
or U7754 (N_7754,N_4342,N_5587);
xor U7755 (N_7755,N_5508,N_4412);
nor U7756 (N_7756,N_5434,N_4168);
nand U7757 (N_7757,N_4314,N_4821);
nor U7758 (N_7758,N_5271,N_5531);
or U7759 (N_7759,N_4240,N_5184);
xor U7760 (N_7760,N_4354,N_4146);
nor U7761 (N_7761,N_4024,N_5377);
nor U7762 (N_7762,N_4240,N_4140);
nand U7763 (N_7763,N_5689,N_5248);
nand U7764 (N_7764,N_5897,N_4788);
or U7765 (N_7765,N_5672,N_4221);
or U7766 (N_7766,N_5973,N_4869);
xnor U7767 (N_7767,N_4789,N_5348);
xor U7768 (N_7768,N_4593,N_4125);
nor U7769 (N_7769,N_4794,N_5531);
xnor U7770 (N_7770,N_4068,N_4001);
or U7771 (N_7771,N_4901,N_5793);
or U7772 (N_7772,N_5366,N_5642);
and U7773 (N_7773,N_4710,N_4907);
and U7774 (N_7774,N_4895,N_4296);
xnor U7775 (N_7775,N_4375,N_4463);
or U7776 (N_7776,N_5413,N_4190);
xor U7777 (N_7777,N_5165,N_4330);
nand U7778 (N_7778,N_5353,N_4921);
and U7779 (N_7779,N_4896,N_5231);
or U7780 (N_7780,N_4907,N_4775);
nand U7781 (N_7781,N_5875,N_5251);
nand U7782 (N_7782,N_5756,N_5438);
nand U7783 (N_7783,N_5007,N_4906);
xor U7784 (N_7784,N_5594,N_4858);
nand U7785 (N_7785,N_4031,N_4775);
nand U7786 (N_7786,N_4184,N_5830);
or U7787 (N_7787,N_5526,N_4139);
and U7788 (N_7788,N_5055,N_4923);
nor U7789 (N_7789,N_5146,N_5832);
nand U7790 (N_7790,N_5394,N_5053);
nand U7791 (N_7791,N_4354,N_5432);
nor U7792 (N_7792,N_4641,N_5355);
or U7793 (N_7793,N_4517,N_4631);
nand U7794 (N_7794,N_4613,N_4932);
and U7795 (N_7795,N_4380,N_5006);
nand U7796 (N_7796,N_5068,N_5363);
nand U7797 (N_7797,N_4602,N_4431);
and U7798 (N_7798,N_4844,N_4783);
nor U7799 (N_7799,N_4860,N_4762);
xnor U7800 (N_7800,N_4559,N_4536);
or U7801 (N_7801,N_4640,N_4012);
xor U7802 (N_7802,N_4261,N_5642);
nand U7803 (N_7803,N_4011,N_4692);
or U7804 (N_7804,N_5452,N_4778);
nand U7805 (N_7805,N_5051,N_4260);
nand U7806 (N_7806,N_4809,N_5632);
or U7807 (N_7807,N_5013,N_5271);
and U7808 (N_7808,N_5884,N_5088);
xnor U7809 (N_7809,N_4245,N_5029);
or U7810 (N_7810,N_5726,N_5405);
nand U7811 (N_7811,N_5957,N_4744);
nand U7812 (N_7812,N_5602,N_5728);
xor U7813 (N_7813,N_4031,N_5095);
xnor U7814 (N_7814,N_4557,N_5915);
xor U7815 (N_7815,N_5501,N_4301);
nor U7816 (N_7816,N_5478,N_4817);
and U7817 (N_7817,N_4594,N_4857);
nand U7818 (N_7818,N_4239,N_5943);
nand U7819 (N_7819,N_5877,N_4820);
nand U7820 (N_7820,N_4661,N_5562);
and U7821 (N_7821,N_4229,N_4417);
nand U7822 (N_7822,N_4677,N_4334);
nor U7823 (N_7823,N_5643,N_5199);
and U7824 (N_7824,N_5620,N_4306);
nand U7825 (N_7825,N_4086,N_4294);
or U7826 (N_7826,N_5019,N_4740);
nor U7827 (N_7827,N_5126,N_5448);
xnor U7828 (N_7828,N_5363,N_4808);
xor U7829 (N_7829,N_5922,N_4392);
nand U7830 (N_7830,N_5570,N_5140);
and U7831 (N_7831,N_5065,N_4268);
nand U7832 (N_7832,N_4934,N_5002);
nand U7833 (N_7833,N_4113,N_5731);
and U7834 (N_7834,N_4234,N_4662);
xnor U7835 (N_7835,N_4577,N_4158);
nand U7836 (N_7836,N_4409,N_4133);
nand U7837 (N_7837,N_4807,N_4851);
nand U7838 (N_7838,N_4429,N_4785);
and U7839 (N_7839,N_4272,N_5234);
nor U7840 (N_7840,N_4819,N_4248);
nor U7841 (N_7841,N_5662,N_4125);
and U7842 (N_7842,N_5004,N_4400);
nand U7843 (N_7843,N_4791,N_4954);
xnor U7844 (N_7844,N_5495,N_4520);
or U7845 (N_7845,N_4202,N_5805);
nand U7846 (N_7846,N_4071,N_4562);
xor U7847 (N_7847,N_4243,N_5405);
nand U7848 (N_7848,N_5504,N_5945);
nand U7849 (N_7849,N_4752,N_5588);
nor U7850 (N_7850,N_4775,N_4250);
xnor U7851 (N_7851,N_4582,N_4326);
nand U7852 (N_7852,N_4920,N_5032);
or U7853 (N_7853,N_4897,N_4685);
nor U7854 (N_7854,N_4920,N_5778);
xnor U7855 (N_7855,N_4853,N_5853);
xor U7856 (N_7856,N_5497,N_5587);
or U7857 (N_7857,N_5714,N_4646);
xor U7858 (N_7858,N_5608,N_4613);
xor U7859 (N_7859,N_4671,N_5697);
nand U7860 (N_7860,N_4516,N_5376);
nand U7861 (N_7861,N_4648,N_5385);
or U7862 (N_7862,N_5173,N_4826);
and U7863 (N_7863,N_5263,N_5679);
nor U7864 (N_7864,N_4660,N_5353);
and U7865 (N_7865,N_5390,N_4500);
or U7866 (N_7866,N_4401,N_5429);
and U7867 (N_7867,N_5584,N_5889);
or U7868 (N_7868,N_5048,N_4909);
nor U7869 (N_7869,N_5907,N_5605);
xor U7870 (N_7870,N_4158,N_5795);
xnor U7871 (N_7871,N_5858,N_4919);
nor U7872 (N_7872,N_4852,N_4913);
nand U7873 (N_7873,N_5189,N_5554);
nor U7874 (N_7874,N_4906,N_4879);
and U7875 (N_7875,N_5954,N_5411);
nand U7876 (N_7876,N_4675,N_5451);
or U7877 (N_7877,N_4158,N_4677);
and U7878 (N_7878,N_4648,N_4806);
and U7879 (N_7879,N_4959,N_4568);
and U7880 (N_7880,N_4479,N_4105);
nand U7881 (N_7881,N_5112,N_5496);
nand U7882 (N_7882,N_4981,N_4139);
nand U7883 (N_7883,N_4372,N_5990);
nand U7884 (N_7884,N_5205,N_5436);
nor U7885 (N_7885,N_4611,N_4778);
nor U7886 (N_7886,N_4412,N_4793);
or U7887 (N_7887,N_5938,N_4688);
nor U7888 (N_7888,N_4044,N_4425);
or U7889 (N_7889,N_4795,N_4107);
and U7890 (N_7890,N_4747,N_5718);
nor U7891 (N_7891,N_4690,N_4656);
nor U7892 (N_7892,N_5624,N_4227);
xor U7893 (N_7893,N_4687,N_4841);
xor U7894 (N_7894,N_4682,N_4351);
xnor U7895 (N_7895,N_5078,N_4615);
xnor U7896 (N_7896,N_4188,N_4245);
or U7897 (N_7897,N_5488,N_5268);
or U7898 (N_7898,N_5374,N_5114);
and U7899 (N_7899,N_4330,N_5523);
nand U7900 (N_7900,N_5172,N_4734);
and U7901 (N_7901,N_4152,N_4633);
nand U7902 (N_7902,N_5863,N_5105);
and U7903 (N_7903,N_5325,N_4087);
and U7904 (N_7904,N_5976,N_5331);
xnor U7905 (N_7905,N_5212,N_5985);
and U7906 (N_7906,N_4282,N_4435);
xnor U7907 (N_7907,N_5929,N_4749);
nor U7908 (N_7908,N_4425,N_5693);
or U7909 (N_7909,N_5489,N_4095);
and U7910 (N_7910,N_4982,N_4065);
and U7911 (N_7911,N_4919,N_5876);
and U7912 (N_7912,N_5454,N_5006);
xor U7913 (N_7913,N_5347,N_5249);
nor U7914 (N_7914,N_5352,N_5666);
nand U7915 (N_7915,N_5397,N_5122);
nand U7916 (N_7916,N_5032,N_5182);
or U7917 (N_7917,N_4834,N_4404);
nand U7918 (N_7918,N_5970,N_4784);
xor U7919 (N_7919,N_4719,N_4383);
xnor U7920 (N_7920,N_5723,N_4369);
nor U7921 (N_7921,N_5607,N_5527);
xnor U7922 (N_7922,N_5350,N_4824);
nor U7923 (N_7923,N_5339,N_4719);
and U7924 (N_7924,N_5056,N_4469);
nor U7925 (N_7925,N_4895,N_5087);
or U7926 (N_7926,N_4340,N_4904);
xnor U7927 (N_7927,N_4228,N_5873);
and U7928 (N_7928,N_5128,N_4024);
or U7929 (N_7929,N_5076,N_5177);
or U7930 (N_7930,N_4794,N_4770);
nand U7931 (N_7931,N_5842,N_4707);
nand U7932 (N_7932,N_4051,N_5903);
nand U7933 (N_7933,N_4032,N_4825);
and U7934 (N_7934,N_5035,N_4684);
xor U7935 (N_7935,N_5142,N_5800);
and U7936 (N_7936,N_4505,N_4995);
or U7937 (N_7937,N_4616,N_5721);
or U7938 (N_7938,N_4532,N_5109);
and U7939 (N_7939,N_4856,N_5332);
nand U7940 (N_7940,N_5810,N_5450);
or U7941 (N_7941,N_4341,N_5891);
nor U7942 (N_7942,N_4494,N_5428);
nand U7943 (N_7943,N_5775,N_4673);
and U7944 (N_7944,N_5373,N_5857);
nand U7945 (N_7945,N_4015,N_5095);
nand U7946 (N_7946,N_4004,N_4618);
and U7947 (N_7947,N_4787,N_4783);
xor U7948 (N_7948,N_4149,N_4669);
nand U7949 (N_7949,N_5160,N_4451);
nand U7950 (N_7950,N_4719,N_5875);
nand U7951 (N_7951,N_5855,N_4037);
xor U7952 (N_7952,N_4085,N_4434);
and U7953 (N_7953,N_4075,N_5540);
nor U7954 (N_7954,N_5496,N_4246);
nor U7955 (N_7955,N_4918,N_5367);
and U7956 (N_7956,N_5685,N_4806);
nor U7957 (N_7957,N_5717,N_5206);
or U7958 (N_7958,N_4771,N_4545);
and U7959 (N_7959,N_5241,N_5774);
xor U7960 (N_7960,N_5003,N_5664);
nand U7961 (N_7961,N_4253,N_4824);
and U7962 (N_7962,N_4916,N_4566);
or U7963 (N_7963,N_4090,N_4251);
nor U7964 (N_7964,N_5350,N_4049);
nand U7965 (N_7965,N_4295,N_5626);
nand U7966 (N_7966,N_4848,N_4519);
nand U7967 (N_7967,N_4575,N_4305);
xor U7968 (N_7968,N_4571,N_5950);
xnor U7969 (N_7969,N_5336,N_4356);
xor U7970 (N_7970,N_4774,N_5075);
and U7971 (N_7971,N_5205,N_5952);
or U7972 (N_7972,N_4925,N_4431);
xor U7973 (N_7973,N_5043,N_4087);
xor U7974 (N_7974,N_4552,N_5475);
nand U7975 (N_7975,N_4725,N_5024);
xor U7976 (N_7976,N_4602,N_5320);
xnor U7977 (N_7977,N_4926,N_5870);
nand U7978 (N_7978,N_5601,N_5545);
xnor U7979 (N_7979,N_5781,N_5343);
and U7980 (N_7980,N_5914,N_4355);
nor U7981 (N_7981,N_4717,N_4977);
xor U7982 (N_7982,N_4246,N_5654);
xnor U7983 (N_7983,N_4329,N_5037);
nand U7984 (N_7984,N_4292,N_5234);
nor U7985 (N_7985,N_5292,N_4881);
or U7986 (N_7986,N_4372,N_4368);
xnor U7987 (N_7987,N_5275,N_4877);
nor U7988 (N_7988,N_5958,N_4857);
and U7989 (N_7989,N_4247,N_4937);
nor U7990 (N_7990,N_4001,N_5816);
or U7991 (N_7991,N_5298,N_5957);
nand U7992 (N_7992,N_5865,N_5401);
or U7993 (N_7993,N_5091,N_4821);
or U7994 (N_7994,N_5970,N_5832);
nand U7995 (N_7995,N_4813,N_5057);
or U7996 (N_7996,N_5826,N_4438);
or U7997 (N_7997,N_5179,N_4240);
and U7998 (N_7998,N_4527,N_5202);
and U7999 (N_7999,N_4971,N_4049);
nor U8000 (N_8000,N_7079,N_6371);
or U8001 (N_8001,N_7023,N_7809);
and U8002 (N_8002,N_7498,N_7125);
nor U8003 (N_8003,N_7010,N_7654);
nand U8004 (N_8004,N_7698,N_7115);
nor U8005 (N_8005,N_6131,N_6378);
and U8006 (N_8006,N_6989,N_7135);
nand U8007 (N_8007,N_6412,N_7148);
or U8008 (N_8008,N_7676,N_7393);
and U8009 (N_8009,N_7949,N_7098);
xor U8010 (N_8010,N_7215,N_7122);
nor U8011 (N_8011,N_7857,N_7780);
xor U8012 (N_8012,N_6260,N_6076);
and U8013 (N_8013,N_6703,N_6618);
nand U8014 (N_8014,N_6704,N_7826);
nand U8015 (N_8015,N_6723,N_7419);
or U8016 (N_8016,N_7439,N_7110);
xnor U8017 (N_8017,N_6708,N_7585);
and U8018 (N_8018,N_7161,N_7308);
and U8019 (N_8019,N_7164,N_6885);
or U8020 (N_8020,N_6475,N_6360);
nor U8021 (N_8021,N_6546,N_6870);
and U8022 (N_8022,N_6971,N_7539);
and U8023 (N_8023,N_7262,N_7845);
and U8024 (N_8024,N_7095,N_6983);
nand U8025 (N_8025,N_7825,N_7877);
nand U8026 (N_8026,N_6092,N_7785);
xor U8027 (N_8027,N_7324,N_7758);
nand U8028 (N_8028,N_6910,N_6702);
nor U8029 (N_8029,N_7211,N_7688);
or U8030 (N_8030,N_7093,N_6447);
nand U8031 (N_8031,N_7740,N_7330);
or U8032 (N_8032,N_6202,N_7796);
nor U8033 (N_8033,N_6537,N_6341);
xor U8034 (N_8034,N_7987,N_7045);
and U8035 (N_8035,N_7918,N_6269);
nor U8036 (N_8036,N_7528,N_6113);
and U8037 (N_8037,N_6856,N_7313);
and U8038 (N_8038,N_7241,N_6329);
or U8039 (N_8039,N_7179,N_6535);
nand U8040 (N_8040,N_6163,N_7423);
nand U8041 (N_8041,N_7936,N_7154);
and U8042 (N_8042,N_6289,N_6459);
nand U8043 (N_8043,N_6957,N_6352);
xor U8044 (N_8044,N_7917,N_7605);
nor U8045 (N_8045,N_6011,N_6886);
xor U8046 (N_8046,N_6993,N_7775);
or U8047 (N_8047,N_6224,N_6650);
nand U8048 (N_8048,N_6351,N_6954);
xnor U8049 (N_8049,N_6848,N_6130);
nand U8050 (N_8050,N_7896,N_7645);
xnor U8051 (N_8051,N_6861,N_7943);
or U8052 (N_8052,N_7513,N_6062);
and U8053 (N_8053,N_6466,N_7805);
xor U8054 (N_8054,N_7881,N_7459);
nand U8055 (N_8055,N_7505,N_6832);
xnor U8056 (N_8056,N_7047,N_6860);
nand U8057 (N_8057,N_7575,N_6917);
nand U8058 (N_8058,N_7409,N_6345);
and U8059 (N_8059,N_7374,N_6323);
nor U8060 (N_8060,N_7819,N_6803);
and U8061 (N_8061,N_7042,N_6806);
nor U8062 (N_8062,N_6476,N_7567);
nand U8063 (N_8063,N_6791,N_7601);
nand U8064 (N_8064,N_6183,N_7523);
xor U8065 (N_8065,N_7352,N_7894);
xor U8066 (N_8066,N_7387,N_7149);
or U8067 (N_8067,N_7248,N_6616);
or U8068 (N_8068,N_7677,N_6127);
xnor U8069 (N_8069,N_7971,N_6544);
xnor U8070 (N_8070,N_6456,N_6668);
or U8071 (N_8071,N_7469,N_6816);
nand U8072 (N_8072,N_6750,N_6500);
and U8073 (N_8073,N_7976,N_7991);
nor U8074 (N_8074,N_6659,N_7369);
or U8075 (N_8075,N_7684,N_7245);
xor U8076 (N_8076,N_6357,N_7472);
nand U8077 (N_8077,N_6242,N_7269);
xor U8078 (N_8078,N_6675,N_7964);
nand U8079 (N_8079,N_7617,N_7680);
or U8080 (N_8080,N_6842,N_6599);
nor U8081 (N_8081,N_7574,N_6373);
and U8082 (N_8082,N_6006,N_7293);
and U8083 (N_8083,N_6140,N_6218);
xnor U8084 (N_8084,N_7221,N_6731);
nand U8085 (N_8085,N_6562,N_7589);
and U8086 (N_8086,N_7531,N_7781);
nor U8087 (N_8087,N_7348,N_7616);
xnor U8088 (N_8088,N_6829,N_6319);
or U8089 (N_8089,N_6013,N_7041);
and U8090 (N_8090,N_6785,N_7163);
or U8091 (N_8091,N_6206,N_6815);
or U8092 (N_8092,N_6729,N_6875);
nor U8093 (N_8093,N_7464,N_7001);
xor U8094 (N_8094,N_7265,N_6233);
xor U8095 (N_8095,N_7033,N_6058);
or U8096 (N_8096,N_6464,N_6307);
nand U8097 (N_8097,N_7365,N_6123);
xor U8098 (N_8098,N_6317,N_6027);
xor U8099 (N_8099,N_6952,N_7608);
nor U8100 (N_8100,N_6980,N_7948);
or U8101 (N_8101,N_7104,N_6024);
or U8102 (N_8102,N_6671,N_7715);
xor U8103 (N_8103,N_6697,N_6580);
xor U8104 (N_8104,N_7633,N_7686);
and U8105 (N_8105,N_7415,N_6448);
xnor U8106 (N_8106,N_7160,N_7279);
nand U8107 (N_8107,N_7870,N_6662);
or U8108 (N_8108,N_7776,N_6947);
nand U8109 (N_8109,N_7711,N_7708);
nor U8110 (N_8110,N_7481,N_6333);
xor U8111 (N_8111,N_6121,N_6590);
or U8112 (N_8112,N_6921,N_7180);
and U8113 (N_8113,N_7206,N_6926);
xnor U8114 (N_8114,N_7418,N_6962);
nand U8115 (N_8115,N_6800,N_7841);
xor U8116 (N_8116,N_7673,N_7290);
or U8117 (N_8117,N_6372,N_6442);
nand U8118 (N_8118,N_7391,N_7468);
nand U8119 (N_8119,N_6724,N_6730);
nor U8120 (N_8120,N_6934,N_6126);
or U8121 (N_8121,N_7128,N_6699);
and U8122 (N_8122,N_7900,N_6304);
nor U8123 (N_8123,N_7882,N_6310);
or U8124 (N_8124,N_7671,N_6541);
nand U8125 (N_8125,N_6502,N_7187);
nor U8126 (N_8126,N_7101,N_7636);
and U8127 (N_8127,N_7925,N_6085);
xnor U8128 (N_8128,N_7013,N_7901);
nand U8129 (N_8129,N_7386,N_6821);
xnor U8130 (N_8130,N_6920,N_6505);
or U8131 (N_8131,N_6690,N_6632);
and U8132 (N_8132,N_6658,N_6843);
and U8133 (N_8133,N_7938,N_7015);
or U8134 (N_8134,N_7621,N_6775);
nor U8135 (N_8135,N_7861,N_6814);
nand U8136 (N_8136,N_6460,N_7962);
and U8137 (N_8137,N_7650,N_7993);
and U8138 (N_8138,N_6823,N_7849);
or U8139 (N_8139,N_6471,N_6879);
nor U8140 (N_8140,N_6779,N_6941);
and U8141 (N_8141,N_7334,N_6570);
or U8142 (N_8142,N_7009,N_7488);
or U8143 (N_8143,N_6474,N_6203);
nor U8144 (N_8144,N_7639,N_7679);
and U8145 (N_8145,N_7413,N_6427);
or U8146 (N_8146,N_6028,N_6367);
and U8147 (N_8147,N_7296,N_6393);
or U8148 (N_8148,N_7099,N_7588);
xnor U8149 (N_8149,N_6630,N_6313);
and U8150 (N_8150,N_6839,N_6030);
nand U8151 (N_8151,N_6066,N_7672);
or U8152 (N_8152,N_7253,N_7565);
xnor U8153 (N_8153,N_6005,N_6654);
nand U8154 (N_8154,N_7937,N_6444);
and U8155 (N_8155,N_7525,N_6802);
nor U8156 (N_8156,N_7297,N_6855);
nand U8157 (N_8157,N_6804,N_7449);
or U8158 (N_8158,N_6913,N_6605);
xnor U8159 (N_8159,N_6764,N_7735);
xnor U8160 (N_8160,N_6905,N_6984);
or U8161 (N_8161,N_6079,N_7689);
nand U8162 (N_8162,N_7966,N_6274);
nand U8163 (N_8163,N_7266,N_7685);
nand U8164 (N_8164,N_6748,N_7152);
nand U8165 (N_8165,N_6350,N_6298);
or U8166 (N_8166,N_6777,N_7100);
nor U8167 (N_8167,N_6540,N_7800);
xor U8168 (N_8168,N_6782,N_6053);
nand U8169 (N_8169,N_6213,N_7871);
and U8170 (N_8170,N_7339,N_6105);
and U8171 (N_8171,N_7126,N_7499);
xnor U8172 (N_8172,N_7768,N_6089);
xnor U8173 (N_8173,N_7664,N_7802);
nand U8174 (N_8174,N_6558,N_7060);
nor U8175 (N_8175,N_7032,N_6208);
xor U8176 (N_8176,N_7345,N_6435);
xor U8177 (N_8177,N_6489,N_7666);
nor U8178 (N_8178,N_6266,N_7076);
nand U8179 (N_8179,N_7842,N_7897);
and U8180 (N_8180,N_6868,N_6472);
or U8181 (N_8181,N_7720,N_7097);
or U8182 (N_8182,N_7371,N_6744);
nand U8183 (N_8183,N_6807,N_7906);
nor U8184 (N_8184,N_6003,N_6596);
or U8185 (N_8185,N_6417,N_6639);
xnor U8186 (N_8186,N_7132,N_6725);
xnor U8187 (N_8187,N_7343,N_7306);
or U8188 (N_8188,N_7764,N_6439);
nand U8189 (N_8189,N_6430,N_6872);
nor U8190 (N_8190,N_7899,N_7862);
or U8191 (N_8191,N_6339,N_6404);
nor U8192 (N_8192,N_6244,N_6152);
nand U8193 (N_8193,N_7500,N_7581);
or U8194 (N_8194,N_7818,N_7695);
or U8195 (N_8195,N_7091,N_7549);
nand U8196 (N_8196,N_6401,N_6965);
nand U8197 (N_8197,N_7361,N_6320);
nor U8198 (N_8198,N_7898,N_7109);
nand U8199 (N_8199,N_6166,N_7668);
xnor U8200 (N_8200,N_6162,N_7744);
nor U8201 (N_8201,N_6933,N_7377);
xor U8202 (N_8202,N_6165,N_6492);
nand U8203 (N_8203,N_7216,N_6239);
or U8204 (N_8204,N_7105,N_6743);
xnor U8205 (N_8205,N_7325,N_6299);
nand U8206 (N_8206,N_7786,N_6916);
nand U8207 (N_8207,N_6286,N_6841);
xor U8208 (N_8208,N_6086,N_7185);
and U8209 (N_8209,N_7420,N_6794);
or U8210 (N_8210,N_6151,N_7738);
or U8211 (N_8211,N_6963,N_6586);
and U8212 (N_8212,N_7311,N_6116);
nor U8213 (N_8213,N_7623,N_7335);
and U8214 (N_8214,N_7425,N_6383);
nor U8215 (N_8215,N_7246,N_7627);
xnor U8216 (N_8216,N_6834,N_7930);
nand U8217 (N_8217,N_7970,N_7598);
and U8218 (N_8218,N_6433,N_6270);
and U8219 (N_8219,N_7159,N_6778);
xnor U8220 (N_8220,N_7475,N_6641);
and U8221 (N_8221,N_6170,N_6238);
and U8222 (N_8222,N_6985,N_6761);
or U8223 (N_8223,N_7697,N_7175);
or U8224 (N_8224,N_6204,N_7840);
and U8225 (N_8225,N_7520,N_6438);
and U8226 (N_8226,N_6523,N_7085);
or U8227 (N_8227,N_6508,N_7869);
nor U8228 (N_8228,N_7515,N_6359);
and U8229 (N_8229,N_7006,N_7493);
nand U8230 (N_8230,N_6824,N_7675);
nor U8231 (N_8231,N_7626,N_6031);
and U8232 (N_8232,N_6566,N_7797);
and U8233 (N_8233,N_6331,N_7144);
and U8234 (N_8234,N_7380,N_6095);
or U8235 (N_8235,N_7106,N_7992);
or U8236 (N_8236,N_7353,N_6177);
or U8237 (N_8237,N_7208,N_7272);
or U8238 (N_8238,N_6626,N_6880);
or U8239 (N_8239,N_6620,N_6629);
or U8240 (N_8240,N_7130,N_7538);
nand U8241 (N_8241,N_6932,N_7207);
and U8242 (N_8242,N_6867,N_6061);
nand U8243 (N_8243,N_7599,N_7568);
xor U8244 (N_8244,N_7059,N_7674);
or U8245 (N_8245,N_6169,N_7162);
nor U8246 (N_8246,N_6882,N_6554);
nand U8247 (N_8247,N_6898,N_6569);
nand U8248 (N_8248,N_6249,N_6607);
xor U8249 (N_8249,N_7312,N_7771);
or U8250 (N_8250,N_6346,N_6161);
nor U8251 (N_8251,N_7368,N_7198);
nor U8252 (N_8252,N_6256,N_6774);
or U8253 (N_8253,N_7620,N_7021);
xor U8254 (N_8254,N_6966,N_6328);
xnor U8255 (N_8255,N_6495,N_6930);
nand U8256 (N_8256,N_7167,N_6042);
nor U8257 (N_8257,N_6532,N_7112);
or U8258 (N_8258,N_6416,N_6407);
or U8259 (N_8259,N_7236,N_7920);
xor U8260 (N_8260,N_7181,N_7234);
nor U8261 (N_8261,N_6595,N_7502);
nand U8262 (N_8262,N_6715,N_7566);
xor U8263 (N_8263,N_6259,N_6827);
nor U8264 (N_8264,N_7350,N_7682);
xor U8265 (N_8265,N_6016,N_6223);
and U8266 (N_8266,N_6463,N_6603);
nand U8267 (N_8267,N_7383,N_7158);
nand U8268 (N_8268,N_7233,N_6117);
or U8269 (N_8269,N_7924,N_7228);
nor U8270 (N_8270,N_6716,N_6263);
and U8271 (N_8271,N_6732,N_6899);
and U8272 (N_8272,N_6052,N_7120);
or U8273 (N_8273,N_6384,N_6343);
and U8274 (N_8274,N_6976,N_6557);
nand U8275 (N_8275,N_7824,N_7746);
and U8276 (N_8276,N_6608,N_7517);
nand U8277 (N_8277,N_6210,N_6581);
xor U8278 (N_8278,N_7237,N_7737);
nor U8279 (N_8279,N_6440,N_6990);
nand U8280 (N_8280,N_6284,N_6970);
or U8281 (N_8281,N_7260,N_7587);
xnor U8282 (N_8282,N_7979,N_7298);
or U8283 (N_8283,N_6901,N_6881);
or U8284 (N_8284,N_6247,N_7954);
nand U8285 (N_8285,N_6720,N_6437);
nor U8286 (N_8286,N_6364,N_6707);
nand U8287 (N_8287,N_6494,N_6009);
or U8288 (N_8288,N_7153,N_7069);
nor U8289 (N_8289,N_6154,N_7745);
nand U8290 (N_8290,N_7532,N_6600);
nand U8291 (N_8291,N_6625,N_7050);
nor U8292 (N_8292,N_6565,N_7641);
xnor U8293 (N_8293,N_6271,N_7670);
or U8294 (N_8294,N_6964,N_6747);
nand U8295 (N_8295,N_6949,N_6040);
nand U8296 (N_8296,N_7850,N_7631);
nor U8297 (N_8297,N_7055,N_6485);
and U8298 (N_8298,N_6619,N_7584);
nand U8299 (N_8299,N_6168,N_7822);
nor U8300 (N_8300,N_7703,N_6470);
or U8301 (N_8301,N_6296,N_6822);
or U8302 (N_8302,N_7321,N_7295);
or U8303 (N_8303,N_6611,N_7958);
xor U8304 (N_8304,N_7838,N_7694);
xnor U8305 (N_8305,N_6986,N_7145);
nor U8306 (N_8306,N_6661,N_7701);
or U8307 (N_8307,N_6628,N_6892);
nor U8308 (N_8308,N_7516,N_7985);
xor U8309 (N_8309,N_7340,N_7726);
xnor U8310 (N_8310,N_6582,N_7611);
xnor U8311 (N_8311,N_7808,N_7466);
nor U8312 (N_8312,N_7398,N_6451);
or U8313 (N_8313,N_6891,N_6267);
and U8314 (N_8314,N_6937,N_6638);
nand U8315 (N_8315,N_6547,N_6897);
xnor U8316 (N_8316,N_7537,N_6395);
xnor U8317 (N_8317,N_7916,N_7750);
nor U8318 (N_8318,N_6303,N_7774);
nand U8319 (N_8319,N_6043,N_7653);
nand U8320 (N_8320,N_6002,N_6428);
nand U8321 (N_8321,N_6129,N_6689);
nor U8322 (N_8322,N_6805,N_7051);
nor U8323 (N_8323,N_7024,N_7662);
and U8324 (N_8324,N_6385,N_6902);
and U8325 (N_8325,N_7288,N_6787);
xnor U8326 (N_8326,N_6374,N_6524);
and U8327 (N_8327,N_7632,N_6446);
xnor U8328 (N_8328,N_6288,N_6694);
or U8329 (N_8329,N_7606,N_7000);
or U8330 (N_8330,N_7509,N_6146);
xnor U8331 (N_8331,N_6230,N_7438);
or U8332 (N_8332,N_7543,N_7082);
and U8333 (N_8333,N_7835,N_6147);
and U8334 (N_8334,N_6773,N_7683);
xor U8335 (N_8335,N_6135,N_7289);
xnor U8336 (N_8336,N_6858,N_7458);
or U8337 (N_8337,N_6865,N_6571);
nor U8338 (N_8338,N_7829,N_7760);
or U8339 (N_8339,N_6845,N_6712);
nor U8340 (N_8340,N_6559,N_6358);
and U8341 (N_8341,N_6680,N_7089);
nor U8342 (N_8342,N_7950,N_7168);
nand U8343 (N_8343,N_7529,N_7124);
nand U8344 (N_8344,N_7156,N_6413);
xnor U8345 (N_8345,N_6065,N_6091);
and U8346 (N_8346,N_6250,N_6959);
nor U8347 (N_8347,N_7141,N_6321);
nor U8348 (N_8348,N_6150,N_7524);
xnor U8349 (N_8349,N_7941,N_6929);
or U8350 (N_8350,N_7362,N_7595);
nand U8351 (N_8351,N_6248,N_6854);
nand U8352 (N_8352,N_7806,N_6096);
xor U8353 (N_8353,N_7430,N_7429);
nor U8354 (N_8354,N_7795,N_6483);
nor U8355 (N_8355,N_7678,N_7790);
nor U8356 (N_8356,N_6332,N_7482);
xor U8357 (N_8357,N_6033,N_7548);
xnor U8358 (N_8358,N_6125,N_7742);
and U8359 (N_8359,N_7777,N_7990);
or U8360 (N_8360,N_7454,N_6604);
xnor U8361 (N_8361,N_6988,N_7129);
nand U8362 (N_8362,N_7336,N_7716);
or U8363 (N_8363,N_6480,N_6128);
or U8364 (N_8364,N_7074,N_7405);
or U8365 (N_8365,N_7880,N_7017);
nor U8366 (N_8366,N_6429,N_7926);
xnor U8367 (N_8367,N_6634,N_6292);
nor U8368 (N_8368,N_7977,N_7772);
nor U8369 (N_8369,N_6810,N_7866);
or U8370 (N_8370,N_6762,N_6232);
or U8371 (N_8371,N_6665,N_7960);
or U8372 (N_8372,N_7721,N_7229);
xnor U8373 (N_8373,N_7463,N_7594);
nor U8374 (N_8374,N_7218,N_7731);
nand U8375 (N_8375,N_7995,N_7830);
nor U8376 (N_8376,N_6691,N_6767);
and U8377 (N_8377,N_6573,N_6869);
or U8378 (N_8378,N_7905,N_6231);
nand U8379 (N_8379,N_6592,N_6567);
xor U8380 (N_8380,N_6961,N_6316);
or U8381 (N_8381,N_7436,N_6000);
xnor U8382 (N_8382,N_6261,N_7657);
or U8383 (N_8383,N_6873,N_6887);
and U8384 (N_8384,N_7793,N_6758);
or U8385 (N_8385,N_6849,N_6759);
and U8386 (N_8386,N_7477,N_7660);
and U8387 (N_8387,N_6171,N_6391);
xnor U8388 (N_8388,N_7728,N_7913);
or U8389 (N_8389,N_7379,N_7367);
nand U8390 (N_8390,N_6379,N_7359);
or U8391 (N_8391,N_7951,N_7111);
or U8392 (N_8392,N_6160,N_6545);
and U8393 (N_8393,N_6115,N_7554);
xnor U8394 (N_8394,N_7717,N_6903);
and U8395 (N_8395,N_7562,N_7471);
xor U8396 (N_8396,N_6196,N_7681);
or U8397 (N_8397,N_6852,N_7552);
nor U8398 (N_8398,N_6888,N_7508);
or U8399 (N_8399,N_7376,N_7604);
nor U8400 (N_8400,N_6104,N_6083);
and U8401 (N_8401,N_7204,N_7778);
xor U8402 (N_8402,N_7615,N_6594);
or U8403 (N_8403,N_7256,N_6575);
xor U8404 (N_8404,N_7848,N_6245);
or U8405 (N_8405,N_6519,N_6830);
or U8406 (N_8406,N_7123,N_7058);
and U8407 (N_8407,N_6458,N_7586);
and U8408 (N_8408,N_7570,N_6035);
xnor U8409 (N_8409,N_6134,N_6473);
nand U8410 (N_8410,N_6553,N_6155);
xor U8411 (N_8411,N_7736,N_6653);
nor U8412 (N_8412,N_6589,N_7358);
and U8413 (N_8413,N_7462,N_6560);
or U8414 (N_8414,N_7012,N_6836);
nor U8415 (N_8415,N_6111,N_6038);
xnor U8416 (N_8416,N_7195,N_7476);
nor U8417 (N_8417,N_7577,N_6572);
nand U8418 (N_8418,N_6578,N_6615);
and U8419 (N_8419,N_7722,N_6193);
xnor U8420 (N_8420,N_7320,N_7887);
or U8421 (N_8421,N_7860,N_7747);
xor U8422 (N_8422,N_6857,N_7270);
xnor U8423 (N_8423,N_6551,N_7618);
or U8424 (N_8424,N_7490,N_7197);
nor U8425 (N_8425,N_7580,N_7384);
xnor U8426 (N_8426,N_6914,N_7174);
nand U8427 (N_8427,N_6176,N_6693);
or U8428 (N_8428,N_6798,N_7705);
nand U8429 (N_8429,N_7912,N_6698);
nor U8430 (N_8430,N_7884,N_6342);
or U8431 (N_8431,N_6370,N_6769);
nor U8432 (N_8432,N_7274,N_6217);
nor U8433 (N_8433,N_6056,N_6499);
nor U8434 (N_8434,N_6484,N_6454);
nand U8435 (N_8435,N_6987,N_7421);
nand U8436 (N_8436,N_6846,N_6106);
nor U8437 (N_8437,N_7434,N_6812);
or U8438 (N_8438,N_7448,N_7784);
nand U8439 (N_8439,N_7108,N_7090);
or U8440 (N_8440,N_6801,N_7375);
or U8441 (N_8441,N_6189,N_7319);
nor U8442 (N_8442,N_6246,N_6039);
xor U8443 (N_8443,N_6940,N_7310);
or U8444 (N_8444,N_6225,N_7530);
or U8445 (N_8445,N_6876,N_6110);
xor U8446 (N_8446,N_7364,N_7318);
and U8447 (N_8447,N_7285,N_7942);
nor U8448 (N_8448,N_6831,N_6666);
and U8449 (N_8449,N_6327,N_6746);
and U8450 (N_8450,N_7903,N_7008);
and U8451 (N_8451,N_6293,N_6612);
or U8452 (N_8452,N_7492,N_6365);
or U8453 (N_8453,N_6669,N_7944);
xnor U8454 (N_8454,N_7299,N_6510);
xor U8455 (N_8455,N_7019,N_6516);
nand U8456 (N_8456,N_6696,N_7267);
nand U8457 (N_8457,N_7724,N_7396);
and U8458 (N_8458,N_6924,N_7065);
nand U8459 (N_8459,N_6449,N_7314);
nor U8460 (N_8460,N_6944,N_7007);
or U8461 (N_8461,N_6706,N_7667);
nand U8462 (N_8462,N_7545,N_7630);
nand U8463 (N_8463,N_6148,N_7064);
or U8464 (N_8464,N_6060,N_7895);
nor U8465 (N_8465,N_7470,N_7355);
nor U8466 (N_8466,N_6120,N_6817);
nor U8467 (N_8467,N_6711,N_7182);
nand U8468 (N_8468,N_6700,N_6182);
xor U8469 (N_8469,N_7972,N_6445);
nand U8470 (N_8470,N_7794,N_6262);
nor U8471 (N_8471,N_7644,N_6141);
or U8472 (N_8472,N_7304,N_7349);
nand U8473 (N_8473,N_7823,N_6953);
and U8474 (N_8474,N_7113,N_7227);
or U8475 (N_8475,N_6398,N_6992);
nor U8476 (N_8476,N_7029,N_7150);
nor U8477 (N_8477,N_6084,N_7249);
and U8478 (N_8478,N_7699,N_7183);
nor U8479 (N_8479,N_6969,N_6420);
or U8480 (N_8480,N_7360,N_6396);
and U8481 (N_8481,N_6536,N_6102);
nand U8482 (N_8482,N_6948,N_6878);
xnor U8483 (N_8483,N_7597,N_7190);
nand U8484 (N_8484,N_6077,N_7373);
nand U8485 (N_8485,N_6504,N_6318);
xnor U8486 (N_8486,N_7184,N_6909);
nand U8487 (N_8487,N_6667,N_6555);
and U8488 (N_8488,N_6563,N_6598);
or U8489 (N_8489,N_6112,N_7214);
nand U8490 (N_8490,N_7390,N_6294);
xor U8491 (N_8491,N_7070,N_6425);
or U8492 (N_8492,N_7663,N_7607);
nor U8493 (N_8493,N_6497,N_7282);
or U8494 (N_8494,N_6048,N_7550);
xnor U8495 (N_8495,N_6904,N_6082);
xor U8496 (N_8496,N_7754,N_6087);
and U8497 (N_8497,N_6044,N_7486);
and U8498 (N_8498,N_6478,N_6025);
and U8499 (N_8499,N_7447,N_6789);
and U8500 (N_8500,N_6465,N_7798);
or U8501 (N_8501,N_7428,N_7613);
nor U8502 (N_8502,N_6766,N_7837);
nor U8503 (N_8503,N_7868,N_6402);
nor U8504 (N_8504,N_7199,N_6414);
nand U8505 (N_8505,N_6745,N_7407);
nor U8506 (N_8506,N_7054,N_6527);
nor U8507 (N_8507,N_7982,N_7629);
xor U8508 (N_8508,N_6525,N_6705);
xor U8509 (N_8509,N_6912,N_7056);
xor U8510 (N_8510,N_7879,N_6265);
and U8511 (N_8511,N_7622,N_7560);
and U8512 (N_8512,N_7507,N_7836);
xor U8513 (N_8513,N_6894,N_7134);
and U8514 (N_8514,N_6277,N_7276);
nand U8515 (N_8515,N_7337,N_6950);
or U8516 (N_8516,N_7072,N_6386);
or U8517 (N_8517,N_7503,N_7268);
and U8518 (N_8518,N_7275,N_6215);
xor U8519 (N_8519,N_7856,N_7404);
nand U8520 (N_8520,N_6844,N_7157);
or U8521 (N_8521,N_6808,N_6682);
and U8522 (N_8522,N_6550,N_7400);
xnor U8523 (N_8523,N_6421,N_7637);
nand U8524 (N_8524,N_6149,N_7250);
xnor U8525 (N_8525,N_7453,N_7933);
and U8526 (N_8526,N_7762,N_6792);
xnor U8527 (N_8527,N_7242,N_7984);
and U8528 (N_8528,N_6734,N_6617);
nor U8529 (N_8529,N_7461,N_6014);
or U8530 (N_8530,N_7049,N_6300);
xnor U8531 (N_8531,N_6185,N_6647);
and U8532 (N_8532,N_7243,N_7593);
or U8533 (N_8533,N_6677,N_7442);
and U8534 (N_8534,N_7437,N_6295);
or U8535 (N_8535,N_6776,N_6864);
or U8536 (N_8536,N_7044,N_6178);
nor U8537 (N_8537,N_6818,N_7980);
nand U8538 (N_8538,N_6991,N_7062);
nand U8539 (N_8539,N_7527,N_7743);
nand U8540 (N_8540,N_7435,N_7381);
or U8541 (N_8541,N_6080,N_7773);
nand U8542 (N_8542,N_6431,N_6585);
and U8543 (N_8543,N_7872,N_7761);
nand U8544 (N_8544,N_7707,N_6190);
nand U8545 (N_8545,N_7709,N_7300);
nor U8546 (N_8546,N_6278,N_7544);
nor U8547 (N_8547,N_6415,N_6996);
nor U8548 (N_8548,N_6408,N_6090);
nand U8549 (N_8549,N_7700,N_7635);
and U8550 (N_8550,N_7338,N_7659);
xnor U8551 (N_8551,N_6064,N_7891);
and U8552 (N_8552,N_6004,N_6198);
and U8553 (N_8553,N_6621,N_6967);
nor U8554 (N_8554,N_7874,N_6399);
nand U8555 (N_8555,N_7263,N_7315);
nor U8556 (N_8556,N_7927,N_6601);
nor U8557 (N_8557,N_7934,N_7025);
and U8558 (N_8558,N_6032,N_7557);
nor U8559 (N_8559,N_7302,N_7426);
and U8560 (N_8560,N_7770,N_7016);
or U8561 (N_8561,N_7753,N_7220);
or U8562 (N_8562,N_7997,N_6850);
nand U8563 (N_8563,N_6229,N_7231);
xor U8564 (N_8564,N_6179,N_7741);
nor U8565 (N_8565,N_7402,N_6772);
nor U8566 (N_8566,N_6008,N_7305);
nand U8567 (N_8567,N_6515,N_7739);
or U8568 (N_8568,N_7235,N_7226);
nor U8569 (N_8569,N_6145,N_6243);
and U8570 (N_8570,N_6692,N_6279);
nor U8571 (N_8571,N_7931,N_7291);
xnor U8572 (N_8572,N_7759,N_7443);
nor U8573 (N_8573,N_6192,N_7536);
nor U8574 (N_8574,N_6649,N_6180);
nor U8575 (N_8575,N_7834,N_6368);
xor U8576 (N_8576,N_7086,N_6741);
or U8577 (N_8577,N_6434,N_7172);
and U8578 (N_8578,N_7102,N_6907);
nor U8579 (N_8579,N_6452,N_6955);
nor U8580 (N_8580,N_6995,N_6678);
xor U8581 (N_8581,N_7628,N_7600);
and U8582 (N_8582,N_7885,N_7392);
nand U8583 (N_8583,N_6651,N_6491);
or U8584 (N_8584,N_6859,N_6254);
and U8585 (N_8585,N_7787,N_7147);
nand U8586 (N_8586,N_6455,N_7316);
nor U8587 (N_8587,N_6037,N_6049);
xor U8588 (N_8588,N_6624,N_6409);
nor U8589 (N_8589,N_6482,N_6159);
and U8590 (N_8590,N_7658,N_6506);
and U8591 (N_8591,N_6919,N_7649);
nand U8592 (N_8592,N_6528,N_6784);
nand U8593 (N_8593,N_6538,N_6685);
and U8594 (N_8594,N_6153,N_6139);
xnor U8595 (N_8595,N_7053,N_6453);
nor U8596 (N_8596,N_6207,N_7087);
nor U8597 (N_8597,N_7978,N_7922);
nand U8598 (N_8598,N_6579,N_6462);
and U8599 (N_8599,N_6101,N_7422);
or U8600 (N_8600,N_6908,N_7357);
xor U8601 (N_8601,N_7945,N_7444);
nand U8602 (N_8602,N_6467,N_6347);
xnor U8603 (N_8603,N_6432,N_7965);
nand U8604 (N_8604,N_6754,N_7080);
and U8605 (N_8605,N_6737,N_6228);
and U8606 (N_8606,N_6157,N_6012);
or U8607 (N_8607,N_6797,N_6768);
and U8608 (N_8608,N_6939,N_6548);
xor U8609 (N_8609,N_7484,N_6394);
and U8610 (N_8610,N_7052,N_7648);
or U8611 (N_8611,N_6825,N_6771);
xnor U8612 (N_8612,N_6330,N_6780);
and U8613 (N_8613,N_6915,N_7139);
and U8614 (N_8614,N_6840,N_7177);
nor U8615 (N_8615,N_6418,N_6522);
or U8616 (N_8616,N_7996,N_6436);
nor U8617 (N_8617,N_6925,N_7031);
xnor U8618 (N_8618,N_6175,N_6640);
nand U8619 (N_8619,N_6670,N_7039);
or U8620 (N_8620,N_6227,N_7232);
nor U8621 (N_8621,N_6119,N_6172);
xnor U8622 (N_8622,N_7833,N_6529);
nor U8623 (N_8623,N_6051,N_6828);
or U8624 (N_8624,N_6376,N_6059);
nor U8625 (N_8625,N_7710,N_7534);
or U8626 (N_8626,N_6055,N_7643);
nor U8627 (N_8627,N_7821,N_6871);
or U8628 (N_8628,N_7075,N_6686);
or U8629 (N_8629,N_7191,N_7576);
and U8630 (N_8630,N_7952,N_6158);
or U8631 (N_8631,N_7751,N_6097);
xor U8632 (N_8632,N_7326,N_7491);
or U8633 (N_8633,N_7424,N_6549);
nand U8634 (N_8634,N_6026,N_6017);
nor U8635 (N_8635,N_7963,N_7445);
nand U8636 (N_8636,N_7494,N_6071);
and U8637 (N_8637,N_7702,N_7212);
or U8638 (N_8638,N_7457,N_7910);
nor U8639 (N_8639,N_7749,N_7765);
or U8640 (N_8640,N_7081,N_6765);
or U8641 (N_8641,N_7939,N_7752);
nor U8642 (N_8642,N_7713,N_6081);
xor U8643 (N_8643,N_7691,N_6340);
and U8644 (N_8644,N_7864,N_7579);
nand U8645 (N_8645,N_6613,N_7037);
nor U8646 (N_8646,N_6835,N_6574);
nor U8647 (N_8647,N_6488,N_7510);
xnor U8648 (N_8648,N_7347,N_6069);
xor U8649 (N_8649,N_6099,N_6974);
nor U8650 (N_8650,N_7501,N_7789);
nand U8651 (N_8651,N_7504,N_6718);
xnor U8652 (N_8652,N_7063,N_7928);
nor U8653 (N_8653,N_7867,N_6663);
nor U8654 (N_8654,N_7655,N_6094);
xnor U8655 (N_8655,N_6752,N_6443);
or U8656 (N_8656,N_6273,N_7327);
and U8657 (N_8657,N_7521,N_6922);
and U8658 (N_8658,N_7328,N_6251);
nand U8659 (N_8659,N_6188,N_6410);
nand U8660 (N_8660,N_7756,N_6297);
nor U8661 (N_8661,N_7914,N_7935);
and U8662 (N_8662,N_7647,N_7999);
nand U8663 (N_8663,N_7446,N_6520);
nor U8664 (N_8664,N_7131,N_7766);
nor U8665 (N_8665,N_6820,N_7388);
and U8666 (N_8666,N_6733,N_7748);
xnor U8667 (N_8667,N_7255,N_7035);
nand U8668 (N_8668,N_6220,N_7209);
xnor U8669 (N_8669,N_7656,N_7088);
xnor U8670 (N_8670,N_7998,N_6972);
nor U8671 (N_8671,N_6282,N_7114);
nor U8672 (N_8672,N_6517,N_6833);
xor U8673 (N_8673,N_6701,N_7955);
nor U8674 (N_8674,N_6866,N_7692);
xnor U8675 (N_8675,N_6623,N_7192);
or U8676 (N_8676,N_6756,N_6450);
nand U8677 (N_8677,N_6045,N_7292);
xnor U8678 (N_8678,N_7610,N_7563);
or U8679 (N_8679,N_7151,N_6073);
or U8680 (N_8680,N_7878,N_7222);
and U8681 (N_8681,N_6397,N_7704);
and U8682 (N_8682,N_7578,N_6688);
and U8683 (N_8683,N_7902,N_7719);
nand U8684 (N_8684,N_6534,N_7416);
and U8685 (N_8685,N_7040,N_7200);
or U8686 (N_8686,N_7450,N_7254);
nand U8687 (N_8687,N_7414,N_6813);
xor U8688 (N_8688,N_7669,N_7981);
or U8689 (N_8689,N_7791,N_7309);
nand U8690 (N_8690,N_6597,N_6973);
and U8691 (N_8691,N_7341,N_7067);
nand U8692 (N_8692,N_7561,N_6664);
nor U8693 (N_8693,N_7876,N_7188);
nand U8694 (N_8694,N_7103,N_7946);
nand U8695 (N_8695,N_6757,N_6338);
nor U8696 (N_8696,N_7078,N_7286);
nor U8697 (N_8697,N_7022,N_7077);
nand U8698 (N_8698,N_7205,N_7351);
and U8699 (N_8699,N_7852,N_6655);
nand U8700 (N_8700,N_6326,N_6552);
nor U8701 (N_8701,N_6366,N_6018);
and U8702 (N_8702,N_7410,N_6576);
nand U8703 (N_8703,N_6311,N_6543);
xor U8704 (N_8704,N_7911,N_6874);
xnor U8705 (N_8705,N_7583,N_7858);
nand U8706 (N_8706,N_6542,N_7121);
or U8707 (N_8707,N_6133,N_7117);
or U8708 (N_8708,N_6375,N_7889);
and U8709 (N_8709,N_7792,N_6790);
or U8710 (N_8710,N_6468,N_6469);
nand U8711 (N_8711,N_7495,N_6740);
xnor U8712 (N_8712,N_6531,N_6205);
nor U8713 (N_8713,N_7556,N_7455);
nor U8714 (N_8714,N_6107,N_7452);
nor U8715 (N_8715,N_6978,N_7474);
or U8716 (N_8716,N_7863,N_6212);
nand U8717 (N_8717,N_6683,N_6673);
nand U8718 (N_8718,N_6635,N_7690);
or U8719 (N_8719,N_7564,N_7143);
xor U8720 (N_8720,N_7284,N_6606);
nand U8721 (N_8721,N_7859,N_6648);
nand U8722 (N_8722,N_6631,N_7073);
nand U8723 (N_8723,N_7696,N_7005);
xnor U8724 (N_8724,N_7252,N_6424);
nor U8725 (N_8725,N_6695,N_7553);
and U8726 (N_8726,N_6561,N_6507);
and U8727 (N_8727,N_7210,N_7892);
xnor U8728 (N_8728,N_7609,N_7890);
and U8729 (N_8729,N_6187,N_6308);
nand U8730 (N_8730,N_7301,N_6609);
xor U8731 (N_8731,N_6602,N_6264);
and U8732 (N_8732,N_7855,N_7411);
and U8733 (N_8733,N_7665,N_7541);
nor U8734 (N_8734,N_7573,N_6068);
and U8735 (N_8735,N_7169,N_7038);
nand U8736 (N_8736,N_7511,N_6660);
xor U8737 (N_8737,N_6377,N_7801);
or U8738 (N_8738,N_7732,N_6108);
or U8739 (N_8739,N_6337,N_6315);
xnor U8740 (N_8740,N_6194,N_7559);
or U8741 (N_8741,N_7714,N_6943);
or U8742 (N_8742,N_6240,N_7514);
nor U8743 (N_8743,N_6403,N_7196);
or U8744 (N_8744,N_6382,N_6290);
or U8745 (N_8745,N_6722,N_6336);
xor U8746 (N_8746,N_6487,N_6199);
and U8747 (N_8747,N_7166,N_6799);
or U8748 (N_8748,N_7465,N_6144);
nor U8749 (N_8749,N_6945,N_6975);
xnor U8750 (N_8750,N_7322,N_6257);
and U8751 (N_8751,N_6124,N_6717);
nor U8752 (N_8752,N_7727,N_6793);
nand U8753 (N_8753,N_7473,N_7202);
nand U8754 (N_8754,N_6796,N_6252);
or U8755 (N_8755,N_7225,N_7026);
xnor U8756 (N_8756,N_7346,N_7755);
and U8757 (N_8757,N_6942,N_7590);
nand U8758 (N_8758,N_6826,N_7483);
and U8759 (N_8759,N_7820,N_6348);
nand U8760 (N_8760,N_7723,N_6509);
nand U8761 (N_8761,N_6610,N_6481);
xnor U8762 (N_8762,N_6007,N_7923);
and U8763 (N_8763,N_7844,N_7591);
nand U8764 (N_8764,N_7083,N_7883);
nor U8765 (N_8765,N_7382,N_6614);
xnor U8766 (N_8766,N_7331,N_6788);
and U8767 (N_8767,N_6118,N_6645);
and U8768 (N_8768,N_7909,N_7395);
nand U8769 (N_8769,N_6362,N_6241);
xor U8770 (N_8770,N_6200,N_6751);
nand U8771 (N_8771,N_6388,N_6291);
or U8772 (N_8772,N_6936,N_7294);
nand U8773 (N_8773,N_7176,N_7155);
and U8774 (N_8774,N_7273,N_7329);
and U8775 (N_8775,N_7847,N_7929);
nand U8776 (N_8776,N_6255,N_7165);
and U8777 (N_8777,N_7014,N_7092);
or U8778 (N_8778,N_7810,N_6490);
or U8779 (N_8779,N_7066,N_7140);
nor U8780 (N_8780,N_7651,N_7027);
nor U8781 (N_8781,N_6305,N_6637);
or U8782 (N_8782,N_6526,N_7146);
nand U8783 (N_8783,N_6591,N_6074);
or U8784 (N_8784,N_7730,N_7264);
nand U8785 (N_8785,N_6272,N_6195);
xnor U8786 (N_8786,N_7441,N_6142);
xor U8787 (N_8787,N_7558,N_6381);
and U8788 (N_8788,N_6067,N_6088);
nor U8789 (N_8789,N_6503,N_7614);
and U8790 (N_8790,N_6726,N_6411);
or U8791 (N_8791,N_6143,N_7767);
nor U8792 (N_8792,N_6356,N_6283);
or U8793 (N_8793,N_6714,N_6981);
xnor U8794 (N_8794,N_6191,N_6900);
nand U8795 (N_8795,N_7240,N_6276);
xor U8796 (N_8796,N_6809,N_7366);
nor U8797 (N_8797,N_7506,N_6457);
or U8798 (N_8798,N_7846,N_7406);
and U8799 (N_8799,N_7440,N_6781);
or U8800 (N_8800,N_7919,N_7068);
or U8801 (N_8801,N_7904,N_7213);
and U8802 (N_8802,N_7986,N_6334);
xnor U8803 (N_8803,N_7733,N_6380);
xor U8804 (N_8804,N_6918,N_7582);
or U8805 (N_8805,N_6029,N_6312);
and U8806 (N_8806,N_6513,N_7460);
or U8807 (N_8807,N_6895,N_7118);
nand U8808 (N_8808,N_6672,N_7947);
nand U8809 (N_8809,N_6075,N_6021);
xor U8810 (N_8810,N_6057,N_7271);
xor U8811 (N_8811,N_7932,N_6174);
xor U8812 (N_8812,N_7854,N_6539);
nand U8813 (N_8813,N_6070,N_6353);
nand U8814 (N_8814,N_7278,N_7142);
nor U8815 (N_8815,N_7342,N_6763);
nor U8816 (N_8816,N_6302,N_7988);
or U8817 (N_8817,N_6911,N_6214);
and U8818 (N_8818,N_6713,N_7953);
and U8819 (N_8819,N_6627,N_7427);
or U8820 (N_8820,N_7011,N_6738);
and U8821 (N_8821,N_7706,N_7661);
or U8822 (N_8822,N_7522,N_6851);
or U8823 (N_8823,N_7317,N_6811);
or U8824 (N_8824,N_7251,N_6521);
and U8825 (N_8825,N_6979,N_6138);
or U8826 (N_8826,N_7815,N_7203);
xor U8827 (N_8827,N_6047,N_6173);
or U8828 (N_8828,N_7687,N_6679);
nand U8829 (N_8829,N_6275,N_6643);
and U8830 (N_8830,N_7186,N_7915);
nand U8831 (N_8831,N_7814,N_7540);
nand U8832 (N_8832,N_6556,N_6946);
or U8833 (N_8833,N_7061,N_7018);
nor U8834 (N_8834,N_6709,N_7432);
xor U8835 (N_8835,N_6186,N_7546);
or U8836 (N_8836,N_6530,N_6046);
or U8837 (N_8837,N_7969,N_6889);
and U8838 (N_8838,N_7729,N_7344);
nand U8839 (N_8839,N_6999,N_6587);
nand U8840 (N_8840,N_6253,N_6324);
nand U8841 (N_8841,N_6132,N_7803);
nor U8842 (N_8842,N_6853,N_6622);
nor U8843 (N_8843,N_6093,N_7596);
xnor U8844 (N_8844,N_6325,N_6387);
or U8845 (N_8845,N_7385,N_6593);
and U8846 (N_8846,N_7603,N_6893);
nand U8847 (N_8847,N_6657,N_7399);
nand U8848 (N_8848,N_7201,N_6258);
nand U8849 (N_8849,N_7831,N_6906);
or U8850 (N_8850,N_6847,N_7989);
nor U8851 (N_8851,N_7034,N_7451);
xor U8852 (N_8852,N_7827,N_6721);
nor U8853 (N_8853,N_7046,N_7956);
or U8854 (N_8854,N_6349,N_6977);
or U8855 (N_8855,N_6486,N_6041);
or U8856 (N_8856,N_6235,N_6533);
or U8857 (N_8857,N_6167,N_6406);
nand U8858 (N_8858,N_6968,N_7370);
and U8859 (N_8859,N_7259,N_6022);
nand U8860 (N_8860,N_7194,N_7718);
or U8861 (N_8861,N_6931,N_7036);
nor U8862 (N_8862,N_7817,N_6389);
nor U8863 (N_8863,N_7048,N_7178);
xor U8864 (N_8864,N_6636,N_7217);
nor U8865 (N_8865,N_7332,N_6181);
or U8866 (N_8866,N_7478,N_7261);
or U8867 (N_8867,N_7569,N_7975);
nor U8868 (N_8868,N_7612,N_6783);
or U8869 (N_8869,N_7480,N_6268);
and U8870 (N_8870,N_7417,N_7020);
xnor U8871 (N_8871,N_6687,N_6819);
nor U8872 (N_8872,N_6795,N_6676);
nand U8873 (N_8873,N_6511,N_6306);
or U8874 (N_8874,N_7519,N_6109);
nand U8875 (N_8875,N_7757,N_7804);
and U8876 (N_8876,N_6355,N_7028);
or U8877 (N_8877,N_7624,N_6285);
or U8878 (N_8878,N_7497,N_6588);
nor U8879 (N_8879,N_7223,N_7287);
and U8880 (N_8880,N_6426,N_7921);
nor U8881 (N_8881,N_6209,N_6222);
nand U8882 (N_8882,N_7378,N_7873);
nand U8883 (N_8883,N_7119,N_6226);
nor U8884 (N_8884,N_7547,N_6890);
nand U8885 (N_8885,N_7959,N_7389);
nor U8886 (N_8886,N_6514,N_6201);
and U8887 (N_8887,N_6063,N_7725);
nor U8888 (N_8888,N_6050,N_7652);
xnor U8889 (N_8889,N_6419,N_7496);
and U8890 (N_8890,N_7363,N_7397);
xor U8891 (N_8891,N_7640,N_7433);
xnor U8892 (N_8892,N_7003,N_6136);
xor U8893 (N_8893,N_7634,N_6400);
nor U8894 (N_8894,N_6335,N_6883);
nand U8895 (N_8895,N_6935,N_7968);
and U8896 (N_8896,N_6493,N_7431);
nand U8897 (N_8897,N_7002,N_6956);
and U8898 (N_8898,N_6642,N_7832);
nand U8899 (N_8899,N_7907,N_7277);
nand U8900 (N_8900,N_6998,N_6838);
nand U8901 (N_8901,N_7853,N_6770);
nor U8902 (N_8902,N_6577,N_7693);
nor U8903 (N_8903,N_7189,N_6512);
nand U8904 (N_8904,N_6736,N_6098);
nor U8905 (N_8905,N_7851,N_7487);
or U8906 (N_8906,N_7394,N_6710);
and U8907 (N_8907,N_6156,N_7171);
xor U8908 (N_8908,N_6314,N_6023);
xor U8909 (N_8909,N_6020,N_7888);
nor U8910 (N_8910,N_6760,N_6652);
nor U8911 (N_8911,N_6280,N_6216);
nand U8912 (N_8912,N_6928,N_7813);
nor U8913 (N_8913,N_7127,N_6719);
nor U8914 (N_8914,N_6344,N_7788);
xor U8915 (N_8915,N_6019,N_7526);
xnor U8916 (N_8916,N_6735,N_7281);
and U8917 (N_8917,N_7843,N_6479);
nor U8918 (N_8918,N_6583,N_6369);
nor U8919 (N_8919,N_6301,N_6078);
xnor U8920 (N_8920,N_7518,N_7456);
nor U8921 (N_8921,N_7280,N_7779);
nor U8922 (N_8922,N_7303,N_7642);
nand U8923 (N_8923,N_7865,N_6633);
nor U8924 (N_8924,N_6564,N_6072);
nor U8925 (N_8925,N_7875,N_6862);
nor U8926 (N_8926,N_7408,N_7839);
or U8927 (N_8927,N_6015,N_6392);
nand U8928 (N_8928,N_6361,N_6674);
and U8929 (N_8929,N_7136,N_6644);
nand U8930 (N_8930,N_6234,N_7323);
or U8931 (N_8931,N_7542,N_7602);
or U8932 (N_8932,N_7096,N_7230);
nor U8933 (N_8933,N_6496,N_6363);
nor U8934 (N_8934,N_6114,N_7057);
nor U8935 (N_8935,N_7812,N_6036);
nand U8936 (N_8936,N_6681,N_6749);
or U8937 (N_8937,N_6405,N_6923);
nand U8938 (N_8938,N_7533,N_7485);
or U8939 (N_8939,N_7625,N_6884);
or U8940 (N_8940,N_7974,N_7799);
nand U8941 (N_8941,N_6164,N_6568);
xnor U8942 (N_8942,N_6184,N_6837);
nand U8943 (N_8943,N_7138,N_6896);
nand U8944 (N_8944,N_6863,N_6137);
and U8945 (N_8945,N_7551,N_6753);
nor U8946 (N_8946,N_7333,N_7712);
and U8947 (N_8947,N_7403,N_6728);
and U8948 (N_8948,N_7973,N_6354);
xnor U8949 (N_8949,N_7734,N_7133);
nor U8950 (N_8950,N_6656,N_6997);
or U8951 (N_8951,N_7354,N_7782);
nor U8952 (N_8952,N_6938,N_7084);
or U8953 (N_8953,N_7107,N_7247);
xor U8954 (N_8954,N_7619,N_7224);
xnor U8955 (N_8955,N_7356,N_6994);
xor U8956 (N_8956,N_7646,N_7467);
nand U8957 (N_8957,N_6498,N_6727);
xnor U8958 (N_8958,N_6684,N_7783);
or U8959 (N_8959,N_7489,N_6211);
xnor U8960 (N_8960,N_6219,N_7555);
or U8961 (N_8961,N_6441,N_7512);
and U8962 (N_8962,N_7908,N_7763);
nand U8963 (N_8963,N_6646,N_6100);
and U8964 (N_8964,N_7170,N_7238);
or U8965 (N_8965,N_7137,N_6877);
nor U8966 (N_8966,N_7886,N_7893);
nand U8967 (N_8967,N_7638,N_7572);
xnor U8968 (N_8968,N_7967,N_7244);
nand U8969 (N_8969,N_7257,N_7479);
nor U8970 (N_8970,N_6477,N_7571);
xnor U8971 (N_8971,N_7994,N_7116);
xor U8972 (N_8972,N_6103,N_6461);
xor U8973 (N_8973,N_7940,N_7283);
xor U8974 (N_8974,N_6982,N_7957);
nand U8975 (N_8975,N_6584,N_6287);
nor U8976 (N_8976,N_6786,N_7412);
nor U8977 (N_8977,N_6237,N_6501);
or U8978 (N_8978,N_6422,N_7401);
xor U8979 (N_8979,N_7372,N_6755);
xnor U8980 (N_8980,N_7769,N_7071);
and U8981 (N_8981,N_7239,N_7258);
nor U8982 (N_8982,N_7828,N_7094);
xor U8983 (N_8983,N_7043,N_7592);
and U8984 (N_8984,N_7807,N_7535);
and U8985 (N_8985,N_6742,N_6958);
nor U8986 (N_8986,N_6034,N_7193);
xor U8987 (N_8987,N_6309,N_7030);
xnor U8988 (N_8988,N_6221,N_6001);
and U8989 (N_8989,N_6054,N_7004);
nand U8990 (N_8990,N_6518,N_6423);
and U8991 (N_8991,N_6197,N_6322);
and U8992 (N_8992,N_7961,N_7173);
and U8993 (N_8993,N_6122,N_6960);
nand U8994 (N_8994,N_6236,N_7811);
xor U8995 (N_8995,N_6390,N_7816);
xor U8996 (N_8996,N_6927,N_7307);
nand U8997 (N_8997,N_6739,N_6281);
xnor U8998 (N_8998,N_6010,N_7983);
nor U8999 (N_8999,N_6951,N_7219);
xnor U9000 (N_9000,N_6782,N_6608);
and U9001 (N_9001,N_7258,N_6090);
or U9002 (N_9002,N_6038,N_6030);
nand U9003 (N_9003,N_7872,N_7828);
nand U9004 (N_9004,N_7873,N_7145);
and U9005 (N_9005,N_7368,N_7719);
nor U9006 (N_9006,N_6320,N_6232);
xnor U9007 (N_9007,N_6656,N_6838);
or U9008 (N_9008,N_6992,N_6118);
xnor U9009 (N_9009,N_7042,N_7738);
xor U9010 (N_9010,N_7726,N_7617);
and U9011 (N_9011,N_7221,N_6426);
or U9012 (N_9012,N_7601,N_7506);
xor U9013 (N_9013,N_7362,N_7578);
nand U9014 (N_9014,N_6306,N_7923);
and U9015 (N_9015,N_6446,N_7110);
nor U9016 (N_9016,N_7858,N_7193);
xnor U9017 (N_9017,N_6100,N_7740);
nand U9018 (N_9018,N_7098,N_7518);
or U9019 (N_9019,N_6134,N_7997);
nand U9020 (N_9020,N_7115,N_6259);
nor U9021 (N_9021,N_7540,N_6233);
nand U9022 (N_9022,N_6092,N_6278);
xnor U9023 (N_9023,N_7296,N_6146);
and U9024 (N_9024,N_6595,N_6178);
nand U9025 (N_9025,N_6574,N_7210);
nor U9026 (N_9026,N_7642,N_7749);
xor U9027 (N_9027,N_7025,N_6695);
nand U9028 (N_9028,N_7297,N_6199);
nor U9029 (N_9029,N_7224,N_7869);
or U9030 (N_9030,N_6529,N_6537);
xor U9031 (N_9031,N_6305,N_6369);
xor U9032 (N_9032,N_7410,N_7271);
and U9033 (N_9033,N_6713,N_6681);
and U9034 (N_9034,N_7077,N_7631);
xnor U9035 (N_9035,N_6543,N_6205);
nand U9036 (N_9036,N_6780,N_6210);
nor U9037 (N_9037,N_6059,N_6714);
and U9038 (N_9038,N_6291,N_6375);
and U9039 (N_9039,N_7760,N_7088);
nand U9040 (N_9040,N_7957,N_7405);
or U9041 (N_9041,N_6466,N_7749);
nand U9042 (N_9042,N_6188,N_7563);
nand U9043 (N_9043,N_7918,N_7226);
nor U9044 (N_9044,N_6904,N_6159);
or U9045 (N_9045,N_7787,N_6428);
nand U9046 (N_9046,N_7024,N_7084);
and U9047 (N_9047,N_7729,N_6539);
nor U9048 (N_9048,N_7490,N_7324);
and U9049 (N_9049,N_6176,N_6430);
nand U9050 (N_9050,N_7334,N_6232);
and U9051 (N_9051,N_7460,N_6869);
and U9052 (N_9052,N_6157,N_7498);
and U9053 (N_9053,N_7872,N_7173);
nor U9054 (N_9054,N_6195,N_6403);
xor U9055 (N_9055,N_6748,N_7342);
or U9056 (N_9056,N_6332,N_7980);
nor U9057 (N_9057,N_6358,N_7602);
xor U9058 (N_9058,N_6982,N_7546);
nand U9059 (N_9059,N_7483,N_7074);
or U9060 (N_9060,N_6551,N_6237);
and U9061 (N_9061,N_6350,N_7042);
or U9062 (N_9062,N_7538,N_6806);
or U9063 (N_9063,N_7846,N_7446);
or U9064 (N_9064,N_6417,N_7740);
nand U9065 (N_9065,N_6708,N_7583);
nand U9066 (N_9066,N_6041,N_6485);
or U9067 (N_9067,N_7947,N_7418);
and U9068 (N_9068,N_7425,N_6583);
nand U9069 (N_9069,N_7714,N_6793);
xor U9070 (N_9070,N_7932,N_7881);
nor U9071 (N_9071,N_7498,N_7127);
nand U9072 (N_9072,N_7497,N_7053);
or U9073 (N_9073,N_7236,N_6711);
nor U9074 (N_9074,N_7276,N_7475);
and U9075 (N_9075,N_7869,N_6045);
nand U9076 (N_9076,N_7904,N_6394);
and U9077 (N_9077,N_6066,N_6022);
and U9078 (N_9078,N_7925,N_7407);
and U9079 (N_9079,N_7192,N_6873);
and U9080 (N_9080,N_6953,N_6700);
nand U9081 (N_9081,N_7794,N_7407);
xor U9082 (N_9082,N_6743,N_7870);
nand U9083 (N_9083,N_7936,N_7164);
nand U9084 (N_9084,N_6253,N_7687);
xor U9085 (N_9085,N_6219,N_6628);
and U9086 (N_9086,N_7150,N_6660);
xor U9087 (N_9087,N_7360,N_6677);
and U9088 (N_9088,N_7817,N_7511);
xnor U9089 (N_9089,N_7986,N_7542);
nand U9090 (N_9090,N_7866,N_6905);
xnor U9091 (N_9091,N_6194,N_6763);
nor U9092 (N_9092,N_6015,N_6974);
nand U9093 (N_9093,N_7038,N_6106);
or U9094 (N_9094,N_6011,N_6464);
nand U9095 (N_9095,N_6989,N_7818);
and U9096 (N_9096,N_7734,N_6208);
nand U9097 (N_9097,N_6882,N_7084);
and U9098 (N_9098,N_6307,N_6644);
or U9099 (N_9099,N_6303,N_7039);
and U9100 (N_9100,N_6712,N_7283);
nor U9101 (N_9101,N_7153,N_6314);
nand U9102 (N_9102,N_6867,N_6749);
nor U9103 (N_9103,N_6608,N_7839);
or U9104 (N_9104,N_7333,N_7305);
xnor U9105 (N_9105,N_6644,N_7646);
and U9106 (N_9106,N_7250,N_7304);
nor U9107 (N_9107,N_6702,N_7023);
nor U9108 (N_9108,N_6945,N_7326);
and U9109 (N_9109,N_6666,N_7061);
nor U9110 (N_9110,N_7770,N_6922);
nor U9111 (N_9111,N_7611,N_7748);
or U9112 (N_9112,N_6200,N_6927);
nand U9113 (N_9113,N_6337,N_6811);
nor U9114 (N_9114,N_6204,N_6404);
nor U9115 (N_9115,N_6213,N_7789);
nor U9116 (N_9116,N_6818,N_7323);
xor U9117 (N_9117,N_7256,N_6410);
nor U9118 (N_9118,N_7198,N_6965);
or U9119 (N_9119,N_6529,N_7525);
nand U9120 (N_9120,N_7939,N_6668);
nand U9121 (N_9121,N_7660,N_7499);
nor U9122 (N_9122,N_6573,N_7545);
or U9123 (N_9123,N_7770,N_6541);
or U9124 (N_9124,N_7781,N_7230);
nor U9125 (N_9125,N_7888,N_7032);
nand U9126 (N_9126,N_7724,N_6386);
nand U9127 (N_9127,N_7976,N_6689);
nand U9128 (N_9128,N_6928,N_7455);
xnor U9129 (N_9129,N_7241,N_7532);
nand U9130 (N_9130,N_7349,N_7592);
and U9131 (N_9131,N_7754,N_6614);
nand U9132 (N_9132,N_7587,N_6600);
and U9133 (N_9133,N_7512,N_6155);
nor U9134 (N_9134,N_6861,N_7396);
nor U9135 (N_9135,N_7675,N_7157);
nor U9136 (N_9136,N_7187,N_7766);
nand U9137 (N_9137,N_6375,N_7055);
xor U9138 (N_9138,N_7847,N_6218);
and U9139 (N_9139,N_7656,N_7390);
nor U9140 (N_9140,N_7941,N_7577);
xor U9141 (N_9141,N_7566,N_6271);
and U9142 (N_9142,N_6953,N_6856);
nor U9143 (N_9143,N_7955,N_7777);
and U9144 (N_9144,N_7383,N_7486);
xnor U9145 (N_9145,N_7526,N_7627);
nand U9146 (N_9146,N_6223,N_6293);
nand U9147 (N_9147,N_7232,N_7562);
nor U9148 (N_9148,N_6209,N_6703);
xor U9149 (N_9149,N_6888,N_6526);
nor U9150 (N_9150,N_7990,N_7831);
xor U9151 (N_9151,N_7637,N_6088);
nand U9152 (N_9152,N_7511,N_6863);
and U9153 (N_9153,N_6148,N_6910);
nand U9154 (N_9154,N_6443,N_7034);
nor U9155 (N_9155,N_6236,N_6985);
or U9156 (N_9156,N_7102,N_7870);
nand U9157 (N_9157,N_6821,N_7712);
xnor U9158 (N_9158,N_7701,N_7968);
nand U9159 (N_9159,N_6582,N_6573);
nor U9160 (N_9160,N_7691,N_7094);
xor U9161 (N_9161,N_7555,N_7835);
and U9162 (N_9162,N_6934,N_7017);
xor U9163 (N_9163,N_7325,N_6587);
nor U9164 (N_9164,N_7957,N_7911);
nor U9165 (N_9165,N_6482,N_7402);
nor U9166 (N_9166,N_7378,N_7287);
and U9167 (N_9167,N_6204,N_6210);
or U9168 (N_9168,N_6744,N_6970);
and U9169 (N_9169,N_7651,N_6548);
xor U9170 (N_9170,N_6169,N_6103);
or U9171 (N_9171,N_7303,N_6303);
xnor U9172 (N_9172,N_6907,N_6521);
nor U9173 (N_9173,N_6157,N_6250);
or U9174 (N_9174,N_6348,N_7890);
xor U9175 (N_9175,N_7222,N_7213);
or U9176 (N_9176,N_6401,N_6209);
and U9177 (N_9177,N_7671,N_6391);
nor U9178 (N_9178,N_7966,N_7514);
or U9179 (N_9179,N_6362,N_7649);
nand U9180 (N_9180,N_7627,N_6990);
nand U9181 (N_9181,N_7304,N_7793);
nand U9182 (N_9182,N_6675,N_7277);
xor U9183 (N_9183,N_6600,N_6833);
or U9184 (N_9184,N_6274,N_6624);
nand U9185 (N_9185,N_6794,N_6125);
nor U9186 (N_9186,N_6737,N_7847);
nand U9187 (N_9187,N_7686,N_6921);
xor U9188 (N_9188,N_7567,N_6958);
xnor U9189 (N_9189,N_6494,N_7269);
nand U9190 (N_9190,N_6598,N_6593);
or U9191 (N_9191,N_7732,N_6203);
xnor U9192 (N_9192,N_6633,N_6970);
or U9193 (N_9193,N_7647,N_6676);
xnor U9194 (N_9194,N_7723,N_7733);
or U9195 (N_9195,N_6528,N_6271);
nor U9196 (N_9196,N_7162,N_6671);
xnor U9197 (N_9197,N_7407,N_6548);
and U9198 (N_9198,N_6448,N_6353);
nor U9199 (N_9199,N_6264,N_6156);
xor U9200 (N_9200,N_6330,N_6656);
nor U9201 (N_9201,N_6279,N_6049);
or U9202 (N_9202,N_6438,N_7491);
or U9203 (N_9203,N_7037,N_6234);
nor U9204 (N_9204,N_7511,N_7971);
nand U9205 (N_9205,N_6672,N_6887);
nand U9206 (N_9206,N_7815,N_6281);
nor U9207 (N_9207,N_6858,N_7810);
or U9208 (N_9208,N_7717,N_7282);
xor U9209 (N_9209,N_6590,N_7653);
xor U9210 (N_9210,N_7610,N_7296);
or U9211 (N_9211,N_7007,N_6371);
and U9212 (N_9212,N_7286,N_6589);
xor U9213 (N_9213,N_7075,N_6041);
nor U9214 (N_9214,N_7789,N_7880);
nor U9215 (N_9215,N_7458,N_7829);
nand U9216 (N_9216,N_7336,N_6241);
and U9217 (N_9217,N_6610,N_7573);
nor U9218 (N_9218,N_7968,N_6477);
or U9219 (N_9219,N_6217,N_7709);
nand U9220 (N_9220,N_6890,N_7762);
nor U9221 (N_9221,N_6119,N_6755);
xnor U9222 (N_9222,N_6431,N_7529);
nand U9223 (N_9223,N_6454,N_6745);
or U9224 (N_9224,N_6413,N_6430);
xor U9225 (N_9225,N_6535,N_7071);
xor U9226 (N_9226,N_6731,N_7926);
and U9227 (N_9227,N_7966,N_6199);
nor U9228 (N_9228,N_7859,N_7235);
or U9229 (N_9229,N_7659,N_7623);
or U9230 (N_9230,N_6821,N_6404);
nand U9231 (N_9231,N_7357,N_6298);
nand U9232 (N_9232,N_7814,N_6445);
nand U9233 (N_9233,N_6099,N_7918);
or U9234 (N_9234,N_6293,N_7896);
nand U9235 (N_9235,N_7483,N_7565);
nand U9236 (N_9236,N_6944,N_7103);
or U9237 (N_9237,N_6083,N_7854);
or U9238 (N_9238,N_7224,N_6202);
nor U9239 (N_9239,N_7494,N_7364);
nand U9240 (N_9240,N_7664,N_6052);
or U9241 (N_9241,N_7296,N_7989);
nor U9242 (N_9242,N_6137,N_6381);
or U9243 (N_9243,N_7362,N_6169);
and U9244 (N_9244,N_6797,N_6603);
xor U9245 (N_9245,N_7962,N_6158);
xnor U9246 (N_9246,N_7523,N_6102);
xnor U9247 (N_9247,N_7245,N_6147);
nor U9248 (N_9248,N_7973,N_6479);
nor U9249 (N_9249,N_6101,N_6380);
and U9250 (N_9250,N_7648,N_7831);
xnor U9251 (N_9251,N_6822,N_7668);
or U9252 (N_9252,N_6018,N_6104);
or U9253 (N_9253,N_7529,N_7804);
nor U9254 (N_9254,N_6343,N_6722);
nand U9255 (N_9255,N_6416,N_7912);
nand U9256 (N_9256,N_7812,N_6140);
nand U9257 (N_9257,N_6206,N_6521);
and U9258 (N_9258,N_7706,N_6258);
nand U9259 (N_9259,N_6143,N_7539);
nor U9260 (N_9260,N_6016,N_6839);
or U9261 (N_9261,N_6320,N_6354);
nor U9262 (N_9262,N_6627,N_6659);
or U9263 (N_9263,N_7422,N_6445);
and U9264 (N_9264,N_6604,N_6045);
nand U9265 (N_9265,N_7319,N_6378);
and U9266 (N_9266,N_6075,N_7643);
and U9267 (N_9267,N_7300,N_7404);
or U9268 (N_9268,N_6653,N_7013);
xnor U9269 (N_9269,N_7068,N_6458);
and U9270 (N_9270,N_7373,N_6682);
nor U9271 (N_9271,N_7376,N_7463);
and U9272 (N_9272,N_7173,N_6882);
and U9273 (N_9273,N_6115,N_7095);
nand U9274 (N_9274,N_6612,N_6851);
or U9275 (N_9275,N_7660,N_7826);
xnor U9276 (N_9276,N_7515,N_6719);
xnor U9277 (N_9277,N_7383,N_7566);
nand U9278 (N_9278,N_7160,N_7748);
or U9279 (N_9279,N_6212,N_6180);
xnor U9280 (N_9280,N_7757,N_6125);
nor U9281 (N_9281,N_7723,N_6219);
or U9282 (N_9282,N_6409,N_7200);
nand U9283 (N_9283,N_7659,N_6468);
and U9284 (N_9284,N_6923,N_7504);
nand U9285 (N_9285,N_7854,N_7141);
or U9286 (N_9286,N_7537,N_6392);
nor U9287 (N_9287,N_7343,N_7164);
xnor U9288 (N_9288,N_6046,N_7912);
and U9289 (N_9289,N_7665,N_6720);
and U9290 (N_9290,N_7236,N_6645);
nor U9291 (N_9291,N_6009,N_6084);
nand U9292 (N_9292,N_7533,N_6599);
nand U9293 (N_9293,N_7509,N_7562);
nor U9294 (N_9294,N_6955,N_7132);
xor U9295 (N_9295,N_7403,N_7724);
and U9296 (N_9296,N_6871,N_7488);
xor U9297 (N_9297,N_7684,N_7092);
and U9298 (N_9298,N_6016,N_6007);
xnor U9299 (N_9299,N_6625,N_6274);
xnor U9300 (N_9300,N_7785,N_6450);
and U9301 (N_9301,N_7741,N_7856);
nand U9302 (N_9302,N_6765,N_7405);
and U9303 (N_9303,N_6785,N_7579);
or U9304 (N_9304,N_6182,N_6490);
xnor U9305 (N_9305,N_6461,N_6176);
nand U9306 (N_9306,N_7399,N_7951);
nor U9307 (N_9307,N_6477,N_7216);
and U9308 (N_9308,N_6720,N_6948);
nor U9309 (N_9309,N_7619,N_6673);
or U9310 (N_9310,N_6615,N_7618);
xnor U9311 (N_9311,N_7971,N_6301);
nor U9312 (N_9312,N_7546,N_6302);
or U9313 (N_9313,N_6810,N_7490);
or U9314 (N_9314,N_6683,N_7627);
nor U9315 (N_9315,N_7836,N_7871);
or U9316 (N_9316,N_7481,N_7476);
nor U9317 (N_9317,N_6660,N_7304);
nor U9318 (N_9318,N_7568,N_7422);
and U9319 (N_9319,N_6709,N_6421);
nor U9320 (N_9320,N_6521,N_7930);
nand U9321 (N_9321,N_6183,N_7155);
nand U9322 (N_9322,N_6510,N_7301);
nor U9323 (N_9323,N_6527,N_7808);
or U9324 (N_9324,N_6475,N_6485);
xor U9325 (N_9325,N_6457,N_6473);
xor U9326 (N_9326,N_7340,N_6287);
nand U9327 (N_9327,N_7001,N_6171);
nor U9328 (N_9328,N_6716,N_7494);
and U9329 (N_9329,N_7929,N_6938);
xor U9330 (N_9330,N_7710,N_6089);
nor U9331 (N_9331,N_7262,N_7473);
nor U9332 (N_9332,N_6612,N_6771);
and U9333 (N_9333,N_7659,N_6121);
xnor U9334 (N_9334,N_7497,N_6662);
or U9335 (N_9335,N_7497,N_6510);
nor U9336 (N_9336,N_7867,N_7660);
nor U9337 (N_9337,N_6298,N_7124);
nor U9338 (N_9338,N_7977,N_6127);
or U9339 (N_9339,N_7518,N_7292);
or U9340 (N_9340,N_7456,N_7833);
nor U9341 (N_9341,N_6145,N_7414);
or U9342 (N_9342,N_7474,N_7781);
nand U9343 (N_9343,N_6846,N_6203);
or U9344 (N_9344,N_6164,N_7792);
nor U9345 (N_9345,N_7598,N_7457);
xor U9346 (N_9346,N_7581,N_7580);
nor U9347 (N_9347,N_7407,N_7124);
xor U9348 (N_9348,N_7968,N_7408);
xnor U9349 (N_9349,N_7901,N_7104);
nor U9350 (N_9350,N_6874,N_6424);
or U9351 (N_9351,N_7345,N_6731);
nand U9352 (N_9352,N_7358,N_7867);
nor U9353 (N_9353,N_6604,N_7642);
nor U9354 (N_9354,N_6717,N_6892);
and U9355 (N_9355,N_6201,N_6168);
xnor U9356 (N_9356,N_7245,N_6526);
or U9357 (N_9357,N_6142,N_6558);
and U9358 (N_9358,N_7193,N_7111);
nor U9359 (N_9359,N_7862,N_6740);
xnor U9360 (N_9360,N_6870,N_6728);
xor U9361 (N_9361,N_7439,N_7413);
nand U9362 (N_9362,N_7429,N_7800);
and U9363 (N_9363,N_7461,N_6873);
or U9364 (N_9364,N_7749,N_7119);
nor U9365 (N_9365,N_7116,N_6589);
nor U9366 (N_9366,N_7712,N_7786);
nand U9367 (N_9367,N_7949,N_6695);
and U9368 (N_9368,N_7782,N_6737);
nand U9369 (N_9369,N_6381,N_6809);
xor U9370 (N_9370,N_6596,N_6893);
nor U9371 (N_9371,N_6015,N_7576);
xnor U9372 (N_9372,N_6367,N_6130);
and U9373 (N_9373,N_7866,N_7741);
and U9374 (N_9374,N_7272,N_6563);
xor U9375 (N_9375,N_6561,N_7263);
and U9376 (N_9376,N_6551,N_6831);
and U9377 (N_9377,N_7278,N_6441);
and U9378 (N_9378,N_7644,N_7154);
and U9379 (N_9379,N_6400,N_6362);
nor U9380 (N_9380,N_7923,N_6145);
xnor U9381 (N_9381,N_6097,N_6526);
nand U9382 (N_9382,N_7105,N_7139);
and U9383 (N_9383,N_6836,N_7340);
nand U9384 (N_9384,N_6406,N_7059);
nand U9385 (N_9385,N_6901,N_6010);
xnor U9386 (N_9386,N_7982,N_6373);
nor U9387 (N_9387,N_6415,N_7387);
xor U9388 (N_9388,N_7396,N_7853);
nor U9389 (N_9389,N_6352,N_6903);
and U9390 (N_9390,N_6766,N_6072);
nand U9391 (N_9391,N_6169,N_6318);
xnor U9392 (N_9392,N_7447,N_7477);
xor U9393 (N_9393,N_6735,N_6515);
or U9394 (N_9394,N_7661,N_7697);
xor U9395 (N_9395,N_6952,N_7105);
or U9396 (N_9396,N_7225,N_7598);
xor U9397 (N_9397,N_6375,N_7156);
nor U9398 (N_9398,N_6035,N_6945);
and U9399 (N_9399,N_7359,N_6445);
and U9400 (N_9400,N_6265,N_6106);
and U9401 (N_9401,N_6932,N_6188);
and U9402 (N_9402,N_6523,N_7305);
and U9403 (N_9403,N_7201,N_6169);
and U9404 (N_9404,N_7013,N_7321);
nor U9405 (N_9405,N_7855,N_7186);
nor U9406 (N_9406,N_6918,N_6757);
xnor U9407 (N_9407,N_6933,N_6424);
xnor U9408 (N_9408,N_7101,N_6483);
nor U9409 (N_9409,N_6090,N_6371);
nor U9410 (N_9410,N_7340,N_7634);
or U9411 (N_9411,N_7888,N_6466);
xor U9412 (N_9412,N_7939,N_6232);
xnor U9413 (N_9413,N_6196,N_6102);
and U9414 (N_9414,N_7855,N_7916);
xor U9415 (N_9415,N_6020,N_6379);
or U9416 (N_9416,N_7782,N_7538);
and U9417 (N_9417,N_7890,N_7855);
nand U9418 (N_9418,N_6028,N_7470);
xnor U9419 (N_9419,N_7255,N_6197);
xnor U9420 (N_9420,N_6656,N_7189);
and U9421 (N_9421,N_7684,N_7272);
nor U9422 (N_9422,N_7409,N_6192);
or U9423 (N_9423,N_6511,N_7359);
or U9424 (N_9424,N_6179,N_6465);
xnor U9425 (N_9425,N_6065,N_7644);
and U9426 (N_9426,N_6469,N_6567);
xnor U9427 (N_9427,N_7916,N_6474);
xnor U9428 (N_9428,N_7985,N_6479);
nand U9429 (N_9429,N_7362,N_7392);
xnor U9430 (N_9430,N_6902,N_6791);
nand U9431 (N_9431,N_6993,N_7890);
and U9432 (N_9432,N_7564,N_7278);
and U9433 (N_9433,N_6444,N_7188);
nand U9434 (N_9434,N_7782,N_6854);
nor U9435 (N_9435,N_7657,N_6572);
nand U9436 (N_9436,N_6027,N_7190);
nand U9437 (N_9437,N_7215,N_7534);
and U9438 (N_9438,N_7925,N_6849);
nand U9439 (N_9439,N_6334,N_6262);
nor U9440 (N_9440,N_7632,N_6462);
and U9441 (N_9441,N_7578,N_6884);
xor U9442 (N_9442,N_6697,N_6743);
and U9443 (N_9443,N_6571,N_7754);
xor U9444 (N_9444,N_6228,N_7349);
or U9445 (N_9445,N_7351,N_7618);
xnor U9446 (N_9446,N_6726,N_7508);
nor U9447 (N_9447,N_6898,N_6521);
xnor U9448 (N_9448,N_7456,N_6147);
or U9449 (N_9449,N_6056,N_6906);
or U9450 (N_9450,N_6226,N_6980);
nor U9451 (N_9451,N_6551,N_7546);
xnor U9452 (N_9452,N_6672,N_6527);
xnor U9453 (N_9453,N_6646,N_7038);
nor U9454 (N_9454,N_6677,N_7222);
and U9455 (N_9455,N_7646,N_6318);
and U9456 (N_9456,N_6507,N_6792);
xnor U9457 (N_9457,N_7300,N_7841);
or U9458 (N_9458,N_6764,N_7414);
or U9459 (N_9459,N_6275,N_6250);
or U9460 (N_9460,N_6237,N_6827);
and U9461 (N_9461,N_7191,N_6427);
xor U9462 (N_9462,N_7032,N_7993);
nor U9463 (N_9463,N_6547,N_7423);
nand U9464 (N_9464,N_6032,N_6619);
nand U9465 (N_9465,N_6417,N_7554);
nand U9466 (N_9466,N_7719,N_6177);
or U9467 (N_9467,N_7203,N_6172);
and U9468 (N_9468,N_6340,N_7139);
nand U9469 (N_9469,N_7356,N_7312);
nand U9470 (N_9470,N_6675,N_7581);
or U9471 (N_9471,N_7653,N_6910);
or U9472 (N_9472,N_7076,N_6939);
nand U9473 (N_9473,N_7354,N_6174);
nor U9474 (N_9474,N_7546,N_7218);
xor U9475 (N_9475,N_6954,N_7178);
xnor U9476 (N_9476,N_6238,N_7977);
nor U9477 (N_9477,N_6745,N_7413);
nor U9478 (N_9478,N_6069,N_6123);
xnor U9479 (N_9479,N_7704,N_6055);
or U9480 (N_9480,N_7509,N_7814);
nand U9481 (N_9481,N_7922,N_6238);
nand U9482 (N_9482,N_6100,N_6006);
or U9483 (N_9483,N_6993,N_7854);
nor U9484 (N_9484,N_6293,N_6203);
xor U9485 (N_9485,N_6299,N_7029);
or U9486 (N_9486,N_7303,N_7518);
nand U9487 (N_9487,N_6603,N_7830);
nand U9488 (N_9488,N_6735,N_6844);
nand U9489 (N_9489,N_6490,N_7298);
nand U9490 (N_9490,N_6154,N_7751);
or U9491 (N_9491,N_6755,N_7573);
nand U9492 (N_9492,N_6752,N_6493);
and U9493 (N_9493,N_6798,N_6347);
and U9494 (N_9494,N_6418,N_6203);
nor U9495 (N_9495,N_6801,N_6425);
xor U9496 (N_9496,N_6124,N_7488);
and U9497 (N_9497,N_7788,N_6377);
nor U9498 (N_9498,N_7814,N_7128);
and U9499 (N_9499,N_6459,N_6807);
and U9500 (N_9500,N_6873,N_7738);
xor U9501 (N_9501,N_7038,N_6400);
nor U9502 (N_9502,N_7287,N_6794);
or U9503 (N_9503,N_6918,N_7805);
nor U9504 (N_9504,N_7118,N_7559);
and U9505 (N_9505,N_7410,N_7941);
nand U9506 (N_9506,N_7274,N_7016);
xnor U9507 (N_9507,N_6915,N_7093);
or U9508 (N_9508,N_7107,N_7265);
nor U9509 (N_9509,N_6243,N_7760);
or U9510 (N_9510,N_6942,N_7838);
and U9511 (N_9511,N_7515,N_6041);
and U9512 (N_9512,N_7892,N_6448);
and U9513 (N_9513,N_6060,N_7825);
and U9514 (N_9514,N_7672,N_6908);
or U9515 (N_9515,N_7055,N_6271);
xor U9516 (N_9516,N_7800,N_7924);
nor U9517 (N_9517,N_7520,N_7637);
nand U9518 (N_9518,N_6814,N_7558);
nor U9519 (N_9519,N_6835,N_6599);
nand U9520 (N_9520,N_6445,N_7934);
xnor U9521 (N_9521,N_7021,N_7645);
xor U9522 (N_9522,N_7719,N_7772);
nand U9523 (N_9523,N_7369,N_7292);
nand U9524 (N_9524,N_6611,N_7351);
or U9525 (N_9525,N_7985,N_6607);
nor U9526 (N_9526,N_6952,N_6115);
nand U9527 (N_9527,N_6112,N_7829);
nor U9528 (N_9528,N_6017,N_7160);
nor U9529 (N_9529,N_6884,N_6545);
xor U9530 (N_9530,N_7242,N_6081);
xnor U9531 (N_9531,N_7206,N_7233);
nor U9532 (N_9532,N_7808,N_7011);
and U9533 (N_9533,N_7942,N_7790);
or U9534 (N_9534,N_7305,N_6473);
and U9535 (N_9535,N_7324,N_6978);
and U9536 (N_9536,N_7805,N_6131);
xnor U9537 (N_9537,N_7805,N_7436);
nor U9538 (N_9538,N_7217,N_6382);
nor U9539 (N_9539,N_6966,N_6363);
xnor U9540 (N_9540,N_7853,N_6005);
xnor U9541 (N_9541,N_7413,N_6629);
or U9542 (N_9542,N_6281,N_7550);
xor U9543 (N_9543,N_7124,N_6981);
and U9544 (N_9544,N_6987,N_6585);
and U9545 (N_9545,N_7177,N_6133);
xnor U9546 (N_9546,N_7757,N_7670);
nor U9547 (N_9547,N_6489,N_6881);
xnor U9548 (N_9548,N_6117,N_7913);
xor U9549 (N_9549,N_7758,N_7121);
and U9550 (N_9550,N_7891,N_6451);
nand U9551 (N_9551,N_6015,N_7073);
nand U9552 (N_9552,N_6670,N_6793);
nand U9553 (N_9553,N_7593,N_6265);
nand U9554 (N_9554,N_6992,N_7535);
nor U9555 (N_9555,N_7823,N_6333);
xnor U9556 (N_9556,N_7595,N_6435);
nor U9557 (N_9557,N_6515,N_7121);
xnor U9558 (N_9558,N_7724,N_7566);
or U9559 (N_9559,N_6940,N_6616);
xnor U9560 (N_9560,N_6746,N_6311);
and U9561 (N_9561,N_6127,N_7365);
or U9562 (N_9562,N_6524,N_7349);
nor U9563 (N_9563,N_7389,N_6304);
and U9564 (N_9564,N_7294,N_6835);
xnor U9565 (N_9565,N_7911,N_7520);
nand U9566 (N_9566,N_6921,N_7618);
nand U9567 (N_9567,N_6592,N_6608);
or U9568 (N_9568,N_6213,N_6647);
nand U9569 (N_9569,N_7530,N_6185);
or U9570 (N_9570,N_6308,N_6352);
or U9571 (N_9571,N_7151,N_6151);
nand U9572 (N_9572,N_7607,N_6177);
nor U9573 (N_9573,N_7892,N_7133);
or U9574 (N_9574,N_6057,N_6555);
and U9575 (N_9575,N_7725,N_6535);
nand U9576 (N_9576,N_7310,N_6663);
xor U9577 (N_9577,N_6351,N_7574);
nor U9578 (N_9578,N_7753,N_7458);
nor U9579 (N_9579,N_7296,N_6931);
xor U9580 (N_9580,N_7084,N_7091);
nor U9581 (N_9581,N_6408,N_7635);
and U9582 (N_9582,N_7547,N_6124);
xor U9583 (N_9583,N_7870,N_7787);
nand U9584 (N_9584,N_6117,N_6593);
and U9585 (N_9585,N_7565,N_7811);
nor U9586 (N_9586,N_6891,N_7249);
and U9587 (N_9587,N_7867,N_6070);
or U9588 (N_9588,N_7221,N_6843);
or U9589 (N_9589,N_7345,N_6709);
or U9590 (N_9590,N_7872,N_6393);
xor U9591 (N_9591,N_7204,N_6878);
or U9592 (N_9592,N_7827,N_6784);
and U9593 (N_9593,N_7470,N_6972);
nand U9594 (N_9594,N_6069,N_6441);
xnor U9595 (N_9595,N_7272,N_7045);
or U9596 (N_9596,N_7064,N_7772);
or U9597 (N_9597,N_7765,N_7498);
nand U9598 (N_9598,N_6733,N_6952);
nor U9599 (N_9599,N_7721,N_7790);
and U9600 (N_9600,N_6953,N_7170);
and U9601 (N_9601,N_6888,N_7673);
xor U9602 (N_9602,N_6176,N_6061);
or U9603 (N_9603,N_7447,N_7094);
nor U9604 (N_9604,N_7972,N_6454);
and U9605 (N_9605,N_6615,N_7563);
and U9606 (N_9606,N_6984,N_6462);
or U9607 (N_9607,N_6935,N_6893);
nand U9608 (N_9608,N_6907,N_6221);
nand U9609 (N_9609,N_6069,N_7538);
nor U9610 (N_9610,N_6557,N_6611);
nand U9611 (N_9611,N_7394,N_6577);
or U9612 (N_9612,N_6038,N_7132);
xor U9613 (N_9613,N_6027,N_7541);
or U9614 (N_9614,N_6629,N_6475);
or U9615 (N_9615,N_7468,N_6092);
nor U9616 (N_9616,N_6576,N_6718);
xor U9617 (N_9617,N_7854,N_6288);
nor U9618 (N_9618,N_7372,N_7446);
xnor U9619 (N_9619,N_6932,N_7261);
nand U9620 (N_9620,N_6987,N_7128);
and U9621 (N_9621,N_7595,N_7570);
and U9622 (N_9622,N_7251,N_7605);
xor U9623 (N_9623,N_6405,N_6828);
or U9624 (N_9624,N_7952,N_7117);
nand U9625 (N_9625,N_6392,N_7275);
nand U9626 (N_9626,N_7840,N_6493);
or U9627 (N_9627,N_7975,N_6645);
xor U9628 (N_9628,N_7043,N_6912);
xor U9629 (N_9629,N_6870,N_6952);
nand U9630 (N_9630,N_7522,N_6664);
nor U9631 (N_9631,N_6724,N_7263);
xnor U9632 (N_9632,N_7848,N_7291);
xor U9633 (N_9633,N_6606,N_6758);
xor U9634 (N_9634,N_7564,N_7177);
or U9635 (N_9635,N_7334,N_7354);
nand U9636 (N_9636,N_7411,N_6263);
or U9637 (N_9637,N_6897,N_6247);
and U9638 (N_9638,N_7085,N_6875);
or U9639 (N_9639,N_7122,N_7480);
nand U9640 (N_9640,N_7296,N_6386);
or U9641 (N_9641,N_7581,N_7349);
xnor U9642 (N_9642,N_7183,N_6920);
xor U9643 (N_9643,N_6403,N_7496);
xnor U9644 (N_9644,N_7785,N_6401);
nor U9645 (N_9645,N_7133,N_7183);
or U9646 (N_9646,N_6520,N_6996);
xnor U9647 (N_9647,N_7909,N_6087);
xnor U9648 (N_9648,N_7349,N_7393);
nor U9649 (N_9649,N_7396,N_7213);
or U9650 (N_9650,N_6705,N_6513);
or U9651 (N_9651,N_6396,N_7536);
or U9652 (N_9652,N_7355,N_6733);
xor U9653 (N_9653,N_6417,N_6434);
or U9654 (N_9654,N_7955,N_7428);
nor U9655 (N_9655,N_7882,N_7751);
xor U9656 (N_9656,N_7527,N_7193);
and U9657 (N_9657,N_6672,N_6388);
nand U9658 (N_9658,N_6600,N_7125);
xor U9659 (N_9659,N_7727,N_6617);
nor U9660 (N_9660,N_7529,N_6104);
and U9661 (N_9661,N_6020,N_6046);
and U9662 (N_9662,N_6948,N_6028);
and U9663 (N_9663,N_7294,N_7917);
xor U9664 (N_9664,N_7249,N_7876);
or U9665 (N_9665,N_6320,N_7008);
nor U9666 (N_9666,N_7036,N_7732);
nor U9667 (N_9667,N_6681,N_7972);
or U9668 (N_9668,N_6447,N_7902);
or U9669 (N_9669,N_7280,N_7315);
or U9670 (N_9670,N_6728,N_7263);
or U9671 (N_9671,N_6512,N_7543);
xnor U9672 (N_9672,N_7997,N_6873);
xnor U9673 (N_9673,N_6081,N_6610);
nor U9674 (N_9674,N_7369,N_6770);
xnor U9675 (N_9675,N_7573,N_7713);
xor U9676 (N_9676,N_7758,N_7952);
nand U9677 (N_9677,N_6510,N_6514);
nand U9678 (N_9678,N_7963,N_6681);
and U9679 (N_9679,N_7894,N_6159);
xnor U9680 (N_9680,N_7580,N_6010);
nand U9681 (N_9681,N_7877,N_7964);
and U9682 (N_9682,N_7313,N_7512);
xor U9683 (N_9683,N_6651,N_6801);
nor U9684 (N_9684,N_6688,N_6706);
nand U9685 (N_9685,N_6440,N_6435);
or U9686 (N_9686,N_6712,N_6472);
nor U9687 (N_9687,N_6554,N_7729);
and U9688 (N_9688,N_6906,N_7557);
nor U9689 (N_9689,N_7662,N_6133);
nor U9690 (N_9690,N_6182,N_7072);
or U9691 (N_9691,N_6641,N_7824);
nand U9692 (N_9692,N_7597,N_6812);
xor U9693 (N_9693,N_7301,N_6441);
nand U9694 (N_9694,N_6325,N_7250);
or U9695 (N_9695,N_6583,N_7125);
or U9696 (N_9696,N_7854,N_7184);
and U9697 (N_9697,N_6238,N_6124);
and U9698 (N_9698,N_7937,N_7505);
and U9699 (N_9699,N_7956,N_7966);
and U9700 (N_9700,N_6953,N_6022);
nor U9701 (N_9701,N_7786,N_6026);
xor U9702 (N_9702,N_7914,N_6754);
xnor U9703 (N_9703,N_7119,N_7706);
or U9704 (N_9704,N_7615,N_7060);
nor U9705 (N_9705,N_7947,N_7301);
and U9706 (N_9706,N_7596,N_7938);
and U9707 (N_9707,N_7114,N_6783);
nor U9708 (N_9708,N_7888,N_7892);
and U9709 (N_9709,N_7110,N_7409);
nand U9710 (N_9710,N_6987,N_6853);
and U9711 (N_9711,N_6758,N_7949);
and U9712 (N_9712,N_6369,N_6089);
or U9713 (N_9713,N_6506,N_7292);
or U9714 (N_9714,N_6380,N_6013);
and U9715 (N_9715,N_7891,N_6915);
nor U9716 (N_9716,N_6530,N_7278);
nor U9717 (N_9717,N_7360,N_6124);
or U9718 (N_9718,N_7916,N_7283);
nand U9719 (N_9719,N_7443,N_7480);
nor U9720 (N_9720,N_6260,N_7141);
xor U9721 (N_9721,N_7397,N_6701);
xor U9722 (N_9722,N_6339,N_7509);
nand U9723 (N_9723,N_7548,N_7585);
nor U9724 (N_9724,N_7924,N_7075);
nand U9725 (N_9725,N_6027,N_6353);
or U9726 (N_9726,N_7577,N_7125);
nand U9727 (N_9727,N_7969,N_6795);
nor U9728 (N_9728,N_7116,N_7073);
nand U9729 (N_9729,N_6526,N_6758);
or U9730 (N_9730,N_7367,N_7093);
nand U9731 (N_9731,N_7795,N_7387);
nor U9732 (N_9732,N_6047,N_6083);
xnor U9733 (N_9733,N_6876,N_6975);
or U9734 (N_9734,N_7369,N_6691);
or U9735 (N_9735,N_6531,N_7043);
nor U9736 (N_9736,N_6667,N_6454);
nor U9737 (N_9737,N_6116,N_6989);
nor U9738 (N_9738,N_7936,N_7114);
and U9739 (N_9739,N_7987,N_7128);
nor U9740 (N_9740,N_7831,N_7390);
xnor U9741 (N_9741,N_7794,N_7641);
or U9742 (N_9742,N_7183,N_6047);
or U9743 (N_9743,N_7496,N_7889);
and U9744 (N_9744,N_6963,N_7310);
nor U9745 (N_9745,N_6191,N_7177);
xor U9746 (N_9746,N_7914,N_6777);
nor U9747 (N_9747,N_7365,N_7226);
xnor U9748 (N_9748,N_6055,N_7138);
or U9749 (N_9749,N_6711,N_6502);
or U9750 (N_9750,N_7117,N_7404);
xnor U9751 (N_9751,N_7619,N_6684);
nand U9752 (N_9752,N_7556,N_7135);
xor U9753 (N_9753,N_6008,N_6374);
and U9754 (N_9754,N_6624,N_7096);
or U9755 (N_9755,N_6538,N_6092);
nor U9756 (N_9756,N_7343,N_7303);
nor U9757 (N_9757,N_7860,N_7420);
nor U9758 (N_9758,N_6239,N_6112);
nand U9759 (N_9759,N_7407,N_6170);
nor U9760 (N_9760,N_6918,N_6917);
nor U9761 (N_9761,N_6071,N_7356);
nand U9762 (N_9762,N_6595,N_6798);
nand U9763 (N_9763,N_6041,N_6934);
xnor U9764 (N_9764,N_7928,N_7337);
xor U9765 (N_9765,N_6564,N_7669);
and U9766 (N_9766,N_6354,N_6936);
nor U9767 (N_9767,N_7044,N_6867);
xor U9768 (N_9768,N_6484,N_7425);
nand U9769 (N_9769,N_6984,N_7580);
or U9770 (N_9770,N_6779,N_7425);
nor U9771 (N_9771,N_7291,N_6350);
and U9772 (N_9772,N_7182,N_6685);
or U9773 (N_9773,N_6648,N_6221);
nor U9774 (N_9774,N_6890,N_6455);
nand U9775 (N_9775,N_7984,N_7022);
xor U9776 (N_9776,N_6279,N_7993);
or U9777 (N_9777,N_6759,N_7437);
nor U9778 (N_9778,N_7003,N_6899);
xnor U9779 (N_9779,N_7915,N_7375);
nor U9780 (N_9780,N_7416,N_7397);
nor U9781 (N_9781,N_6686,N_6275);
or U9782 (N_9782,N_6420,N_7134);
nor U9783 (N_9783,N_6298,N_7069);
and U9784 (N_9784,N_6530,N_7859);
xnor U9785 (N_9785,N_7280,N_7858);
xnor U9786 (N_9786,N_6937,N_7253);
or U9787 (N_9787,N_7910,N_7126);
nor U9788 (N_9788,N_7711,N_6401);
and U9789 (N_9789,N_7482,N_7093);
xnor U9790 (N_9790,N_7430,N_7241);
xor U9791 (N_9791,N_6769,N_7448);
nand U9792 (N_9792,N_7382,N_7754);
xor U9793 (N_9793,N_7049,N_7510);
nor U9794 (N_9794,N_6348,N_6435);
xor U9795 (N_9795,N_6225,N_6047);
nand U9796 (N_9796,N_7678,N_7937);
nand U9797 (N_9797,N_7408,N_7446);
nor U9798 (N_9798,N_7953,N_6393);
nor U9799 (N_9799,N_6826,N_7035);
xnor U9800 (N_9800,N_7145,N_6977);
nor U9801 (N_9801,N_6549,N_6668);
or U9802 (N_9802,N_6791,N_7403);
xor U9803 (N_9803,N_6390,N_6479);
nand U9804 (N_9804,N_6246,N_6712);
nor U9805 (N_9805,N_6783,N_7434);
nor U9806 (N_9806,N_7623,N_6159);
and U9807 (N_9807,N_7715,N_7535);
xor U9808 (N_9808,N_6533,N_7860);
nor U9809 (N_9809,N_6500,N_6969);
or U9810 (N_9810,N_6070,N_6056);
and U9811 (N_9811,N_6534,N_7173);
nand U9812 (N_9812,N_6767,N_7910);
or U9813 (N_9813,N_6909,N_6792);
nor U9814 (N_9814,N_6403,N_7186);
or U9815 (N_9815,N_6781,N_7278);
nand U9816 (N_9816,N_6172,N_7318);
and U9817 (N_9817,N_6426,N_7061);
nor U9818 (N_9818,N_6740,N_6090);
and U9819 (N_9819,N_7574,N_7199);
nor U9820 (N_9820,N_7878,N_6861);
and U9821 (N_9821,N_6567,N_7791);
or U9822 (N_9822,N_6282,N_7245);
nor U9823 (N_9823,N_7288,N_7617);
or U9824 (N_9824,N_7765,N_6860);
nand U9825 (N_9825,N_6655,N_7668);
nand U9826 (N_9826,N_7014,N_6777);
nor U9827 (N_9827,N_6590,N_7234);
xor U9828 (N_9828,N_6007,N_6794);
nor U9829 (N_9829,N_7237,N_7321);
xor U9830 (N_9830,N_6929,N_7727);
and U9831 (N_9831,N_6858,N_6172);
nand U9832 (N_9832,N_6611,N_7990);
and U9833 (N_9833,N_7152,N_6686);
nor U9834 (N_9834,N_7967,N_7532);
nor U9835 (N_9835,N_7116,N_6012);
nand U9836 (N_9836,N_6649,N_6294);
xor U9837 (N_9837,N_7414,N_6827);
nand U9838 (N_9838,N_7963,N_7697);
nor U9839 (N_9839,N_7574,N_6047);
and U9840 (N_9840,N_7652,N_6578);
and U9841 (N_9841,N_7353,N_6476);
nor U9842 (N_9842,N_6760,N_7032);
nand U9843 (N_9843,N_7018,N_6415);
nor U9844 (N_9844,N_6071,N_6596);
or U9845 (N_9845,N_6090,N_7398);
and U9846 (N_9846,N_6901,N_6036);
xor U9847 (N_9847,N_7660,N_6741);
xor U9848 (N_9848,N_6322,N_7838);
nand U9849 (N_9849,N_7100,N_6908);
or U9850 (N_9850,N_6135,N_7217);
xnor U9851 (N_9851,N_7157,N_7135);
nor U9852 (N_9852,N_6753,N_6595);
nand U9853 (N_9853,N_7615,N_7532);
xnor U9854 (N_9854,N_6723,N_7936);
nor U9855 (N_9855,N_6846,N_6670);
and U9856 (N_9856,N_6576,N_6640);
and U9857 (N_9857,N_7371,N_7287);
and U9858 (N_9858,N_6588,N_7678);
xnor U9859 (N_9859,N_7517,N_7188);
and U9860 (N_9860,N_6580,N_6226);
or U9861 (N_9861,N_7828,N_7883);
or U9862 (N_9862,N_7775,N_7245);
or U9863 (N_9863,N_7184,N_7222);
nand U9864 (N_9864,N_6422,N_6759);
or U9865 (N_9865,N_7386,N_6151);
or U9866 (N_9866,N_7399,N_7416);
nand U9867 (N_9867,N_7418,N_7553);
xnor U9868 (N_9868,N_6451,N_6435);
xnor U9869 (N_9869,N_6058,N_7812);
or U9870 (N_9870,N_7821,N_7928);
xor U9871 (N_9871,N_7057,N_7944);
and U9872 (N_9872,N_6798,N_6686);
or U9873 (N_9873,N_6865,N_7842);
or U9874 (N_9874,N_6462,N_6765);
xnor U9875 (N_9875,N_6234,N_7929);
or U9876 (N_9876,N_6280,N_6774);
xor U9877 (N_9877,N_6557,N_6444);
nand U9878 (N_9878,N_6227,N_6345);
nor U9879 (N_9879,N_6538,N_7256);
or U9880 (N_9880,N_6669,N_6562);
xor U9881 (N_9881,N_7841,N_6876);
or U9882 (N_9882,N_6885,N_6082);
and U9883 (N_9883,N_6003,N_7164);
or U9884 (N_9884,N_6226,N_7623);
nor U9885 (N_9885,N_6407,N_6327);
nor U9886 (N_9886,N_7172,N_6221);
nand U9887 (N_9887,N_7638,N_7531);
and U9888 (N_9888,N_6427,N_6232);
xor U9889 (N_9889,N_6866,N_6223);
xor U9890 (N_9890,N_7671,N_7903);
or U9891 (N_9891,N_6689,N_7377);
nand U9892 (N_9892,N_7818,N_6068);
nor U9893 (N_9893,N_7346,N_7155);
nand U9894 (N_9894,N_7551,N_7047);
or U9895 (N_9895,N_7228,N_6366);
nand U9896 (N_9896,N_7139,N_6515);
nor U9897 (N_9897,N_6630,N_6565);
xnor U9898 (N_9898,N_7910,N_6186);
nand U9899 (N_9899,N_7017,N_7640);
nor U9900 (N_9900,N_6021,N_6659);
nand U9901 (N_9901,N_7100,N_6254);
nor U9902 (N_9902,N_6971,N_7089);
xor U9903 (N_9903,N_7190,N_7738);
nand U9904 (N_9904,N_6411,N_6312);
and U9905 (N_9905,N_6637,N_7402);
xor U9906 (N_9906,N_6179,N_7724);
and U9907 (N_9907,N_7187,N_7184);
or U9908 (N_9908,N_6098,N_6184);
or U9909 (N_9909,N_7625,N_7809);
nand U9910 (N_9910,N_7025,N_7688);
nand U9911 (N_9911,N_6618,N_7980);
xor U9912 (N_9912,N_6200,N_7428);
and U9913 (N_9913,N_7303,N_7212);
nand U9914 (N_9914,N_7206,N_6770);
and U9915 (N_9915,N_7730,N_6054);
or U9916 (N_9916,N_7192,N_6712);
nor U9917 (N_9917,N_6478,N_6002);
nor U9918 (N_9918,N_7451,N_6211);
nand U9919 (N_9919,N_7265,N_6275);
and U9920 (N_9920,N_6921,N_6880);
and U9921 (N_9921,N_7981,N_6741);
and U9922 (N_9922,N_7983,N_6938);
or U9923 (N_9923,N_6422,N_7310);
nor U9924 (N_9924,N_7081,N_6294);
nand U9925 (N_9925,N_7625,N_7315);
and U9926 (N_9926,N_6792,N_7572);
nand U9927 (N_9927,N_6381,N_6711);
xor U9928 (N_9928,N_7850,N_6443);
and U9929 (N_9929,N_6075,N_7191);
xnor U9930 (N_9930,N_7466,N_7594);
nand U9931 (N_9931,N_6647,N_7343);
nor U9932 (N_9932,N_7086,N_6534);
or U9933 (N_9933,N_7493,N_7251);
and U9934 (N_9934,N_7678,N_7340);
and U9935 (N_9935,N_6523,N_6683);
xor U9936 (N_9936,N_7307,N_7350);
xnor U9937 (N_9937,N_7840,N_6801);
nand U9938 (N_9938,N_6322,N_6302);
xor U9939 (N_9939,N_6330,N_7843);
nor U9940 (N_9940,N_6286,N_7296);
xnor U9941 (N_9941,N_6790,N_6658);
or U9942 (N_9942,N_7121,N_6497);
xnor U9943 (N_9943,N_7406,N_7852);
or U9944 (N_9944,N_6639,N_7999);
nand U9945 (N_9945,N_6546,N_7614);
or U9946 (N_9946,N_6965,N_6987);
nand U9947 (N_9947,N_6929,N_6435);
xnor U9948 (N_9948,N_6413,N_6526);
nand U9949 (N_9949,N_6617,N_7114);
nor U9950 (N_9950,N_6565,N_6504);
nand U9951 (N_9951,N_6181,N_7474);
xor U9952 (N_9952,N_6542,N_7464);
or U9953 (N_9953,N_6822,N_6921);
and U9954 (N_9954,N_6615,N_6111);
or U9955 (N_9955,N_6245,N_7459);
nor U9956 (N_9956,N_7068,N_6813);
or U9957 (N_9957,N_6585,N_6744);
nor U9958 (N_9958,N_7661,N_7430);
or U9959 (N_9959,N_6023,N_6298);
xor U9960 (N_9960,N_6552,N_6383);
nor U9961 (N_9961,N_7420,N_6126);
nand U9962 (N_9962,N_6312,N_7173);
nor U9963 (N_9963,N_7821,N_7200);
nor U9964 (N_9964,N_6168,N_7933);
nor U9965 (N_9965,N_6547,N_6838);
xor U9966 (N_9966,N_6849,N_7930);
and U9967 (N_9967,N_6548,N_6226);
nor U9968 (N_9968,N_7162,N_6829);
or U9969 (N_9969,N_6356,N_6709);
xnor U9970 (N_9970,N_6267,N_7267);
nor U9971 (N_9971,N_6023,N_7081);
nor U9972 (N_9972,N_6407,N_6881);
nand U9973 (N_9973,N_6635,N_6729);
or U9974 (N_9974,N_6456,N_6740);
xnor U9975 (N_9975,N_6247,N_6645);
and U9976 (N_9976,N_6133,N_7192);
or U9977 (N_9977,N_6816,N_7574);
and U9978 (N_9978,N_7905,N_7086);
or U9979 (N_9979,N_6720,N_7228);
nor U9980 (N_9980,N_7722,N_7002);
nor U9981 (N_9981,N_7582,N_6004);
or U9982 (N_9982,N_6055,N_6065);
or U9983 (N_9983,N_6706,N_6716);
and U9984 (N_9984,N_6112,N_7109);
or U9985 (N_9985,N_6900,N_7831);
and U9986 (N_9986,N_7119,N_6575);
or U9987 (N_9987,N_6279,N_6826);
xor U9988 (N_9988,N_7142,N_6655);
nand U9989 (N_9989,N_6367,N_7964);
xor U9990 (N_9990,N_7340,N_7970);
xnor U9991 (N_9991,N_6643,N_7676);
or U9992 (N_9992,N_6344,N_6462);
and U9993 (N_9993,N_6483,N_6171);
and U9994 (N_9994,N_6392,N_7794);
nor U9995 (N_9995,N_7555,N_7829);
nand U9996 (N_9996,N_7759,N_6669);
nand U9997 (N_9997,N_7059,N_6881);
xor U9998 (N_9998,N_7263,N_6892);
and U9999 (N_9999,N_7953,N_7177);
nor UO_0 (O_0,N_9886,N_9829);
nand UO_1 (O_1,N_9071,N_8072);
and UO_2 (O_2,N_8869,N_9279);
xnor UO_3 (O_3,N_9780,N_9882);
xnor UO_4 (O_4,N_8957,N_8434);
nor UO_5 (O_5,N_9718,N_8371);
and UO_6 (O_6,N_8192,N_8805);
xor UO_7 (O_7,N_8606,N_9660);
nand UO_8 (O_8,N_8472,N_8587);
xor UO_9 (O_9,N_8683,N_9356);
and UO_10 (O_10,N_8402,N_9327);
nor UO_11 (O_11,N_9685,N_8874);
nand UO_12 (O_12,N_8373,N_9234);
and UO_13 (O_13,N_8208,N_9790);
nand UO_14 (O_14,N_8172,N_8635);
xor UO_15 (O_15,N_9306,N_8995);
xor UO_16 (O_16,N_8568,N_9117);
nand UO_17 (O_17,N_9012,N_8761);
nand UO_18 (O_18,N_8582,N_9486);
or UO_19 (O_19,N_8897,N_8969);
nand UO_20 (O_20,N_8253,N_9241);
and UO_21 (O_21,N_9011,N_8425);
nor UO_22 (O_22,N_9971,N_8230);
nand UO_23 (O_23,N_9382,N_8421);
xnor UO_24 (O_24,N_8065,N_9345);
nand UO_25 (O_25,N_8609,N_8457);
nor UO_26 (O_26,N_8640,N_9165);
or UO_27 (O_27,N_8348,N_8738);
xnor UO_28 (O_28,N_9768,N_9263);
and UO_29 (O_29,N_9361,N_9126);
nand UO_30 (O_30,N_9713,N_8436);
and UO_31 (O_31,N_8357,N_8614);
nor UO_32 (O_32,N_9495,N_9357);
xor UO_33 (O_33,N_9462,N_9468);
nand UO_34 (O_34,N_9587,N_8814);
and UO_35 (O_35,N_8464,N_8615);
xnor UO_36 (O_36,N_9365,N_8682);
or UO_37 (O_37,N_9329,N_9593);
and UO_38 (O_38,N_8714,N_8727);
nor UO_39 (O_39,N_9230,N_8409);
xor UO_40 (O_40,N_8537,N_9251);
or UO_41 (O_41,N_9802,N_8119);
nand UO_42 (O_42,N_9852,N_9175);
or UO_43 (O_43,N_8277,N_8104);
xor UO_44 (O_44,N_8842,N_8400);
or UO_45 (O_45,N_9646,N_8859);
nor UO_46 (O_46,N_9027,N_8234);
nor UO_47 (O_47,N_8223,N_8908);
nand UO_48 (O_48,N_8783,N_8573);
or UO_49 (O_49,N_8315,N_9205);
xnor UO_50 (O_50,N_8649,N_9250);
xor UO_51 (O_51,N_9597,N_9368);
and UO_52 (O_52,N_8024,N_8204);
and UO_53 (O_53,N_8058,N_9615);
and UO_54 (O_54,N_8231,N_9331);
nor UO_55 (O_55,N_9400,N_8032);
nand UO_56 (O_56,N_9804,N_9019);
nand UO_57 (O_57,N_8066,N_9322);
nand UO_58 (O_58,N_9262,N_8796);
nand UO_59 (O_59,N_9044,N_8834);
nor UO_60 (O_60,N_8951,N_9152);
or UO_61 (O_61,N_8292,N_8790);
and UO_62 (O_62,N_8403,N_8379);
nor UO_63 (O_63,N_9995,N_9135);
and UO_64 (O_64,N_8644,N_9967);
nand UO_65 (O_65,N_8828,N_9679);
xor UO_66 (O_66,N_9063,N_8144);
xor UO_67 (O_67,N_9556,N_9808);
and UO_68 (O_68,N_8012,N_8651);
or UO_69 (O_69,N_9036,N_9417);
or UO_70 (O_70,N_9539,N_8362);
nor UO_71 (O_71,N_9403,N_8675);
nor UO_72 (O_72,N_9313,N_9483);
xnor UO_73 (O_73,N_9481,N_9965);
nand UO_74 (O_74,N_9692,N_8955);
or UO_75 (O_75,N_9610,N_8516);
or UO_76 (O_76,N_8732,N_8465);
nand UO_77 (O_77,N_9979,N_8755);
and UO_78 (O_78,N_8327,N_8647);
xor UO_79 (O_79,N_9138,N_9396);
or UO_80 (O_80,N_8345,N_9281);
nor UO_81 (O_81,N_9809,N_8343);
nand UO_82 (O_82,N_8171,N_8132);
or UO_83 (O_83,N_8366,N_9437);
nor UO_84 (O_84,N_9887,N_9835);
and UO_85 (O_85,N_8496,N_8070);
and UO_86 (O_86,N_9976,N_9687);
nand UO_87 (O_87,N_8607,N_8210);
nand UO_88 (O_88,N_8762,N_9451);
nor UO_89 (O_89,N_9163,N_8535);
nand UO_90 (O_90,N_9889,N_9140);
xnor UO_91 (O_91,N_9114,N_8905);
or UO_92 (O_92,N_8827,N_9649);
or UO_93 (O_93,N_8736,N_8696);
or UO_94 (O_94,N_9560,N_9868);
nand UO_95 (O_95,N_8351,N_9757);
nor UO_96 (O_96,N_8795,N_8939);
nor UO_97 (O_97,N_9208,N_9733);
and UO_98 (O_98,N_8456,N_9499);
nand UO_99 (O_99,N_9161,N_8352);
and UO_100 (O_100,N_8475,N_9880);
and UO_101 (O_101,N_9116,N_9360);
nand UO_102 (O_102,N_9332,N_8341);
or UO_103 (O_103,N_9201,N_9007);
xor UO_104 (O_104,N_9469,N_9746);
xor UO_105 (O_105,N_8140,N_8863);
nand UO_106 (O_106,N_8497,N_9876);
xnor UO_107 (O_107,N_8947,N_8554);
nor UO_108 (O_108,N_8984,N_9452);
nand UO_109 (O_109,N_8510,N_9002);
and UO_110 (O_110,N_9515,N_8722);
nand UO_111 (O_111,N_8663,N_9910);
xnor UO_112 (O_112,N_9257,N_9682);
xor UO_113 (O_113,N_9187,N_9789);
nor UO_114 (O_114,N_8639,N_9245);
nand UO_115 (O_115,N_9708,N_8617);
nand UO_116 (O_116,N_8260,N_9303);
and UO_117 (O_117,N_9869,N_9551);
xor UO_118 (O_118,N_9725,N_9270);
xor UO_119 (O_119,N_8128,N_8438);
and UO_120 (O_120,N_8093,N_9912);
nor UO_121 (O_121,N_9634,N_9355);
nand UO_122 (O_122,N_9778,N_8536);
nor UO_123 (O_123,N_8094,N_8023);
or UO_124 (O_124,N_8700,N_8306);
nand UO_125 (O_125,N_8698,N_8643);
xor UO_126 (O_126,N_8099,N_9045);
nand UO_127 (O_127,N_9944,N_8356);
or UO_128 (O_128,N_8953,N_9978);
nand UO_129 (O_129,N_8173,N_8062);
nor UO_130 (O_130,N_9948,N_8757);
nand UO_131 (O_131,N_9893,N_8278);
and UO_132 (O_132,N_9423,N_8913);
or UO_133 (O_133,N_8441,N_9074);
and UO_134 (O_134,N_8583,N_9955);
or UO_135 (O_135,N_9870,N_8848);
xor UO_136 (O_136,N_9238,N_9420);
nand UO_137 (O_137,N_8196,N_8887);
and UO_138 (O_138,N_9825,N_9534);
nand UO_139 (O_139,N_8991,N_9859);
xnor UO_140 (O_140,N_8177,N_8712);
nand UO_141 (O_141,N_9670,N_9716);
nand UO_142 (O_142,N_8322,N_8089);
and UO_143 (O_143,N_8836,N_9061);
or UO_144 (O_144,N_8560,N_9781);
nor UO_145 (O_145,N_9543,N_9213);
and UO_146 (O_146,N_9047,N_8669);
nor UO_147 (O_147,N_9374,N_9686);
or UO_148 (O_148,N_9337,N_8598);
nand UO_149 (O_149,N_9378,N_8988);
or UO_150 (O_150,N_9709,N_8120);
or UO_151 (O_151,N_9028,N_8867);
nand UO_152 (O_152,N_8075,N_9164);
nor UO_153 (O_153,N_8511,N_8862);
and UO_154 (O_154,N_9878,N_9542);
xnor UO_155 (O_155,N_8340,N_9226);
nor UO_156 (O_156,N_9305,N_8801);
or UO_157 (O_157,N_9093,N_8195);
and UO_158 (O_158,N_8390,N_9448);
nor UO_159 (O_159,N_9038,N_8243);
and UO_160 (O_160,N_9972,N_8244);
nand UO_161 (O_161,N_9179,N_8593);
or UO_162 (O_162,N_8746,N_8934);
or UO_163 (O_163,N_9631,N_8449);
xnor UO_164 (O_164,N_9252,N_8729);
and UO_165 (O_165,N_9980,N_8973);
xnor UO_166 (O_166,N_8518,N_9494);
and UO_167 (O_167,N_9983,N_9676);
and UO_168 (O_168,N_9017,N_8423);
nand UO_169 (O_169,N_8324,N_8215);
and UO_170 (O_170,N_8517,N_9970);
xor UO_171 (O_171,N_8291,N_8816);
nand UO_172 (O_172,N_8702,N_8300);
nor UO_173 (O_173,N_8183,N_9957);
xor UO_174 (O_174,N_9066,N_9029);
nor UO_175 (O_175,N_8787,N_9700);
or UO_176 (O_176,N_8227,N_8730);
and UO_177 (O_177,N_8671,N_9512);
nand UO_178 (O_178,N_8164,N_8478);
xnor UO_179 (O_179,N_8452,N_9703);
xor UO_180 (O_180,N_8445,N_8622);
nor UO_181 (O_181,N_8206,N_8558);
nand UO_182 (O_182,N_9237,N_8569);
xor UO_183 (O_183,N_8916,N_8411);
nor UO_184 (O_184,N_9376,N_9862);
xnor UO_185 (O_185,N_9614,N_8036);
and UO_186 (O_186,N_9656,N_8169);
and UO_187 (O_187,N_8604,N_8800);
and UO_188 (O_188,N_9411,N_8935);
or UO_189 (O_189,N_8274,N_9606);
nand UO_190 (O_190,N_8804,N_9582);
nor UO_191 (O_191,N_8338,N_9786);
and UO_192 (O_192,N_9056,N_8525);
and UO_193 (O_193,N_8484,N_9750);
xnor UO_194 (O_194,N_9561,N_9581);
xnor UO_195 (O_195,N_9013,N_9014);
nand UO_196 (O_196,N_8739,N_9212);
and UO_197 (O_197,N_8364,N_8613);
nand UO_198 (O_198,N_8228,N_9247);
or UO_199 (O_199,N_8754,N_8301);
and UO_200 (O_200,N_9603,N_9792);
nand UO_201 (O_201,N_9959,N_9583);
nor UO_202 (O_202,N_8067,N_9339);
nand UO_203 (O_203,N_8764,N_9974);
nand UO_204 (O_204,N_8384,N_8311);
or UO_205 (O_205,N_9295,N_8427);
and UO_206 (O_206,N_9744,N_8581);
and UO_207 (O_207,N_9570,N_9046);
xnor UO_208 (O_208,N_8589,N_9460);
nor UO_209 (O_209,N_9067,N_8822);
and UO_210 (O_210,N_9643,N_8061);
and UO_211 (O_211,N_8176,N_9850);
xnor UO_212 (O_212,N_8970,N_9892);
and UO_213 (O_213,N_8741,N_9898);
xnor UO_214 (O_214,N_8728,N_9325);
nor UO_215 (O_215,N_9635,N_8992);
nand UO_216 (O_216,N_9373,N_8817);
nor UO_217 (O_217,N_9349,N_9964);
or UO_218 (O_218,N_8131,N_9287);
and UO_219 (O_219,N_9544,N_9210);
nand UO_220 (O_220,N_8308,N_9775);
xor UO_221 (O_221,N_8634,N_8840);
xor UO_222 (O_222,N_8595,N_8653);
xor UO_223 (O_223,N_9573,N_9215);
nand UO_224 (O_224,N_8367,N_8711);
and UO_225 (O_225,N_9180,N_8027);
xnor UO_226 (O_226,N_8380,N_8232);
and UO_227 (O_227,N_8150,N_8470);
and UO_228 (O_228,N_9999,N_8632);
xor UO_229 (O_229,N_8295,N_9756);
or UO_230 (O_230,N_9253,N_8860);
xnor UO_231 (O_231,N_8624,N_8601);
nand UO_232 (O_232,N_9291,N_8413);
nor UO_233 (O_233,N_8830,N_8962);
or UO_234 (O_234,N_9271,N_8126);
and UO_235 (O_235,N_8856,N_9981);
or UO_236 (O_236,N_8261,N_8219);
nor UO_237 (O_237,N_8055,N_8326);
or UO_238 (O_238,N_9842,N_8699);
nor UO_239 (O_239,N_9697,N_9352);
xnor UO_240 (O_240,N_8538,N_9391);
and UO_241 (O_241,N_8268,N_8629);
or UO_242 (O_242,N_9266,N_8694);
or UO_243 (O_243,N_9729,N_8287);
nor UO_244 (O_244,N_8927,N_8378);
and UO_245 (O_245,N_9820,N_9485);
or UO_246 (O_246,N_9776,N_9504);
nor UO_247 (O_247,N_9232,N_9509);
nor UO_248 (O_248,N_9688,N_9769);
and UO_249 (O_249,N_8059,N_9344);
nor UO_250 (O_250,N_8855,N_8302);
or UO_251 (O_251,N_9070,N_9550);
nor UO_252 (O_252,N_8618,N_8799);
nor UO_253 (O_253,N_8545,N_9602);
or UO_254 (O_254,N_9977,N_8866);
xnor UO_255 (O_255,N_9795,N_9939);
or UO_256 (O_256,N_9919,N_9458);
nand UO_257 (O_257,N_9085,N_8846);
xnor UO_258 (O_258,N_9370,N_9567);
nand UO_259 (O_259,N_9752,N_8245);
nor UO_260 (O_260,N_8431,N_9655);
or UO_261 (O_261,N_8980,N_9951);
or UO_262 (O_262,N_8788,N_8668);
or UO_263 (O_263,N_8317,N_9846);
nor UO_264 (O_264,N_9025,N_9916);
xor UO_265 (O_265,N_8946,N_8494);
nor UO_266 (O_266,N_9115,N_9301);
or UO_267 (O_267,N_9267,N_8487);
or UO_268 (O_268,N_9320,N_9463);
nand UO_269 (O_269,N_9591,N_9720);
or UO_270 (O_270,N_9255,N_8959);
or UO_271 (O_271,N_8266,N_9815);
and UO_272 (O_272,N_9347,N_9906);
xnor UO_273 (O_273,N_9600,N_9755);
and UO_274 (O_274,N_8832,N_9943);
and UO_275 (O_275,N_9538,N_9121);
and UO_276 (O_276,N_8851,N_8523);
nor UO_277 (O_277,N_8542,N_9529);
xnor UO_278 (O_278,N_9146,N_9535);
or UO_279 (O_279,N_9759,N_8994);
nand UO_280 (O_280,N_8363,N_9734);
nor UO_281 (O_281,N_9903,N_9508);
xnor UO_282 (O_282,N_8388,N_8592);
or UO_283 (O_283,N_9623,N_9613);
nand UO_284 (O_284,N_9741,N_9847);
and UO_285 (O_285,N_8599,N_9285);
xor UO_286 (O_286,N_8031,N_8282);
and UO_287 (O_287,N_8680,N_8337);
or UO_288 (O_288,N_8267,N_8975);
and UO_289 (O_289,N_9217,N_8708);
nand UO_290 (O_290,N_8255,N_9107);
xor UO_291 (O_291,N_9521,N_9527);
or UO_292 (O_292,N_9407,N_9861);
or UO_293 (O_293,N_9541,N_8721);
nand UO_294 (O_294,N_9182,N_8765);
and UO_295 (O_295,N_8829,N_9397);
or UO_296 (O_296,N_8648,N_8299);
nand UO_297 (O_297,N_9137,N_8903);
nor UO_298 (O_298,N_9779,N_9207);
nand UO_299 (O_299,N_8336,N_9991);
or UO_300 (O_300,N_9005,N_8824);
or UO_301 (O_301,N_9162,N_9385);
or UO_302 (O_302,N_8419,N_8047);
nor UO_303 (O_303,N_8972,N_8925);
xnor UO_304 (O_304,N_8270,N_8839);
or UO_305 (O_305,N_8759,N_8474);
nand UO_306 (O_306,N_8987,N_8288);
or UO_307 (O_307,N_8110,N_9268);
and UO_308 (O_308,N_9280,N_8563);
nand UO_309 (O_309,N_9585,N_8147);
nand UO_310 (O_310,N_9645,N_9689);
nor UO_311 (O_311,N_8782,N_8165);
and UO_312 (O_312,N_8513,N_9197);
xnor UO_313 (O_313,N_8784,N_9466);
or UO_314 (O_314,N_9911,N_9930);
and UO_315 (O_315,N_9654,N_9900);
or UO_316 (O_316,N_8479,N_8166);
nand UO_317 (O_317,N_9143,N_9100);
nor UO_318 (O_318,N_8768,N_9575);
nor UO_319 (O_319,N_8557,N_8365);
nor UO_320 (O_320,N_8807,N_9805);
xor UO_321 (O_321,N_8007,N_9653);
nand UO_322 (O_322,N_8137,N_9844);
and UO_323 (O_323,N_9942,N_9599);
and UO_324 (O_324,N_9735,N_9824);
nand UO_325 (O_325,N_8087,N_8610);
and UO_326 (O_326,N_8415,N_9502);
nand UO_327 (O_327,N_8477,N_9770);
nand UO_328 (O_328,N_8395,N_8949);
nor UO_329 (O_329,N_8529,N_8213);
xnor UO_330 (O_330,N_9419,N_8802);
nor UO_331 (O_331,N_8401,N_9897);
nor UO_332 (O_332,N_9387,N_8279);
and UO_333 (O_333,N_8942,N_8064);
nand UO_334 (O_334,N_8314,N_9326);
and UO_335 (O_335,N_9219,N_9726);
and UO_336 (O_336,N_8872,N_8003);
nor UO_337 (O_337,N_8578,N_8667);
and UO_338 (O_338,N_9579,N_8238);
or UO_339 (O_339,N_9711,N_8369);
or UO_340 (O_340,N_9202,N_9321);
xor UO_341 (O_341,N_8543,N_9547);
and UO_342 (O_342,N_9435,N_9907);
nor UO_343 (O_343,N_9669,N_8981);
and UO_344 (O_344,N_8507,N_9545);
nor UO_345 (O_345,N_8685,N_8028);
nand UO_346 (O_346,N_8155,N_9418);
and UO_347 (O_347,N_8963,N_9554);
and UO_348 (O_348,N_8893,N_9838);
xor UO_349 (O_349,N_9380,N_8342);
nand UO_350 (O_350,N_9772,N_8316);
nor UO_351 (O_351,N_8319,N_8141);
or UO_352 (O_352,N_8202,N_8051);
and UO_353 (O_353,N_8052,N_8133);
nor UO_354 (O_354,N_9517,N_9961);
nand UO_355 (O_355,N_8015,N_9584);
xor UO_356 (O_356,N_8019,N_9612);
xnor UO_357 (O_357,N_9958,N_9855);
or UO_358 (O_358,N_8999,N_8530);
nand UO_359 (O_359,N_9909,N_8442);
and UO_360 (O_360,N_9514,N_8008);
or UO_361 (O_361,N_8548,N_9160);
and UO_362 (O_362,N_8000,N_9133);
nand UO_363 (O_363,N_8914,N_9873);
xor UO_364 (O_364,N_9422,N_9472);
xnor UO_365 (O_365,N_8081,N_8719);
or UO_366 (O_366,N_9284,N_8620);
nor UO_367 (O_367,N_8713,N_9638);
xnor UO_368 (O_368,N_8100,N_9715);
nand UO_369 (O_369,N_8843,N_8381);
nand UO_370 (O_370,N_8033,N_8226);
or UO_371 (O_371,N_8778,N_8552);
nor UO_372 (O_372,N_8293,N_8567);
xor UO_373 (O_373,N_8666,N_9806);
or UO_374 (O_374,N_9004,N_8844);
nor UO_375 (O_375,N_8102,N_8361);
xor UO_376 (O_376,N_9921,N_8286);
nand UO_377 (O_377,N_9191,N_9754);
or UO_378 (O_378,N_8600,N_9181);
nor UO_379 (O_379,N_8333,N_8174);
nor UO_380 (O_380,N_9698,N_8191);
or UO_381 (O_381,N_8284,N_8786);
and UO_382 (O_382,N_9302,N_8997);
nor UO_383 (O_383,N_9552,N_9470);
nand UO_384 (O_384,N_8248,N_8845);
and UO_385 (O_385,N_9350,N_8193);
nand UO_386 (O_386,N_9608,N_9106);
nor UO_387 (O_387,N_8321,N_8794);
xnor UO_388 (O_388,N_8043,N_8789);
or UO_389 (O_389,N_8383,N_8272);
and UO_390 (O_390,N_8242,N_8701);
or UO_391 (O_391,N_9125,N_9398);
xnor UO_392 (O_392,N_9343,N_9946);
nor UO_393 (O_393,N_9712,N_8376);
xnor UO_394 (O_394,N_8359,N_9925);
nand UO_395 (O_395,N_9783,N_9185);
xnor UO_396 (O_396,N_9057,N_8198);
or UO_397 (O_397,N_8793,N_9490);
or UO_398 (O_398,N_9722,N_9184);
nand UO_399 (O_399,N_8937,N_8930);
xor UO_400 (O_400,N_8684,N_9088);
nand UO_401 (O_401,N_8547,N_9129);
and UO_402 (O_402,N_8948,N_8920);
nand UO_403 (O_403,N_8430,N_8993);
nand UO_404 (O_404,N_9092,N_9934);
xor UO_405 (O_405,N_9340,N_8646);
nor UO_406 (O_406,N_8919,N_8309);
nand UO_407 (O_407,N_9956,N_9323);
xnor UO_408 (O_408,N_8041,N_9474);
and UO_409 (O_409,N_8527,N_8382);
nor UO_410 (O_410,N_8360,N_9335);
nor UO_411 (O_411,N_8188,N_8090);
nor UO_412 (O_412,N_8854,N_9721);
nor UO_413 (O_413,N_8113,N_9000);
nor UO_414 (O_414,N_8806,N_8857);
nor UO_415 (O_415,N_9764,N_9520);
and UO_416 (O_416,N_8978,N_9381);
nand UO_417 (O_417,N_9225,N_8160);
nand UO_418 (O_418,N_9630,N_9426);
nor UO_419 (O_419,N_8850,N_8899);
nand UO_420 (O_420,N_8506,N_8670);
or UO_421 (O_421,N_9199,N_8655);
xnor UO_422 (O_422,N_8825,N_8428);
and UO_423 (O_423,N_9500,N_9745);
xor UO_424 (O_424,N_9299,N_9113);
nor UO_425 (O_425,N_8142,N_9665);
and UO_426 (O_426,N_9875,N_9863);
nor UO_427 (O_427,N_8285,N_8310);
or UO_428 (O_428,N_8304,N_8275);
xnor UO_429 (O_429,N_8892,N_8416);
nand UO_430 (O_430,N_9392,N_8161);
xnor UO_431 (O_431,N_9216,N_9446);
and UO_432 (O_432,N_8108,N_8018);
or UO_433 (O_433,N_8950,N_9707);
xor UO_434 (O_434,N_9389,N_9001);
nand UO_435 (O_435,N_9173,N_8217);
and UO_436 (O_436,N_9644,N_8485);
nor UO_437 (O_437,N_9018,N_8965);
and UO_438 (O_438,N_9590,N_8810);
and UO_439 (O_439,N_8940,N_8898);
nor UO_440 (O_440,N_9839,N_8922);
xnor UO_441 (O_441,N_8092,N_8665);
nand UO_442 (O_442,N_8086,N_9791);
and UO_443 (O_443,N_8909,N_8115);
nor UO_444 (O_444,N_8344,N_9139);
or UO_445 (O_445,N_8580,N_8774);
and UO_446 (O_446,N_9566,N_8943);
xnor UO_447 (O_447,N_8350,N_9997);
nor UO_448 (O_448,N_8290,N_8358);
or UO_449 (O_449,N_8753,N_8519);
xnor UO_450 (O_450,N_8742,N_8901);
and UO_451 (O_451,N_9147,N_9696);
xnor UO_452 (O_452,N_9960,N_9523);
nand UO_453 (O_453,N_9103,N_9156);
and UO_454 (O_454,N_8303,N_9292);
nand UO_455 (O_455,N_9177,N_8054);
nand UO_456 (O_456,N_9680,N_8986);
and UO_457 (O_457,N_8044,N_8868);
and UO_458 (O_458,N_8254,N_8005);
and UO_459 (O_459,N_8178,N_9837);
or UO_460 (O_460,N_9275,N_9098);
nor UO_461 (O_461,N_9231,N_9395);
nand UO_462 (O_462,N_9062,N_9799);
xor UO_463 (O_463,N_9857,N_9158);
or UO_464 (O_464,N_8002,N_9249);
and UO_465 (O_465,N_9796,N_9672);
xor UO_466 (O_466,N_9917,N_9658);
nand UO_467 (O_467,N_8770,N_8156);
nor UO_468 (O_468,N_9127,N_8691);
xor UO_469 (O_469,N_9401,N_8627);
nor UO_470 (O_470,N_9940,N_9642);
xnor UO_471 (O_471,N_9577,N_9498);
xnor UO_472 (O_472,N_9084,N_9578);
xnor UO_473 (O_473,N_9760,N_8945);
nand UO_474 (O_474,N_9065,N_9341);
or UO_475 (O_475,N_8748,N_9763);
and UO_476 (O_476,N_8123,N_8546);
xor UO_477 (O_477,N_8257,N_8515);
or UO_478 (O_478,N_8185,N_8503);
and UO_479 (O_479,N_9338,N_9982);
xnor UO_480 (O_480,N_8813,N_8262);
and UO_481 (O_481,N_9915,N_8247);
or UO_482 (O_482,N_9124,N_9020);
and UO_483 (O_483,N_9445,N_9626);
or UO_484 (O_484,N_9950,N_8453);
nor UO_485 (O_485,N_9973,N_8076);
nor UO_486 (O_486,N_9920,N_9414);
xor UO_487 (O_487,N_9883,N_9918);
or UO_488 (O_488,N_9657,N_8071);
nand UO_489 (O_489,N_9108,N_8715);
nor UO_490 (O_490,N_9895,N_9167);
nand UO_491 (O_491,N_9831,N_8264);
and UO_492 (O_492,N_8392,N_8389);
and UO_493 (O_493,N_9072,N_9024);
or UO_494 (O_494,N_8038,N_8852);
nand UO_495 (O_495,N_8386,N_8399);
and UO_496 (O_496,N_8096,N_8731);
nand UO_497 (O_497,N_8049,N_9914);
and UO_498 (O_498,N_9442,N_9487);
and UO_499 (O_499,N_8502,N_9988);
and UO_500 (O_500,N_8677,N_8835);
xor UO_501 (O_501,N_8977,N_9297);
xnor UO_502 (O_502,N_9986,N_8283);
xnor UO_503 (O_503,N_8124,N_9639);
or UO_504 (O_504,N_9492,N_8404);
or UO_505 (O_505,N_8692,N_9571);
nand UO_506 (O_506,N_9596,N_8201);
nor UO_507 (O_507,N_8486,N_9496);
xnor UO_508 (O_508,N_8785,N_9843);
xnor UO_509 (O_509,N_9902,N_8769);
nor UO_510 (O_510,N_8117,N_9877);
nand UO_511 (O_511,N_9186,N_8410);
or UO_512 (O_512,N_8564,N_8060);
nand UO_513 (O_513,N_8512,N_9968);
nor UO_514 (O_514,N_9966,N_8956);
nor UO_515 (O_515,N_9736,N_9307);
or UO_516 (O_516,N_9166,N_8885);
and UO_517 (O_517,N_9823,N_8405);
nor UO_518 (O_518,N_9239,N_9827);
xnor UO_519 (O_519,N_8216,N_8882);
and UO_520 (O_520,N_9324,N_8127);
or UO_521 (O_521,N_9812,N_9064);
and UO_522 (O_522,N_8037,N_9773);
xor UO_523 (O_523,N_8705,N_9094);
nor UO_524 (O_524,N_8444,N_8833);
nand UO_525 (O_525,N_8085,N_9701);
xor UO_526 (O_526,N_9924,N_8849);
xor UO_527 (O_527,N_9204,N_9574);
nand UO_528 (O_528,N_8658,N_9454);
xnor UO_529 (O_529,N_9037,N_9762);
xnor UO_530 (O_530,N_9176,N_9198);
and UO_531 (O_531,N_8803,N_8281);
or UO_532 (O_532,N_8697,N_9728);
nand UO_533 (O_533,N_8775,N_8853);
or UO_534 (O_534,N_8289,N_9730);
nand UO_535 (O_535,N_9743,N_8911);
and UO_536 (O_536,N_8717,N_8744);
or UO_537 (O_537,N_9432,N_9264);
nor UO_538 (O_538,N_9536,N_9652);
and UO_539 (O_539,N_8565,N_8101);
xor UO_540 (O_540,N_8074,N_8531);
and UO_541 (O_541,N_9434,N_9039);
nand UO_542 (O_542,N_9293,N_8229);
or UO_543 (O_543,N_8374,N_9714);
nand UO_544 (O_544,N_9935,N_8056);
and UO_545 (O_545,N_9371,N_8664);
or UO_546 (O_546,N_9822,N_9800);
nor UO_547 (O_547,N_8902,N_8422);
nor UO_548 (O_548,N_8689,N_8528);
and UO_549 (O_549,N_9963,N_8710);
nand UO_550 (O_550,N_8831,N_8740);
or UO_551 (O_551,N_8190,N_9647);
nand UO_552 (O_552,N_9366,N_9719);
or UO_553 (O_553,N_8203,N_9505);
xor UO_554 (O_554,N_9798,N_8894);
or UO_555 (O_555,N_8417,N_9817);
xor UO_556 (O_556,N_9351,N_8504);
xnor UO_557 (O_557,N_9931,N_8616);
or UO_558 (O_558,N_9890,N_8205);
nand UO_559 (O_559,N_9724,N_8463);
xnor UO_560 (O_560,N_8724,N_9611);
and UO_561 (O_561,N_8555,N_8186);
nor UO_562 (O_562,N_8661,N_9482);
or UO_563 (O_563,N_9304,N_8619);
nor UO_564 (O_564,N_9661,N_8406);
nand UO_565 (O_565,N_8676,N_9168);
and UO_566 (O_566,N_9229,N_8116);
xor UO_567 (O_567,N_8209,N_9932);
nand UO_568 (O_568,N_8091,N_8162);
nand UO_569 (O_569,N_8200,N_9609);
or UO_570 (O_570,N_8473,N_9415);
nand UO_571 (O_571,N_9040,N_9461);
xor UO_572 (O_572,N_9947,N_9702);
and UO_573 (O_573,N_9455,N_9851);
nand UO_574 (O_574,N_8873,N_8004);
nand UO_575 (O_575,N_8251,N_8584);
or UO_576 (O_576,N_8912,N_8335);
nor UO_577 (O_577,N_9079,N_9927);
or UO_578 (O_578,N_9819,N_8153);
and UO_579 (O_579,N_9265,N_8910);
and UO_580 (O_580,N_9962,N_8760);
or UO_581 (O_581,N_8212,N_8181);
xor UO_582 (O_582,N_8347,N_8320);
and UO_583 (O_583,N_8883,N_9739);
nor UO_584 (O_584,N_8521,N_8077);
nand UO_585 (O_585,N_9501,N_8612);
nor UO_586 (O_586,N_9990,N_8396);
and UO_587 (O_587,N_9258,N_9375);
nor UO_588 (O_588,N_8888,N_9929);
xor UO_589 (O_589,N_8109,N_9393);
and UO_590 (O_590,N_9690,N_9616);
xor UO_591 (O_591,N_8630,N_8998);
or UO_592 (O_592,N_9674,N_8798);
xor UO_593 (O_593,N_9888,N_8797);
or UO_594 (O_594,N_9840,N_9695);
and UO_595 (O_595,N_8941,N_9849);
or UO_596 (O_596,N_9041,N_9236);
and UO_597 (O_597,N_8602,N_9926);
nand UO_598 (O_598,N_8134,N_9938);
xor UO_599 (O_599,N_8034,N_8621);
nor UO_600 (O_600,N_8570,N_9975);
nand UO_601 (O_601,N_8952,N_8989);
xnor UO_602 (O_602,N_9807,N_8650);
and UO_603 (O_603,N_9518,N_9283);
and UO_604 (O_604,N_8098,N_8020);
and UO_605 (O_605,N_8642,N_9195);
xnor UO_606 (O_606,N_8447,N_8674);
xnor UO_607 (O_607,N_8541,N_8756);
or UO_608 (O_608,N_8346,N_9082);
and UO_609 (O_609,N_9936,N_9369);
nor UO_610 (O_610,N_9478,N_8328);
and UO_611 (O_611,N_8735,N_9174);
or UO_612 (O_612,N_8039,N_8576);
or UO_613 (O_613,N_8391,N_9148);
nor UO_614 (O_614,N_9131,N_9751);
nand UO_615 (O_615,N_9433,N_9221);
nor UO_616 (O_616,N_9102,N_9399);
nand UO_617 (O_617,N_9663,N_8221);
and UO_618 (O_618,N_9354,N_9705);
or UO_619 (O_619,N_9937,N_9580);
nor UO_620 (O_620,N_8837,N_8522);
nand UO_621 (O_621,N_9640,N_8847);
or UO_622 (O_622,N_9112,N_9119);
nor UO_623 (O_623,N_8826,N_8218);
nor UO_624 (O_624,N_9747,N_8561);
xnor UO_625 (O_625,N_9476,N_8652);
or UO_626 (O_626,N_9410,N_8111);
xnor UO_627 (O_627,N_9059,N_8149);
nor UO_628 (O_628,N_9531,N_8559);
nor UO_629 (O_629,N_9416,N_9488);
nand UO_630 (O_630,N_8819,N_9785);
xnor UO_631 (O_631,N_9300,N_8660);
or UO_632 (O_632,N_9830,N_8779);
xnor UO_633 (O_633,N_9170,N_9540);
nor UO_634 (O_634,N_8408,N_9475);
or UO_635 (O_635,N_8106,N_9440);
and UO_636 (O_636,N_9601,N_9787);
or UO_637 (O_637,N_9096,N_9172);
xnor UO_638 (O_638,N_8046,N_8439);
or UO_639 (O_639,N_8679,N_9671);
xnor UO_640 (O_640,N_8152,N_9503);
and UO_641 (O_641,N_8571,N_8050);
xnor UO_642 (O_642,N_8143,N_9627);
nand UO_643 (O_643,N_8146,N_9788);
xnor UO_644 (O_644,N_9526,N_8907);
xnor UO_645 (O_645,N_9122,N_9144);
xor UO_646 (O_646,N_8418,N_8329);
nor UO_647 (O_647,N_9318,N_9588);
nand UO_648 (O_648,N_9192,N_9342);
xor UO_649 (O_649,N_9564,N_8968);
or UO_650 (O_650,N_9086,N_9899);
nand UO_651 (O_651,N_9945,N_9867);
nor UO_652 (O_652,N_8011,N_9404);
nand UO_653 (O_653,N_9016,N_8118);
xnor UO_654 (O_654,N_8476,N_8490);
nand UO_655 (O_655,N_9406,N_8645);
or UO_656 (O_656,N_9068,N_9425);
nor UO_657 (O_657,N_9553,N_9651);
nand UO_658 (O_658,N_8088,N_9771);
xnor UO_659 (O_659,N_9153,N_8112);
nor UO_660 (O_660,N_9042,N_9390);
and UO_661 (O_661,N_9049,N_8918);
nor UO_662 (O_662,N_9572,N_9196);
or UO_663 (O_663,N_9150,N_8398);
and UO_664 (O_664,N_9511,N_9871);
and UO_665 (O_665,N_8771,N_9742);
and UO_666 (O_666,N_8508,N_8349);
nand UO_667 (O_667,N_9949,N_8097);
or UO_668 (O_668,N_9473,N_9864);
nand UO_669 (O_669,N_8733,N_9622);
nand UO_670 (O_670,N_9048,N_9256);
nor UO_671 (O_671,N_9159,N_8443);
xor UO_672 (O_672,N_9078,N_9922);
xor UO_673 (O_673,N_9314,N_8876);
or UO_674 (O_674,N_9675,N_9439);
and UO_675 (O_675,N_9528,N_8752);
and UO_676 (O_676,N_9200,N_8585);
nor UO_677 (O_677,N_8500,N_8574);
or UO_678 (O_678,N_8820,N_9120);
nand UO_679 (O_679,N_8370,N_8180);
or UO_680 (O_680,N_8656,N_9479);
or UO_681 (O_681,N_9286,N_9814);
and UO_682 (O_682,N_8662,N_9189);
or UO_683 (O_683,N_9621,N_9394);
nand UO_684 (O_684,N_9289,N_9826);
nand UO_685 (O_685,N_9984,N_9362);
or UO_686 (O_686,N_9683,N_9569);
nor UO_687 (O_687,N_9969,N_9209);
or UO_688 (O_688,N_8594,N_8471);
nand UO_689 (O_689,N_8057,N_9227);
nand UO_690 (O_690,N_8591,N_9203);
or UO_691 (O_691,N_8623,N_9813);
nor UO_692 (O_692,N_9154,N_9853);
nand UO_693 (O_693,N_9668,N_8225);
nand UO_694 (O_694,N_8886,N_8079);
xnor UO_695 (O_695,N_9811,N_8276);
xor UO_696 (O_696,N_8534,N_8236);
and UO_697 (O_697,N_9111,N_8259);
nand UO_698 (O_698,N_8514,N_9034);
nand UO_699 (O_699,N_8633,N_9077);
or UO_700 (O_700,N_9261,N_8672);
or UO_701 (O_701,N_8532,N_9678);
or UO_702 (O_702,N_9141,N_8597);
and UO_703 (O_703,N_9510,N_9151);
and UO_704 (O_704,N_9858,N_9053);
or UO_705 (O_705,N_8870,N_8129);
nand UO_706 (O_706,N_8394,N_8809);
nor UO_707 (O_707,N_9834,N_8772);
nand UO_708 (O_708,N_8021,N_8063);
or UO_709 (O_709,N_9793,N_9254);
nand UO_710 (O_710,N_9364,N_9087);
and UO_711 (O_711,N_9142,N_9110);
and UO_712 (O_712,N_8540,N_8014);
nand UO_713 (O_713,N_8590,N_9562);
or UO_714 (O_714,N_8488,N_9308);
and UO_715 (O_715,N_9328,N_8122);
or UO_716 (O_716,N_8460,N_9684);
and UO_717 (O_717,N_9363,N_9624);
nor UO_718 (O_718,N_8187,N_9319);
or UO_719 (O_719,N_8001,N_9130);
nor UO_720 (O_720,N_8743,N_8904);
nand UO_721 (O_721,N_9522,N_8235);
or UO_722 (O_722,N_8368,N_9060);
and UO_723 (O_723,N_9625,N_9372);
xor UO_724 (O_724,N_8461,N_8189);
or UO_725 (O_725,N_8211,N_8318);
nor UO_726 (O_726,N_8084,N_9905);
or UO_727 (O_727,N_9856,N_9894);
or UO_728 (O_728,N_8891,N_8353);
xnor UO_729 (O_729,N_8469,N_8884);
and UO_730 (O_730,N_8566,N_8432);
nor UO_731 (O_731,N_8271,N_8331);
nand UO_732 (O_732,N_8467,N_8073);
and UO_733 (O_733,N_9277,N_8654);
nand UO_734 (O_734,N_8875,N_8440);
or UO_735 (O_735,N_8214,N_8974);
nand UO_736 (O_736,N_8372,N_9309);
nand UO_737 (O_737,N_9533,N_9290);
and UO_738 (O_738,N_9928,N_8815);
or UO_739 (O_739,N_9879,N_8625);
and UO_740 (O_740,N_8220,N_9818);
xnor UO_741 (O_741,N_9413,N_9294);
nand UO_742 (O_742,N_9480,N_9749);
nand UO_743 (O_743,N_9157,N_9828);
and UO_744 (O_744,N_8982,N_9134);
nor UO_745 (O_745,N_8114,N_8737);
and UO_746 (O_746,N_9633,N_9023);
nand UO_747 (O_747,N_8224,N_9105);
and UO_748 (O_748,N_8325,N_9704);
xnor UO_749 (O_749,N_8312,N_9032);
or UO_750 (O_750,N_8313,N_8553);
and UO_751 (O_751,N_8889,N_9589);
nand UO_752 (O_752,N_8944,N_9444);
nand UO_753 (O_753,N_9832,N_8572);
nand UO_754 (O_754,N_8256,N_9563);
xnor UO_755 (O_755,N_8010,N_8083);
and UO_756 (O_756,N_9233,N_9441);
xor UO_757 (O_757,N_9081,N_8455);
nand UO_758 (O_758,N_8194,N_9008);
xnor UO_759 (O_759,N_8138,N_9447);
nand UO_760 (O_760,N_8767,N_9524);
or UO_761 (O_761,N_9666,N_8107);
xor UO_762 (O_762,N_8323,N_8426);
nand UO_763 (O_763,N_9190,N_8577);
or UO_764 (O_764,N_9604,N_8269);
or UO_765 (O_765,N_8121,N_8841);
nor UO_766 (O_766,N_9178,N_8967);
xnor UO_767 (O_767,N_9881,N_8906);
xor UO_768 (O_768,N_8163,N_8971);
nand UO_769 (O_769,N_8641,N_9274);
or UO_770 (O_770,N_8781,N_8976);
or UO_771 (O_771,N_9717,N_9421);
or UO_772 (O_772,N_8029,N_8450);
and UO_773 (O_773,N_8068,N_8481);
nor UO_774 (O_774,N_9259,N_9408);
nor UO_775 (O_775,N_9901,N_8509);
and UO_776 (O_776,N_8009,N_8491);
and UO_777 (O_777,N_9009,N_8136);
nor UO_778 (O_778,N_9617,N_9794);
nand UO_779 (O_779,N_8462,N_8526);
xnor UO_780 (O_780,N_8154,N_9090);
nor UO_781 (O_781,N_8720,N_8678);
or UO_782 (O_782,N_8926,N_8179);
or UO_783 (O_783,N_8878,N_8979);
xnor UO_784 (O_784,N_9055,N_8222);
nor UO_785 (O_785,N_9453,N_9218);
or UO_786 (O_786,N_8960,N_9761);
xor UO_787 (O_787,N_8628,N_9033);
and UO_788 (O_788,N_9021,N_9691);
xor UO_789 (O_789,N_9222,N_8407);
nand UO_790 (O_790,N_9636,N_9095);
nor UO_791 (O_791,N_8924,N_8792);
nand UO_792 (O_792,N_8928,N_9097);
xor UO_793 (O_793,N_9118,N_9430);
xor UO_794 (O_794,N_8749,N_8638);
nand UO_795 (O_795,N_8550,N_9506);
nor UO_796 (O_796,N_8148,N_8961);
nand UO_797 (O_797,N_8249,N_8280);
and UO_798 (O_798,N_8890,N_8958);
and UO_799 (O_799,N_9428,N_9737);
and UO_800 (O_800,N_8042,N_9629);
or UO_801 (O_801,N_9194,N_9379);
xnor UO_802 (O_802,N_8158,N_8758);
or UO_803 (O_803,N_9211,N_9637);
nand UO_804 (O_804,N_9051,N_8482);
xnor UO_805 (O_805,N_9359,N_9330);
nor UO_806 (O_806,N_8611,N_8035);
nor UO_807 (O_807,N_8750,N_9311);
and UO_808 (O_808,N_8808,N_8659);
nor UO_809 (O_809,N_9052,N_8709);
nand UO_810 (O_810,N_9183,N_8233);
xnor UO_811 (O_811,N_9836,N_8048);
nor UO_812 (O_812,N_9885,N_8505);
xor UO_813 (O_813,N_8501,N_9782);
nand UO_814 (O_814,N_9664,N_8562);
nor UO_815 (O_815,N_8921,N_8448);
and UO_816 (O_816,N_9594,N_9188);
or UO_817 (O_817,N_8688,N_8258);
or UO_818 (O_818,N_9091,N_9954);
nor UO_819 (O_819,N_9555,N_9913);
xor UO_820 (O_820,N_9841,N_9628);
or UO_821 (O_821,N_9089,N_8695);
and UO_822 (O_822,N_8864,N_8298);
or UO_823 (O_823,N_9242,N_9641);
and UO_824 (O_824,N_9568,N_9592);
xnor UO_825 (O_825,N_8480,N_8985);
xor UO_826 (O_826,N_8170,N_9662);
or UO_827 (O_827,N_8466,N_9224);
nand UO_828 (O_828,N_8397,N_9450);
and UO_829 (O_829,N_8240,N_9424);
or UO_830 (O_830,N_9101,N_9228);
and UO_831 (O_831,N_9030,N_9619);
nand UO_832 (O_832,N_9803,N_9748);
nor UO_833 (O_833,N_8823,N_9821);
or UO_834 (O_834,N_9050,N_9031);
or UO_835 (O_835,N_9989,N_9532);
or UO_836 (O_836,N_8080,N_9288);
nor UO_837 (O_837,N_9235,N_8556);
xor UO_838 (O_838,N_8130,N_9558);
and UO_839 (O_839,N_9035,N_9003);
nor UO_840 (O_840,N_8896,N_9833);
xnor UO_841 (O_841,N_9992,N_9797);
xnor UO_842 (O_842,N_9043,N_8716);
or UO_843 (O_843,N_8626,N_9586);
xor UO_844 (O_844,N_9276,N_8858);
nor UO_845 (O_845,N_9402,N_9109);
or UO_846 (O_846,N_9516,N_9699);
xnor UO_847 (O_847,N_9484,N_9456);
and UO_848 (O_848,N_8703,N_8175);
or UO_849 (O_849,N_8747,N_9348);
nand UO_850 (O_850,N_9872,N_9316);
and UO_851 (O_851,N_8006,N_9412);
xnor UO_852 (O_852,N_9334,N_9214);
or UO_853 (O_853,N_9015,N_8167);
or UO_854 (O_854,N_8139,N_8693);
or UO_855 (O_855,N_9618,N_9240);
nor UO_856 (O_856,N_8544,N_9694);
nor UO_857 (O_857,N_9367,N_8588);
or UO_858 (O_858,N_8915,N_8726);
and UO_859 (O_859,N_9801,N_9477);
xnor UO_860 (O_860,N_8412,N_9278);
nor UO_861 (O_861,N_9123,N_8420);
xor UO_862 (O_862,N_9282,N_8377);
nor UO_863 (O_863,N_8734,N_8812);
and UO_864 (O_864,N_8296,N_8745);
or UO_865 (O_865,N_9993,N_9953);
and UO_866 (O_866,N_9244,N_9467);
xor UO_867 (O_867,N_8673,N_8263);
and UO_868 (O_868,N_9459,N_9427);
nand UO_869 (O_869,N_8936,N_9438);
or UO_870 (O_870,N_8933,N_8135);
nor UO_871 (O_871,N_9732,N_8657);
nor UO_872 (O_872,N_9272,N_9816);
nor UO_873 (O_873,N_9904,N_9358);
xnor UO_874 (O_874,N_9312,N_9464);
nor UO_875 (O_875,N_8492,N_9632);
or UO_876 (O_876,N_9667,N_9559);
xnor UO_877 (O_877,N_8103,N_8025);
xnor UO_878 (O_878,N_9998,N_9388);
or UO_879 (O_879,N_8082,N_8932);
nand UO_880 (O_880,N_8468,N_9383);
xor UO_881 (O_881,N_9952,N_8437);
nor UO_882 (O_882,N_9866,N_8706);
nor UO_883 (O_883,N_9767,N_8493);
xor UO_884 (O_884,N_8330,N_8895);
nor UO_885 (O_885,N_9193,N_8923);
or UO_886 (O_886,N_9650,N_8983);
nand UO_887 (O_887,N_9073,N_8687);
xor UO_888 (O_888,N_8931,N_9409);
xor UO_889 (O_889,N_9457,N_9519);
nor UO_890 (O_890,N_8520,N_8339);
and UO_891 (O_891,N_8533,N_9336);
nand UO_892 (O_892,N_9659,N_8917);
xnor UO_893 (O_893,N_9507,N_8751);
nor UO_894 (O_894,N_9136,N_8105);
nor UO_895 (O_895,N_8030,N_9537);
and UO_896 (O_896,N_8636,N_8877);
or UO_897 (O_897,N_9080,N_8053);
nor UO_898 (O_898,N_8355,N_9576);
xnor UO_899 (O_899,N_8294,N_9248);
and UO_900 (O_900,N_8879,N_8246);
or UO_901 (O_901,N_9315,N_8429);
and UO_902 (O_902,N_9884,N_9145);
and UO_903 (O_903,N_8184,N_8723);
nand UO_904 (O_904,N_9774,N_8579);
or UO_905 (O_905,N_9994,N_9099);
nand UO_906 (O_906,N_8575,N_9865);
xnor UO_907 (O_907,N_8207,N_9436);
and UO_908 (O_908,N_9710,N_9565);
nand UO_909 (O_909,N_8603,N_9557);
or UO_910 (O_910,N_9607,N_9860);
xnor UO_911 (O_911,N_9810,N_8375);
nand UO_912 (O_912,N_8838,N_9298);
xnor UO_913 (O_913,N_9384,N_8637);
xor UO_914 (O_914,N_8393,N_8495);
and UO_915 (O_915,N_8549,N_8017);
nand UO_916 (O_916,N_8780,N_9784);
xnor UO_917 (O_917,N_8250,N_9269);
nand UO_918 (O_918,N_9548,N_9738);
nand UO_919 (O_919,N_8168,N_9753);
xor UO_920 (O_920,N_9489,N_9987);
or UO_921 (O_921,N_9169,N_9766);
nor UO_922 (O_922,N_9530,N_8446);
and UO_923 (O_923,N_9731,N_9525);
or UO_924 (O_924,N_8551,N_8725);
nand UO_925 (O_925,N_9310,N_9845);
or UO_926 (O_926,N_8881,N_8777);
and UO_927 (O_927,N_9353,N_9681);
and UO_928 (O_928,N_9206,N_9648);
and UO_929 (O_929,N_8424,N_8069);
or UO_930 (O_930,N_9727,N_8966);
nand UO_931 (O_931,N_9598,N_9620);
or UO_932 (O_932,N_8307,N_8016);
xor UO_933 (O_933,N_8483,N_9493);
nand UO_934 (O_934,N_8305,N_8199);
nor UO_935 (O_935,N_9405,N_9243);
nor UO_936 (O_936,N_9443,N_8354);
and UO_937 (O_937,N_9854,N_9549);
nand UO_938 (O_938,N_9223,N_8145);
nor UO_939 (O_939,N_8454,N_9605);
nand UO_940 (O_940,N_9333,N_9941);
xnor UO_941 (O_941,N_8681,N_8414);
or UO_942 (O_942,N_8990,N_9923);
nor UO_943 (O_943,N_9777,N_9465);
xnor UO_944 (O_944,N_9723,N_9083);
nor UO_945 (O_945,N_8499,N_8197);
nor UO_946 (O_946,N_9006,N_9497);
nor UO_947 (O_947,N_8938,N_8766);
nand UO_948 (O_948,N_8704,N_8996);
and UO_949 (O_949,N_8458,N_8013);
or UO_950 (O_950,N_8605,N_9429);
xnor UO_951 (O_951,N_8297,N_9758);
nor UO_952 (O_952,N_8524,N_9104);
nor UO_953 (O_953,N_8045,N_9171);
or UO_954 (O_954,N_8821,N_9220);
nand UO_955 (O_955,N_9054,N_8818);
nand UO_956 (O_956,N_9246,N_8265);
and UO_957 (O_957,N_9346,N_9075);
xnor UO_958 (O_958,N_9874,N_9449);
and UO_959 (O_959,N_8539,N_8773);
nand UO_960 (O_960,N_8586,N_9026);
or UO_961 (O_961,N_9155,N_8237);
nand UO_962 (O_962,N_8334,N_8880);
and UO_963 (O_963,N_9076,N_9677);
nand UO_964 (O_964,N_9010,N_8159);
xor UO_965 (O_965,N_8763,N_9693);
and UO_966 (O_966,N_9058,N_8865);
or UO_967 (O_967,N_9891,N_8459);
and UO_968 (O_968,N_8489,N_9706);
or UO_969 (O_969,N_9128,N_9377);
and UO_970 (O_970,N_8332,N_8811);
nor UO_971 (O_971,N_8451,N_8776);
and UO_972 (O_972,N_9296,N_8498);
and UO_973 (O_973,N_8252,N_8631);
xnor UO_974 (O_974,N_9022,N_9386);
and UO_975 (O_975,N_8040,N_9132);
and UO_976 (O_976,N_8435,N_9069);
and UO_977 (O_977,N_9471,N_8182);
xnor UO_978 (O_978,N_8929,N_8125);
nand UO_979 (O_979,N_9513,N_8686);
or UO_980 (O_980,N_8241,N_9491);
nor UO_981 (O_981,N_8964,N_8387);
nand UO_982 (O_982,N_8385,N_9431);
nand UO_983 (O_983,N_9765,N_9149);
nor UO_984 (O_984,N_8239,N_8095);
xnor UO_985 (O_985,N_9996,N_8157);
nand UO_986 (O_986,N_8273,N_8078);
xnor UO_987 (O_987,N_9933,N_9908);
or UO_988 (O_988,N_8861,N_8608);
xnor UO_989 (O_989,N_8791,N_8151);
nand UO_990 (O_990,N_8690,N_9848);
and UO_991 (O_991,N_8871,N_8596);
nor UO_992 (O_992,N_8954,N_8718);
and UO_993 (O_993,N_9260,N_8900);
nand UO_994 (O_994,N_9896,N_9673);
or UO_995 (O_995,N_9595,N_9985);
or UO_996 (O_996,N_9273,N_8022);
and UO_997 (O_997,N_9317,N_9740);
xor UO_998 (O_998,N_9546,N_8707);
or UO_999 (O_999,N_8026,N_8433);
and UO_1000 (O_1000,N_9311,N_8754);
nor UO_1001 (O_1001,N_9155,N_9966);
nand UO_1002 (O_1002,N_8315,N_8337);
nand UO_1003 (O_1003,N_8575,N_8357);
nor UO_1004 (O_1004,N_8837,N_9349);
and UO_1005 (O_1005,N_8744,N_8840);
or UO_1006 (O_1006,N_8908,N_8228);
nand UO_1007 (O_1007,N_9998,N_8553);
nand UO_1008 (O_1008,N_8553,N_9184);
xor UO_1009 (O_1009,N_8464,N_9448);
and UO_1010 (O_1010,N_8646,N_9476);
and UO_1011 (O_1011,N_8359,N_9442);
xnor UO_1012 (O_1012,N_8931,N_8842);
nor UO_1013 (O_1013,N_8836,N_9556);
nand UO_1014 (O_1014,N_9788,N_8859);
xor UO_1015 (O_1015,N_8454,N_9813);
nand UO_1016 (O_1016,N_8614,N_9814);
nand UO_1017 (O_1017,N_8801,N_9290);
nor UO_1018 (O_1018,N_9771,N_8454);
or UO_1019 (O_1019,N_9129,N_9213);
nor UO_1020 (O_1020,N_9337,N_9739);
or UO_1021 (O_1021,N_9563,N_8016);
and UO_1022 (O_1022,N_8407,N_8071);
xor UO_1023 (O_1023,N_9373,N_9187);
nand UO_1024 (O_1024,N_9859,N_8353);
xor UO_1025 (O_1025,N_9098,N_8524);
xnor UO_1026 (O_1026,N_8894,N_9981);
nor UO_1027 (O_1027,N_8100,N_8564);
or UO_1028 (O_1028,N_9787,N_8028);
nor UO_1029 (O_1029,N_8356,N_9878);
xnor UO_1030 (O_1030,N_8245,N_9994);
and UO_1031 (O_1031,N_9029,N_9978);
xor UO_1032 (O_1032,N_9990,N_8886);
nor UO_1033 (O_1033,N_8860,N_8410);
and UO_1034 (O_1034,N_9347,N_8207);
or UO_1035 (O_1035,N_8525,N_8188);
nand UO_1036 (O_1036,N_8182,N_9997);
and UO_1037 (O_1037,N_9272,N_8598);
xor UO_1038 (O_1038,N_9587,N_9296);
and UO_1039 (O_1039,N_8003,N_8095);
or UO_1040 (O_1040,N_8563,N_9984);
xnor UO_1041 (O_1041,N_9917,N_8317);
nand UO_1042 (O_1042,N_9798,N_9829);
nor UO_1043 (O_1043,N_9924,N_9910);
nor UO_1044 (O_1044,N_9212,N_8438);
xor UO_1045 (O_1045,N_8946,N_9375);
or UO_1046 (O_1046,N_9427,N_9486);
and UO_1047 (O_1047,N_8890,N_8512);
and UO_1048 (O_1048,N_9976,N_8181);
nor UO_1049 (O_1049,N_8779,N_8275);
nor UO_1050 (O_1050,N_9177,N_8350);
and UO_1051 (O_1051,N_8723,N_8946);
or UO_1052 (O_1052,N_9965,N_9649);
or UO_1053 (O_1053,N_8387,N_8646);
xor UO_1054 (O_1054,N_8116,N_9834);
xor UO_1055 (O_1055,N_8101,N_8882);
or UO_1056 (O_1056,N_8968,N_9043);
xnor UO_1057 (O_1057,N_8409,N_8298);
and UO_1058 (O_1058,N_9585,N_9301);
or UO_1059 (O_1059,N_8422,N_8861);
xor UO_1060 (O_1060,N_9257,N_8170);
and UO_1061 (O_1061,N_8230,N_8388);
nand UO_1062 (O_1062,N_9585,N_9253);
nand UO_1063 (O_1063,N_8720,N_8776);
nor UO_1064 (O_1064,N_8021,N_8414);
nand UO_1065 (O_1065,N_9751,N_9560);
nand UO_1066 (O_1066,N_8286,N_8811);
or UO_1067 (O_1067,N_9222,N_9072);
or UO_1068 (O_1068,N_9244,N_9405);
and UO_1069 (O_1069,N_8183,N_9958);
nand UO_1070 (O_1070,N_8682,N_8229);
nand UO_1071 (O_1071,N_8283,N_9932);
or UO_1072 (O_1072,N_9114,N_8929);
or UO_1073 (O_1073,N_9260,N_8686);
nor UO_1074 (O_1074,N_9905,N_8918);
nand UO_1075 (O_1075,N_9405,N_9610);
nand UO_1076 (O_1076,N_9621,N_9327);
xnor UO_1077 (O_1077,N_8704,N_8810);
nand UO_1078 (O_1078,N_8665,N_8361);
nand UO_1079 (O_1079,N_9343,N_9439);
and UO_1080 (O_1080,N_9178,N_9853);
nor UO_1081 (O_1081,N_9926,N_9828);
or UO_1082 (O_1082,N_9679,N_9172);
nand UO_1083 (O_1083,N_9512,N_8944);
and UO_1084 (O_1084,N_8156,N_9431);
and UO_1085 (O_1085,N_9949,N_9641);
nor UO_1086 (O_1086,N_9850,N_9067);
nor UO_1087 (O_1087,N_8085,N_8589);
nor UO_1088 (O_1088,N_8280,N_9148);
and UO_1089 (O_1089,N_9119,N_9976);
or UO_1090 (O_1090,N_8706,N_9007);
nand UO_1091 (O_1091,N_8540,N_8028);
or UO_1092 (O_1092,N_9095,N_9989);
nand UO_1093 (O_1093,N_8504,N_9315);
nand UO_1094 (O_1094,N_9167,N_9611);
nand UO_1095 (O_1095,N_8632,N_8111);
and UO_1096 (O_1096,N_8427,N_9349);
nor UO_1097 (O_1097,N_9400,N_8904);
xor UO_1098 (O_1098,N_8467,N_9462);
xor UO_1099 (O_1099,N_9639,N_9689);
xnor UO_1100 (O_1100,N_8329,N_9792);
nor UO_1101 (O_1101,N_8509,N_8090);
nor UO_1102 (O_1102,N_8893,N_8425);
nand UO_1103 (O_1103,N_8797,N_8985);
and UO_1104 (O_1104,N_8218,N_8201);
xnor UO_1105 (O_1105,N_8578,N_9917);
and UO_1106 (O_1106,N_9510,N_9026);
nand UO_1107 (O_1107,N_9765,N_8285);
and UO_1108 (O_1108,N_9311,N_8293);
xor UO_1109 (O_1109,N_8270,N_9077);
and UO_1110 (O_1110,N_9655,N_9182);
or UO_1111 (O_1111,N_8268,N_9115);
or UO_1112 (O_1112,N_9731,N_9076);
xor UO_1113 (O_1113,N_9910,N_8242);
and UO_1114 (O_1114,N_8282,N_9114);
and UO_1115 (O_1115,N_9692,N_8669);
and UO_1116 (O_1116,N_9862,N_9988);
and UO_1117 (O_1117,N_8478,N_8479);
nand UO_1118 (O_1118,N_8785,N_9886);
and UO_1119 (O_1119,N_8440,N_9278);
xnor UO_1120 (O_1120,N_9738,N_9455);
xnor UO_1121 (O_1121,N_9464,N_9809);
or UO_1122 (O_1122,N_9424,N_8580);
nor UO_1123 (O_1123,N_8674,N_9225);
nor UO_1124 (O_1124,N_8261,N_8028);
xnor UO_1125 (O_1125,N_9807,N_9895);
nor UO_1126 (O_1126,N_9580,N_8387);
xor UO_1127 (O_1127,N_9030,N_9303);
nand UO_1128 (O_1128,N_9063,N_8918);
nor UO_1129 (O_1129,N_8606,N_9065);
xnor UO_1130 (O_1130,N_9026,N_9793);
xor UO_1131 (O_1131,N_8539,N_8152);
or UO_1132 (O_1132,N_8401,N_8986);
nand UO_1133 (O_1133,N_9335,N_8815);
and UO_1134 (O_1134,N_8425,N_9570);
nand UO_1135 (O_1135,N_9973,N_9621);
or UO_1136 (O_1136,N_9750,N_8100);
nand UO_1137 (O_1137,N_9421,N_8600);
or UO_1138 (O_1138,N_8427,N_9911);
and UO_1139 (O_1139,N_9966,N_8368);
and UO_1140 (O_1140,N_9891,N_9723);
xnor UO_1141 (O_1141,N_9059,N_8650);
nor UO_1142 (O_1142,N_8961,N_9401);
nor UO_1143 (O_1143,N_8721,N_9148);
and UO_1144 (O_1144,N_8599,N_8509);
xnor UO_1145 (O_1145,N_9576,N_9240);
nand UO_1146 (O_1146,N_8512,N_8752);
and UO_1147 (O_1147,N_8478,N_9080);
and UO_1148 (O_1148,N_8722,N_8896);
and UO_1149 (O_1149,N_8848,N_8669);
or UO_1150 (O_1150,N_9465,N_8616);
nor UO_1151 (O_1151,N_9866,N_8917);
and UO_1152 (O_1152,N_9956,N_9989);
nand UO_1153 (O_1153,N_8001,N_9291);
nor UO_1154 (O_1154,N_9568,N_8596);
nand UO_1155 (O_1155,N_8460,N_9346);
nor UO_1156 (O_1156,N_8983,N_9922);
nor UO_1157 (O_1157,N_9631,N_9683);
or UO_1158 (O_1158,N_8675,N_8352);
or UO_1159 (O_1159,N_9753,N_8769);
xor UO_1160 (O_1160,N_8756,N_9188);
and UO_1161 (O_1161,N_8797,N_9718);
nand UO_1162 (O_1162,N_9113,N_9582);
nand UO_1163 (O_1163,N_8662,N_8780);
and UO_1164 (O_1164,N_9806,N_9261);
nor UO_1165 (O_1165,N_9369,N_8054);
or UO_1166 (O_1166,N_8530,N_9516);
and UO_1167 (O_1167,N_9117,N_9796);
xor UO_1168 (O_1168,N_8940,N_8671);
and UO_1169 (O_1169,N_8448,N_9630);
nor UO_1170 (O_1170,N_9344,N_8600);
and UO_1171 (O_1171,N_9286,N_8859);
xnor UO_1172 (O_1172,N_9626,N_9232);
and UO_1173 (O_1173,N_9601,N_8510);
or UO_1174 (O_1174,N_9710,N_9147);
or UO_1175 (O_1175,N_8224,N_8027);
and UO_1176 (O_1176,N_8434,N_8733);
nand UO_1177 (O_1177,N_9616,N_9807);
or UO_1178 (O_1178,N_8661,N_8532);
or UO_1179 (O_1179,N_8724,N_9265);
and UO_1180 (O_1180,N_8311,N_9946);
and UO_1181 (O_1181,N_9282,N_9881);
or UO_1182 (O_1182,N_9901,N_9027);
nand UO_1183 (O_1183,N_9140,N_9152);
or UO_1184 (O_1184,N_8164,N_8012);
nor UO_1185 (O_1185,N_8642,N_9606);
nand UO_1186 (O_1186,N_8714,N_9898);
and UO_1187 (O_1187,N_9586,N_8721);
nor UO_1188 (O_1188,N_8336,N_8862);
nor UO_1189 (O_1189,N_8802,N_9591);
nor UO_1190 (O_1190,N_8353,N_9066);
nand UO_1191 (O_1191,N_9488,N_8864);
nor UO_1192 (O_1192,N_9668,N_8014);
or UO_1193 (O_1193,N_8766,N_9985);
xnor UO_1194 (O_1194,N_8116,N_8745);
xor UO_1195 (O_1195,N_9629,N_9324);
nor UO_1196 (O_1196,N_8423,N_8399);
xnor UO_1197 (O_1197,N_9210,N_9556);
nor UO_1198 (O_1198,N_9237,N_8977);
and UO_1199 (O_1199,N_9564,N_9158);
xnor UO_1200 (O_1200,N_8499,N_8111);
xor UO_1201 (O_1201,N_8335,N_8456);
or UO_1202 (O_1202,N_8162,N_8293);
nand UO_1203 (O_1203,N_8387,N_9390);
nor UO_1204 (O_1204,N_9292,N_9231);
xnor UO_1205 (O_1205,N_9280,N_9739);
nor UO_1206 (O_1206,N_8141,N_8052);
xnor UO_1207 (O_1207,N_8154,N_9445);
and UO_1208 (O_1208,N_9021,N_9250);
or UO_1209 (O_1209,N_9274,N_9138);
nand UO_1210 (O_1210,N_8949,N_8327);
xnor UO_1211 (O_1211,N_9522,N_8574);
xor UO_1212 (O_1212,N_8447,N_8516);
nand UO_1213 (O_1213,N_8248,N_9182);
or UO_1214 (O_1214,N_8531,N_8205);
nor UO_1215 (O_1215,N_9279,N_9878);
xnor UO_1216 (O_1216,N_9910,N_9236);
or UO_1217 (O_1217,N_9806,N_9540);
xnor UO_1218 (O_1218,N_8633,N_8262);
and UO_1219 (O_1219,N_8459,N_9247);
nor UO_1220 (O_1220,N_8434,N_9420);
or UO_1221 (O_1221,N_9267,N_8683);
and UO_1222 (O_1222,N_8070,N_9600);
or UO_1223 (O_1223,N_8067,N_9495);
nor UO_1224 (O_1224,N_8858,N_9864);
xor UO_1225 (O_1225,N_8708,N_8652);
or UO_1226 (O_1226,N_9389,N_9370);
nand UO_1227 (O_1227,N_9000,N_8932);
xor UO_1228 (O_1228,N_9383,N_8208);
nor UO_1229 (O_1229,N_8484,N_8718);
nand UO_1230 (O_1230,N_9800,N_8968);
nand UO_1231 (O_1231,N_8800,N_8112);
and UO_1232 (O_1232,N_9871,N_9749);
nand UO_1233 (O_1233,N_8070,N_8274);
nand UO_1234 (O_1234,N_8308,N_8772);
nand UO_1235 (O_1235,N_8161,N_8071);
and UO_1236 (O_1236,N_9009,N_9859);
or UO_1237 (O_1237,N_8416,N_8087);
or UO_1238 (O_1238,N_8980,N_8949);
xnor UO_1239 (O_1239,N_8735,N_9340);
xnor UO_1240 (O_1240,N_9179,N_9401);
nand UO_1241 (O_1241,N_9839,N_8490);
and UO_1242 (O_1242,N_8010,N_8883);
nand UO_1243 (O_1243,N_9493,N_9719);
nor UO_1244 (O_1244,N_8476,N_9843);
nand UO_1245 (O_1245,N_8535,N_9113);
nand UO_1246 (O_1246,N_9756,N_8309);
nand UO_1247 (O_1247,N_8474,N_8334);
nor UO_1248 (O_1248,N_8498,N_9948);
or UO_1249 (O_1249,N_9525,N_9986);
nor UO_1250 (O_1250,N_9124,N_9451);
and UO_1251 (O_1251,N_9342,N_9509);
xnor UO_1252 (O_1252,N_8242,N_9062);
and UO_1253 (O_1253,N_9087,N_8361);
nor UO_1254 (O_1254,N_9032,N_9257);
or UO_1255 (O_1255,N_8384,N_9779);
or UO_1256 (O_1256,N_9812,N_9611);
or UO_1257 (O_1257,N_9862,N_8594);
nand UO_1258 (O_1258,N_8532,N_8556);
nor UO_1259 (O_1259,N_8660,N_9725);
xnor UO_1260 (O_1260,N_9134,N_8559);
xor UO_1261 (O_1261,N_8436,N_8789);
and UO_1262 (O_1262,N_8657,N_8938);
xnor UO_1263 (O_1263,N_9407,N_8721);
nor UO_1264 (O_1264,N_8560,N_8734);
nor UO_1265 (O_1265,N_8588,N_8566);
nand UO_1266 (O_1266,N_9574,N_8322);
and UO_1267 (O_1267,N_8222,N_9316);
nor UO_1268 (O_1268,N_8065,N_8558);
and UO_1269 (O_1269,N_8128,N_9280);
or UO_1270 (O_1270,N_9768,N_9400);
xnor UO_1271 (O_1271,N_8704,N_8897);
nand UO_1272 (O_1272,N_9089,N_8988);
xnor UO_1273 (O_1273,N_8180,N_9005);
nand UO_1274 (O_1274,N_9759,N_8298);
nor UO_1275 (O_1275,N_8667,N_9392);
xnor UO_1276 (O_1276,N_8969,N_8812);
and UO_1277 (O_1277,N_8700,N_8720);
or UO_1278 (O_1278,N_9229,N_9875);
xor UO_1279 (O_1279,N_8811,N_9749);
xnor UO_1280 (O_1280,N_8997,N_9982);
xor UO_1281 (O_1281,N_9268,N_9774);
nand UO_1282 (O_1282,N_8928,N_8993);
xnor UO_1283 (O_1283,N_8647,N_9879);
xor UO_1284 (O_1284,N_9910,N_9822);
xnor UO_1285 (O_1285,N_9059,N_9699);
or UO_1286 (O_1286,N_8442,N_8939);
nor UO_1287 (O_1287,N_9545,N_9746);
nor UO_1288 (O_1288,N_8678,N_8567);
or UO_1289 (O_1289,N_9793,N_9506);
and UO_1290 (O_1290,N_9967,N_9635);
and UO_1291 (O_1291,N_9157,N_9089);
nand UO_1292 (O_1292,N_9864,N_8091);
or UO_1293 (O_1293,N_9745,N_8818);
and UO_1294 (O_1294,N_9583,N_9469);
xnor UO_1295 (O_1295,N_8440,N_9866);
nand UO_1296 (O_1296,N_9292,N_9153);
nand UO_1297 (O_1297,N_9592,N_9763);
xnor UO_1298 (O_1298,N_9927,N_8948);
nor UO_1299 (O_1299,N_8031,N_8058);
or UO_1300 (O_1300,N_9223,N_8302);
or UO_1301 (O_1301,N_8852,N_9086);
nand UO_1302 (O_1302,N_9234,N_8615);
nand UO_1303 (O_1303,N_8896,N_9375);
nand UO_1304 (O_1304,N_8999,N_9980);
or UO_1305 (O_1305,N_8610,N_8185);
xor UO_1306 (O_1306,N_9546,N_8643);
nand UO_1307 (O_1307,N_9483,N_8203);
and UO_1308 (O_1308,N_9821,N_9685);
xor UO_1309 (O_1309,N_9658,N_9526);
nor UO_1310 (O_1310,N_9784,N_8957);
nor UO_1311 (O_1311,N_9099,N_9664);
and UO_1312 (O_1312,N_8161,N_9187);
xnor UO_1313 (O_1313,N_8556,N_8231);
xnor UO_1314 (O_1314,N_9432,N_9677);
nand UO_1315 (O_1315,N_8639,N_9071);
xnor UO_1316 (O_1316,N_9168,N_8900);
xnor UO_1317 (O_1317,N_8308,N_8127);
nor UO_1318 (O_1318,N_9087,N_9915);
xnor UO_1319 (O_1319,N_9935,N_9776);
xnor UO_1320 (O_1320,N_9088,N_9719);
and UO_1321 (O_1321,N_9867,N_9482);
and UO_1322 (O_1322,N_8910,N_8426);
nor UO_1323 (O_1323,N_9269,N_8288);
nand UO_1324 (O_1324,N_9262,N_9166);
or UO_1325 (O_1325,N_8145,N_8175);
xnor UO_1326 (O_1326,N_9479,N_9517);
xnor UO_1327 (O_1327,N_8183,N_9426);
or UO_1328 (O_1328,N_9670,N_9252);
and UO_1329 (O_1329,N_9975,N_8601);
or UO_1330 (O_1330,N_8729,N_8656);
nand UO_1331 (O_1331,N_8282,N_8175);
or UO_1332 (O_1332,N_9296,N_9903);
and UO_1333 (O_1333,N_9717,N_8621);
xor UO_1334 (O_1334,N_9369,N_8284);
and UO_1335 (O_1335,N_8611,N_8008);
and UO_1336 (O_1336,N_8588,N_9587);
nor UO_1337 (O_1337,N_8706,N_9109);
xnor UO_1338 (O_1338,N_9801,N_8015);
nor UO_1339 (O_1339,N_8418,N_9979);
and UO_1340 (O_1340,N_9729,N_9528);
and UO_1341 (O_1341,N_9914,N_8115);
nor UO_1342 (O_1342,N_8336,N_9783);
or UO_1343 (O_1343,N_8631,N_9917);
or UO_1344 (O_1344,N_9368,N_8803);
nor UO_1345 (O_1345,N_9532,N_9531);
nand UO_1346 (O_1346,N_9363,N_9162);
nand UO_1347 (O_1347,N_8441,N_8997);
or UO_1348 (O_1348,N_9274,N_8861);
xnor UO_1349 (O_1349,N_9471,N_8212);
nand UO_1350 (O_1350,N_8437,N_9049);
xnor UO_1351 (O_1351,N_9407,N_8485);
and UO_1352 (O_1352,N_9281,N_9176);
nand UO_1353 (O_1353,N_8579,N_8827);
and UO_1354 (O_1354,N_8200,N_9700);
nand UO_1355 (O_1355,N_8048,N_9903);
nand UO_1356 (O_1356,N_9667,N_8052);
xnor UO_1357 (O_1357,N_9225,N_8181);
nand UO_1358 (O_1358,N_8855,N_8103);
and UO_1359 (O_1359,N_9794,N_8398);
or UO_1360 (O_1360,N_9992,N_9262);
nand UO_1361 (O_1361,N_9466,N_8443);
nand UO_1362 (O_1362,N_9233,N_8260);
nor UO_1363 (O_1363,N_8978,N_9084);
nand UO_1364 (O_1364,N_9450,N_9365);
and UO_1365 (O_1365,N_9247,N_8530);
nand UO_1366 (O_1366,N_8079,N_8462);
xnor UO_1367 (O_1367,N_8512,N_8369);
nand UO_1368 (O_1368,N_9817,N_8394);
and UO_1369 (O_1369,N_8094,N_8074);
or UO_1370 (O_1370,N_8019,N_9676);
nand UO_1371 (O_1371,N_9918,N_9447);
nor UO_1372 (O_1372,N_9104,N_9699);
nor UO_1373 (O_1373,N_8487,N_9296);
or UO_1374 (O_1374,N_9891,N_9084);
nand UO_1375 (O_1375,N_8517,N_8610);
nor UO_1376 (O_1376,N_8553,N_8679);
nor UO_1377 (O_1377,N_8248,N_8386);
and UO_1378 (O_1378,N_8146,N_8275);
or UO_1379 (O_1379,N_8331,N_8470);
and UO_1380 (O_1380,N_8827,N_8277);
or UO_1381 (O_1381,N_8491,N_9903);
xnor UO_1382 (O_1382,N_9589,N_9157);
nand UO_1383 (O_1383,N_8088,N_9768);
nor UO_1384 (O_1384,N_8792,N_8168);
and UO_1385 (O_1385,N_9789,N_8301);
and UO_1386 (O_1386,N_8770,N_9901);
nand UO_1387 (O_1387,N_8527,N_8479);
nand UO_1388 (O_1388,N_9687,N_9400);
or UO_1389 (O_1389,N_8025,N_9632);
xnor UO_1390 (O_1390,N_9284,N_9462);
nand UO_1391 (O_1391,N_9199,N_8705);
and UO_1392 (O_1392,N_8090,N_9731);
nor UO_1393 (O_1393,N_9366,N_8888);
xnor UO_1394 (O_1394,N_8282,N_8746);
or UO_1395 (O_1395,N_9242,N_8289);
xor UO_1396 (O_1396,N_8558,N_9005);
and UO_1397 (O_1397,N_9372,N_8903);
and UO_1398 (O_1398,N_9008,N_8963);
nand UO_1399 (O_1399,N_9049,N_9477);
or UO_1400 (O_1400,N_8341,N_8914);
nor UO_1401 (O_1401,N_9821,N_8783);
and UO_1402 (O_1402,N_9482,N_9068);
and UO_1403 (O_1403,N_9443,N_8662);
nand UO_1404 (O_1404,N_9967,N_9535);
nand UO_1405 (O_1405,N_8434,N_9205);
and UO_1406 (O_1406,N_8968,N_9075);
and UO_1407 (O_1407,N_8077,N_9647);
and UO_1408 (O_1408,N_9377,N_8732);
nor UO_1409 (O_1409,N_8853,N_9282);
or UO_1410 (O_1410,N_9229,N_8337);
or UO_1411 (O_1411,N_9107,N_8944);
nand UO_1412 (O_1412,N_8002,N_9404);
xnor UO_1413 (O_1413,N_8669,N_9642);
nor UO_1414 (O_1414,N_9428,N_8118);
or UO_1415 (O_1415,N_9783,N_8229);
xor UO_1416 (O_1416,N_8857,N_9548);
nor UO_1417 (O_1417,N_9971,N_8528);
nand UO_1418 (O_1418,N_8435,N_9749);
and UO_1419 (O_1419,N_9364,N_8197);
xnor UO_1420 (O_1420,N_8074,N_9679);
and UO_1421 (O_1421,N_8545,N_9777);
xnor UO_1422 (O_1422,N_8417,N_9128);
nor UO_1423 (O_1423,N_8622,N_9434);
or UO_1424 (O_1424,N_8410,N_8311);
or UO_1425 (O_1425,N_8940,N_9193);
and UO_1426 (O_1426,N_9099,N_9764);
xnor UO_1427 (O_1427,N_8625,N_8744);
xnor UO_1428 (O_1428,N_8433,N_8079);
nor UO_1429 (O_1429,N_9429,N_9555);
xnor UO_1430 (O_1430,N_9713,N_9211);
nand UO_1431 (O_1431,N_8603,N_9350);
and UO_1432 (O_1432,N_8917,N_9449);
nand UO_1433 (O_1433,N_9840,N_9963);
nor UO_1434 (O_1434,N_9066,N_9246);
xor UO_1435 (O_1435,N_9946,N_8429);
xnor UO_1436 (O_1436,N_9780,N_8356);
nand UO_1437 (O_1437,N_9893,N_8119);
nand UO_1438 (O_1438,N_9568,N_9473);
xnor UO_1439 (O_1439,N_8105,N_8236);
and UO_1440 (O_1440,N_9265,N_9277);
nand UO_1441 (O_1441,N_9017,N_9605);
nand UO_1442 (O_1442,N_9543,N_9044);
and UO_1443 (O_1443,N_9617,N_8954);
nand UO_1444 (O_1444,N_8387,N_8984);
or UO_1445 (O_1445,N_9590,N_9207);
nand UO_1446 (O_1446,N_9846,N_8973);
xor UO_1447 (O_1447,N_9606,N_8208);
xor UO_1448 (O_1448,N_9707,N_9957);
xor UO_1449 (O_1449,N_8178,N_9090);
nor UO_1450 (O_1450,N_8005,N_8019);
or UO_1451 (O_1451,N_9722,N_8306);
nor UO_1452 (O_1452,N_9893,N_8382);
nor UO_1453 (O_1453,N_9172,N_9592);
or UO_1454 (O_1454,N_8319,N_8637);
xor UO_1455 (O_1455,N_8177,N_9364);
and UO_1456 (O_1456,N_9411,N_9644);
nor UO_1457 (O_1457,N_8960,N_8496);
nand UO_1458 (O_1458,N_8590,N_8619);
nor UO_1459 (O_1459,N_8438,N_8281);
xor UO_1460 (O_1460,N_8680,N_8595);
or UO_1461 (O_1461,N_9315,N_9693);
and UO_1462 (O_1462,N_8647,N_8757);
nor UO_1463 (O_1463,N_8223,N_9166);
and UO_1464 (O_1464,N_8068,N_9050);
or UO_1465 (O_1465,N_9382,N_9538);
nor UO_1466 (O_1466,N_8478,N_8804);
nand UO_1467 (O_1467,N_8890,N_8552);
or UO_1468 (O_1468,N_9613,N_8309);
nor UO_1469 (O_1469,N_8017,N_9620);
nand UO_1470 (O_1470,N_9755,N_8808);
xor UO_1471 (O_1471,N_9515,N_9888);
and UO_1472 (O_1472,N_8249,N_9192);
nand UO_1473 (O_1473,N_9296,N_8781);
nand UO_1474 (O_1474,N_9844,N_9716);
and UO_1475 (O_1475,N_8923,N_8505);
nand UO_1476 (O_1476,N_9577,N_9018);
xor UO_1477 (O_1477,N_9920,N_9734);
nand UO_1478 (O_1478,N_9210,N_8895);
or UO_1479 (O_1479,N_8759,N_9720);
nor UO_1480 (O_1480,N_8640,N_9352);
and UO_1481 (O_1481,N_9845,N_9810);
nand UO_1482 (O_1482,N_8314,N_8249);
and UO_1483 (O_1483,N_8987,N_8210);
xor UO_1484 (O_1484,N_8010,N_9964);
nand UO_1485 (O_1485,N_9047,N_8111);
and UO_1486 (O_1486,N_9090,N_8957);
nand UO_1487 (O_1487,N_9269,N_9424);
nand UO_1488 (O_1488,N_9831,N_8774);
and UO_1489 (O_1489,N_9241,N_9696);
and UO_1490 (O_1490,N_9883,N_8081);
nor UO_1491 (O_1491,N_8971,N_9274);
xor UO_1492 (O_1492,N_8227,N_9901);
xor UO_1493 (O_1493,N_8885,N_8014);
and UO_1494 (O_1494,N_8619,N_9020);
or UO_1495 (O_1495,N_8751,N_8278);
nor UO_1496 (O_1496,N_8726,N_8204);
or UO_1497 (O_1497,N_9811,N_8461);
and UO_1498 (O_1498,N_9046,N_8538);
nand UO_1499 (O_1499,N_9023,N_8608);
endmodule