module basic_500_3000_500_3_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_382,In_29);
xor U1 (N_1,In_79,In_442);
and U2 (N_2,In_192,In_331);
xor U3 (N_3,In_314,In_313);
and U4 (N_4,In_438,In_159);
or U5 (N_5,In_279,In_16);
nor U6 (N_6,In_145,In_398);
nor U7 (N_7,In_104,In_483);
or U8 (N_8,In_247,In_440);
and U9 (N_9,In_168,In_453);
nand U10 (N_10,In_183,In_93);
or U11 (N_11,In_189,In_372);
or U12 (N_12,In_295,In_307);
and U13 (N_13,In_221,In_134);
or U14 (N_14,In_232,In_81);
nor U15 (N_15,In_243,In_156);
or U16 (N_16,In_369,In_188);
nor U17 (N_17,In_470,In_20);
nand U18 (N_18,In_437,In_178);
nand U19 (N_19,In_139,In_444);
or U20 (N_20,In_405,In_57);
and U21 (N_21,In_268,In_153);
xor U22 (N_22,In_388,In_476);
nand U23 (N_23,In_36,In_4);
and U24 (N_24,In_43,In_51);
and U25 (N_25,In_258,In_259);
or U26 (N_26,In_105,In_190);
or U27 (N_27,In_435,In_276);
xor U28 (N_28,In_263,In_161);
xnor U29 (N_29,In_454,In_69);
xor U30 (N_30,In_137,In_141);
xnor U31 (N_31,In_466,In_434);
or U32 (N_32,In_127,In_327);
nand U33 (N_33,In_200,In_24);
nor U34 (N_34,In_339,In_455);
nand U35 (N_35,In_167,In_251);
xor U36 (N_36,In_391,In_408);
nand U37 (N_37,In_499,In_102);
xor U38 (N_38,In_410,In_230);
nor U39 (N_39,In_30,In_478);
and U40 (N_40,In_462,In_321);
nand U41 (N_41,In_163,In_9);
nor U42 (N_42,In_103,In_487);
and U43 (N_43,In_275,In_155);
nor U44 (N_44,In_273,In_17);
or U45 (N_45,In_42,In_54);
xor U46 (N_46,In_312,In_334);
or U47 (N_47,In_254,In_427);
and U48 (N_48,In_267,In_73);
nor U49 (N_49,In_330,In_174);
and U50 (N_50,In_208,In_315);
or U51 (N_51,In_459,In_237);
xnor U52 (N_52,In_86,In_471);
and U53 (N_53,In_65,In_431);
xnor U54 (N_54,In_337,In_257);
nor U55 (N_55,In_371,In_429);
and U56 (N_56,In_458,In_222);
nand U57 (N_57,In_266,In_357);
xnor U58 (N_58,In_203,In_432);
xor U59 (N_59,In_162,In_414);
nand U60 (N_60,In_58,In_236);
or U61 (N_61,In_497,In_402);
or U62 (N_62,In_92,In_345);
or U63 (N_63,In_246,In_443);
xnor U64 (N_64,In_277,In_446);
nand U65 (N_65,In_389,In_212);
xor U66 (N_66,In_305,In_165);
and U67 (N_67,In_120,In_304);
nor U68 (N_68,In_172,In_71);
nor U69 (N_69,In_48,In_472);
nor U70 (N_70,In_490,In_456);
nor U71 (N_71,In_412,In_248);
nor U72 (N_72,In_264,In_385);
and U73 (N_73,In_419,In_113);
xor U74 (N_74,In_56,In_194);
and U75 (N_75,In_201,In_219);
nand U76 (N_76,In_352,In_491);
or U77 (N_77,In_169,In_220);
nor U78 (N_78,In_116,In_299);
xnor U79 (N_79,In_40,In_138);
xor U80 (N_80,In_89,In_433);
xor U81 (N_81,In_477,In_400);
nand U82 (N_82,In_235,In_475);
and U83 (N_83,In_34,In_50);
xor U84 (N_84,In_368,In_317);
nand U85 (N_85,In_216,In_481);
nand U86 (N_86,In_355,In_326);
xor U87 (N_87,In_423,In_347);
nand U88 (N_88,In_322,In_393);
nand U89 (N_89,In_302,In_255);
xor U90 (N_90,In_395,In_366);
xor U91 (N_91,In_150,In_492);
nand U92 (N_92,In_108,In_27);
xor U93 (N_93,In_333,In_238);
xnor U94 (N_94,In_467,In_84);
and U95 (N_95,In_319,In_328);
nor U96 (N_96,In_479,In_265);
xor U97 (N_97,In_346,In_341);
or U98 (N_98,In_70,In_82);
nand U99 (N_99,In_316,In_485);
nor U100 (N_100,In_128,In_480);
nor U101 (N_101,In_233,In_298);
or U102 (N_102,In_131,In_125);
and U103 (N_103,In_8,In_160);
and U104 (N_104,In_363,In_482);
or U105 (N_105,In_23,In_436);
and U106 (N_106,In_114,In_362);
nand U107 (N_107,In_494,In_31);
nor U108 (N_108,In_342,In_118);
nand U109 (N_109,In_488,In_404);
nand U110 (N_110,In_424,In_142);
xor U111 (N_111,In_60,In_68);
and U112 (N_112,In_223,In_375);
or U113 (N_113,In_381,In_293);
xor U114 (N_114,In_38,In_180);
nor U115 (N_115,In_422,In_1);
xor U116 (N_116,In_463,In_28);
nand U117 (N_117,In_19,In_310);
and U118 (N_118,In_226,In_418);
or U119 (N_119,In_75,In_380);
nor U120 (N_120,In_77,In_280);
nor U121 (N_121,In_452,In_354);
and U122 (N_122,In_348,In_415);
nand U123 (N_123,In_173,In_52);
and U124 (N_124,In_367,In_270);
nor U125 (N_125,In_45,In_44);
nand U126 (N_126,In_409,In_278);
or U127 (N_127,In_465,In_303);
and U128 (N_128,In_249,In_239);
or U129 (N_129,In_122,In_364);
or U130 (N_130,In_256,In_252);
nand U131 (N_131,In_394,In_241);
nand U132 (N_132,In_461,In_324);
nor U133 (N_133,In_421,In_3);
or U134 (N_134,In_164,In_66);
or U135 (N_135,In_225,In_450);
nand U136 (N_136,In_83,In_63);
and U137 (N_137,In_136,In_181);
nand U138 (N_138,In_360,In_218);
xor U139 (N_139,In_464,In_32);
xnor U140 (N_140,In_101,In_130);
nand U141 (N_141,In_109,In_379);
nand U142 (N_142,In_115,In_498);
or U143 (N_143,In_285,In_148);
nand U144 (N_144,In_90,In_336);
nand U145 (N_145,In_445,In_495);
and U146 (N_146,In_484,In_126);
and U147 (N_147,In_140,In_62);
nor U148 (N_148,In_175,In_300);
xor U149 (N_149,In_320,In_143);
nor U150 (N_150,In_343,In_119);
xor U151 (N_151,In_290,In_99);
xor U152 (N_152,In_98,In_107);
nand U153 (N_153,In_416,In_297);
xor U154 (N_154,In_274,In_7);
xor U155 (N_155,In_74,In_383);
and U156 (N_156,In_338,In_411);
xor U157 (N_157,In_151,In_396);
nor U158 (N_158,In_213,In_413);
or U159 (N_159,In_407,In_111);
and U160 (N_160,In_217,In_154);
xnor U161 (N_161,In_234,In_185);
or U162 (N_162,In_401,In_11);
nand U163 (N_163,In_387,In_95);
or U164 (N_164,In_291,In_323);
or U165 (N_165,In_392,In_365);
nand U166 (N_166,In_425,In_117);
and U167 (N_167,In_59,In_250);
and U168 (N_168,In_349,In_193);
nor U169 (N_169,In_198,In_430);
or U170 (N_170,In_417,In_85);
xnor U171 (N_171,In_26,In_78);
nand U172 (N_172,In_428,In_350);
and U173 (N_173,In_441,In_282);
nand U174 (N_174,In_309,In_97);
and U175 (N_175,In_439,In_353);
nand U176 (N_176,In_96,In_76);
nor U177 (N_177,In_376,In_157);
or U178 (N_178,In_187,In_344);
or U179 (N_179,In_384,In_426);
nor U180 (N_180,In_158,In_170);
or U181 (N_181,In_356,In_244);
or U182 (N_182,In_325,In_202);
and U183 (N_183,In_53,In_378);
nor U184 (N_184,In_493,In_449);
nand U185 (N_185,In_340,In_473);
xor U186 (N_186,In_332,In_6);
xnor U187 (N_187,In_41,In_489);
xnor U188 (N_188,In_253,In_215);
nor U189 (N_189,In_469,In_88);
nor U190 (N_190,In_260,In_123);
nand U191 (N_191,In_179,In_296);
nand U192 (N_192,In_46,In_39);
or U193 (N_193,In_5,In_289);
xnor U194 (N_194,In_373,In_205);
nand U195 (N_195,In_196,In_474);
nand U196 (N_196,In_359,In_10);
or U197 (N_197,In_308,In_242);
nand U198 (N_198,In_460,In_288);
nand U199 (N_199,In_55,In_318);
and U200 (N_200,In_448,In_152);
xor U201 (N_201,In_195,In_207);
xnor U202 (N_202,In_224,In_447);
nand U203 (N_203,In_361,In_133);
and U204 (N_204,In_49,In_420);
or U205 (N_205,In_397,In_35);
and U206 (N_206,In_147,In_149);
or U207 (N_207,In_377,In_294);
nor U208 (N_208,In_15,In_206);
nand U209 (N_209,In_272,In_186);
xor U210 (N_210,In_287,In_100);
nand U211 (N_211,In_21,In_197);
nor U212 (N_212,In_245,In_129);
xor U213 (N_213,In_144,In_12);
nor U214 (N_214,In_211,In_229);
xor U215 (N_215,In_61,In_191);
nor U216 (N_216,In_269,In_406);
xnor U217 (N_217,In_329,In_204);
nand U218 (N_218,In_335,In_214);
or U219 (N_219,In_358,In_110);
or U220 (N_220,In_457,In_261);
and U221 (N_221,In_390,In_112);
nor U222 (N_222,In_171,In_403);
and U223 (N_223,In_399,In_496);
nor U224 (N_224,In_14,In_262);
xor U225 (N_225,In_284,In_2);
nand U226 (N_226,In_351,In_184);
nand U227 (N_227,In_87,In_292);
nand U228 (N_228,In_281,In_121);
xor U229 (N_229,In_306,In_486);
nand U230 (N_230,In_370,In_146);
nand U231 (N_231,In_64,In_227);
nor U232 (N_232,In_13,In_374);
or U233 (N_233,In_166,In_132);
xnor U234 (N_234,In_386,In_22);
and U235 (N_235,In_283,In_468);
xnor U236 (N_236,In_33,In_124);
and U237 (N_237,In_210,In_199);
nand U238 (N_238,In_209,In_286);
or U239 (N_239,In_311,In_37);
and U240 (N_240,In_182,In_135);
and U241 (N_241,In_231,In_451);
nor U242 (N_242,In_240,In_228);
nand U243 (N_243,In_0,In_94);
nand U244 (N_244,In_106,In_176);
nor U245 (N_245,In_47,In_67);
nor U246 (N_246,In_177,In_72);
nand U247 (N_247,In_25,In_91);
nor U248 (N_248,In_80,In_271);
xnor U249 (N_249,In_301,In_18);
or U250 (N_250,In_410,In_417);
xor U251 (N_251,In_200,In_132);
xnor U252 (N_252,In_79,In_370);
nor U253 (N_253,In_410,In_72);
nor U254 (N_254,In_161,In_312);
nor U255 (N_255,In_214,In_380);
xor U256 (N_256,In_178,In_270);
nor U257 (N_257,In_473,In_110);
or U258 (N_258,In_295,In_140);
nor U259 (N_259,In_183,In_455);
nand U260 (N_260,In_491,In_458);
or U261 (N_261,In_301,In_381);
nor U262 (N_262,In_171,In_216);
and U263 (N_263,In_20,In_463);
and U264 (N_264,In_484,In_282);
nand U265 (N_265,In_202,In_279);
xnor U266 (N_266,In_318,In_331);
and U267 (N_267,In_73,In_438);
or U268 (N_268,In_291,In_364);
xnor U269 (N_269,In_252,In_98);
nand U270 (N_270,In_370,In_289);
or U271 (N_271,In_318,In_75);
and U272 (N_272,In_491,In_272);
nor U273 (N_273,In_107,In_371);
and U274 (N_274,In_155,In_400);
and U275 (N_275,In_409,In_19);
and U276 (N_276,In_84,In_221);
or U277 (N_277,In_54,In_57);
xnor U278 (N_278,In_234,In_406);
and U279 (N_279,In_53,In_387);
xnor U280 (N_280,In_366,In_305);
xnor U281 (N_281,In_441,In_259);
or U282 (N_282,In_150,In_230);
nand U283 (N_283,In_186,In_196);
nand U284 (N_284,In_395,In_224);
or U285 (N_285,In_319,In_446);
nand U286 (N_286,In_294,In_497);
or U287 (N_287,In_74,In_280);
or U288 (N_288,In_382,In_113);
xor U289 (N_289,In_340,In_423);
nand U290 (N_290,In_207,In_413);
xor U291 (N_291,In_242,In_422);
xnor U292 (N_292,In_203,In_237);
and U293 (N_293,In_322,In_26);
or U294 (N_294,In_112,In_429);
nor U295 (N_295,In_338,In_345);
nor U296 (N_296,In_355,In_140);
or U297 (N_297,In_424,In_464);
nor U298 (N_298,In_341,In_479);
and U299 (N_299,In_75,In_86);
or U300 (N_300,In_222,In_292);
nor U301 (N_301,In_281,In_51);
nand U302 (N_302,In_164,In_152);
xnor U303 (N_303,In_351,In_284);
nand U304 (N_304,In_129,In_369);
xor U305 (N_305,In_289,In_499);
xor U306 (N_306,In_93,In_175);
or U307 (N_307,In_170,In_101);
xnor U308 (N_308,In_233,In_318);
xnor U309 (N_309,In_462,In_124);
or U310 (N_310,In_130,In_285);
nor U311 (N_311,In_389,In_482);
xor U312 (N_312,In_198,In_82);
or U313 (N_313,In_15,In_116);
xor U314 (N_314,In_269,In_167);
xnor U315 (N_315,In_211,In_26);
or U316 (N_316,In_143,In_38);
nand U317 (N_317,In_88,In_391);
xnor U318 (N_318,In_21,In_18);
nor U319 (N_319,In_360,In_180);
and U320 (N_320,In_140,In_377);
or U321 (N_321,In_164,In_404);
and U322 (N_322,In_179,In_122);
and U323 (N_323,In_86,In_369);
nor U324 (N_324,In_452,In_256);
and U325 (N_325,In_399,In_253);
xor U326 (N_326,In_114,In_145);
xnor U327 (N_327,In_164,In_189);
xor U328 (N_328,In_447,In_93);
nor U329 (N_329,In_257,In_343);
xor U330 (N_330,In_444,In_415);
and U331 (N_331,In_256,In_180);
nor U332 (N_332,In_291,In_112);
or U333 (N_333,In_218,In_375);
nor U334 (N_334,In_283,In_399);
nor U335 (N_335,In_273,In_145);
nand U336 (N_336,In_45,In_206);
nand U337 (N_337,In_362,In_497);
xnor U338 (N_338,In_231,In_442);
xnor U339 (N_339,In_351,In_495);
or U340 (N_340,In_418,In_376);
and U341 (N_341,In_358,In_270);
nor U342 (N_342,In_33,In_332);
nand U343 (N_343,In_124,In_449);
nand U344 (N_344,In_100,In_354);
xor U345 (N_345,In_206,In_278);
nor U346 (N_346,In_353,In_271);
and U347 (N_347,In_95,In_351);
and U348 (N_348,In_239,In_201);
and U349 (N_349,In_326,In_71);
or U350 (N_350,In_176,In_320);
and U351 (N_351,In_327,In_254);
nand U352 (N_352,In_134,In_126);
or U353 (N_353,In_5,In_320);
and U354 (N_354,In_187,In_346);
and U355 (N_355,In_125,In_472);
and U356 (N_356,In_177,In_62);
nand U357 (N_357,In_237,In_198);
xnor U358 (N_358,In_121,In_275);
and U359 (N_359,In_92,In_0);
or U360 (N_360,In_156,In_391);
or U361 (N_361,In_240,In_365);
xnor U362 (N_362,In_161,In_373);
and U363 (N_363,In_485,In_361);
xor U364 (N_364,In_90,In_179);
nand U365 (N_365,In_208,In_199);
nand U366 (N_366,In_448,In_167);
or U367 (N_367,In_415,In_174);
and U368 (N_368,In_218,In_316);
and U369 (N_369,In_388,In_38);
or U370 (N_370,In_172,In_223);
and U371 (N_371,In_51,In_223);
and U372 (N_372,In_284,In_389);
and U373 (N_373,In_492,In_411);
or U374 (N_374,In_226,In_113);
xor U375 (N_375,In_304,In_29);
nand U376 (N_376,In_246,In_140);
or U377 (N_377,In_130,In_306);
and U378 (N_378,In_384,In_474);
and U379 (N_379,In_164,In_431);
or U380 (N_380,In_440,In_470);
and U381 (N_381,In_183,In_240);
and U382 (N_382,In_157,In_349);
nor U383 (N_383,In_131,In_208);
or U384 (N_384,In_373,In_248);
and U385 (N_385,In_450,In_131);
and U386 (N_386,In_284,In_465);
nand U387 (N_387,In_336,In_433);
or U388 (N_388,In_141,In_217);
nand U389 (N_389,In_410,In_321);
and U390 (N_390,In_459,In_322);
nor U391 (N_391,In_142,In_111);
nand U392 (N_392,In_78,In_485);
nor U393 (N_393,In_63,In_475);
nand U394 (N_394,In_225,In_38);
and U395 (N_395,In_448,In_145);
nor U396 (N_396,In_449,In_375);
or U397 (N_397,In_354,In_148);
nand U398 (N_398,In_499,In_369);
xor U399 (N_399,In_120,In_118);
xor U400 (N_400,In_470,In_195);
xor U401 (N_401,In_142,In_120);
xor U402 (N_402,In_496,In_380);
nand U403 (N_403,In_179,In_144);
nor U404 (N_404,In_192,In_317);
xor U405 (N_405,In_421,In_263);
and U406 (N_406,In_240,In_320);
or U407 (N_407,In_16,In_430);
and U408 (N_408,In_396,In_325);
and U409 (N_409,In_318,In_340);
or U410 (N_410,In_100,In_446);
and U411 (N_411,In_326,In_185);
nor U412 (N_412,In_430,In_252);
and U413 (N_413,In_478,In_12);
nor U414 (N_414,In_356,In_428);
nor U415 (N_415,In_11,In_129);
xnor U416 (N_416,In_181,In_299);
and U417 (N_417,In_340,In_463);
or U418 (N_418,In_183,In_8);
nand U419 (N_419,In_198,In_23);
xnor U420 (N_420,In_90,In_334);
or U421 (N_421,In_495,In_53);
nor U422 (N_422,In_203,In_172);
or U423 (N_423,In_178,In_287);
and U424 (N_424,In_130,In_384);
or U425 (N_425,In_492,In_305);
or U426 (N_426,In_493,In_454);
nand U427 (N_427,In_122,In_230);
xnor U428 (N_428,In_473,In_25);
nand U429 (N_429,In_477,In_277);
and U430 (N_430,In_150,In_82);
or U431 (N_431,In_117,In_375);
nor U432 (N_432,In_155,In_357);
nand U433 (N_433,In_7,In_56);
xor U434 (N_434,In_138,In_113);
nand U435 (N_435,In_494,In_444);
or U436 (N_436,In_455,In_120);
and U437 (N_437,In_209,In_57);
and U438 (N_438,In_112,In_129);
nor U439 (N_439,In_237,In_294);
xor U440 (N_440,In_290,In_364);
or U441 (N_441,In_224,In_145);
xor U442 (N_442,In_56,In_395);
nand U443 (N_443,In_26,In_425);
nand U444 (N_444,In_389,In_226);
nor U445 (N_445,In_137,In_491);
nor U446 (N_446,In_182,In_42);
or U447 (N_447,In_174,In_270);
nor U448 (N_448,In_52,In_97);
nor U449 (N_449,In_320,In_341);
nand U450 (N_450,In_253,In_71);
and U451 (N_451,In_395,In_17);
or U452 (N_452,In_121,In_22);
and U453 (N_453,In_370,In_1);
or U454 (N_454,In_4,In_188);
nor U455 (N_455,In_484,In_160);
or U456 (N_456,In_434,In_270);
or U457 (N_457,In_472,In_289);
or U458 (N_458,In_132,In_103);
nand U459 (N_459,In_16,In_318);
nand U460 (N_460,In_85,In_4);
nand U461 (N_461,In_418,In_242);
and U462 (N_462,In_21,In_239);
or U463 (N_463,In_40,In_1);
nand U464 (N_464,In_465,In_245);
or U465 (N_465,In_403,In_377);
xnor U466 (N_466,In_360,In_356);
xnor U467 (N_467,In_497,In_125);
nand U468 (N_468,In_311,In_282);
nor U469 (N_469,In_139,In_198);
nand U470 (N_470,In_422,In_79);
or U471 (N_471,In_365,In_204);
nor U472 (N_472,In_278,In_464);
nor U473 (N_473,In_398,In_497);
nor U474 (N_474,In_21,In_14);
xnor U475 (N_475,In_222,In_264);
nand U476 (N_476,In_35,In_258);
xor U477 (N_477,In_190,In_198);
or U478 (N_478,In_266,In_474);
and U479 (N_479,In_175,In_352);
nor U480 (N_480,In_359,In_390);
xor U481 (N_481,In_273,In_178);
nor U482 (N_482,In_310,In_234);
xor U483 (N_483,In_20,In_297);
nor U484 (N_484,In_92,In_81);
nor U485 (N_485,In_67,In_111);
nor U486 (N_486,In_110,In_483);
or U487 (N_487,In_354,In_89);
and U488 (N_488,In_498,In_72);
or U489 (N_489,In_163,In_191);
nor U490 (N_490,In_206,In_163);
nand U491 (N_491,In_61,In_38);
and U492 (N_492,In_332,In_430);
or U493 (N_493,In_404,In_460);
nor U494 (N_494,In_187,In_96);
and U495 (N_495,In_340,In_47);
xor U496 (N_496,In_280,In_32);
nor U497 (N_497,In_155,In_93);
nand U498 (N_498,In_475,In_223);
nand U499 (N_499,In_156,In_141);
and U500 (N_500,In_368,In_29);
nand U501 (N_501,In_451,In_413);
nand U502 (N_502,In_284,In_390);
and U503 (N_503,In_459,In_170);
or U504 (N_504,In_293,In_125);
and U505 (N_505,In_205,In_30);
nand U506 (N_506,In_154,In_222);
or U507 (N_507,In_224,In_210);
nand U508 (N_508,In_314,In_368);
and U509 (N_509,In_417,In_327);
xnor U510 (N_510,In_194,In_80);
nand U511 (N_511,In_371,In_299);
nand U512 (N_512,In_294,In_6);
nor U513 (N_513,In_436,In_327);
and U514 (N_514,In_352,In_120);
or U515 (N_515,In_346,In_115);
xor U516 (N_516,In_112,In_148);
and U517 (N_517,In_387,In_71);
or U518 (N_518,In_481,In_82);
nand U519 (N_519,In_55,In_386);
or U520 (N_520,In_233,In_66);
or U521 (N_521,In_179,In_20);
xnor U522 (N_522,In_162,In_215);
and U523 (N_523,In_384,In_485);
or U524 (N_524,In_136,In_149);
or U525 (N_525,In_85,In_481);
nor U526 (N_526,In_473,In_69);
or U527 (N_527,In_362,In_86);
xor U528 (N_528,In_178,In_439);
nand U529 (N_529,In_461,In_113);
or U530 (N_530,In_274,In_418);
or U531 (N_531,In_230,In_437);
and U532 (N_532,In_273,In_365);
or U533 (N_533,In_241,In_221);
and U534 (N_534,In_384,In_222);
nand U535 (N_535,In_254,In_156);
xor U536 (N_536,In_357,In_160);
nor U537 (N_537,In_332,In_165);
and U538 (N_538,In_90,In_257);
or U539 (N_539,In_187,In_410);
and U540 (N_540,In_461,In_277);
or U541 (N_541,In_418,In_299);
nor U542 (N_542,In_381,In_181);
nand U543 (N_543,In_464,In_192);
and U544 (N_544,In_459,In_50);
xnor U545 (N_545,In_389,In_293);
or U546 (N_546,In_382,In_42);
and U547 (N_547,In_290,In_418);
or U548 (N_548,In_481,In_130);
xnor U549 (N_549,In_197,In_443);
xnor U550 (N_550,In_177,In_289);
nor U551 (N_551,In_218,In_470);
nor U552 (N_552,In_213,In_269);
nor U553 (N_553,In_335,In_108);
or U554 (N_554,In_480,In_185);
nor U555 (N_555,In_392,In_280);
nand U556 (N_556,In_476,In_145);
xnor U557 (N_557,In_14,In_180);
and U558 (N_558,In_32,In_258);
nand U559 (N_559,In_363,In_83);
and U560 (N_560,In_452,In_258);
or U561 (N_561,In_164,In_228);
or U562 (N_562,In_290,In_230);
nand U563 (N_563,In_298,In_293);
or U564 (N_564,In_9,In_486);
and U565 (N_565,In_309,In_216);
or U566 (N_566,In_448,In_187);
or U567 (N_567,In_168,In_152);
nand U568 (N_568,In_88,In_18);
nor U569 (N_569,In_146,In_144);
and U570 (N_570,In_449,In_92);
and U571 (N_571,In_298,In_69);
or U572 (N_572,In_16,In_218);
nand U573 (N_573,In_86,In_183);
or U574 (N_574,In_1,In_383);
and U575 (N_575,In_355,In_164);
nor U576 (N_576,In_244,In_485);
or U577 (N_577,In_374,In_46);
xor U578 (N_578,In_357,In_380);
xnor U579 (N_579,In_182,In_2);
nor U580 (N_580,In_482,In_405);
nand U581 (N_581,In_162,In_241);
and U582 (N_582,In_73,In_163);
nand U583 (N_583,In_268,In_317);
and U584 (N_584,In_116,In_249);
or U585 (N_585,In_325,In_214);
xnor U586 (N_586,In_436,In_215);
xnor U587 (N_587,In_143,In_331);
xor U588 (N_588,In_81,In_95);
or U589 (N_589,In_28,In_496);
xor U590 (N_590,In_432,In_142);
xnor U591 (N_591,In_138,In_233);
xnor U592 (N_592,In_354,In_344);
nor U593 (N_593,In_98,In_340);
nor U594 (N_594,In_247,In_256);
or U595 (N_595,In_25,In_99);
nand U596 (N_596,In_271,In_63);
nand U597 (N_597,In_390,In_172);
nor U598 (N_598,In_46,In_321);
and U599 (N_599,In_203,In_62);
or U600 (N_600,In_363,In_436);
nand U601 (N_601,In_437,In_239);
and U602 (N_602,In_492,In_156);
xor U603 (N_603,In_415,In_419);
nand U604 (N_604,In_127,In_112);
and U605 (N_605,In_344,In_449);
and U606 (N_606,In_93,In_433);
nor U607 (N_607,In_370,In_362);
or U608 (N_608,In_466,In_187);
xnor U609 (N_609,In_145,In_5);
xnor U610 (N_610,In_230,In_261);
nand U611 (N_611,In_190,In_214);
or U612 (N_612,In_216,In_35);
or U613 (N_613,In_343,In_498);
and U614 (N_614,In_45,In_254);
and U615 (N_615,In_256,In_199);
or U616 (N_616,In_113,In_257);
xnor U617 (N_617,In_148,In_336);
xnor U618 (N_618,In_179,In_32);
nand U619 (N_619,In_11,In_421);
nor U620 (N_620,In_313,In_168);
and U621 (N_621,In_258,In_382);
nand U622 (N_622,In_231,In_96);
nand U623 (N_623,In_349,In_190);
and U624 (N_624,In_310,In_225);
or U625 (N_625,In_387,In_128);
nor U626 (N_626,In_87,In_11);
or U627 (N_627,In_389,In_251);
nor U628 (N_628,In_96,In_86);
xor U629 (N_629,In_417,In_389);
or U630 (N_630,In_60,In_193);
or U631 (N_631,In_341,In_495);
nor U632 (N_632,In_230,In_249);
nand U633 (N_633,In_72,In_482);
and U634 (N_634,In_466,In_378);
and U635 (N_635,In_397,In_350);
xnor U636 (N_636,In_241,In_185);
nand U637 (N_637,In_142,In_267);
or U638 (N_638,In_406,In_312);
nor U639 (N_639,In_328,In_102);
nor U640 (N_640,In_42,In_222);
nand U641 (N_641,In_71,In_77);
or U642 (N_642,In_443,In_387);
and U643 (N_643,In_360,In_412);
nor U644 (N_644,In_431,In_481);
and U645 (N_645,In_228,In_272);
nand U646 (N_646,In_323,In_118);
xor U647 (N_647,In_403,In_290);
nor U648 (N_648,In_388,In_296);
nand U649 (N_649,In_365,In_241);
nor U650 (N_650,In_174,In_232);
xnor U651 (N_651,In_478,In_335);
nor U652 (N_652,In_145,In_75);
and U653 (N_653,In_418,In_40);
or U654 (N_654,In_160,In_436);
nand U655 (N_655,In_495,In_402);
and U656 (N_656,In_140,In_67);
xnor U657 (N_657,In_263,In_496);
nand U658 (N_658,In_299,In_13);
nand U659 (N_659,In_418,In_43);
xnor U660 (N_660,In_432,In_232);
or U661 (N_661,In_261,In_249);
or U662 (N_662,In_132,In_268);
and U663 (N_663,In_411,In_452);
xor U664 (N_664,In_348,In_324);
and U665 (N_665,In_23,In_170);
nor U666 (N_666,In_117,In_385);
xor U667 (N_667,In_80,In_317);
xor U668 (N_668,In_55,In_148);
or U669 (N_669,In_385,In_279);
or U670 (N_670,In_17,In_164);
and U671 (N_671,In_209,In_126);
or U672 (N_672,In_301,In_172);
nor U673 (N_673,In_171,In_473);
nand U674 (N_674,In_362,In_155);
nand U675 (N_675,In_177,In_357);
nor U676 (N_676,In_490,In_301);
and U677 (N_677,In_498,In_187);
or U678 (N_678,In_163,In_77);
nor U679 (N_679,In_258,In_386);
nand U680 (N_680,In_76,In_228);
nand U681 (N_681,In_361,In_283);
nor U682 (N_682,In_9,In_196);
nand U683 (N_683,In_259,In_360);
xnor U684 (N_684,In_360,In_40);
and U685 (N_685,In_412,In_252);
or U686 (N_686,In_213,In_302);
xor U687 (N_687,In_198,In_340);
nand U688 (N_688,In_24,In_159);
xor U689 (N_689,In_293,In_319);
xor U690 (N_690,In_477,In_229);
xor U691 (N_691,In_147,In_122);
nor U692 (N_692,In_403,In_336);
or U693 (N_693,In_394,In_246);
and U694 (N_694,In_430,In_469);
xnor U695 (N_695,In_136,In_492);
or U696 (N_696,In_89,In_67);
nor U697 (N_697,In_261,In_14);
nand U698 (N_698,In_229,In_108);
and U699 (N_699,In_149,In_122);
nand U700 (N_700,In_275,In_498);
nor U701 (N_701,In_19,In_10);
nand U702 (N_702,In_38,In_110);
or U703 (N_703,In_300,In_14);
xnor U704 (N_704,In_158,In_13);
xor U705 (N_705,In_291,In_410);
nor U706 (N_706,In_469,In_193);
nand U707 (N_707,In_65,In_497);
and U708 (N_708,In_0,In_198);
nor U709 (N_709,In_227,In_287);
or U710 (N_710,In_396,In_479);
xor U711 (N_711,In_68,In_76);
nor U712 (N_712,In_77,In_245);
and U713 (N_713,In_432,In_495);
and U714 (N_714,In_372,In_76);
or U715 (N_715,In_87,In_284);
and U716 (N_716,In_480,In_265);
xor U717 (N_717,In_480,In_320);
and U718 (N_718,In_452,In_466);
or U719 (N_719,In_459,In_287);
nor U720 (N_720,In_46,In_349);
xor U721 (N_721,In_369,In_427);
xor U722 (N_722,In_156,In_358);
xor U723 (N_723,In_18,In_429);
nand U724 (N_724,In_452,In_39);
nand U725 (N_725,In_4,In_467);
and U726 (N_726,In_437,In_127);
nand U727 (N_727,In_43,In_143);
nand U728 (N_728,In_175,In_159);
or U729 (N_729,In_364,In_345);
nor U730 (N_730,In_122,In_362);
nor U731 (N_731,In_438,In_131);
nand U732 (N_732,In_65,In_130);
and U733 (N_733,In_477,In_107);
nor U734 (N_734,In_382,In_377);
xor U735 (N_735,In_320,In_22);
or U736 (N_736,In_325,In_0);
nand U737 (N_737,In_403,In_25);
xor U738 (N_738,In_319,In_178);
nor U739 (N_739,In_69,In_291);
nand U740 (N_740,In_495,In_270);
and U741 (N_741,In_8,In_304);
or U742 (N_742,In_40,In_8);
and U743 (N_743,In_286,In_438);
or U744 (N_744,In_316,In_377);
or U745 (N_745,In_203,In_255);
nor U746 (N_746,In_21,In_29);
xnor U747 (N_747,In_424,In_439);
or U748 (N_748,In_51,In_167);
and U749 (N_749,In_10,In_50);
nand U750 (N_750,In_119,In_427);
xnor U751 (N_751,In_389,In_445);
xnor U752 (N_752,In_176,In_78);
or U753 (N_753,In_157,In_483);
xor U754 (N_754,In_4,In_143);
nor U755 (N_755,In_481,In_140);
nand U756 (N_756,In_181,In_25);
xor U757 (N_757,In_364,In_275);
nand U758 (N_758,In_70,In_10);
or U759 (N_759,In_24,In_336);
and U760 (N_760,In_142,In_105);
nand U761 (N_761,In_236,In_124);
xor U762 (N_762,In_393,In_495);
xor U763 (N_763,In_418,In_85);
xor U764 (N_764,In_319,In_36);
xor U765 (N_765,In_232,In_445);
nor U766 (N_766,In_68,In_399);
nor U767 (N_767,In_100,In_202);
xor U768 (N_768,In_182,In_396);
or U769 (N_769,In_339,In_163);
or U770 (N_770,In_458,In_94);
nand U771 (N_771,In_140,In_301);
xnor U772 (N_772,In_28,In_493);
and U773 (N_773,In_124,In_308);
nand U774 (N_774,In_139,In_491);
and U775 (N_775,In_281,In_113);
xor U776 (N_776,In_431,In_88);
nor U777 (N_777,In_164,In_380);
and U778 (N_778,In_62,In_366);
xor U779 (N_779,In_146,In_322);
or U780 (N_780,In_411,In_462);
nand U781 (N_781,In_98,In_48);
nor U782 (N_782,In_300,In_368);
nand U783 (N_783,In_171,In_209);
xor U784 (N_784,In_296,In_306);
or U785 (N_785,In_99,In_470);
xor U786 (N_786,In_172,In_121);
xor U787 (N_787,In_448,In_234);
and U788 (N_788,In_247,In_151);
xnor U789 (N_789,In_101,In_63);
xnor U790 (N_790,In_459,In_388);
nor U791 (N_791,In_297,In_72);
nor U792 (N_792,In_388,In_178);
xnor U793 (N_793,In_290,In_188);
nand U794 (N_794,In_357,In_410);
and U795 (N_795,In_438,In_229);
xnor U796 (N_796,In_274,In_29);
and U797 (N_797,In_222,In_345);
xnor U798 (N_798,In_185,In_79);
and U799 (N_799,In_416,In_198);
or U800 (N_800,In_494,In_224);
nor U801 (N_801,In_86,In_66);
and U802 (N_802,In_323,In_329);
and U803 (N_803,In_410,In_106);
or U804 (N_804,In_314,In_19);
xor U805 (N_805,In_405,In_410);
nand U806 (N_806,In_99,In_161);
and U807 (N_807,In_253,In_279);
nor U808 (N_808,In_188,In_124);
nand U809 (N_809,In_21,In_351);
nand U810 (N_810,In_394,In_150);
nor U811 (N_811,In_222,In_373);
nor U812 (N_812,In_202,In_330);
and U813 (N_813,In_489,In_16);
or U814 (N_814,In_367,In_386);
or U815 (N_815,In_46,In_415);
and U816 (N_816,In_320,In_92);
or U817 (N_817,In_376,In_210);
nand U818 (N_818,In_53,In_203);
nand U819 (N_819,In_18,In_364);
nor U820 (N_820,In_57,In_239);
and U821 (N_821,In_449,In_244);
nand U822 (N_822,In_187,In_486);
or U823 (N_823,In_285,In_340);
nor U824 (N_824,In_165,In_122);
nor U825 (N_825,In_50,In_35);
nor U826 (N_826,In_396,In_162);
xnor U827 (N_827,In_146,In_51);
or U828 (N_828,In_163,In_199);
nor U829 (N_829,In_50,In_214);
nor U830 (N_830,In_266,In_231);
nor U831 (N_831,In_483,In_139);
and U832 (N_832,In_95,In_252);
and U833 (N_833,In_158,In_336);
or U834 (N_834,In_334,In_344);
or U835 (N_835,In_256,In_109);
nand U836 (N_836,In_433,In_157);
nand U837 (N_837,In_351,In_411);
or U838 (N_838,In_31,In_202);
or U839 (N_839,In_294,In_491);
xor U840 (N_840,In_476,In_420);
nor U841 (N_841,In_180,In_194);
nor U842 (N_842,In_477,In_152);
nor U843 (N_843,In_447,In_103);
or U844 (N_844,In_63,In_122);
or U845 (N_845,In_39,In_0);
nand U846 (N_846,In_430,In_114);
and U847 (N_847,In_275,In_85);
xnor U848 (N_848,In_194,In_461);
and U849 (N_849,In_334,In_25);
or U850 (N_850,In_45,In_386);
or U851 (N_851,In_87,In_248);
or U852 (N_852,In_123,In_408);
xnor U853 (N_853,In_141,In_274);
and U854 (N_854,In_318,In_40);
or U855 (N_855,In_294,In_49);
or U856 (N_856,In_237,In_31);
and U857 (N_857,In_435,In_97);
nor U858 (N_858,In_453,In_100);
xor U859 (N_859,In_250,In_291);
or U860 (N_860,In_114,In_101);
nand U861 (N_861,In_224,In_343);
or U862 (N_862,In_491,In_126);
or U863 (N_863,In_222,In_281);
xnor U864 (N_864,In_185,In_208);
nor U865 (N_865,In_154,In_63);
xnor U866 (N_866,In_341,In_380);
and U867 (N_867,In_280,In_243);
and U868 (N_868,In_264,In_27);
xnor U869 (N_869,In_71,In_78);
xnor U870 (N_870,In_195,In_206);
xnor U871 (N_871,In_378,In_271);
or U872 (N_872,In_196,In_268);
nor U873 (N_873,In_332,In_359);
nor U874 (N_874,In_305,In_455);
and U875 (N_875,In_85,In_264);
or U876 (N_876,In_481,In_385);
and U877 (N_877,In_50,In_64);
or U878 (N_878,In_465,In_300);
and U879 (N_879,In_439,In_88);
and U880 (N_880,In_303,In_99);
nand U881 (N_881,In_115,In_199);
and U882 (N_882,In_72,In_318);
or U883 (N_883,In_48,In_86);
xor U884 (N_884,In_27,In_365);
nor U885 (N_885,In_468,In_68);
nor U886 (N_886,In_441,In_486);
and U887 (N_887,In_245,In_362);
nor U888 (N_888,In_499,In_375);
or U889 (N_889,In_403,In_459);
xnor U890 (N_890,In_437,In_160);
nand U891 (N_891,In_20,In_358);
nand U892 (N_892,In_417,In_76);
xnor U893 (N_893,In_379,In_367);
nor U894 (N_894,In_327,In_70);
and U895 (N_895,In_251,In_20);
and U896 (N_896,In_43,In_58);
or U897 (N_897,In_46,In_435);
or U898 (N_898,In_258,In_13);
and U899 (N_899,In_221,In_175);
and U900 (N_900,In_100,In_293);
nand U901 (N_901,In_199,In_323);
nor U902 (N_902,In_297,In_272);
nor U903 (N_903,In_55,In_371);
xor U904 (N_904,In_496,In_315);
nand U905 (N_905,In_122,In_281);
xnor U906 (N_906,In_313,In_33);
nor U907 (N_907,In_167,In_449);
and U908 (N_908,In_6,In_26);
nor U909 (N_909,In_276,In_436);
nor U910 (N_910,In_77,In_4);
or U911 (N_911,In_261,In_120);
or U912 (N_912,In_113,In_199);
xnor U913 (N_913,In_337,In_50);
nand U914 (N_914,In_85,In_462);
nand U915 (N_915,In_239,In_479);
or U916 (N_916,In_288,In_267);
and U917 (N_917,In_346,In_297);
xor U918 (N_918,In_201,In_326);
and U919 (N_919,In_324,In_403);
nand U920 (N_920,In_302,In_401);
nor U921 (N_921,In_371,In_432);
xnor U922 (N_922,In_263,In_482);
nor U923 (N_923,In_358,In_200);
xnor U924 (N_924,In_473,In_253);
nand U925 (N_925,In_232,In_80);
nand U926 (N_926,In_307,In_102);
xor U927 (N_927,In_176,In_161);
nand U928 (N_928,In_416,In_61);
nor U929 (N_929,In_271,In_398);
and U930 (N_930,In_228,In_229);
or U931 (N_931,In_57,In_234);
nand U932 (N_932,In_277,In_259);
xnor U933 (N_933,In_209,In_54);
and U934 (N_934,In_452,In_66);
nor U935 (N_935,In_208,In_279);
or U936 (N_936,In_364,In_470);
and U937 (N_937,In_1,In_291);
xnor U938 (N_938,In_119,In_321);
nor U939 (N_939,In_51,In_333);
or U940 (N_940,In_210,In_77);
and U941 (N_941,In_464,In_85);
or U942 (N_942,In_465,In_399);
or U943 (N_943,In_177,In_136);
or U944 (N_944,In_232,In_11);
xor U945 (N_945,In_110,In_492);
or U946 (N_946,In_437,In_17);
or U947 (N_947,In_105,In_78);
and U948 (N_948,In_497,In_299);
xor U949 (N_949,In_487,In_371);
xor U950 (N_950,In_53,In_288);
xor U951 (N_951,In_354,In_217);
nor U952 (N_952,In_180,In_291);
nor U953 (N_953,In_381,In_242);
and U954 (N_954,In_326,In_63);
or U955 (N_955,In_390,In_141);
nand U956 (N_956,In_169,In_289);
xnor U957 (N_957,In_340,In_3);
and U958 (N_958,In_341,In_49);
or U959 (N_959,In_252,In_142);
or U960 (N_960,In_421,In_118);
nor U961 (N_961,In_150,In_351);
nand U962 (N_962,In_458,In_443);
and U963 (N_963,In_60,In_330);
nor U964 (N_964,In_174,In_463);
nand U965 (N_965,In_31,In_105);
nand U966 (N_966,In_445,In_370);
nand U967 (N_967,In_405,In_150);
xnor U968 (N_968,In_112,In_357);
nor U969 (N_969,In_326,In_357);
nor U970 (N_970,In_363,In_290);
and U971 (N_971,In_385,In_386);
and U972 (N_972,In_29,In_261);
and U973 (N_973,In_122,In_0);
or U974 (N_974,In_107,In_300);
and U975 (N_975,In_379,In_186);
nand U976 (N_976,In_378,In_383);
or U977 (N_977,In_68,In_425);
and U978 (N_978,In_105,In_461);
xnor U979 (N_979,In_307,In_442);
nor U980 (N_980,In_168,In_297);
or U981 (N_981,In_370,In_465);
xnor U982 (N_982,In_233,In_368);
xnor U983 (N_983,In_245,In_66);
nor U984 (N_984,In_239,In_224);
nor U985 (N_985,In_85,In_239);
xor U986 (N_986,In_462,In_325);
or U987 (N_987,In_223,In_312);
nor U988 (N_988,In_50,In_149);
nor U989 (N_989,In_111,In_471);
or U990 (N_990,In_51,In_367);
xor U991 (N_991,In_334,In_461);
xnor U992 (N_992,In_369,In_415);
nor U993 (N_993,In_119,In_76);
nand U994 (N_994,In_89,In_225);
nor U995 (N_995,In_360,In_166);
nand U996 (N_996,In_353,In_396);
or U997 (N_997,In_287,In_196);
or U998 (N_998,In_371,In_320);
and U999 (N_999,In_154,In_12);
and U1000 (N_1000,N_339,N_66);
nor U1001 (N_1001,N_861,N_615);
and U1002 (N_1002,N_34,N_602);
nor U1003 (N_1003,N_797,N_459);
nand U1004 (N_1004,N_305,N_848);
nand U1005 (N_1005,N_824,N_439);
xnor U1006 (N_1006,N_450,N_357);
nand U1007 (N_1007,N_814,N_639);
and U1008 (N_1008,N_990,N_867);
nand U1009 (N_1009,N_191,N_88);
xnor U1010 (N_1010,N_839,N_581);
xor U1011 (N_1011,N_226,N_155);
xnor U1012 (N_1012,N_908,N_500);
nor U1013 (N_1013,N_181,N_886);
nor U1014 (N_1014,N_99,N_370);
xor U1015 (N_1015,N_249,N_711);
and U1016 (N_1016,N_426,N_457);
xnor U1017 (N_1017,N_464,N_510);
nor U1018 (N_1018,N_919,N_157);
nor U1019 (N_1019,N_698,N_25);
nor U1020 (N_1020,N_768,N_134);
xor U1021 (N_1021,N_781,N_918);
or U1022 (N_1022,N_140,N_132);
xnor U1023 (N_1023,N_75,N_383);
nor U1024 (N_1024,N_692,N_350);
nand U1025 (N_1025,N_379,N_763);
or U1026 (N_1026,N_505,N_913);
or U1027 (N_1027,N_153,N_72);
xnor U1028 (N_1028,N_588,N_926);
or U1029 (N_1029,N_605,N_810);
nand U1030 (N_1030,N_257,N_179);
nand U1031 (N_1031,N_770,N_558);
nand U1032 (N_1032,N_633,N_598);
nor U1033 (N_1033,N_45,N_859);
nor U1034 (N_1034,N_219,N_338);
nand U1035 (N_1035,N_858,N_67);
nand U1036 (N_1036,N_728,N_309);
nand U1037 (N_1037,N_182,N_233);
xnor U1038 (N_1038,N_991,N_80);
xor U1039 (N_1039,N_653,N_934);
xnor U1040 (N_1040,N_941,N_661);
xnor U1041 (N_1041,N_300,N_917);
nor U1042 (N_1042,N_241,N_963);
nor U1043 (N_1043,N_599,N_611);
nand U1044 (N_1044,N_463,N_489);
xnor U1045 (N_1045,N_641,N_819);
nor U1046 (N_1046,N_275,N_499);
xnor U1047 (N_1047,N_180,N_374);
and U1048 (N_1048,N_168,N_947);
xor U1049 (N_1049,N_929,N_16);
and U1050 (N_1050,N_703,N_263);
nand U1051 (N_1051,N_412,N_937);
or U1052 (N_1052,N_590,N_519);
xor U1053 (N_1053,N_630,N_758);
or U1054 (N_1054,N_877,N_667);
or U1055 (N_1055,N_892,N_515);
or U1056 (N_1056,N_416,N_900);
xnor U1057 (N_1057,N_609,N_248);
and U1058 (N_1058,N_407,N_22);
or U1059 (N_1059,N_230,N_662);
or U1060 (N_1060,N_212,N_869);
nand U1061 (N_1061,N_465,N_396);
nand U1062 (N_1062,N_358,N_643);
xor U1063 (N_1063,N_816,N_44);
nor U1064 (N_1064,N_793,N_488);
or U1065 (N_1065,N_328,N_552);
or U1066 (N_1066,N_835,N_749);
xnor U1067 (N_1067,N_687,N_190);
nor U1068 (N_1068,N_647,N_906);
xnor U1069 (N_1069,N_264,N_894);
or U1070 (N_1070,N_270,N_887);
nor U1071 (N_1071,N_635,N_85);
nand U1072 (N_1072,N_691,N_575);
and U1073 (N_1073,N_211,N_924);
and U1074 (N_1074,N_844,N_452);
and U1075 (N_1075,N_369,N_845);
and U1076 (N_1076,N_149,N_502);
xnor U1077 (N_1077,N_923,N_889);
nand U1078 (N_1078,N_112,N_659);
xnor U1079 (N_1079,N_145,N_138);
nand U1080 (N_1080,N_517,N_534);
nand U1081 (N_1081,N_652,N_367);
nor U1082 (N_1082,N_785,N_24);
nand U1083 (N_1083,N_621,N_490);
nor U1084 (N_1084,N_291,N_612);
nand U1085 (N_1085,N_930,N_764);
and U1086 (N_1086,N_429,N_782);
or U1087 (N_1087,N_314,N_569);
xor U1088 (N_1088,N_658,N_259);
nor U1089 (N_1089,N_999,N_366);
and U1090 (N_1090,N_8,N_880);
and U1091 (N_1091,N_156,N_953);
or U1092 (N_1092,N_716,N_289);
xnor U1093 (N_1093,N_444,N_287);
xnor U1094 (N_1094,N_94,N_121);
xor U1095 (N_1095,N_495,N_55);
xor U1096 (N_1096,N_343,N_221);
or U1097 (N_1097,N_903,N_745);
nand U1098 (N_1098,N_318,N_513);
and U1099 (N_1099,N_165,N_595);
xnor U1100 (N_1100,N_755,N_122);
nor U1101 (N_1101,N_574,N_281);
xor U1102 (N_1102,N_821,N_205);
and U1103 (N_1103,N_316,N_954);
and U1104 (N_1104,N_158,N_202);
nor U1105 (N_1105,N_430,N_402);
nor U1106 (N_1106,N_117,N_881);
nand U1107 (N_1107,N_127,N_719);
xor U1108 (N_1108,N_696,N_532);
xor U1109 (N_1109,N_186,N_177);
and U1110 (N_1110,N_722,N_110);
nand U1111 (N_1111,N_812,N_794);
and U1112 (N_1112,N_584,N_600);
nor U1113 (N_1113,N_362,N_272);
xnor U1114 (N_1114,N_497,N_123);
and U1115 (N_1115,N_503,N_129);
or U1116 (N_1116,N_139,N_415);
xor U1117 (N_1117,N_298,N_322);
and U1118 (N_1118,N_256,N_284);
or U1119 (N_1119,N_160,N_458);
xnor U1120 (N_1120,N_980,N_167);
nor U1121 (N_1121,N_218,N_262);
xor U1122 (N_1122,N_619,N_627);
xor U1123 (N_1123,N_258,N_818);
and U1124 (N_1124,N_509,N_104);
xnor U1125 (N_1125,N_724,N_232);
nor U1126 (N_1126,N_660,N_949);
or U1127 (N_1127,N_688,N_111);
and U1128 (N_1128,N_432,N_494);
nor U1129 (N_1129,N_17,N_62);
nand U1130 (N_1130,N_341,N_196);
or U1131 (N_1131,N_637,N_141);
nand U1132 (N_1132,N_280,N_209);
and U1133 (N_1133,N_197,N_484);
or U1134 (N_1134,N_418,N_455);
nand U1135 (N_1135,N_670,N_86);
nand U1136 (N_1136,N_936,N_411);
nand U1137 (N_1137,N_786,N_713);
nor U1138 (N_1138,N_622,N_740);
or U1139 (N_1139,N_486,N_796);
and U1140 (N_1140,N_390,N_706);
and U1141 (N_1141,N_337,N_545);
and U1142 (N_1142,N_126,N_538);
or U1143 (N_1143,N_817,N_52);
and U1144 (N_1144,N_617,N_580);
nand U1145 (N_1145,N_119,N_285);
nand U1146 (N_1146,N_260,N_556);
nor U1147 (N_1147,N_616,N_512);
or U1148 (N_1148,N_384,N_474);
xnor U1149 (N_1149,N_0,N_741);
or U1150 (N_1150,N_335,N_511);
or U1151 (N_1151,N_92,N_884);
xnor U1152 (N_1152,N_29,N_53);
or U1153 (N_1153,N_323,N_224);
xnor U1154 (N_1154,N_345,N_32);
nand U1155 (N_1155,N_665,N_524);
nor U1156 (N_1156,N_307,N_475);
or U1157 (N_1157,N_888,N_787);
and U1158 (N_1158,N_142,N_244);
nand U1159 (N_1159,N_840,N_225);
and U1160 (N_1160,N_433,N_471);
nand U1161 (N_1161,N_700,N_736);
and U1162 (N_1162,N_306,N_21);
nor U1163 (N_1163,N_482,N_557);
nor U1164 (N_1164,N_792,N_685);
or U1165 (N_1165,N_65,N_295);
xor U1166 (N_1166,N_163,N_666);
xor U1167 (N_1167,N_297,N_240);
and U1168 (N_1168,N_456,N_978);
nor U1169 (N_1169,N_276,N_128);
or U1170 (N_1170,N_431,N_613);
or U1171 (N_1171,N_638,N_472);
nor U1172 (N_1172,N_7,N_864);
nor U1173 (N_1173,N_152,N_251);
or U1174 (N_1174,N_820,N_576);
or U1175 (N_1175,N_645,N_583);
xor U1176 (N_1176,N_485,N_811);
xnor U1177 (N_1177,N_198,N_71);
nand U1178 (N_1178,N_996,N_108);
nand U1179 (N_1179,N_995,N_164);
and U1180 (N_1180,N_435,N_169);
nor U1181 (N_1181,N_773,N_981);
or U1182 (N_1182,N_721,N_823);
nor U1183 (N_1183,N_118,N_399);
nor U1184 (N_1184,N_800,N_705);
nand U1185 (N_1185,N_247,N_909);
or U1186 (N_1186,N_380,N_33);
nor U1187 (N_1187,N_321,N_46);
or U1188 (N_1188,N_237,N_84);
xnor U1189 (N_1189,N_730,N_945);
xnor U1190 (N_1190,N_77,N_765);
nand U1191 (N_1191,N_354,N_253);
xnor U1192 (N_1192,N_234,N_971);
nor U1193 (N_1193,N_842,N_742);
and U1194 (N_1194,N_695,N_359);
nor U1195 (N_1195,N_650,N_686);
nor U1196 (N_1196,N_833,N_625);
nand U1197 (N_1197,N_353,N_697);
nor U1198 (N_1198,N_543,N_912);
nor U1199 (N_1199,N_408,N_680);
and U1200 (N_1200,N_105,N_493);
xnor U1201 (N_1201,N_352,N_663);
and U1202 (N_1202,N_571,N_363);
nor U1203 (N_1203,N_883,N_18);
nor U1204 (N_1204,N_831,N_9);
nor U1205 (N_1205,N_231,N_201);
and U1206 (N_1206,N_970,N_739);
xnor U1207 (N_1207,N_674,N_644);
or U1208 (N_1208,N_438,N_355);
nand U1209 (N_1209,N_228,N_100);
or U1210 (N_1210,N_572,N_213);
nand U1211 (N_1211,N_563,N_434);
and U1212 (N_1212,N_63,N_549);
xnor U1213 (N_1213,N_546,N_172);
and U1214 (N_1214,N_422,N_95);
nor U1215 (N_1215,N_31,N_677);
nor U1216 (N_1216,N_397,N_273);
and U1217 (N_1217,N_531,N_114);
or U1218 (N_1218,N_451,N_732);
and U1219 (N_1219,N_51,N_246);
and U1220 (N_1220,N_43,N_116);
xnor U1221 (N_1221,N_540,N_162);
nand U1222 (N_1222,N_690,N_346);
nand U1223 (N_1223,N_807,N_907);
and U1224 (N_1224,N_317,N_746);
and U1225 (N_1225,N_520,N_57);
and U1226 (N_1226,N_320,N_943);
or U1227 (N_1227,N_351,N_671);
nor U1228 (N_1228,N_938,N_561);
nand U1229 (N_1229,N_12,N_548);
nor U1230 (N_1230,N_97,N_301);
nand U1231 (N_1231,N_725,N_39);
nor U1232 (N_1232,N_239,N_441);
or U1233 (N_1233,N_368,N_330);
nor U1234 (N_1234,N_727,N_928);
and U1235 (N_1235,N_395,N_3);
nand U1236 (N_1236,N_70,N_206);
nand U1237 (N_1237,N_476,N_767);
xnor U1238 (N_1238,N_779,N_398);
xor U1239 (N_1239,N_185,N_878);
nand U1240 (N_1240,N_752,N_468);
nand U1241 (N_1241,N_526,N_506);
and U1242 (N_1242,N_400,N_589);
xnor U1243 (N_1243,N_536,N_76);
xnor U1244 (N_1244,N_784,N_679);
nand U1245 (N_1245,N_203,N_13);
and U1246 (N_1246,N_81,N_757);
and U1247 (N_1247,N_579,N_89);
nand U1248 (N_1248,N_529,N_603);
nand U1249 (N_1249,N_657,N_216);
and U1250 (N_1250,N_559,N_299);
nand U1251 (N_1251,N_853,N_731);
and U1252 (N_1252,N_414,N_646);
nor U1253 (N_1253,N_377,N_290);
nand U1254 (N_1254,N_601,N_738);
or U1255 (N_1255,N_699,N_857);
or U1256 (N_1256,N_766,N_189);
nand U1257 (N_1257,N_146,N_274);
nand U1258 (N_1258,N_340,N_326);
or U1259 (N_1259,N_760,N_669);
xnor U1260 (N_1260,N_446,N_480);
or U1261 (N_1261,N_882,N_501);
or U1262 (N_1262,N_542,N_150);
nand U1263 (N_1263,N_154,N_860);
xor U1264 (N_1264,N_523,N_735);
nand U1265 (N_1265,N_242,N_743);
or U1266 (N_1266,N_235,N_516);
xnor U1267 (N_1267,N_82,N_130);
xnor U1268 (N_1268,N_238,N_870);
xnor U1269 (N_1269,N_626,N_11);
and U1270 (N_1270,N_23,N_445);
nand U1271 (N_1271,N_243,N_496);
or U1272 (N_1272,N_885,N_762);
or U1273 (N_1273,N_401,N_729);
nor U1274 (N_1274,N_440,N_855);
nand U1275 (N_1275,N_608,N_544);
nor U1276 (N_1276,N_862,N_998);
nand U1277 (N_1277,N_950,N_944);
nand U1278 (N_1278,N_606,N_958);
nor U1279 (N_1279,N_261,N_40);
xor U1280 (N_1280,N_905,N_560);
nor U1281 (N_1281,N_460,N_10);
and U1282 (N_1282,N_871,N_946);
and U1283 (N_1283,N_829,N_902);
nor U1284 (N_1284,N_443,N_592);
nand U1285 (N_1285,N_843,N_772);
xor U1286 (N_1286,N_19,N_360);
or U1287 (N_1287,N_148,N_504);
nor U1288 (N_1288,N_551,N_492);
xnor U1289 (N_1289,N_610,N_992);
and U1290 (N_1290,N_550,N_268);
or U1291 (N_1291,N_775,N_419);
nor U1292 (N_1292,N_751,N_789);
and U1293 (N_1293,N_267,N_979);
xnor U1294 (N_1294,N_537,N_147);
xnor U1295 (N_1295,N_56,N_329);
nor U1296 (N_1296,N_804,N_702);
or U1297 (N_1297,N_447,N_364);
and U1298 (N_1298,N_710,N_873);
nor U1299 (N_1299,N_910,N_708);
nor U1300 (N_1300,N_356,N_994);
xnor U1301 (N_1301,N_73,N_997);
xnor U1302 (N_1302,N_125,N_327);
xnor U1303 (N_1303,N_522,N_678);
and U1304 (N_1304,N_373,N_808);
xor U1305 (N_1305,N_391,N_204);
or U1306 (N_1306,N_106,N_54);
nor U1307 (N_1307,N_777,N_521);
and U1308 (N_1308,N_838,N_801);
nand U1309 (N_1309,N_596,N_651);
xnor U1310 (N_1310,N_325,N_932);
nand U1311 (N_1311,N_208,N_896);
or U1312 (N_1312,N_969,N_254);
or U1313 (N_1313,N_931,N_668);
or U1314 (N_1314,N_311,N_308);
nand U1315 (N_1315,N_491,N_962);
and U1316 (N_1316,N_107,N_378);
or U1317 (N_1317,N_294,N_675);
nor U1318 (N_1318,N_895,N_279);
and U1319 (N_1319,N_826,N_734);
and U1320 (N_1320,N_282,N_361);
xnor U1321 (N_1321,N_915,N_101);
nand U1322 (N_1322,N_642,N_1);
nand U1323 (N_1323,N_974,N_554);
or U1324 (N_1324,N_791,N_587);
nor U1325 (N_1325,N_957,N_649);
xor U1326 (N_1326,N_539,N_682);
xnor U1327 (N_1327,N_737,N_847);
xor U1328 (N_1328,N_577,N_709);
nand U1329 (N_1329,N_803,N_683);
and U1330 (N_1330,N_283,N_334);
or U1331 (N_1331,N_866,N_161);
and U1332 (N_1332,N_229,N_223);
xor U1333 (N_1333,N_614,N_69);
xor U1334 (N_1334,N_759,N_87);
or U1335 (N_1335,N_41,N_850);
and U1336 (N_1336,N_109,N_806);
nand U1337 (N_1337,N_776,N_20);
and U1338 (N_1338,N_78,N_215);
nor U1339 (N_1339,N_98,N_222);
and U1340 (N_1340,N_347,N_640);
nand U1341 (N_1341,N_966,N_333);
nand U1342 (N_1342,N_933,N_79);
or U1343 (N_1343,N_113,N_591);
and U1344 (N_1344,N_720,N_977);
xor U1345 (N_1345,N_133,N_406);
nand U1346 (N_1346,N_483,N_175);
nand U1347 (N_1347,N_959,N_193);
xnor U1348 (N_1348,N_916,N_856);
nand U1349 (N_1349,N_310,N_813);
or U1350 (N_1350,N_712,N_976);
or U1351 (N_1351,N_940,N_195);
or U1352 (N_1352,N_61,N_879);
xor U1353 (N_1353,N_684,N_891);
nor U1354 (N_1354,N_304,N_47);
nand U1355 (N_1355,N_942,N_948);
or U1356 (N_1356,N_344,N_467);
and U1357 (N_1357,N_780,N_96);
nand U1358 (N_1358,N_771,N_255);
and U1359 (N_1359,N_952,N_135);
and U1360 (N_1360,N_372,N_849);
and U1361 (N_1361,N_939,N_371);
xor U1362 (N_1362,N_137,N_6);
and U1363 (N_1363,N_473,N_562);
and U1364 (N_1364,N_982,N_876);
and U1365 (N_1365,N_58,N_704);
nor U1366 (N_1366,N_836,N_236);
nand U1367 (N_1367,N_487,N_90);
nand U1368 (N_1368,N_35,N_809);
xnor U1369 (N_1369,N_798,N_171);
or U1370 (N_1370,N_220,N_393);
xor U1371 (N_1371,N_694,N_424);
xnor U1372 (N_1372,N_783,N_960);
nor U1373 (N_1373,N_2,N_754);
or U1374 (N_1374,N_693,N_717);
xor U1375 (N_1375,N_897,N_744);
nand U1376 (N_1376,N_597,N_846);
xor U1377 (N_1377,N_832,N_348);
or U1378 (N_1378,N_893,N_921);
nand U1379 (N_1379,N_968,N_403);
and U1380 (N_1380,N_387,N_750);
xor U1381 (N_1381,N_631,N_336);
nand U1382 (N_1382,N_528,N_927);
and U1383 (N_1383,N_586,N_381);
or U1384 (N_1384,N_324,N_795);
xnor U1385 (N_1385,N_541,N_565);
nor U1386 (N_1386,N_673,N_269);
nand U1387 (N_1387,N_629,N_604);
nand U1388 (N_1388,N_394,N_296);
nor U1389 (N_1389,N_64,N_618);
nand U1390 (N_1390,N_173,N_115);
nand U1391 (N_1391,N_530,N_664);
nor U1392 (N_1392,N_250,N_555);
or U1393 (N_1393,N_124,N_922);
xnor U1394 (N_1394,N_707,N_187);
xor U1395 (N_1395,N_428,N_382);
xor U1396 (N_1396,N_830,N_200);
nand U1397 (N_1397,N_131,N_527);
nand U1398 (N_1398,N_176,N_961);
nor U1399 (N_1399,N_533,N_170);
xnor U1400 (N_1400,N_478,N_413);
and U1401 (N_1401,N_26,N_989);
xnor U1402 (N_1402,N_50,N_827);
xor U1403 (N_1403,N_5,N_28);
nor U1404 (N_1404,N_747,N_761);
and U1405 (N_1405,N_453,N_194);
xor U1406 (N_1406,N_508,N_648);
or U1407 (N_1407,N_214,N_975);
nand U1408 (N_1408,N_210,N_822);
xnor U1409 (N_1409,N_828,N_442);
xnor U1410 (N_1410,N_967,N_634);
nand U1411 (N_1411,N_837,N_68);
or U1412 (N_1412,N_834,N_143);
nor U1413 (N_1413,N_983,N_376);
nor U1414 (N_1414,N_993,N_37);
and U1415 (N_1415,N_514,N_748);
or U1416 (N_1416,N_436,N_38);
nand U1417 (N_1417,N_964,N_778);
nand U1418 (N_1418,N_547,N_449);
nand U1419 (N_1419,N_217,N_417);
nor U1420 (N_1420,N_375,N_278);
or U1421 (N_1421,N_715,N_872);
xor U1422 (N_1422,N_911,N_689);
and U1423 (N_1423,N_462,N_404);
nor U1424 (N_1424,N_753,N_525);
or U1425 (N_1425,N_14,N_349);
xor U1426 (N_1426,N_973,N_578);
or U1427 (N_1427,N_899,N_410);
xor U1428 (N_1428,N_568,N_315);
or U1429 (N_1429,N_986,N_965);
xor U1430 (N_1430,N_42,N_423);
or U1431 (N_1431,N_723,N_607);
and U1432 (N_1432,N_799,N_188);
nand U1433 (N_1433,N_265,N_466);
or U1434 (N_1434,N_620,N_286);
or U1435 (N_1435,N_477,N_288);
or U1436 (N_1436,N_628,N_988);
and U1437 (N_1437,N_166,N_570);
nor U1438 (N_1438,N_718,N_585);
or U1439 (N_1439,N_479,N_178);
or U1440 (N_1440,N_518,N_392);
or U1441 (N_1441,N_507,N_470);
and U1442 (N_1442,N_498,N_469);
and U1443 (N_1443,N_388,N_15);
nor U1444 (N_1444,N_681,N_854);
nor U1445 (N_1445,N_863,N_632);
nor U1446 (N_1446,N_461,N_365);
nand U1447 (N_1447,N_676,N_409);
nor U1448 (N_1448,N_769,N_245);
and U1449 (N_1449,N_935,N_91);
nand U1450 (N_1450,N_802,N_898);
nor U1451 (N_1451,N_920,N_868);
nand U1452 (N_1452,N_136,N_207);
xnor U1453 (N_1453,N_30,N_159);
xnor U1454 (N_1454,N_654,N_672);
or U1455 (N_1455,N_955,N_144);
nand U1456 (N_1456,N_553,N_481);
or U1457 (N_1457,N_48,N_852);
or U1458 (N_1458,N_567,N_985);
xnor U1459 (N_1459,N_302,N_313);
nor U1460 (N_1460,N_331,N_623);
and U1461 (N_1461,N_726,N_448);
or U1462 (N_1462,N_192,N_184);
xor U1463 (N_1463,N_421,N_851);
or U1464 (N_1464,N_593,N_594);
and U1465 (N_1465,N_266,N_151);
and U1466 (N_1466,N_385,N_427);
and U1467 (N_1467,N_342,N_733);
nor U1468 (N_1468,N_36,N_904);
xnor U1469 (N_1469,N_987,N_972);
xnor U1470 (N_1470,N_788,N_774);
xor U1471 (N_1471,N_636,N_582);
xor U1472 (N_1472,N_790,N_60);
or U1473 (N_1473,N_252,N_174);
xor U1474 (N_1474,N_292,N_890);
nor U1475 (N_1475,N_293,N_319);
and U1476 (N_1476,N_756,N_925);
xnor U1477 (N_1477,N_102,N_83);
and U1478 (N_1478,N_277,N_656);
nor U1479 (N_1479,N_564,N_841);
xnor U1480 (N_1480,N_183,N_825);
xnor U1481 (N_1481,N_199,N_624);
xor U1482 (N_1482,N_951,N_389);
and U1483 (N_1483,N_227,N_303);
and U1484 (N_1484,N_4,N_332);
xnor U1485 (N_1485,N_535,N_956);
xnor U1486 (N_1486,N_271,N_27);
and U1487 (N_1487,N_103,N_120);
nand U1488 (N_1488,N_566,N_701);
or U1489 (N_1489,N_437,N_875);
nor U1490 (N_1490,N_93,N_74);
and U1491 (N_1491,N_914,N_312);
and U1492 (N_1492,N_454,N_59);
xor U1493 (N_1493,N_49,N_901);
xor U1494 (N_1494,N_573,N_420);
and U1495 (N_1495,N_815,N_386);
xnor U1496 (N_1496,N_714,N_874);
or U1497 (N_1497,N_655,N_805);
xor U1498 (N_1498,N_405,N_425);
nor U1499 (N_1499,N_984,N_865);
nand U1500 (N_1500,N_550,N_300);
nor U1501 (N_1501,N_442,N_54);
xnor U1502 (N_1502,N_352,N_452);
or U1503 (N_1503,N_132,N_246);
nor U1504 (N_1504,N_561,N_876);
nor U1505 (N_1505,N_272,N_7);
nor U1506 (N_1506,N_177,N_649);
nor U1507 (N_1507,N_763,N_770);
nor U1508 (N_1508,N_474,N_335);
nor U1509 (N_1509,N_331,N_729);
nand U1510 (N_1510,N_434,N_666);
xnor U1511 (N_1511,N_529,N_588);
or U1512 (N_1512,N_14,N_519);
and U1513 (N_1513,N_775,N_527);
xnor U1514 (N_1514,N_286,N_806);
nor U1515 (N_1515,N_13,N_424);
and U1516 (N_1516,N_124,N_924);
or U1517 (N_1517,N_737,N_627);
nor U1518 (N_1518,N_617,N_794);
xor U1519 (N_1519,N_976,N_160);
xor U1520 (N_1520,N_871,N_716);
xnor U1521 (N_1521,N_97,N_550);
and U1522 (N_1522,N_186,N_234);
nand U1523 (N_1523,N_347,N_857);
xnor U1524 (N_1524,N_652,N_868);
or U1525 (N_1525,N_388,N_202);
and U1526 (N_1526,N_395,N_561);
and U1527 (N_1527,N_820,N_707);
xor U1528 (N_1528,N_167,N_112);
xnor U1529 (N_1529,N_707,N_796);
xor U1530 (N_1530,N_127,N_492);
xor U1531 (N_1531,N_5,N_81);
and U1532 (N_1532,N_425,N_568);
xnor U1533 (N_1533,N_395,N_69);
xor U1534 (N_1534,N_671,N_712);
or U1535 (N_1535,N_297,N_921);
and U1536 (N_1536,N_230,N_876);
nor U1537 (N_1537,N_470,N_120);
nand U1538 (N_1538,N_570,N_162);
nand U1539 (N_1539,N_692,N_411);
nor U1540 (N_1540,N_814,N_453);
nand U1541 (N_1541,N_911,N_161);
or U1542 (N_1542,N_430,N_241);
or U1543 (N_1543,N_161,N_263);
nand U1544 (N_1544,N_415,N_533);
nor U1545 (N_1545,N_872,N_585);
and U1546 (N_1546,N_551,N_323);
and U1547 (N_1547,N_88,N_27);
and U1548 (N_1548,N_636,N_924);
or U1549 (N_1549,N_118,N_546);
nand U1550 (N_1550,N_917,N_17);
nand U1551 (N_1551,N_18,N_646);
nor U1552 (N_1552,N_428,N_481);
and U1553 (N_1553,N_929,N_32);
nor U1554 (N_1554,N_110,N_586);
nor U1555 (N_1555,N_542,N_157);
nor U1556 (N_1556,N_575,N_146);
or U1557 (N_1557,N_0,N_609);
nor U1558 (N_1558,N_963,N_578);
nand U1559 (N_1559,N_56,N_160);
and U1560 (N_1560,N_707,N_675);
or U1561 (N_1561,N_707,N_450);
and U1562 (N_1562,N_450,N_530);
and U1563 (N_1563,N_902,N_65);
xnor U1564 (N_1564,N_405,N_936);
and U1565 (N_1565,N_824,N_423);
xnor U1566 (N_1566,N_974,N_483);
xor U1567 (N_1567,N_955,N_658);
or U1568 (N_1568,N_465,N_982);
xnor U1569 (N_1569,N_235,N_878);
xor U1570 (N_1570,N_410,N_839);
nand U1571 (N_1571,N_212,N_10);
or U1572 (N_1572,N_924,N_815);
xnor U1573 (N_1573,N_368,N_196);
xnor U1574 (N_1574,N_756,N_428);
and U1575 (N_1575,N_502,N_635);
and U1576 (N_1576,N_417,N_480);
nor U1577 (N_1577,N_186,N_260);
nor U1578 (N_1578,N_411,N_773);
or U1579 (N_1579,N_739,N_440);
xor U1580 (N_1580,N_782,N_388);
xnor U1581 (N_1581,N_893,N_670);
or U1582 (N_1582,N_142,N_792);
nor U1583 (N_1583,N_101,N_533);
and U1584 (N_1584,N_315,N_902);
nand U1585 (N_1585,N_100,N_547);
xnor U1586 (N_1586,N_569,N_964);
nand U1587 (N_1587,N_817,N_129);
nor U1588 (N_1588,N_613,N_966);
xor U1589 (N_1589,N_412,N_244);
nor U1590 (N_1590,N_775,N_159);
xor U1591 (N_1591,N_118,N_724);
and U1592 (N_1592,N_528,N_855);
and U1593 (N_1593,N_855,N_635);
nand U1594 (N_1594,N_386,N_310);
or U1595 (N_1595,N_760,N_80);
nor U1596 (N_1596,N_891,N_576);
nor U1597 (N_1597,N_863,N_99);
or U1598 (N_1598,N_752,N_711);
and U1599 (N_1599,N_803,N_107);
or U1600 (N_1600,N_627,N_944);
or U1601 (N_1601,N_289,N_712);
nand U1602 (N_1602,N_134,N_204);
nor U1603 (N_1603,N_95,N_72);
and U1604 (N_1604,N_497,N_136);
nor U1605 (N_1605,N_812,N_834);
nand U1606 (N_1606,N_224,N_41);
nand U1607 (N_1607,N_94,N_680);
and U1608 (N_1608,N_953,N_830);
or U1609 (N_1609,N_721,N_594);
xor U1610 (N_1610,N_733,N_627);
and U1611 (N_1611,N_487,N_216);
nor U1612 (N_1612,N_929,N_194);
nand U1613 (N_1613,N_791,N_28);
xnor U1614 (N_1614,N_337,N_926);
nand U1615 (N_1615,N_544,N_753);
nand U1616 (N_1616,N_862,N_99);
or U1617 (N_1617,N_438,N_554);
nor U1618 (N_1618,N_138,N_161);
xor U1619 (N_1619,N_408,N_15);
nand U1620 (N_1620,N_552,N_198);
xnor U1621 (N_1621,N_69,N_434);
xor U1622 (N_1622,N_733,N_656);
or U1623 (N_1623,N_190,N_800);
or U1624 (N_1624,N_537,N_812);
and U1625 (N_1625,N_975,N_808);
nand U1626 (N_1626,N_393,N_100);
or U1627 (N_1627,N_754,N_140);
nand U1628 (N_1628,N_688,N_215);
nand U1629 (N_1629,N_431,N_35);
nand U1630 (N_1630,N_433,N_316);
nand U1631 (N_1631,N_115,N_694);
xnor U1632 (N_1632,N_425,N_784);
and U1633 (N_1633,N_601,N_243);
or U1634 (N_1634,N_29,N_828);
xor U1635 (N_1635,N_358,N_666);
or U1636 (N_1636,N_103,N_748);
nor U1637 (N_1637,N_703,N_655);
nor U1638 (N_1638,N_469,N_286);
nand U1639 (N_1639,N_297,N_861);
or U1640 (N_1640,N_998,N_738);
or U1641 (N_1641,N_136,N_429);
or U1642 (N_1642,N_4,N_579);
xor U1643 (N_1643,N_970,N_769);
and U1644 (N_1644,N_995,N_741);
nand U1645 (N_1645,N_759,N_873);
nand U1646 (N_1646,N_839,N_604);
xor U1647 (N_1647,N_279,N_850);
nand U1648 (N_1648,N_666,N_893);
nand U1649 (N_1649,N_938,N_854);
and U1650 (N_1650,N_16,N_383);
xnor U1651 (N_1651,N_506,N_934);
xnor U1652 (N_1652,N_252,N_546);
nor U1653 (N_1653,N_249,N_794);
nor U1654 (N_1654,N_66,N_311);
xnor U1655 (N_1655,N_267,N_522);
nand U1656 (N_1656,N_432,N_572);
xnor U1657 (N_1657,N_333,N_446);
nand U1658 (N_1658,N_485,N_973);
nand U1659 (N_1659,N_95,N_931);
and U1660 (N_1660,N_846,N_201);
xor U1661 (N_1661,N_781,N_775);
nor U1662 (N_1662,N_733,N_986);
xor U1663 (N_1663,N_971,N_967);
nand U1664 (N_1664,N_843,N_660);
and U1665 (N_1665,N_722,N_123);
nand U1666 (N_1666,N_838,N_906);
or U1667 (N_1667,N_677,N_205);
and U1668 (N_1668,N_456,N_39);
and U1669 (N_1669,N_886,N_378);
nand U1670 (N_1670,N_807,N_184);
xnor U1671 (N_1671,N_1,N_792);
and U1672 (N_1672,N_593,N_859);
and U1673 (N_1673,N_134,N_156);
nand U1674 (N_1674,N_789,N_311);
nand U1675 (N_1675,N_422,N_124);
and U1676 (N_1676,N_355,N_557);
nor U1677 (N_1677,N_121,N_364);
nand U1678 (N_1678,N_119,N_367);
and U1679 (N_1679,N_384,N_729);
xnor U1680 (N_1680,N_298,N_189);
nor U1681 (N_1681,N_983,N_203);
or U1682 (N_1682,N_105,N_458);
and U1683 (N_1683,N_437,N_979);
nand U1684 (N_1684,N_224,N_510);
nor U1685 (N_1685,N_422,N_338);
nor U1686 (N_1686,N_243,N_716);
and U1687 (N_1687,N_544,N_984);
nand U1688 (N_1688,N_592,N_726);
nand U1689 (N_1689,N_230,N_646);
and U1690 (N_1690,N_771,N_696);
or U1691 (N_1691,N_608,N_231);
xor U1692 (N_1692,N_758,N_458);
nor U1693 (N_1693,N_964,N_458);
nor U1694 (N_1694,N_437,N_179);
xor U1695 (N_1695,N_102,N_235);
or U1696 (N_1696,N_389,N_304);
and U1697 (N_1697,N_496,N_126);
or U1698 (N_1698,N_979,N_387);
and U1699 (N_1699,N_641,N_156);
nand U1700 (N_1700,N_205,N_820);
nor U1701 (N_1701,N_647,N_406);
nand U1702 (N_1702,N_311,N_142);
and U1703 (N_1703,N_45,N_270);
nand U1704 (N_1704,N_531,N_977);
or U1705 (N_1705,N_351,N_117);
or U1706 (N_1706,N_440,N_686);
nor U1707 (N_1707,N_995,N_563);
and U1708 (N_1708,N_334,N_551);
xor U1709 (N_1709,N_302,N_903);
nand U1710 (N_1710,N_223,N_262);
or U1711 (N_1711,N_5,N_342);
nand U1712 (N_1712,N_532,N_356);
nand U1713 (N_1713,N_872,N_856);
or U1714 (N_1714,N_764,N_584);
and U1715 (N_1715,N_627,N_3);
or U1716 (N_1716,N_747,N_435);
nor U1717 (N_1717,N_855,N_780);
nand U1718 (N_1718,N_93,N_165);
or U1719 (N_1719,N_140,N_949);
nor U1720 (N_1720,N_955,N_921);
xor U1721 (N_1721,N_674,N_139);
nor U1722 (N_1722,N_727,N_943);
nand U1723 (N_1723,N_175,N_513);
xnor U1724 (N_1724,N_906,N_600);
nand U1725 (N_1725,N_258,N_358);
xor U1726 (N_1726,N_937,N_988);
nor U1727 (N_1727,N_998,N_51);
xor U1728 (N_1728,N_587,N_912);
and U1729 (N_1729,N_95,N_290);
or U1730 (N_1730,N_525,N_604);
or U1731 (N_1731,N_876,N_911);
xor U1732 (N_1732,N_939,N_515);
nand U1733 (N_1733,N_707,N_22);
or U1734 (N_1734,N_615,N_503);
nor U1735 (N_1735,N_416,N_732);
nand U1736 (N_1736,N_507,N_796);
or U1737 (N_1737,N_833,N_427);
or U1738 (N_1738,N_339,N_566);
and U1739 (N_1739,N_630,N_436);
xor U1740 (N_1740,N_226,N_268);
xnor U1741 (N_1741,N_857,N_36);
nor U1742 (N_1742,N_480,N_995);
or U1743 (N_1743,N_268,N_983);
nor U1744 (N_1744,N_829,N_851);
and U1745 (N_1745,N_48,N_684);
nand U1746 (N_1746,N_210,N_225);
nand U1747 (N_1747,N_268,N_670);
or U1748 (N_1748,N_283,N_534);
nand U1749 (N_1749,N_347,N_269);
or U1750 (N_1750,N_784,N_685);
and U1751 (N_1751,N_799,N_555);
nand U1752 (N_1752,N_232,N_217);
nand U1753 (N_1753,N_406,N_254);
xor U1754 (N_1754,N_72,N_806);
and U1755 (N_1755,N_453,N_788);
and U1756 (N_1756,N_728,N_218);
nand U1757 (N_1757,N_196,N_566);
xnor U1758 (N_1758,N_207,N_504);
or U1759 (N_1759,N_711,N_997);
xnor U1760 (N_1760,N_300,N_707);
and U1761 (N_1761,N_354,N_405);
or U1762 (N_1762,N_191,N_509);
nor U1763 (N_1763,N_634,N_269);
nand U1764 (N_1764,N_976,N_305);
nor U1765 (N_1765,N_901,N_73);
and U1766 (N_1766,N_255,N_152);
and U1767 (N_1767,N_832,N_85);
nor U1768 (N_1768,N_595,N_289);
and U1769 (N_1769,N_358,N_958);
or U1770 (N_1770,N_456,N_628);
nor U1771 (N_1771,N_700,N_807);
or U1772 (N_1772,N_82,N_68);
xnor U1773 (N_1773,N_931,N_38);
xnor U1774 (N_1774,N_917,N_480);
nand U1775 (N_1775,N_44,N_903);
nand U1776 (N_1776,N_383,N_440);
xnor U1777 (N_1777,N_516,N_380);
nand U1778 (N_1778,N_905,N_96);
nand U1779 (N_1779,N_686,N_297);
nand U1780 (N_1780,N_203,N_878);
or U1781 (N_1781,N_983,N_14);
or U1782 (N_1782,N_591,N_359);
nor U1783 (N_1783,N_559,N_369);
nand U1784 (N_1784,N_760,N_341);
xor U1785 (N_1785,N_13,N_683);
and U1786 (N_1786,N_41,N_186);
and U1787 (N_1787,N_674,N_22);
xnor U1788 (N_1788,N_185,N_50);
nand U1789 (N_1789,N_399,N_25);
nor U1790 (N_1790,N_157,N_252);
xnor U1791 (N_1791,N_605,N_589);
or U1792 (N_1792,N_371,N_279);
or U1793 (N_1793,N_258,N_173);
or U1794 (N_1794,N_578,N_863);
nor U1795 (N_1795,N_925,N_598);
or U1796 (N_1796,N_851,N_341);
xor U1797 (N_1797,N_672,N_20);
or U1798 (N_1798,N_399,N_189);
or U1799 (N_1799,N_785,N_403);
nand U1800 (N_1800,N_935,N_274);
nand U1801 (N_1801,N_184,N_156);
or U1802 (N_1802,N_515,N_10);
or U1803 (N_1803,N_446,N_147);
or U1804 (N_1804,N_450,N_938);
xnor U1805 (N_1805,N_945,N_947);
nor U1806 (N_1806,N_194,N_726);
or U1807 (N_1807,N_459,N_53);
nand U1808 (N_1808,N_465,N_728);
or U1809 (N_1809,N_26,N_933);
nand U1810 (N_1810,N_546,N_83);
xnor U1811 (N_1811,N_477,N_94);
nand U1812 (N_1812,N_286,N_473);
and U1813 (N_1813,N_607,N_849);
and U1814 (N_1814,N_402,N_797);
nand U1815 (N_1815,N_124,N_211);
nor U1816 (N_1816,N_451,N_614);
and U1817 (N_1817,N_528,N_755);
xnor U1818 (N_1818,N_997,N_220);
or U1819 (N_1819,N_318,N_726);
and U1820 (N_1820,N_551,N_279);
nand U1821 (N_1821,N_155,N_7);
xnor U1822 (N_1822,N_507,N_381);
nor U1823 (N_1823,N_853,N_761);
and U1824 (N_1824,N_445,N_449);
xor U1825 (N_1825,N_283,N_778);
and U1826 (N_1826,N_238,N_580);
and U1827 (N_1827,N_171,N_222);
and U1828 (N_1828,N_458,N_808);
nand U1829 (N_1829,N_398,N_206);
xor U1830 (N_1830,N_867,N_675);
nor U1831 (N_1831,N_757,N_54);
or U1832 (N_1832,N_831,N_403);
and U1833 (N_1833,N_904,N_613);
and U1834 (N_1834,N_983,N_469);
nand U1835 (N_1835,N_268,N_660);
xor U1836 (N_1836,N_513,N_856);
and U1837 (N_1837,N_626,N_750);
xnor U1838 (N_1838,N_456,N_485);
xnor U1839 (N_1839,N_472,N_877);
and U1840 (N_1840,N_69,N_694);
and U1841 (N_1841,N_210,N_245);
xnor U1842 (N_1842,N_878,N_93);
and U1843 (N_1843,N_710,N_25);
xor U1844 (N_1844,N_593,N_804);
and U1845 (N_1845,N_784,N_637);
nand U1846 (N_1846,N_527,N_170);
and U1847 (N_1847,N_665,N_746);
nor U1848 (N_1848,N_959,N_837);
and U1849 (N_1849,N_132,N_637);
xor U1850 (N_1850,N_664,N_612);
xnor U1851 (N_1851,N_507,N_784);
nand U1852 (N_1852,N_247,N_778);
xnor U1853 (N_1853,N_537,N_621);
or U1854 (N_1854,N_879,N_333);
nand U1855 (N_1855,N_650,N_372);
or U1856 (N_1856,N_919,N_262);
and U1857 (N_1857,N_735,N_938);
and U1858 (N_1858,N_394,N_191);
and U1859 (N_1859,N_649,N_668);
or U1860 (N_1860,N_987,N_346);
nor U1861 (N_1861,N_718,N_609);
xnor U1862 (N_1862,N_792,N_738);
xnor U1863 (N_1863,N_820,N_334);
xnor U1864 (N_1864,N_906,N_57);
and U1865 (N_1865,N_371,N_519);
or U1866 (N_1866,N_203,N_582);
and U1867 (N_1867,N_226,N_782);
xnor U1868 (N_1868,N_362,N_325);
xor U1869 (N_1869,N_71,N_317);
xor U1870 (N_1870,N_657,N_508);
nor U1871 (N_1871,N_966,N_298);
and U1872 (N_1872,N_573,N_160);
nor U1873 (N_1873,N_244,N_254);
or U1874 (N_1874,N_131,N_35);
or U1875 (N_1875,N_854,N_133);
and U1876 (N_1876,N_599,N_76);
and U1877 (N_1877,N_12,N_913);
or U1878 (N_1878,N_321,N_491);
nand U1879 (N_1879,N_865,N_382);
and U1880 (N_1880,N_602,N_319);
nand U1881 (N_1881,N_450,N_661);
and U1882 (N_1882,N_682,N_943);
xor U1883 (N_1883,N_482,N_832);
and U1884 (N_1884,N_841,N_755);
xnor U1885 (N_1885,N_606,N_453);
nor U1886 (N_1886,N_939,N_925);
nor U1887 (N_1887,N_380,N_394);
and U1888 (N_1888,N_921,N_670);
nor U1889 (N_1889,N_613,N_111);
nor U1890 (N_1890,N_657,N_650);
xnor U1891 (N_1891,N_93,N_528);
and U1892 (N_1892,N_118,N_418);
and U1893 (N_1893,N_821,N_101);
and U1894 (N_1894,N_921,N_958);
xor U1895 (N_1895,N_871,N_724);
nand U1896 (N_1896,N_341,N_319);
xnor U1897 (N_1897,N_385,N_851);
nor U1898 (N_1898,N_377,N_380);
and U1899 (N_1899,N_771,N_79);
nor U1900 (N_1900,N_988,N_478);
or U1901 (N_1901,N_70,N_164);
nand U1902 (N_1902,N_798,N_598);
nor U1903 (N_1903,N_752,N_664);
or U1904 (N_1904,N_401,N_326);
or U1905 (N_1905,N_416,N_616);
nand U1906 (N_1906,N_310,N_373);
and U1907 (N_1907,N_905,N_637);
nand U1908 (N_1908,N_457,N_397);
and U1909 (N_1909,N_479,N_728);
or U1910 (N_1910,N_321,N_417);
nand U1911 (N_1911,N_597,N_398);
and U1912 (N_1912,N_494,N_153);
nor U1913 (N_1913,N_496,N_67);
nor U1914 (N_1914,N_468,N_365);
nand U1915 (N_1915,N_57,N_790);
or U1916 (N_1916,N_853,N_288);
nor U1917 (N_1917,N_590,N_574);
and U1918 (N_1918,N_380,N_392);
nand U1919 (N_1919,N_353,N_26);
or U1920 (N_1920,N_711,N_996);
and U1921 (N_1921,N_710,N_358);
xnor U1922 (N_1922,N_84,N_739);
xnor U1923 (N_1923,N_813,N_11);
xor U1924 (N_1924,N_70,N_615);
xnor U1925 (N_1925,N_292,N_750);
and U1926 (N_1926,N_931,N_732);
or U1927 (N_1927,N_870,N_293);
nand U1928 (N_1928,N_413,N_209);
nor U1929 (N_1929,N_630,N_505);
nor U1930 (N_1930,N_800,N_708);
xnor U1931 (N_1931,N_724,N_739);
xnor U1932 (N_1932,N_181,N_497);
nor U1933 (N_1933,N_837,N_47);
nor U1934 (N_1934,N_668,N_64);
xor U1935 (N_1935,N_555,N_851);
nand U1936 (N_1936,N_580,N_246);
nand U1937 (N_1937,N_747,N_334);
xor U1938 (N_1938,N_21,N_847);
nor U1939 (N_1939,N_206,N_879);
and U1940 (N_1940,N_43,N_514);
or U1941 (N_1941,N_759,N_932);
nand U1942 (N_1942,N_360,N_124);
nand U1943 (N_1943,N_446,N_41);
nand U1944 (N_1944,N_830,N_79);
xnor U1945 (N_1945,N_738,N_635);
and U1946 (N_1946,N_60,N_639);
xor U1947 (N_1947,N_680,N_338);
nand U1948 (N_1948,N_466,N_223);
or U1949 (N_1949,N_229,N_882);
or U1950 (N_1950,N_618,N_763);
and U1951 (N_1951,N_619,N_672);
nand U1952 (N_1952,N_38,N_917);
xor U1953 (N_1953,N_389,N_839);
and U1954 (N_1954,N_3,N_278);
nor U1955 (N_1955,N_63,N_983);
or U1956 (N_1956,N_837,N_763);
nor U1957 (N_1957,N_487,N_133);
xor U1958 (N_1958,N_241,N_871);
and U1959 (N_1959,N_744,N_687);
nand U1960 (N_1960,N_163,N_47);
or U1961 (N_1961,N_577,N_453);
nor U1962 (N_1962,N_289,N_466);
and U1963 (N_1963,N_812,N_103);
nor U1964 (N_1964,N_793,N_316);
nand U1965 (N_1965,N_849,N_93);
nand U1966 (N_1966,N_162,N_85);
xor U1967 (N_1967,N_994,N_287);
or U1968 (N_1968,N_48,N_410);
and U1969 (N_1969,N_85,N_56);
xor U1970 (N_1970,N_989,N_777);
or U1971 (N_1971,N_214,N_310);
nor U1972 (N_1972,N_854,N_164);
and U1973 (N_1973,N_792,N_310);
xor U1974 (N_1974,N_623,N_373);
or U1975 (N_1975,N_564,N_90);
nand U1976 (N_1976,N_61,N_699);
xor U1977 (N_1977,N_798,N_655);
nand U1978 (N_1978,N_645,N_102);
xor U1979 (N_1979,N_32,N_74);
xor U1980 (N_1980,N_665,N_686);
nor U1981 (N_1981,N_793,N_426);
nor U1982 (N_1982,N_837,N_329);
xor U1983 (N_1983,N_494,N_484);
nor U1984 (N_1984,N_629,N_347);
and U1985 (N_1985,N_890,N_394);
nor U1986 (N_1986,N_778,N_576);
or U1987 (N_1987,N_161,N_727);
xnor U1988 (N_1988,N_571,N_258);
nor U1989 (N_1989,N_775,N_618);
xor U1990 (N_1990,N_689,N_518);
or U1991 (N_1991,N_45,N_118);
and U1992 (N_1992,N_345,N_86);
xor U1993 (N_1993,N_710,N_410);
nand U1994 (N_1994,N_162,N_720);
xnor U1995 (N_1995,N_91,N_14);
or U1996 (N_1996,N_721,N_927);
nand U1997 (N_1997,N_36,N_834);
nor U1998 (N_1998,N_721,N_412);
or U1999 (N_1999,N_812,N_89);
and U2000 (N_2000,N_1887,N_1493);
nor U2001 (N_2001,N_1741,N_1667);
xor U2002 (N_2002,N_1475,N_1484);
or U2003 (N_2003,N_1432,N_1967);
or U2004 (N_2004,N_1441,N_1610);
xor U2005 (N_2005,N_1474,N_1378);
nand U2006 (N_2006,N_1770,N_1899);
nor U2007 (N_2007,N_1535,N_1628);
nor U2008 (N_2008,N_1406,N_1306);
xor U2009 (N_2009,N_1212,N_1750);
nand U2010 (N_2010,N_1897,N_1877);
or U2011 (N_2011,N_1332,N_1532);
xor U2012 (N_2012,N_1708,N_1066);
nor U2013 (N_2013,N_1629,N_1787);
nor U2014 (N_2014,N_1419,N_1187);
or U2015 (N_2015,N_1883,N_1876);
xor U2016 (N_2016,N_1706,N_1530);
xor U2017 (N_2017,N_1505,N_1926);
nor U2018 (N_2018,N_1684,N_1573);
or U2019 (N_2019,N_1796,N_1941);
nand U2020 (N_2020,N_1570,N_1117);
nor U2021 (N_2021,N_1330,N_1756);
nor U2022 (N_2022,N_1546,N_1590);
nor U2023 (N_2023,N_1416,N_1291);
or U2024 (N_2024,N_1646,N_1295);
nand U2025 (N_2025,N_1501,N_1140);
and U2026 (N_2026,N_1259,N_1184);
or U2027 (N_2027,N_1367,N_1659);
nor U2028 (N_2028,N_1949,N_1278);
or U2029 (N_2029,N_1625,N_1989);
and U2030 (N_2030,N_1359,N_1286);
and U2031 (N_2031,N_1845,N_1404);
and U2032 (N_2032,N_1614,N_1998);
and U2033 (N_2033,N_1107,N_1634);
or U2034 (N_2034,N_1267,N_1285);
nor U2035 (N_2035,N_1736,N_1690);
or U2036 (N_2036,N_1049,N_1992);
xnor U2037 (N_2037,N_1930,N_1450);
xor U2038 (N_2038,N_1811,N_1743);
nor U2039 (N_2039,N_1551,N_1592);
or U2040 (N_2040,N_1601,N_1520);
or U2041 (N_2041,N_1084,N_1409);
xor U2042 (N_2042,N_1898,N_1950);
nor U2043 (N_2043,N_1124,N_1793);
or U2044 (N_2044,N_1673,N_1995);
nand U2045 (N_2045,N_1933,N_1449);
nand U2046 (N_2046,N_1408,N_1759);
or U2047 (N_2047,N_1376,N_1622);
or U2048 (N_2048,N_1670,N_1913);
nand U2049 (N_2049,N_1236,N_1361);
xnor U2050 (N_2050,N_1269,N_1348);
xor U2051 (N_2051,N_1808,N_1956);
xor U2052 (N_2052,N_1082,N_1166);
and U2053 (N_2053,N_1645,N_1446);
nor U2054 (N_2054,N_1412,N_1313);
nor U2055 (N_2055,N_1963,N_1307);
xnor U2056 (N_2056,N_1296,N_1241);
and U2057 (N_2057,N_1596,N_1973);
or U2058 (N_2058,N_1886,N_1232);
or U2059 (N_2059,N_1215,N_1487);
xnor U2060 (N_2060,N_1794,N_1397);
nand U2061 (N_2061,N_1068,N_1746);
nor U2062 (N_2062,N_1867,N_1856);
nand U2063 (N_2063,N_1960,N_1198);
nand U2064 (N_2064,N_1597,N_1315);
or U2065 (N_2065,N_1586,N_1025);
nor U2066 (N_2066,N_1022,N_1067);
xnor U2067 (N_2067,N_1885,N_1693);
xor U2068 (N_2068,N_1060,N_1948);
or U2069 (N_2069,N_1177,N_1439);
xnor U2070 (N_2070,N_1909,N_1627);
xnor U2071 (N_2071,N_1402,N_1220);
nand U2072 (N_2072,N_1511,N_1425);
nor U2073 (N_2073,N_1577,N_1228);
and U2074 (N_2074,N_1213,N_1040);
and U2075 (N_2075,N_1660,N_1059);
or U2076 (N_2076,N_1704,N_1410);
nor U2077 (N_2077,N_1012,N_1105);
xor U2078 (N_2078,N_1769,N_1422);
or U2079 (N_2079,N_1339,N_1118);
nor U2080 (N_2080,N_1097,N_1130);
or U2081 (N_2081,N_1906,N_1418);
nor U2082 (N_2082,N_1093,N_1942);
or U2083 (N_2083,N_1765,N_1245);
nor U2084 (N_2084,N_1002,N_1832);
and U2085 (N_2085,N_1462,N_1128);
and U2086 (N_2086,N_1823,N_1932);
and U2087 (N_2087,N_1078,N_1202);
nand U2088 (N_2088,N_1635,N_1112);
nand U2089 (N_2089,N_1043,N_1063);
or U2090 (N_2090,N_1677,N_1194);
xor U2091 (N_2091,N_1133,N_1185);
nor U2092 (N_2092,N_1672,N_1777);
nor U2093 (N_2093,N_1509,N_1862);
nand U2094 (N_2094,N_1749,N_1261);
or U2095 (N_2095,N_1700,N_1533);
nor U2096 (N_2096,N_1553,N_1141);
or U2097 (N_2097,N_1587,N_1004);
xor U2098 (N_2098,N_1195,N_1694);
or U2099 (N_2099,N_1248,N_1270);
xnor U2100 (N_2100,N_1497,N_1606);
and U2101 (N_2101,N_1683,N_1090);
and U2102 (N_2102,N_1905,N_1954);
xnor U2103 (N_2103,N_1934,N_1287);
or U2104 (N_2104,N_1781,N_1009);
and U2105 (N_2105,N_1007,N_1768);
or U2106 (N_2106,N_1256,N_1400);
and U2107 (N_2107,N_1035,N_1020);
nor U2108 (N_2108,N_1846,N_1653);
and U2109 (N_2109,N_1253,N_1340);
nand U2110 (N_2110,N_1583,N_1156);
xnor U2111 (N_2111,N_1921,N_1051);
and U2112 (N_2112,N_1154,N_1952);
xor U2113 (N_2113,N_1526,N_1303);
or U2114 (N_2114,N_1208,N_1196);
or U2115 (N_2115,N_1804,N_1589);
and U2116 (N_2116,N_1486,N_1254);
xnor U2117 (N_2117,N_1103,N_1438);
or U2118 (N_2118,N_1807,N_1502);
xnor U2119 (N_2119,N_1150,N_1182);
or U2120 (N_2120,N_1473,N_1901);
and U2121 (N_2121,N_1203,N_1356);
xor U2122 (N_2122,N_1783,N_1233);
nor U2123 (N_2123,N_1041,N_1516);
nand U2124 (N_2124,N_1802,N_1753);
nand U2125 (N_2125,N_1000,N_1758);
xor U2126 (N_2126,N_1797,N_1556);
xor U2127 (N_2127,N_1541,N_1938);
and U2128 (N_2128,N_1210,N_1651);
nand U2129 (N_2129,N_1776,N_1585);
nor U2130 (N_2130,N_1874,N_1873);
nor U2131 (N_2131,N_1944,N_1172);
or U2132 (N_2132,N_1352,N_1120);
nor U2133 (N_2133,N_1958,N_1461);
nor U2134 (N_2134,N_1737,N_1837);
xor U2135 (N_2135,N_1679,N_1292);
xnor U2136 (N_2136,N_1388,N_1274);
nor U2137 (N_2137,N_1735,N_1987);
nor U2138 (N_2138,N_1917,N_1578);
nor U2139 (N_2139,N_1310,N_1841);
xnor U2140 (N_2140,N_1317,N_1994);
xor U2141 (N_2141,N_1016,N_1231);
nor U2142 (N_2142,N_1642,N_1031);
and U2143 (N_2143,N_1908,N_1222);
and U2144 (N_2144,N_1162,N_1483);
xnor U2145 (N_2145,N_1631,N_1716);
nor U2146 (N_2146,N_1563,N_1293);
or U2147 (N_2147,N_1174,N_1600);
nor U2148 (N_2148,N_1861,N_1658);
nor U2149 (N_2149,N_1544,N_1143);
and U2150 (N_2150,N_1834,N_1073);
xor U2151 (N_2151,N_1146,N_1676);
xnor U2152 (N_2152,N_1572,N_1365);
nand U2153 (N_2153,N_1358,N_1003);
or U2154 (N_2154,N_1545,N_1104);
xor U2155 (N_2155,N_1386,N_1217);
and U2156 (N_2156,N_1347,N_1255);
or U2157 (N_2157,N_1817,N_1984);
or U2158 (N_2158,N_1054,N_1978);
nor U2159 (N_2159,N_1852,N_1246);
nor U2160 (N_2160,N_1844,N_1454);
xor U2161 (N_2161,N_1393,N_1273);
nor U2162 (N_2162,N_1403,N_1380);
nor U2163 (N_2163,N_1430,N_1214);
xor U2164 (N_2164,N_1453,N_1966);
nand U2165 (N_2165,N_1763,N_1875);
nor U2166 (N_2166,N_1053,N_1478);
or U2167 (N_2167,N_1311,N_1440);
or U2168 (N_2168,N_1263,N_1703);
and U2169 (N_2169,N_1641,N_1519);
nand U2170 (N_2170,N_1757,N_1464);
nor U2171 (N_2171,N_1223,N_1385);
nand U2172 (N_2172,N_1827,N_1689);
nand U2173 (N_2173,N_1218,N_1580);
nor U2174 (N_2174,N_1072,N_1711);
nand U2175 (N_2175,N_1924,N_1224);
nor U2176 (N_2176,N_1163,N_1329);
and U2177 (N_2177,N_1458,N_1316);
nand U2178 (N_2178,N_1126,N_1387);
and U2179 (N_2179,N_1648,N_1742);
and U2180 (N_2180,N_1148,N_1970);
xor U2181 (N_2181,N_1615,N_1238);
or U2182 (N_2182,N_1021,N_1109);
nand U2183 (N_2183,N_1904,N_1325);
nand U2184 (N_2184,N_1680,N_1980);
nor U2185 (N_2185,N_1319,N_1001);
and U2186 (N_2186,N_1019,N_1713);
and U2187 (N_2187,N_1032,N_1131);
and U2188 (N_2188,N_1034,N_1395);
and U2189 (N_2189,N_1153,N_1803);
xor U2190 (N_2190,N_1328,N_1023);
nor U2191 (N_2191,N_1671,N_1106);
xnor U2192 (N_2192,N_1122,N_1854);
xnor U2193 (N_2193,N_1160,N_1552);
xor U2194 (N_2194,N_1363,N_1108);
or U2195 (N_2195,N_1571,N_1857);
nor U2196 (N_2196,N_1565,N_1086);
nor U2197 (N_2197,N_1165,N_1528);
and U2198 (N_2198,N_1014,N_1939);
or U2199 (N_2199,N_1968,N_1953);
xor U2200 (N_2200,N_1981,N_1907);
nor U2201 (N_2201,N_1624,N_1279);
nor U2202 (N_2202,N_1836,N_1975);
nor U2203 (N_2203,N_1864,N_1152);
nand U2204 (N_2204,N_1959,N_1969);
and U2205 (N_2205,N_1420,N_1180);
or U2206 (N_2206,N_1529,N_1824);
xnor U2207 (N_2207,N_1161,N_1173);
nor U2208 (N_2208,N_1943,N_1335);
nor U2209 (N_2209,N_1575,N_1445);
and U2210 (N_2210,N_1448,N_1865);
or U2211 (N_2211,N_1494,N_1850);
or U2212 (N_2212,N_1351,N_1434);
xnor U2213 (N_2213,N_1476,N_1209);
xor U2214 (N_2214,N_1452,N_1705);
or U2215 (N_2215,N_1879,N_1423);
xor U2216 (N_2216,N_1721,N_1201);
nor U2217 (N_2217,N_1472,N_1566);
nand U2218 (N_2218,N_1134,N_1633);
nand U2219 (N_2219,N_1536,N_1373);
xnor U2220 (N_2220,N_1755,N_1559);
nor U2221 (N_2221,N_1136,N_1499);
nand U2222 (N_2222,N_1788,N_1115);
or U2223 (N_2223,N_1028,N_1186);
nor U2224 (N_2224,N_1123,N_1164);
nor U2225 (N_2225,N_1355,N_1243);
nand U2226 (N_2226,N_1221,N_1518);
or U2227 (N_2227,N_1427,N_1192);
and U2228 (N_2228,N_1691,N_1888);
nor U2229 (N_2229,N_1647,N_1979);
and U2230 (N_2230,N_1595,N_1436);
nand U2231 (N_2231,N_1983,N_1927);
xor U2232 (N_2232,N_1900,N_1377);
nand U2233 (N_2233,N_1961,N_1849);
xnor U2234 (N_2234,N_1923,N_1534);
and U2235 (N_2235,N_1613,N_1451);
and U2236 (N_2236,N_1816,N_1251);
nor U2237 (N_2237,N_1181,N_1819);
nand U2238 (N_2238,N_1076,N_1539);
nor U2239 (N_2239,N_1678,N_1695);
nor U2240 (N_2240,N_1853,N_1620);
nor U2241 (N_2241,N_1304,N_1460);
and U2242 (N_2242,N_1492,N_1142);
or U2243 (N_2243,N_1760,N_1280);
nor U2244 (N_2244,N_1542,N_1345);
nand U2245 (N_2245,N_1798,N_1785);
nor U2246 (N_2246,N_1780,N_1398);
and U2247 (N_2247,N_1752,N_1723);
or U2248 (N_2248,N_1443,N_1096);
and U2249 (N_2249,N_1955,N_1264);
and U2250 (N_2250,N_1047,N_1155);
and U2251 (N_2251,N_1982,N_1940);
nor U2252 (N_2252,N_1537,N_1290);
xor U2253 (N_2253,N_1974,N_1276);
nor U2254 (N_2254,N_1971,N_1362);
and U2255 (N_2255,N_1698,N_1421);
or U2256 (N_2256,N_1297,N_1724);
xor U2257 (N_2257,N_1603,N_1190);
or U2258 (N_2258,N_1080,N_1379);
nand U2259 (N_2259,N_1301,N_1230);
nand U2260 (N_2260,N_1821,N_1730);
xnor U2261 (N_2261,N_1892,N_1343);
and U2262 (N_2262,N_1922,N_1838);
and U2263 (N_2263,N_1814,N_1878);
nor U2264 (N_2264,N_1822,N_1557);
or U2265 (N_2265,N_1851,N_1341);
nand U2266 (N_2266,N_1947,N_1384);
xnor U2267 (N_2267,N_1320,N_1829);
or U2268 (N_2268,N_1074,N_1401);
nand U2269 (N_2269,N_1789,N_1331);
nand U2270 (N_2270,N_1262,N_1026);
or U2271 (N_2271,N_1030,N_1717);
nor U2272 (N_2272,N_1588,N_1169);
xnor U2273 (N_2273,N_1866,N_1119);
nand U2274 (N_2274,N_1881,N_1644);
xor U2275 (N_2275,N_1976,N_1091);
and U2276 (N_2276,N_1626,N_1810);
nand U2277 (N_2277,N_1158,N_1986);
and U2278 (N_2278,N_1413,N_1847);
or U2279 (N_2279,N_1479,N_1496);
or U2280 (N_2280,N_1687,N_1099);
xnor U2281 (N_2281,N_1271,N_1206);
and U2282 (N_2282,N_1411,N_1444);
nor U2283 (N_2283,N_1521,N_1372);
and U2284 (N_2284,N_1069,N_1751);
nor U2285 (N_2285,N_1548,N_1465);
and U2286 (N_2286,N_1715,N_1733);
or U2287 (N_2287,N_1268,N_1540);
nor U2288 (N_2288,N_1092,N_1349);
nand U2289 (N_2289,N_1931,N_1058);
xor U2290 (N_2290,N_1965,N_1782);
and U2291 (N_2291,N_1524,N_1481);
nand U2292 (N_2292,N_1985,N_1281);
nor U2293 (N_2293,N_1795,N_1191);
or U2294 (N_2294,N_1820,N_1294);
or U2295 (N_2295,N_1506,N_1480);
xnor U2296 (N_2296,N_1747,N_1490);
or U2297 (N_2297,N_1726,N_1719);
nor U2298 (N_2298,N_1071,N_1636);
nand U2299 (N_2299,N_1350,N_1889);
or U2300 (N_2300,N_1662,N_1692);
nand U2301 (N_2301,N_1801,N_1249);
and U2302 (N_2302,N_1065,N_1050);
and U2303 (N_2303,N_1972,N_1247);
or U2304 (N_2304,N_1562,N_1116);
nand U2305 (N_2305,N_1013,N_1664);
or U2306 (N_2306,N_1951,N_1786);
nand U2307 (N_2307,N_1655,N_1110);
or U2308 (N_2308,N_1561,N_1175);
and U2309 (N_2309,N_1178,N_1669);
nor U2310 (N_2310,N_1024,N_1707);
and U2311 (N_2311,N_1712,N_1284);
nor U2312 (N_2312,N_1568,N_1812);
nor U2313 (N_2313,N_1946,N_1010);
xnor U2314 (N_2314,N_1179,N_1630);
xor U2315 (N_2315,N_1792,N_1079);
and U2316 (N_2316,N_1504,N_1468);
nor U2317 (N_2317,N_1729,N_1991);
or U2318 (N_2318,N_1869,N_1127);
nand U2319 (N_2319,N_1652,N_1237);
nor U2320 (N_2320,N_1993,N_1697);
nand U2321 (N_2321,N_1925,N_1144);
or U2322 (N_2322,N_1265,N_1722);
and U2323 (N_2323,N_1895,N_1621);
xor U2324 (N_2324,N_1375,N_1015);
nor U2325 (N_2325,N_1366,N_1455);
and U2326 (N_2326,N_1560,N_1369);
nand U2327 (N_2327,N_1738,N_1466);
xor U2328 (N_2328,N_1574,N_1999);
or U2329 (N_2329,N_1207,N_1396);
nand U2330 (N_2330,N_1346,N_1353);
nand U2331 (N_2331,N_1714,N_1381);
nand U2332 (N_2332,N_1517,N_1945);
nand U2333 (N_2333,N_1197,N_1048);
nand U2334 (N_2334,N_1157,N_1370);
nor U2335 (N_2335,N_1205,N_1391);
and U2336 (N_2336,N_1159,N_1818);
nand U2337 (N_2337,N_1064,N_1042);
xor U2338 (N_2338,N_1342,N_1593);
xnor U2339 (N_2339,N_1863,N_1477);
nor U2340 (N_2340,N_1088,N_1772);
and U2341 (N_2341,N_1732,N_1008);
nand U2342 (N_2342,N_1102,N_1428);
or U2343 (N_2343,N_1299,N_1338);
and U2344 (N_2344,N_1594,N_1188);
and U2345 (N_2345,N_1790,N_1579);
and U2346 (N_2346,N_1168,N_1326);
and U2347 (N_2347,N_1011,N_1305);
nor U2348 (N_2348,N_1919,N_1761);
or U2349 (N_2349,N_1129,N_1200);
nor U2350 (N_2350,N_1139,N_1211);
nand U2351 (N_2351,N_1368,N_1006);
nand U2352 (N_2352,N_1283,N_1489);
or U2353 (N_2353,N_1469,N_1607);
xnor U2354 (N_2354,N_1145,N_1360);
nand U2355 (N_2355,N_1426,N_1773);
xor U2356 (N_2356,N_1855,N_1833);
nand U2357 (N_2357,N_1137,N_1503);
xor U2358 (N_2358,N_1914,N_1550);
and U2359 (N_2359,N_1514,N_1216);
nand U2360 (N_2360,N_1649,N_1848);
nor U2361 (N_2361,N_1219,N_1928);
nand U2362 (N_2362,N_1061,N_1056);
or U2363 (N_2363,N_1062,N_1605);
xnor U2364 (N_2364,N_1498,N_1429);
nor U2365 (N_2365,N_1962,N_1657);
or U2366 (N_2366,N_1623,N_1882);
xor U2367 (N_2367,N_1800,N_1744);
nor U2368 (N_2368,N_1766,N_1831);
or U2369 (N_2369,N_1858,N_1675);
and U2370 (N_2370,N_1725,N_1229);
xnor U2371 (N_2371,N_1235,N_1070);
xnor U2372 (N_2372,N_1903,N_1656);
nand U2373 (N_2373,N_1643,N_1513);
nor U2374 (N_2374,N_1151,N_1915);
nand U2375 (N_2375,N_1463,N_1027);
and U2376 (N_2376,N_1567,N_1260);
nor U2377 (N_2377,N_1809,N_1609);
xor U2378 (N_2378,N_1558,N_1244);
nand U2379 (N_2379,N_1132,N_1718);
and U2380 (N_2380,N_1531,N_1300);
nand U2381 (N_2381,N_1839,N_1910);
and U2382 (N_2382,N_1522,N_1762);
and U2383 (N_2383,N_1791,N_1005);
xnor U2384 (N_2384,N_1323,N_1147);
and U2385 (N_2385,N_1696,N_1916);
xor U2386 (N_2386,N_1257,N_1665);
or U2387 (N_2387,N_1666,N_1170);
or U2388 (N_2388,N_1239,N_1616);
xor U2389 (N_2389,N_1599,N_1618);
nor U2390 (N_2390,N_1392,N_1988);
xor U2391 (N_2391,N_1549,N_1471);
nor U2392 (N_2392,N_1891,N_1602);
and U2393 (N_2393,N_1842,N_1417);
xor U2394 (N_2394,N_1884,N_1394);
nor U2395 (N_2395,N_1495,N_1470);
or U2396 (N_2396,N_1569,N_1227);
nor U2397 (N_2397,N_1997,N_1491);
or U2398 (N_2398,N_1674,N_1250);
and U2399 (N_2399,N_1407,N_1488);
or U2400 (N_2400,N_1564,N_1324);
xnor U2401 (N_2401,N_1859,N_1668);
and U2402 (N_2402,N_1523,N_1456);
xor U2403 (N_2403,N_1138,N_1242);
or U2404 (N_2404,N_1996,N_1893);
nand U2405 (N_2405,N_1405,N_1880);
nor U2406 (N_2406,N_1282,N_1442);
nor U2407 (N_2407,N_1619,N_1314);
or U2408 (N_2408,N_1114,N_1374);
or U2409 (N_2409,N_1632,N_1964);
and U2410 (N_2410,N_1390,N_1183);
xor U2411 (N_2411,N_1252,N_1654);
or U2412 (N_2412,N_1977,N_1547);
xor U2413 (N_2413,N_1508,N_1754);
xnor U2414 (N_2414,N_1312,N_1843);
xnor U2415 (N_2415,N_1322,N_1389);
or U2416 (N_2416,N_1189,N_1081);
xnor U2417 (N_2417,N_1507,N_1640);
or U2418 (N_2418,N_1581,N_1937);
or U2419 (N_2419,N_1095,N_1709);
xnor U2420 (N_2420,N_1825,N_1611);
and U2421 (N_2421,N_1435,N_1840);
or U2422 (N_2422,N_1688,N_1344);
and U2423 (N_2423,N_1101,N_1617);
or U2424 (N_2424,N_1935,N_1036);
nor U2425 (N_2425,N_1771,N_1135);
nand U2426 (N_2426,N_1052,N_1815);
nor U2427 (N_2427,N_1371,N_1739);
and U2428 (N_2428,N_1467,N_1918);
or U2429 (N_2429,N_1336,N_1591);
or U2430 (N_2430,N_1868,N_1525);
xnor U2431 (N_2431,N_1289,N_1149);
nor U2432 (N_2432,N_1748,N_1527);
nor U2433 (N_2433,N_1920,N_1176);
xnor U2434 (N_2434,N_1045,N_1382);
or U2435 (N_2435,N_1424,N_1038);
or U2436 (N_2436,N_1699,N_1298);
and U2437 (N_2437,N_1258,N_1702);
nand U2438 (N_2438,N_1100,N_1055);
and U2439 (N_2439,N_1872,N_1740);
nor U2440 (N_2440,N_1774,N_1046);
and U2441 (N_2441,N_1612,N_1686);
nand U2442 (N_2442,N_1685,N_1538);
and U2443 (N_2443,N_1085,N_1234);
xnor U2444 (N_2444,N_1929,N_1327);
xnor U2445 (N_2445,N_1275,N_1598);
xor U2446 (N_2446,N_1302,N_1767);
and U2447 (N_2447,N_1663,N_1582);
and U2448 (N_2448,N_1226,N_1277);
nand U2449 (N_2449,N_1826,N_1321);
xor U2450 (N_2450,N_1399,N_1745);
nand U2451 (N_2451,N_1272,N_1337);
or U2452 (N_2452,N_1113,N_1057);
xor U2453 (N_2453,N_1637,N_1902);
xnor U2454 (N_2454,N_1870,N_1308);
nor U2455 (N_2455,N_1457,N_1779);
xor U2456 (N_2456,N_1018,N_1240);
nand U2457 (N_2457,N_1701,N_1334);
or U2458 (N_2458,N_1734,N_1167);
xnor U2459 (N_2459,N_1784,N_1459);
or U2460 (N_2460,N_1576,N_1912);
nor U2461 (N_2461,N_1650,N_1835);
xor U2462 (N_2462,N_1728,N_1333);
nor U2463 (N_2463,N_1681,N_1309);
xor U2464 (N_2464,N_1288,N_1098);
or U2465 (N_2465,N_1111,N_1894);
and U2466 (N_2466,N_1087,N_1083);
and U2467 (N_2467,N_1584,N_1543);
nor U2468 (N_2468,N_1830,N_1813);
nand U2469 (N_2469,N_1775,N_1383);
and U2470 (N_2470,N_1731,N_1661);
or U2471 (N_2471,N_1515,N_1482);
or U2472 (N_2472,N_1764,N_1828);
nor U2473 (N_2473,N_1193,N_1437);
nand U2474 (N_2474,N_1414,N_1044);
and U2475 (N_2475,N_1510,N_1017);
and U2476 (N_2476,N_1199,N_1554);
nand U2477 (N_2477,N_1485,N_1720);
nor U2478 (N_2478,N_1512,N_1896);
or U2479 (N_2479,N_1037,N_1936);
xor U2480 (N_2480,N_1033,N_1957);
and U2481 (N_2481,N_1029,N_1415);
xnor U2482 (N_2482,N_1125,N_1075);
xor U2483 (N_2483,N_1171,N_1225);
xor U2484 (N_2484,N_1710,N_1604);
and U2485 (N_2485,N_1077,N_1354);
nand U2486 (N_2486,N_1500,N_1911);
or U2487 (N_2487,N_1431,N_1860);
xor U2488 (N_2488,N_1094,N_1089);
xnor U2489 (N_2489,N_1778,N_1799);
xnor U2490 (N_2490,N_1639,N_1364);
or U2491 (N_2491,N_1805,N_1318);
and U2492 (N_2492,N_1121,N_1638);
and U2493 (N_2493,N_1039,N_1806);
or U2494 (N_2494,N_1871,N_1682);
nor U2495 (N_2495,N_1266,N_1433);
and U2496 (N_2496,N_1890,N_1357);
and U2497 (N_2497,N_1608,N_1204);
nor U2498 (N_2498,N_1727,N_1447);
and U2499 (N_2499,N_1555,N_1990);
nand U2500 (N_2500,N_1104,N_1282);
and U2501 (N_2501,N_1302,N_1173);
and U2502 (N_2502,N_1270,N_1809);
nor U2503 (N_2503,N_1158,N_1943);
nor U2504 (N_2504,N_1532,N_1622);
nand U2505 (N_2505,N_1164,N_1348);
xor U2506 (N_2506,N_1169,N_1820);
nor U2507 (N_2507,N_1405,N_1162);
xor U2508 (N_2508,N_1069,N_1869);
and U2509 (N_2509,N_1663,N_1738);
nand U2510 (N_2510,N_1675,N_1866);
xor U2511 (N_2511,N_1853,N_1935);
nand U2512 (N_2512,N_1404,N_1871);
xor U2513 (N_2513,N_1388,N_1049);
and U2514 (N_2514,N_1024,N_1887);
nand U2515 (N_2515,N_1048,N_1652);
xor U2516 (N_2516,N_1625,N_1319);
or U2517 (N_2517,N_1685,N_1630);
and U2518 (N_2518,N_1501,N_1692);
nand U2519 (N_2519,N_1809,N_1395);
nand U2520 (N_2520,N_1940,N_1793);
nand U2521 (N_2521,N_1267,N_1724);
nand U2522 (N_2522,N_1482,N_1404);
xor U2523 (N_2523,N_1166,N_1423);
nor U2524 (N_2524,N_1210,N_1424);
or U2525 (N_2525,N_1109,N_1113);
nand U2526 (N_2526,N_1382,N_1384);
or U2527 (N_2527,N_1438,N_1651);
nand U2528 (N_2528,N_1841,N_1847);
nand U2529 (N_2529,N_1664,N_1039);
or U2530 (N_2530,N_1644,N_1888);
or U2531 (N_2531,N_1968,N_1031);
xor U2532 (N_2532,N_1540,N_1745);
nor U2533 (N_2533,N_1969,N_1790);
and U2534 (N_2534,N_1153,N_1093);
xnor U2535 (N_2535,N_1222,N_1822);
nor U2536 (N_2536,N_1208,N_1809);
nand U2537 (N_2537,N_1915,N_1681);
and U2538 (N_2538,N_1899,N_1562);
nor U2539 (N_2539,N_1245,N_1262);
nand U2540 (N_2540,N_1964,N_1970);
nand U2541 (N_2541,N_1594,N_1449);
or U2542 (N_2542,N_1671,N_1287);
or U2543 (N_2543,N_1602,N_1519);
xnor U2544 (N_2544,N_1566,N_1990);
xor U2545 (N_2545,N_1961,N_1344);
or U2546 (N_2546,N_1965,N_1658);
nor U2547 (N_2547,N_1821,N_1893);
xnor U2548 (N_2548,N_1112,N_1386);
nand U2549 (N_2549,N_1836,N_1238);
nor U2550 (N_2550,N_1651,N_1811);
nand U2551 (N_2551,N_1976,N_1374);
nor U2552 (N_2552,N_1104,N_1632);
nand U2553 (N_2553,N_1134,N_1672);
nor U2554 (N_2554,N_1368,N_1388);
nand U2555 (N_2555,N_1504,N_1479);
nor U2556 (N_2556,N_1772,N_1251);
or U2557 (N_2557,N_1774,N_1601);
nand U2558 (N_2558,N_1518,N_1399);
nand U2559 (N_2559,N_1383,N_1759);
and U2560 (N_2560,N_1367,N_1716);
and U2561 (N_2561,N_1090,N_1828);
xnor U2562 (N_2562,N_1115,N_1791);
nor U2563 (N_2563,N_1851,N_1089);
and U2564 (N_2564,N_1974,N_1804);
nor U2565 (N_2565,N_1593,N_1905);
or U2566 (N_2566,N_1289,N_1793);
nor U2567 (N_2567,N_1794,N_1281);
nor U2568 (N_2568,N_1679,N_1992);
or U2569 (N_2569,N_1162,N_1995);
and U2570 (N_2570,N_1346,N_1757);
and U2571 (N_2571,N_1563,N_1451);
nor U2572 (N_2572,N_1944,N_1624);
nand U2573 (N_2573,N_1444,N_1787);
nor U2574 (N_2574,N_1812,N_1718);
nand U2575 (N_2575,N_1786,N_1099);
and U2576 (N_2576,N_1159,N_1801);
nor U2577 (N_2577,N_1891,N_1723);
xnor U2578 (N_2578,N_1495,N_1030);
nor U2579 (N_2579,N_1543,N_1106);
xor U2580 (N_2580,N_1973,N_1654);
or U2581 (N_2581,N_1996,N_1513);
nand U2582 (N_2582,N_1920,N_1455);
or U2583 (N_2583,N_1704,N_1726);
and U2584 (N_2584,N_1742,N_1689);
nand U2585 (N_2585,N_1270,N_1843);
or U2586 (N_2586,N_1820,N_1291);
and U2587 (N_2587,N_1460,N_1318);
nand U2588 (N_2588,N_1213,N_1081);
or U2589 (N_2589,N_1871,N_1007);
xnor U2590 (N_2590,N_1168,N_1856);
nor U2591 (N_2591,N_1128,N_1333);
and U2592 (N_2592,N_1115,N_1232);
xor U2593 (N_2593,N_1703,N_1220);
and U2594 (N_2594,N_1660,N_1726);
nand U2595 (N_2595,N_1346,N_1061);
nor U2596 (N_2596,N_1626,N_1392);
nor U2597 (N_2597,N_1337,N_1030);
and U2598 (N_2598,N_1219,N_1750);
xnor U2599 (N_2599,N_1754,N_1279);
xor U2600 (N_2600,N_1833,N_1918);
nand U2601 (N_2601,N_1790,N_1160);
or U2602 (N_2602,N_1924,N_1897);
or U2603 (N_2603,N_1156,N_1820);
xor U2604 (N_2604,N_1487,N_1801);
and U2605 (N_2605,N_1462,N_1254);
or U2606 (N_2606,N_1154,N_1253);
and U2607 (N_2607,N_1054,N_1551);
nand U2608 (N_2608,N_1446,N_1836);
or U2609 (N_2609,N_1668,N_1431);
nor U2610 (N_2610,N_1510,N_1941);
nand U2611 (N_2611,N_1756,N_1639);
or U2612 (N_2612,N_1632,N_1500);
xnor U2613 (N_2613,N_1960,N_1043);
nor U2614 (N_2614,N_1884,N_1301);
nand U2615 (N_2615,N_1294,N_1214);
or U2616 (N_2616,N_1321,N_1565);
nand U2617 (N_2617,N_1113,N_1899);
nor U2618 (N_2618,N_1009,N_1310);
and U2619 (N_2619,N_1818,N_1284);
or U2620 (N_2620,N_1256,N_1737);
nand U2621 (N_2621,N_1449,N_1238);
and U2622 (N_2622,N_1651,N_1702);
xnor U2623 (N_2623,N_1836,N_1447);
nor U2624 (N_2624,N_1470,N_1034);
nor U2625 (N_2625,N_1350,N_1916);
or U2626 (N_2626,N_1714,N_1142);
and U2627 (N_2627,N_1900,N_1208);
xor U2628 (N_2628,N_1862,N_1569);
or U2629 (N_2629,N_1497,N_1124);
nor U2630 (N_2630,N_1464,N_1482);
xnor U2631 (N_2631,N_1218,N_1936);
xor U2632 (N_2632,N_1173,N_1367);
nor U2633 (N_2633,N_1585,N_1264);
nor U2634 (N_2634,N_1329,N_1269);
xor U2635 (N_2635,N_1933,N_1270);
nor U2636 (N_2636,N_1259,N_1774);
xor U2637 (N_2637,N_1648,N_1546);
nand U2638 (N_2638,N_1427,N_1508);
nand U2639 (N_2639,N_1598,N_1352);
xor U2640 (N_2640,N_1766,N_1880);
and U2641 (N_2641,N_1498,N_1573);
nor U2642 (N_2642,N_1651,N_1099);
xor U2643 (N_2643,N_1400,N_1520);
xnor U2644 (N_2644,N_1958,N_1732);
nand U2645 (N_2645,N_1801,N_1244);
nor U2646 (N_2646,N_1513,N_1534);
or U2647 (N_2647,N_1172,N_1910);
or U2648 (N_2648,N_1262,N_1445);
xnor U2649 (N_2649,N_1285,N_1649);
or U2650 (N_2650,N_1913,N_1051);
xnor U2651 (N_2651,N_1936,N_1153);
nor U2652 (N_2652,N_1088,N_1686);
nand U2653 (N_2653,N_1255,N_1857);
xor U2654 (N_2654,N_1519,N_1119);
xnor U2655 (N_2655,N_1872,N_1616);
nor U2656 (N_2656,N_1154,N_1061);
or U2657 (N_2657,N_1923,N_1475);
nor U2658 (N_2658,N_1969,N_1365);
or U2659 (N_2659,N_1229,N_1070);
and U2660 (N_2660,N_1254,N_1647);
xnor U2661 (N_2661,N_1441,N_1216);
and U2662 (N_2662,N_1312,N_1721);
or U2663 (N_2663,N_1922,N_1986);
or U2664 (N_2664,N_1362,N_1698);
or U2665 (N_2665,N_1754,N_1267);
nor U2666 (N_2666,N_1794,N_1706);
or U2667 (N_2667,N_1742,N_1626);
and U2668 (N_2668,N_1606,N_1403);
nor U2669 (N_2669,N_1547,N_1161);
nand U2670 (N_2670,N_1749,N_1636);
and U2671 (N_2671,N_1872,N_1881);
or U2672 (N_2672,N_1712,N_1016);
and U2673 (N_2673,N_1976,N_1740);
and U2674 (N_2674,N_1025,N_1165);
and U2675 (N_2675,N_1076,N_1321);
or U2676 (N_2676,N_1376,N_1391);
nor U2677 (N_2677,N_1150,N_1214);
xor U2678 (N_2678,N_1596,N_1241);
nor U2679 (N_2679,N_1299,N_1193);
or U2680 (N_2680,N_1194,N_1390);
and U2681 (N_2681,N_1259,N_1477);
or U2682 (N_2682,N_1222,N_1940);
or U2683 (N_2683,N_1079,N_1681);
nand U2684 (N_2684,N_1651,N_1381);
nand U2685 (N_2685,N_1372,N_1844);
nand U2686 (N_2686,N_1882,N_1964);
nand U2687 (N_2687,N_1607,N_1481);
and U2688 (N_2688,N_1257,N_1798);
nor U2689 (N_2689,N_1358,N_1731);
and U2690 (N_2690,N_1405,N_1128);
nor U2691 (N_2691,N_1030,N_1600);
and U2692 (N_2692,N_1796,N_1075);
xnor U2693 (N_2693,N_1390,N_1102);
and U2694 (N_2694,N_1034,N_1392);
xnor U2695 (N_2695,N_1278,N_1317);
nand U2696 (N_2696,N_1994,N_1977);
nand U2697 (N_2697,N_1683,N_1398);
or U2698 (N_2698,N_1164,N_1468);
nand U2699 (N_2699,N_1972,N_1695);
or U2700 (N_2700,N_1436,N_1366);
nand U2701 (N_2701,N_1858,N_1538);
and U2702 (N_2702,N_1689,N_1181);
and U2703 (N_2703,N_1421,N_1236);
or U2704 (N_2704,N_1691,N_1940);
nand U2705 (N_2705,N_1635,N_1206);
nor U2706 (N_2706,N_1657,N_1889);
xnor U2707 (N_2707,N_1625,N_1808);
xor U2708 (N_2708,N_1557,N_1553);
nand U2709 (N_2709,N_1638,N_1945);
and U2710 (N_2710,N_1416,N_1353);
or U2711 (N_2711,N_1805,N_1611);
or U2712 (N_2712,N_1615,N_1491);
nand U2713 (N_2713,N_1415,N_1242);
or U2714 (N_2714,N_1767,N_1020);
xor U2715 (N_2715,N_1555,N_1970);
nor U2716 (N_2716,N_1657,N_1513);
xor U2717 (N_2717,N_1934,N_1641);
nor U2718 (N_2718,N_1093,N_1178);
or U2719 (N_2719,N_1924,N_1173);
and U2720 (N_2720,N_1124,N_1836);
or U2721 (N_2721,N_1042,N_1883);
and U2722 (N_2722,N_1096,N_1565);
nor U2723 (N_2723,N_1537,N_1349);
nand U2724 (N_2724,N_1252,N_1308);
or U2725 (N_2725,N_1741,N_1948);
nor U2726 (N_2726,N_1401,N_1993);
nor U2727 (N_2727,N_1409,N_1018);
nand U2728 (N_2728,N_1882,N_1192);
or U2729 (N_2729,N_1578,N_1018);
nand U2730 (N_2730,N_1784,N_1448);
xnor U2731 (N_2731,N_1980,N_1097);
or U2732 (N_2732,N_1024,N_1774);
or U2733 (N_2733,N_1624,N_1807);
and U2734 (N_2734,N_1439,N_1925);
nor U2735 (N_2735,N_1068,N_1892);
nand U2736 (N_2736,N_1633,N_1940);
or U2737 (N_2737,N_1129,N_1303);
and U2738 (N_2738,N_1277,N_1456);
and U2739 (N_2739,N_1216,N_1892);
nor U2740 (N_2740,N_1393,N_1333);
nor U2741 (N_2741,N_1098,N_1298);
and U2742 (N_2742,N_1665,N_1533);
xnor U2743 (N_2743,N_1402,N_1742);
nor U2744 (N_2744,N_1301,N_1751);
or U2745 (N_2745,N_1573,N_1448);
and U2746 (N_2746,N_1869,N_1397);
or U2747 (N_2747,N_1194,N_1002);
xor U2748 (N_2748,N_1182,N_1882);
and U2749 (N_2749,N_1467,N_1000);
nor U2750 (N_2750,N_1763,N_1234);
xor U2751 (N_2751,N_1241,N_1862);
nand U2752 (N_2752,N_1005,N_1371);
nor U2753 (N_2753,N_1276,N_1456);
nand U2754 (N_2754,N_1620,N_1800);
nor U2755 (N_2755,N_1090,N_1363);
and U2756 (N_2756,N_1349,N_1787);
and U2757 (N_2757,N_1764,N_1153);
nand U2758 (N_2758,N_1040,N_1710);
nand U2759 (N_2759,N_1765,N_1594);
or U2760 (N_2760,N_1717,N_1761);
or U2761 (N_2761,N_1616,N_1849);
nand U2762 (N_2762,N_1772,N_1958);
or U2763 (N_2763,N_1375,N_1327);
and U2764 (N_2764,N_1050,N_1018);
or U2765 (N_2765,N_1222,N_1339);
nor U2766 (N_2766,N_1155,N_1202);
and U2767 (N_2767,N_1294,N_1205);
and U2768 (N_2768,N_1262,N_1177);
nor U2769 (N_2769,N_1852,N_1391);
nor U2770 (N_2770,N_1792,N_1311);
or U2771 (N_2771,N_1078,N_1027);
xor U2772 (N_2772,N_1122,N_1338);
or U2773 (N_2773,N_1663,N_1063);
or U2774 (N_2774,N_1928,N_1329);
xor U2775 (N_2775,N_1251,N_1048);
or U2776 (N_2776,N_1862,N_1001);
and U2777 (N_2777,N_1611,N_1039);
xnor U2778 (N_2778,N_1768,N_1373);
nor U2779 (N_2779,N_1200,N_1928);
xnor U2780 (N_2780,N_1379,N_1467);
and U2781 (N_2781,N_1735,N_1879);
nor U2782 (N_2782,N_1220,N_1163);
and U2783 (N_2783,N_1267,N_1897);
nor U2784 (N_2784,N_1263,N_1753);
xor U2785 (N_2785,N_1089,N_1222);
nor U2786 (N_2786,N_1457,N_1946);
and U2787 (N_2787,N_1088,N_1435);
nand U2788 (N_2788,N_1591,N_1768);
nand U2789 (N_2789,N_1074,N_1396);
or U2790 (N_2790,N_1789,N_1471);
nand U2791 (N_2791,N_1490,N_1049);
xor U2792 (N_2792,N_1368,N_1135);
xor U2793 (N_2793,N_1575,N_1822);
and U2794 (N_2794,N_1171,N_1735);
and U2795 (N_2795,N_1203,N_1525);
and U2796 (N_2796,N_1522,N_1590);
and U2797 (N_2797,N_1932,N_1255);
or U2798 (N_2798,N_1613,N_1794);
or U2799 (N_2799,N_1445,N_1133);
and U2800 (N_2800,N_1360,N_1924);
xor U2801 (N_2801,N_1361,N_1556);
or U2802 (N_2802,N_1174,N_1710);
or U2803 (N_2803,N_1435,N_1297);
xnor U2804 (N_2804,N_1693,N_1119);
nor U2805 (N_2805,N_1904,N_1348);
or U2806 (N_2806,N_1490,N_1131);
and U2807 (N_2807,N_1095,N_1240);
nand U2808 (N_2808,N_1354,N_1696);
and U2809 (N_2809,N_1688,N_1669);
and U2810 (N_2810,N_1676,N_1217);
or U2811 (N_2811,N_1388,N_1395);
nand U2812 (N_2812,N_1697,N_1554);
or U2813 (N_2813,N_1174,N_1403);
or U2814 (N_2814,N_1067,N_1621);
nor U2815 (N_2815,N_1601,N_1800);
and U2816 (N_2816,N_1789,N_1065);
nand U2817 (N_2817,N_1655,N_1892);
nor U2818 (N_2818,N_1882,N_1525);
and U2819 (N_2819,N_1844,N_1371);
xor U2820 (N_2820,N_1929,N_1164);
xor U2821 (N_2821,N_1784,N_1382);
nand U2822 (N_2822,N_1984,N_1359);
nand U2823 (N_2823,N_1952,N_1713);
and U2824 (N_2824,N_1695,N_1909);
and U2825 (N_2825,N_1384,N_1636);
nor U2826 (N_2826,N_1454,N_1873);
nor U2827 (N_2827,N_1001,N_1265);
nand U2828 (N_2828,N_1896,N_1063);
and U2829 (N_2829,N_1367,N_1605);
xnor U2830 (N_2830,N_1676,N_1448);
nor U2831 (N_2831,N_1776,N_1676);
nor U2832 (N_2832,N_1191,N_1256);
nand U2833 (N_2833,N_1874,N_1454);
nand U2834 (N_2834,N_1146,N_1027);
xor U2835 (N_2835,N_1452,N_1207);
nor U2836 (N_2836,N_1685,N_1437);
nor U2837 (N_2837,N_1690,N_1140);
nor U2838 (N_2838,N_1069,N_1389);
and U2839 (N_2839,N_1524,N_1587);
and U2840 (N_2840,N_1526,N_1868);
and U2841 (N_2841,N_1849,N_1667);
nand U2842 (N_2842,N_1291,N_1382);
or U2843 (N_2843,N_1452,N_1277);
nor U2844 (N_2844,N_1539,N_1297);
or U2845 (N_2845,N_1837,N_1656);
or U2846 (N_2846,N_1394,N_1437);
and U2847 (N_2847,N_1669,N_1908);
or U2848 (N_2848,N_1309,N_1777);
nand U2849 (N_2849,N_1665,N_1996);
and U2850 (N_2850,N_1611,N_1880);
nand U2851 (N_2851,N_1108,N_1490);
nand U2852 (N_2852,N_1283,N_1600);
nand U2853 (N_2853,N_1387,N_1881);
or U2854 (N_2854,N_1917,N_1719);
and U2855 (N_2855,N_1627,N_1348);
nor U2856 (N_2856,N_1427,N_1481);
or U2857 (N_2857,N_1249,N_1125);
and U2858 (N_2858,N_1595,N_1873);
or U2859 (N_2859,N_1541,N_1827);
and U2860 (N_2860,N_1378,N_1232);
and U2861 (N_2861,N_1358,N_1118);
xnor U2862 (N_2862,N_1586,N_1200);
and U2863 (N_2863,N_1133,N_1502);
nor U2864 (N_2864,N_1793,N_1333);
or U2865 (N_2865,N_1613,N_1386);
nor U2866 (N_2866,N_1138,N_1274);
or U2867 (N_2867,N_1880,N_1668);
nor U2868 (N_2868,N_1223,N_1501);
nor U2869 (N_2869,N_1447,N_1748);
or U2870 (N_2870,N_1993,N_1082);
nand U2871 (N_2871,N_1467,N_1857);
and U2872 (N_2872,N_1945,N_1758);
or U2873 (N_2873,N_1821,N_1872);
xor U2874 (N_2874,N_1359,N_1914);
xnor U2875 (N_2875,N_1166,N_1121);
and U2876 (N_2876,N_1683,N_1650);
and U2877 (N_2877,N_1837,N_1755);
nand U2878 (N_2878,N_1837,N_1991);
nor U2879 (N_2879,N_1447,N_1432);
nand U2880 (N_2880,N_1823,N_1864);
and U2881 (N_2881,N_1378,N_1787);
xnor U2882 (N_2882,N_1220,N_1863);
nor U2883 (N_2883,N_1422,N_1246);
and U2884 (N_2884,N_1936,N_1877);
xnor U2885 (N_2885,N_1336,N_1182);
nor U2886 (N_2886,N_1009,N_1184);
or U2887 (N_2887,N_1130,N_1667);
xor U2888 (N_2888,N_1359,N_1136);
or U2889 (N_2889,N_1466,N_1959);
nor U2890 (N_2890,N_1180,N_1108);
or U2891 (N_2891,N_1683,N_1861);
or U2892 (N_2892,N_1550,N_1927);
xor U2893 (N_2893,N_1269,N_1090);
nand U2894 (N_2894,N_1612,N_1085);
or U2895 (N_2895,N_1673,N_1957);
xnor U2896 (N_2896,N_1332,N_1612);
xnor U2897 (N_2897,N_1432,N_1824);
nand U2898 (N_2898,N_1784,N_1855);
nand U2899 (N_2899,N_1656,N_1818);
and U2900 (N_2900,N_1469,N_1885);
nand U2901 (N_2901,N_1374,N_1789);
xor U2902 (N_2902,N_1712,N_1596);
or U2903 (N_2903,N_1380,N_1492);
nand U2904 (N_2904,N_1133,N_1719);
or U2905 (N_2905,N_1369,N_1011);
nand U2906 (N_2906,N_1502,N_1137);
and U2907 (N_2907,N_1440,N_1218);
or U2908 (N_2908,N_1851,N_1516);
xor U2909 (N_2909,N_1348,N_1811);
xor U2910 (N_2910,N_1887,N_1175);
xnor U2911 (N_2911,N_1810,N_1518);
nor U2912 (N_2912,N_1123,N_1031);
nor U2913 (N_2913,N_1721,N_1667);
or U2914 (N_2914,N_1953,N_1842);
xnor U2915 (N_2915,N_1290,N_1295);
or U2916 (N_2916,N_1185,N_1747);
or U2917 (N_2917,N_1672,N_1584);
xnor U2918 (N_2918,N_1979,N_1806);
nor U2919 (N_2919,N_1825,N_1896);
and U2920 (N_2920,N_1491,N_1883);
and U2921 (N_2921,N_1438,N_1214);
and U2922 (N_2922,N_1038,N_1567);
nand U2923 (N_2923,N_1190,N_1058);
and U2924 (N_2924,N_1245,N_1951);
nand U2925 (N_2925,N_1919,N_1039);
nand U2926 (N_2926,N_1092,N_1920);
nand U2927 (N_2927,N_1870,N_1548);
or U2928 (N_2928,N_1057,N_1283);
nand U2929 (N_2929,N_1226,N_1186);
nor U2930 (N_2930,N_1541,N_1725);
or U2931 (N_2931,N_1057,N_1108);
or U2932 (N_2932,N_1290,N_1545);
xnor U2933 (N_2933,N_1827,N_1444);
nand U2934 (N_2934,N_1886,N_1219);
or U2935 (N_2935,N_1770,N_1247);
nor U2936 (N_2936,N_1144,N_1277);
or U2937 (N_2937,N_1273,N_1361);
nor U2938 (N_2938,N_1641,N_1937);
xnor U2939 (N_2939,N_1676,N_1684);
nor U2940 (N_2940,N_1294,N_1536);
and U2941 (N_2941,N_1507,N_1193);
xor U2942 (N_2942,N_1142,N_1876);
nor U2943 (N_2943,N_1002,N_1872);
nor U2944 (N_2944,N_1017,N_1337);
nand U2945 (N_2945,N_1639,N_1795);
nor U2946 (N_2946,N_1714,N_1260);
or U2947 (N_2947,N_1718,N_1954);
nor U2948 (N_2948,N_1553,N_1501);
xor U2949 (N_2949,N_1941,N_1101);
nand U2950 (N_2950,N_1705,N_1536);
or U2951 (N_2951,N_1329,N_1034);
and U2952 (N_2952,N_1567,N_1957);
and U2953 (N_2953,N_1697,N_1430);
or U2954 (N_2954,N_1694,N_1331);
nand U2955 (N_2955,N_1246,N_1079);
nand U2956 (N_2956,N_1599,N_1107);
xnor U2957 (N_2957,N_1943,N_1583);
or U2958 (N_2958,N_1766,N_1170);
and U2959 (N_2959,N_1755,N_1724);
xnor U2960 (N_2960,N_1391,N_1416);
nor U2961 (N_2961,N_1398,N_1377);
nor U2962 (N_2962,N_1361,N_1522);
xor U2963 (N_2963,N_1317,N_1206);
nand U2964 (N_2964,N_1072,N_1576);
nand U2965 (N_2965,N_1601,N_1885);
nand U2966 (N_2966,N_1582,N_1065);
xnor U2967 (N_2967,N_1266,N_1412);
nand U2968 (N_2968,N_1741,N_1275);
or U2969 (N_2969,N_1031,N_1962);
xnor U2970 (N_2970,N_1200,N_1423);
nor U2971 (N_2971,N_1468,N_1351);
nand U2972 (N_2972,N_1495,N_1606);
nor U2973 (N_2973,N_1065,N_1522);
nand U2974 (N_2974,N_1575,N_1931);
xor U2975 (N_2975,N_1002,N_1670);
nor U2976 (N_2976,N_1766,N_1481);
or U2977 (N_2977,N_1160,N_1404);
nor U2978 (N_2978,N_1760,N_1985);
and U2979 (N_2979,N_1612,N_1705);
xor U2980 (N_2980,N_1495,N_1044);
and U2981 (N_2981,N_1683,N_1599);
and U2982 (N_2982,N_1804,N_1877);
nand U2983 (N_2983,N_1756,N_1307);
nor U2984 (N_2984,N_1096,N_1823);
xor U2985 (N_2985,N_1105,N_1490);
or U2986 (N_2986,N_1437,N_1311);
or U2987 (N_2987,N_1092,N_1141);
nand U2988 (N_2988,N_1538,N_1306);
or U2989 (N_2989,N_1587,N_1679);
or U2990 (N_2990,N_1563,N_1683);
xor U2991 (N_2991,N_1943,N_1311);
xnor U2992 (N_2992,N_1352,N_1913);
nand U2993 (N_2993,N_1795,N_1457);
nand U2994 (N_2994,N_1229,N_1120);
and U2995 (N_2995,N_1149,N_1673);
and U2996 (N_2996,N_1896,N_1734);
nand U2997 (N_2997,N_1791,N_1677);
and U2998 (N_2998,N_1072,N_1124);
xor U2999 (N_2999,N_1680,N_1157);
xnor UO_0 (O_0,N_2841,N_2506);
nor UO_1 (O_1,N_2082,N_2544);
and UO_2 (O_2,N_2677,N_2864);
and UO_3 (O_3,N_2803,N_2287);
nand UO_4 (O_4,N_2407,N_2592);
nand UO_5 (O_5,N_2169,N_2831);
or UO_6 (O_6,N_2545,N_2116);
nor UO_7 (O_7,N_2092,N_2572);
nor UO_8 (O_8,N_2563,N_2852);
nor UO_9 (O_9,N_2203,N_2997);
nor UO_10 (O_10,N_2651,N_2960);
xor UO_11 (O_11,N_2080,N_2775);
xnor UO_12 (O_12,N_2576,N_2182);
nand UO_13 (O_13,N_2488,N_2389);
xnor UO_14 (O_14,N_2976,N_2018);
nand UO_15 (O_15,N_2917,N_2707);
or UO_16 (O_16,N_2396,N_2041);
nand UO_17 (O_17,N_2773,N_2345);
xnor UO_18 (O_18,N_2424,N_2905);
or UO_19 (O_19,N_2955,N_2685);
nand UO_20 (O_20,N_2713,N_2186);
and UO_21 (O_21,N_2224,N_2916);
nand UO_22 (O_22,N_2950,N_2821);
or UO_23 (O_23,N_2722,N_2484);
or UO_24 (O_24,N_2428,N_2109);
or UO_25 (O_25,N_2516,N_2822);
and UO_26 (O_26,N_2137,N_2240);
and UO_27 (O_27,N_2285,N_2688);
and UO_28 (O_28,N_2218,N_2341);
nand UO_29 (O_29,N_2062,N_2176);
nor UO_30 (O_30,N_2717,N_2533);
nand UO_31 (O_31,N_2930,N_2634);
xnor UO_32 (O_32,N_2799,N_2689);
xnor UO_33 (O_33,N_2724,N_2269);
nand UO_34 (O_34,N_2877,N_2543);
nor UO_35 (O_35,N_2476,N_2764);
xnor UO_36 (O_36,N_2995,N_2649);
xnor UO_37 (O_37,N_2358,N_2001);
and UO_38 (O_38,N_2144,N_2902);
nand UO_39 (O_39,N_2479,N_2475);
or UO_40 (O_40,N_2440,N_2032);
xnor UO_41 (O_41,N_2455,N_2589);
nor UO_42 (O_42,N_2007,N_2469);
xnor UO_43 (O_43,N_2142,N_2560);
nor UO_44 (O_44,N_2352,N_2417);
xnor UO_45 (O_45,N_2798,N_2855);
and UO_46 (O_46,N_2541,N_2264);
or UO_47 (O_47,N_2151,N_2656);
or UO_48 (O_48,N_2662,N_2122);
nor UO_49 (O_49,N_2650,N_2067);
and UO_50 (O_50,N_2261,N_2205);
xor UO_51 (O_51,N_2553,N_2118);
nand UO_52 (O_52,N_2781,N_2395);
nor UO_53 (O_53,N_2865,N_2800);
nand UO_54 (O_54,N_2549,N_2719);
nor UO_55 (O_55,N_2840,N_2616);
or UO_56 (O_56,N_2197,N_2654);
or UO_57 (O_57,N_2536,N_2655);
or UO_58 (O_58,N_2777,N_2190);
and UO_59 (O_59,N_2675,N_2747);
xnor UO_60 (O_60,N_2814,N_2384);
or UO_61 (O_61,N_2382,N_2404);
and UO_62 (O_62,N_2665,N_2077);
nor UO_63 (O_63,N_2568,N_2737);
and UO_64 (O_64,N_2486,N_2385);
and UO_65 (O_65,N_2646,N_2839);
or UO_66 (O_66,N_2879,N_2272);
and UO_67 (O_67,N_2982,N_2350);
and UO_68 (O_68,N_2127,N_2988);
xnor UO_69 (O_69,N_2823,N_2910);
xor UO_70 (O_70,N_2355,N_2757);
and UO_71 (O_71,N_2079,N_2083);
xor UO_72 (O_72,N_2220,N_2241);
nand UO_73 (O_73,N_2490,N_2827);
or UO_74 (O_74,N_2219,N_2157);
nand UO_75 (O_75,N_2256,N_2253);
nor UO_76 (O_76,N_2554,N_2327);
xnor UO_77 (O_77,N_2056,N_2935);
or UO_78 (O_78,N_2808,N_2332);
nand UO_79 (O_79,N_2045,N_2557);
nor UO_80 (O_80,N_2146,N_2502);
nand UO_81 (O_81,N_2415,N_2254);
and UO_82 (O_82,N_2198,N_2051);
and UO_83 (O_83,N_2913,N_2565);
xor UO_84 (O_84,N_2704,N_2785);
and UO_85 (O_85,N_2282,N_2990);
nand UO_86 (O_86,N_2586,N_2487);
nand UO_87 (O_87,N_2892,N_2088);
nand UO_88 (O_88,N_2199,N_2668);
and UO_89 (O_89,N_2830,N_2555);
nor UO_90 (O_90,N_2222,N_2787);
and UO_91 (O_91,N_2323,N_2267);
nor UO_92 (O_92,N_2661,N_2732);
nor UO_93 (O_93,N_2965,N_2094);
xnor UO_94 (O_94,N_2063,N_2848);
or UO_95 (O_95,N_2375,N_2537);
xor UO_96 (O_96,N_2333,N_2005);
nor UO_97 (O_97,N_2577,N_2867);
xor UO_98 (O_98,N_2213,N_2108);
xnor UO_99 (O_99,N_2882,N_2615);
xnor UO_100 (O_100,N_2356,N_2028);
nand UO_101 (O_101,N_2816,N_2055);
nand UO_102 (O_102,N_2097,N_2414);
xor UO_103 (O_103,N_2683,N_2521);
nand UO_104 (O_104,N_2299,N_2701);
and UO_105 (O_105,N_2979,N_2165);
nor UO_106 (O_106,N_2226,N_2311);
xor UO_107 (O_107,N_2635,N_2904);
xor UO_108 (O_108,N_2614,N_2809);
nand UO_109 (O_109,N_2061,N_2164);
nor UO_110 (O_110,N_2697,N_2187);
or UO_111 (O_111,N_2262,N_2334);
or UO_112 (O_112,N_2595,N_2054);
nand UO_113 (O_113,N_2302,N_2755);
and UO_114 (O_114,N_2002,N_2664);
xnor UO_115 (O_115,N_2695,N_2340);
and UO_116 (O_116,N_2354,N_2412);
nand UO_117 (O_117,N_2035,N_2344);
and UO_118 (O_118,N_2143,N_2221);
nand UO_119 (O_119,N_2338,N_2449);
nor UO_120 (O_120,N_2590,N_2064);
nand UO_121 (O_121,N_2049,N_2379);
xor UO_122 (O_122,N_2166,N_2914);
nor UO_123 (O_123,N_2192,N_2248);
or UO_124 (O_124,N_2700,N_2547);
nor UO_125 (O_125,N_2147,N_2971);
nand UO_126 (O_126,N_2270,N_2131);
nand UO_127 (O_127,N_2495,N_2657);
xnor UO_128 (O_128,N_2891,N_2394);
nand UO_129 (O_129,N_2617,N_2251);
xor UO_130 (O_130,N_2086,N_2893);
and UO_131 (O_131,N_2884,N_2929);
nand UO_132 (O_132,N_2312,N_2813);
and UO_133 (O_133,N_2017,N_2731);
and UO_134 (O_134,N_2343,N_2485);
xor UO_135 (O_135,N_2692,N_2819);
nand UO_136 (O_136,N_2956,N_2939);
xnor UO_137 (O_137,N_2733,N_2607);
and UO_138 (O_138,N_2567,N_2605);
or UO_139 (O_139,N_2741,N_2501);
or UO_140 (O_140,N_2712,N_2753);
nor UO_141 (O_141,N_2377,N_2445);
xnor UO_142 (O_142,N_2519,N_2837);
and UO_143 (O_143,N_2033,N_2423);
nand UO_144 (O_144,N_2968,N_2693);
nand UO_145 (O_145,N_2638,N_2335);
nor UO_146 (O_146,N_2535,N_2391);
nor UO_147 (O_147,N_2569,N_2801);
and UO_148 (O_148,N_2820,N_2128);
nand UO_149 (O_149,N_2783,N_2509);
nor UO_150 (O_150,N_2825,N_2497);
or UO_151 (O_151,N_2030,N_2772);
nand UO_152 (O_152,N_2648,N_2957);
xnor UO_153 (O_153,N_2575,N_2628);
nand UO_154 (O_154,N_2274,N_2585);
nand UO_155 (O_155,N_2769,N_2696);
nor UO_156 (O_156,N_2750,N_2708);
nand UO_157 (O_157,N_2744,N_2690);
nor UO_158 (O_158,N_2460,N_2471);
or UO_159 (O_159,N_2993,N_2066);
nand UO_160 (O_160,N_2301,N_2550);
and UO_161 (O_161,N_2673,N_2684);
nand UO_162 (O_162,N_2168,N_2387);
and UO_163 (O_163,N_2925,N_2161);
nand UO_164 (O_164,N_2120,N_2959);
or UO_165 (O_165,N_2975,N_2602);
nor UO_166 (O_166,N_2637,N_2255);
and UO_167 (O_167,N_2175,N_2718);
or UO_168 (O_168,N_2046,N_2687);
nor UO_169 (O_169,N_2915,N_2736);
xnor UO_170 (O_170,N_2158,N_2996);
and UO_171 (O_171,N_2752,N_2667);
nor UO_172 (O_172,N_2721,N_2257);
nand UO_173 (O_173,N_2791,N_2771);
nand UO_174 (O_174,N_2989,N_2659);
xnor UO_175 (O_175,N_2784,N_2492);
or UO_176 (O_176,N_2511,N_2564);
and UO_177 (O_177,N_2869,N_2991);
nor UO_178 (O_178,N_2829,N_2928);
and UO_179 (O_179,N_2400,N_2847);
or UO_180 (O_180,N_2778,N_2672);
and UO_181 (O_181,N_2815,N_2949);
or UO_182 (O_182,N_2843,N_2729);
xor UO_183 (O_183,N_2580,N_2038);
xnor UO_184 (O_184,N_2691,N_2402);
nand UO_185 (O_185,N_2053,N_2139);
nand UO_186 (O_186,N_2907,N_2876);
nand UO_187 (O_187,N_2624,N_2438);
and UO_188 (O_188,N_2973,N_2320);
nor UO_189 (O_189,N_2348,N_2851);
or UO_190 (O_190,N_2326,N_2838);
nor UO_191 (O_191,N_2003,N_2606);
and UO_192 (O_192,N_2994,N_2878);
nor UO_193 (O_193,N_2101,N_2406);
and UO_194 (O_194,N_2517,N_2068);
or UO_195 (O_195,N_2709,N_2277);
or UO_196 (O_196,N_2948,N_2011);
xor UO_197 (O_197,N_2467,N_2705);
nand UO_198 (O_198,N_2503,N_2663);
nor UO_199 (O_199,N_2181,N_2482);
xnor UO_200 (O_200,N_2232,N_2618);
and UO_201 (O_201,N_2933,N_2266);
or UO_202 (O_202,N_2797,N_2857);
xor UO_203 (O_203,N_2281,N_2728);
or UO_204 (O_204,N_2639,N_2875);
nor UO_205 (O_205,N_2317,N_2748);
and UO_206 (O_206,N_2818,N_2401);
nand UO_207 (O_207,N_2514,N_2100);
nor UO_208 (O_208,N_2325,N_2444);
or UO_209 (O_209,N_2858,N_2940);
xnor UO_210 (O_210,N_2026,N_2716);
xor UO_211 (O_211,N_2610,N_2529);
nand UO_212 (O_212,N_2314,N_2870);
nor UO_213 (O_213,N_2546,N_2505);
and UO_214 (O_214,N_2494,N_2461);
nor UO_215 (O_215,N_2022,N_2945);
and UO_216 (O_216,N_2745,N_2459);
and UO_217 (O_217,N_2245,N_2518);
and UO_218 (O_218,N_2899,N_2571);
nor UO_219 (O_219,N_2641,N_2084);
nand UO_220 (O_220,N_2008,N_2652);
nand UO_221 (O_221,N_2739,N_2596);
nand UO_222 (O_222,N_2633,N_2980);
or UO_223 (O_223,N_2193,N_2725);
nor UO_224 (O_224,N_2574,N_2040);
nor UO_225 (O_225,N_2630,N_2632);
or UO_226 (O_226,N_2433,N_2235);
xor UO_227 (O_227,N_2981,N_2179);
and UO_228 (O_228,N_2102,N_2360);
nand UO_229 (O_229,N_2278,N_2970);
xor UO_230 (O_230,N_2742,N_2888);
xor UO_231 (O_231,N_2896,N_2145);
or UO_232 (O_232,N_2489,N_2920);
xnor UO_233 (O_233,N_2817,N_2020);
and UO_234 (O_234,N_2075,N_2794);
or UO_235 (O_235,N_2496,N_2200);
nor UO_236 (O_236,N_2983,N_2763);
nor UO_237 (O_237,N_2622,N_2156);
or UO_238 (O_238,N_2135,N_2322);
or UO_239 (O_239,N_2059,N_2034);
nor UO_240 (O_240,N_2448,N_2362);
and UO_241 (O_241,N_2629,N_2790);
xor UO_242 (O_242,N_2951,N_2405);
nor UO_243 (O_243,N_2862,N_2367);
and UO_244 (O_244,N_2582,N_2873);
nor UO_245 (O_245,N_2263,N_2531);
xor UO_246 (O_246,N_2740,N_2016);
xor UO_247 (O_247,N_2863,N_2499);
or UO_248 (O_248,N_2242,N_2845);
nand UO_249 (O_249,N_2609,N_2726);
nor UO_250 (O_250,N_2604,N_2942);
nor UO_251 (O_251,N_2296,N_2283);
nor UO_252 (O_252,N_2608,N_2227);
xnor UO_253 (O_253,N_2528,N_2887);
or UO_254 (O_254,N_2021,N_2252);
nand UO_255 (O_255,N_2964,N_2627);
and UO_256 (O_256,N_2105,N_2336);
nor UO_257 (O_257,N_2670,N_2280);
xor UO_258 (O_258,N_2805,N_2937);
or UO_259 (O_259,N_2149,N_2029);
xnor UO_260 (O_260,N_2500,N_2019);
nor UO_261 (O_261,N_2416,N_2774);
nor UO_262 (O_262,N_2793,N_2749);
xor UO_263 (O_263,N_2099,N_2076);
xor UO_264 (O_264,N_2714,N_2447);
or UO_265 (O_265,N_2163,N_2986);
and UO_266 (O_266,N_2903,N_2954);
nor UO_267 (O_267,N_2620,N_2504);
and UO_268 (O_268,N_2436,N_2160);
or UO_269 (O_269,N_2006,N_2756);
nand UO_270 (O_270,N_2998,N_2611);
and UO_271 (O_271,N_2559,N_2191);
nand UO_272 (O_272,N_2653,N_2470);
xnor UO_273 (O_273,N_2969,N_2095);
nand UO_274 (O_274,N_2050,N_2408);
xnor UO_275 (O_275,N_2478,N_2710);
nor UO_276 (O_276,N_2472,N_2594);
xor UO_277 (O_277,N_2573,N_2908);
and UO_278 (O_278,N_2601,N_2947);
nor UO_279 (O_279,N_2702,N_2273);
xnor UO_280 (O_280,N_2674,N_2081);
or UO_281 (O_281,N_2792,N_2309);
xnor UO_282 (O_282,N_2824,N_2432);
nand UO_283 (O_283,N_2515,N_2846);
xnor UO_284 (O_284,N_2295,N_2443);
and UO_285 (O_285,N_2890,N_2390);
or UO_286 (O_286,N_2625,N_2353);
nor UO_287 (O_287,N_2259,N_2932);
xnor UO_288 (O_288,N_2883,N_2374);
and UO_289 (O_289,N_2435,N_2682);
nor UO_290 (O_290,N_2934,N_2856);
nor UO_291 (O_291,N_2631,N_2216);
nand UO_292 (O_292,N_2359,N_2860);
nand UO_293 (O_293,N_2392,N_2473);
xor UO_294 (O_294,N_2539,N_2419);
xor UO_295 (O_295,N_2786,N_2125);
nand UO_296 (O_296,N_2681,N_2881);
xor UO_297 (O_297,N_2978,N_2897);
and UO_298 (O_298,N_2119,N_2369);
nor UO_299 (O_299,N_2397,N_2480);
xor UO_300 (O_300,N_2331,N_2307);
or UO_301 (O_301,N_2922,N_2944);
and UO_302 (O_302,N_2526,N_2911);
xnor UO_303 (O_303,N_2085,N_2579);
nor UO_304 (O_304,N_2894,N_2393);
nor UO_305 (O_305,N_2581,N_2676);
xnor UO_306 (O_306,N_2446,N_2421);
and UO_307 (O_307,N_2104,N_2315);
or UO_308 (O_308,N_2812,N_2645);
or UO_309 (O_309,N_2244,N_2291);
nand UO_310 (O_310,N_2727,N_2807);
and UO_311 (O_311,N_2154,N_2715);
nand UO_312 (O_312,N_2588,N_2265);
and UO_313 (O_313,N_2351,N_2136);
or UO_314 (O_314,N_2779,N_2880);
xor UO_315 (O_315,N_2538,N_2210);
nand UO_316 (O_316,N_2861,N_2130);
xnor UO_317 (O_317,N_2201,N_2698);
xnor UO_318 (O_318,N_2530,N_2089);
or UO_319 (O_319,N_2140,N_2184);
nand UO_320 (O_320,N_2542,N_2931);
xor UO_321 (O_321,N_2962,N_2188);
and UO_322 (O_322,N_2422,N_2699);
nor UO_323 (O_323,N_2765,N_2303);
nand UO_324 (O_324,N_2039,N_2508);
xnor UO_325 (O_325,N_2174,N_2121);
nor UO_326 (O_326,N_2720,N_2318);
nor UO_327 (O_327,N_2398,N_2238);
and UO_328 (O_328,N_2074,N_2172);
nor UO_329 (O_329,N_2173,N_2308);
or UO_330 (O_330,N_2912,N_2426);
nand UO_331 (O_331,N_2464,N_2427);
or UO_332 (O_332,N_2313,N_2211);
nand UO_333 (O_333,N_2498,N_2298);
and UO_334 (O_334,N_2346,N_2598);
xor UO_335 (O_335,N_2376,N_2552);
nand UO_336 (O_336,N_2069,N_2096);
and UO_337 (O_337,N_2152,N_2548);
xor UO_338 (O_338,N_2886,N_2743);
nand UO_339 (O_339,N_2758,N_2091);
or UO_340 (O_340,N_2292,N_2523);
nor UO_341 (O_341,N_2974,N_2431);
xor UO_342 (O_342,N_2456,N_2371);
xnor UO_343 (O_343,N_2249,N_2520);
and UO_344 (O_344,N_2112,N_2413);
or UO_345 (O_345,N_2561,N_2963);
or UO_346 (O_346,N_2047,N_2826);
nand UO_347 (O_347,N_2621,N_2465);
or UO_348 (O_348,N_2409,N_2678);
xnor UO_349 (O_349,N_2058,N_2111);
xor UO_350 (O_350,N_2671,N_2802);
nand UO_351 (O_351,N_2992,N_2977);
xor UO_352 (O_352,N_2027,N_2070);
nand UO_353 (O_353,N_2759,N_2872);
and UO_354 (O_354,N_2834,N_2735);
xor UO_355 (O_355,N_2065,N_2462);
or UO_356 (O_356,N_2189,N_2150);
nand UO_357 (O_357,N_2780,N_2760);
nand UO_358 (O_358,N_2450,N_2388);
and UO_359 (O_359,N_2098,N_2031);
or UO_360 (O_360,N_2583,N_2153);
xor UO_361 (O_361,N_2789,N_2167);
nand UO_362 (O_362,N_2430,N_2177);
or UO_363 (O_363,N_2329,N_2386);
nor UO_364 (O_364,N_2636,N_2507);
xor UO_365 (O_365,N_2178,N_2669);
or UO_366 (O_366,N_2525,N_2215);
nand UO_367 (O_367,N_2999,N_2042);
nand UO_368 (O_368,N_2349,N_2703);
or UO_369 (O_369,N_2686,N_2953);
nand UO_370 (O_370,N_2279,N_2048);
nand UO_371 (O_371,N_2037,N_2694);
xnor UO_372 (O_372,N_2305,N_2293);
xnor UO_373 (O_373,N_2171,N_2613);
nor UO_374 (O_374,N_2987,N_2403);
xor UO_375 (O_375,N_2828,N_2584);
nor UO_376 (O_376,N_2593,N_2090);
and UO_377 (O_377,N_2310,N_2558);
nand UO_378 (O_378,N_2036,N_2660);
or UO_379 (O_379,N_2357,N_2556);
or UO_380 (O_380,N_2836,N_2746);
nand UO_381 (O_381,N_2228,N_2952);
nand UO_382 (O_382,N_2434,N_2938);
nor UO_383 (O_383,N_2477,N_2300);
nor UO_384 (O_384,N_2463,N_2366);
nand UO_385 (O_385,N_2373,N_2025);
and UO_386 (O_386,N_2113,N_2788);
nand UO_387 (O_387,N_2365,N_2347);
nand UO_388 (O_388,N_2383,N_2231);
and UO_389 (O_389,N_2207,N_2276);
xnor UO_390 (O_390,N_2513,N_2943);
or UO_391 (O_391,N_2866,N_2591);
xnor UO_392 (O_392,N_2212,N_2304);
nor UO_393 (O_393,N_2138,N_2141);
or UO_394 (O_394,N_2324,N_2015);
nor UO_395 (O_395,N_2439,N_2853);
nor UO_396 (O_396,N_2418,N_2597);
nand UO_397 (O_397,N_2243,N_2919);
and UO_398 (O_398,N_2871,N_2849);
or UO_399 (O_399,N_2967,N_2399);
nand UO_400 (O_400,N_2004,N_2380);
nand UO_401 (O_401,N_2206,N_2562);
xor UO_402 (O_402,N_2159,N_2132);
nor UO_403 (O_403,N_2734,N_2319);
xor UO_404 (O_404,N_2924,N_2425);
nand UO_405 (O_405,N_2457,N_2233);
xor UO_406 (O_406,N_2372,N_2208);
nand UO_407 (O_407,N_2420,N_2895);
xnor UO_408 (O_408,N_2850,N_2306);
nand UO_409 (O_409,N_2225,N_2901);
nor UO_410 (O_410,N_2600,N_2466);
nor UO_411 (O_411,N_2115,N_2009);
or UO_412 (O_412,N_2795,N_2289);
nand UO_413 (O_413,N_2124,N_2275);
nand UO_414 (O_414,N_2658,N_2442);
xor UO_415 (O_415,N_2183,N_2854);
and UO_416 (O_416,N_2885,N_2180);
or UO_417 (O_417,N_2468,N_2918);
nor UO_418 (O_418,N_2437,N_2014);
and UO_419 (O_419,N_2195,N_2024);
nand UO_420 (O_420,N_2532,N_2217);
nand UO_421 (O_421,N_2288,N_2129);
or UO_422 (O_422,N_2134,N_2804);
and UO_423 (O_423,N_2117,N_2644);
and UO_424 (O_424,N_2776,N_2483);
or UO_425 (O_425,N_2761,N_2052);
and UO_426 (O_426,N_2859,N_2512);
and UO_427 (O_427,N_2770,N_2204);
nand UO_428 (O_428,N_2972,N_2909);
nor UO_429 (O_429,N_2844,N_2522);
and UO_430 (O_430,N_2321,N_2566);
nor UO_431 (O_431,N_2474,N_2551);
xnor UO_432 (O_432,N_2454,N_2711);
nand UO_433 (O_433,N_2923,N_2209);
xnor UO_434 (O_434,N_2540,N_2679);
nor UO_435 (O_435,N_2491,N_2268);
or UO_436 (O_436,N_2411,N_2599);
nand UO_437 (O_437,N_2078,N_2762);
xnor UO_438 (O_438,N_2236,N_2453);
nand UO_439 (O_439,N_2754,N_2961);
xor UO_440 (O_440,N_2044,N_2337);
nor UO_441 (O_441,N_2010,N_2107);
and UO_442 (O_442,N_2106,N_2229);
or UO_443 (O_443,N_2133,N_2316);
nor UO_444 (O_444,N_2093,N_2832);
nand UO_445 (O_445,N_2868,N_2271);
xor UO_446 (O_446,N_2185,N_2363);
xor UO_447 (O_447,N_2230,N_2666);
xor UO_448 (O_448,N_2429,N_2835);
nor UO_449 (O_449,N_2643,N_2239);
or UO_450 (O_450,N_2330,N_2114);
or UO_451 (O_451,N_2730,N_2946);
or UO_452 (O_452,N_2234,N_2647);
xor UO_453 (O_453,N_2570,N_2510);
xor UO_454 (O_454,N_2043,N_2623);
or UO_455 (O_455,N_2072,N_2361);
or UO_456 (O_456,N_2452,N_2294);
nand UO_457 (O_457,N_2767,N_2906);
nand UO_458 (O_458,N_2926,N_2196);
nor UO_459 (O_459,N_2612,N_2833);
xnor UO_460 (O_460,N_2260,N_2214);
nor UO_461 (O_461,N_2162,N_2441);
or UO_462 (O_462,N_2481,N_2364);
xor UO_463 (O_463,N_2000,N_2984);
and UO_464 (O_464,N_2768,N_2073);
nor UO_465 (O_465,N_2921,N_2368);
nor UO_466 (O_466,N_2527,N_2071);
or UO_467 (O_467,N_2619,N_2958);
nor UO_468 (O_468,N_2342,N_2706);
and UO_469 (O_469,N_2898,N_2202);
nor UO_470 (O_470,N_2806,N_2126);
and UO_471 (O_471,N_2810,N_2782);
or UO_472 (O_472,N_2023,N_2286);
nand UO_473 (O_473,N_2258,N_2603);
nor UO_474 (O_474,N_2451,N_2493);
or UO_475 (O_475,N_2587,N_2123);
nor UO_476 (O_476,N_2889,N_2738);
nand UO_477 (O_477,N_2900,N_2766);
and UO_478 (O_478,N_2534,N_2370);
nor UO_479 (O_479,N_2328,N_2148);
and UO_480 (O_480,N_2087,N_2223);
or UO_481 (O_481,N_2642,N_2284);
or UO_482 (O_482,N_2796,N_2842);
and UO_483 (O_483,N_2723,N_2640);
nand UO_484 (O_484,N_2013,N_2811);
or UO_485 (O_485,N_2250,N_2290);
and UO_486 (O_486,N_2626,N_2936);
nor UO_487 (O_487,N_2874,N_2060);
xor UO_488 (O_488,N_2378,N_2012);
and UO_489 (O_489,N_2103,N_2524);
and UO_490 (O_490,N_2170,N_2966);
nor UO_491 (O_491,N_2155,N_2751);
xor UO_492 (O_492,N_2246,N_2339);
nor UO_493 (O_493,N_2110,N_2410);
xor UO_494 (O_494,N_2941,N_2237);
and UO_495 (O_495,N_2985,N_2247);
nor UO_496 (O_496,N_2927,N_2680);
xor UO_497 (O_497,N_2381,N_2297);
nand UO_498 (O_498,N_2194,N_2057);
xnor UO_499 (O_499,N_2458,N_2578);
endmodule