module basic_1000_10000_1500_5_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_187,In_272);
nand U1 (N_1,In_719,In_121);
nor U2 (N_2,In_401,In_33);
and U3 (N_3,In_425,In_836);
nand U4 (N_4,In_704,In_235);
nand U5 (N_5,In_708,In_580);
or U6 (N_6,In_981,In_296);
and U7 (N_7,In_735,In_157);
nor U8 (N_8,In_30,In_18);
and U9 (N_9,In_684,In_163);
and U10 (N_10,In_206,In_636);
or U11 (N_11,In_584,In_522);
and U12 (N_12,In_91,In_196);
and U13 (N_13,In_88,In_55);
or U14 (N_14,In_601,In_267);
nor U15 (N_15,In_850,In_883);
and U16 (N_16,In_35,In_644);
nor U17 (N_17,In_410,In_338);
nand U18 (N_18,In_518,In_640);
and U19 (N_19,In_377,In_268);
nand U20 (N_20,In_71,In_602);
xor U21 (N_21,In_537,In_552);
nand U22 (N_22,In_889,In_86);
nand U23 (N_23,In_42,In_100);
nor U24 (N_24,In_955,In_178);
nor U25 (N_25,In_585,In_515);
nand U26 (N_26,In_242,In_882);
or U27 (N_27,In_558,In_360);
and U28 (N_28,In_11,In_737);
or U29 (N_29,In_185,In_723);
or U30 (N_30,In_97,In_613);
or U31 (N_31,In_551,In_978);
nand U32 (N_32,In_765,In_226);
nor U33 (N_33,In_824,In_49);
or U34 (N_34,In_872,In_17);
and U35 (N_35,In_311,In_966);
and U36 (N_36,In_230,In_921);
nor U37 (N_37,In_470,In_307);
nor U38 (N_38,In_670,In_36);
or U39 (N_39,In_700,In_96);
nand U40 (N_40,In_788,In_867);
nand U41 (N_41,In_404,In_925);
nand U42 (N_42,In_133,In_176);
nand U43 (N_43,In_958,In_860);
and U44 (N_44,In_817,In_615);
and U45 (N_45,In_977,In_650);
or U46 (N_46,In_729,In_171);
nand U47 (N_47,In_648,In_856);
nor U48 (N_48,In_713,In_645);
or U49 (N_49,In_498,In_174);
nor U50 (N_50,In_46,In_864);
nand U51 (N_51,In_895,In_420);
or U52 (N_52,In_571,In_341);
nand U53 (N_53,In_626,In_510);
nand U54 (N_54,In_592,In_288);
or U55 (N_55,In_682,In_778);
and U56 (N_56,In_767,In_172);
and U57 (N_57,In_878,In_707);
or U58 (N_58,In_766,In_691);
nand U59 (N_59,In_203,In_374);
nor U60 (N_60,In_52,In_660);
nand U61 (N_61,In_790,In_982);
and U62 (N_62,In_800,In_450);
nand U63 (N_63,In_590,In_509);
and U64 (N_64,In_451,In_1);
or U65 (N_65,In_538,In_932);
nand U66 (N_66,In_136,In_173);
or U67 (N_67,In_475,In_198);
nor U68 (N_68,In_968,In_953);
nand U69 (N_69,In_458,In_68);
nand U70 (N_70,In_480,In_622);
or U71 (N_71,In_880,In_317);
nand U72 (N_72,In_284,In_854);
or U73 (N_73,In_581,In_167);
or U74 (N_74,In_78,In_671);
and U75 (N_75,In_210,In_367);
nand U76 (N_76,In_933,In_297);
nand U77 (N_77,In_840,In_327);
nand U78 (N_78,In_140,In_389);
nor U79 (N_79,In_569,In_438);
and U80 (N_80,In_144,In_370);
and U81 (N_81,In_714,In_653);
or U82 (N_82,In_663,In_734);
nor U83 (N_83,In_429,In_718);
nand U84 (N_84,In_436,In_110);
or U85 (N_85,In_48,In_869);
nor U86 (N_86,In_833,In_138);
or U87 (N_87,In_959,In_190);
nor U88 (N_88,In_989,In_384);
nor U89 (N_89,In_668,In_629);
nand U90 (N_90,In_314,In_278);
or U91 (N_91,In_524,In_616);
nand U92 (N_92,In_447,In_417);
nor U93 (N_93,In_768,In_744);
or U94 (N_94,In_479,In_63);
or U95 (N_95,In_95,In_464);
or U96 (N_96,In_208,In_852);
nand U97 (N_97,In_545,In_620);
or U98 (N_98,In_784,In_4);
and U99 (N_99,In_987,In_356);
or U100 (N_100,In_870,In_383);
nand U101 (N_101,In_935,In_435);
or U102 (N_102,In_694,In_114);
nand U103 (N_103,In_930,In_686);
nand U104 (N_104,In_712,In_459);
nand U105 (N_105,In_40,In_281);
nand U106 (N_106,In_302,In_504);
and U107 (N_107,In_603,In_80);
and U108 (N_108,In_868,In_485);
nand U109 (N_109,In_624,In_974);
nand U110 (N_110,In_466,In_74);
or U111 (N_111,In_915,In_588);
or U112 (N_112,In_927,In_559);
and U113 (N_113,In_323,In_760);
nand U114 (N_114,In_117,In_546);
or U115 (N_115,In_407,In_655);
and U116 (N_116,In_597,In_802);
or U117 (N_117,In_28,In_320);
nor U118 (N_118,In_433,In_240);
and U119 (N_119,In_773,In_491);
and U120 (N_120,In_627,In_848);
or U121 (N_121,In_593,In_460);
or U122 (N_122,In_26,In_248);
and U123 (N_123,In_938,In_416);
nor U124 (N_124,In_967,In_53);
or U125 (N_125,In_637,In_610);
nor U126 (N_126,In_813,In_570);
and U127 (N_127,In_853,In_654);
or U128 (N_128,In_876,In_999);
nor U129 (N_129,In_358,In_123);
or U130 (N_130,In_432,In_646);
or U131 (N_131,In_238,In_446);
nand U132 (N_132,In_772,In_961);
and U133 (N_133,In_501,In_24);
nand U134 (N_134,In_168,In_994);
nor U135 (N_135,In_596,In_85);
and U136 (N_136,In_422,In_595);
nor U137 (N_137,In_471,In_200);
and U138 (N_138,In_962,In_505);
nor U139 (N_139,In_411,In_62);
or U140 (N_140,In_695,In_126);
and U141 (N_141,In_231,In_984);
nand U142 (N_142,In_224,In_32);
or U143 (N_143,In_56,In_263);
and U144 (N_144,In_403,In_722);
nand U145 (N_145,In_359,In_947);
or U146 (N_146,In_991,In_201);
nand U147 (N_147,In_0,In_348);
nor U148 (N_148,In_112,In_855);
nand U149 (N_149,In_717,In_738);
or U150 (N_150,In_942,In_764);
or U151 (N_151,In_441,In_742);
or U152 (N_152,In_412,In_562);
nand U153 (N_153,In_652,In_271);
and U154 (N_154,In_154,In_69);
and U155 (N_155,In_779,In_222);
and U156 (N_156,In_631,In_806);
and U157 (N_157,In_667,In_607);
nor U158 (N_158,In_844,In_34);
and U159 (N_159,In_57,In_65);
nor U160 (N_160,In_478,In_945);
nand U161 (N_161,In_553,In_177);
nand U162 (N_162,In_762,In_642);
or U163 (N_163,In_67,In_783);
nand U164 (N_164,In_948,In_818);
nor U165 (N_165,In_757,In_493);
nor U166 (N_166,In_365,In_221);
and U167 (N_167,In_294,In_748);
nor U168 (N_168,In_688,In_687);
or U169 (N_169,In_90,In_547);
and U170 (N_170,In_555,In_794);
nand U171 (N_171,In_262,In_771);
nor U172 (N_172,In_419,In_336);
and U173 (N_173,In_679,In_319);
nor U174 (N_174,In_996,In_59);
nand U175 (N_175,In_634,In_134);
or U176 (N_176,In_488,In_874);
nand U177 (N_177,In_260,In_431);
xor U178 (N_178,In_290,In_58);
nand U179 (N_179,In_649,In_430);
nor U180 (N_180,In_361,In_674);
or U181 (N_181,In_741,In_128);
and U182 (N_182,In_342,In_328);
or U183 (N_183,In_499,In_892);
or U184 (N_184,In_37,In_143);
nand U185 (N_185,In_202,In_863);
nor U186 (N_186,In_199,In_27);
nor U187 (N_187,In_651,In_347);
and U188 (N_188,In_672,In_931);
nor U189 (N_189,In_375,In_261);
and U190 (N_190,In_727,In_259);
nor U191 (N_191,In_194,In_286);
or U192 (N_192,In_720,In_378);
nand U193 (N_193,In_600,In_258);
xor U194 (N_194,In_904,In_252);
nor U195 (N_195,In_386,In_903);
and U196 (N_196,In_693,In_770);
or U197 (N_197,In_612,In_265);
and U198 (N_198,In_151,In_685);
nor U199 (N_199,In_937,In_690);
or U200 (N_200,In_983,In_905);
and U201 (N_201,In_703,In_155);
or U202 (N_202,In_705,In_912);
nand U203 (N_203,In_979,In_84);
or U204 (N_204,In_246,In_835);
nor U205 (N_205,In_591,In_796);
nand U206 (N_206,In_897,In_975);
nand U207 (N_207,In_149,In_807);
nor U208 (N_208,In_696,In_139);
or U209 (N_209,In_124,In_211);
nand U210 (N_210,In_6,In_541);
or U211 (N_211,In_639,In_871);
nor U212 (N_212,In_357,In_396);
or U213 (N_213,In_98,In_763);
or U214 (N_214,In_500,In_725);
or U215 (N_215,In_301,In_158);
nand U216 (N_216,In_564,In_456);
or U217 (N_217,In_264,In_287);
nor U218 (N_218,In_387,In_379);
and U219 (N_219,In_815,In_598);
or U220 (N_220,In_236,In_186);
or U221 (N_221,In_957,In_408);
nand U222 (N_222,In_502,In_204);
nand U223 (N_223,In_469,In_249);
nor U224 (N_224,In_223,In_822);
nand U225 (N_225,In_195,In_656);
nand U226 (N_226,In_527,In_998);
and U227 (N_227,In_544,In_661);
nor U228 (N_228,In_944,In_842);
nand U229 (N_229,In_809,In_119);
and U230 (N_230,In_461,In_291);
nor U231 (N_231,In_680,In_891);
nand U232 (N_232,In_971,In_299);
or U233 (N_233,In_520,In_216);
and U234 (N_234,In_94,In_623);
nand U235 (N_235,In_665,In_87);
or U236 (N_236,In_218,In_215);
nand U237 (N_237,In_758,In_929);
or U238 (N_238,In_392,In_219);
or U239 (N_239,In_535,In_394);
nor U240 (N_240,In_93,In_303);
nand U241 (N_241,In_164,In_350);
nor U242 (N_242,In_829,In_355);
nor U243 (N_243,In_183,In_332);
nand U244 (N_244,In_956,In_746);
or U245 (N_245,In_799,In_519);
or U246 (N_246,In_756,In_513);
or U247 (N_247,In_599,In_706);
or U248 (N_248,In_170,In_289);
nor U249 (N_249,In_339,In_542);
nor U250 (N_250,In_711,In_279);
nand U251 (N_251,In_821,In_300);
or U252 (N_252,In_823,In_572);
or U253 (N_253,In_362,In_440);
or U254 (N_254,In_462,In_827);
nor U255 (N_255,In_819,In_709);
or U256 (N_256,In_954,In_740);
and U257 (N_257,In_873,In_621);
or U258 (N_258,In_344,In_77);
and U259 (N_259,In_251,In_269);
and U260 (N_260,In_345,In_483);
nor U261 (N_261,In_442,In_120);
and U262 (N_262,In_795,In_917);
nand U263 (N_263,In_244,In_506);
nand U264 (N_264,In_14,In_255);
and U265 (N_265,In_15,In_638);
nand U266 (N_266,In_521,In_313);
nand U267 (N_267,In_181,In_503);
and U268 (N_268,In_23,In_614);
nand U269 (N_269,In_988,In_277);
and U270 (N_270,In_184,In_111);
or U271 (N_271,In_549,In_444);
nand U272 (N_272,In_769,In_609);
nor U273 (N_273,In_79,In_141);
nor U274 (N_274,In_561,In_516);
nor U275 (N_275,In_632,In_970);
and U276 (N_276,In_793,In_51);
nor U277 (N_277,In_791,In_894);
and U278 (N_278,In_888,In_494);
or U279 (N_279,In_828,In_424);
and U280 (N_280,In_101,In_241);
nand U281 (N_281,In_220,In_192);
nor U282 (N_282,In_625,In_454);
nand U283 (N_283,In_229,In_885);
nand U284 (N_284,In_212,In_566);
nand U285 (N_285,In_617,In_382);
nor U286 (N_286,In_877,In_577);
nor U287 (N_287,In_16,In_761);
nor U288 (N_288,In_750,In_38);
or U289 (N_289,In_161,In_107);
and U290 (N_290,In_759,In_664);
and U291 (N_291,In_926,In_225);
nor U292 (N_292,In_608,In_463);
nand U293 (N_293,In_465,In_841);
nand U294 (N_294,In_305,In_39);
and U295 (N_295,In_391,In_116);
or U296 (N_296,In_12,In_274);
and U297 (N_297,In_354,In_804);
and U298 (N_298,In_658,In_531);
and U299 (N_299,In_973,In_330);
and U300 (N_300,In_364,In_125);
nand U301 (N_301,In_31,In_232);
and U302 (N_302,In_534,In_207);
nand U303 (N_303,In_413,In_749);
or U304 (N_304,In_409,In_924);
nand U305 (N_305,In_142,In_605);
xor U306 (N_306,In_7,In_312);
nand U307 (N_307,In_29,In_292);
nand U308 (N_308,In_960,In_745);
nor U309 (N_309,In_865,In_539);
or U310 (N_310,In_434,In_439);
nand U311 (N_311,In_775,In_283);
or U312 (N_312,In_697,In_659);
and U313 (N_313,In_227,In_82);
and U314 (N_314,In_568,In_474);
nor U315 (N_315,In_54,In_326);
nor U316 (N_316,In_847,In_512);
nand U317 (N_317,In_105,In_393);
or U318 (N_318,In_487,In_875);
and U319 (N_319,In_754,In_940);
and U320 (N_320,In_633,In_369);
or U321 (N_321,In_346,In_941);
or U322 (N_322,In_557,In_657);
nand U323 (N_323,In_191,In_898);
nor U324 (N_324,In_721,In_239);
or U325 (N_325,In_579,In_736);
nand U326 (N_326,In_820,In_148);
nor U327 (N_327,In_985,In_702);
and U328 (N_328,In_395,In_563);
nor U329 (N_329,In_776,In_366);
and U330 (N_330,In_641,In_963);
nand U331 (N_331,In_965,In_373);
or U332 (N_332,In_913,In_368);
nor U333 (N_333,In_152,In_145);
nor U334 (N_334,In_21,In_310);
and U335 (N_335,In_402,In_669);
and U336 (N_336,In_481,In_254);
nand U337 (N_337,In_60,In_182);
nand U338 (N_338,In_901,In_293);
nor U339 (N_339,In_445,In_489);
or U340 (N_340,In_245,In_851);
and U341 (N_341,In_604,In_160);
and U342 (N_342,In_256,In_922);
and U343 (N_343,In_179,In_677);
or U344 (N_344,In_911,In_131);
nor U345 (N_345,In_472,In_525);
and U346 (N_346,In_934,In_811);
nand U347 (N_347,In_747,In_335);
or U348 (N_348,In_381,In_106);
nor U349 (N_349,In_859,In_540);
or U350 (N_350,In_780,In_692);
or U351 (N_351,In_532,In_846);
nand U352 (N_352,In_397,In_906);
nor U353 (N_353,In_507,In_666);
nor U354 (N_354,In_83,In_986);
and U355 (N_355,In_298,In_914);
nand U356 (N_356,In_837,In_9);
nor U357 (N_357,In_550,In_122);
nand U358 (N_358,In_951,In_834);
or U359 (N_359,In_826,In_529);
nand U360 (N_360,In_533,In_919);
nor U361 (N_361,In_421,In_743);
nand U362 (N_362,In_405,In_406);
or U363 (N_363,In_275,In_990);
or U364 (N_364,In_839,In_890);
nor U365 (N_365,In_887,In_468);
or U366 (N_366,In_964,In_751);
nor U367 (N_367,In_969,In_70);
nor U368 (N_368,In_511,In_270);
nand U369 (N_369,In_118,In_643);
and U370 (N_370,In_673,In_388);
and U371 (N_371,In_589,In_103);
xor U372 (N_372,In_188,In_418);
and U373 (N_373,In_233,In_162);
nand U374 (N_374,In_526,In_156);
nand U375 (N_375,In_782,In_611);
or U376 (N_376,In_75,In_5);
or U377 (N_377,In_20,In_318);
or U378 (N_378,In_536,In_331);
and U379 (N_379,In_61,In_340);
and U380 (N_380,In_496,In_13);
and U381 (N_381,In_731,In_936);
or U382 (N_382,In_497,In_304);
nand U383 (N_383,In_415,In_884);
nor U384 (N_384,In_785,In_399);
or U385 (N_385,In_467,In_8);
and U386 (N_386,In_699,In_881);
or U387 (N_387,In_862,In_414);
and U388 (N_388,In_113,In_726);
nand U389 (N_389,In_213,In_363);
nand U390 (N_390,In_353,In_575);
or U391 (N_391,In_972,In_324);
and U392 (N_392,In_893,In_755);
or U393 (N_393,In_477,In_315);
nor U394 (N_394,In_443,In_337);
nand U395 (N_395,In_250,In_578);
nor U396 (N_396,In_939,In_701);
nor U397 (N_397,In_849,In_99);
nor U398 (N_398,In_322,In_343);
or U399 (N_399,In_838,In_180);
and U400 (N_400,In_455,In_193);
nor U401 (N_401,In_567,In_845);
and U402 (N_402,In_349,In_169);
and U403 (N_403,In_732,In_789);
xnor U404 (N_404,In_683,In_385);
and U405 (N_405,In_321,In_333);
nor U406 (N_406,In_427,In_452);
nand U407 (N_407,In_618,In_528);
nor U408 (N_408,In_517,In_214);
or U409 (N_409,In_995,In_560);
xor U410 (N_410,In_234,In_457);
nor U411 (N_411,In_66,In_132);
nor U412 (N_412,In_918,In_282);
or U413 (N_413,In_285,In_587);
nand U414 (N_414,In_710,In_473);
nor U415 (N_415,In_554,In_698);
nand U416 (N_416,In_43,In_376);
and U417 (N_417,In_316,In_166);
nor U418 (N_418,In_325,In_41);
nand U419 (N_419,In_801,In_19);
nor U420 (N_420,In_582,In_606);
and U421 (N_421,In_266,In_879);
or U422 (N_422,In_805,In_25);
and U423 (N_423,In_130,In_594);
and U424 (N_424,In_486,In_334);
and U425 (N_425,In_681,In_390);
and U426 (N_426,In_825,In_950);
nor U427 (N_427,In_980,In_72);
and U428 (N_428,In_647,In_543);
nand U429 (N_429,In_733,In_946);
nor U430 (N_430,In_89,In_159);
nand U431 (N_431,In_137,In_352);
or U432 (N_432,In_273,In_997);
and U433 (N_433,In_803,In_423);
or U434 (N_434,In_900,In_437);
nand U435 (N_435,In_739,In_380);
nor U436 (N_436,In_109,In_197);
and U437 (N_437,In_73,In_689);
nor U438 (N_438,In_400,In_175);
nand U439 (N_439,In_716,In_781);
nor U440 (N_440,In_792,In_724);
and U441 (N_441,In_514,In_426);
and U442 (N_442,In_276,In_22);
or U443 (N_443,In_129,In_484);
nor U444 (N_444,In_910,In_928);
or U445 (N_445,In_952,In_372);
nand U446 (N_446,In_64,In_102);
nand U447 (N_447,In_574,In_47);
and U448 (N_448,In_530,In_787);
and U449 (N_449,In_115,In_976);
nand U450 (N_450,In_371,In_428);
and U451 (N_451,In_448,In_992);
nand U452 (N_452,In_831,In_81);
and U453 (N_453,In_886,In_150);
and U454 (N_454,In_449,In_135);
nand U455 (N_455,In_243,In_147);
nand U456 (N_456,In_492,In_548);
and U457 (N_457,In_797,In_556);
nor U458 (N_458,In_257,In_830);
nand U459 (N_459,In_923,In_50);
or U460 (N_460,In_730,In_857);
nand U461 (N_461,In_3,In_715);
nor U462 (N_462,In_816,In_153);
nor U463 (N_463,In_586,In_165);
nor U464 (N_464,In_810,In_866);
and U465 (N_465,In_351,In_44);
nor U466 (N_466,In_482,In_490);
nor U467 (N_467,In_576,In_943);
or U468 (N_468,In_306,In_678);
or U469 (N_469,In_993,In_774);
or U470 (N_470,In_752,In_902);
or U471 (N_471,In_861,In_453);
nor U472 (N_472,In_676,In_217);
and U473 (N_473,In_908,In_205);
nor U474 (N_474,In_247,In_45);
nor U475 (N_475,In_329,In_127);
and U476 (N_476,In_104,In_573);
or U477 (N_477,In_843,In_619);
or U478 (N_478,In_10,In_92);
nor U479 (N_479,In_565,In_896);
and U480 (N_480,In_253,In_786);
nor U481 (N_481,In_662,In_808);
nor U482 (N_482,In_308,In_812);
or U483 (N_483,In_295,In_523);
and U484 (N_484,In_495,In_907);
or U485 (N_485,In_508,In_309);
nor U486 (N_486,In_916,In_228);
and U487 (N_487,In_920,In_108);
and U488 (N_488,In_476,In_777);
and U489 (N_489,In_635,In_675);
or U490 (N_490,In_899,In_146);
xor U491 (N_491,In_2,In_798);
nand U492 (N_492,In_858,In_280);
nor U493 (N_493,In_728,In_832);
or U494 (N_494,In_76,In_630);
and U495 (N_495,In_398,In_814);
nor U496 (N_496,In_628,In_189);
nor U497 (N_497,In_949,In_237);
or U498 (N_498,In_209,In_909);
nand U499 (N_499,In_583,In_753);
nand U500 (N_500,In_55,In_595);
nor U501 (N_501,In_340,In_928);
nand U502 (N_502,In_871,In_323);
nor U503 (N_503,In_364,In_768);
and U504 (N_504,In_124,In_129);
nor U505 (N_505,In_45,In_828);
or U506 (N_506,In_487,In_184);
nor U507 (N_507,In_428,In_595);
and U508 (N_508,In_229,In_947);
or U509 (N_509,In_198,In_952);
and U510 (N_510,In_592,In_208);
or U511 (N_511,In_499,In_62);
and U512 (N_512,In_371,In_862);
nor U513 (N_513,In_261,In_96);
or U514 (N_514,In_323,In_884);
and U515 (N_515,In_844,In_341);
nor U516 (N_516,In_645,In_584);
nand U517 (N_517,In_168,In_140);
nand U518 (N_518,In_879,In_588);
and U519 (N_519,In_500,In_576);
or U520 (N_520,In_614,In_414);
and U521 (N_521,In_226,In_590);
or U522 (N_522,In_223,In_679);
xnor U523 (N_523,In_42,In_564);
and U524 (N_524,In_969,In_271);
or U525 (N_525,In_250,In_179);
nor U526 (N_526,In_306,In_20);
nand U527 (N_527,In_833,In_999);
nor U528 (N_528,In_788,In_344);
or U529 (N_529,In_851,In_313);
and U530 (N_530,In_365,In_721);
and U531 (N_531,In_766,In_162);
nor U532 (N_532,In_537,In_940);
nor U533 (N_533,In_891,In_965);
or U534 (N_534,In_29,In_624);
nand U535 (N_535,In_239,In_264);
nor U536 (N_536,In_470,In_269);
nand U537 (N_537,In_33,In_640);
or U538 (N_538,In_217,In_283);
nand U539 (N_539,In_587,In_946);
nor U540 (N_540,In_610,In_26);
nor U541 (N_541,In_621,In_117);
or U542 (N_542,In_409,In_431);
nor U543 (N_543,In_503,In_516);
or U544 (N_544,In_318,In_39);
and U545 (N_545,In_601,In_575);
nand U546 (N_546,In_355,In_621);
and U547 (N_547,In_714,In_463);
and U548 (N_548,In_9,In_65);
xor U549 (N_549,In_768,In_915);
and U550 (N_550,In_553,In_960);
nand U551 (N_551,In_851,In_531);
and U552 (N_552,In_298,In_647);
nand U553 (N_553,In_907,In_844);
nor U554 (N_554,In_791,In_828);
or U555 (N_555,In_311,In_443);
nand U556 (N_556,In_784,In_317);
and U557 (N_557,In_352,In_11);
or U558 (N_558,In_548,In_522);
or U559 (N_559,In_783,In_834);
nand U560 (N_560,In_889,In_721);
nand U561 (N_561,In_693,In_677);
nor U562 (N_562,In_345,In_944);
and U563 (N_563,In_178,In_629);
and U564 (N_564,In_202,In_601);
and U565 (N_565,In_822,In_361);
and U566 (N_566,In_769,In_422);
and U567 (N_567,In_283,In_279);
and U568 (N_568,In_602,In_857);
or U569 (N_569,In_40,In_262);
nand U570 (N_570,In_207,In_36);
and U571 (N_571,In_508,In_461);
or U572 (N_572,In_24,In_20);
or U573 (N_573,In_143,In_227);
nor U574 (N_574,In_893,In_275);
and U575 (N_575,In_961,In_62);
and U576 (N_576,In_288,In_587);
and U577 (N_577,In_483,In_931);
nor U578 (N_578,In_7,In_390);
nor U579 (N_579,In_371,In_145);
or U580 (N_580,In_211,In_581);
nand U581 (N_581,In_214,In_901);
or U582 (N_582,In_202,In_948);
nand U583 (N_583,In_451,In_729);
nor U584 (N_584,In_472,In_762);
nor U585 (N_585,In_965,In_19);
nor U586 (N_586,In_111,In_568);
and U587 (N_587,In_603,In_537);
and U588 (N_588,In_894,In_226);
and U589 (N_589,In_238,In_744);
nand U590 (N_590,In_880,In_377);
nand U591 (N_591,In_1,In_219);
or U592 (N_592,In_686,In_116);
nor U593 (N_593,In_348,In_861);
nand U594 (N_594,In_601,In_612);
nand U595 (N_595,In_422,In_499);
and U596 (N_596,In_594,In_10);
nor U597 (N_597,In_400,In_928);
and U598 (N_598,In_394,In_267);
or U599 (N_599,In_745,In_768);
nand U600 (N_600,In_341,In_96);
and U601 (N_601,In_67,In_710);
nor U602 (N_602,In_57,In_306);
and U603 (N_603,In_709,In_584);
and U604 (N_604,In_59,In_404);
nor U605 (N_605,In_857,In_656);
nor U606 (N_606,In_362,In_338);
nor U607 (N_607,In_620,In_437);
nor U608 (N_608,In_273,In_643);
nand U609 (N_609,In_914,In_810);
or U610 (N_610,In_703,In_930);
nor U611 (N_611,In_598,In_574);
nand U612 (N_612,In_87,In_228);
nor U613 (N_613,In_248,In_122);
xnor U614 (N_614,In_135,In_304);
nor U615 (N_615,In_192,In_208);
and U616 (N_616,In_261,In_780);
nor U617 (N_617,In_727,In_771);
and U618 (N_618,In_642,In_204);
or U619 (N_619,In_274,In_406);
nor U620 (N_620,In_578,In_471);
and U621 (N_621,In_816,In_830);
nor U622 (N_622,In_374,In_322);
nor U623 (N_623,In_510,In_30);
nor U624 (N_624,In_630,In_749);
nand U625 (N_625,In_792,In_159);
nor U626 (N_626,In_206,In_642);
nand U627 (N_627,In_282,In_299);
and U628 (N_628,In_164,In_209);
nor U629 (N_629,In_339,In_432);
nand U630 (N_630,In_60,In_825);
nor U631 (N_631,In_759,In_793);
nand U632 (N_632,In_750,In_942);
and U633 (N_633,In_404,In_119);
nand U634 (N_634,In_790,In_795);
and U635 (N_635,In_594,In_241);
or U636 (N_636,In_211,In_110);
nand U637 (N_637,In_954,In_854);
or U638 (N_638,In_634,In_742);
nor U639 (N_639,In_917,In_785);
and U640 (N_640,In_221,In_308);
nand U641 (N_641,In_206,In_104);
nand U642 (N_642,In_730,In_118);
nor U643 (N_643,In_110,In_485);
nand U644 (N_644,In_436,In_90);
nor U645 (N_645,In_428,In_597);
nand U646 (N_646,In_486,In_568);
nand U647 (N_647,In_933,In_673);
and U648 (N_648,In_876,In_25);
nor U649 (N_649,In_700,In_754);
and U650 (N_650,In_256,In_666);
or U651 (N_651,In_903,In_925);
or U652 (N_652,In_756,In_325);
nor U653 (N_653,In_326,In_722);
or U654 (N_654,In_255,In_174);
nand U655 (N_655,In_115,In_701);
or U656 (N_656,In_968,In_39);
and U657 (N_657,In_30,In_554);
nand U658 (N_658,In_389,In_185);
nand U659 (N_659,In_191,In_251);
nor U660 (N_660,In_50,In_87);
nand U661 (N_661,In_697,In_698);
and U662 (N_662,In_745,In_393);
or U663 (N_663,In_867,In_131);
nand U664 (N_664,In_225,In_434);
and U665 (N_665,In_134,In_63);
nor U666 (N_666,In_74,In_401);
nor U667 (N_667,In_556,In_552);
nand U668 (N_668,In_943,In_574);
and U669 (N_669,In_996,In_375);
xnor U670 (N_670,In_663,In_519);
or U671 (N_671,In_847,In_634);
and U672 (N_672,In_601,In_872);
and U673 (N_673,In_445,In_750);
or U674 (N_674,In_500,In_518);
or U675 (N_675,In_605,In_740);
nand U676 (N_676,In_504,In_175);
or U677 (N_677,In_126,In_465);
nand U678 (N_678,In_91,In_646);
nor U679 (N_679,In_682,In_345);
or U680 (N_680,In_453,In_47);
and U681 (N_681,In_561,In_942);
nor U682 (N_682,In_113,In_66);
or U683 (N_683,In_241,In_453);
nor U684 (N_684,In_450,In_517);
or U685 (N_685,In_847,In_7);
or U686 (N_686,In_847,In_44);
nor U687 (N_687,In_75,In_696);
or U688 (N_688,In_650,In_660);
xor U689 (N_689,In_482,In_385);
or U690 (N_690,In_62,In_860);
and U691 (N_691,In_123,In_917);
and U692 (N_692,In_264,In_485);
or U693 (N_693,In_33,In_166);
nand U694 (N_694,In_649,In_871);
or U695 (N_695,In_50,In_451);
and U696 (N_696,In_998,In_892);
or U697 (N_697,In_880,In_393);
nor U698 (N_698,In_670,In_175);
nor U699 (N_699,In_247,In_521);
or U700 (N_700,In_29,In_743);
nand U701 (N_701,In_368,In_856);
nand U702 (N_702,In_151,In_880);
and U703 (N_703,In_419,In_840);
nor U704 (N_704,In_42,In_957);
or U705 (N_705,In_949,In_540);
nand U706 (N_706,In_527,In_233);
nand U707 (N_707,In_403,In_707);
or U708 (N_708,In_193,In_21);
nor U709 (N_709,In_657,In_306);
nand U710 (N_710,In_485,In_824);
nand U711 (N_711,In_706,In_489);
or U712 (N_712,In_5,In_906);
nand U713 (N_713,In_573,In_909);
nor U714 (N_714,In_652,In_781);
nand U715 (N_715,In_972,In_158);
or U716 (N_716,In_754,In_456);
nor U717 (N_717,In_745,In_926);
nor U718 (N_718,In_503,In_447);
nand U719 (N_719,In_148,In_763);
nand U720 (N_720,In_681,In_30);
or U721 (N_721,In_878,In_151);
nor U722 (N_722,In_946,In_758);
nor U723 (N_723,In_258,In_245);
and U724 (N_724,In_72,In_981);
or U725 (N_725,In_86,In_277);
or U726 (N_726,In_377,In_828);
or U727 (N_727,In_700,In_545);
nor U728 (N_728,In_445,In_840);
nor U729 (N_729,In_667,In_359);
nor U730 (N_730,In_94,In_585);
or U731 (N_731,In_621,In_314);
nor U732 (N_732,In_95,In_11);
and U733 (N_733,In_745,In_365);
or U734 (N_734,In_377,In_327);
or U735 (N_735,In_451,In_509);
xor U736 (N_736,In_104,In_948);
nand U737 (N_737,In_296,In_203);
or U738 (N_738,In_567,In_837);
nand U739 (N_739,In_357,In_104);
nand U740 (N_740,In_825,In_171);
and U741 (N_741,In_90,In_792);
nor U742 (N_742,In_107,In_983);
or U743 (N_743,In_789,In_866);
or U744 (N_744,In_907,In_76);
or U745 (N_745,In_933,In_921);
nor U746 (N_746,In_332,In_341);
or U747 (N_747,In_749,In_704);
nand U748 (N_748,In_700,In_35);
or U749 (N_749,In_51,In_299);
or U750 (N_750,In_978,In_231);
nor U751 (N_751,In_901,In_34);
nand U752 (N_752,In_58,In_98);
and U753 (N_753,In_362,In_332);
nand U754 (N_754,In_254,In_801);
and U755 (N_755,In_193,In_935);
or U756 (N_756,In_72,In_510);
and U757 (N_757,In_870,In_115);
and U758 (N_758,In_114,In_213);
nand U759 (N_759,In_270,In_996);
or U760 (N_760,In_877,In_431);
nor U761 (N_761,In_377,In_288);
and U762 (N_762,In_927,In_403);
or U763 (N_763,In_929,In_86);
or U764 (N_764,In_537,In_350);
nor U765 (N_765,In_923,In_873);
and U766 (N_766,In_944,In_576);
or U767 (N_767,In_201,In_649);
nor U768 (N_768,In_300,In_362);
and U769 (N_769,In_67,In_243);
nor U770 (N_770,In_149,In_88);
nor U771 (N_771,In_68,In_920);
nand U772 (N_772,In_912,In_944);
nor U773 (N_773,In_625,In_279);
nand U774 (N_774,In_459,In_752);
nor U775 (N_775,In_639,In_67);
or U776 (N_776,In_202,In_331);
nand U777 (N_777,In_765,In_871);
or U778 (N_778,In_320,In_375);
or U779 (N_779,In_352,In_169);
and U780 (N_780,In_335,In_780);
and U781 (N_781,In_795,In_86);
or U782 (N_782,In_790,In_226);
or U783 (N_783,In_435,In_675);
nand U784 (N_784,In_216,In_118);
and U785 (N_785,In_891,In_747);
nor U786 (N_786,In_667,In_824);
nor U787 (N_787,In_648,In_686);
and U788 (N_788,In_744,In_978);
or U789 (N_789,In_199,In_377);
and U790 (N_790,In_279,In_169);
nand U791 (N_791,In_368,In_748);
nor U792 (N_792,In_880,In_684);
and U793 (N_793,In_671,In_856);
and U794 (N_794,In_939,In_678);
or U795 (N_795,In_564,In_474);
nand U796 (N_796,In_442,In_499);
or U797 (N_797,In_183,In_970);
and U798 (N_798,In_292,In_250);
nor U799 (N_799,In_442,In_112);
nand U800 (N_800,In_425,In_457);
nand U801 (N_801,In_662,In_387);
nor U802 (N_802,In_704,In_71);
nor U803 (N_803,In_792,In_770);
nand U804 (N_804,In_942,In_29);
nor U805 (N_805,In_114,In_564);
nor U806 (N_806,In_567,In_356);
nand U807 (N_807,In_984,In_337);
or U808 (N_808,In_706,In_756);
and U809 (N_809,In_813,In_355);
nand U810 (N_810,In_209,In_64);
nor U811 (N_811,In_317,In_497);
or U812 (N_812,In_155,In_470);
and U813 (N_813,In_967,In_346);
nand U814 (N_814,In_892,In_486);
and U815 (N_815,In_594,In_813);
or U816 (N_816,In_921,In_814);
or U817 (N_817,In_64,In_277);
nor U818 (N_818,In_954,In_876);
or U819 (N_819,In_936,In_29);
or U820 (N_820,In_809,In_348);
and U821 (N_821,In_369,In_612);
and U822 (N_822,In_620,In_495);
or U823 (N_823,In_759,In_81);
nor U824 (N_824,In_126,In_312);
and U825 (N_825,In_177,In_362);
or U826 (N_826,In_5,In_253);
or U827 (N_827,In_484,In_713);
and U828 (N_828,In_57,In_881);
nand U829 (N_829,In_545,In_398);
nor U830 (N_830,In_964,In_111);
nand U831 (N_831,In_295,In_62);
nor U832 (N_832,In_928,In_535);
nor U833 (N_833,In_333,In_538);
nor U834 (N_834,In_174,In_773);
or U835 (N_835,In_361,In_806);
or U836 (N_836,In_940,In_110);
or U837 (N_837,In_915,In_781);
nand U838 (N_838,In_78,In_898);
nor U839 (N_839,In_175,In_959);
nor U840 (N_840,In_0,In_356);
nand U841 (N_841,In_522,In_966);
and U842 (N_842,In_665,In_371);
xor U843 (N_843,In_303,In_884);
and U844 (N_844,In_214,In_838);
and U845 (N_845,In_677,In_863);
xnor U846 (N_846,In_964,In_88);
and U847 (N_847,In_955,In_551);
and U848 (N_848,In_878,In_540);
and U849 (N_849,In_459,In_864);
nor U850 (N_850,In_121,In_177);
or U851 (N_851,In_543,In_133);
nor U852 (N_852,In_230,In_81);
nor U853 (N_853,In_763,In_139);
nand U854 (N_854,In_715,In_165);
and U855 (N_855,In_358,In_413);
nor U856 (N_856,In_640,In_753);
or U857 (N_857,In_447,In_441);
and U858 (N_858,In_723,In_969);
or U859 (N_859,In_1,In_730);
and U860 (N_860,In_23,In_637);
or U861 (N_861,In_946,In_998);
nand U862 (N_862,In_718,In_210);
nor U863 (N_863,In_976,In_152);
nand U864 (N_864,In_130,In_288);
or U865 (N_865,In_839,In_993);
nor U866 (N_866,In_396,In_563);
nand U867 (N_867,In_777,In_292);
and U868 (N_868,In_615,In_767);
nand U869 (N_869,In_81,In_432);
and U870 (N_870,In_167,In_576);
and U871 (N_871,In_404,In_899);
or U872 (N_872,In_595,In_207);
nor U873 (N_873,In_635,In_480);
nor U874 (N_874,In_556,In_393);
or U875 (N_875,In_6,In_343);
or U876 (N_876,In_723,In_899);
and U877 (N_877,In_693,In_681);
nor U878 (N_878,In_289,In_247);
and U879 (N_879,In_55,In_36);
nand U880 (N_880,In_898,In_96);
or U881 (N_881,In_201,In_81);
nor U882 (N_882,In_543,In_331);
nand U883 (N_883,In_532,In_820);
or U884 (N_884,In_327,In_767);
or U885 (N_885,In_291,In_737);
or U886 (N_886,In_707,In_818);
nand U887 (N_887,In_264,In_634);
and U888 (N_888,In_952,In_846);
or U889 (N_889,In_430,In_784);
and U890 (N_890,In_609,In_664);
nand U891 (N_891,In_937,In_345);
nor U892 (N_892,In_877,In_582);
nand U893 (N_893,In_97,In_570);
or U894 (N_894,In_988,In_138);
nand U895 (N_895,In_511,In_39);
or U896 (N_896,In_220,In_32);
and U897 (N_897,In_39,In_862);
or U898 (N_898,In_945,In_399);
nand U899 (N_899,In_89,In_617);
or U900 (N_900,In_752,In_678);
or U901 (N_901,In_972,In_484);
nor U902 (N_902,In_479,In_550);
nand U903 (N_903,In_875,In_698);
nand U904 (N_904,In_802,In_919);
and U905 (N_905,In_320,In_200);
nand U906 (N_906,In_153,In_544);
nor U907 (N_907,In_769,In_269);
and U908 (N_908,In_144,In_624);
and U909 (N_909,In_619,In_31);
and U910 (N_910,In_272,In_745);
and U911 (N_911,In_203,In_938);
nor U912 (N_912,In_538,In_281);
and U913 (N_913,In_373,In_45);
and U914 (N_914,In_616,In_21);
nor U915 (N_915,In_87,In_555);
nand U916 (N_916,In_251,In_118);
or U917 (N_917,In_78,In_528);
or U918 (N_918,In_249,In_922);
nor U919 (N_919,In_662,In_945);
or U920 (N_920,In_864,In_482);
nand U921 (N_921,In_836,In_219);
and U922 (N_922,In_603,In_261);
or U923 (N_923,In_630,In_140);
nand U924 (N_924,In_281,In_713);
nand U925 (N_925,In_482,In_870);
and U926 (N_926,In_177,In_179);
nor U927 (N_927,In_959,In_493);
nor U928 (N_928,In_431,In_331);
or U929 (N_929,In_790,In_764);
and U930 (N_930,In_410,In_904);
nand U931 (N_931,In_532,In_495);
or U932 (N_932,In_957,In_175);
nor U933 (N_933,In_109,In_210);
or U934 (N_934,In_768,In_682);
nor U935 (N_935,In_948,In_244);
nor U936 (N_936,In_793,In_3);
nor U937 (N_937,In_960,In_859);
and U938 (N_938,In_8,In_330);
nand U939 (N_939,In_710,In_575);
nor U940 (N_940,In_307,In_956);
nor U941 (N_941,In_24,In_215);
nor U942 (N_942,In_61,In_455);
and U943 (N_943,In_160,In_261);
or U944 (N_944,In_56,In_536);
or U945 (N_945,In_298,In_507);
xnor U946 (N_946,In_817,In_70);
and U947 (N_947,In_29,In_345);
or U948 (N_948,In_792,In_639);
nand U949 (N_949,In_603,In_291);
nor U950 (N_950,In_12,In_188);
and U951 (N_951,In_737,In_799);
nand U952 (N_952,In_708,In_201);
or U953 (N_953,In_157,In_277);
or U954 (N_954,In_461,In_385);
or U955 (N_955,In_864,In_297);
nor U956 (N_956,In_466,In_154);
or U957 (N_957,In_745,In_698);
and U958 (N_958,In_391,In_290);
nor U959 (N_959,In_672,In_815);
nand U960 (N_960,In_230,In_645);
nor U961 (N_961,In_150,In_120);
nor U962 (N_962,In_397,In_336);
and U963 (N_963,In_98,In_249);
and U964 (N_964,In_562,In_126);
nand U965 (N_965,In_419,In_907);
nor U966 (N_966,In_967,In_618);
nor U967 (N_967,In_861,In_881);
and U968 (N_968,In_815,In_230);
nor U969 (N_969,In_753,In_818);
and U970 (N_970,In_462,In_114);
and U971 (N_971,In_962,In_440);
nand U972 (N_972,In_777,In_712);
nor U973 (N_973,In_631,In_228);
nand U974 (N_974,In_807,In_859);
nand U975 (N_975,In_585,In_468);
nor U976 (N_976,In_211,In_371);
or U977 (N_977,In_814,In_322);
and U978 (N_978,In_519,In_829);
nor U979 (N_979,In_208,In_819);
nand U980 (N_980,In_336,In_258);
and U981 (N_981,In_147,In_21);
and U982 (N_982,In_859,In_100);
and U983 (N_983,In_323,In_333);
or U984 (N_984,In_223,In_193);
or U985 (N_985,In_775,In_458);
nor U986 (N_986,In_744,In_137);
and U987 (N_987,In_146,In_314);
or U988 (N_988,In_907,In_340);
and U989 (N_989,In_226,In_347);
and U990 (N_990,In_943,In_722);
nor U991 (N_991,In_917,In_847);
nand U992 (N_992,In_511,In_801);
and U993 (N_993,In_176,In_663);
or U994 (N_994,In_360,In_168);
or U995 (N_995,In_818,In_351);
nand U996 (N_996,In_831,In_251);
nor U997 (N_997,In_740,In_981);
nor U998 (N_998,In_441,In_299);
or U999 (N_999,In_852,In_250);
or U1000 (N_1000,In_319,In_415);
nand U1001 (N_1001,In_809,In_697);
nand U1002 (N_1002,In_752,In_865);
or U1003 (N_1003,In_536,In_860);
and U1004 (N_1004,In_482,In_207);
or U1005 (N_1005,In_785,In_955);
or U1006 (N_1006,In_946,In_718);
or U1007 (N_1007,In_485,In_270);
nand U1008 (N_1008,In_80,In_677);
nand U1009 (N_1009,In_443,In_88);
nand U1010 (N_1010,In_102,In_301);
nor U1011 (N_1011,In_156,In_491);
nor U1012 (N_1012,In_442,In_638);
nand U1013 (N_1013,In_789,In_366);
nor U1014 (N_1014,In_912,In_713);
nor U1015 (N_1015,In_141,In_509);
or U1016 (N_1016,In_561,In_825);
and U1017 (N_1017,In_29,In_32);
or U1018 (N_1018,In_550,In_928);
or U1019 (N_1019,In_341,In_123);
nor U1020 (N_1020,In_580,In_551);
nor U1021 (N_1021,In_634,In_481);
and U1022 (N_1022,In_351,In_252);
or U1023 (N_1023,In_687,In_641);
nand U1024 (N_1024,In_446,In_898);
or U1025 (N_1025,In_781,In_859);
nor U1026 (N_1026,In_817,In_104);
nand U1027 (N_1027,In_779,In_878);
nor U1028 (N_1028,In_566,In_29);
nand U1029 (N_1029,In_673,In_903);
and U1030 (N_1030,In_12,In_292);
nand U1031 (N_1031,In_786,In_661);
or U1032 (N_1032,In_962,In_688);
nand U1033 (N_1033,In_892,In_393);
nand U1034 (N_1034,In_879,In_511);
or U1035 (N_1035,In_681,In_527);
nand U1036 (N_1036,In_126,In_326);
nor U1037 (N_1037,In_43,In_649);
and U1038 (N_1038,In_316,In_593);
xnor U1039 (N_1039,In_58,In_697);
xor U1040 (N_1040,In_107,In_862);
and U1041 (N_1041,In_87,In_267);
and U1042 (N_1042,In_165,In_886);
and U1043 (N_1043,In_334,In_154);
nor U1044 (N_1044,In_526,In_896);
nor U1045 (N_1045,In_87,In_471);
and U1046 (N_1046,In_594,In_201);
nor U1047 (N_1047,In_472,In_603);
and U1048 (N_1048,In_62,In_148);
or U1049 (N_1049,In_136,In_543);
or U1050 (N_1050,In_912,In_135);
or U1051 (N_1051,In_698,In_408);
xnor U1052 (N_1052,In_70,In_122);
and U1053 (N_1053,In_303,In_163);
nand U1054 (N_1054,In_66,In_251);
or U1055 (N_1055,In_178,In_715);
nand U1056 (N_1056,In_571,In_799);
or U1057 (N_1057,In_144,In_426);
nand U1058 (N_1058,In_2,In_222);
or U1059 (N_1059,In_224,In_497);
nand U1060 (N_1060,In_612,In_911);
nor U1061 (N_1061,In_27,In_334);
or U1062 (N_1062,In_666,In_613);
nor U1063 (N_1063,In_897,In_633);
or U1064 (N_1064,In_338,In_830);
nand U1065 (N_1065,In_279,In_168);
and U1066 (N_1066,In_533,In_357);
nand U1067 (N_1067,In_89,In_616);
or U1068 (N_1068,In_771,In_980);
and U1069 (N_1069,In_335,In_592);
nor U1070 (N_1070,In_694,In_7);
and U1071 (N_1071,In_533,In_475);
and U1072 (N_1072,In_825,In_296);
or U1073 (N_1073,In_415,In_501);
and U1074 (N_1074,In_415,In_389);
or U1075 (N_1075,In_709,In_796);
nor U1076 (N_1076,In_448,In_912);
and U1077 (N_1077,In_92,In_349);
or U1078 (N_1078,In_873,In_217);
and U1079 (N_1079,In_859,In_414);
or U1080 (N_1080,In_487,In_733);
or U1081 (N_1081,In_609,In_98);
and U1082 (N_1082,In_364,In_841);
or U1083 (N_1083,In_342,In_549);
nand U1084 (N_1084,In_590,In_787);
and U1085 (N_1085,In_328,In_749);
nor U1086 (N_1086,In_568,In_989);
nor U1087 (N_1087,In_162,In_980);
nor U1088 (N_1088,In_771,In_382);
and U1089 (N_1089,In_370,In_103);
nand U1090 (N_1090,In_717,In_120);
or U1091 (N_1091,In_102,In_498);
or U1092 (N_1092,In_408,In_308);
nor U1093 (N_1093,In_454,In_840);
nand U1094 (N_1094,In_345,In_558);
or U1095 (N_1095,In_609,In_932);
or U1096 (N_1096,In_873,In_220);
nor U1097 (N_1097,In_800,In_0);
or U1098 (N_1098,In_217,In_73);
and U1099 (N_1099,In_454,In_308);
xor U1100 (N_1100,In_997,In_763);
or U1101 (N_1101,In_104,In_176);
nand U1102 (N_1102,In_815,In_315);
and U1103 (N_1103,In_527,In_497);
nor U1104 (N_1104,In_274,In_759);
nand U1105 (N_1105,In_849,In_115);
nor U1106 (N_1106,In_889,In_34);
or U1107 (N_1107,In_870,In_561);
nor U1108 (N_1108,In_577,In_342);
nor U1109 (N_1109,In_418,In_146);
nor U1110 (N_1110,In_853,In_463);
or U1111 (N_1111,In_419,In_42);
nor U1112 (N_1112,In_645,In_531);
and U1113 (N_1113,In_448,In_913);
nor U1114 (N_1114,In_528,In_307);
nor U1115 (N_1115,In_675,In_926);
or U1116 (N_1116,In_290,In_305);
nor U1117 (N_1117,In_785,In_209);
nand U1118 (N_1118,In_742,In_275);
nand U1119 (N_1119,In_417,In_59);
or U1120 (N_1120,In_659,In_89);
nand U1121 (N_1121,In_550,In_967);
or U1122 (N_1122,In_107,In_659);
nor U1123 (N_1123,In_694,In_559);
or U1124 (N_1124,In_633,In_415);
or U1125 (N_1125,In_807,In_707);
and U1126 (N_1126,In_424,In_156);
or U1127 (N_1127,In_227,In_727);
nor U1128 (N_1128,In_790,In_103);
or U1129 (N_1129,In_90,In_209);
nor U1130 (N_1130,In_881,In_963);
nand U1131 (N_1131,In_561,In_327);
xor U1132 (N_1132,In_737,In_493);
nand U1133 (N_1133,In_539,In_682);
nand U1134 (N_1134,In_155,In_459);
and U1135 (N_1135,In_311,In_645);
nand U1136 (N_1136,In_436,In_168);
or U1137 (N_1137,In_932,In_981);
and U1138 (N_1138,In_760,In_213);
nand U1139 (N_1139,In_79,In_891);
nor U1140 (N_1140,In_435,In_947);
or U1141 (N_1141,In_791,In_433);
and U1142 (N_1142,In_36,In_879);
nor U1143 (N_1143,In_613,In_207);
or U1144 (N_1144,In_47,In_855);
or U1145 (N_1145,In_298,In_728);
and U1146 (N_1146,In_502,In_861);
or U1147 (N_1147,In_911,In_751);
nand U1148 (N_1148,In_988,In_463);
nand U1149 (N_1149,In_682,In_775);
nand U1150 (N_1150,In_961,In_170);
nor U1151 (N_1151,In_418,In_60);
or U1152 (N_1152,In_700,In_195);
and U1153 (N_1153,In_159,In_633);
or U1154 (N_1154,In_894,In_425);
and U1155 (N_1155,In_250,In_271);
nor U1156 (N_1156,In_329,In_435);
nor U1157 (N_1157,In_928,In_886);
or U1158 (N_1158,In_993,In_27);
or U1159 (N_1159,In_483,In_911);
and U1160 (N_1160,In_959,In_839);
nand U1161 (N_1161,In_269,In_761);
and U1162 (N_1162,In_592,In_609);
and U1163 (N_1163,In_206,In_269);
or U1164 (N_1164,In_272,In_414);
nand U1165 (N_1165,In_215,In_443);
nand U1166 (N_1166,In_417,In_878);
and U1167 (N_1167,In_16,In_460);
and U1168 (N_1168,In_857,In_792);
or U1169 (N_1169,In_288,In_771);
nand U1170 (N_1170,In_545,In_327);
nand U1171 (N_1171,In_940,In_708);
xnor U1172 (N_1172,In_864,In_878);
or U1173 (N_1173,In_456,In_784);
or U1174 (N_1174,In_132,In_170);
nor U1175 (N_1175,In_377,In_308);
or U1176 (N_1176,In_455,In_338);
nor U1177 (N_1177,In_61,In_992);
nand U1178 (N_1178,In_712,In_561);
or U1179 (N_1179,In_129,In_477);
or U1180 (N_1180,In_372,In_979);
nor U1181 (N_1181,In_449,In_759);
nand U1182 (N_1182,In_683,In_289);
nor U1183 (N_1183,In_13,In_408);
or U1184 (N_1184,In_370,In_636);
nand U1185 (N_1185,In_872,In_758);
nand U1186 (N_1186,In_920,In_613);
or U1187 (N_1187,In_213,In_574);
nor U1188 (N_1188,In_706,In_289);
nor U1189 (N_1189,In_954,In_536);
nand U1190 (N_1190,In_606,In_510);
nand U1191 (N_1191,In_19,In_968);
nand U1192 (N_1192,In_143,In_870);
nand U1193 (N_1193,In_422,In_336);
and U1194 (N_1194,In_97,In_86);
nand U1195 (N_1195,In_112,In_134);
nand U1196 (N_1196,In_238,In_489);
nor U1197 (N_1197,In_797,In_921);
and U1198 (N_1198,In_461,In_740);
or U1199 (N_1199,In_992,In_317);
nand U1200 (N_1200,In_794,In_81);
nor U1201 (N_1201,In_325,In_734);
nor U1202 (N_1202,In_820,In_547);
or U1203 (N_1203,In_813,In_246);
or U1204 (N_1204,In_361,In_149);
nor U1205 (N_1205,In_105,In_474);
and U1206 (N_1206,In_580,In_86);
nand U1207 (N_1207,In_958,In_972);
nand U1208 (N_1208,In_944,In_634);
or U1209 (N_1209,In_14,In_944);
or U1210 (N_1210,In_689,In_491);
nor U1211 (N_1211,In_309,In_81);
nand U1212 (N_1212,In_943,In_331);
and U1213 (N_1213,In_818,In_584);
nor U1214 (N_1214,In_43,In_946);
nor U1215 (N_1215,In_343,In_790);
or U1216 (N_1216,In_933,In_655);
xnor U1217 (N_1217,In_130,In_49);
nor U1218 (N_1218,In_393,In_894);
and U1219 (N_1219,In_639,In_796);
nand U1220 (N_1220,In_717,In_720);
or U1221 (N_1221,In_578,In_518);
nand U1222 (N_1222,In_668,In_127);
nand U1223 (N_1223,In_105,In_430);
and U1224 (N_1224,In_841,In_171);
and U1225 (N_1225,In_155,In_635);
or U1226 (N_1226,In_623,In_97);
nand U1227 (N_1227,In_276,In_320);
or U1228 (N_1228,In_280,In_775);
and U1229 (N_1229,In_517,In_715);
and U1230 (N_1230,In_651,In_324);
xor U1231 (N_1231,In_850,In_930);
nor U1232 (N_1232,In_126,In_711);
nand U1233 (N_1233,In_745,In_537);
nor U1234 (N_1234,In_217,In_377);
nor U1235 (N_1235,In_570,In_581);
and U1236 (N_1236,In_793,In_900);
nand U1237 (N_1237,In_519,In_947);
or U1238 (N_1238,In_61,In_403);
and U1239 (N_1239,In_630,In_2);
or U1240 (N_1240,In_166,In_459);
nor U1241 (N_1241,In_183,In_150);
nand U1242 (N_1242,In_509,In_900);
and U1243 (N_1243,In_727,In_439);
and U1244 (N_1244,In_137,In_832);
nand U1245 (N_1245,In_786,In_654);
and U1246 (N_1246,In_482,In_945);
nand U1247 (N_1247,In_313,In_775);
or U1248 (N_1248,In_366,In_131);
or U1249 (N_1249,In_108,In_558);
and U1250 (N_1250,In_914,In_875);
or U1251 (N_1251,In_371,In_158);
nor U1252 (N_1252,In_367,In_878);
and U1253 (N_1253,In_303,In_809);
and U1254 (N_1254,In_709,In_705);
nor U1255 (N_1255,In_21,In_366);
nor U1256 (N_1256,In_367,In_159);
or U1257 (N_1257,In_522,In_334);
and U1258 (N_1258,In_357,In_365);
nand U1259 (N_1259,In_98,In_771);
xnor U1260 (N_1260,In_232,In_478);
nor U1261 (N_1261,In_855,In_689);
and U1262 (N_1262,In_193,In_444);
and U1263 (N_1263,In_301,In_31);
nand U1264 (N_1264,In_570,In_190);
nor U1265 (N_1265,In_225,In_436);
nor U1266 (N_1266,In_17,In_758);
and U1267 (N_1267,In_869,In_183);
nand U1268 (N_1268,In_699,In_819);
nor U1269 (N_1269,In_895,In_348);
nor U1270 (N_1270,In_177,In_194);
nor U1271 (N_1271,In_808,In_618);
or U1272 (N_1272,In_671,In_300);
or U1273 (N_1273,In_622,In_142);
nand U1274 (N_1274,In_896,In_101);
or U1275 (N_1275,In_527,In_576);
nand U1276 (N_1276,In_393,In_921);
or U1277 (N_1277,In_567,In_686);
and U1278 (N_1278,In_71,In_275);
and U1279 (N_1279,In_424,In_255);
or U1280 (N_1280,In_215,In_634);
and U1281 (N_1281,In_660,In_407);
and U1282 (N_1282,In_861,In_199);
nor U1283 (N_1283,In_236,In_798);
nor U1284 (N_1284,In_740,In_860);
and U1285 (N_1285,In_160,In_25);
or U1286 (N_1286,In_37,In_266);
nand U1287 (N_1287,In_811,In_472);
nor U1288 (N_1288,In_515,In_170);
nand U1289 (N_1289,In_156,In_90);
or U1290 (N_1290,In_435,In_855);
nor U1291 (N_1291,In_954,In_949);
nand U1292 (N_1292,In_305,In_767);
nand U1293 (N_1293,In_836,In_533);
and U1294 (N_1294,In_29,In_337);
and U1295 (N_1295,In_229,In_665);
nand U1296 (N_1296,In_133,In_419);
or U1297 (N_1297,In_816,In_801);
nand U1298 (N_1298,In_910,In_907);
or U1299 (N_1299,In_840,In_463);
nor U1300 (N_1300,In_202,In_5);
xnor U1301 (N_1301,In_718,In_342);
and U1302 (N_1302,In_48,In_767);
nand U1303 (N_1303,In_63,In_28);
or U1304 (N_1304,In_133,In_95);
nor U1305 (N_1305,In_802,In_868);
and U1306 (N_1306,In_868,In_979);
nand U1307 (N_1307,In_814,In_496);
or U1308 (N_1308,In_848,In_275);
nand U1309 (N_1309,In_565,In_536);
nor U1310 (N_1310,In_391,In_820);
or U1311 (N_1311,In_934,In_575);
nor U1312 (N_1312,In_515,In_736);
nand U1313 (N_1313,In_255,In_893);
nand U1314 (N_1314,In_492,In_29);
and U1315 (N_1315,In_376,In_759);
or U1316 (N_1316,In_2,In_638);
or U1317 (N_1317,In_55,In_570);
and U1318 (N_1318,In_408,In_261);
nand U1319 (N_1319,In_858,In_599);
and U1320 (N_1320,In_912,In_215);
and U1321 (N_1321,In_920,In_522);
nand U1322 (N_1322,In_7,In_500);
nor U1323 (N_1323,In_534,In_797);
nor U1324 (N_1324,In_70,In_58);
nor U1325 (N_1325,In_647,In_755);
nand U1326 (N_1326,In_882,In_112);
or U1327 (N_1327,In_884,In_525);
nand U1328 (N_1328,In_494,In_797);
nor U1329 (N_1329,In_130,In_705);
and U1330 (N_1330,In_125,In_584);
nand U1331 (N_1331,In_664,In_409);
and U1332 (N_1332,In_473,In_980);
nand U1333 (N_1333,In_31,In_34);
or U1334 (N_1334,In_932,In_164);
nand U1335 (N_1335,In_532,In_109);
or U1336 (N_1336,In_786,In_738);
nor U1337 (N_1337,In_258,In_406);
nor U1338 (N_1338,In_362,In_305);
nand U1339 (N_1339,In_498,In_705);
or U1340 (N_1340,In_130,In_107);
nand U1341 (N_1341,In_570,In_535);
or U1342 (N_1342,In_693,In_464);
nor U1343 (N_1343,In_62,In_893);
and U1344 (N_1344,In_494,In_191);
nand U1345 (N_1345,In_105,In_464);
or U1346 (N_1346,In_6,In_280);
nor U1347 (N_1347,In_928,In_568);
or U1348 (N_1348,In_685,In_164);
or U1349 (N_1349,In_487,In_766);
nand U1350 (N_1350,In_855,In_37);
and U1351 (N_1351,In_169,In_791);
and U1352 (N_1352,In_520,In_172);
nor U1353 (N_1353,In_501,In_366);
nand U1354 (N_1354,In_893,In_721);
or U1355 (N_1355,In_640,In_440);
nand U1356 (N_1356,In_837,In_450);
or U1357 (N_1357,In_136,In_732);
nor U1358 (N_1358,In_376,In_11);
or U1359 (N_1359,In_530,In_716);
xnor U1360 (N_1360,In_550,In_916);
or U1361 (N_1361,In_266,In_111);
nand U1362 (N_1362,In_993,In_293);
and U1363 (N_1363,In_87,In_335);
nand U1364 (N_1364,In_335,In_32);
or U1365 (N_1365,In_425,In_220);
and U1366 (N_1366,In_498,In_759);
nand U1367 (N_1367,In_908,In_689);
and U1368 (N_1368,In_841,In_333);
or U1369 (N_1369,In_349,In_882);
nor U1370 (N_1370,In_634,In_784);
or U1371 (N_1371,In_875,In_181);
nor U1372 (N_1372,In_763,In_89);
and U1373 (N_1373,In_749,In_191);
nand U1374 (N_1374,In_244,In_672);
and U1375 (N_1375,In_641,In_420);
and U1376 (N_1376,In_101,In_748);
or U1377 (N_1377,In_516,In_200);
nor U1378 (N_1378,In_154,In_779);
nor U1379 (N_1379,In_956,In_364);
nand U1380 (N_1380,In_48,In_817);
and U1381 (N_1381,In_892,In_162);
nor U1382 (N_1382,In_243,In_834);
nor U1383 (N_1383,In_977,In_243);
nand U1384 (N_1384,In_133,In_879);
and U1385 (N_1385,In_528,In_731);
and U1386 (N_1386,In_442,In_674);
nand U1387 (N_1387,In_156,In_474);
or U1388 (N_1388,In_23,In_228);
nor U1389 (N_1389,In_615,In_109);
or U1390 (N_1390,In_514,In_696);
nor U1391 (N_1391,In_684,In_606);
and U1392 (N_1392,In_237,In_738);
or U1393 (N_1393,In_700,In_491);
and U1394 (N_1394,In_28,In_624);
xnor U1395 (N_1395,In_53,In_939);
or U1396 (N_1396,In_891,In_336);
nand U1397 (N_1397,In_548,In_737);
nor U1398 (N_1398,In_213,In_318);
nand U1399 (N_1399,In_758,In_937);
nor U1400 (N_1400,In_982,In_517);
nor U1401 (N_1401,In_38,In_417);
nand U1402 (N_1402,In_754,In_334);
nor U1403 (N_1403,In_352,In_583);
or U1404 (N_1404,In_812,In_20);
nor U1405 (N_1405,In_555,In_45);
or U1406 (N_1406,In_584,In_27);
nand U1407 (N_1407,In_619,In_465);
and U1408 (N_1408,In_667,In_858);
or U1409 (N_1409,In_707,In_307);
or U1410 (N_1410,In_597,In_910);
or U1411 (N_1411,In_578,In_757);
nor U1412 (N_1412,In_606,In_3);
or U1413 (N_1413,In_824,In_842);
nand U1414 (N_1414,In_270,In_563);
nand U1415 (N_1415,In_821,In_452);
nand U1416 (N_1416,In_28,In_926);
and U1417 (N_1417,In_80,In_896);
nand U1418 (N_1418,In_139,In_635);
or U1419 (N_1419,In_163,In_105);
and U1420 (N_1420,In_652,In_220);
nand U1421 (N_1421,In_710,In_68);
and U1422 (N_1422,In_390,In_46);
nor U1423 (N_1423,In_701,In_127);
nand U1424 (N_1424,In_674,In_267);
nand U1425 (N_1425,In_837,In_323);
or U1426 (N_1426,In_982,In_509);
and U1427 (N_1427,In_907,In_459);
nor U1428 (N_1428,In_56,In_649);
nand U1429 (N_1429,In_307,In_791);
nor U1430 (N_1430,In_967,In_421);
nor U1431 (N_1431,In_397,In_216);
and U1432 (N_1432,In_666,In_311);
nor U1433 (N_1433,In_988,In_882);
nand U1434 (N_1434,In_605,In_69);
nor U1435 (N_1435,In_359,In_542);
and U1436 (N_1436,In_219,In_363);
or U1437 (N_1437,In_552,In_703);
or U1438 (N_1438,In_349,In_669);
or U1439 (N_1439,In_406,In_112);
and U1440 (N_1440,In_847,In_616);
nor U1441 (N_1441,In_94,In_276);
nand U1442 (N_1442,In_684,In_552);
or U1443 (N_1443,In_797,In_615);
nor U1444 (N_1444,In_677,In_184);
nor U1445 (N_1445,In_54,In_337);
nor U1446 (N_1446,In_729,In_936);
or U1447 (N_1447,In_633,In_795);
or U1448 (N_1448,In_552,In_557);
or U1449 (N_1449,In_241,In_228);
and U1450 (N_1450,In_989,In_377);
nand U1451 (N_1451,In_692,In_512);
and U1452 (N_1452,In_632,In_838);
and U1453 (N_1453,In_98,In_323);
nor U1454 (N_1454,In_585,In_904);
and U1455 (N_1455,In_20,In_722);
and U1456 (N_1456,In_391,In_454);
or U1457 (N_1457,In_218,In_748);
or U1458 (N_1458,In_952,In_378);
nor U1459 (N_1459,In_264,In_985);
and U1460 (N_1460,In_62,In_706);
nor U1461 (N_1461,In_140,In_892);
xor U1462 (N_1462,In_28,In_374);
nand U1463 (N_1463,In_232,In_364);
or U1464 (N_1464,In_902,In_889);
nor U1465 (N_1465,In_543,In_548);
and U1466 (N_1466,In_362,In_108);
and U1467 (N_1467,In_998,In_174);
or U1468 (N_1468,In_281,In_945);
nand U1469 (N_1469,In_320,In_422);
nor U1470 (N_1470,In_305,In_944);
and U1471 (N_1471,In_158,In_552);
nand U1472 (N_1472,In_437,In_431);
nor U1473 (N_1473,In_103,In_822);
and U1474 (N_1474,In_607,In_344);
nor U1475 (N_1475,In_418,In_504);
nand U1476 (N_1476,In_85,In_338);
nand U1477 (N_1477,In_332,In_479);
or U1478 (N_1478,In_900,In_780);
nor U1479 (N_1479,In_883,In_877);
or U1480 (N_1480,In_775,In_477);
nand U1481 (N_1481,In_742,In_361);
and U1482 (N_1482,In_886,In_568);
nand U1483 (N_1483,In_647,In_996);
and U1484 (N_1484,In_648,In_115);
and U1485 (N_1485,In_849,In_402);
xor U1486 (N_1486,In_837,In_591);
nand U1487 (N_1487,In_587,In_500);
nor U1488 (N_1488,In_281,In_907);
or U1489 (N_1489,In_914,In_414);
or U1490 (N_1490,In_157,In_184);
nand U1491 (N_1491,In_694,In_232);
and U1492 (N_1492,In_795,In_218);
nand U1493 (N_1493,In_659,In_521);
nand U1494 (N_1494,In_852,In_100);
xnor U1495 (N_1495,In_477,In_893);
or U1496 (N_1496,In_10,In_83);
nor U1497 (N_1497,In_430,In_322);
and U1498 (N_1498,In_872,In_185);
and U1499 (N_1499,In_72,In_459);
and U1500 (N_1500,In_462,In_432);
and U1501 (N_1501,In_898,In_320);
nand U1502 (N_1502,In_987,In_333);
nor U1503 (N_1503,In_202,In_62);
or U1504 (N_1504,In_442,In_648);
and U1505 (N_1505,In_568,In_625);
and U1506 (N_1506,In_977,In_434);
or U1507 (N_1507,In_104,In_491);
nor U1508 (N_1508,In_3,In_547);
nand U1509 (N_1509,In_722,In_58);
and U1510 (N_1510,In_977,In_601);
nor U1511 (N_1511,In_437,In_405);
and U1512 (N_1512,In_331,In_646);
nor U1513 (N_1513,In_860,In_763);
or U1514 (N_1514,In_299,In_61);
or U1515 (N_1515,In_42,In_532);
nand U1516 (N_1516,In_706,In_986);
and U1517 (N_1517,In_25,In_268);
and U1518 (N_1518,In_78,In_902);
nand U1519 (N_1519,In_953,In_869);
nor U1520 (N_1520,In_659,In_2);
nor U1521 (N_1521,In_484,In_553);
and U1522 (N_1522,In_220,In_771);
and U1523 (N_1523,In_165,In_822);
or U1524 (N_1524,In_164,In_379);
nand U1525 (N_1525,In_361,In_86);
nor U1526 (N_1526,In_556,In_100);
or U1527 (N_1527,In_814,In_924);
nand U1528 (N_1528,In_335,In_432);
nand U1529 (N_1529,In_142,In_599);
nand U1530 (N_1530,In_609,In_631);
and U1531 (N_1531,In_81,In_660);
nor U1532 (N_1532,In_740,In_912);
nand U1533 (N_1533,In_486,In_659);
and U1534 (N_1534,In_596,In_779);
or U1535 (N_1535,In_770,In_873);
nor U1536 (N_1536,In_979,In_762);
nor U1537 (N_1537,In_947,In_574);
nand U1538 (N_1538,In_73,In_486);
nand U1539 (N_1539,In_613,In_110);
or U1540 (N_1540,In_651,In_662);
and U1541 (N_1541,In_21,In_214);
nand U1542 (N_1542,In_10,In_692);
nand U1543 (N_1543,In_712,In_120);
and U1544 (N_1544,In_142,In_82);
nand U1545 (N_1545,In_775,In_65);
nand U1546 (N_1546,In_253,In_734);
and U1547 (N_1547,In_137,In_363);
and U1548 (N_1548,In_278,In_656);
and U1549 (N_1549,In_440,In_995);
nor U1550 (N_1550,In_89,In_531);
nor U1551 (N_1551,In_854,In_62);
or U1552 (N_1552,In_963,In_855);
nor U1553 (N_1553,In_960,In_563);
or U1554 (N_1554,In_786,In_896);
and U1555 (N_1555,In_604,In_928);
and U1556 (N_1556,In_256,In_187);
and U1557 (N_1557,In_205,In_979);
or U1558 (N_1558,In_536,In_119);
nor U1559 (N_1559,In_512,In_860);
or U1560 (N_1560,In_631,In_796);
nor U1561 (N_1561,In_685,In_186);
nor U1562 (N_1562,In_692,In_61);
and U1563 (N_1563,In_290,In_751);
nor U1564 (N_1564,In_225,In_709);
and U1565 (N_1565,In_348,In_620);
nor U1566 (N_1566,In_48,In_993);
nor U1567 (N_1567,In_490,In_171);
and U1568 (N_1568,In_850,In_100);
or U1569 (N_1569,In_499,In_33);
nor U1570 (N_1570,In_602,In_103);
and U1571 (N_1571,In_54,In_280);
and U1572 (N_1572,In_373,In_726);
and U1573 (N_1573,In_638,In_538);
nor U1574 (N_1574,In_364,In_322);
nand U1575 (N_1575,In_178,In_475);
and U1576 (N_1576,In_703,In_273);
nand U1577 (N_1577,In_888,In_585);
or U1578 (N_1578,In_891,In_875);
nor U1579 (N_1579,In_458,In_19);
nand U1580 (N_1580,In_680,In_51);
nand U1581 (N_1581,In_405,In_892);
nand U1582 (N_1582,In_755,In_386);
nand U1583 (N_1583,In_608,In_719);
nor U1584 (N_1584,In_357,In_150);
and U1585 (N_1585,In_99,In_78);
nor U1586 (N_1586,In_722,In_570);
nand U1587 (N_1587,In_867,In_92);
nor U1588 (N_1588,In_736,In_566);
and U1589 (N_1589,In_120,In_72);
nand U1590 (N_1590,In_492,In_542);
or U1591 (N_1591,In_150,In_153);
and U1592 (N_1592,In_622,In_348);
nand U1593 (N_1593,In_169,In_65);
and U1594 (N_1594,In_159,In_279);
nand U1595 (N_1595,In_284,In_670);
or U1596 (N_1596,In_651,In_484);
nand U1597 (N_1597,In_480,In_39);
or U1598 (N_1598,In_885,In_223);
or U1599 (N_1599,In_695,In_100);
nor U1600 (N_1600,In_651,In_956);
and U1601 (N_1601,In_383,In_86);
nor U1602 (N_1602,In_298,In_141);
or U1603 (N_1603,In_330,In_786);
and U1604 (N_1604,In_834,In_435);
or U1605 (N_1605,In_651,In_357);
nand U1606 (N_1606,In_666,In_100);
nor U1607 (N_1607,In_690,In_339);
nor U1608 (N_1608,In_315,In_690);
and U1609 (N_1609,In_754,In_908);
nand U1610 (N_1610,In_622,In_841);
or U1611 (N_1611,In_791,In_82);
nand U1612 (N_1612,In_824,In_759);
xor U1613 (N_1613,In_265,In_417);
nor U1614 (N_1614,In_524,In_105);
or U1615 (N_1615,In_634,In_687);
nand U1616 (N_1616,In_91,In_11);
nor U1617 (N_1617,In_385,In_854);
and U1618 (N_1618,In_151,In_675);
nor U1619 (N_1619,In_84,In_883);
or U1620 (N_1620,In_875,In_867);
nor U1621 (N_1621,In_77,In_25);
nor U1622 (N_1622,In_21,In_838);
and U1623 (N_1623,In_171,In_6);
nor U1624 (N_1624,In_911,In_53);
and U1625 (N_1625,In_447,In_709);
nor U1626 (N_1626,In_876,In_225);
and U1627 (N_1627,In_322,In_681);
or U1628 (N_1628,In_143,In_886);
nor U1629 (N_1629,In_310,In_500);
nor U1630 (N_1630,In_606,In_322);
nand U1631 (N_1631,In_172,In_247);
or U1632 (N_1632,In_33,In_536);
and U1633 (N_1633,In_611,In_818);
nand U1634 (N_1634,In_590,In_131);
or U1635 (N_1635,In_872,In_389);
and U1636 (N_1636,In_647,In_443);
nor U1637 (N_1637,In_804,In_824);
or U1638 (N_1638,In_821,In_225);
or U1639 (N_1639,In_620,In_286);
or U1640 (N_1640,In_97,In_364);
nor U1641 (N_1641,In_265,In_555);
and U1642 (N_1642,In_6,In_71);
or U1643 (N_1643,In_369,In_357);
nor U1644 (N_1644,In_397,In_347);
and U1645 (N_1645,In_995,In_104);
nand U1646 (N_1646,In_992,In_779);
nor U1647 (N_1647,In_3,In_864);
and U1648 (N_1648,In_457,In_605);
or U1649 (N_1649,In_497,In_683);
and U1650 (N_1650,In_668,In_157);
nand U1651 (N_1651,In_908,In_377);
nor U1652 (N_1652,In_101,In_605);
xor U1653 (N_1653,In_442,In_173);
and U1654 (N_1654,In_967,In_681);
nor U1655 (N_1655,In_402,In_714);
and U1656 (N_1656,In_207,In_539);
or U1657 (N_1657,In_603,In_882);
or U1658 (N_1658,In_333,In_273);
nand U1659 (N_1659,In_990,In_390);
and U1660 (N_1660,In_795,In_698);
or U1661 (N_1661,In_247,In_965);
and U1662 (N_1662,In_496,In_580);
nor U1663 (N_1663,In_918,In_594);
nand U1664 (N_1664,In_324,In_589);
nand U1665 (N_1665,In_756,In_336);
or U1666 (N_1666,In_657,In_290);
nor U1667 (N_1667,In_452,In_779);
and U1668 (N_1668,In_311,In_816);
xor U1669 (N_1669,In_569,In_146);
nand U1670 (N_1670,In_780,In_374);
nor U1671 (N_1671,In_350,In_767);
and U1672 (N_1672,In_824,In_673);
or U1673 (N_1673,In_209,In_955);
nor U1674 (N_1674,In_151,In_584);
nor U1675 (N_1675,In_39,In_474);
and U1676 (N_1676,In_283,In_583);
nor U1677 (N_1677,In_216,In_880);
or U1678 (N_1678,In_554,In_210);
nor U1679 (N_1679,In_739,In_726);
or U1680 (N_1680,In_840,In_190);
and U1681 (N_1681,In_674,In_277);
or U1682 (N_1682,In_464,In_641);
or U1683 (N_1683,In_880,In_467);
nor U1684 (N_1684,In_510,In_411);
nor U1685 (N_1685,In_56,In_48);
nor U1686 (N_1686,In_431,In_575);
or U1687 (N_1687,In_518,In_706);
nand U1688 (N_1688,In_895,In_597);
or U1689 (N_1689,In_859,In_419);
nor U1690 (N_1690,In_406,In_740);
nand U1691 (N_1691,In_986,In_368);
nand U1692 (N_1692,In_46,In_169);
or U1693 (N_1693,In_519,In_214);
and U1694 (N_1694,In_800,In_164);
and U1695 (N_1695,In_367,In_657);
and U1696 (N_1696,In_484,In_409);
nand U1697 (N_1697,In_125,In_315);
nand U1698 (N_1698,In_730,In_520);
nor U1699 (N_1699,In_891,In_586);
nand U1700 (N_1700,In_357,In_678);
nand U1701 (N_1701,In_730,In_825);
nand U1702 (N_1702,In_169,In_332);
nor U1703 (N_1703,In_272,In_501);
and U1704 (N_1704,In_587,In_153);
nand U1705 (N_1705,In_805,In_676);
or U1706 (N_1706,In_142,In_918);
or U1707 (N_1707,In_691,In_942);
or U1708 (N_1708,In_372,In_91);
or U1709 (N_1709,In_708,In_96);
and U1710 (N_1710,In_608,In_902);
and U1711 (N_1711,In_405,In_345);
nor U1712 (N_1712,In_62,In_330);
nand U1713 (N_1713,In_569,In_44);
xnor U1714 (N_1714,In_448,In_834);
and U1715 (N_1715,In_375,In_148);
nor U1716 (N_1716,In_982,In_93);
and U1717 (N_1717,In_285,In_677);
nand U1718 (N_1718,In_304,In_681);
nor U1719 (N_1719,In_890,In_501);
and U1720 (N_1720,In_148,In_704);
and U1721 (N_1721,In_467,In_23);
nor U1722 (N_1722,In_391,In_626);
and U1723 (N_1723,In_924,In_821);
xor U1724 (N_1724,In_552,In_50);
or U1725 (N_1725,In_246,In_244);
nand U1726 (N_1726,In_983,In_90);
nand U1727 (N_1727,In_404,In_985);
and U1728 (N_1728,In_533,In_718);
nand U1729 (N_1729,In_966,In_113);
or U1730 (N_1730,In_829,In_544);
nand U1731 (N_1731,In_198,In_419);
and U1732 (N_1732,In_387,In_303);
nor U1733 (N_1733,In_832,In_202);
or U1734 (N_1734,In_899,In_408);
nand U1735 (N_1735,In_238,In_709);
nand U1736 (N_1736,In_890,In_496);
nand U1737 (N_1737,In_599,In_638);
or U1738 (N_1738,In_484,In_737);
or U1739 (N_1739,In_178,In_341);
nor U1740 (N_1740,In_70,In_726);
nor U1741 (N_1741,In_955,In_990);
or U1742 (N_1742,In_943,In_315);
nand U1743 (N_1743,In_719,In_243);
or U1744 (N_1744,In_591,In_248);
and U1745 (N_1745,In_440,In_536);
or U1746 (N_1746,In_959,In_705);
nand U1747 (N_1747,In_316,In_108);
or U1748 (N_1748,In_815,In_695);
and U1749 (N_1749,In_608,In_884);
nand U1750 (N_1750,In_115,In_327);
nor U1751 (N_1751,In_873,In_323);
and U1752 (N_1752,In_315,In_293);
nand U1753 (N_1753,In_28,In_734);
and U1754 (N_1754,In_467,In_802);
and U1755 (N_1755,In_952,In_435);
nand U1756 (N_1756,In_506,In_612);
nor U1757 (N_1757,In_193,In_518);
nor U1758 (N_1758,In_519,In_669);
nor U1759 (N_1759,In_346,In_329);
or U1760 (N_1760,In_567,In_86);
nand U1761 (N_1761,In_281,In_153);
and U1762 (N_1762,In_664,In_734);
nand U1763 (N_1763,In_320,In_380);
or U1764 (N_1764,In_426,In_888);
or U1765 (N_1765,In_230,In_221);
or U1766 (N_1766,In_626,In_625);
nor U1767 (N_1767,In_545,In_109);
or U1768 (N_1768,In_523,In_937);
nor U1769 (N_1769,In_371,In_704);
nand U1770 (N_1770,In_65,In_906);
nand U1771 (N_1771,In_528,In_595);
nor U1772 (N_1772,In_489,In_97);
nor U1773 (N_1773,In_482,In_35);
and U1774 (N_1774,In_947,In_346);
nor U1775 (N_1775,In_577,In_602);
and U1776 (N_1776,In_202,In_638);
nor U1777 (N_1777,In_681,In_656);
and U1778 (N_1778,In_654,In_742);
nor U1779 (N_1779,In_288,In_834);
and U1780 (N_1780,In_480,In_179);
nor U1781 (N_1781,In_439,In_336);
nand U1782 (N_1782,In_406,In_35);
nand U1783 (N_1783,In_602,In_428);
and U1784 (N_1784,In_808,In_644);
nor U1785 (N_1785,In_227,In_195);
and U1786 (N_1786,In_523,In_80);
xnor U1787 (N_1787,In_946,In_664);
and U1788 (N_1788,In_161,In_69);
nor U1789 (N_1789,In_838,In_824);
nand U1790 (N_1790,In_717,In_173);
or U1791 (N_1791,In_176,In_448);
or U1792 (N_1792,In_50,In_148);
or U1793 (N_1793,In_574,In_795);
nand U1794 (N_1794,In_862,In_7);
nor U1795 (N_1795,In_884,In_691);
nor U1796 (N_1796,In_430,In_461);
or U1797 (N_1797,In_450,In_382);
nor U1798 (N_1798,In_878,In_397);
and U1799 (N_1799,In_786,In_638);
or U1800 (N_1800,In_588,In_559);
nor U1801 (N_1801,In_255,In_789);
nor U1802 (N_1802,In_604,In_231);
or U1803 (N_1803,In_103,In_445);
nor U1804 (N_1804,In_596,In_285);
nand U1805 (N_1805,In_95,In_64);
nand U1806 (N_1806,In_211,In_750);
or U1807 (N_1807,In_52,In_217);
nand U1808 (N_1808,In_495,In_35);
and U1809 (N_1809,In_191,In_462);
and U1810 (N_1810,In_184,In_871);
nor U1811 (N_1811,In_292,In_826);
or U1812 (N_1812,In_326,In_859);
or U1813 (N_1813,In_675,In_862);
nor U1814 (N_1814,In_431,In_387);
or U1815 (N_1815,In_928,In_332);
and U1816 (N_1816,In_126,In_621);
or U1817 (N_1817,In_394,In_353);
nand U1818 (N_1818,In_822,In_245);
nor U1819 (N_1819,In_65,In_770);
or U1820 (N_1820,In_295,In_565);
or U1821 (N_1821,In_591,In_309);
and U1822 (N_1822,In_148,In_949);
nor U1823 (N_1823,In_347,In_529);
nand U1824 (N_1824,In_184,In_719);
or U1825 (N_1825,In_560,In_941);
or U1826 (N_1826,In_112,In_375);
nand U1827 (N_1827,In_180,In_47);
and U1828 (N_1828,In_950,In_433);
nand U1829 (N_1829,In_789,In_10);
or U1830 (N_1830,In_330,In_123);
and U1831 (N_1831,In_908,In_347);
nand U1832 (N_1832,In_794,In_760);
nor U1833 (N_1833,In_83,In_191);
or U1834 (N_1834,In_421,In_367);
and U1835 (N_1835,In_906,In_97);
and U1836 (N_1836,In_282,In_568);
nand U1837 (N_1837,In_860,In_258);
or U1838 (N_1838,In_624,In_650);
nor U1839 (N_1839,In_295,In_513);
nand U1840 (N_1840,In_541,In_690);
nor U1841 (N_1841,In_824,In_142);
and U1842 (N_1842,In_449,In_552);
and U1843 (N_1843,In_717,In_553);
nor U1844 (N_1844,In_508,In_149);
nor U1845 (N_1845,In_449,In_806);
nor U1846 (N_1846,In_216,In_160);
nand U1847 (N_1847,In_774,In_35);
nand U1848 (N_1848,In_861,In_657);
nand U1849 (N_1849,In_352,In_157);
nor U1850 (N_1850,In_715,In_227);
nand U1851 (N_1851,In_787,In_2);
and U1852 (N_1852,In_589,In_28);
nor U1853 (N_1853,In_103,In_199);
and U1854 (N_1854,In_254,In_484);
nor U1855 (N_1855,In_6,In_294);
and U1856 (N_1856,In_620,In_640);
or U1857 (N_1857,In_532,In_345);
and U1858 (N_1858,In_345,In_194);
or U1859 (N_1859,In_976,In_56);
or U1860 (N_1860,In_564,In_68);
and U1861 (N_1861,In_116,In_896);
and U1862 (N_1862,In_728,In_296);
and U1863 (N_1863,In_877,In_482);
or U1864 (N_1864,In_410,In_794);
or U1865 (N_1865,In_666,In_379);
and U1866 (N_1866,In_534,In_667);
and U1867 (N_1867,In_978,In_853);
or U1868 (N_1868,In_88,In_954);
or U1869 (N_1869,In_643,In_199);
xor U1870 (N_1870,In_244,In_818);
or U1871 (N_1871,In_560,In_12);
or U1872 (N_1872,In_262,In_211);
nand U1873 (N_1873,In_233,In_144);
and U1874 (N_1874,In_635,In_40);
and U1875 (N_1875,In_358,In_321);
nor U1876 (N_1876,In_929,In_145);
or U1877 (N_1877,In_654,In_632);
or U1878 (N_1878,In_256,In_990);
nand U1879 (N_1879,In_381,In_497);
nor U1880 (N_1880,In_594,In_333);
or U1881 (N_1881,In_203,In_583);
nor U1882 (N_1882,In_264,In_11);
nand U1883 (N_1883,In_198,In_457);
nand U1884 (N_1884,In_834,In_66);
and U1885 (N_1885,In_696,In_782);
nor U1886 (N_1886,In_183,In_938);
nand U1887 (N_1887,In_309,In_222);
and U1888 (N_1888,In_861,In_141);
and U1889 (N_1889,In_235,In_109);
nor U1890 (N_1890,In_900,In_740);
or U1891 (N_1891,In_394,In_456);
nor U1892 (N_1892,In_615,In_936);
nor U1893 (N_1893,In_959,In_173);
or U1894 (N_1894,In_920,In_154);
nand U1895 (N_1895,In_786,In_403);
nand U1896 (N_1896,In_20,In_605);
or U1897 (N_1897,In_153,In_370);
nor U1898 (N_1898,In_397,In_825);
nor U1899 (N_1899,In_824,In_698);
nor U1900 (N_1900,In_914,In_217);
nor U1901 (N_1901,In_388,In_887);
nand U1902 (N_1902,In_904,In_530);
nor U1903 (N_1903,In_314,In_567);
nor U1904 (N_1904,In_332,In_459);
and U1905 (N_1905,In_735,In_520);
or U1906 (N_1906,In_498,In_77);
or U1907 (N_1907,In_85,In_159);
or U1908 (N_1908,In_837,In_289);
nor U1909 (N_1909,In_304,In_983);
nor U1910 (N_1910,In_479,In_798);
nor U1911 (N_1911,In_506,In_626);
nand U1912 (N_1912,In_810,In_561);
and U1913 (N_1913,In_624,In_873);
nand U1914 (N_1914,In_454,In_661);
and U1915 (N_1915,In_607,In_929);
or U1916 (N_1916,In_339,In_232);
and U1917 (N_1917,In_176,In_55);
nor U1918 (N_1918,In_191,In_740);
nor U1919 (N_1919,In_474,In_308);
nor U1920 (N_1920,In_188,In_536);
and U1921 (N_1921,In_175,In_958);
or U1922 (N_1922,In_769,In_452);
or U1923 (N_1923,In_555,In_206);
or U1924 (N_1924,In_683,In_85);
nor U1925 (N_1925,In_794,In_776);
xor U1926 (N_1926,In_3,In_247);
nor U1927 (N_1927,In_157,In_58);
and U1928 (N_1928,In_308,In_531);
nor U1929 (N_1929,In_282,In_604);
nand U1930 (N_1930,In_627,In_876);
and U1931 (N_1931,In_205,In_728);
nor U1932 (N_1932,In_640,In_856);
nand U1933 (N_1933,In_323,In_974);
and U1934 (N_1934,In_289,In_254);
nand U1935 (N_1935,In_184,In_110);
and U1936 (N_1936,In_598,In_327);
nand U1937 (N_1937,In_646,In_653);
nand U1938 (N_1938,In_827,In_57);
and U1939 (N_1939,In_42,In_276);
nor U1940 (N_1940,In_496,In_702);
nand U1941 (N_1941,In_769,In_41);
nor U1942 (N_1942,In_215,In_711);
or U1943 (N_1943,In_387,In_614);
and U1944 (N_1944,In_424,In_361);
nor U1945 (N_1945,In_688,In_625);
nand U1946 (N_1946,In_630,In_941);
and U1947 (N_1947,In_970,In_891);
or U1948 (N_1948,In_981,In_367);
nand U1949 (N_1949,In_421,In_571);
nand U1950 (N_1950,In_677,In_648);
nor U1951 (N_1951,In_213,In_694);
and U1952 (N_1952,In_831,In_476);
nand U1953 (N_1953,In_640,In_967);
nand U1954 (N_1954,In_944,In_716);
nor U1955 (N_1955,In_938,In_822);
nor U1956 (N_1956,In_246,In_926);
nand U1957 (N_1957,In_516,In_724);
nor U1958 (N_1958,In_190,In_43);
or U1959 (N_1959,In_181,In_802);
nand U1960 (N_1960,In_168,In_675);
nand U1961 (N_1961,In_102,In_900);
nand U1962 (N_1962,In_522,In_74);
and U1963 (N_1963,In_622,In_427);
or U1964 (N_1964,In_702,In_552);
nand U1965 (N_1965,In_407,In_390);
nand U1966 (N_1966,In_61,In_614);
nor U1967 (N_1967,In_182,In_763);
nor U1968 (N_1968,In_41,In_151);
and U1969 (N_1969,In_543,In_688);
and U1970 (N_1970,In_324,In_443);
nor U1971 (N_1971,In_980,In_469);
xor U1972 (N_1972,In_218,In_338);
and U1973 (N_1973,In_864,In_359);
and U1974 (N_1974,In_945,In_64);
nor U1975 (N_1975,In_544,In_327);
and U1976 (N_1976,In_356,In_629);
and U1977 (N_1977,In_676,In_207);
nor U1978 (N_1978,In_614,In_500);
nand U1979 (N_1979,In_94,In_507);
nor U1980 (N_1980,In_942,In_153);
and U1981 (N_1981,In_245,In_292);
and U1982 (N_1982,In_891,In_787);
or U1983 (N_1983,In_205,In_288);
nor U1984 (N_1984,In_137,In_800);
nor U1985 (N_1985,In_664,In_146);
or U1986 (N_1986,In_255,In_485);
or U1987 (N_1987,In_734,In_598);
and U1988 (N_1988,In_808,In_777);
or U1989 (N_1989,In_417,In_444);
and U1990 (N_1990,In_487,In_697);
or U1991 (N_1991,In_25,In_449);
or U1992 (N_1992,In_208,In_229);
nor U1993 (N_1993,In_559,In_68);
nor U1994 (N_1994,In_446,In_393);
nand U1995 (N_1995,In_809,In_963);
and U1996 (N_1996,In_928,In_87);
nand U1997 (N_1997,In_801,In_928);
nor U1998 (N_1998,In_968,In_6);
and U1999 (N_1999,In_124,In_497);
nor U2000 (N_2000,N_1457,N_1510);
and U2001 (N_2001,N_1057,N_305);
nor U2002 (N_2002,N_34,N_747);
xor U2003 (N_2003,N_734,N_1490);
nor U2004 (N_2004,N_1259,N_392);
or U2005 (N_2005,N_648,N_1115);
nand U2006 (N_2006,N_1901,N_1884);
nor U2007 (N_2007,N_1565,N_1448);
and U2008 (N_2008,N_1232,N_1599);
and U2009 (N_2009,N_168,N_1846);
and U2010 (N_2010,N_1610,N_117);
nand U2011 (N_2011,N_363,N_1217);
or U2012 (N_2012,N_457,N_1325);
nor U2013 (N_2013,N_1416,N_1204);
or U2014 (N_2014,N_315,N_1093);
or U2015 (N_2015,N_207,N_1076);
or U2016 (N_2016,N_812,N_252);
nand U2017 (N_2017,N_1297,N_1552);
nor U2018 (N_2018,N_1776,N_281);
nor U2019 (N_2019,N_380,N_817);
nor U2020 (N_2020,N_947,N_1066);
nand U2021 (N_2021,N_192,N_257);
and U2022 (N_2022,N_1827,N_1538);
or U2023 (N_2023,N_224,N_1332);
and U2024 (N_2024,N_1673,N_1265);
nor U2025 (N_2025,N_543,N_396);
and U2026 (N_2026,N_1581,N_880);
nand U2027 (N_2027,N_1624,N_791);
and U2028 (N_2028,N_631,N_1589);
or U2029 (N_2029,N_1108,N_1878);
or U2030 (N_2030,N_1166,N_1110);
and U2031 (N_2031,N_1869,N_1503);
nand U2032 (N_2032,N_495,N_1413);
or U2033 (N_2033,N_194,N_826);
nand U2034 (N_2034,N_1560,N_567);
and U2035 (N_2035,N_1568,N_1453);
nor U2036 (N_2036,N_1592,N_885);
nor U2037 (N_2037,N_1524,N_438);
nor U2038 (N_2038,N_411,N_1939);
and U2039 (N_2039,N_1251,N_1263);
nand U2040 (N_2040,N_1426,N_1);
nor U2041 (N_2041,N_1993,N_470);
nor U2042 (N_2042,N_1190,N_299);
or U2043 (N_2043,N_309,N_787);
or U2044 (N_2044,N_733,N_1770);
nor U2045 (N_2045,N_659,N_499);
nand U2046 (N_2046,N_882,N_1918);
nor U2047 (N_2047,N_187,N_706);
and U2048 (N_2048,N_9,N_629);
nor U2049 (N_2049,N_1506,N_243);
nand U2050 (N_2050,N_70,N_1912);
nand U2051 (N_2051,N_1656,N_1079);
nand U2052 (N_2052,N_1123,N_1346);
nand U2053 (N_2053,N_242,N_852);
or U2054 (N_2054,N_398,N_1023);
nor U2055 (N_2055,N_1248,N_1586);
or U2056 (N_2056,N_278,N_135);
or U2057 (N_2057,N_133,N_483);
or U2058 (N_2058,N_318,N_1147);
nand U2059 (N_2059,N_1484,N_1629);
nor U2060 (N_2060,N_754,N_1222);
or U2061 (N_2061,N_1087,N_456);
or U2062 (N_2062,N_1400,N_1742);
or U2063 (N_2063,N_1098,N_476);
or U2064 (N_2064,N_131,N_1529);
nor U2065 (N_2065,N_1981,N_48);
or U2066 (N_2066,N_1614,N_1854);
or U2067 (N_2067,N_1406,N_1192);
nor U2068 (N_2068,N_1310,N_1021);
nand U2069 (N_2069,N_1420,N_707);
xnor U2070 (N_2070,N_710,N_1582);
or U2071 (N_2071,N_3,N_1208);
nor U2072 (N_2072,N_855,N_186);
nor U2073 (N_2073,N_1055,N_307);
nor U2074 (N_2074,N_14,N_1155);
and U2075 (N_2075,N_1486,N_12);
and U2076 (N_2076,N_1316,N_1702);
and U2077 (N_2077,N_92,N_1831);
and U2078 (N_2078,N_1006,N_121);
and U2079 (N_2079,N_1301,N_85);
and U2080 (N_2080,N_1188,N_7);
and U2081 (N_2081,N_858,N_1684);
or U2082 (N_2082,N_81,N_237);
or U2083 (N_2083,N_1101,N_175);
and U2084 (N_2084,N_777,N_612);
nor U2085 (N_2085,N_1362,N_1694);
nor U2086 (N_2086,N_27,N_147);
and U2087 (N_2087,N_416,N_1580);
nor U2088 (N_2088,N_1397,N_1893);
or U2089 (N_2089,N_1293,N_794);
and U2090 (N_2090,N_1683,N_1547);
nor U2091 (N_2091,N_1607,N_1233);
nor U2092 (N_2092,N_1498,N_1883);
or U2093 (N_2093,N_216,N_1951);
nor U2094 (N_2094,N_1441,N_189);
and U2095 (N_2095,N_1758,N_414);
nor U2096 (N_2096,N_1862,N_1478);
nor U2097 (N_2097,N_1177,N_870);
nor U2098 (N_2098,N_519,N_1813);
and U2099 (N_2099,N_1680,N_1491);
and U2100 (N_2100,N_291,N_902);
and U2101 (N_2101,N_282,N_690);
nand U2102 (N_2102,N_864,N_1775);
nor U2103 (N_2103,N_399,N_42);
nand U2104 (N_2104,N_424,N_645);
and U2105 (N_2105,N_1083,N_1711);
or U2106 (N_2106,N_539,N_1964);
and U2107 (N_2107,N_1660,N_113);
or U2108 (N_2108,N_1184,N_1823);
or U2109 (N_2109,N_1170,N_1917);
and U2110 (N_2110,N_1008,N_425);
and U2111 (N_2111,N_1324,N_1916);
nand U2112 (N_2112,N_332,N_1932);
and U2113 (N_2113,N_1142,N_1320);
and U2114 (N_2114,N_1289,N_91);
and U2115 (N_2115,N_1877,N_1246);
nand U2116 (N_2116,N_1200,N_481);
and U2117 (N_2117,N_540,N_1096);
nor U2118 (N_2118,N_1176,N_595);
or U2119 (N_2119,N_1421,N_960);
or U2120 (N_2120,N_508,N_621);
and U2121 (N_2121,N_793,N_21);
or U2122 (N_2122,N_1850,N_169);
nand U2123 (N_2123,N_767,N_576);
nor U2124 (N_2124,N_150,N_638);
or U2125 (N_2125,N_790,N_301);
nand U2126 (N_2126,N_1034,N_1214);
and U2127 (N_2127,N_1151,N_1318);
nor U2128 (N_2128,N_1399,N_30);
and U2129 (N_2129,N_836,N_692);
and U2130 (N_2130,N_449,N_1871);
and U2131 (N_2131,N_634,N_401);
nand U2132 (N_2132,N_918,N_494);
or U2133 (N_2133,N_1226,N_592);
and U2134 (N_2134,N_430,N_763);
and U2135 (N_2135,N_890,N_1097);
or U2136 (N_2136,N_1111,N_1579);
nand U2137 (N_2137,N_1438,N_1493);
or U2138 (N_2138,N_1525,N_651);
and U2139 (N_2139,N_343,N_1608);
nand U2140 (N_2140,N_1873,N_542);
nor U2141 (N_2141,N_179,N_1764);
nor U2142 (N_2142,N_1252,N_1187);
nor U2143 (N_2143,N_570,N_927);
and U2144 (N_2144,N_1002,N_323);
or U2145 (N_2145,N_872,N_770);
or U2146 (N_2146,N_1109,N_1569);
nand U2147 (N_2147,N_1256,N_57);
and U2148 (N_2148,N_784,N_349);
nand U2149 (N_2149,N_879,N_1085);
and U2150 (N_2150,N_579,N_1132);
or U2151 (N_2151,N_1695,N_1521);
nand U2152 (N_2152,N_442,N_832);
or U2153 (N_2153,N_376,N_588);
or U2154 (N_2154,N_501,N_503);
or U2155 (N_2155,N_1300,N_827);
and U2156 (N_2156,N_602,N_663);
nand U2157 (N_2157,N_816,N_909);
nand U2158 (N_2158,N_46,N_1311);
nor U2159 (N_2159,N_350,N_1752);
xor U2160 (N_2160,N_156,N_577);
nand U2161 (N_2161,N_964,N_1531);
nand U2162 (N_2162,N_861,N_51);
nand U2163 (N_2163,N_1800,N_1621);
xnor U2164 (N_2164,N_134,N_962);
or U2165 (N_2165,N_1613,N_838);
nand U2166 (N_2166,N_1836,N_163);
or U2167 (N_2167,N_1548,N_279);
or U2168 (N_2168,N_439,N_584);
or U2169 (N_2169,N_1218,N_1969);
nand U2170 (N_2170,N_1042,N_272);
or U2171 (N_2171,N_1726,N_1830);
and U2172 (N_2172,N_1161,N_1329);
and U2173 (N_2173,N_725,N_983);
and U2174 (N_2174,N_1175,N_208);
nand U2175 (N_2175,N_1848,N_1904);
or U2176 (N_2176,N_1632,N_1743);
or U2177 (N_2177,N_1140,N_1210);
or U2178 (N_2178,N_285,N_1975);
and U2179 (N_2179,N_1052,N_1304);
nor U2180 (N_2180,N_1215,N_86);
and U2181 (N_2181,N_1956,N_923);
or U2182 (N_2182,N_1555,N_249);
nor U2183 (N_2183,N_1460,N_1211);
nor U2184 (N_2184,N_1383,N_726);
nor U2185 (N_2185,N_1106,N_1496);
nor U2186 (N_2186,N_1221,N_361);
or U2187 (N_2187,N_344,N_1388);
nand U2188 (N_2188,N_876,N_1386);
nor U2189 (N_2189,N_566,N_844);
nand U2190 (N_2190,N_1982,N_1874);
or U2191 (N_2191,N_1908,N_1045);
and U2192 (N_2192,N_1001,N_937);
and U2193 (N_2193,N_1889,N_1323);
and U2194 (N_2194,N_41,N_1996);
nand U2195 (N_2195,N_158,N_1985);
and U2196 (N_2196,N_1016,N_792);
nand U2197 (N_2197,N_991,N_959);
and U2198 (N_2198,N_25,N_491);
nand U2199 (N_2199,N_296,N_1302);
or U2200 (N_2200,N_996,N_524);
or U2201 (N_2201,N_831,N_765);
or U2202 (N_2202,N_1801,N_119);
nor U2203 (N_2203,N_1707,N_977);
nand U2204 (N_2204,N_796,N_1987);
or U2205 (N_2205,N_1044,N_1870);
nand U2206 (N_2206,N_1699,N_357);
xnor U2207 (N_2207,N_955,N_840);
nor U2208 (N_2208,N_544,N_1428);
and U2209 (N_2209,N_1077,N_1442);
nand U2210 (N_2210,N_1082,N_247);
and U2211 (N_2211,N_18,N_1365);
or U2212 (N_2212,N_1267,N_1239);
or U2213 (N_2213,N_1279,N_590);
nor U2214 (N_2214,N_1454,N_298);
or U2215 (N_2215,N_729,N_1907);
or U2216 (N_2216,N_772,N_1266);
nor U2217 (N_2217,N_1692,N_903);
nor U2218 (N_2218,N_1024,N_1938);
or U2219 (N_2219,N_1007,N_1567);
or U2220 (N_2220,N_1746,N_1745);
nand U2221 (N_2221,N_334,N_297);
or U2222 (N_2222,N_1043,N_1998);
nand U2223 (N_2223,N_409,N_1157);
and U2224 (N_2224,N_968,N_1104);
or U2225 (N_2225,N_10,N_455);
nand U2226 (N_2226,N_1799,N_926);
or U2227 (N_2227,N_1720,N_1025);
and U2228 (N_2228,N_1872,N_397);
or U2229 (N_2229,N_312,N_308);
nand U2230 (N_2230,N_721,N_1857);
nor U2231 (N_2231,N_1644,N_230);
or U2232 (N_2232,N_1462,N_582);
and U2233 (N_2233,N_1906,N_1336);
nor U2234 (N_2234,N_1288,N_1299);
nor U2235 (N_2235,N_412,N_1773);
and U2236 (N_2236,N_1797,N_1852);
and U2237 (N_2237,N_466,N_1920);
and U2238 (N_2238,N_53,N_1231);
or U2239 (N_2239,N_671,N_1131);
nor U2240 (N_2240,N_166,N_417);
and U2241 (N_2241,N_875,N_549);
and U2242 (N_2242,N_1706,N_461);
nand U2243 (N_2243,N_1509,N_884);
nand U2244 (N_2244,N_408,N_120);
or U2245 (N_2245,N_821,N_933);
and U2246 (N_2246,N_698,N_568);
nor U2247 (N_2247,N_1691,N_869);
nand U2248 (N_2248,N_1639,N_714);
nor U2249 (N_2249,N_1662,N_1084);
and U2250 (N_2250,N_1380,N_1769);
and U2251 (N_2251,N_1507,N_1735);
nor U2252 (N_2252,N_1227,N_1359);
nand U2253 (N_2253,N_84,N_126);
nor U2254 (N_2254,N_1787,N_1331);
nor U2255 (N_2255,N_1103,N_165);
nor U2256 (N_2256,N_984,N_1461);
and U2257 (N_2257,N_1130,N_130);
nand U2258 (N_2258,N_1348,N_775);
nand U2259 (N_2259,N_1747,N_673);
nor U2260 (N_2260,N_160,N_1991);
and U2261 (N_2261,N_1881,N_1716);
nand U2262 (N_2262,N_33,N_686);
and U2263 (N_2263,N_586,N_1526);
or U2264 (N_2264,N_443,N_1688);
nand U2265 (N_2265,N_190,N_1844);
and U2266 (N_2266,N_697,N_1820);
or U2267 (N_2267,N_1867,N_1689);
nand U2268 (N_2268,N_273,N_1499);
nor U2269 (N_2269,N_1180,N_1622);
and U2270 (N_2270,N_1995,N_1431);
and U2271 (N_2271,N_1159,N_541);
and U2272 (N_2272,N_1790,N_972);
nand U2273 (N_2273,N_650,N_1005);
nor U2274 (N_2274,N_201,N_195);
or U2275 (N_2275,N_713,N_109);
and U2276 (N_2276,N_637,N_1968);
or U2277 (N_2277,N_1739,N_153);
or U2278 (N_2278,N_1378,N_521);
nor U2279 (N_2279,N_1564,N_1763);
nand U2280 (N_2280,N_124,N_319);
and U2281 (N_2281,N_1627,N_1254);
nor U2282 (N_2282,N_1062,N_1863);
nor U2283 (N_2283,N_758,N_1150);
or U2284 (N_2284,N_75,N_802);
nor U2285 (N_2285,N_625,N_1887);
nor U2286 (N_2286,N_205,N_322);
and U2287 (N_2287,N_658,N_1843);
nand U2288 (N_2288,N_1946,N_1886);
nor U2289 (N_2289,N_755,N_665);
xor U2290 (N_2290,N_1812,N_1407);
and U2291 (N_2291,N_1468,N_448);
and U2292 (N_2292,N_1027,N_1139);
and U2293 (N_2293,N_504,N_59);
and U2294 (N_2294,N_1339,N_222);
or U2295 (N_2295,N_1961,N_1544);
nand U2296 (N_2296,N_1149,N_788);
or U2297 (N_2297,N_1069,N_354);
or U2298 (N_2298,N_1980,N_1258);
and U2299 (N_2299,N_240,N_83);
or U2300 (N_2300,N_306,N_182);
or U2301 (N_2301,N_771,N_709);
nand U2302 (N_2302,N_250,N_1053);
or U2303 (N_2303,N_1741,N_63);
nand U2304 (N_2304,N_258,N_1269);
nor U2305 (N_2305,N_871,N_768);
nand U2306 (N_2306,N_351,N_1875);
xnor U2307 (N_2307,N_320,N_1591);
nand U2308 (N_2308,N_825,N_532);
nor U2309 (N_2309,N_857,N_472);
nand U2310 (N_2310,N_1390,N_623);
nand U2311 (N_2311,N_437,N_1120);
and U2312 (N_2312,N_685,N_1409);
nand U2313 (N_2313,N_1663,N_1402);
nand U2314 (N_2314,N_58,N_1168);
nor U2315 (N_2315,N_529,N_159);
nand U2316 (N_2316,N_730,N_1755);
or U2317 (N_2317,N_1196,N_467);
nor U2318 (N_2318,N_911,N_464);
xnor U2319 (N_2319,N_1395,N_778);
nor U2320 (N_2320,N_1137,N_701);
nand U2321 (N_2321,N_1974,N_525);
or U2322 (N_2322,N_1911,N_1306);
and U2323 (N_2323,N_256,N_894);
or U2324 (N_2324,N_564,N_641);
nand U2325 (N_2325,N_61,N_391);
and U2326 (N_2326,N_445,N_1281);
or U2327 (N_2327,N_1921,N_1642);
or U2328 (N_2328,N_1670,N_652);
and U2329 (N_2329,N_386,N_1179);
and U2330 (N_2330,N_1636,N_38);
or U2331 (N_2331,N_516,N_125);
nand U2332 (N_2332,N_141,N_118);
nand U2333 (N_2333,N_1225,N_1379);
or U2334 (N_2334,N_295,N_1253);
or U2335 (N_2335,N_337,N_786);
nand U2336 (N_2336,N_845,N_333);
nand U2337 (N_2337,N_795,N_1681);
xnor U2338 (N_2338,N_1282,N_1377);
nor U2339 (N_2339,N_173,N_1558);
or U2340 (N_2340,N_490,N_1437);
and U2341 (N_2341,N_624,N_547);
xor U2342 (N_2342,N_1469,N_565);
and U2343 (N_2343,N_992,N_269);
or U2344 (N_2344,N_1909,N_1709);
nand U2345 (N_2345,N_1892,N_446);
nor U2346 (N_2346,N_407,N_687);
and U2347 (N_2347,N_1577,N_776);
or U2348 (N_2348,N_822,N_610);
and U2349 (N_2349,N_1896,N_948);
nor U2350 (N_2350,N_1730,N_723);
and U2351 (N_2351,N_1305,N_1923);
or U2352 (N_2352,N_1516,N_387);
nor U2353 (N_2353,N_666,N_915);
and U2354 (N_2354,N_1136,N_860);
or U2355 (N_2355,N_1434,N_807);
and U2356 (N_2356,N_1038,N_679);
and U2357 (N_2357,N_904,N_1385);
nor U2358 (N_2358,N_609,N_78);
and U2359 (N_2359,N_711,N_198);
xor U2360 (N_2360,N_1994,N_980);
nor U2361 (N_2361,N_1209,N_1479);
or U2362 (N_2362,N_824,N_1537);
and U2363 (N_2363,N_413,N_1924);
nor U2364 (N_2364,N_988,N_1286);
nand U2365 (N_2365,N_183,N_227);
nor U2366 (N_2366,N_669,N_1174);
nor U2367 (N_2367,N_47,N_535);
and U2368 (N_2368,N_1374,N_626);
nor U2369 (N_2369,N_1126,N_1578);
nand U2370 (N_2370,N_1962,N_1808);
and U2371 (N_2371,N_670,N_560);
nand U2372 (N_2372,N_1721,N_608);
or U2373 (N_2373,N_967,N_917);
nand U2374 (N_2374,N_1633,N_1733);
and U2375 (N_2375,N_1795,N_152);
nor U2376 (N_2376,N_1124,N_1321);
and U2377 (N_2377,N_1056,N_1668);
nor U2378 (N_2378,N_1774,N_1542);
nor U2379 (N_2379,N_1655,N_480);
nand U2380 (N_2380,N_447,N_1957);
nand U2381 (N_2381,N_1207,N_731);
nand U2382 (N_2382,N_874,N_559);
and U2383 (N_2383,N_1925,N_897);
nand U2384 (N_2384,N_290,N_1063);
nand U2385 (N_2385,N_1765,N_799);
nor U2386 (N_2386,N_454,N_810);
and U2387 (N_2387,N_1158,N_1809);
or U2388 (N_2388,N_1172,N_963);
xor U2389 (N_2389,N_1556,N_773);
nand U2390 (N_2390,N_217,N_1117);
and U2391 (N_2391,N_520,N_883);
or U2392 (N_2392,N_803,N_762);
and U2393 (N_2393,N_1890,N_288);
nor U2394 (N_2394,N_1811,N_1929);
nand U2395 (N_2395,N_639,N_1815);
nor U2396 (N_2396,N_1520,N_428);
xor U2397 (N_2397,N_1658,N_1144);
nand U2398 (N_2398,N_1532,N_1292);
nand U2399 (N_2399,N_1659,N_509);
nand U2400 (N_2400,N_1017,N_1156);
xor U2401 (N_2401,N_1476,N_1864);
nand U2402 (N_2402,N_97,N_505);
nor U2403 (N_2403,N_1999,N_1433);
nand U2404 (N_2404,N_944,N_847);
or U2405 (N_2405,N_1145,N_1554);
nand U2406 (N_2406,N_1349,N_1724);
or U2407 (N_2407,N_779,N_1489);
nand U2408 (N_2408,N_1430,N_677);
nor U2409 (N_2409,N_1230,N_1540);
nor U2410 (N_2410,N_1127,N_1612);
and U2411 (N_2411,N_1944,N_1094);
nor U2412 (N_2412,N_170,N_1429);
nand U2413 (N_2413,N_1018,N_1549);
and U2414 (N_2414,N_1467,N_502);
nand U2415 (N_2415,N_1687,N_451);
and U2416 (N_2416,N_325,N_1347);
or U2417 (N_2417,N_1370,N_1832);
nor U2418 (N_2418,N_575,N_1181);
and U2419 (N_2419,N_1766,N_901);
nor U2420 (N_2420,N_1086,N_475);
and U2421 (N_2421,N_1250,N_1640);
and U2422 (N_2422,N_218,N_1480);
or U2423 (N_2423,N_932,N_410);
or U2424 (N_2424,N_1118,N_694);
nand U2425 (N_2425,N_1527,N_229);
nor U2426 (N_2426,N_717,N_700);
or U2427 (N_2427,N_533,N_1700);
or U2428 (N_2428,N_618,N_1167);
and U2429 (N_2429,N_1242,N_1272);
nand U2430 (N_2430,N_1833,N_756);
and U2431 (N_2431,N_1060,N_1223);
nand U2432 (N_2432,N_693,N_164);
nor U2433 (N_2433,N_60,N_931);
nor U2434 (N_2434,N_1326,N_1114);
and U2435 (N_2435,N_1444,N_675);
and U2436 (N_2436,N_934,N_1501);
and U2437 (N_2437,N_489,N_674);
nor U2438 (N_2438,N_1340,N_1802);
and U2439 (N_2439,N_613,N_953);
or U2440 (N_2440,N_142,N_819);
nor U2441 (N_2441,N_1708,N_154);
or U2442 (N_2442,N_1371,N_1492);
nand U2443 (N_2443,N_1842,N_1665);
nor U2444 (N_2444,N_206,N_1403);
nor U2445 (N_2445,N_11,N_1536);
nor U2446 (N_2446,N_1219,N_203);
and U2447 (N_2447,N_1652,N_925);
nor U2448 (N_2448,N_1583,N_1337);
and U2449 (N_2449,N_1585,N_1031);
nor U2450 (N_2450,N_93,N_716);
and U2451 (N_2451,N_881,N_1678);
or U2452 (N_2452,N_1853,N_534);
nor U2453 (N_2453,N_268,N_287);
or U2454 (N_2454,N_157,N_1308);
nor U2455 (N_2455,N_1675,N_916);
or U2456 (N_2456,N_1605,N_1634);
and U2457 (N_2457,N_761,N_493);
and U2458 (N_2458,N_1679,N_174);
xor U2459 (N_2459,N_1081,N_1930);
xor U2460 (N_2460,N_1330,N_1910);
and U2461 (N_2461,N_1826,N_672);
nor U2462 (N_2462,N_1731,N_24);
nor U2463 (N_2463,N_751,N_303);
and U2464 (N_2464,N_1012,N_688);
or U2465 (N_2465,N_418,N_104);
nor U2466 (N_2466,N_906,N_110);
nand U2467 (N_2467,N_328,N_359);
or U2468 (N_2468,N_748,N_1860);
and U2469 (N_2469,N_1705,N_251);
xnor U2470 (N_2470,N_536,N_1539);
or U2471 (N_2471,N_867,N_851);
nor U2472 (N_2472,N_221,N_1352);
nand U2473 (N_2473,N_1905,N_1417);
nand U2474 (N_2474,N_1112,N_1105);
nor U2475 (N_2475,N_558,N_712);
nand U2476 (N_2476,N_1414,N_1973);
nand U2477 (N_2477,N_813,N_69);
nand U2478 (N_2478,N_805,N_512);
or U2479 (N_2479,N_1997,N_531);
and U2480 (N_2480,N_1472,N_1819);
nor U2481 (N_2481,N_45,N_782);
nand U2482 (N_2482,N_554,N_1979);
or U2483 (N_2483,N_603,N_1628);
and U2484 (N_2484,N_1317,N_488);
nand U2485 (N_2485,N_1903,N_339);
or U2486 (N_2486,N_1926,N_384);
nand U2487 (N_2487,N_127,N_1839);
and U2488 (N_2488,N_1792,N_809);
or U2489 (N_2489,N_1354,N_76);
nand U2490 (N_2490,N_193,N_849);
nand U2491 (N_2491,N_1241,N_848);
and U2492 (N_2492,N_64,N_1671);
and U2493 (N_2493,N_732,N_1319);
nand U2494 (N_2494,N_54,N_1424);
and U2495 (N_2495,N_441,N_589);
nor U2496 (N_2496,N_1654,N_1779);
nand U2497 (N_2497,N_66,N_115);
nand U2498 (N_2498,N_274,N_1477);
or U2499 (N_2499,N_997,N_1757);
and U2500 (N_2500,N_681,N_1646);
and U2501 (N_2501,N_420,N_601);
and U2502 (N_2502,N_1781,N_199);
nor U2503 (N_2503,N_978,N_1296);
nand U2504 (N_2504,N_830,N_20);
or U2505 (N_2505,N_974,N_950);
nor U2506 (N_2506,N_327,N_171);
nor U2507 (N_2507,N_1271,N_653);
nor U2508 (N_2508,N_971,N_530);
nand U2509 (N_2509,N_275,N_789);
or U2510 (N_2510,N_460,N_1427);
or U2511 (N_2511,N_1235,N_1364);
and U2512 (N_2512,N_144,N_105);
nand U2513 (N_2513,N_528,N_936);
nand U2514 (N_2514,N_1197,N_1888);
and U2515 (N_2515,N_140,N_908);
and U2516 (N_2516,N_1091,N_738);
and U2517 (N_2517,N_68,N_1748);
and U2518 (N_2518,N_661,N_1977);
and U2519 (N_2519,N_1356,N_667);
and U2520 (N_2520,N_1229,N_620);
nor U2521 (N_2521,N_887,N_545);
and U2522 (N_2522,N_1497,N_178);
and U2523 (N_2523,N_185,N_1343);
nor U2524 (N_2524,N_998,N_400);
or U2525 (N_2525,N_1382,N_468);
and U2526 (N_2526,N_77,N_373);
and U2527 (N_2527,N_1682,N_814);
nor U2528 (N_2528,N_347,N_1361);
nor U2529 (N_2529,N_1000,N_1717);
nand U2530 (N_2530,N_1309,N_31);
or U2531 (N_2531,N_231,N_1948);
or U2532 (N_2532,N_1919,N_1028);
and U2533 (N_2533,N_1153,N_28);
nand U2534 (N_2534,N_854,N_728);
and U2535 (N_2535,N_957,N_500);
and U2536 (N_2536,N_6,N_742);
and U2537 (N_2537,N_1804,N_1715);
nand U2538 (N_2538,N_346,N_1794);
nor U2539 (N_2539,N_599,N_1391);
nor U2540 (N_2540,N_1935,N_1270);
nand U2541 (N_2541,N_498,N_1523);
and U2542 (N_2542,N_1791,N_1070);
and U2543 (N_2543,N_1471,N_999);
nor U2544 (N_2544,N_823,N_1059);
nand U2545 (N_2545,N_1135,N_146);
and U2546 (N_2546,N_750,N_394);
nor U2547 (N_2547,N_116,N_1143);
and U2548 (N_2548,N_1749,N_946);
and U2549 (N_2549,N_850,N_1154);
nand U2550 (N_2550,N_804,N_1805);
nor U2551 (N_2551,N_1519,N_56);
nand U2552 (N_2552,N_302,N_1412);
and U2553 (N_2553,N_1089,N_829);
or U2554 (N_2554,N_1713,N_703);
nor U2555 (N_2555,N_181,N_655);
nor U2556 (N_2556,N_292,N_924);
nand U2557 (N_2557,N_606,N_1753);
or U2558 (N_2558,N_783,N_1494);
and U2559 (N_2559,N_62,N_103);
or U2560 (N_2560,N_1897,N_100);
or U2561 (N_2561,N_197,N_188);
or U2562 (N_2562,N_979,N_640);
nand U2563 (N_2563,N_583,N_73);
and U2564 (N_2564,N_691,N_1806);
or U2565 (N_2565,N_4,N_71);
or U2566 (N_2566,N_1914,N_1759);
or U2567 (N_2567,N_1729,N_89);
nand U2568 (N_2568,N_1314,N_1619);
or U2569 (N_2569,N_1162,N_1095);
nor U2570 (N_2570,N_96,N_1037);
nor U2571 (N_2571,N_1933,N_1936);
nand U2572 (N_2572,N_1334,N_383);
and U2573 (N_2573,N_1559,N_1446);
or U2574 (N_2574,N_106,N_212);
nand U2575 (N_2575,N_149,N_145);
nand U2576 (N_2576,N_1363,N_16);
or U2577 (N_2577,N_317,N_1100);
nor U2578 (N_2578,N_1845,N_1945);
or U2579 (N_2579,N_1814,N_764);
nor U2580 (N_2580,N_220,N_1573);
or U2581 (N_2581,N_1988,N_1788);
nand U2582 (N_2582,N_1954,N_662);
nor U2583 (N_2583,N_1756,N_405);
nand U2584 (N_2584,N_572,N_1931);
xnor U2585 (N_2585,N_1934,N_1697);
nor U2586 (N_2586,N_1061,N_1672);
nor U2587 (N_2587,N_1366,N_654);
nand U2588 (N_2588,N_1401,N_1740);
or U2589 (N_2589,N_1966,N_615);
and U2590 (N_2590,N_1880,N_371);
or U2591 (N_2591,N_55,N_151);
nor U2592 (N_2592,N_1847,N_719);
nor U2593 (N_2593,N_737,N_1772);
nand U2594 (N_2594,N_553,N_1732);
and U2595 (N_2595,N_684,N_482);
nand U2596 (N_2596,N_1835,N_1950);
or U2597 (N_2597,N_617,N_956);
or U2598 (N_2598,N_1648,N_368);
and U2599 (N_2599,N_527,N_1313);
and U2600 (N_2600,N_1022,N_1015);
or U2601 (N_2601,N_1030,N_1032);
nand U2602 (N_2602,N_1796,N_1899);
or U2603 (N_2603,N_390,N_797);
or U2604 (N_2604,N_806,N_1182);
or U2605 (N_2605,N_555,N_1450);
and U2606 (N_2606,N_8,N_1793);
nand U2607 (N_2607,N_1009,N_1952);
nor U2608 (N_2608,N_1965,N_421);
or U2609 (N_2609,N_444,N_244);
nor U2610 (N_2610,N_263,N_1635);
and U2611 (N_2611,N_236,N_1690);
nor U2612 (N_2612,N_1571,N_569);
nand U2613 (N_2613,N_895,N_1262);
or U2614 (N_2614,N_1078,N_239);
or U2615 (N_2615,N_961,N_161);
or U2616 (N_2616,N_1268,N_1593);
and U2617 (N_2617,N_966,N_226);
and U2618 (N_2618,N_1609,N_235);
or U2619 (N_2619,N_246,N_1572);
nor U2620 (N_2620,N_1643,N_1840);
or U2621 (N_2621,N_372,N_1322);
nor U2622 (N_2622,N_74,N_1898);
and U2623 (N_2623,N_1465,N_1206);
nand U2624 (N_2624,N_604,N_981);
or U2625 (N_2625,N_492,N_65);
nand U2626 (N_2626,N_1338,N_1389);
nor U2627 (N_2627,N_1976,N_260);
nor U2628 (N_2628,N_1576,N_1128);
or U2629 (N_2629,N_935,N_1458);
and U2630 (N_2630,N_1515,N_184);
nor U2631 (N_2631,N_1102,N_1891);
and U2632 (N_2632,N_316,N_1119);
nor U2633 (N_2633,N_422,N_985);
nand U2634 (N_2634,N_989,N_1373);
nor U2635 (N_2635,N_952,N_1657);
nor U2636 (N_2636,N_1148,N_664);
and U2637 (N_2637,N_1602,N_352);
nand U2638 (N_2638,N_1512,N_1195);
nor U2639 (N_2639,N_513,N_1727);
or U2640 (N_2640,N_1483,N_598);
nor U2641 (N_2641,N_1594,N_1029);
nand U2642 (N_2642,N_1287,N_459);
or U2643 (N_2643,N_1274,N_1895);
and U2644 (N_2644,N_431,N_1327);
nand U2645 (N_2645,N_1620,N_646);
nand U2646 (N_2646,N_1333,N_360);
nor U2647 (N_2647,N_1452,N_1129);
nand U2648 (N_2648,N_261,N_1367);
nand U2649 (N_2649,N_1355,N_264);
or U2650 (N_2650,N_1734,N_474);
and U2651 (N_2651,N_892,N_1398);
nor U2652 (N_2652,N_329,N_23);
and U2653 (N_2653,N_1464,N_1394);
or U2654 (N_2654,N_365,N_940);
nand U2655 (N_2655,N_402,N_735);
nand U2656 (N_2656,N_311,N_1518);
nand U2657 (N_2657,N_1990,N_1344);
nand U2658 (N_2658,N_95,N_1821);
and U2659 (N_2659,N_1653,N_497);
nor U2660 (N_2660,N_757,N_1942);
or U2661 (N_2661,N_1470,N_853);
nand U2662 (N_2662,N_280,N_1216);
and U2663 (N_2663,N_1943,N_67);
and U2664 (N_2664,N_1152,N_1121);
and U2665 (N_2665,N_1199,N_943);
nor U2666 (N_2666,N_1169,N_1003);
and U2667 (N_2667,N_35,N_699);
nand U2668 (N_2668,N_1125,N_1513);
nor U2669 (N_2669,N_1807,N_1185);
and U2670 (N_2670,N_1744,N_868);
or U2671 (N_2671,N_196,N_1626);
nand U2672 (N_2672,N_313,N_580);
nand U2673 (N_2673,N_1396,N_238);
nand U2674 (N_2674,N_563,N_50);
or U2675 (N_2675,N_453,N_1178);
nand U2676 (N_2676,N_389,N_1782);
or U2677 (N_2677,N_1368,N_215);
nor U2678 (N_2678,N_642,N_1075);
or U2679 (N_2679,N_1351,N_1777);
or U2680 (N_2680,N_1505,N_1958);
nor U2681 (N_2681,N_26,N_435);
nor U2682 (N_2682,N_507,N_87);
nor U2683 (N_2683,N_1261,N_1970);
nand U2684 (N_2684,N_607,N_1280);
and U2685 (N_2685,N_1183,N_1487);
and U2686 (N_2686,N_326,N_616);
or U2687 (N_2687,N_1290,N_1381);
nand U2688 (N_2688,N_1528,N_614);
nand U2689 (N_2689,N_1463,N_1859);
nor U2690 (N_2690,N_1666,N_913);
nor U2691 (N_2691,N_1283,N_1439);
or U2692 (N_2692,N_740,N_914);
and U2693 (N_2693,N_1133,N_1530);
and U2694 (N_2694,N_1885,N_1611);
or U2695 (N_2695,N_1701,N_1134);
and U2696 (N_2696,N_1198,N_1041);
nand U2697 (N_2697,N_370,N_1392);
or U2698 (N_2698,N_111,N_353);
nor U2699 (N_2699,N_877,N_878);
nor U2700 (N_2700,N_689,N_605);
nor U2701 (N_2701,N_1737,N_801);
xnor U2702 (N_2702,N_1960,N_1545);
and U2703 (N_2703,N_627,N_1312);
and U2704 (N_2704,N_600,N_265);
or U2705 (N_2705,N_1050,N_37);
nand U2706 (N_2706,N_766,N_1203);
nor U2707 (N_2707,N_1255,N_382);
nand U2708 (N_2708,N_211,N_452);
nor U2709 (N_2709,N_656,N_1989);
nand U2710 (N_2710,N_341,N_213);
nand U2711 (N_2711,N_176,N_286);
nand U2712 (N_2712,N_835,N_1436);
nand U2713 (N_2713,N_1408,N_1677);
nand U2714 (N_2714,N_1224,N_910);
or U2715 (N_2715,N_886,N_433);
nor U2716 (N_2716,N_1963,N_485);
nand U2717 (N_2717,N_587,N_1723);
nand U2718 (N_2718,N_866,N_1562);
or U2719 (N_2719,N_107,N_1984);
nor U2720 (N_2720,N_1650,N_1829);
nand U2721 (N_2721,N_1243,N_993);
nand U2722 (N_2722,N_907,N_374);
nor U2723 (N_2723,N_1767,N_1033);
and U2724 (N_2724,N_43,N_1570);
and U2725 (N_2725,N_1551,N_1882);
nand U2726 (N_2726,N_128,N_1455);
nor U2727 (N_2727,N_1074,N_284);
nand U2728 (N_2728,N_1419,N_636);
and U2729 (N_2729,N_1474,N_484);
or U2730 (N_2730,N_774,N_1482);
or U2731 (N_2731,N_930,N_1597);
or U2732 (N_2732,N_1341,N_1618);
nand U2733 (N_2733,N_1202,N_88);
or U2734 (N_2734,N_760,N_833);
and U2735 (N_2735,N_1107,N_1816);
or U2736 (N_2736,N_1298,N_702);
or U2737 (N_2737,N_1947,N_1818);
nor U2738 (N_2738,N_1164,N_458);
and U2739 (N_2739,N_994,N_596);
and U2740 (N_2740,N_348,N_377);
and U2741 (N_2741,N_293,N_632);
or U2742 (N_2742,N_1789,N_1278);
nor U2743 (N_2743,N_214,N_808);
and U2744 (N_2744,N_1116,N_715);
nor U2745 (N_2745,N_155,N_1574);
nand U2746 (N_2746,N_949,N_1247);
nand U2747 (N_2747,N_1387,N_1238);
or U2748 (N_2748,N_1785,N_1553);
nor U2749 (N_2749,N_367,N_1533);
or U2750 (N_2750,N_1588,N_611);
nor U2751 (N_2751,N_1550,N_1937);
nor U2752 (N_2752,N_294,N_1803);
nand U2753 (N_2753,N_769,N_556);
and U2754 (N_2754,N_633,N_276);
nor U2755 (N_2755,N_1879,N_1955);
and U2756 (N_2756,N_310,N_815);
or U2757 (N_2757,N_1141,N_1584);
and U2758 (N_2758,N_1783,N_94);
or U2759 (N_2759,N_1761,N_1014);
and U2760 (N_2760,N_635,N_1485);
and U2761 (N_2761,N_143,N_1445);
or U2762 (N_2762,N_1466,N_538);
or U2763 (N_2763,N_1189,N_1587);
nand U2764 (N_2764,N_358,N_496);
nor U2765 (N_2765,N_888,N_5);
nor U2766 (N_2766,N_958,N_1786);
and U2767 (N_2767,N_345,N_1273);
or U2768 (N_2768,N_139,N_1495);
nor U2769 (N_2769,N_643,N_225);
nand U2770 (N_2770,N_746,N_210);
and U2771 (N_2771,N_122,N_1704);
nand U2772 (N_2772,N_17,N_463);
nor U2773 (N_2773,N_1201,N_13);
or U2774 (N_2774,N_136,N_1099);
and U2775 (N_2775,N_342,N_375);
nor U2776 (N_2776,N_1649,N_1623);
and U2777 (N_2777,N_1967,N_486);
and U2778 (N_2778,N_331,N_1696);
nor U2779 (N_2779,N_842,N_362);
nand U2780 (N_2780,N_1601,N_330);
nand U2781 (N_2781,N_233,N_1257);
and U2782 (N_2782,N_1146,N_1500);
nand U2783 (N_2783,N_517,N_1068);
nand U2784 (N_2784,N_515,N_1855);
or U2785 (N_2785,N_395,N_1067);
nand U2786 (N_2786,N_912,N_929);
or U2787 (N_2787,N_1335,N_1345);
nor U2788 (N_2788,N_551,N_1674);
or U2789 (N_2789,N_270,N_1443);
or U2790 (N_2790,N_1511,N_619);
nand U2791 (N_2791,N_941,N_378);
or U2792 (N_2792,N_1113,N_552);
nor U2793 (N_2793,N_510,N_423);
or U2794 (N_2794,N_432,N_80);
and U2795 (N_2795,N_969,N_1165);
and U2796 (N_2796,N_818,N_340);
nor U2797 (N_2797,N_1504,N_593);
nand U2798 (N_2798,N_267,N_259);
and U2799 (N_2799,N_19,N_1598);
nand U2800 (N_2800,N_102,N_743);
and U2801 (N_2801,N_856,N_1534);
nand U2802 (N_2802,N_578,N_1817);
and U2803 (N_2803,N_820,N_1736);
or U2804 (N_2804,N_982,N_112);
and U2805 (N_2805,N_537,N_1828);
and U2806 (N_2806,N_1291,N_1928);
and U2807 (N_2807,N_1048,N_40);
or U2808 (N_2808,N_1425,N_523);
and U2809 (N_2809,N_123,N_1762);
xnor U2810 (N_2810,N_2,N_557);
or U2811 (N_2811,N_1810,N_1771);
nand U2812 (N_2812,N_1861,N_1194);
and U2813 (N_2813,N_506,N_1393);
nand U2814 (N_2814,N_1350,N_1600);
nand U2815 (N_2815,N_1244,N_162);
and U2816 (N_2816,N_1719,N_1851);
or U2817 (N_2817,N_1277,N_1435);
nor U2818 (N_2818,N_628,N_1240);
nand U2819 (N_2819,N_1404,N_1236);
xnor U2820 (N_2820,N_1838,N_253);
nand U2821 (N_2821,N_1940,N_36);
nand U2822 (N_2822,N_1557,N_1010);
and U2823 (N_2823,N_304,N_1451);
nor U2824 (N_2824,N_1971,N_1186);
nor U2825 (N_2825,N_1054,N_1051);
nor U2826 (N_2826,N_1013,N_336);
and U2827 (N_2827,N_942,N_893);
nand U2828 (N_2828,N_1561,N_976);
and U2829 (N_2829,N_546,N_951);
and U2830 (N_2830,N_597,N_1798);
or U2831 (N_2831,N_1615,N_973);
or U2832 (N_2832,N_741,N_1423);
and U2833 (N_2833,N_1972,N_366);
nor U2834 (N_2834,N_1384,N_138);
nand U2835 (N_2835,N_905,N_862);
and U2836 (N_2836,N_415,N_99);
nand U2837 (N_2837,N_1625,N_1508);
and U2838 (N_2838,N_49,N_1171);
nand U2839 (N_2839,N_680,N_1725);
and U2840 (N_2840,N_1865,N_1191);
nor U2841 (N_2841,N_708,N_647);
nand U2842 (N_2842,N_465,N_1522);
nor U2843 (N_2843,N_1080,N_1058);
or U2844 (N_2844,N_1514,N_1703);
nand U2845 (N_2845,N_271,N_1986);
and U2846 (N_2846,N_891,N_355);
or U2847 (N_2847,N_1375,N_574);
and U2848 (N_2848,N_381,N_1047);
nand U2849 (N_2849,N_1049,N_585);
nor U2850 (N_2850,N_683,N_1019);
and U2851 (N_2851,N_427,N_678);
and U2852 (N_2852,N_1447,N_450);
or U2853 (N_2853,N_1606,N_101);
nand U2854 (N_2854,N_1303,N_736);
nor U2855 (N_2855,N_1693,N_800);
nor U2856 (N_2856,N_954,N_369);
nor U2857 (N_2857,N_1011,N_753);
nand U2858 (N_2858,N_865,N_1638);
and U2859 (N_2859,N_1641,N_0);
or U2860 (N_2860,N_29,N_338);
or U2861 (N_2861,N_1750,N_314);
xnor U2862 (N_2862,N_1473,N_1315);
nor U2863 (N_2863,N_1590,N_254);
and U2864 (N_2864,N_965,N_1566);
nor U2865 (N_2865,N_473,N_1422);
and U2866 (N_2866,N_1849,N_571);
nor U2867 (N_2867,N_1418,N_573);
nor U2868 (N_2868,N_970,N_1822);
or U2869 (N_2869,N_899,N_1754);
nand U2870 (N_2870,N_834,N_462);
nand U2871 (N_2871,N_630,N_1372);
and U2872 (N_2872,N_1825,N_1415);
nor U2873 (N_2873,N_1228,N_223);
nand U2874 (N_2874,N_749,N_1275);
nor U2875 (N_2875,N_403,N_148);
nor U2876 (N_2876,N_739,N_1205);
and U2877 (N_2877,N_828,N_1212);
or U2878 (N_2878,N_1264,N_986);
xnor U2879 (N_2879,N_204,N_1004);
and U2880 (N_2880,N_469,N_1978);
nand U2881 (N_2881,N_1405,N_1738);
or U2882 (N_2882,N_1603,N_718);
nand U2883 (N_2883,N_262,N_919);
or U2884 (N_2884,N_724,N_1073);
and U2885 (N_2885,N_704,N_1284);
nor U2886 (N_2886,N_1071,N_1090);
and U2887 (N_2887,N_419,N_1122);
nor U2888 (N_2888,N_324,N_990);
and U2889 (N_2889,N_478,N_429);
nor U2890 (N_2890,N_1630,N_406);
or U2891 (N_2891,N_1837,N_1360);
or U2892 (N_2892,N_1369,N_1712);
nor U2893 (N_2893,N_1722,N_745);
nor U2894 (N_2894,N_644,N_232);
nor U2895 (N_2895,N_1502,N_938);
or U2896 (N_2896,N_1616,N_900);
nor U2897 (N_2897,N_177,N_39);
nand U2898 (N_2898,N_859,N_1440);
nand U2899 (N_2899,N_898,N_1535);
or U2900 (N_2900,N_98,N_1285);
xnor U2901 (N_2901,N_1834,N_1449);
nand U2902 (N_2902,N_1307,N_785);
nand U2903 (N_2903,N_248,N_1481);
and U2904 (N_2904,N_1245,N_1546);
or U2905 (N_2905,N_1651,N_780);
and U2906 (N_2906,N_920,N_32);
nand U2907 (N_2907,N_837,N_811);
or U2908 (N_2908,N_1714,N_622);
or U2909 (N_2909,N_129,N_550);
and U2910 (N_2910,N_1876,N_720);
nor U2911 (N_2911,N_1676,N_1751);
and U2912 (N_2912,N_1949,N_479);
nor U2913 (N_2913,N_1459,N_526);
or U2914 (N_2914,N_436,N_385);
nor U2915 (N_2915,N_660,N_1065);
or U2916 (N_2916,N_727,N_300);
nand U2917 (N_2917,N_90,N_277);
or U2918 (N_2918,N_843,N_873);
and U2919 (N_2919,N_1868,N_1661);
nor U2920 (N_2920,N_471,N_1517);
nor U2921 (N_2921,N_1163,N_1088);
and U2922 (N_2922,N_283,N_1160);
and U2923 (N_2923,N_657,N_44);
or U2924 (N_2924,N_1543,N_798);
nor U2925 (N_2925,N_108,N_889);
nor U2926 (N_2926,N_1915,N_200);
nand U2927 (N_2927,N_1617,N_514);
nor U2928 (N_2928,N_1072,N_335);
or U2929 (N_2929,N_266,N_191);
nor U2930 (N_2930,N_1866,N_1784);
and U2931 (N_2931,N_695,N_440);
nor U2932 (N_2932,N_1342,N_676);
nor U2933 (N_2933,N_1760,N_591);
nor U2934 (N_2934,N_682,N_1358);
nor U2935 (N_2935,N_752,N_1718);
nand U2936 (N_2936,N_180,N_379);
and U2937 (N_2937,N_1902,N_1685);
nand U2938 (N_2938,N_321,N_202);
nor U2939 (N_2939,N_1669,N_1992);
and U2940 (N_2940,N_1092,N_219);
nand U2941 (N_2941,N_1631,N_1922);
or U2942 (N_2942,N_1953,N_1841);
nor U2943 (N_2943,N_594,N_696);
nand U2944 (N_2944,N_581,N_1220);
nor U2945 (N_2945,N_1856,N_1039);
nand U2946 (N_2946,N_172,N_1036);
nor U2947 (N_2947,N_1686,N_404);
and U2948 (N_2948,N_1411,N_1596);
nand U2949 (N_2949,N_1410,N_1710);
nor U2950 (N_2950,N_1035,N_1894);
and U2951 (N_2951,N_393,N_1357);
nor U2952 (N_2952,N_1213,N_22);
and U2953 (N_2953,N_759,N_137);
and U2954 (N_2954,N_781,N_1294);
and U2955 (N_2955,N_241,N_1637);
nor U2956 (N_2956,N_255,N_1276);
nand U2957 (N_2957,N_82,N_1858);
nand U2958 (N_2958,N_1173,N_388);
nand U2959 (N_2959,N_1664,N_846);
nand U2960 (N_2960,N_863,N_987);
nand U2961 (N_2961,N_52,N_1645);
nand U2962 (N_2962,N_1563,N_72);
or U2963 (N_2963,N_705,N_132);
nand U2964 (N_2964,N_561,N_995);
and U2965 (N_2965,N_1983,N_364);
nor U2966 (N_2966,N_426,N_975);
nand U2967 (N_2967,N_548,N_511);
and U2968 (N_2968,N_945,N_167);
nor U2969 (N_2969,N_1026,N_1432);
and U2970 (N_2970,N_928,N_245);
nor U2971 (N_2971,N_1604,N_1328);
nor U2972 (N_2972,N_522,N_79);
or U2973 (N_2973,N_114,N_1237);
nor U2974 (N_2974,N_1020,N_722);
nor U2975 (N_2975,N_1824,N_1913);
nand U2976 (N_2976,N_939,N_1959);
or U2977 (N_2977,N_234,N_921);
nor U2978 (N_2978,N_1376,N_518);
nor U2979 (N_2979,N_1941,N_1900);
and U2980 (N_2980,N_1595,N_1046);
or U2981 (N_2981,N_839,N_1575);
nand U2982 (N_2982,N_1353,N_1295);
and U2983 (N_2983,N_1927,N_1040);
and U2984 (N_2984,N_356,N_487);
and U2985 (N_2985,N_434,N_1541);
nand U2986 (N_2986,N_289,N_15);
nand U2987 (N_2987,N_562,N_1260);
nor U2988 (N_2988,N_1698,N_1647);
and U2989 (N_2989,N_1780,N_1475);
nand U2990 (N_2990,N_1667,N_668);
or U2991 (N_2991,N_1768,N_1193);
nor U2992 (N_2992,N_744,N_1138);
nor U2993 (N_2993,N_1249,N_649);
and U2994 (N_2994,N_1488,N_1456);
and U2995 (N_2995,N_841,N_1778);
nand U2996 (N_2996,N_1234,N_896);
nor U2997 (N_2997,N_228,N_1064);
nand U2998 (N_2998,N_477,N_922);
nand U2999 (N_2999,N_1728,N_209);
or U3000 (N_3000,N_1553,N_179);
and U3001 (N_3001,N_1259,N_424);
and U3002 (N_3002,N_491,N_1680);
and U3003 (N_3003,N_1,N_391);
nand U3004 (N_3004,N_226,N_510);
nor U3005 (N_3005,N_1047,N_69);
nand U3006 (N_3006,N_1682,N_151);
or U3007 (N_3007,N_354,N_1086);
and U3008 (N_3008,N_72,N_1590);
nand U3009 (N_3009,N_943,N_1354);
or U3010 (N_3010,N_894,N_1599);
or U3011 (N_3011,N_1795,N_658);
nor U3012 (N_3012,N_1788,N_34);
and U3013 (N_3013,N_1428,N_307);
and U3014 (N_3014,N_560,N_240);
and U3015 (N_3015,N_388,N_1309);
nor U3016 (N_3016,N_922,N_953);
nor U3017 (N_3017,N_528,N_963);
and U3018 (N_3018,N_633,N_1258);
xor U3019 (N_3019,N_41,N_866);
nor U3020 (N_3020,N_587,N_1016);
or U3021 (N_3021,N_1326,N_1156);
or U3022 (N_3022,N_444,N_1906);
nor U3023 (N_3023,N_1562,N_1717);
and U3024 (N_3024,N_155,N_702);
nand U3025 (N_3025,N_346,N_990);
or U3026 (N_3026,N_1436,N_549);
nor U3027 (N_3027,N_229,N_279);
nand U3028 (N_3028,N_987,N_243);
nand U3029 (N_3029,N_1893,N_105);
nor U3030 (N_3030,N_427,N_782);
nor U3031 (N_3031,N_702,N_1161);
nor U3032 (N_3032,N_552,N_1260);
and U3033 (N_3033,N_28,N_147);
and U3034 (N_3034,N_1572,N_149);
nor U3035 (N_3035,N_1843,N_295);
nor U3036 (N_3036,N_532,N_1031);
or U3037 (N_3037,N_875,N_1507);
and U3038 (N_3038,N_909,N_543);
and U3039 (N_3039,N_1599,N_1348);
or U3040 (N_3040,N_1205,N_1625);
nor U3041 (N_3041,N_1962,N_763);
or U3042 (N_3042,N_1279,N_983);
and U3043 (N_3043,N_1735,N_1803);
or U3044 (N_3044,N_1474,N_650);
or U3045 (N_3045,N_154,N_1010);
nand U3046 (N_3046,N_379,N_615);
or U3047 (N_3047,N_1191,N_1704);
or U3048 (N_3048,N_46,N_1436);
nand U3049 (N_3049,N_495,N_1573);
nand U3050 (N_3050,N_1672,N_343);
nor U3051 (N_3051,N_512,N_303);
and U3052 (N_3052,N_1046,N_1881);
nand U3053 (N_3053,N_751,N_201);
or U3054 (N_3054,N_733,N_691);
nor U3055 (N_3055,N_1796,N_1223);
nor U3056 (N_3056,N_1410,N_1131);
and U3057 (N_3057,N_1973,N_914);
or U3058 (N_3058,N_611,N_1102);
or U3059 (N_3059,N_1553,N_1358);
and U3060 (N_3060,N_1090,N_1139);
and U3061 (N_3061,N_943,N_923);
nor U3062 (N_3062,N_1995,N_90);
or U3063 (N_3063,N_550,N_504);
or U3064 (N_3064,N_613,N_864);
nand U3065 (N_3065,N_1925,N_24);
nand U3066 (N_3066,N_903,N_1633);
nand U3067 (N_3067,N_837,N_1475);
xnor U3068 (N_3068,N_1211,N_501);
nor U3069 (N_3069,N_1642,N_244);
nand U3070 (N_3070,N_1104,N_1596);
and U3071 (N_3071,N_1244,N_1266);
or U3072 (N_3072,N_1833,N_1264);
nand U3073 (N_3073,N_855,N_1262);
and U3074 (N_3074,N_354,N_1644);
nand U3075 (N_3075,N_1039,N_740);
and U3076 (N_3076,N_549,N_1339);
nor U3077 (N_3077,N_940,N_1449);
nand U3078 (N_3078,N_1338,N_1693);
nor U3079 (N_3079,N_1880,N_405);
xnor U3080 (N_3080,N_1138,N_1467);
nor U3081 (N_3081,N_1030,N_80);
nand U3082 (N_3082,N_1299,N_664);
or U3083 (N_3083,N_1049,N_24);
nand U3084 (N_3084,N_1129,N_1237);
or U3085 (N_3085,N_861,N_1388);
or U3086 (N_3086,N_1432,N_1679);
or U3087 (N_3087,N_1743,N_371);
nand U3088 (N_3088,N_52,N_1978);
or U3089 (N_3089,N_322,N_1305);
or U3090 (N_3090,N_69,N_1821);
and U3091 (N_3091,N_18,N_1869);
or U3092 (N_3092,N_1419,N_1528);
and U3093 (N_3093,N_1883,N_1349);
nor U3094 (N_3094,N_1256,N_504);
nand U3095 (N_3095,N_938,N_719);
nor U3096 (N_3096,N_154,N_1288);
nor U3097 (N_3097,N_1647,N_213);
or U3098 (N_3098,N_1538,N_682);
and U3099 (N_3099,N_1483,N_1450);
nand U3100 (N_3100,N_763,N_1068);
or U3101 (N_3101,N_1373,N_1523);
nand U3102 (N_3102,N_496,N_629);
nand U3103 (N_3103,N_1430,N_835);
nand U3104 (N_3104,N_148,N_1123);
nor U3105 (N_3105,N_1567,N_322);
and U3106 (N_3106,N_1147,N_1661);
nor U3107 (N_3107,N_239,N_1233);
nor U3108 (N_3108,N_139,N_387);
and U3109 (N_3109,N_204,N_1139);
nand U3110 (N_3110,N_284,N_633);
and U3111 (N_3111,N_710,N_719);
and U3112 (N_3112,N_365,N_1152);
and U3113 (N_3113,N_408,N_913);
and U3114 (N_3114,N_713,N_1618);
or U3115 (N_3115,N_114,N_354);
nor U3116 (N_3116,N_1075,N_1134);
nor U3117 (N_3117,N_1855,N_1620);
nor U3118 (N_3118,N_391,N_1556);
nand U3119 (N_3119,N_431,N_1221);
and U3120 (N_3120,N_900,N_1439);
nand U3121 (N_3121,N_1777,N_1315);
nand U3122 (N_3122,N_229,N_352);
nand U3123 (N_3123,N_1691,N_66);
or U3124 (N_3124,N_994,N_8);
and U3125 (N_3125,N_1636,N_1257);
nand U3126 (N_3126,N_1944,N_342);
nand U3127 (N_3127,N_1805,N_1469);
or U3128 (N_3128,N_1966,N_1209);
or U3129 (N_3129,N_274,N_848);
or U3130 (N_3130,N_458,N_755);
nor U3131 (N_3131,N_1387,N_1566);
or U3132 (N_3132,N_412,N_1612);
nor U3133 (N_3133,N_969,N_387);
and U3134 (N_3134,N_926,N_275);
nand U3135 (N_3135,N_1133,N_475);
or U3136 (N_3136,N_1142,N_556);
and U3137 (N_3137,N_1741,N_1006);
nor U3138 (N_3138,N_1489,N_10);
or U3139 (N_3139,N_918,N_1545);
and U3140 (N_3140,N_1611,N_377);
and U3141 (N_3141,N_434,N_1616);
nand U3142 (N_3142,N_687,N_729);
or U3143 (N_3143,N_614,N_547);
and U3144 (N_3144,N_1035,N_1807);
and U3145 (N_3145,N_41,N_531);
nor U3146 (N_3146,N_783,N_1379);
and U3147 (N_3147,N_1972,N_37);
and U3148 (N_3148,N_1716,N_24);
and U3149 (N_3149,N_726,N_1941);
nor U3150 (N_3150,N_1340,N_1398);
or U3151 (N_3151,N_1484,N_766);
and U3152 (N_3152,N_1896,N_1153);
nor U3153 (N_3153,N_1182,N_617);
and U3154 (N_3154,N_969,N_1271);
nor U3155 (N_3155,N_491,N_533);
nand U3156 (N_3156,N_110,N_528);
nor U3157 (N_3157,N_532,N_1584);
nor U3158 (N_3158,N_921,N_1402);
or U3159 (N_3159,N_1781,N_922);
nor U3160 (N_3160,N_1221,N_1677);
nand U3161 (N_3161,N_335,N_485);
nand U3162 (N_3162,N_867,N_761);
nor U3163 (N_3163,N_1401,N_1720);
or U3164 (N_3164,N_1265,N_1342);
or U3165 (N_3165,N_1662,N_1062);
and U3166 (N_3166,N_1754,N_366);
nor U3167 (N_3167,N_1042,N_236);
and U3168 (N_3168,N_1612,N_1000);
or U3169 (N_3169,N_1425,N_441);
or U3170 (N_3170,N_916,N_781);
and U3171 (N_3171,N_1025,N_170);
nor U3172 (N_3172,N_1242,N_1103);
and U3173 (N_3173,N_223,N_1257);
and U3174 (N_3174,N_1087,N_1504);
or U3175 (N_3175,N_1921,N_523);
nand U3176 (N_3176,N_1772,N_282);
nor U3177 (N_3177,N_50,N_1961);
nor U3178 (N_3178,N_634,N_1791);
and U3179 (N_3179,N_185,N_736);
nor U3180 (N_3180,N_447,N_1045);
nor U3181 (N_3181,N_467,N_810);
and U3182 (N_3182,N_754,N_1356);
and U3183 (N_3183,N_836,N_1331);
and U3184 (N_3184,N_552,N_1078);
and U3185 (N_3185,N_1791,N_308);
nand U3186 (N_3186,N_44,N_1791);
and U3187 (N_3187,N_1949,N_1437);
nand U3188 (N_3188,N_581,N_419);
or U3189 (N_3189,N_301,N_750);
or U3190 (N_3190,N_168,N_1831);
nor U3191 (N_3191,N_1957,N_1195);
and U3192 (N_3192,N_1081,N_1846);
or U3193 (N_3193,N_401,N_1657);
nand U3194 (N_3194,N_1662,N_1816);
and U3195 (N_3195,N_465,N_876);
or U3196 (N_3196,N_1142,N_819);
or U3197 (N_3197,N_1111,N_727);
and U3198 (N_3198,N_1327,N_1823);
or U3199 (N_3199,N_161,N_1877);
or U3200 (N_3200,N_733,N_1498);
and U3201 (N_3201,N_455,N_1793);
nor U3202 (N_3202,N_1241,N_482);
or U3203 (N_3203,N_1612,N_175);
nand U3204 (N_3204,N_105,N_1220);
and U3205 (N_3205,N_996,N_1321);
and U3206 (N_3206,N_136,N_863);
or U3207 (N_3207,N_210,N_819);
nand U3208 (N_3208,N_76,N_620);
nor U3209 (N_3209,N_1712,N_1968);
or U3210 (N_3210,N_471,N_1625);
nand U3211 (N_3211,N_1208,N_486);
and U3212 (N_3212,N_1691,N_1354);
nand U3213 (N_3213,N_1325,N_1221);
nand U3214 (N_3214,N_581,N_387);
or U3215 (N_3215,N_763,N_1497);
or U3216 (N_3216,N_32,N_401);
and U3217 (N_3217,N_410,N_881);
and U3218 (N_3218,N_741,N_1642);
or U3219 (N_3219,N_1195,N_1727);
nor U3220 (N_3220,N_1082,N_132);
nor U3221 (N_3221,N_805,N_1409);
nand U3222 (N_3222,N_197,N_1830);
nand U3223 (N_3223,N_347,N_219);
xor U3224 (N_3224,N_1481,N_76);
and U3225 (N_3225,N_525,N_825);
and U3226 (N_3226,N_185,N_558);
nand U3227 (N_3227,N_1645,N_1377);
xnor U3228 (N_3228,N_199,N_857);
nand U3229 (N_3229,N_365,N_1562);
nor U3230 (N_3230,N_1381,N_1546);
nor U3231 (N_3231,N_1991,N_534);
or U3232 (N_3232,N_1697,N_1142);
nor U3233 (N_3233,N_904,N_1743);
or U3234 (N_3234,N_47,N_687);
or U3235 (N_3235,N_1050,N_1241);
and U3236 (N_3236,N_1176,N_1638);
or U3237 (N_3237,N_350,N_1503);
nor U3238 (N_3238,N_1241,N_1866);
and U3239 (N_3239,N_895,N_665);
and U3240 (N_3240,N_327,N_95);
or U3241 (N_3241,N_1605,N_1979);
nor U3242 (N_3242,N_1211,N_1193);
or U3243 (N_3243,N_1955,N_715);
and U3244 (N_3244,N_410,N_432);
or U3245 (N_3245,N_1483,N_1733);
nand U3246 (N_3246,N_1666,N_1047);
or U3247 (N_3247,N_282,N_316);
or U3248 (N_3248,N_1236,N_1193);
nor U3249 (N_3249,N_1527,N_61);
or U3250 (N_3250,N_450,N_1361);
and U3251 (N_3251,N_1837,N_133);
nand U3252 (N_3252,N_108,N_277);
nand U3253 (N_3253,N_1085,N_1445);
nand U3254 (N_3254,N_164,N_1055);
and U3255 (N_3255,N_1996,N_1807);
or U3256 (N_3256,N_721,N_1159);
nor U3257 (N_3257,N_915,N_1634);
nor U3258 (N_3258,N_1407,N_631);
or U3259 (N_3259,N_346,N_1880);
or U3260 (N_3260,N_1070,N_739);
nand U3261 (N_3261,N_1401,N_1977);
nor U3262 (N_3262,N_1053,N_1444);
nand U3263 (N_3263,N_1105,N_458);
or U3264 (N_3264,N_1805,N_2);
nor U3265 (N_3265,N_531,N_1800);
nand U3266 (N_3266,N_1764,N_1072);
and U3267 (N_3267,N_1252,N_220);
nand U3268 (N_3268,N_481,N_593);
nand U3269 (N_3269,N_236,N_696);
and U3270 (N_3270,N_56,N_701);
and U3271 (N_3271,N_1619,N_959);
nand U3272 (N_3272,N_398,N_762);
nor U3273 (N_3273,N_1348,N_1880);
nand U3274 (N_3274,N_1919,N_919);
and U3275 (N_3275,N_1396,N_1761);
nor U3276 (N_3276,N_250,N_548);
nor U3277 (N_3277,N_744,N_1117);
nand U3278 (N_3278,N_1514,N_1856);
and U3279 (N_3279,N_1236,N_1567);
nor U3280 (N_3280,N_422,N_1228);
and U3281 (N_3281,N_1775,N_807);
nor U3282 (N_3282,N_82,N_1768);
and U3283 (N_3283,N_358,N_1708);
nand U3284 (N_3284,N_1766,N_725);
and U3285 (N_3285,N_313,N_1036);
nand U3286 (N_3286,N_1330,N_887);
and U3287 (N_3287,N_713,N_1733);
and U3288 (N_3288,N_605,N_1851);
nand U3289 (N_3289,N_327,N_906);
or U3290 (N_3290,N_833,N_1069);
nor U3291 (N_3291,N_967,N_1746);
nor U3292 (N_3292,N_1965,N_281);
and U3293 (N_3293,N_1468,N_1056);
or U3294 (N_3294,N_1139,N_1288);
or U3295 (N_3295,N_1270,N_1803);
nand U3296 (N_3296,N_1309,N_552);
nand U3297 (N_3297,N_555,N_202);
and U3298 (N_3298,N_1675,N_1359);
or U3299 (N_3299,N_2,N_1583);
nor U3300 (N_3300,N_1599,N_864);
nor U3301 (N_3301,N_1992,N_550);
nor U3302 (N_3302,N_1248,N_1638);
and U3303 (N_3303,N_375,N_1947);
nor U3304 (N_3304,N_244,N_1896);
nand U3305 (N_3305,N_1503,N_1145);
or U3306 (N_3306,N_470,N_1473);
nand U3307 (N_3307,N_1478,N_1643);
or U3308 (N_3308,N_1716,N_595);
nor U3309 (N_3309,N_1290,N_1739);
or U3310 (N_3310,N_1460,N_123);
nor U3311 (N_3311,N_1025,N_1861);
nand U3312 (N_3312,N_1690,N_353);
and U3313 (N_3313,N_236,N_527);
nand U3314 (N_3314,N_166,N_562);
nor U3315 (N_3315,N_1624,N_108);
nor U3316 (N_3316,N_1731,N_556);
nor U3317 (N_3317,N_1510,N_1283);
and U3318 (N_3318,N_62,N_378);
or U3319 (N_3319,N_1961,N_16);
or U3320 (N_3320,N_830,N_1839);
nor U3321 (N_3321,N_263,N_727);
or U3322 (N_3322,N_102,N_1168);
nor U3323 (N_3323,N_851,N_496);
or U3324 (N_3324,N_690,N_834);
or U3325 (N_3325,N_1495,N_900);
nand U3326 (N_3326,N_606,N_322);
nand U3327 (N_3327,N_588,N_18);
nand U3328 (N_3328,N_88,N_689);
nand U3329 (N_3329,N_614,N_1824);
nor U3330 (N_3330,N_1538,N_513);
nand U3331 (N_3331,N_1826,N_1298);
or U3332 (N_3332,N_1867,N_631);
nor U3333 (N_3333,N_852,N_527);
or U3334 (N_3334,N_844,N_350);
nand U3335 (N_3335,N_402,N_1336);
nand U3336 (N_3336,N_964,N_1286);
nor U3337 (N_3337,N_1032,N_507);
xnor U3338 (N_3338,N_800,N_1022);
nor U3339 (N_3339,N_817,N_166);
nor U3340 (N_3340,N_295,N_904);
or U3341 (N_3341,N_690,N_1096);
nand U3342 (N_3342,N_1892,N_376);
and U3343 (N_3343,N_609,N_138);
nor U3344 (N_3344,N_1124,N_1049);
nor U3345 (N_3345,N_1926,N_1976);
and U3346 (N_3346,N_1549,N_11);
or U3347 (N_3347,N_1548,N_627);
nand U3348 (N_3348,N_489,N_381);
nor U3349 (N_3349,N_437,N_1738);
and U3350 (N_3350,N_502,N_1866);
nor U3351 (N_3351,N_378,N_1288);
nand U3352 (N_3352,N_268,N_184);
nor U3353 (N_3353,N_1065,N_1731);
nand U3354 (N_3354,N_1007,N_1508);
or U3355 (N_3355,N_1550,N_968);
nor U3356 (N_3356,N_1907,N_161);
and U3357 (N_3357,N_887,N_1014);
nand U3358 (N_3358,N_172,N_214);
and U3359 (N_3359,N_946,N_775);
and U3360 (N_3360,N_1266,N_1898);
nor U3361 (N_3361,N_1777,N_414);
or U3362 (N_3362,N_1599,N_1289);
or U3363 (N_3363,N_1519,N_886);
nand U3364 (N_3364,N_652,N_1483);
or U3365 (N_3365,N_1866,N_643);
nor U3366 (N_3366,N_139,N_968);
nand U3367 (N_3367,N_1631,N_1714);
and U3368 (N_3368,N_453,N_1511);
nor U3369 (N_3369,N_1142,N_502);
nand U3370 (N_3370,N_1624,N_1332);
nand U3371 (N_3371,N_1801,N_1209);
nor U3372 (N_3372,N_1638,N_548);
nor U3373 (N_3373,N_788,N_1918);
nor U3374 (N_3374,N_1270,N_501);
or U3375 (N_3375,N_1525,N_935);
or U3376 (N_3376,N_1927,N_1414);
or U3377 (N_3377,N_1334,N_544);
and U3378 (N_3378,N_1501,N_1487);
or U3379 (N_3379,N_956,N_82);
or U3380 (N_3380,N_12,N_817);
nand U3381 (N_3381,N_956,N_1256);
and U3382 (N_3382,N_693,N_1963);
and U3383 (N_3383,N_1606,N_376);
nor U3384 (N_3384,N_371,N_724);
xor U3385 (N_3385,N_104,N_115);
and U3386 (N_3386,N_1711,N_31);
and U3387 (N_3387,N_1790,N_118);
and U3388 (N_3388,N_144,N_1499);
and U3389 (N_3389,N_1025,N_814);
or U3390 (N_3390,N_914,N_1309);
nor U3391 (N_3391,N_1017,N_424);
nor U3392 (N_3392,N_364,N_519);
nor U3393 (N_3393,N_816,N_930);
and U3394 (N_3394,N_1238,N_238);
and U3395 (N_3395,N_1316,N_298);
nor U3396 (N_3396,N_1833,N_1331);
or U3397 (N_3397,N_378,N_1767);
nand U3398 (N_3398,N_1272,N_1346);
or U3399 (N_3399,N_1657,N_1854);
nand U3400 (N_3400,N_1510,N_721);
or U3401 (N_3401,N_674,N_905);
and U3402 (N_3402,N_1086,N_777);
or U3403 (N_3403,N_169,N_906);
xnor U3404 (N_3404,N_1084,N_116);
nand U3405 (N_3405,N_961,N_573);
or U3406 (N_3406,N_933,N_1299);
and U3407 (N_3407,N_26,N_383);
or U3408 (N_3408,N_1999,N_1158);
nand U3409 (N_3409,N_389,N_1358);
or U3410 (N_3410,N_24,N_444);
nand U3411 (N_3411,N_37,N_1775);
nor U3412 (N_3412,N_346,N_1036);
and U3413 (N_3413,N_676,N_1822);
or U3414 (N_3414,N_1331,N_673);
nor U3415 (N_3415,N_352,N_982);
and U3416 (N_3416,N_453,N_1722);
nor U3417 (N_3417,N_1558,N_1432);
xnor U3418 (N_3418,N_925,N_31);
nor U3419 (N_3419,N_847,N_1041);
nor U3420 (N_3420,N_1454,N_369);
and U3421 (N_3421,N_511,N_65);
or U3422 (N_3422,N_1466,N_1045);
and U3423 (N_3423,N_928,N_1682);
or U3424 (N_3424,N_430,N_582);
or U3425 (N_3425,N_230,N_1186);
nand U3426 (N_3426,N_685,N_894);
or U3427 (N_3427,N_372,N_1148);
and U3428 (N_3428,N_373,N_517);
and U3429 (N_3429,N_1266,N_1770);
nor U3430 (N_3430,N_47,N_1142);
nand U3431 (N_3431,N_831,N_1115);
nand U3432 (N_3432,N_957,N_784);
nor U3433 (N_3433,N_799,N_399);
or U3434 (N_3434,N_1472,N_394);
or U3435 (N_3435,N_509,N_1608);
and U3436 (N_3436,N_554,N_61);
nor U3437 (N_3437,N_685,N_1199);
nand U3438 (N_3438,N_1445,N_1808);
and U3439 (N_3439,N_1608,N_1048);
nand U3440 (N_3440,N_1005,N_432);
nand U3441 (N_3441,N_1001,N_30);
or U3442 (N_3442,N_250,N_1666);
and U3443 (N_3443,N_1658,N_1746);
nor U3444 (N_3444,N_1054,N_1648);
nor U3445 (N_3445,N_344,N_1254);
or U3446 (N_3446,N_1022,N_1125);
and U3447 (N_3447,N_980,N_808);
or U3448 (N_3448,N_105,N_553);
nand U3449 (N_3449,N_1455,N_255);
nand U3450 (N_3450,N_1410,N_1362);
and U3451 (N_3451,N_1863,N_1949);
nor U3452 (N_3452,N_346,N_167);
nand U3453 (N_3453,N_673,N_941);
nor U3454 (N_3454,N_1692,N_1408);
or U3455 (N_3455,N_1407,N_530);
or U3456 (N_3456,N_1379,N_397);
nor U3457 (N_3457,N_1124,N_674);
and U3458 (N_3458,N_906,N_1205);
and U3459 (N_3459,N_834,N_1307);
nor U3460 (N_3460,N_1486,N_848);
nor U3461 (N_3461,N_318,N_1486);
nor U3462 (N_3462,N_999,N_748);
nand U3463 (N_3463,N_60,N_208);
or U3464 (N_3464,N_1198,N_229);
nand U3465 (N_3465,N_1486,N_232);
nand U3466 (N_3466,N_218,N_1428);
nor U3467 (N_3467,N_97,N_1309);
nand U3468 (N_3468,N_659,N_117);
and U3469 (N_3469,N_1104,N_1277);
nor U3470 (N_3470,N_1012,N_744);
xor U3471 (N_3471,N_511,N_1529);
and U3472 (N_3472,N_637,N_1258);
nor U3473 (N_3473,N_37,N_1467);
nor U3474 (N_3474,N_294,N_996);
nand U3475 (N_3475,N_1648,N_1736);
or U3476 (N_3476,N_1107,N_1579);
or U3477 (N_3477,N_1760,N_1474);
nor U3478 (N_3478,N_1357,N_923);
nand U3479 (N_3479,N_912,N_1358);
nand U3480 (N_3480,N_543,N_1190);
and U3481 (N_3481,N_574,N_311);
and U3482 (N_3482,N_1914,N_1271);
nand U3483 (N_3483,N_1674,N_1837);
nand U3484 (N_3484,N_161,N_638);
or U3485 (N_3485,N_1995,N_1301);
or U3486 (N_3486,N_988,N_409);
or U3487 (N_3487,N_947,N_1036);
nand U3488 (N_3488,N_613,N_1855);
nor U3489 (N_3489,N_1074,N_1060);
or U3490 (N_3490,N_1626,N_67);
nand U3491 (N_3491,N_744,N_1986);
nand U3492 (N_3492,N_218,N_105);
nand U3493 (N_3493,N_760,N_1720);
nand U3494 (N_3494,N_1727,N_1673);
nand U3495 (N_3495,N_795,N_1478);
xnor U3496 (N_3496,N_1609,N_1612);
nand U3497 (N_3497,N_1889,N_1826);
nand U3498 (N_3498,N_1166,N_1157);
or U3499 (N_3499,N_1159,N_632);
nor U3500 (N_3500,N_1469,N_1445);
or U3501 (N_3501,N_1661,N_292);
or U3502 (N_3502,N_1506,N_378);
or U3503 (N_3503,N_1564,N_1131);
or U3504 (N_3504,N_386,N_95);
xor U3505 (N_3505,N_172,N_536);
or U3506 (N_3506,N_819,N_31);
and U3507 (N_3507,N_301,N_119);
and U3508 (N_3508,N_1445,N_1974);
nor U3509 (N_3509,N_1617,N_265);
nor U3510 (N_3510,N_1693,N_1295);
or U3511 (N_3511,N_1582,N_937);
nand U3512 (N_3512,N_1710,N_31);
nor U3513 (N_3513,N_1611,N_1736);
nor U3514 (N_3514,N_1658,N_861);
and U3515 (N_3515,N_1262,N_656);
nand U3516 (N_3516,N_1288,N_269);
nand U3517 (N_3517,N_1592,N_1339);
or U3518 (N_3518,N_1569,N_1464);
nand U3519 (N_3519,N_435,N_69);
nand U3520 (N_3520,N_1390,N_1060);
or U3521 (N_3521,N_737,N_1125);
or U3522 (N_3522,N_772,N_1464);
nor U3523 (N_3523,N_823,N_625);
or U3524 (N_3524,N_1102,N_542);
nand U3525 (N_3525,N_1168,N_744);
or U3526 (N_3526,N_704,N_669);
nor U3527 (N_3527,N_1833,N_1261);
or U3528 (N_3528,N_1289,N_151);
or U3529 (N_3529,N_641,N_111);
nand U3530 (N_3530,N_1860,N_451);
and U3531 (N_3531,N_280,N_1309);
and U3532 (N_3532,N_1238,N_1778);
nand U3533 (N_3533,N_1892,N_1344);
nand U3534 (N_3534,N_952,N_462);
and U3535 (N_3535,N_504,N_1419);
and U3536 (N_3536,N_1436,N_4);
nand U3537 (N_3537,N_517,N_1211);
nor U3538 (N_3538,N_1128,N_1331);
and U3539 (N_3539,N_1162,N_1367);
nor U3540 (N_3540,N_224,N_667);
and U3541 (N_3541,N_1870,N_1159);
or U3542 (N_3542,N_57,N_1601);
or U3543 (N_3543,N_1332,N_110);
nand U3544 (N_3544,N_357,N_1035);
or U3545 (N_3545,N_367,N_810);
and U3546 (N_3546,N_522,N_618);
or U3547 (N_3547,N_1447,N_1068);
and U3548 (N_3548,N_129,N_1234);
or U3549 (N_3549,N_1880,N_174);
and U3550 (N_3550,N_343,N_231);
nand U3551 (N_3551,N_904,N_1563);
nand U3552 (N_3552,N_1341,N_492);
or U3553 (N_3553,N_1262,N_1937);
and U3554 (N_3554,N_172,N_1389);
nor U3555 (N_3555,N_1349,N_49);
or U3556 (N_3556,N_1482,N_982);
or U3557 (N_3557,N_563,N_375);
or U3558 (N_3558,N_1561,N_83);
and U3559 (N_3559,N_319,N_1180);
nor U3560 (N_3560,N_1944,N_1075);
nor U3561 (N_3561,N_713,N_1873);
or U3562 (N_3562,N_918,N_451);
nand U3563 (N_3563,N_970,N_116);
and U3564 (N_3564,N_203,N_718);
nor U3565 (N_3565,N_223,N_554);
and U3566 (N_3566,N_1328,N_1822);
nand U3567 (N_3567,N_65,N_271);
nand U3568 (N_3568,N_1636,N_284);
nor U3569 (N_3569,N_158,N_355);
or U3570 (N_3570,N_1686,N_1591);
and U3571 (N_3571,N_986,N_625);
nand U3572 (N_3572,N_1534,N_792);
nor U3573 (N_3573,N_1582,N_1656);
and U3574 (N_3574,N_1219,N_199);
or U3575 (N_3575,N_1754,N_49);
and U3576 (N_3576,N_1280,N_1215);
nand U3577 (N_3577,N_775,N_1849);
nor U3578 (N_3578,N_978,N_1270);
and U3579 (N_3579,N_976,N_1368);
or U3580 (N_3580,N_1771,N_1629);
nand U3581 (N_3581,N_1053,N_208);
nor U3582 (N_3582,N_1089,N_1739);
nand U3583 (N_3583,N_1621,N_662);
and U3584 (N_3584,N_1889,N_1146);
or U3585 (N_3585,N_1820,N_1905);
nor U3586 (N_3586,N_395,N_538);
or U3587 (N_3587,N_1873,N_910);
nand U3588 (N_3588,N_159,N_156);
nor U3589 (N_3589,N_40,N_1779);
and U3590 (N_3590,N_461,N_1505);
or U3591 (N_3591,N_1790,N_1181);
nand U3592 (N_3592,N_358,N_295);
or U3593 (N_3593,N_1214,N_1964);
nor U3594 (N_3594,N_1888,N_828);
or U3595 (N_3595,N_1050,N_1017);
nor U3596 (N_3596,N_1064,N_848);
or U3597 (N_3597,N_1033,N_83);
nand U3598 (N_3598,N_479,N_1888);
nor U3599 (N_3599,N_33,N_552);
nand U3600 (N_3600,N_786,N_76);
or U3601 (N_3601,N_1407,N_1918);
nand U3602 (N_3602,N_398,N_770);
and U3603 (N_3603,N_1836,N_889);
and U3604 (N_3604,N_299,N_1266);
nand U3605 (N_3605,N_719,N_1146);
or U3606 (N_3606,N_1292,N_1410);
and U3607 (N_3607,N_521,N_1381);
and U3608 (N_3608,N_262,N_776);
nand U3609 (N_3609,N_1647,N_728);
and U3610 (N_3610,N_549,N_173);
or U3611 (N_3611,N_1914,N_1924);
or U3612 (N_3612,N_1678,N_1723);
nor U3613 (N_3613,N_307,N_1950);
nand U3614 (N_3614,N_1382,N_596);
nor U3615 (N_3615,N_1881,N_1954);
nor U3616 (N_3616,N_1658,N_477);
and U3617 (N_3617,N_1252,N_418);
and U3618 (N_3618,N_206,N_438);
nand U3619 (N_3619,N_95,N_255);
or U3620 (N_3620,N_726,N_652);
nand U3621 (N_3621,N_575,N_1568);
or U3622 (N_3622,N_1817,N_1482);
or U3623 (N_3623,N_1186,N_1299);
nand U3624 (N_3624,N_96,N_1688);
and U3625 (N_3625,N_1764,N_1238);
nand U3626 (N_3626,N_226,N_1562);
nand U3627 (N_3627,N_1692,N_1535);
nor U3628 (N_3628,N_1665,N_712);
nor U3629 (N_3629,N_1425,N_1662);
nand U3630 (N_3630,N_1632,N_302);
nand U3631 (N_3631,N_1936,N_391);
or U3632 (N_3632,N_601,N_462);
and U3633 (N_3633,N_1070,N_253);
or U3634 (N_3634,N_1085,N_160);
nand U3635 (N_3635,N_82,N_15);
nand U3636 (N_3636,N_1443,N_1056);
and U3637 (N_3637,N_1735,N_926);
nor U3638 (N_3638,N_342,N_502);
and U3639 (N_3639,N_751,N_1641);
nand U3640 (N_3640,N_1721,N_1648);
and U3641 (N_3641,N_661,N_538);
or U3642 (N_3642,N_1970,N_1681);
or U3643 (N_3643,N_133,N_1376);
or U3644 (N_3644,N_586,N_1299);
or U3645 (N_3645,N_195,N_63);
or U3646 (N_3646,N_927,N_460);
or U3647 (N_3647,N_313,N_1433);
or U3648 (N_3648,N_939,N_28);
nand U3649 (N_3649,N_1262,N_1338);
nor U3650 (N_3650,N_1839,N_473);
nor U3651 (N_3651,N_205,N_1357);
and U3652 (N_3652,N_1372,N_1079);
or U3653 (N_3653,N_80,N_726);
and U3654 (N_3654,N_1954,N_949);
or U3655 (N_3655,N_1818,N_128);
nand U3656 (N_3656,N_1511,N_1871);
or U3657 (N_3657,N_877,N_138);
nand U3658 (N_3658,N_1934,N_1424);
or U3659 (N_3659,N_1013,N_540);
nor U3660 (N_3660,N_240,N_175);
and U3661 (N_3661,N_186,N_1463);
nor U3662 (N_3662,N_1056,N_672);
nor U3663 (N_3663,N_708,N_1967);
and U3664 (N_3664,N_636,N_1134);
nor U3665 (N_3665,N_224,N_1469);
nor U3666 (N_3666,N_1626,N_481);
and U3667 (N_3667,N_449,N_181);
or U3668 (N_3668,N_997,N_1041);
and U3669 (N_3669,N_518,N_1720);
or U3670 (N_3670,N_496,N_1928);
nand U3671 (N_3671,N_1304,N_1804);
or U3672 (N_3672,N_366,N_1877);
nand U3673 (N_3673,N_1972,N_679);
nor U3674 (N_3674,N_790,N_755);
nor U3675 (N_3675,N_1293,N_310);
nor U3676 (N_3676,N_182,N_588);
and U3677 (N_3677,N_12,N_1131);
or U3678 (N_3678,N_214,N_784);
or U3679 (N_3679,N_868,N_1299);
or U3680 (N_3680,N_48,N_1630);
or U3681 (N_3681,N_1662,N_752);
nor U3682 (N_3682,N_1660,N_372);
nand U3683 (N_3683,N_851,N_709);
or U3684 (N_3684,N_1578,N_232);
or U3685 (N_3685,N_148,N_1353);
or U3686 (N_3686,N_136,N_91);
nor U3687 (N_3687,N_1867,N_350);
and U3688 (N_3688,N_1329,N_1106);
nor U3689 (N_3689,N_762,N_109);
and U3690 (N_3690,N_43,N_1631);
and U3691 (N_3691,N_1906,N_628);
nand U3692 (N_3692,N_743,N_1469);
nor U3693 (N_3693,N_1935,N_957);
and U3694 (N_3694,N_211,N_1583);
and U3695 (N_3695,N_141,N_1142);
nor U3696 (N_3696,N_1139,N_1921);
or U3697 (N_3697,N_630,N_640);
or U3698 (N_3698,N_371,N_1917);
or U3699 (N_3699,N_225,N_1593);
nand U3700 (N_3700,N_803,N_1591);
nand U3701 (N_3701,N_873,N_1739);
nor U3702 (N_3702,N_218,N_709);
nand U3703 (N_3703,N_794,N_1602);
nand U3704 (N_3704,N_438,N_1571);
nor U3705 (N_3705,N_942,N_1347);
nor U3706 (N_3706,N_1349,N_75);
and U3707 (N_3707,N_832,N_881);
or U3708 (N_3708,N_1849,N_1893);
nand U3709 (N_3709,N_1106,N_1173);
or U3710 (N_3710,N_1641,N_1487);
and U3711 (N_3711,N_1963,N_1079);
and U3712 (N_3712,N_193,N_947);
nor U3713 (N_3713,N_179,N_1452);
or U3714 (N_3714,N_845,N_574);
and U3715 (N_3715,N_278,N_1639);
or U3716 (N_3716,N_1166,N_541);
and U3717 (N_3717,N_936,N_54);
and U3718 (N_3718,N_252,N_5);
nand U3719 (N_3719,N_424,N_1012);
nor U3720 (N_3720,N_977,N_562);
nand U3721 (N_3721,N_1099,N_383);
or U3722 (N_3722,N_1803,N_975);
or U3723 (N_3723,N_1208,N_469);
or U3724 (N_3724,N_597,N_479);
nand U3725 (N_3725,N_1843,N_361);
nor U3726 (N_3726,N_1970,N_1996);
nor U3727 (N_3727,N_1361,N_43);
or U3728 (N_3728,N_737,N_1518);
nor U3729 (N_3729,N_1758,N_962);
nand U3730 (N_3730,N_1862,N_644);
and U3731 (N_3731,N_1333,N_1773);
and U3732 (N_3732,N_757,N_1415);
nor U3733 (N_3733,N_1673,N_1045);
and U3734 (N_3734,N_1887,N_1135);
or U3735 (N_3735,N_526,N_42);
or U3736 (N_3736,N_1084,N_566);
and U3737 (N_3737,N_627,N_1594);
or U3738 (N_3738,N_35,N_925);
nor U3739 (N_3739,N_1659,N_59);
nor U3740 (N_3740,N_785,N_190);
nor U3741 (N_3741,N_711,N_1082);
nor U3742 (N_3742,N_997,N_1746);
nor U3743 (N_3743,N_1127,N_1533);
or U3744 (N_3744,N_498,N_299);
or U3745 (N_3745,N_1486,N_120);
nor U3746 (N_3746,N_1941,N_202);
nand U3747 (N_3747,N_137,N_1282);
nand U3748 (N_3748,N_1201,N_1700);
nor U3749 (N_3749,N_1431,N_1574);
and U3750 (N_3750,N_332,N_47);
or U3751 (N_3751,N_1766,N_1735);
nand U3752 (N_3752,N_1214,N_499);
nor U3753 (N_3753,N_1450,N_854);
nor U3754 (N_3754,N_270,N_1244);
or U3755 (N_3755,N_979,N_587);
nand U3756 (N_3756,N_817,N_395);
and U3757 (N_3757,N_1350,N_1143);
nand U3758 (N_3758,N_674,N_705);
nand U3759 (N_3759,N_1430,N_1171);
nand U3760 (N_3760,N_1504,N_1899);
nand U3761 (N_3761,N_270,N_1573);
or U3762 (N_3762,N_1673,N_997);
or U3763 (N_3763,N_1366,N_311);
or U3764 (N_3764,N_1797,N_584);
or U3765 (N_3765,N_118,N_1324);
or U3766 (N_3766,N_258,N_581);
or U3767 (N_3767,N_1050,N_1354);
or U3768 (N_3768,N_1729,N_648);
or U3769 (N_3769,N_1207,N_904);
nand U3770 (N_3770,N_1067,N_20);
nor U3771 (N_3771,N_1563,N_1810);
and U3772 (N_3772,N_833,N_375);
nand U3773 (N_3773,N_337,N_1716);
nand U3774 (N_3774,N_1498,N_1370);
nor U3775 (N_3775,N_551,N_666);
nor U3776 (N_3776,N_1736,N_748);
nor U3777 (N_3777,N_539,N_139);
and U3778 (N_3778,N_82,N_168);
or U3779 (N_3779,N_1333,N_530);
nand U3780 (N_3780,N_207,N_1948);
nor U3781 (N_3781,N_48,N_1104);
nor U3782 (N_3782,N_1939,N_128);
nand U3783 (N_3783,N_529,N_939);
and U3784 (N_3784,N_1183,N_880);
nor U3785 (N_3785,N_904,N_1527);
nor U3786 (N_3786,N_1407,N_438);
and U3787 (N_3787,N_183,N_161);
nor U3788 (N_3788,N_809,N_687);
or U3789 (N_3789,N_1811,N_1359);
nor U3790 (N_3790,N_163,N_599);
or U3791 (N_3791,N_1512,N_270);
or U3792 (N_3792,N_956,N_211);
nand U3793 (N_3793,N_134,N_595);
and U3794 (N_3794,N_693,N_778);
or U3795 (N_3795,N_487,N_603);
nand U3796 (N_3796,N_1489,N_1730);
nand U3797 (N_3797,N_157,N_1160);
or U3798 (N_3798,N_581,N_585);
and U3799 (N_3799,N_1453,N_293);
nand U3800 (N_3800,N_120,N_630);
and U3801 (N_3801,N_421,N_478);
nor U3802 (N_3802,N_618,N_270);
nor U3803 (N_3803,N_1702,N_727);
and U3804 (N_3804,N_1209,N_121);
nor U3805 (N_3805,N_331,N_1893);
nor U3806 (N_3806,N_575,N_1532);
xnor U3807 (N_3807,N_684,N_1950);
or U3808 (N_3808,N_625,N_1016);
and U3809 (N_3809,N_1394,N_1043);
nor U3810 (N_3810,N_1545,N_1511);
and U3811 (N_3811,N_1932,N_537);
or U3812 (N_3812,N_477,N_1580);
nor U3813 (N_3813,N_1658,N_1499);
and U3814 (N_3814,N_194,N_554);
or U3815 (N_3815,N_745,N_282);
and U3816 (N_3816,N_637,N_1334);
or U3817 (N_3817,N_760,N_1484);
or U3818 (N_3818,N_764,N_33);
and U3819 (N_3819,N_718,N_90);
or U3820 (N_3820,N_1794,N_1815);
or U3821 (N_3821,N_463,N_1864);
nand U3822 (N_3822,N_1962,N_537);
nand U3823 (N_3823,N_1044,N_130);
and U3824 (N_3824,N_1154,N_1832);
or U3825 (N_3825,N_1353,N_1263);
nand U3826 (N_3826,N_1692,N_1126);
nor U3827 (N_3827,N_946,N_420);
and U3828 (N_3828,N_1009,N_416);
nor U3829 (N_3829,N_1856,N_1872);
nand U3830 (N_3830,N_880,N_1403);
or U3831 (N_3831,N_801,N_1464);
and U3832 (N_3832,N_1321,N_1367);
nor U3833 (N_3833,N_1573,N_1);
and U3834 (N_3834,N_1101,N_534);
and U3835 (N_3835,N_742,N_782);
or U3836 (N_3836,N_1746,N_1481);
and U3837 (N_3837,N_1443,N_641);
and U3838 (N_3838,N_1533,N_1209);
nand U3839 (N_3839,N_629,N_1206);
nand U3840 (N_3840,N_878,N_1196);
and U3841 (N_3841,N_1736,N_1927);
and U3842 (N_3842,N_1081,N_132);
nor U3843 (N_3843,N_967,N_440);
and U3844 (N_3844,N_1941,N_1356);
and U3845 (N_3845,N_271,N_516);
nor U3846 (N_3846,N_278,N_1068);
nor U3847 (N_3847,N_463,N_1097);
and U3848 (N_3848,N_1132,N_1337);
or U3849 (N_3849,N_328,N_769);
and U3850 (N_3850,N_1495,N_797);
nor U3851 (N_3851,N_1566,N_1593);
nor U3852 (N_3852,N_446,N_1104);
nor U3853 (N_3853,N_701,N_156);
and U3854 (N_3854,N_163,N_1700);
and U3855 (N_3855,N_539,N_1259);
and U3856 (N_3856,N_1422,N_538);
nor U3857 (N_3857,N_1190,N_1402);
and U3858 (N_3858,N_926,N_820);
nand U3859 (N_3859,N_1292,N_1908);
nor U3860 (N_3860,N_1090,N_298);
and U3861 (N_3861,N_415,N_568);
xor U3862 (N_3862,N_251,N_1754);
or U3863 (N_3863,N_662,N_391);
nand U3864 (N_3864,N_428,N_137);
and U3865 (N_3865,N_1073,N_1117);
nor U3866 (N_3866,N_321,N_184);
and U3867 (N_3867,N_488,N_1408);
or U3868 (N_3868,N_313,N_1889);
and U3869 (N_3869,N_442,N_1025);
nor U3870 (N_3870,N_130,N_79);
nor U3871 (N_3871,N_1002,N_1896);
and U3872 (N_3872,N_121,N_1719);
nor U3873 (N_3873,N_1898,N_1458);
nor U3874 (N_3874,N_1303,N_700);
nor U3875 (N_3875,N_1961,N_727);
nor U3876 (N_3876,N_454,N_1977);
nand U3877 (N_3877,N_1594,N_724);
nor U3878 (N_3878,N_937,N_688);
nand U3879 (N_3879,N_269,N_520);
and U3880 (N_3880,N_571,N_224);
and U3881 (N_3881,N_1328,N_1773);
nand U3882 (N_3882,N_681,N_13);
and U3883 (N_3883,N_518,N_1152);
or U3884 (N_3884,N_524,N_1110);
nor U3885 (N_3885,N_1276,N_301);
and U3886 (N_3886,N_477,N_1813);
or U3887 (N_3887,N_1698,N_1928);
nor U3888 (N_3888,N_1637,N_618);
and U3889 (N_3889,N_1680,N_549);
nor U3890 (N_3890,N_1830,N_274);
and U3891 (N_3891,N_20,N_1807);
or U3892 (N_3892,N_295,N_2);
or U3893 (N_3893,N_1307,N_420);
nand U3894 (N_3894,N_856,N_1101);
or U3895 (N_3895,N_1924,N_1220);
or U3896 (N_3896,N_1326,N_1521);
and U3897 (N_3897,N_1545,N_1567);
nor U3898 (N_3898,N_1290,N_328);
and U3899 (N_3899,N_466,N_1596);
nor U3900 (N_3900,N_176,N_302);
nand U3901 (N_3901,N_882,N_309);
nand U3902 (N_3902,N_1580,N_1995);
and U3903 (N_3903,N_1155,N_21);
nand U3904 (N_3904,N_1210,N_1660);
nor U3905 (N_3905,N_1807,N_1999);
and U3906 (N_3906,N_1263,N_189);
nand U3907 (N_3907,N_996,N_1711);
nand U3908 (N_3908,N_894,N_1303);
and U3909 (N_3909,N_14,N_182);
nand U3910 (N_3910,N_1756,N_1961);
nor U3911 (N_3911,N_1045,N_1694);
or U3912 (N_3912,N_87,N_1166);
nor U3913 (N_3913,N_1029,N_1824);
nor U3914 (N_3914,N_1081,N_772);
nand U3915 (N_3915,N_662,N_1845);
nand U3916 (N_3916,N_587,N_3);
or U3917 (N_3917,N_539,N_908);
or U3918 (N_3918,N_1912,N_812);
or U3919 (N_3919,N_1324,N_241);
or U3920 (N_3920,N_1207,N_1423);
and U3921 (N_3921,N_1964,N_747);
nand U3922 (N_3922,N_507,N_769);
nand U3923 (N_3923,N_982,N_953);
nand U3924 (N_3924,N_1142,N_543);
nand U3925 (N_3925,N_430,N_1454);
and U3926 (N_3926,N_516,N_1366);
nand U3927 (N_3927,N_929,N_1755);
nor U3928 (N_3928,N_1275,N_1598);
nand U3929 (N_3929,N_1715,N_1371);
xnor U3930 (N_3930,N_1733,N_1636);
and U3931 (N_3931,N_1532,N_197);
nor U3932 (N_3932,N_1914,N_858);
and U3933 (N_3933,N_1676,N_1244);
and U3934 (N_3934,N_1627,N_226);
nor U3935 (N_3935,N_1979,N_1512);
nand U3936 (N_3936,N_1893,N_1503);
xnor U3937 (N_3937,N_1149,N_107);
or U3938 (N_3938,N_216,N_1029);
and U3939 (N_3939,N_1921,N_1747);
nand U3940 (N_3940,N_59,N_881);
nand U3941 (N_3941,N_430,N_729);
or U3942 (N_3942,N_1656,N_631);
and U3943 (N_3943,N_1823,N_12);
nor U3944 (N_3944,N_1696,N_1565);
or U3945 (N_3945,N_1453,N_1880);
and U3946 (N_3946,N_1954,N_844);
nor U3947 (N_3947,N_121,N_919);
or U3948 (N_3948,N_498,N_1995);
or U3949 (N_3949,N_42,N_1664);
nand U3950 (N_3950,N_1840,N_648);
or U3951 (N_3951,N_1366,N_1852);
and U3952 (N_3952,N_898,N_1256);
and U3953 (N_3953,N_182,N_321);
nor U3954 (N_3954,N_409,N_72);
nand U3955 (N_3955,N_458,N_1886);
nor U3956 (N_3956,N_44,N_613);
or U3957 (N_3957,N_61,N_1302);
and U3958 (N_3958,N_904,N_376);
nor U3959 (N_3959,N_1490,N_1820);
or U3960 (N_3960,N_215,N_523);
nand U3961 (N_3961,N_288,N_1652);
or U3962 (N_3962,N_1759,N_1827);
or U3963 (N_3963,N_1522,N_1868);
or U3964 (N_3964,N_1987,N_1813);
or U3965 (N_3965,N_1920,N_430);
nor U3966 (N_3966,N_734,N_1638);
nor U3967 (N_3967,N_338,N_224);
nor U3968 (N_3968,N_1872,N_1626);
nor U3969 (N_3969,N_143,N_1493);
nand U3970 (N_3970,N_376,N_8);
and U3971 (N_3971,N_563,N_1393);
nor U3972 (N_3972,N_14,N_87);
and U3973 (N_3973,N_1744,N_385);
nor U3974 (N_3974,N_1541,N_1619);
nor U3975 (N_3975,N_602,N_921);
nand U3976 (N_3976,N_1420,N_186);
or U3977 (N_3977,N_957,N_136);
or U3978 (N_3978,N_400,N_782);
and U3979 (N_3979,N_103,N_981);
nand U3980 (N_3980,N_262,N_1167);
and U3981 (N_3981,N_1593,N_1416);
nor U3982 (N_3982,N_944,N_374);
or U3983 (N_3983,N_230,N_72);
and U3984 (N_3984,N_603,N_1682);
nand U3985 (N_3985,N_863,N_1438);
or U3986 (N_3986,N_869,N_820);
nor U3987 (N_3987,N_312,N_1256);
and U3988 (N_3988,N_1268,N_1550);
nand U3989 (N_3989,N_1208,N_1247);
and U3990 (N_3990,N_979,N_1781);
nor U3991 (N_3991,N_512,N_1362);
or U3992 (N_3992,N_714,N_661);
nand U3993 (N_3993,N_876,N_191);
or U3994 (N_3994,N_5,N_1332);
nor U3995 (N_3995,N_1983,N_660);
nor U3996 (N_3996,N_287,N_1411);
nor U3997 (N_3997,N_1367,N_1482);
nor U3998 (N_3998,N_792,N_598);
and U3999 (N_3999,N_1923,N_1979);
and U4000 (N_4000,N_2396,N_3172);
nor U4001 (N_4001,N_3984,N_3994);
nor U4002 (N_4002,N_3910,N_3461);
or U4003 (N_4003,N_2470,N_2581);
and U4004 (N_4004,N_2656,N_2799);
or U4005 (N_4005,N_2196,N_3249);
nor U4006 (N_4006,N_3872,N_2640);
and U4007 (N_4007,N_2797,N_2791);
nor U4008 (N_4008,N_3733,N_3008);
nand U4009 (N_4009,N_3606,N_3478);
and U4010 (N_4010,N_2431,N_3218);
nand U4011 (N_4011,N_3529,N_2503);
and U4012 (N_4012,N_3625,N_2966);
and U4013 (N_4013,N_2343,N_3770);
or U4014 (N_4014,N_2864,N_3064);
nand U4015 (N_4015,N_3438,N_3221);
and U4016 (N_4016,N_2734,N_2949);
or U4017 (N_4017,N_2385,N_2993);
nand U4018 (N_4018,N_2555,N_3775);
and U4019 (N_4019,N_3947,N_3630);
nor U4020 (N_4020,N_2435,N_3569);
nor U4021 (N_4021,N_2001,N_2533);
nor U4022 (N_4022,N_3639,N_3035);
nand U4023 (N_4023,N_3016,N_3869);
and U4024 (N_4024,N_2678,N_2342);
nand U4025 (N_4025,N_2378,N_3112);
nand U4026 (N_4026,N_2861,N_3978);
or U4027 (N_4027,N_2724,N_2243);
nor U4028 (N_4028,N_2605,N_3295);
nor U4029 (N_4029,N_2440,N_3620);
nor U4030 (N_4030,N_2651,N_2843);
nand U4031 (N_4031,N_3245,N_3051);
nand U4032 (N_4032,N_2401,N_2422);
and U4033 (N_4033,N_3576,N_3931);
nor U4034 (N_4034,N_3126,N_3704);
nand U4035 (N_4035,N_3017,N_2505);
nor U4036 (N_4036,N_3073,N_3122);
and U4037 (N_4037,N_3673,N_3379);
nor U4038 (N_4038,N_3259,N_3214);
nand U4039 (N_4039,N_2455,N_2982);
nor U4040 (N_4040,N_2082,N_2271);
or U4041 (N_4041,N_3099,N_3604);
and U4042 (N_4042,N_2839,N_3049);
nand U4043 (N_4043,N_2663,N_2523);
nand U4044 (N_4044,N_2316,N_2967);
nand U4045 (N_4045,N_3347,N_2235);
nor U4046 (N_4046,N_2331,N_2357);
and U4047 (N_4047,N_3414,N_3916);
nand U4048 (N_4048,N_3061,N_3581);
and U4049 (N_4049,N_2450,N_2252);
nand U4050 (N_4050,N_3136,N_2836);
nor U4051 (N_4051,N_3642,N_3325);
and U4052 (N_4052,N_2356,N_2705);
nor U4053 (N_4053,N_2617,N_2475);
nand U4054 (N_4054,N_2746,N_3742);
nor U4055 (N_4055,N_2382,N_2841);
or U4056 (N_4056,N_2425,N_2075);
nor U4057 (N_4057,N_3324,N_3083);
or U4058 (N_4058,N_2491,N_3210);
and U4059 (N_4059,N_3441,N_2832);
and U4060 (N_4060,N_2265,N_3213);
nor U4061 (N_4061,N_3101,N_3434);
or U4062 (N_4062,N_3993,N_2124);
or U4063 (N_4063,N_2907,N_2403);
or U4064 (N_4064,N_3314,N_2155);
and U4065 (N_4065,N_2901,N_2911);
xor U4066 (N_4066,N_2738,N_3148);
nor U4067 (N_4067,N_3048,N_2681);
or U4068 (N_4068,N_3619,N_3496);
or U4069 (N_4069,N_3244,N_3431);
or U4070 (N_4070,N_2960,N_2969);
or U4071 (N_4071,N_2943,N_2349);
and U4072 (N_4072,N_3151,N_3740);
nand U4073 (N_4073,N_2257,N_2583);
nor U4074 (N_4074,N_2168,N_3066);
or U4075 (N_4075,N_2115,N_3342);
or U4076 (N_4076,N_3175,N_3656);
nor U4077 (N_4077,N_2245,N_2906);
nand U4078 (N_4078,N_2748,N_2856);
or U4079 (N_4079,N_3404,N_3076);
or U4080 (N_4080,N_3121,N_3201);
and U4081 (N_4081,N_3095,N_2441);
nor U4082 (N_4082,N_2613,N_2545);
or U4083 (N_4083,N_3447,N_2217);
and U4084 (N_4084,N_3472,N_2180);
and U4085 (N_4085,N_3290,N_2892);
and U4086 (N_4086,N_3802,N_2706);
or U4087 (N_4087,N_3147,N_2273);
nand U4088 (N_4088,N_3729,N_3392);
and U4089 (N_4089,N_2573,N_2910);
nand U4090 (N_4090,N_2379,N_3373);
and U4091 (N_4091,N_3158,N_2080);
nor U4092 (N_4092,N_3155,N_2372);
or U4093 (N_4093,N_3231,N_3788);
and U4094 (N_4094,N_3777,N_2567);
and U4095 (N_4095,N_2940,N_2668);
and U4096 (N_4096,N_2103,N_3394);
nand U4097 (N_4097,N_3592,N_3306);
and U4098 (N_4098,N_2049,N_2091);
and U4099 (N_4099,N_3677,N_2473);
and U4100 (N_4100,N_2823,N_3469);
nor U4101 (N_4101,N_2310,N_2069);
and U4102 (N_4102,N_3475,N_2042);
and U4103 (N_4103,N_3498,N_3763);
nand U4104 (N_4104,N_3250,N_3806);
or U4105 (N_4105,N_3833,N_2768);
nor U4106 (N_4106,N_3145,N_2603);
nand U4107 (N_4107,N_3545,N_3730);
nand U4108 (N_4108,N_2635,N_3856);
and U4109 (N_4109,N_2673,N_3281);
and U4110 (N_4110,N_2057,N_2500);
or U4111 (N_4111,N_3071,N_3480);
and U4112 (N_4112,N_2474,N_2804);
nand U4113 (N_4113,N_3299,N_3355);
nor U4114 (N_4114,N_3786,N_2903);
and U4115 (N_4115,N_2661,N_2436);
and U4116 (N_4116,N_2953,N_3990);
nand U4117 (N_4117,N_2991,N_3334);
or U4118 (N_4118,N_2530,N_2751);
nand U4119 (N_4119,N_3242,N_3425);
or U4120 (N_4120,N_2323,N_3018);
or U4121 (N_4121,N_3042,N_3901);
nand U4122 (N_4122,N_2383,N_2974);
and U4123 (N_4123,N_3583,N_3188);
nor U4124 (N_4124,N_2809,N_3486);
nor U4125 (N_4125,N_2822,N_2896);
nor U4126 (N_4126,N_2007,N_2850);
nor U4127 (N_4127,N_3701,N_3227);
nand U4128 (N_4128,N_3019,N_2132);
and U4129 (N_4129,N_3060,N_3055);
and U4130 (N_4130,N_3900,N_2044);
nor U4131 (N_4131,N_3636,N_3944);
nor U4132 (N_4132,N_3430,N_3720);
or U4133 (N_4133,N_2774,N_3671);
or U4134 (N_4134,N_3068,N_2464);
and U4135 (N_4135,N_3321,N_2418);
nor U4136 (N_4136,N_2954,N_3455);
nand U4137 (N_4137,N_3666,N_2112);
nand U4138 (N_4138,N_3700,N_3270);
nand U4139 (N_4139,N_2386,N_2912);
or U4140 (N_4140,N_2979,N_2339);
nand U4141 (N_4141,N_2831,N_3542);
and U4142 (N_4142,N_2185,N_3089);
nor U4143 (N_4143,N_3971,N_3141);
nand U4144 (N_4144,N_2139,N_3118);
or U4145 (N_4145,N_2835,N_2690);
and U4146 (N_4146,N_3252,N_2032);
nand U4147 (N_4147,N_2818,N_2306);
and U4148 (N_4148,N_2411,N_2058);
or U4149 (N_4149,N_2702,N_2789);
nor U4150 (N_4150,N_2990,N_2758);
or U4151 (N_4151,N_3494,N_2506);
nand U4152 (N_4152,N_2716,N_2658);
or U4153 (N_4153,N_2744,N_3813);
nor U4154 (N_4154,N_3522,N_3138);
or U4155 (N_4155,N_3832,N_3587);
and U4156 (N_4156,N_3100,N_2236);
nand U4157 (N_4157,N_2695,N_2041);
nand U4158 (N_4158,N_3409,N_3877);
and U4159 (N_4159,N_3109,N_2096);
xnor U4160 (N_4160,N_3376,N_2522);
or U4161 (N_4161,N_3865,N_3711);
nand U4162 (N_4162,N_2565,N_2520);
or U4163 (N_4163,N_2294,N_2468);
nand U4164 (N_4164,N_2723,N_3760);
nor U4165 (N_4165,N_2694,N_3951);
nand U4166 (N_4166,N_2607,N_3313);
and U4167 (N_4167,N_2360,N_2097);
nor U4168 (N_4168,N_2146,N_3670);
and U4169 (N_4169,N_3652,N_3897);
and U4170 (N_4170,N_3146,N_3505);
or U4171 (N_4171,N_3021,N_3364);
and U4172 (N_4172,N_3115,N_3489);
nand U4173 (N_4173,N_3692,N_2055);
nor U4174 (N_4174,N_2697,N_3600);
nand U4175 (N_4175,N_2699,N_2169);
and U4176 (N_4176,N_3482,N_3599);
nand U4177 (N_4177,N_3086,N_2054);
nor U4178 (N_4178,N_2215,N_3933);
and U4179 (N_4179,N_3950,N_3908);
nor U4180 (N_4180,N_2384,N_2325);
or U4181 (N_4181,N_3593,N_3220);
nand U4182 (N_4182,N_2721,N_2736);
or U4183 (N_4183,N_2003,N_3710);
nand U4184 (N_4184,N_3568,N_2917);
and U4185 (N_4185,N_2191,N_3398);
or U4186 (N_4186,N_2704,N_2345);
nor U4187 (N_4187,N_2233,N_2394);
nor U4188 (N_4188,N_2486,N_2085);
and U4189 (N_4189,N_2996,N_3193);
nor U4190 (N_4190,N_3075,N_2921);
nand U4191 (N_4191,N_3986,N_3714);
nand U4192 (N_4192,N_2076,N_3517);
nor U4193 (N_4193,N_3429,N_3030);
or U4194 (N_4194,N_2609,N_3418);
and U4195 (N_4195,N_2687,N_2072);
nand U4196 (N_4196,N_2959,N_3928);
and U4197 (N_4197,N_2117,N_2632);
nor U4198 (N_4198,N_3597,N_3144);
or U4199 (N_4199,N_3663,N_2052);
or U4200 (N_4200,N_2493,N_3911);
nand U4201 (N_4201,N_3331,N_3256);
nor U4202 (N_4202,N_2575,N_2251);
or U4203 (N_4203,N_2941,N_2188);
xnor U4204 (N_4204,N_2918,N_3456);
and U4205 (N_4205,N_3874,N_3436);
nor U4206 (N_4206,N_2140,N_3919);
nor U4207 (N_4207,N_3561,N_2011);
and U4208 (N_4208,N_2534,N_2402);
xor U4209 (N_4209,N_2249,N_3724);
nor U4210 (N_4210,N_3407,N_2871);
and U4211 (N_4211,N_3871,N_3989);
and U4212 (N_4212,N_2869,N_2919);
and U4213 (N_4213,N_2174,N_3185);
and U4214 (N_4214,N_3672,N_3820);
nand U4215 (N_4215,N_3289,N_2181);
nand U4216 (N_4216,N_2879,N_2526);
and U4217 (N_4217,N_2867,N_3209);
nand U4218 (N_4218,N_3938,N_3857);
nand U4219 (N_4219,N_2037,N_3696);
nand U4220 (N_4220,N_2754,N_2773);
or U4221 (N_4221,N_3124,N_2264);
nor U4222 (N_4222,N_2584,N_2494);
and U4223 (N_4223,N_2204,N_2988);
and U4224 (N_4224,N_3834,N_2028);
nor U4225 (N_4225,N_2457,N_2580);
or U4226 (N_4226,N_3782,N_2176);
nand U4227 (N_4227,N_2490,N_2665);
nand U4228 (N_4228,N_3552,N_2570);
nor U4229 (N_4229,N_3559,N_3632);
or U4230 (N_4230,N_3098,N_2100);
or U4231 (N_4231,N_3554,N_3003);
nand U4232 (N_4232,N_3844,N_3891);
and U4233 (N_4233,N_3241,N_3359);
or U4234 (N_4234,N_2269,N_3570);
or U4235 (N_4235,N_2387,N_3257);
nor U4236 (N_4236,N_2410,N_2838);
and U4237 (N_4237,N_2718,N_3847);
nor U4238 (N_4238,N_2680,N_2105);
and U4239 (N_4239,N_3421,N_3683);
nor U4240 (N_4240,N_2853,N_3007);
and U4241 (N_4241,N_2891,N_3512);
nand U4242 (N_4242,N_2398,N_3163);
and U4243 (N_4243,N_3131,N_3387);
nor U4244 (N_4244,N_2266,N_3992);
or U4245 (N_4245,N_3894,N_3825);
or U4246 (N_4246,N_2281,N_2501);
nand U4247 (N_4247,N_2925,N_3205);
and U4248 (N_4248,N_2932,N_3647);
nand U4249 (N_4249,N_2980,N_3174);
and U4250 (N_4250,N_2309,N_2419);
nor U4251 (N_4251,N_2299,N_3337);
nor U4252 (N_4252,N_2391,N_3527);
or U4253 (N_4253,N_3664,N_2674);
nand U4254 (N_4254,N_2444,N_2201);
and U4255 (N_4255,N_3932,N_2604);
or U4256 (N_4256,N_2556,N_2561);
nor U4257 (N_4257,N_3826,N_3859);
and U4258 (N_4258,N_3178,N_2312);
or U4259 (N_4259,N_3699,N_3694);
nor U4260 (N_4260,N_3279,N_2035);
or U4261 (N_4261,N_2027,N_3917);
nor U4262 (N_4262,N_2578,N_2562);
or U4263 (N_4263,N_2779,N_3767);
and U4264 (N_4264,N_2992,N_2554);
nand U4265 (N_4265,N_2307,N_3814);
and U4266 (N_4266,N_3792,N_3203);
nand U4267 (N_4267,N_3190,N_2270);
or U4268 (N_4268,N_3236,N_2770);
or U4269 (N_4269,N_2361,N_3794);
nand U4270 (N_4270,N_3892,N_2890);
or U4271 (N_4271,N_2446,N_2899);
and U4272 (N_4272,N_2909,N_2764);
nor U4273 (N_4273,N_3180,N_3899);
or U4274 (N_4274,N_3361,N_3765);
nand U4275 (N_4275,N_2225,N_3646);
nand U4276 (N_4276,N_3156,N_2676);
nand U4277 (N_4277,N_2727,N_2336);
nor U4278 (N_4278,N_3548,N_3854);
or U4279 (N_4279,N_2825,N_2412);
nor U4280 (N_4280,N_3260,N_2467);
or U4281 (N_4281,N_2998,N_3332);
nor U4282 (N_4282,N_3949,N_2184);
or U4283 (N_4283,N_3852,N_2178);
and U4284 (N_4284,N_2606,N_2487);
and U4285 (N_4285,N_3886,N_3798);
and U4286 (N_4286,N_2111,N_3764);
or U4287 (N_4287,N_3362,N_2426);
and U4288 (N_4288,N_3644,N_2034);
and U4289 (N_4289,N_2078,N_3963);
and U4290 (N_4290,N_3015,N_2795);
and U4291 (N_4291,N_3608,N_3996);
or U4292 (N_4292,N_3152,N_2152);
nand U4293 (N_4293,N_3222,N_2395);
xor U4294 (N_4294,N_3779,N_3878);
nand U4295 (N_4295,N_3127,N_3336);
nand U4296 (N_4296,N_2375,N_2870);
nor U4297 (N_4297,N_3232,N_3102);
nand U4298 (N_4298,N_3598,N_2594);
or U4299 (N_4299,N_3735,N_3166);
and U4300 (N_4300,N_2187,N_2848);
and U4301 (N_4301,N_2951,N_3219);
and U4302 (N_4302,N_2905,N_2755);
and U4303 (N_4303,N_2893,N_3631);
nor U4304 (N_4304,N_3437,N_3459);
nand U4305 (N_4305,N_3053,N_3006);
nand U4306 (N_4306,N_2489,N_2136);
nand U4307 (N_4307,N_3697,N_2707);
nor U4308 (N_4308,N_2945,N_2449);
nor U4309 (N_4309,N_3339,N_3153);
nand U4310 (N_4310,N_2023,N_2715);
nor U4311 (N_4311,N_2195,N_2756);
nand U4312 (N_4312,N_2127,N_3493);
nor U4313 (N_4313,N_3465,N_2552);
or U4314 (N_4314,N_2710,N_2485);
and U4315 (N_4315,N_3104,N_3474);
nand U4316 (N_4316,N_2591,N_2048);
or U4317 (N_4317,N_3516,N_2897);
nor U4318 (N_4318,N_3553,N_3285);
and U4319 (N_4319,N_2840,N_3893);
and U4320 (N_4320,N_3640,N_2456);
nand U4321 (N_4321,N_2043,N_3964);
nand U4322 (N_4322,N_3778,N_2047);
nor U4323 (N_4323,N_3261,N_3371);
and U4324 (N_4324,N_2083,N_2301);
nor U4325 (N_4325,N_3424,N_3695);
and U4326 (N_4326,N_2737,N_2952);
nand U4327 (N_4327,N_3275,N_2863);
and U4328 (N_4328,N_3405,N_2589);
nand U4329 (N_4329,N_3399,N_3889);
and U4330 (N_4330,N_2826,N_3199);
or U4331 (N_4331,N_2691,N_2972);
and U4332 (N_4332,N_2778,N_3582);
and U4333 (N_4333,N_2511,N_3246);
or U4334 (N_4334,N_2753,N_2504);
or U4335 (N_4335,N_2194,N_2421);
and U4336 (N_4336,N_2660,N_2865);
and U4337 (N_4337,N_2794,N_2013);
nand U4338 (N_4338,N_2305,N_3584);
and U4339 (N_4339,N_2559,N_2571);
nand U4340 (N_4340,N_3797,N_3954);
and U4341 (N_4341,N_3268,N_2373);
nand U4342 (N_4342,N_2209,N_3579);
or U4343 (N_4343,N_3707,N_2370);
nand U4344 (N_4344,N_2439,N_2012);
or U4345 (N_4345,N_2389,N_2407);
nor U4346 (N_4346,N_2612,N_2783);
or U4347 (N_4347,N_2232,N_3351);
and U4348 (N_4348,N_2937,N_2645);
nor U4349 (N_4349,N_2040,N_2471);
nand U4350 (N_4350,N_2685,N_2302);
or U4351 (N_4351,N_3052,N_2569);
nor U4352 (N_4352,N_2062,N_3948);
nor U4353 (N_4353,N_2693,N_2700);
or U4354 (N_4354,N_2004,N_3687);
and U4355 (N_4355,N_3036,N_2133);
and U4356 (N_4356,N_2518,N_3654);
and U4357 (N_4357,N_2484,N_3966);
or U4358 (N_4358,N_2247,N_3801);
nor U4359 (N_4359,N_3759,N_3848);
nand U4360 (N_4360,N_2689,N_2543);
or U4361 (N_4361,N_2406,N_3041);
nor U4362 (N_4362,N_3410,N_3396);
or U4363 (N_4363,N_3501,N_3223);
nand U4364 (N_4364,N_2759,N_3183);
nand U4365 (N_4365,N_3452,N_2800);
nand U4366 (N_4366,N_3416,N_3123);
nand U4367 (N_4367,N_2197,N_2122);
nand U4368 (N_4368,N_3614,N_2495);
nand U4369 (N_4369,N_3385,N_2397);
nor U4370 (N_4370,N_2855,N_3291);
and U4371 (N_4371,N_3097,N_3078);
or U4372 (N_4372,N_2303,N_2156);
nand U4373 (N_4373,N_2742,N_3173);
nor U4374 (N_4374,N_2983,N_2173);
and U4375 (N_4375,N_2120,N_3084);
nand U4376 (N_4376,N_2999,N_2478);
or U4377 (N_4377,N_3182,N_2255);
nor U4378 (N_4378,N_3574,N_2296);
nand U4379 (N_4379,N_2150,N_3386);
or U4380 (N_4380,N_3217,N_2365);
and U4381 (N_4381,N_2984,N_3525);
nand U4382 (N_4382,N_2792,N_2297);
or U4383 (N_4383,N_2994,N_3590);
nor U4384 (N_4384,N_2527,N_2145);
nand U4385 (N_4385,N_3335,N_2817);
nand U4386 (N_4386,N_3762,N_2788);
and U4387 (N_4387,N_3974,N_2333);
nand U4388 (N_4388,N_2894,N_2280);
nor U4389 (N_4389,N_2885,N_2611);
or U4390 (N_4390,N_2948,N_2106);
and U4391 (N_4391,N_2913,N_2017);
and U4392 (N_4392,N_3411,N_3358);
nor U4393 (N_4393,N_3698,N_3315);
and U4394 (N_4394,N_3812,N_2638);
or U4395 (N_4395,N_2094,N_3069);
and U4396 (N_4396,N_3717,N_2392);
or U4397 (N_4397,N_2199,N_3116);
and U4398 (N_4398,N_3085,N_3863);
and U4399 (N_4399,N_2557,N_3939);
or U4400 (N_4400,N_3432,N_3688);
or U4401 (N_4401,N_2098,N_2986);
nand U4402 (N_4402,N_3164,N_2517);
nand U4403 (N_4403,N_2944,N_2560);
and U4404 (N_4404,N_2733,N_2417);
or U4405 (N_4405,N_3689,N_2061);
and U4406 (N_4406,N_3945,N_3354);
nor U4407 (N_4407,N_3179,N_2653);
and U4408 (N_4408,N_2498,N_3028);
nor U4409 (N_4409,N_3823,N_3288);
xor U4410 (N_4410,N_3239,N_3623);
nand U4411 (N_4411,N_2851,N_3506);
nand U4412 (N_4412,N_2977,N_3756);
and U4413 (N_4413,N_3237,N_3918);
nand U4414 (N_4414,N_3079,N_3790);
nor U4415 (N_4415,N_2344,N_2241);
xnor U4416 (N_4416,N_2368,N_2338);
and U4417 (N_4417,N_2424,N_2670);
nand U4418 (N_4418,N_2981,N_2908);
nor U4419 (N_4419,N_2588,N_2364);
nor U4420 (N_4420,N_3967,N_2709);
nand U4421 (N_4421,N_3423,N_3566);
nor U4422 (N_4422,N_3556,N_2847);
and U4423 (N_4423,N_3960,N_2542);
and U4424 (N_4424,N_3384,N_2071);
nor U4425 (N_4425,N_3535,N_2837);
nand U4426 (N_4426,N_2268,N_3278);
or U4427 (N_4427,N_3780,N_3463);
or U4428 (N_4428,N_2428,N_2144);
nand U4429 (N_4429,N_3845,N_3067);
nand U4430 (N_4430,N_2123,N_2975);
nand U4431 (N_4431,N_3617,N_3880);
nand U4432 (N_4432,N_3749,N_2790);
nor U4433 (N_4433,N_2546,N_2730);
or U4434 (N_4434,N_3715,N_2359);
nand U4435 (N_4435,N_3422,N_3171);
or U4436 (N_4436,N_2803,N_2363);
or U4437 (N_4437,N_3706,N_2154);
and U4438 (N_4438,N_3057,N_2317);
nor U4439 (N_4439,N_3748,N_3374);
nand U4440 (N_4440,N_3024,N_2240);
nor U4441 (N_4441,N_3923,N_3280);
nor U4442 (N_4442,N_3026,N_3616);
or U4443 (N_4443,N_3370,N_3282);
nand U4444 (N_4444,N_2291,N_2806);
nand U4445 (N_4445,N_3613,N_3649);
nor U4446 (N_4446,N_3703,N_2246);
nand U4447 (N_4447,N_3283,N_3137);
or U4448 (N_4448,N_2973,N_2347);
or U4449 (N_4449,N_2447,N_2568);
and U4450 (N_4450,N_3681,N_2722);
or U4451 (N_4451,N_3500,N_2295);
or U4452 (N_4452,N_3995,N_3739);
nand U4453 (N_4453,N_2572,N_2340);
nor U4454 (N_4454,N_2477,N_3540);
or U4455 (N_4455,N_3113,N_2978);
nor U4456 (N_4456,N_3734,N_3233);
nand U4457 (N_4457,N_2880,N_3920);
and U4458 (N_4458,N_3367,N_2161);
xnor U4459 (N_4459,N_3310,N_3108);
or U4460 (N_4460,N_2502,N_3816);
nand U4461 (N_4461,N_2212,N_2362);
or U4462 (N_4462,N_3867,N_2077);
or U4463 (N_4463,N_3303,N_3010);
or U4464 (N_4464,N_2579,N_3272);
or U4465 (N_4465,N_2278,N_2947);
nand U4466 (N_4466,N_3327,N_2203);
nor U4467 (N_4467,N_2207,N_2285);
nor U4468 (N_4468,N_3307,N_3976);
nand U4469 (N_4469,N_3473,N_2516);
or U4470 (N_4470,N_3541,N_3909);
or U4471 (N_4471,N_3316,N_3783);
or U4472 (N_4472,N_3955,N_2633);
nand U4473 (N_4473,N_2654,N_3032);
and U4474 (N_4474,N_2987,N_3921);
nor U4475 (N_4475,N_2740,N_3000);
nor U4476 (N_4476,N_3389,N_2816);
nand U4477 (N_4477,N_2961,N_3722);
or U4478 (N_4478,N_2766,N_3135);
nor U4479 (N_4479,N_2131,N_3718);
nand U4480 (N_4480,N_3194,N_2714);
and U4481 (N_4481,N_3157,N_2538);
or U4482 (N_4482,N_2015,N_3420);
nor U4483 (N_4483,N_3904,N_3412);
or U4484 (N_4484,N_2683,N_3345);
or U4485 (N_4485,N_2427,N_2314);
or U4486 (N_4486,N_3243,N_2808);
nand U4487 (N_4487,N_2210,N_3226);
or U4488 (N_4488,N_3882,N_3685);
and U4489 (N_4489,N_2731,N_2989);
or U4490 (N_4490,N_3139,N_3382);
and U4491 (N_4491,N_2084,N_3661);
nor U4492 (N_4492,N_3111,N_3216);
and U4493 (N_4493,N_2143,N_2846);
nor U4494 (N_4494,N_3723,N_2741);
nand U4495 (N_4495,N_3274,N_3002);
or U4496 (N_4496,N_3843,N_2262);
or U4497 (N_4497,N_3676,N_3023);
nand U4498 (N_4498,N_2067,N_3519);
and U4499 (N_4499,N_2128,N_3070);
xnor U4500 (N_4500,N_2786,N_3589);
nor U4501 (N_4501,N_3952,N_3497);
nor U4502 (N_4502,N_2942,N_2760);
xor U4503 (N_4503,N_3262,N_2289);
nand U4504 (N_4504,N_2448,N_2479);
nor U4505 (N_4505,N_3513,N_3150);
and U4506 (N_4506,N_3741,N_2443);
nand U4507 (N_4507,N_3269,N_2073);
and U4508 (N_4508,N_2587,N_3077);
nand U4509 (N_4509,N_3906,N_3328);
nor U4510 (N_4510,N_3523,N_3712);
and U4511 (N_4511,N_3815,N_3479);
and U4512 (N_4512,N_2798,N_3657);
nor U4513 (N_4513,N_3502,N_3413);
or U4514 (N_4514,N_3969,N_3839);
nand U4515 (N_4515,N_2682,N_3483);
and U4516 (N_4516,N_2657,N_2828);
or U4517 (N_4517,N_3453,N_2537);
or U4518 (N_4518,N_2713,N_2963);
or U4519 (N_4519,N_3490,N_2414);
xor U4520 (N_4520,N_3159,N_3440);
nor U4521 (N_4521,N_3368,N_3031);
nand U4522 (N_4522,N_2636,N_2824);
or U4523 (N_4523,N_2956,N_3716);
or U4524 (N_4524,N_2749,N_3014);
nor U4525 (N_4525,N_2274,N_2765);
nand U4526 (N_4526,N_2887,N_2283);
or U4527 (N_4527,N_2782,N_3961);
nand U4528 (N_4528,N_2922,N_2684);
nand U4529 (N_4529,N_3298,N_3302);
nor U4530 (N_4530,N_2099,N_2253);
nand U4531 (N_4531,N_2872,N_2433);
and U4532 (N_4532,N_2025,N_3853);
and U4533 (N_4533,N_2416,N_2728);
or U4534 (N_4534,N_3907,N_2182);
nand U4535 (N_4535,N_3215,N_2862);
nor U4536 (N_4536,N_3340,N_3129);
or U4537 (N_4537,N_3383,N_2540);
or U4538 (N_4538,N_3341,N_3959);
and U4539 (N_4539,N_3884,N_3817);
nor U4540 (N_4540,N_2171,N_2107);
nor U4541 (N_4541,N_3755,N_2022);
nand U4542 (N_4542,N_3503,N_3248);
or U4543 (N_4543,N_3093,N_3787);
nor U4544 (N_4544,N_2876,N_3726);
and U4545 (N_4545,N_3207,N_3705);
and U4546 (N_4546,N_3660,N_3356);
nor U4547 (N_4547,N_3862,N_3022);
nor U4548 (N_4548,N_2350,N_3725);
and U4549 (N_4549,N_2820,N_2703);
nor U4550 (N_4550,N_2224,N_2650);
and U4551 (N_4551,N_2686,N_2877);
and U4552 (N_4552,N_3133,N_3868);
and U4553 (N_4553,N_2219,N_2459);
and U4554 (N_4554,N_3758,N_3091);
or U4555 (N_4555,N_2964,N_2400);
or U4556 (N_4556,N_3251,N_2648);
and U4557 (N_4557,N_3444,N_2634);
or U4558 (N_4558,N_3271,N_3543);
and U4559 (N_4559,N_3477,N_2237);
or U4560 (N_4560,N_2159,N_3267);
and U4561 (N_4561,N_3595,N_3196);
or U4562 (N_4562,N_3047,N_3881);
nand U4563 (N_4563,N_3514,N_2926);
nor U4564 (N_4564,N_3352,N_2884);
nand U4565 (N_4565,N_2050,N_2192);
or U4566 (N_4566,N_3338,N_2810);
or U4567 (N_4567,N_2166,N_3732);
nor U4568 (N_4568,N_2873,N_2962);
or U4569 (N_4569,N_3883,N_2666);
or U4570 (N_4570,N_2104,N_3451);
and U4571 (N_4571,N_3835,N_2321);
or U4572 (N_4572,N_2776,N_3988);
nand U4573 (N_4573,N_3038,N_3276);
nor U4574 (N_4574,N_3629,N_3029);
nand U4575 (N_4575,N_2933,N_2177);
nor U4576 (N_4576,N_3333,N_3800);
nand U4577 (N_4577,N_2248,N_2558);
nand U4578 (N_4578,N_3846,N_3571);
and U4579 (N_4579,N_3012,N_3119);
and U4580 (N_4580,N_2202,N_3610);
nand U4581 (N_4581,N_2213,N_3309);
or U4582 (N_4582,N_2056,N_3528);
nor U4583 (N_4583,N_3641,N_3308);
and U4584 (N_4584,N_3184,N_2198);
nand U4585 (N_4585,N_3462,N_2881);
nand U4586 (N_4586,N_3090,N_2600);
nand U4587 (N_4587,N_2598,N_3011);
xnor U4588 (N_4588,N_3426,N_2318);
or U4589 (N_4589,N_2830,N_3074);
and U4590 (N_4590,N_2130,N_2777);
nand U4591 (N_4591,N_3557,N_2254);
nand U4592 (N_4592,N_3979,N_3958);
nand U4593 (N_4593,N_2514,N_3300);
nor U4594 (N_4594,N_3128,N_3743);
and U4595 (N_4595,N_2854,N_2329);
nand U4596 (N_4596,N_3981,N_3924);
nor U4597 (N_4597,N_3821,N_2172);
or U4598 (N_4598,N_3972,N_2539);
and U4599 (N_4599,N_3751,N_2320);
and U4600 (N_4600,N_2811,N_3349);
and U4601 (N_4601,N_3192,N_2618);
and U4602 (N_4602,N_3668,N_3005);
and U4603 (N_4603,N_3390,N_2258);
and U4604 (N_4604,N_3913,N_3264);
and U4605 (N_4605,N_2081,N_2927);
nor U4606 (N_4606,N_3962,N_3234);
nor U4607 (N_4607,N_2593,N_2087);
nand U4608 (N_4608,N_2528,N_3940);
and U4609 (N_4609,N_2644,N_2292);
nor U4610 (N_4610,N_2110,N_2590);
or U4611 (N_4611,N_2290,N_2550);
nand U4612 (N_4612,N_3789,N_2564);
and U4613 (N_4613,N_2955,N_3555);
or U4614 (N_4614,N_2672,N_2548);
nor U4615 (N_4615,N_2045,N_3140);
or U4616 (N_4616,N_3653,N_3605);
and U4617 (N_4617,N_3935,N_3896);
nand U4618 (N_4618,N_2874,N_2186);
nand U4619 (N_4619,N_3769,N_2698);
and U4620 (N_4620,N_3682,N_2965);
or U4621 (N_4621,N_3936,N_3082);
and U4622 (N_4622,N_3258,N_3296);
and U4623 (N_4623,N_2802,N_2513);
nor U4624 (N_4624,N_3615,N_2655);
nand U4625 (N_4625,N_3750,N_3346);
or U4626 (N_4626,N_3350,N_2335);
and U4627 (N_4627,N_2574,N_3905);
or U4628 (N_4628,N_2827,N_2646);
or U4629 (N_4629,N_2608,N_3160);
xor U4630 (N_4630,N_3925,N_2938);
and U4631 (N_4631,N_2857,N_3861);
nand U4632 (N_4632,N_3027,N_3902);
or U4633 (N_4633,N_2620,N_2630);
or U4634 (N_4634,N_2381,N_2793);
nor U4635 (N_4635,N_2669,N_3684);
or U4636 (N_4636,N_3621,N_2623);
or U4637 (N_4637,N_3344,N_3643);
or U4638 (N_4638,N_3065,N_2946);
or U4639 (N_4639,N_3433,N_3406);
and U4640 (N_4640,N_2355,N_2599);
and U4641 (N_4641,N_2348,N_3766);
nor U4642 (N_4642,N_3601,N_3809);
and U4643 (N_4643,N_3588,N_3212);
nand U4644 (N_4644,N_3637,N_3890);
nor U4645 (N_4645,N_3277,N_3402);
nand U4646 (N_4646,N_2529,N_3204);
or U4647 (N_4647,N_2208,N_2293);
and U4648 (N_4648,N_2627,N_2282);
nand U4649 (N_4649,N_3117,N_3973);
or U4650 (N_4650,N_2002,N_2234);
or U4651 (N_4651,N_3985,N_3922);
and U4652 (N_4652,N_2476,N_2374);
or U4653 (N_4653,N_2842,N_3435);
nor U4654 (N_4654,N_3197,N_2429);
nand U4655 (N_4655,N_3317,N_3879);
or U4656 (N_4656,N_3230,N_3403);
nor U4657 (N_4657,N_2442,N_2308);
and U4658 (N_4658,N_3004,N_3651);
and U4659 (N_4659,N_2934,N_3547);
nand U4660 (N_4660,N_3488,N_3120);
or U4661 (N_4661,N_2813,N_2059);
or U4662 (N_4662,N_2134,N_3521);
nand U4663 (N_4663,N_3575,N_3106);
nand U4664 (N_4664,N_3558,N_2735);
or U4665 (N_4665,N_2068,N_2997);
or U4666 (N_4666,N_3980,N_2807);
nand U4667 (N_4667,N_3975,N_3544);
nor U4668 (N_4668,N_2968,N_3533);
and U4669 (N_4669,N_3388,N_2093);
or U4670 (N_4670,N_2875,N_2995);
or U4671 (N_4671,N_2971,N_2719);
nor U4672 (N_4672,N_3591,N_2351);
or U4673 (N_4673,N_2629,N_2126);
or U4674 (N_4674,N_2931,N_2775);
nor U4675 (N_4675,N_3757,N_3791);
nand U4676 (N_4676,N_2463,N_3784);
and U4677 (N_4677,N_2129,N_3747);
and U4678 (N_4678,N_2566,N_2679);
nand U4679 (N_4679,N_2019,N_3808);
and U4680 (N_4680,N_3752,N_2860);
and U4681 (N_4681,N_3793,N_2160);
or U4682 (N_4682,N_2089,N_2162);
nor U4683 (N_4683,N_2183,N_2016);
nor U4684 (N_4684,N_2785,N_3287);
nand U4685 (N_4685,N_2510,N_2218);
nor U4686 (N_4686,N_3266,N_3567);
or U4687 (N_4687,N_3603,N_2267);
nand U4688 (N_4688,N_3058,N_2920);
or U4689 (N_4689,N_2157,N_2829);
and U4690 (N_4690,N_3796,N_3785);
and U4691 (N_4691,N_2353,N_3046);
and U4692 (N_4692,N_2415,N_2497);
or U4693 (N_4693,N_3648,N_3492);
or U4694 (N_4694,N_2677,N_3001);
nor U4695 (N_4695,N_2277,N_3162);
nand U4696 (N_4696,N_2063,N_3596);
nor U4697 (N_4697,N_3235,N_3546);
nand U4698 (N_4698,N_3130,N_2821);
and U4699 (N_4699,N_3467,N_3305);
and U4700 (N_4700,N_3737,N_3062);
and U4701 (N_4701,N_2720,N_2729);
nand U4702 (N_4702,N_3134,N_2915);
and U4703 (N_4703,N_3050,N_2211);
nand U4704 (N_4704,N_3025,N_3736);
and U4705 (N_4705,N_3365,N_2761);
or U4706 (N_4706,N_3611,N_2551);
or U4707 (N_4707,N_3840,N_3929);
nor U4708 (N_4708,N_2595,N_3536);
nand U4709 (N_4709,N_3464,N_2596);
nand U4710 (N_4710,N_2615,N_2408);
nand U4711 (N_4711,N_3563,N_3721);
nor U4712 (N_4712,N_2957,N_3020);
or U4713 (N_4713,N_3225,N_3511);
nor U4714 (N_4714,N_3957,N_2671);
nor U4715 (N_4715,N_3056,N_3810);
and U4716 (N_4716,N_2405,N_3191);
or U4717 (N_4717,N_2509,N_3208);
nand U4718 (N_4718,N_3448,N_3125);
and U4719 (N_4719,N_3585,N_3391);
and U4720 (N_4720,N_3838,N_3189);
or U4721 (N_4721,N_3982,N_3240);
nor U4722 (N_4722,N_2046,N_2747);
nand U4723 (N_4723,N_2652,N_2101);
or U4724 (N_4724,N_3168,N_2031);
and U4725 (N_4725,N_2222,N_2214);
or U4726 (N_4726,N_2667,N_2116);
and U4727 (N_4727,N_3167,N_2223);
and U4728 (N_4728,N_3914,N_3484);
or U4729 (N_4729,N_2228,N_2483);
nor U4730 (N_4730,N_3059,N_2882);
nand U4731 (N_4731,N_3375,N_2014);
nor U4732 (N_4732,N_2958,N_3943);
nor U4733 (N_4733,N_2420,N_3864);
and U4734 (N_4734,N_2142,N_2888);
and U4735 (N_4735,N_2515,N_3033);
and U4736 (N_4736,N_3508,N_2844);
or U4737 (N_4737,N_3633,N_3460);
nor U4738 (N_4738,N_3470,N_2563);
xor U4739 (N_4739,N_2576,N_3466);
nor U4740 (N_4740,N_2026,N_2985);
nand U4741 (N_4741,N_3515,N_3369);
nand U4742 (N_4742,N_3690,N_2227);
and U4743 (N_4743,N_2626,N_3322);
or U4744 (N_4744,N_2460,N_2586);
and U4745 (N_4745,N_3255,N_2279);
nand U4746 (N_4746,N_2259,N_3818);
and U4747 (N_4747,N_3560,N_3999);
nor U4748 (N_4748,N_2849,N_2322);
or U4749 (N_4749,N_2065,N_3415);
or U4750 (N_4750,N_2231,N_3044);
and U4751 (N_4751,N_3819,N_3518);
and U4752 (N_4752,N_3753,N_2597);
and U4753 (N_4753,N_3937,N_3530);
or U4754 (N_4754,N_2300,N_2276);
and U4755 (N_4755,N_2275,N_2423);
nand U4756 (N_4756,N_3154,N_2544);
or U4757 (N_4757,N_2763,N_2701);
nand U4758 (N_4758,N_2664,N_3594);
or U4759 (N_4759,N_2796,N_2970);
or U4760 (N_4760,N_3343,N_2610);
or U4761 (N_4761,N_2135,N_3565);
and U4762 (N_4762,N_3088,N_3363);
and U4763 (N_4763,N_3669,N_3678);
and U4764 (N_4764,N_3708,N_3319);
nand U4765 (N_4765,N_3039,N_3442);
xor U4766 (N_4766,N_2769,N_2151);
and U4767 (N_4767,N_2053,N_3326);
or U4768 (N_4768,N_3427,N_3495);
nor U4769 (N_4769,N_2206,N_2313);
and U4770 (N_4770,N_3941,N_2936);
and U4771 (N_4771,N_3439,N_2834);
and U4772 (N_4772,N_3054,N_2090);
nor U4773 (N_4773,N_3691,N_3034);
and U4774 (N_4774,N_3956,N_2833);
nor U4775 (N_4775,N_3037,N_3468);
nand U4776 (N_4776,N_3609,N_3377);
and U4777 (N_4777,N_2328,N_3577);
nor U4778 (N_4778,N_3850,N_2547);
nor U4779 (N_4779,N_2643,N_2261);
and U4780 (N_4780,N_2148,N_3824);
nand U4781 (N_4781,N_3228,N_3926);
nand U4782 (N_4782,N_2010,N_3094);
nand U4783 (N_4783,N_3849,N_2390);
nor U4784 (N_4784,N_2762,N_3446);
nor U4785 (N_4785,N_2622,N_2036);
nor U4786 (N_4786,N_3181,N_2018);
and U4787 (N_4787,N_2923,N_3401);
and U4788 (N_4788,N_2845,N_3417);
nand U4789 (N_4789,N_3997,N_2801);
and U4790 (N_4790,N_3265,N_3942);
or U4791 (N_4791,N_3224,N_3628);
nor U4792 (N_4792,N_3573,N_2601);
nor U4793 (N_4793,N_3238,N_3761);
nor U4794 (N_4794,N_2508,N_3009);
nor U4795 (N_4795,N_3105,N_2327);
nor U4796 (N_4796,N_3635,N_2928);
nand U4797 (N_4797,N_3781,N_2889);
and U4798 (N_4798,N_2000,N_3507);
nand U4799 (N_4799,N_3887,N_2006);
nand U4800 (N_4800,N_2229,N_3829);
or U4801 (N_4801,N_3254,N_2413);
or U4802 (N_4802,N_2193,N_2409);
nand U4803 (N_4803,N_2939,N_3487);
nand U4804 (N_4804,N_2163,N_2260);
nor U4805 (N_4805,N_3858,N_3301);
and U4806 (N_4806,N_2167,N_3161);
nor U4807 (N_4807,N_3679,N_3110);
nor U4808 (N_4808,N_2725,N_3072);
nand U4809 (N_4809,N_2767,N_3538);
nand U4810 (N_4810,N_3360,N_3719);
nor U4811 (N_4811,N_2138,N_3562);
and U4812 (N_4812,N_3476,N_2469);
and U4813 (N_4813,N_2326,N_3202);
or U4814 (N_4814,N_3532,N_3428);
nand U4815 (N_4815,N_2070,N_2221);
nand U4816 (N_4816,N_2708,N_3293);
and U4817 (N_4817,N_2868,N_2369);
and U4818 (N_4818,N_2886,N_3400);
nor U4819 (N_4819,N_2238,N_2315);
nand U4820 (N_4820,N_3602,N_3103);
and U4821 (N_4821,N_3658,N_2095);
nand U4822 (N_4822,N_2883,N_3572);
or U4823 (N_4823,N_3638,N_3040);
or U4824 (N_4824,N_2750,N_3771);
or U4825 (N_4825,N_2614,N_2029);
nand U4826 (N_4826,N_2149,N_3499);
or U4827 (N_4827,N_3754,N_2242);
nor U4828 (N_4828,N_2189,N_2458);
and U4829 (N_4829,N_2437,N_2038);
or U4830 (N_4830,N_3286,N_2165);
and U4831 (N_4831,N_3965,N_3107);
nor U4832 (N_4832,N_2354,N_3991);
or U4833 (N_4833,N_3866,N_3827);
or U4834 (N_4834,N_3539,N_2088);
nand U4835 (N_4835,N_2319,N_2772);
and U4836 (N_4836,N_3667,N_2929);
and U4837 (N_4837,N_2480,N_3142);
or U4838 (N_4838,N_3165,N_2481);
nor U4839 (N_4839,N_2377,N_3294);
nand U4840 (N_4840,N_3807,N_3318);
or U4841 (N_4841,N_3680,N_2592);
nor U4842 (N_4842,N_3551,N_2220);
nor U4843 (N_4843,N_2051,N_3176);
or U4844 (N_4844,N_3968,N_3169);
nor U4845 (N_4845,N_2472,N_3912);
or U4846 (N_4846,N_3526,N_2164);
and U4847 (N_4847,N_2621,N_2743);
or U4848 (N_4848,N_2519,N_2541);
or U4849 (N_4849,N_3330,N_2284);
and U4850 (N_4850,N_2461,N_2628);
nor U4851 (N_4851,N_2649,N_3397);
or U4852 (N_4852,N_3728,N_3366);
nor U4853 (N_4853,N_2205,N_2158);
nand U4854 (N_4854,N_2147,N_3092);
or U4855 (N_4855,N_3087,N_3450);
xnor U4856 (N_4856,N_2930,N_3727);
or U4857 (N_4857,N_2141,N_2367);
nor U4858 (N_4858,N_3774,N_3851);
nor U4859 (N_4859,N_3443,N_3987);
and U4860 (N_4860,N_2914,N_2637);
nand U4861 (N_4861,N_3132,N_3953);
nand U4862 (N_4862,N_3471,N_3323);
nor U4863 (N_4863,N_2119,N_3655);
and U4864 (N_4864,N_3311,N_3195);
and U4865 (N_4865,N_3607,N_2745);
nor U4866 (N_4866,N_3504,N_2039);
nand U4867 (N_4867,N_2507,N_3096);
or U4868 (N_4868,N_3915,N_2462);
or U4869 (N_4869,N_2118,N_3510);
and U4870 (N_4870,N_2066,N_2324);
nor U4871 (N_4871,N_3903,N_3895);
and U4872 (N_4872,N_3081,N_2692);
or U4873 (N_4873,N_3693,N_2239);
and U4874 (N_4874,N_3043,N_2226);
nand U4875 (N_4875,N_2814,N_3509);
nand U4876 (N_4876,N_2244,N_2631);
nand U4877 (N_4877,N_2784,N_3930);
nand U4878 (N_4878,N_2757,N_3713);
or U4879 (N_4879,N_3662,N_3888);
or U4880 (N_4880,N_3149,N_3772);
or U4881 (N_4881,N_3013,N_2009);
nor U4882 (N_4882,N_2711,N_2525);
nor U4883 (N_4883,N_2900,N_2371);
or U4884 (N_4884,N_2585,N_3454);
or U4885 (N_4885,N_2005,N_3738);
or U4886 (N_4886,N_2898,N_3799);
nand U4887 (N_4887,N_3292,N_2092);
or U4888 (N_4888,N_2878,N_2465);
nand U4889 (N_4889,N_2200,N_3645);
nand U4890 (N_4890,N_3650,N_3457);
or U4891 (N_4891,N_3998,N_3970);
xnor U4892 (N_4892,N_2662,N_3934);
or U4893 (N_4893,N_3378,N_2924);
nand U4894 (N_4894,N_2286,N_2404);
and U4895 (N_4895,N_2376,N_3393);
nand U4896 (N_4896,N_2021,N_2787);
or U4897 (N_4897,N_2805,N_3170);
and U4898 (N_4898,N_2976,N_3674);
and U4899 (N_4899,N_2675,N_2358);
and U4900 (N_4900,N_2512,N_3273);
nand U4901 (N_4901,N_3618,N_2732);
nor U4902 (N_4902,N_2393,N_2380);
nand U4903 (N_4903,N_2688,N_2341);
nor U4904 (N_4904,N_3841,N_3665);
and U4905 (N_4905,N_2726,N_3773);
nor U4906 (N_4906,N_3045,N_2064);
or U4907 (N_4907,N_3357,N_3348);
or U4908 (N_4908,N_2175,N_3855);
nand U4909 (N_4909,N_2430,N_3586);
and U4910 (N_4910,N_2272,N_2717);
nand U4911 (N_4911,N_3198,N_2492);
nand U4912 (N_4912,N_3485,N_2739);
and U4913 (N_4913,N_2496,N_3206);
or U4914 (N_4914,N_2311,N_3263);
and U4915 (N_4915,N_2866,N_2113);
nand U4916 (N_4916,N_2153,N_2532);
or U4917 (N_4917,N_3247,N_2288);
and U4918 (N_4918,N_3550,N_3186);
or U4919 (N_4919,N_3837,N_3578);
and U4920 (N_4920,N_3537,N_2366);
and U4921 (N_4921,N_3080,N_2399);
and U4922 (N_4922,N_3445,N_3746);
and U4923 (N_4923,N_2895,N_3634);
nand U4924 (N_4924,N_3312,N_2712);
or U4925 (N_4925,N_3580,N_3626);
nor U4926 (N_4926,N_3320,N_3885);
nand U4927 (N_4927,N_3200,N_3229);
or U4928 (N_4928,N_2780,N_3187);
nand U4929 (N_4929,N_2642,N_3297);
nand U4930 (N_4930,N_2781,N_2179);
or U4931 (N_4931,N_2109,N_3745);
and U4932 (N_4932,N_2250,N_3380);
or U4933 (N_4933,N_3177,N_2812);
and U4934 (N_4934,N_3564,N_3830);
nor U4935 (N_4935,N_2334,N_2190);
and U4936 (N_4936,N_2216,N_2524);
and U4937 (N_4937,N_2535,N_2819);
nor U4938 (N_4938,N_3491,N_2287);
nand U4939 (N_4939,N_2582,N_3805);
or U4940 (N_4940,N_3927,N_2060);
nor U4941 (N_4941,N_3675,N_3372);
nor U4942 (N_4942,N_2434,N_2536);
and U4943 (N_4943,N_3776,N_3524);
and U4944 (N_4944,N_3946,N_2256);
nand U4945 (N_4945,N_3520,N_3811);
and U4946 (N_4946,N_2432,N_2752);
and U4947 (N_4947,N_3977,N_3114);
and U4948 (N_4948,N_3686,N_3531);
and U4949 (N_4949,N_3842,N_3983);
and U4950 (N_4950,N_3768,N_3836);
or U4951 (N_4951,N_3063,N_3481);
or U4952 (N_4952,N_2170,N_2024);
or U4953 (N_4953,N_2074,N_2935);
nand U4954 (N_4954,N_2641,N_3627);
nand U4955 (N_4955,N_2453,N_2647);
or U4956 (N_4956,N_2488,N_3873);
and U4957 (N_4957,N_3870,N_3549);
nor U4958 (N_4958,N_2619,N_3211);
or U4959 (N_4959,N_2549,N_2696);
nand U4960 (N_4960,N_2577,N_3804);
nor U4961 (N_4961,N_3860,N_3875);
nand U4962 (N_4962,N_2352,N_2102);
nand U4963 (N_4963,N_3353,N_2625);
and U4964 (N_4964,N_2332,N_2659);
nand U4965 (N_4965,N_3329,N_2454);
nor U4966 (N_4966,N_2125,N_3624);
nand U4967 (N_4967,N_2452,N_2451);
nor U4968 (N_4968,N_3898,N_3731);
or U4969 (N_4969,N_2521,N_3795);
and U4970 (N_4970,N_2298,N_2904);
nor U4971 (N_4971,N_3831,N_2008);
nor U4972 (N_4972,N_2137,N_2020);
and U4973 (N_4973,N_2771,N_2033);
nor U4974 (N_4974,N_3381,N_2639);
and U4975 (N_4975,N_3612,N_3284);
nand U4976 (N_4976,N_3822,N_2230);
and U4977 (N_4977,N_2902,N_2499);
nor U4978 (N_4978,N_3534,N_2553);
or U4979 (N_4979,N_3419,N_3876);
nor U4980 (N_4980,N_3449,N_2445);
nand U4981 (N_4981,N_2950,N_2114);
nor U4982 (N_4982,N_3803,N_2337);
xor U4983 (N_4983,N_2815,N_3253);
nand U4984 (N_4984,N_2916,N_2482);
and U4985 (N_4985,N_2030,N_3395);
or U4986 (N_4986,N_2304,N_2079);
nor U4987 (N_4987,N_3709,N_2388);
and U4988 (N_4988,N_2438,N_2466);
nand U4989 (N_4989,N_2108,N_2121);
or U4990 (N_4990,N_2852,N_3622);
or U4991 (N_4991,N_3143,N_2616);
nor U4992 (N_4992,N_3408,N_3458);
and U4993 (N_4993,N_3304,N_2602);
or U4994 (N_4994,N_3702,N_2086);
or U4995 (N_4995,N_3828,N_2330);
nand U4996 (N_4996,N_2346,N_3659);
and U4997 (N_4997,N_2859,N_2263);
nand U4998 (N_4998,N_2531,N_3744);
or U4999 (N_4999,N_2858,N_2624);
nand U5000 (N_5000,N_2907,N_2564);
nor U5001 (N_5001,N_2771,N_2808);
nand U5002 (N_5002,N_3179,N_3483);
or U5003 (N_5003,N_3085,N_3850);
nand U5004 (N_5004,N_2170,N_3148);
or U5005 (N_5005,N_2413,N_3627);
and U5006 (N_5006,N_2009,N_3151);
nand U5007 (N_5007,N_3627,N_2564);
xnor U5008 (N_5008,N_2259,N_3222);
and U5009 (N_5009,N_2416,N_3117);
or U5010 (N_5010,N_2218,N_2453);
or U5011 (N_5011,N_3228,N_2004);
nor U5012 (N_5012,N_2499,N_3932);
and U5013 (N_5013,N_3239,N_3540);
xor U5014 (N_5014,N_2570,N_3752);
or U5015 (N_5015,N_3361,N_3462);
or U5016 (N_5016,N_2530,N_2234);
or U5017 (N_5017,N_2954,N_2407);
and U5018 (N_5018,N_2198,N_2654);
nand U5019 (N_5019,N_3265,N_3877);
nor U5020 (N_5020,N_2963,N_2600);
nand U5021 (N_5021,N_2271,N_3595);
or U5022 (N_5022,N_3882,N_2316);
nand U5023 (N_5023,N_2189,N_2667);
and U5024 (N_5024,N_2536,N_2773);
and U5025 (N_5025,N_2659,N_3417);
and U5026 (N_5026,N_3660,N_3947);
or U5027 (N_5027,N_3719,N_3814);
nor U5028 (N_5028,N_3143,N_2786);
nor U5029 (N_5029,N_2661,N_3540);
nor U5030 (N_5030,N_3028,N_2082);
and U5031 (N_5031,N_3531,N_3056);
and U5032 (N_5032,N_2650,N_2261);
xor U5033 (N_5033,N_2711,N_3173);
or U5034 (N_5034,N_2950,N_3506);
nor U5035 (N_5035,N_3973,N_3682);
or U5036 (N_5036,N_2824,N_3758);
or U5037 (N_5037,N_3583,N_2244);
nand U5038 (N_5038,N_3832,N_3489);
nand U5039 (N_5039,N_3398,N_3327);
and U5040 (N_5040,N_2366,N_3363);
nor U5041 (N_5041,N_2539,N_2200);
or U5042 (N_5042,N_3460,N_2430);
or U5043 (N_5043,N_3473,N_3983);
or U5044 (N_5044,N_3709,N_3818);
nor U5045 (N_5045,N_3435,N_2670);
nor U5046 (N_5046,N_3104,N_2453);
nor U5047 (N_5047,N_2866,N_3905);
and U5048 (N_5048,N_2497,N_3744);
or U5049 (N_5049,N_2991,N_3813);
and U5050 (N_5050,N_2870,N_3161);
nor U5051 (N_5051,N_3272,N_2114);
or U5052 (N_5052,N_3044,N_3696);
xnor U5053 (N_5053,N_3229,N_2249);
and U5054 (N_5054,N_2678,N_2485);
nand U5055 (N_5055,N_3621,N_3238);
and U5056 (N_5056,N_3794,N_2307);
and U5057 (N_5057,N_2627,N_3942);
or U5058 (N_5058,N_3377,N_3486);
or U5059 (N_5059,N_2429,N_3906);
or U5060 (N_5060,N_3863,N_2959);
nor U5061 (N_5061,N_3049,N_3441);
and U5062 (N_5062,N_2304,N_2369);
or U5063 (N_5063,N_2027,N_3426);
nand U5064 (N_5064,N_2998,N_2905);
nor U5065 (N_5065,N_2760,N_2136);
and U5066 (N_5066,N_3452,N_3860);
nand U5067 (N_5067,N_2733,N_3155);
and U5068 (N_5068,N_3877,N_2025);
nor U5069 (N_5069,N_2377,N_2455);
and U5070 (N_5070,N_3984,N_3475);
or U5071 (N_5071,N_2447,N_3532);
and U5072 (N_5072,N_3160,N_2433);
and U5073 (N_5073,N_2678,N_3560);
or U5074 (N_5074,N_3024,N_2271);
nor U5075 (N_5075,N_3756,N_3683);
and U5076 (N_5076,N_3973,N_3816);
or U5077 (N_5077,N_3220,N_3730);
xnor U5078 (N_5078,N_3907,N_3348);
nor U5079 (N_5079,N_3658,N_2815);
nand U5080 (N_5080,N_3536,N_3007);
and U5081 (N_5081,N_3643,N_2997);
nand U5082 (N_5082,N_3424,N_3616);
and U5083 (N_5083,N_2533,N_3447);
or U5084 (N_5084,N_3803,N_2831);
and U5085 (N_5085,N_3250,N_3842);
nand U5086 (N_5086,N_2007,N_2360);
nor U5087 (N_5087,N_3328,N_2240);
nor U5088 (N_5088,N_3629,N_3902);
or U5089 (N_5089,N_2414,N_2596);
or U5090 (N_5090,N_3189,N_3808);
nor U5091 (N_5091,N_3529,N_3597);
and U5092 (N_5092,N_2657,N_2347);
or U5093 (N_5093,N_2635,N_2834);
or U5094 (N_5094,N_3487,N_2538);
nor U5095 (N_5095,N_3780,N_2805);
or U5096 (N_5096,N_3560,N_2461);
nor U5097 (N_5097,N_2091,N_3120);
nor U5098 (N_5098,N_2921,N_2284);
nand U5099 (N_5099,N_3430,N_2491);
nor U5100 (N_5100,N_3333,N_2818);
and U5101 (N_5101,N_3144,N_3863);
nand U5102 (N_5102,N_3411,N_2722);
nor U5103 (N_5103,N_3077,N_3278);
or U5104 (N_5104,N_2799,N_3391);
nand U5105 (N_5105,N_2301,N_3794);
or U5106 (N_5106,N_2739,N_3451);
and U5107 (N_5107,N_2232,N_3865);
nor U5108 (N_5108,N_2974,N_3069);
or U5109 (N_5109,N_3001,N_2889);
nor U5110 (N_5110,N_2858,N_2742);
nand U5111 (N_5111,N_3658,N_2919);
nand U5112 (N_5112,N_3567,N_3506);
and U5113 (N_5113,N_3618,N_3728);
xor U5114 (N_5114,N_3290,N_2784);
and U5115 (N_5115,N_2686,N_3689);
and U5116 (N_5116,N_2415,N_2426);
or U5117 (N_5117,N_2357,N_2885);
nor U5118 (N_5118,N_3697,N_3214);
or U5119 (N_5119,N_2564,N_2608);
and U5120 (N_5120,N_3723,N_2982);
nand U5121 (N_5121,N_3301,N_2967);
nor U5122 (N_5122,N_3586,N_3398);
nor U5123 (N_5123,N_3313,N_2666);
nor U5124 (N_5124,N_3027,N_3390);
nand U5125 (N_5125,N_3147,N_3463);
or U5126 (N_5126,N_3804,N_3334);
nand U5127 (N_5127,N_3093,N_3575);
nand U5128 (N_5128,N_2274,N_2240);
or U5129 (N_5129,N_2798,N_2592);
or U5130 (N_5130,N_2185,N_3991);
or U5131 (N_5131,N_2834,N_3849);
and U5132 (N_5132,N_3683,N_3642);
and U5133 (N_5133,N_3574,N_2025);
and U5134 (N_5134,N_3994,N_2008);
and U5135 (N_5135,N_3546,N_3507);
nand U5136 (N_5136,N_3390,N_3407);
nand U5137 (N_5137,N_2374,N_2115);
nand U5138 (N_5138,N_3412,N_2499);
nor U5139 (N_5139,N_3752,N_2957);
and U5140 (N_5140,N_2905,N_3042);
nor U5141 (N_5141,N_3264,N_3331);
or U5142 (N_5142,N_3878,N_3234);
nor U5143 (N_5143,N_3824,N_3632);
nand U5144 (N_5144,N_2854,N_3232);
nor U5145 (N_5145,N_3179,N_3378);
or U5146 (N_5146,N_2416,N_3425);
nor U5147 (N_5147,N_2934,N_2923);
and U5148 (N_5148,N_2852,N_2160);
nand U5149 (N_5149,N_3399,N_3030);
nor U5150 (N_5150,N_2250,N_3825);
and U5151 (N_5151,N_2492,N_2813);
nand U5152 (N_5152,N_3889,N_2976);
nand U5153 (N_5153,N_3042,N_3511);
nor U5154 (N_5154,N_3359,N_2401);
nor U5155 (N_5155,N_3294,N_3470);
and U5156 (N_5156,N_2212,N_2996);
nor U5157 (N_5157,N_3522,N_3914);
nor U5158 (N_5158,N_2020,N_2379);
and U5159 (N_5159,N_2668,N_3094);
and U5160 (N_5160,N_2096,N_3653);
and U5161 (N_5161,N_3350,N_3948);
nor U5162 (N_5162,N_2084,N_3783);
or U5163 (N_5163,N_3334,N_2119);
and U5164 (N_5164,N_3874,N_2983);
nand U5165 (N_5165,N_2727,N_2389);
nand U5166 (N_5166,N_3509,N_2413);
nand U5167 (N_5167,N_2995,N_3217);
nor U5168 (N_5168,N_3307,N_3670);
nor U5169 (N_5169,N_3017,N_2169);
nand U5170 (N_5170,N_2507,N_3166);
nand U5171 (N_5171,N_3211,N_2735);
nor U5172 (N_5172,N_2221,N_2209);
nor U5173 (N_5173,N_2888,N_3553);
nand U5174 (N_5174,N_2293,N_3968);
or U5175 (N_5175,N_3088,N_3986);
nor U5176 (N_5176,N_2372,N_2205);
or U5177 (N_5177,N_3632,N_3962);
nor U5178 (N_5178,N_3974,N_2813);
nand U5179 (N_5179,N_3604,N_2514);
or U5180 (N_5180,N_2794,N_3555);
nor U5181 (N_5181,N_3701,N_3032);
or U5182 (N_5182,N_2826,N_2519);
or U5183 (N_5183,N_3723,N_3131);
nand U5184 (N_5184,N_2324,N_3401);
or U5185 (N_5185,N_3218,N_3215);
nor U5186 (N_5186,N_3642,N_2492);
and U5187 (N_5187,N_2932,N_3964);
nor U5188 (N_5188,N_3775,N_2152);
or U5189 (N_5189,N_2926,N_3008);
nor U5190 (N_5190,N_3173,N_3701);
nand U5191 (N_5191,N_3168,N_2884);
or U5192 (N_5192,N_3641,N_3945);
or U5193 (N_5193,N_2706,N_2625);
or U5194 (N_5194,N_3378,N_3474);
nand U5195 (N_5195,N_2856,N_2513);
nor U5196 (N_5196,N_3820,N_2415);
or U5197 (N_5197,N_2757,N_3873);
nand U5198 (N_5198,N_3993,N_2018);
nor U5199 (N_5199,N_3496,N_3783);
or U5200 (N_5200,N_3356,N_3362);
and U5201 (N_5201,N_2924,N_3374);
or U5202 (N_5202,N_3118,N_3150);
and U5203 (N_5203,N_2830,N_3209);
and U5204 (N_5204,N_3514,N_2493);
nand U5205 (N_5205,N_2934,N_3115);
nor U5206 (N_5206,N_3798,N_2538);
nand U5207 (N_5207,N_3956,N_2988);
nand U5208 (N_5208,N_3013,N_3106);
nor U5209 (N_5209,N_3822,N_3663);
or U5210 (N_5210,N_3375,N_2737);
nor U5211 (N_5211,N_2320,N_2668);
nand U5212 (N_5212,N_2840,N_2114);
nor U5213 (N_5213,N_2126,N_2412);
nand U5214 (N_5214,N_3870,N_2873);
nor U5215 (N_5215,N_2987,N_3600);
nand U5216 (N_5216,N_3384,N_2581);
nand U5217 (N_5217,N_3735,N_3395);
nand U5218 (N_5218,N_3949,N_3192);
and U5219 (N_5219,N_3197,N_3154);
and U5220 (N_5220,N_2572,N_3148);
nor U5221 (N_5221,N_2166,N_3044);
and U5222 (N_5222,N_3512,N_2108);
or U5223 (N_5223,N_3274,N_3973);
nor U5224 (N_5224,N_2439,N_3525);
nor U5225 (N_5225,N_3620,N_2035);
nor U5226 (N_5226,N_2994,N_2874);
and U5227 (N_5227,N_2886,N_3240);
and U5228 (N_5228,N_3294,N_2935);
nor U5229 (N_5229,N_3506,N_3529);
nand U5230 (N_5230,N_2429,N_2514);
and U5231 (N_5231,N_2764,N_3815);
or U5232 (N_5232,N_2065,N_3590);
and U5233 (N_5233,N_3218,N_2786);
nor U5234 (N_5234,N_2447,N_2653);
or U5235 (N_5235,N_2329,N_2650);
nor U5236 (N_5236,N_2159,N_2661);
and U5237 (N_5237,N_3932,N_3633);
nor U5238 (N_5238,N_2685,N_2197);
nand U5239 (N_5239,N_2893,N_2289);
nor U5240 (N_5240,N_2223,N_3517);
nand U5241 (N_5241,N_2297,N_3977);
nand U5242 (N_5242,N_2357,N_2894);
or U5243 (N_5243,N_3529,N_2198);
or U5244 (N_5244,N_2823,N_2850);
or U5245 (N_5245,N_2994,N_3175);
or U5246 (N_5246,N_3841,N_3475);
and U5247 (N_5247,N_2767,N_3143);
and U5248 (N_5248,N_3539,N_2585);
and U5249 (N_5249,N_3738,N_2800);
nor U5250 (N_5250,N_3070,N_3246);
nor U5251 (N_5251,N_2244,N_2158);
or U5252 (N_5252,N_3294,N_3222);
or U5253 (N_5253,N_3451,N_2540);
or U5254 (N_5254,N_3130,N_2881);
nand U5255 (N_5255,N_3930,N_3782);
and U5256 (N_5256,N_2297,N_2363);
nor U5257 (N_5257,N_2757,N_2573);
or U5258 (N_5258,N_3620,N_2053);
nand U5259 (N_5259,N_3886,N_3425);
nor U5260 (N_5260,N_2141,N_2519);
nand U5261 (N_5261,N_3345,N_2250);
nor U5262 (N_5262,N_3885,N_2913);
nor U5263 (N_5263,N_2912,N_2056);
or U5264 (N_5264,N_2037,N_3470);
nor U5265 (N_5265,N_2923,N_2399);
or U5266 (N_5266,N_3378,N_2786);
or U5267 (N_5267,N_3077,N_3522);
and U5268 (N_5268,N_3217,N_2659);
nor U5269 (N_5269,N_3179,N_2675);
and U5270 (N_5270,N_3802,N_2257);
or U5271 (N_5271,N_2816,N_3605);
or U5272 (N_5272,N_3310,N_2571);
and U5273 (N_5273,N_3527,N_2862);
and U5274 (N_5274,N_3072,N_3643);
and U5275 (N_5275,N_2552,N_2475);
nand U5276 (N_5276,N_2014,N_2308);
and U5277 (N_5277,N_3417,N_3744);
and U5278 (N_5278,N_3464,N_3289);
nor U5279 (N_5279,N_3770,N_3671);
nor U5280 (N_5280,N_3872,N_3670);
and U5281 (N_5281,N_3823,N_3307);
or U5282 (N_5282,N_3433,N_3787);
nand U5283 (N_5283,N_3009,N_3467);
nor U5284 (N_5284,N_3901,N_3637);
and U5285 (N_5285,N_3751,N_3149);
or U5286 (N_5286,N_2684,N_3366);
nand U5287 (N_5287,N_2740,N_2923);
and U5288 (N_5288,N_3865,N_3967);
nor U5289 (N_5289,N_3231,N_3592);
and U5290 (N_5290,N_2745,N_3203);
nand U5291 (N_5291,N_3473,N_3217);
and U5292 (N_5292,N_2139,N_3710);
nand U5293 (N_5293,N_2039,N_2890);
and U5294 (N_5294,N_3558,N_3888);
nand U5295 (N_5295,N_2531,N_2415);
nand U5296 (N_5296,N_3807,N_3770);
and U5297 (N_5297,N_3888,N_3222);
nor U5298 (N_5298,N_3250,N_3033);
nand U5299 (N_5299,N_3356,N_2614);
nor U5300 (N_5300,N_2428,N_2657);
nor U5301 (N_5301,N_3791,N_3914);
nor U5302 (N_5302,N_2273,N_3261);
and U5303 (N_5303,N_2040,N_2948);
or U5304 (N_5304,N_3801,N_2559);
nor U5305 (N_5305,N_2297,N_2431);
or U5306 (N_5306,N_2068,N_3399);
or U5307 (N_5307,N_3180,N_2974);
nand U5308 (N_5308,N_2101,N_3505);
nand U5309 (N_5309,N_2520,N_2972);
nand U5310 (N_5310,N_2990,N_3391);
nor U5311 (N_5311,N_2992,N_2636);
or U5312 (N_5312,N_3456,N_2092);
and U5313 (N_5313,N_2986,N_3625);
or U5314 (N_5314,N_2247,N_3195);
nand U5315 (N_5315,N_2759,N_3646);
nor U5316 (N_5316,N_2839,N_3908);
or U5317 (N_5317,N_3242,N_2388);
nand U5318 (N_5318,N_3930,N_2666);
nor U5319 (N_5319,N_3660,N_2956);
and U5320 (N_5320,N_2280,N_2265);
and U5321 (N_5321,N_2967,N_3775);
nand U5322 (N_5322,N_3718,N_3732);
or U5323 (N_5323,N_2912,N_2518);
or U5324 (N_5324,N_2600,N_2147);
nand U5325 (N_5325,N_2526,N_2267);
nor U5326 (N_5326,N_2299,N_2228);
nand U5327 (N_5327,N_3171,N_2821);
nand U5328 (N_5328,N_2554,N_3034);
nand U5329 (N_5329,N_3638,N_2045);
nand U5330 (N_5330,N_2579,N_3910);
nor U5331 (N_5331,N_3555,N_2795);
or U5332 (N_5332,N_3953,N_3252);
or U5333 (N_5333,N_2552,N_2960);
nand U5334 (N_5334,N_3355,N_3944);
and U5335 (N_5335,N_3801,N_2158);
or U5336 (N_5336,N_2072,N_3581);
nor U5337 (N_5337,N_3889,N_3632);
nor U5338 (N_5338,N_3842,N_2288);
nor U5339 (N_5339,N_2901,N_3660);
or U5340 (N_5340,N_3077,N_3828);
nand U5341 (N_5341,N_3374,N_2858);
and U5342 (N_5342,N_2060,N_3430);
nand U5343 (N_5343,N_3522,N_2058);
or U5344 (N_5344,N_2404,N_3509);
nor U5345 (N_5345,N_2662,N_3182);
and U5346 (N_5346,N_3895,N_3314);
nand U5347 (N_5347,N_3584,N_3697);
or U5348 (N_5348,N_2172,N_3054);
and U5349 (N_5349,N_2678,N_3981);
nand U5350 (N_5350,N_3320,N_3787);
and U5351 (N_5351,N_2157,N_2347);
nor U5352 (N_5352,N_2961,N_3807);
or U5353 (N_5353,N_2239,N_2537);
or U5354 (N_5354,N_2169,N_3577);
and U5355 (N_5355,N_2909,N_3292);
or U5356 (N_5356,N_2144,N_3459);
or U5357 (N_5357,N_2390,N_3517);
or U5358 (N_5358,N_2387,N_3973);
and U5359 (N_5359,N_2506,N_2652);
nand U5360 (N_5360,N_2185,N_3738);
nand U5361 (N_5361,N_2559,N_2795);
xor U5362 (N_5362,N_3055,N_3828);
nor U5363 (N_5363,N_2882,N_3391);
or U5364 (N_5364,N_2724,N_2137);
nand U5365 (N_5365,N_3535,N_2405);
nand U5366 (N_5366,N_3441,N_3185);
or U5367 (N_5367,N_2929,N_2562);
and U5368 (N_5368,N_2191,N_3804);
nand U5369 (N_5369,N_3802,N_3537);
nor U5370 (N_5370,N_2912,N_2789);
nor U5371 (N_5371,N_2615,N_2180);
and U5372 (N_5372,N_3240,N_2188);
nand U5373 (N_5373,N_2911,N_2733);
or U5374 (N_5374,N_2598,N_3192);
and U5375 (N_5375,N_2026,N_2917);
or U5376 (N_5376,N_2786,N_3995);
or U5377 (N_5377,N_2364,N_2294);
and U5378 (N_5378,N_3958,N_2720);
or U5379 (N_5379,N_2627,N_2160);
or U5380 (N_5380,N_3509,N_3294);
and U5381 (N_5381,N_2579,N_2141);
and U5382 (N_5382,N_2619,N_3156);
nor U5383 (N_5383,N_2842,N_3734);
and U5384 (N_5384,N_2413,N_2556);
and U5385 (N_5385,N_2419,N_2124);
or U5386 (N_5386,N_3486,N_2943);
or U5387 (N_5387,N_2207,N_2951);
nand U5388 (N_5388,N_2081,N_2611);
nor U5389 (N_5389,N_2509,N_2187);
and U5390 (N_5390,N_3547,N_3652);
or U5391 (N_5391,N_3774,N_2267);
nand U5392 (N_5392,N_2019,N_2179);
nor U5393 (N_5393,N_2932,N_2123);
and U5394 (N_5394,N_2596,N_2954);
or U5395 (N_5395,N_3023,N_2566);
nor U5396 (N_5396,N_3187,N_2653);
nand U5397 (N_5397,N_3033,N_3225);
or U5398 (N_5398,N_2106,N_3635);
and U5399 (N_5399,N_2278,N_3613);
nand U5400 (N_5400,N_3459,N_2560);
or U5401 (N_5401,N_3494,N_2241);
nand U5402 (N_5402,N_3335,N_3219);
nor U5403 (N_5403,N_3923,N_3974);
or U5404 (N_5404,N_2030,N_3523);
or U5405 (N_5405,N_2559,N_3552);
nor U5406 (N_5406,N_3199,N_3901);
nor U5407 (N_5407,N_2636,N_2564);
or U5408 (N_5408,N_3984,N_3166);
nand U5409 (N_5409,N_3555,N_3658);
or U5410 (N_5410,N_2215,N_2493);
nand U5411 (N_5411,N_3054,N_2548);
or U5412 (N_5412,N_2631,N_3215);
and U5413 (N_5413,N_2118,N_3528);
nor U5414 (N_5414,N_2999,N_2871);
or U5415 (N_5415,N_2230,N_2599);
or U5416 (N_5416,N_3717,N_2946);
nor U5417 (N_5417,N_3872,N_3487);
and U5418 (N_5418,N_2870,N_2111);
nor U5419 (N_5419,N_3153,N_2188);
or U5420 (N_5420,N_2541,N_2906);
nand U5421 (N_5421,N_2592,N_3751);
or U5422 (N_5422,N_2177,N_2403);
nor U5423 (N_5423,N_3285,N_2908);
or U5424 (N_5424,N_2495,N_3099);
and U5425 (N_5425,N_2957,N_2329);
and U5426 (N_5426,N_3940,N_2141);
nor U5427 (N_5427,N_2170,N_2007);
and U5428 (N_5428,N_3212,N_3930);
nor U5429 (N_5429,N_2549,N_3302);
nand U5430 (N_5430,N_2852,N_3858);
nor U5431 (N_5431,N_3761,N_2866);
nor U5432 (N_5432,N_2951,N_3744);
nand U5433 (N_5433,N_3830,N_3340);
nor U5434 (N_5434,N_3210,N_2506);
or U5435 (N_5435,N_3632,N_2617);
or U5436 (N_5436,N_3854,N_3047);
and U5437 (N_5437,N_2295,N_2799);
or U5438 (N_5438,N_3084,N_3582);
nor U5439 (N_5439,N_3586,N_3624);
and U5440 (N_5440,N_2343,N_3778);
or U5441 (N_5441,N_2488,N_3567);
or U5442 (N_5442,N_3206,N_2926);
or U5443 (N_5443,N_3559,N_3285);
nor U5444 (N_5444,N_3423,N_3354);
or U5445 (N_5445,N_2211,N_2571);
or U5446 (N_5446,N_3052,N_2959);
or U5447 (N_5447,N_3770,N_3391);
nand U5448 (N_5448,N_2199,N_3956);
nor U5449 (N_5449,N_3532,N_2588);
and U5450 (N_5450,N_3499,N_2663);
nand U5451 (N_5451,N_2602,N_3740);
or U5452 (N_5452,N_3490,N_2962);
nand U5453 (N_5453,N_3460,N_3420);
or U5454 (N_5454,N_3410,N_2516);
nor U5455 (N_5455,N_3552,N_3275);
nand U5456 (N_5456,N_3560,N_3516);
and U5457 (N_5457,N_2208,N_3802);
nand U5458 (N_5458,N_3829,N_2939);
or U5459 (N_5459,N_2657,N_2750);
or U5460 (N_5460,N_3661,N_3259);
and U5461 (N_5461,N_2241,N_3856);
nor U5462 (N_5462,N_2547,N_3563);
and U5463 (N_5463,N_3908,N_2511);
nor U5464 (N_5464,N_3347,N_2018);
xor U5465 (N_5465,N_3520,N_2198);
nand U5466 (N_5466,N_2956,N_2624);
and U5467 (N_5467,N_2946,N_3894);
nor U5468 (N_5468,N_3932,N_2421);
nor U5469 (N_5469,N_3029,N_2953);
or U5470 (N_5470,N_2844,N_2755);
and U5471 (N_5471,N_3408,N_2883);
nor U5472 (N_5472,N_2381,N_2245);
and U5473 (N_5473,N_3822,N_2491);
and U5474 (N_5474,N_3987,N_3620);
and U5475 (N_5475,N_2357,N_3698);
nor U5476 (N_5476,N_3383,N_2352);
or U5477 (N_5477,N_3317,N_2164);
nand U5478 (N_5478,N_2640,N_3655);
nor U5479 (N_5479,N_2768,N_3703);
or U5480 (N_5480,N_2007,N_3919);
and U5481 (N_5481,N_2314,N_3764);
or U5482 (N_5482,N_2523,N_2470);
nand U5483 (N_5483,N_3337,N_2735);
nand U5484 (N_5484,N_3415,N_3679);
and U5485 (N_5485,N_2487,N_3584);
and U5486 (N_5486,N_2578,N_3403);
nor U5487 (N_5487,N_2853,N_2227);
nand U5488 (N_5488,N_3536,N_3213);
nor U5489 (N_5489,N_2325,N_3515);
or U5490 (N_5490,N_3621,N_3643);
and U5491 (N_5491,N_2673,N_3673);
nand U5492 (N_5492,N_3307,N_2094);
and U5493 (N_5493,N_2369,N_3566);
nor U5494 (N_5494,N_2876,N_2164);
nand U5495 (N_5495,N_3993,N_3625);
and U5496 (N_5496,N_3741,N_3305);
nand U5497 (N_5497,N_3611,N_3206);
or U5498 (N_5498,N_2999,N_3508);
nand U5499 (N_5499,N_3430,N_3759);
nand U5500 (N_5500,N_3882,N_3859);
nand U5501 (N_5501,N_2691,N_2018);
nand U5502 (N_5502,N_2043,N_3885);
and U5503 (N_5503,N_3504,N_3403);
and U5504 (N_5504,N_3313,N_2709);
nand U5505 (N_5505,N_3560,N_3893);
nand U5506 (N_5506,N_3122,N_2675);
nor U5507 (N_5507,N_2351,N_3332);
and U5508 (N_5508,N_2460,N_3369);
or U5509 (N_5509,N_3420,N_2652);
nor U5510 (N_5510,N_3639,N_2657);
nor U5511 (N_5511,N_2694,N_2972);
nor U5512 (N_5512,N_3163,N_3230);
and U5513 (N_5513,N_3289,N_2963);
nand U5514 (N_5514,N_2389,N_2431);
nand U5515 (N_5515,N_3704,N_2178);
and U5516 (N_5516,N_2683,N_2231);
or U5517 (N_5517,N_3625,N_2347);
or U5518 (N_5518,N_2811,N_2034);
and U5519 (N_5519,N_3280,N_3588);
nand U5520 (N_5520,N_2832,N_3128);
and U5521 (N_5521,N_3739,N_2269);
nand U5522 (N_5522,N_2951,N_3269);
nand U5523 (N_5523,N_2992,N_3193);
or U5524 (N_5524,N_2172,N_3174);
or U5525 (N_5525,N_3107,N_2783);
nand U5526 (N_5526,N_3962,N_2261);
nand U5527 (N_5527,N_3532,N_2577);
nor U5528 (N_5528,N_2084,N_3050);
or U5529 (N_5529,N_2525,N_2989);
and U5530 (N_5530,N_2912,N_3167);
nand U5531 (N_5531,N_3252,N_2146);
or U5532 (N_5532,N_3945,N_3216);
and U5533 (N_5533,N_2711,N_3852);
nand U5534 (N_5534,N_2218,N_2291);
nand U5535 (N_5535,N_2201,N_3679);
nand U5536 (N_5536,N_3137,N_2425);
and U5537 (N_5537,N_3071,N_3464);
or U5538 (N_5538,N_3837,N_2726);
or U5539 (N_5539,N_2243,N_3376);
nand U5540 (N_5540,N_3206,N_2392);
nand U5541 (N_5541,N_2263,N_3521);
nand U5542 (N_5542,N_2359,N_3642);
and U5543 (N_5543,N_2174,N_2484);
and U5544 (N_5544,N_2022,N_2483);
nor U5545 (N_5545,N_2316,N_2895);
nor U5546 (N_5546,N_3775,N_3235);
nor U5547 (N_5547,N_2309,N_3722);
nor U5548 (N_5548,N_2646,N_2711);
nand U5549 (N_5549,N_3109,N_2188);
nand U5550 (N_5550,N_3112,N_3023);
or U5551 (N_5551,N_2560,N_3784);
and U5552 (N_5552,N_3984,N_2496);
or U5553 (N_5553,N_2355,N_2111);
nand U5554 (N_5554,N_3997,N_2757);
nor U5555 (N_5555,N_3847,N_3064);
and U5556 (N_5556,N_2080,N_2958);
and U5557 (N_5557,N_3797,N_2161);
nor U5558 (N_5558,N_3499,N_2342);
nor U5559 (N_5559,N_3548,N_3126);
nand U5560 (N_5560,N_2227,N_3540);
or U5561 (N_5561,N_3239,N_2384);
nor U5562 (N_5562,N_2836,N_2952);
nor U5563 (N_5563,N_3093,N_2444);
and U5564 (N_5564,N_2269,N_2090);
and U5565 (N_5565,N_3816,N_3080);
or U5566 (N_5566,N_3800,N_2581);
nor U5567 (N_5567,N_2569,N_3268);
or U5568 (N_5568,N_2870,N_2276);
nor U5569 (N_5569,N_2159,N_2333);
nand U5570 (N_5570,N_3398,N_3315);
nand U5571 (N_5571,N_2703,N_2850);
or U5572 (N_5572,N_3222,N_2505);
and U5573 (N_5573,N_3967,N_2515);
or U5574 (N_5574,N_2392,N_2102);
xnor U5575 (N_5575,N_3739,N_3124);
or U5576 (N_5576,N_2768,N_2790);
nor U5577 (N_5577,N_3927,N_2471);
nand U5578 (N_5578,N_2649,N_3589);
or U5579 (N_5579,N_3125,N_3955);
nand U5580 (N_5580,N_3105,N_3643);
nor U5581 (N_5581,N_3632,N_2090);
or U5582 (N_5582,N_3541,N_3171);
and U5583 (N_5583,N_2741,N_2033);
or U5584 (N_5584,N_3904,N_2019);
nand U5585 (N_5585,N_3741,N_3393);
nand U5586 (N_5586,N_2991,N_3442);
and U5587 (N_5587,N_2507,N_3612);
or U5588 (N_5588,N_3281,N_3343);
xor U5589 (N_5589,N_3652,N_2134);
or U5590 (N_5590,N_2820,N_3021);
nor U5591 (N_5591,N_3440,N_2344);
or U5592 (N_5592,N_3298,N_2056);
and U5593 (N_5593,N_2752,N_3612);
or U5594 (N_5594,N_2117,N_2935);
nand U5595 (N_5595,N_3848,N_3744);
and U5596 (N_5596,N_3672,N_3081);
or U5597 (N_5597,N_3012,N_3014);
nand U5598 (N_5598,N_3415,N_2158);
or U5599 (N_5599,N_2597,N_3201);
or U5600 (N_5600,N_3751,N_3463);
nand U5601 (N_5601,N_2142,N_2879);
nor U5602 (N_5602,N_2678,N_3667);
and U5603 (N_5603,N_3506,N_2821);
and U5604 (N_5604,N_2175,N_2051);
and U5605 (N_5605,N_3559,N_2777);
or U5606 (N_5606,N_3899,N_2520);
nand U5607 (N_5607,N_2595,N_2237);
or U5608 (N_5608,N_2319,N_2545);
or U5609 (N_5609,N_2502,N_2423);
nand U5610 (N_5610,N_3071,N_2788);
or U5611 (N_5611,N_3413,N_3030);
and U5612 (N_5612,N_3819,N_3911);
nor U5613 (N_5613,N_2124,N_2036);
and U5614 (N_5614,N_2054,N_3466);
and U5615 (N_5615,N_2256,N_2434);
or U5616 (N_5616,N_2194,N_2782);
and U5617 (N_5617,N_3464,N_2189);
nand U5618 (N_5618,N_3346,N_2018);
or U5619 (N_5619,N_2449,N_2360);
nor U5620 (N_5620,N_2280,N_3594);
and U5621 (N_5621,N_3810,N_2281);
or U5622 (N_5622,N_3280,N_2305);
nor U5623 (N_5623,N_2109,N_2922);
and U5624 (N_5624,N_2264,N_2540);
nor U5625 (N_5625,N_3273,N_2918);
nor U5626 (N_5626,N_2562,N_2097);
or U5627 (N_5627,N_2921,N_3761);
nor U5628 (N_5628,N_3326,N_3955);
and U5629 (N_5629,N_3727,N_3195);
nor U5630 (N_5630,N_2267,N_3842);
nand U5631 (N_5631,N_2587,N_2565);
nand U5632 (N_5632,N_2823,N_2886);
nor U5633 (N_5633,N_2983,N_3327);
and U5634 (N_5634,N_3930,N_3592);
nand U5635 (N_5635,N_2582,N_3430);
nor U5636 (N_5636,N_2306,N_3701);
nand U5637 (N_5637,N_2494,N_3240);
nor U5638 (N_5638,N_3377,N_2940);
nor U5639 (N_5639,N_3286,N_2813);
and U5640 (N_5640,N_3825,N_3645);
nor U5641 (N_5641,N_3497,N_2419);
and U5642 (N_5642,N_3829,N_3645);
or U5643 (N_5643,N_2811,N_2824);
nand U5644 (N_5644,N_3101,N_3329);
and U5645 (N_5645,N_2667,N_3889);
nand U5646 (N_5646,N_3864,N_2000);
nand U5647 (N_5647,N_2594,N_3886);
nor U5648 (N_5648,N_3652,N_3210);
and U5649 (N_5649,N_3980,N_3173);
nand U5650 (N_5650,N_2408,N_3885);
or U5651 (N_5651,N_3895,N_3749);
and U5652 (N_5652,N_2493,N_3011);
or U5653 (N_5653,N_2850,N_3263);
or U5654 (N_5654,N_2274,N_2737);
nand U5655 (N_5655,N_3911,N_3317);
nand U5656 (N_5656,N_2592,N_3286);
nor U5657 (N_5657,N_3589,N_3763);
or U5658 (N_5658,N_3113,N_2987);
nor U5659 (N_5659,N_3407,N_3705);
or U5660 (N_5660,N_3717,N_2630);
or U5661 (N_5661,N_3409,N_2328);
or U5662 (N_5662,N_2306,N_3367);
nor U5663 (N_5663,N_2296,N_2816);
or U5664 (N_5664,N_3335,N_3467);
and U5665 (N_5665,N_3073,N_2840);
nor U5666 (N_5666,N_3025,N_2225);
nor U5667 (N_5667,N_2636,N_2573);
or U5668 (N_5668,N_3267,N_2244);
and U5669 (N_5669,N_2987,N_3049);
nand U5670 (N_5670,N_3248,N_3663);
or U5671 (N_5671,N_2673,N_2605);
or U5672 (N_5672,N_2178,N_2626);
nor U5673 (N_5673,N_3312,N_2289);
xnor U5674 (N_5674,N_2984,N_2431);
nand U5675 (N_5675,N_2705,N_2005);
nor U5676 (N_5676,N_2223,N_3337);
nor U5677 (N_5677,N_3217,N_2151);
and U5678 (N_5678,N_2414,N_2420);
or U5679 (N_5679,N_3742,N_3394);
and U5680 (N_5680,N_2111,N_3625);
nand U5681 (N_5681,N_3653,N_3981);
or U5682 (N_5682,N_2535,N_3143);
or U5683 (N_5683,N_3359,N_3189);
or U5684 (N_5684,N_3787,N_3806);
nor U5685 (N_5685,N_2378,N_2301);
nor U5686 (N_5686,N_2393,N_2217);
or U5687 (N_5687,N_2121,N_2510);
and U5688 (N_5688,N_2734,N_2958);
or U5689 (N_5689,N_2414,N_2382);
and U5690 (N_5690,N_2020,N_2127);
nor U5691 (N_5691,N_3475,N_2573);
nor U5692 (N_5692,N_2559,N_2943);
nor U5693 (N_5693,N_3877,N_3650);
or U5694 (N_5694,N_3158,N_3383);
nand U5695 (N_5695,N_2332,N_2996);
or U5696 (N_5696,N_2239,N_3061);
nand U5697 (N_5697,N_3411,N_3474);
nand U5698 (N_5698,N_3642,N_2078);
or U5699 (N_5699,N_3025,N_2699);
nor U5700 (N_5700,N_2543,N_3041);
nor U5701 (N_5701,N_2559,N_2488);
or U5702 (N_5702,N_3077,N_3326);
nor U5703 (N_5703,N_2582,N_2360);
nor U5704 (N_5704,N_3349,N_3026);
nor U5705 (N_5705,N_3755,N_3443);
or U5706 (N_5706,N_3690,N_2551);
and U5707 (N_5707,N_3204,N_3656);
nor U5708 (N_5708,N_3928,N_2894);
or U5709 (N_5709,N_2345,N_3186);
nand U5710 (N_5710,N_2787,N_2784);
nor U5711 (N_5711,N_3373,N_3699);
nand U5712 (N_5712,N_2430,N_2023);
nand U5713 (N_5713,N_3141,N_3071);
nor U5714 (N_5714,N_2876,N_2545);
or U5715 (N_5715,N_3273,N_3830);
nand U5716 (N_5716,N_3827,N_2291);
nor U5717 (N_5717,N_3487,N_2692);
or U5718 (N_5718,N_2952,N_2209);
or U5719 (N_5719,N_2532,N_3281);
and U5720 (N_5720,N_3325,N_3908);
nand U5721 (N_5721,N_3449,N_3341);
or U5722 (N_5722,N_2223,N_3250);
nor U5723 (N_5723,N_3666,N_2979);
nand U5724 (N_5724,N_3200,N_2295);
and U5725 (N_5725,N_2846,N_3412);
and U5726 (N_5726,N_3676,N_3174);
nor U5727 (N_5727,N_3259,N_3401);
nand U5728 (N_5728,N_2250,N_3454);
nor U5729 (N_5729,N_3729,N_3173);
or U5730 (N_5730,N_3836,N_3965);
or U5731 (N_5731,N_2785,N_2496);
nor U5732 (N_5732,N_2466,N_2015);
nor U5733 (N_5733,N_2553,N_2515);
nand U5734 (N_5734,N_2091,N_3089);
nand U5735 (N_5735,N_3841,N_2161);
or U5736 (N_5736,N_2514,N_2024);
or U5737 (N_5737,N_2815,N_3404);
nor U5738 (N_5738,N_3357,N_3875);
or U5739 (N_5739,N_2107,N_2935);
or U5740 (N_5740,N_2665,N_3901);
or U5741 (N_5741,N_2369,N_3475);
or U5742 (N_5742,N_3093,N_3952);
nor U5743 (N_5743,N_2247,N_2605);
or U5744 (N_5744,N_2255,N_3949);
nand U5745 (N_5745,N_3807,N_3250);
xnor U5746 (N_5746,N_3820,N_3734);
or U5747 (N_5747,N_3639,N_2158);
and U5748 (N_5748,N_3066,N_2205);
nor U5749 (N_5749,N_3143,N_2070);
nor U5750 (N_5750,N_2748,N_2171);
and U5751 (N_5751,N_2011,N_2730);
nand U5752 (N_5752,N_3510,N_2264);
or U5753 (N_5753,N_2326,N_2760);
and U5754 (N_5754,N_2839,N_3005);
and U5755 (N_5755,N_3410,N_3711);
or U5756 (N_5756,N_3476,N_3872);
and U5757 (N_5757,N_2507,N_2833);
or U5758 (N_5758,N_2977,N_3666);
and U5759 (N_5759,N_2032,N_2035);
nor U5760 (N_5760,N_3365,N_3645);
or U5761 (N_5761,N_3918,N_3611);
or U5762 (N_5762,N_2288,N_3514);
nor U5763 (N_5763,N_3392,N_3617);
nor U5764 (N_5764,N_2926,N_3942);
nor U5765 (N_5765,N_3782,N_2324);
nand U5766 (N_5766,N_2962,N_3058);
nor U5767 (N_5767,N_2150,N_3859);
and U5768 (N_5768,N_2260,N_2578);
and U5769 (N_5769,N_3365,N_3259);
nand U5770 (N_5770,N_2653,N_3378);
and U5771 (N_5771,N_2278,N_2717);
and U5772 (N_5772,N_3683,N_3882);
and U5773 (N_5773,N_3103,N_2430);
or U5774 (N_5774,N_2804,N_3145);
and U5775 (N_5775,N_3084,N_2232);
or U5776 (N_5776,N_3277,N_2331);
or U5777 (N_5777,N_3043,N_2313);
nand U5778 (N_5778,N_2346,N_2064);
or U5779 (N_5779,N_3742,N_2485);
and U5780 (N_5780,N_3635,N_2704);
and U5781 (N_5781,N_3794,N_3022);
nand U5782 (N_5782,N_2001,N_2759);
and U5783 (N_5783,N_3768,N_2562);
or U5784 (N_5784,N_2476,N_3014);
nand U5785 (N_5785,N_2190,N_2080);
and U5786 (N_5786,N_2682,N_2740);
and U5787 (N_5787,N_3193,N_3367);
nand U5788 (N_5788,N_2309,N_3445);
nor U5789 (N_5789,N_2515,N_3739);
nand U5790 (N_5790,N_3062,N_3056);
or U5791 (N_5791,N_3554,N_3462);
nand U5792 (N_5792,N_2683,N_2338);
nand U5793 (N_5793,N_3548,N_3239);
nor U5794 (N_5794,N_3262,N_2546);
nor U5795 (N_5795,N_3587,N_3227);
and U5796 (N_5796,N_2017,N_3910);
or U5797 (N_5797,N_2909,N_3699);
nor U5798 (N_5798,N_2156,N_3600);
or U5799 (N_5799,N_3751,N_3969);
nand U5800 (N_5800,N_3367,N_2729);
xnor U5801 (N_5801,N_2715,N_2321);
or U5802 (N_5802,N_2619,N_2207);
and U5803 (N_5803,N_2564,N_3376);
nand U5804 (N_5804,N_3452,N_2101);
or U5805 (N_5805,N_3495,N_3995);
nand U5806 (N_5806,N_3453,N_3533);
or U5807 (N_5807,N_3200,N_2073);
nand U5808 (N_5808,N_3694,N_3843);
xor U5809 (N_5809,N_3220,N_3007);
and U5810 (N_5810,N_3383,N_3862);
or U5811 (N_5811,N_3362,N_3261);
or U5812 (N_5812,N_3660,N_3409);
nand U5813 (N_5813,N_2441,N_3361);
nand U5814 (N_5814,N_3948,N_3198);
xor U5815 (N_5815,N_3577,N_3712);
nand U5816 (N_5816,N_3677,N_3178);
and U5817 (N_5817,N_3041,N_2260);
nor U5818 (N_5818,N_2166,N_3811);
nor U5819 (N_5819,N_2307,N_3875);
or U5820 (N_5820,N_2761,N_2967);
nand U5821 (N_5821,N_2952,N_2344);
and U5822 (N_5822,N_3965,N_3723);
and U5823 (N_5823,N_3380,N_2028);
nor U5824 (N_5824,N_3641,N_3610);
nor U5825 (N_5825,N_3390,N_3226);
nor U5826 (N_5826,N_3572,N_2944);
nand U5827 (N_5827,N_3324,N_3045);
nand U5828 (N_5828,N_2901,N_3010);
nor U5829 (N_5829,N_3932,N_3670);
nand U5830 (N_5830,N_3245,N_3078);
or U5831 (N_5831,N_2670,N_3855);
nand U5832 (N_5832,N_3806,N_2110);
nand U5833 (N_5833,N_2946,N_2793);
and U5834 (N_5834,N_3675,N_3086);
and U5835 (N_5835,N_3462,N_3655);
nand U5836 (N_5836,N_3920,N_2406);
xnor U5837 (N_5837,N_3567,N_2615);
nand U5838 (N_5838,N_3036,N_3038);
or U5839 (N_5839,N_2851,N_3721);
nor U5840 (N_5840,N_2016,N_3341);
nand U5841 (N_5841,N_3235,N_2690);
and U5842 (N_5842,N_2139,N_2645);
nand U5843 (N_5843,N_2659,N_3044);
and U5844 (N_5844,N_3501,N_2534);
or U5845 (N_5845,N_2865,N_3882);
and U5846 (N_5846,N_2305,N_2259);
or U5847 (N_5847,N_3064,N_3087);
nor U5848 (N_5848,N_2812,N_3595);
or U5849 (N_5849,N_2118,N_2576);
nand U5850 (N_5850,N_3799,N_2272);
or U5851 (N_5851,N_2264,N_3896);
nand U5852 (N_5852,N_2857,N_3727);
nand U5853 (N_5853,N_2267,N_2152);
or U5854 (N_5854,N_2413,N_2721);
nor U5855 (N_5855,N_3002,N_3429);
and U5856 (N_5856,N_2630,N_2094);
nor U5857 (N_5857,N_2982,N_2401);
nor U5858 (N_5858,N_3592,N_2074);
and U5859 (N_5859,N_2760,N_2749);
nand U5860 (N_5860,N_2590,N_2442);
or U5861 (N_5861,N_2267,N_3189);
nor U5862 (N_5862,N_2985,N_3312);
or U5863 (N_5863,N_3396,N_2868);
and U5864 (N_5864,N_3506,N_3167);
and U5865 (N_5865,N_3911,N_3367);
or U5866 (N_5866,N_3952,N_3596);
nor U5867 (N_5867,N_2706,N_2199);
and U5868 (N_5868,N_3228,N_2612);
and U5869 (N_5869,N_3933,N_3523);
nand U5870 (N_5870,N_3500,N_3249);
nand U5871 (N_5871,N_3977,N_2764);
nand U5872 (N_5872,N_2409,N_3916);
nor U5873 (N_5873,N_2726,N_2684);
and U5874 (N_5874,N_3692,N_3190);
nor U5875 (N_5875,N_2228,N_2720);
or U5876 (N_5876,N_2917,N_3940);
xor U5877 (N_5877,N_3689,N_2229);
or U5878 (N_5878,N_3129,N_2837);
and U5879 (N_5879,N_3829,N_3901);
and U5880 (N_5880,N_2982,N_2276);
and U5881 (N_5881,N_2198,N_3418);
nand U5882 (N_5882,N_2767,N_2273);
and U5883 (N_5883,N_2470,N_2851);
or U5884 (N_5884,N_2235,N_3398);
nand U5885 (N_5885,N_2602,N_2094);
or U5886 (N_5886,N_2302,N_2569);
and U5887 (N_5887,N_2880,N_2039);
nand U5888 (N_5888,N_3548,N_3131);
nand U5889 (N_5889,N_2261,N_2399);
and U5890 (N_5890,N_2589,N_2843);
nand U5891 (N_5891,N_2607,N_3555);
or U5892 (N_5892,N_3870,N_3580);
or U5893 (N_5893,N_3021,N_3411);
or U5894 (N_5894,N_3406,N_2728);
and U5895 (N_5895,N_3979,N_3409);
and U5896 (N_5896,N_3188,N_3885);
nand U5897 (N_5897,N_3642,N_3981);
or U5898 (N_5898,N_3592,N_2008);
and U5899 (N_5899,N_2210,N_2884);
nand U5900 (N_5900,N_3488,N_2960);
or U5901 (N_5901,N_2365,N_2344);
and U5902 (N_5902,N_2041,N_2834);
and U5903 (N_5903,N_3957,N_3949);
nor U5904 (N_5904,N_2126,N_3727);
and U5905 (N_5905,N_3584,N_3703);
nor U5906 (N_5906,N_2529,N_2772);
nor U5907 (N_5907,N_2930,N_3165);
and U5908 (N_5908,N_3229,N_3114);
nand U5909 (N_5909,N_2172,N_3994);
or U5910 (N_5910,N_2007,N_3158);
nand U5911 (N_5911,N_2238,N_2196);
nand U5912 (N_5912,N_2536,N_2751);
and U5913 (N_5913,N_2727,N_3869);
nor U5914 (N_5914,N_2365,N_2190);
or U5915 (N_5915,N_3912,N_2449);
or U5916 (N_5916,N_2266,N_3184);
nand U5917 (N_5917,N_3697,N_3946);
nand U5918 (N_5918,N_3345,N_3890);
and U5919 (N_5919,N_2734,N_2184);
nor U5920 (N_5920,N_3512,N_3789);
and U5921 (N_5921,N_2233,N_3113);
or U5922 (N_5922,N_2709,N_3829);
nor U5923 (N_5923,N_2995,N_2799);
nand U5924 (N_5924,N_3984,N_2037);
nor U5925 (N_5925,N_2150,N_2307);
nand U5926 (N_5926,N_3003,N_3272);
and U5927 (N_5927,N_2942,N_3091);
and U5928 (N_5928,N_2196,N_2363);
or U5929 (N_5929,N_3273,N_3269);
nand U5930 (N_5930,N_2258,N_2567);
nand U5931 (N_5931,N_2806,N_3780);
nand U5932 (N_5932,N_2792,N_2332);
or U5933 (N_5933,N_3491,N_2694);
or U5934 (N_5934,N_2066,N_3443);
nand U5935 (N_5935,N_3370,N_2064);
or U5936 (N_5936,N_2731,N_3287);
and U5937 (N_5937,N_3017,N_2139);
xnor U5938 (N_5938,N_3681,N_2133);
and U5939 (N_5939,N_3993,N_2366);
and U5940 (N_5940,N_2849,N_2997);
and U5941 (N_5941,N_2289,N_2717);
xnor U5942 (N_5942,N_3862,N_3088);
or U5943 (N_5943,N_2120,N_3658);
nor U5944 (N_5944,N_2869,N_3337);
and U5945 (N_5945,N_3675,N_2373);
nand U5946 (N_5946,N_3179,N_3885);
nand U5947 (N_5947,N_2915,N_3065);
or U5948 (N_5948,N_3042,N_3097);
or U5949 (N_5949,N_2825,N_2298);
or U5950 (N_5950,N_3598,N_2264);
nand U5951 (N_5951,N_2969,N_2076);
nand U5952 (N_5952,N_3356,N_3334);
nand U5953 (N_5953,N_3646,N_3711);
nand U5954 (N_5954,N_2456,N_3988);
nor U5955 (N_5955,N_3893,N_3188);
nor U5956 (N_5956,N_3068,N_3027);
and U5957 (N_5957,N_3197,N_3275);
nor U5958 (N_5958,N_3718,N_3325);
nor U5959 (N_5959,N_2596,N_3519);
nand U5960 (N_5960,N_3848,N_3751);
nor U5961 (N_5961,N_3617,N_3656);
or U5962 (N_5962,N_3777,N_2217);
nand U5963 (N_5963,N_3002,N_2907);
and U5964 (N_5964,N_2769,N_2315);
nor U5965 (N_5965,N_2517,N_2231);
or U5966 (N_5966,N_3993,N_3219);
or U5967 (N_5967,N_2588,N_3799);
nand U5968 (N_5968,N_3421,N_3394);
nand U5969 (N_5969,N_3275,N_3593);
and U5970 (N_5970,N_2731,N_3799);
nor U5971 (N_5971,N_2537,N_3055);
or U5972 (N_5972,N_3868,N_3200);
and U5973 (N_5973,N_2075,N_2364);
nor U5974 (N_5974,N_3080,N_2834);
nor U5975 (N_5975,N_3208,N_3670);
and U5976 (N_5976,N_2023,N_3451);
or U5977 (N_5977,N_2453,N_3219);
and U5978 (N_5978,N_2095,N_3293);
or U5979 (N_5979,N_3999,N_3042);
or U5980 (N_5980,N_2994,N_2608);
xor U5981 (N_5981,N_3653,N_2802);
or U5982 (N_5982,N_3676,N_2374);
nor U5983 (N_5983,N_2404,N_2903);
nor U5984 (N_5984,N_2018,N_3672);
and U5985 (N_5985,N_3560,N_2457);
or U5986 (N_5986,N_3744,N_3020);
and U5987 (N_5987,N_3168,N_3913);
nor U5988 (N_5988,N_3647,N_2277);
xor U5989 (N_5989,N_2924,N_2520);
nor U5990 (N_5990,N_2910,N_3036);
nor U5991 (N_5991,N_3799,N_2275);
or U5992 (N_5992,N_3199,N_2425);
nand U5993 (N_5993,N_2171,N_2531);
and U5994 (N_5994,N_2784,N_3374);
nand U5995 (N_5995,N_3696,N_3617);
nand U5996 (N_5996,N_3080,N_2816);
and U5997 (N_5997,N_3054,N_3823);
and U5998 (N_5998,N_2352,N_2453);
and U5999 (N_5999,N_3750,N_2799);
and U6000 (N_6000,N_4150,N_4951);
and U6001 (N_6001,N_5985,N_5391);
or U6002 (N_6002,N_4971,N_4461);
and U6003 (N_6003,N_4518,N_4015);
and U6004 (N_6004,N_5368,N_5856);
and U6005 (N_6005,N_5175,N_4705);
nor U6006 (N_6006,N_5589,N_4254);
nand U6007 (N_6007,N_5786,N_4277);
and U6008 (N_6008,N_4391,N_4716);
and U6009 (N_6009,N_5653,N_4526);
or U6010 (N_6010,N_5663,N_5204);
or U6011 (N_6011,N_5143,N_4649);
nor U6012 (N_6012,N_5327,N_4365);
nor U6013 (N_6013,N_5693,N_4779);
and U6014 (N_6014,N_4039,N_4650);
nand U6015 (N_6015,N_5684,N_5138);
and U6016 (N_6016,N_4556,N_5615);
nand U6017 (N_6017,N_4463,N_4354);
nand U6018 (N_6018,N_5257,N_4542);
and U6019 (N_6019,N_4845,N_4214);
nand U6020 (N_6020,N_4814,N_5506);
and U6021 (N_6021,N_4071,N_4078);
and U6022 (N_6022,N_4298,N_4351);
or U6023 (N_6023,N_5283,N_4812);
or U6024 (N_6024,N_4108,N_4822);
and U6025 (N_6025,N_5632,N_4265);
and U6026 (N_6026,N_4737,N_4367);
or U6027 (N_6027,N_4068,N_5962);
nand U6028 (N_6028,N_4771,N_4429);
and U6029 (N_6029,N_4188,N_5490);
or U6030 (N_6030,N_5963,N_4464);
or U6031 (N_6031,N_5101,N_5484);
nor U6032 (N_6032,N_4861,N_5137);
nand U6033 (N_6033,N_5937,N_5209);
or U6034 (N_6034,N_5690,N_5075);
and U6035 (N_6035,N_4191,N_4739);
or U6036 (N_6036,N_4131,N_4567);
and U6037 (N_6037,N_5661,N_5650);
and U6038 (N_6038,N_4043,N_5124);
and U6039 (N_6039,N_5772,N_4968);
and U6040 (N_6040,N_5636,N_5657);
nor U6041 (N_6041,N_4212,N_4830);
and U6042 (N_6042,N_4230,N_5215);
or U6043 (N_6043,N_5775,N_5286);
and U6044 (N_6044,N_4081,N_4720);
or U6045 (N_6045,N_5505,N_4439);
or U6046 (N_6046,N_5904,N_5940);
and U6047 (N_6047,N_5377,N_5617);
nor U6048 (N_6048,N_4988,N_4501);
nand U6049 (N_6049,N_4566,N_5167);
or U6050 (N_6050,N_4061,N_5970);
or U6051 (N_6051,N_5934,N_4754);
nor U6052 (N_6052,N_4255,N_5005);
and U6053 (N_6053,N_4079,N_4408);
or U6054 (N_6054,N_5964,N_5968);
and U6055 (N_6055,N_5202,N_5475);
nand U6056 (N_6056,N_4905,N_5773);
or U6057 (N_6057,N_4472,N_4616);
nand U6058 (N_6058,N_4892,N_4162);
or U6059 (N_6059,N_5106,N_4019);
nand U6060 (N_6060,N_5523,N_5777);
nor U6061 (N_6061,N_4655,N_4453);
and U6062 (N_6062,N_4925,N_4625);
and U6063 (N_6063,N_4028,N_4687);
nor U6064 (N_6064,N_4602,N_4980);
or U6065 (N_6065,N_4732,N_4883);
nand U6066 (N_6066,N_5725,N_5876);
and U6067 (N_6067,N_5910,N_5706);
or U6068 (N_6068,N_4163,N_5805);
nor U6069 (N_6069,N_4099,N_5037);
and U6070 (N_6070,N_4889,N_4490);
xor U6071 (N_6071,N_5884,N_4201);
nor U6072 (N_6072,N_5294,N_4864);
nand U6073 (N_6073,N_5015,N_4857);
nor U6074 (N_6074,N_4138,N_5079);
or U6075 (N_6075,N_4420,N_5251);
nor U6076 (N_6076,N_4316,N_4247);
nand U6077 (N_6077,N_4603,N_5983);
or U6078 (N_6078,N_4090,N_4972);
and U6079 (N_6079,N_4746,N_5715);
nand U6080 (N_6080,N_5580,N_4995);
and U6081 (N_6081,N_4522,N_5383);
nor U6082 (N_6082,N_5556,N_4406);
nand U6083 (N_6083,N_5356,N_4854);
and U6084 (N_6084,N_5945,N_5051);
and U6085 (N_6085,N_5102,N_4363);
and U6086 (N_6086,N_5266,N_4381);
or U6087 (N_6087,N_5601,N_4016);
nor U6088 (N_6088,N_4799,N_4340);
nor U6089 (N_6089,N_4719,N_5752);
and U6090 (N_6090,N_5526,N_4173);
or U6091 (N_6091,N_4009,N_5221);
or U6092 (N_6092,N_5062,N_4535);
and U6093 (N_6093,N_5927,N_4317);
nor U6094 (N_6094,N_4881,N_4144);
nand U6095 (N_6095,N_4303,N_5882);
nor U6096 (N_6096,N_4760,N_4103);
and U6097 (N_6097,N_4748,N_5905);
nor U6098 (N_6098,N_5990,N_5564);
and U6099 (N_6099,N_5742,N_5265);
or U6100 (N_6100,N_5982,N_5360);
nor U6101 (N_6101,N_5868,N_4145);
or U6102 (N_6102,N_4738,N_5729);
and U6103 (N_6103,N_4233,N_5282);
and U6104 (N_6104,N_4614,N_4879);
nor U6105 (N_6105,N_5486,N_4693);
or U6106 (N_6106,N_4778,N_5400);
nand U6107 (N_6107,N_4253,N_5222);
and U6108 (N_6108,N_4989,N_4803);
nor U6109 (N_6109,N_5536,N_4880);
or U6110 (N_6110,N_5631,N_4949);
or U6111 (N_6111,N_5353,N_4390);
and U6112 (N_6112,N_5069,N_4249);
and U6113 (N_6113,N_4063,N_4853);
or U6114 (N_6114,N_5198,N_5507);
and U6115 (N_6115,N_4281,N_4528);
and U6116 (N_6116,N_4809,N_5158);
and U6117 (N_6117,N_5764,N_5685);
and U6118 (N_6118,N_4920,N_5100);
or U6119 (N_6119,N_5673,N_5528);
nand U6120 (N_6120,N_4338,N_4919);
or U6121 (N_6121,N_4441,N_4032);
or U6122 (N_6122,N_4985,N_5097);
and U6123 (N_6123,N_4558,N_5719);
and U6124 (N_6124,N_4591,N_4442);
nand U6125 (N_6125,N_4701,N_4805);
or U6126 (N_6126,N_4942,N_4733);
nor U6127 (N_6127,N_4624,N_4675);
nand U6128 (N_6128,N_4195,N_4940);
nand U6129 (N_6129,N_4300,N_4574);
nor U6130 (N_6130,N_5355,N_4280);
and U6131 (N_6131,N_5066,N_4156);
or U6132 (N_6132,N_5361,N_4547);
nand U6133 (N_6133,N_5487,N_5852);
or U6134 (N_6134,N_5913,N_5966);
nor U6135 (N_6135,N_4537,N_4048);
or U6136 (N_6136,N_4877,N_5369);
nand U6137 (N_6137,N_5907,N_4307);
nor U6138 (N_6138,N_4576,N_4346);
or U6139 (N_6139,N_5770,N_5297);
nor U6140 (N_6140,N_4914,N_4118);
and U6141 (N_6141,N_4952,N_4313);
and U6142 (N_6142,N_4120,N_5861);
or U6143 (N_6143,N_4428,N_5841);
or U6144 (N_6144,N_5925,N_4608);
or U6145 (N_6145,N_5020,N_4674);
and U6146 (N_6146,N_5229,N_5425);
nor U6147 (N_6147,N_4256,N_4884);
and U6148 (N_6148,N_4355,N_5738);
nor U6149 (N_6149,N_5943,N_4187);
nor U6150 (N_6150,N_5183,N_5073);
and U6151 (N_6151,N_5223,N_4456);
and U6152 (N_6152,N_4597,N_4924);
or U6153 (N_6153,N_4035,N_4486);
or U6154 (N_6154,N_5558,N_4415);
or U6155 (N_6155,N_4318,N_4396);
nand U6156 (N_6156,N_4105,N_4296);
nand U6157 (N_6157,N_4699,N_4757);
nand U6158 (N_6158,N_5165,N_5734);
nor U6159 (N_6159,N_5116,N_5978);
nor U6160 (N_6160,N_5396,N_4452);
nand U6161 (N_6161,N_5431,N_5878);
or U6162 (N_6162,N_5093,N_5277);
and U6163 (N_6163,N_5417,N_5248);
or U6164 (N_6164,N_4218,N_4475);
nor U6165 (N_6165,N_4841,N_4412);
or U6166 (N_6166,N_4262,N_5195);
nor U6167 (N_6167,N_5036,N_5393);
nor U6168 (N_6168,N_5967,N_5917);
or U6169 (N_6169,N_5394,N_4888);
nand U6170 (N_6170,N_5768,N_4729);
or U6171 (N_6171,N_5163,N_5622);
nand U6172 (N_6172,N_5351,N_4813);
or U6173 (N_6173,N_5224,N_5287);
and U6174 (N_6174,N_4332,N_5781);
nand U6175 (N_6175,N_5214,N_4835);
nor U6176 (N_6176,N_4374,N_4948);
or U6177 (N_6177,N_4088,N_5515);
nor U6178 (N_6178,N_5040,N_5688);
or U6179 (N_6179,N_4859,N_5960);
nor U6180 (N_6180,N_4477,N_5552);
nor U6181 (N_6181,N_4593,N_5291);
and U6182 (N_6182,N_5578,N_4246);
or U6183 (N_6183,N_5847,N_5821);
and U6184 (N_6184,N_4764,N_4728);
or U6185 (N_6185,N_4447,N_5362);
nor U6186 (N_6186,N_4774,N_4494);
and U6187 (N_6187,N_5780,N_4661);
nand U6188 (N_6188,N_5250,N_4506);
nand U6189 (N_6189,N_5241,N_5687);
and U6190 (N_6190,N_5347,N_5419);
and U6191 (N_6191,N_5359,N_5906);
nand U6192 (N_6192,N_5550,N_5077);
and U6193 (N_6193,N_4197,N_4207);
nor U6194 (N_6194,N_5415,N_4736);
nand U6195 (N_6195,N_5348,N_5111);
or U6196 (N_6196,N_5771,N_5334);
or U6197 (N_6197,N_4270,N_5496);
nor U6198 (N_6198,N_5833,N_5305);
nor U6199 (N_6199,N_5076,N_4302);
or U6200 (N_6200,N_4658,N_4389);
nor U6201 (N_6201,N_4806,N_5041);
xor U6202 (N_6202,N_5030,N_5999);
and U6203 (N_6203,N_4259,N_4020);
or U6204 (N_6204,N_5587,N_4692);
and U6205 (N_6205,N_5923,N_5125);
and U6206 (N_6206,N_4777,N_4828);
nand U6207 (N_6207,N_5412,N_4983);
nand U6208 (N_6208,N_5226,N_5518);
or U6209 (N_6209,N_5270,N_5918);
nand U6210 (N_6210,N_4050,N_5261);
xor U6211 (N_6211,N_4975,N_4264);
nand U6212 (N_6212,N_5743,N_4802);
nand U6213 (N_6213,N_4632,N_5682);
nor U6214 (N_6214,N_4178,N_4876);
and U6215 (N_6215,N_4663,N_5629);
xor U6216 (N_6216,N_5953,N_5732);
nor U6217 (N_6217,N_5479,N_5254);
nand U6218 (N_6218,N_5464,N_5538);
nor U6219 (N_6219,N_4273,N_5338);
nand U6220 (N_6220,N_4798,N_4936);
nand U6221 (N_6221,N_4765,N_4421);
nor U6222 (N_6222,N_4445,N_4610);
nor U6223 (N_6223,N_4184,N_5445);
nand U6224 (N_6224,N_5897,N_5726);
or U6225 (N_6225,N_4029,N_5542);
or U6226 (N_6226,N_5851,N_5310);
and U6227 (N_6227,N_4315,N_5300);
nor U6228 (N_6228,N_5104,N_5790);
or U6229 (N_6229,N_5798,N_4304);
nand U6230 (N_6230,N_4808,N_4769);
and U6231 (N_6231,N_5500,N_4606);
or U6232 (N_6232,N_4213,N_5171);
and U6233 (N_6233,N_4397,N_4267);
nor U6234 (N_6234,N_5367,N_4559);
nand U6235 (N_6235,N_4329,N_4536);
nand U6236 (N_6236,N_5669,N_4770);
or U6237 (N_6237,N_4375,N_4935);
nor U6238 (N_6238,N_5271,N_5474);
or U6239 (N_6239,N_4125,N_5186);
and U6240 (N_6240,N_5932,N_4846);
nand U6241 (N_6241,N_5007,N_5748);
or U6242 (N_6242,N_5689,N_4906);
xor U6243 (N_6243,N_5440,N_4164);
nand U6244 (N_6244,N_4023,N_5366);
or U6245 (N_6245,N_4394,N_4731);
xor U6246 (N_6246,N_5994,N_5634);
or U6247 (N_6247,N_5447,N_4492);
and U6248 (N_6248,N_5707,N_4311);
nor U6249 (N_6249,N_4185,N_4897);
or U6250 (N_6250,N_5900,N_4104);
nor U6251 (N_6251,N_5705,N_4843);
and U6252 (N_6252,N_4279,N_5674);
or U6253 (N_6253,N_5399,N_5581);
nand U6254 (N_6254,N_4660,N_5547);
xor U6255 (N_6255,N_4875,N_4932);
or U6256 (N_6256,N_5295,N_5830);
and U6257 (N_6257,N_4143,N_4966);
nand U6258 (N_6258,N_5446,N_4697);
nor U6259 (N_6259,N_5976,N_5233);
nand U6260 (N_6260,N_4823,N_4040);
nor U6261 (N_6261,N_5956,N_5374);
nor U6262 (N_6262,N_5267,N_4372);
nor U6263 (N_6263,N_4014,N_5845);
or U6264 (N_6264,N_5647,N_4783);
and U6265 (N_6265,N_5021,N_4766);
and U6266 (N_6266,N_4585,N_5262);
nand U6267 (N_6267,N_4672,N_5889);
or U6268 (N_6268,N_4101,N_4349);
nand U6269 (N_6269,N_4545,N_5071);
and U6270 (N_6270,N_5909,N_4106);
nand U6271 (N_6271,N_5627,N_4947);
nor U6272 (N_6272,N_5946,N_4570);
and U6273 (N_6273,N_4226,N_5680);
or U6274 (N_6274,N_5784,N_4782);
or U6275 (N_6275,N_4758,N_4664);
xor U6276 (N_6276,N_5324,N_4721);
or U6277 (N_6277,N_5624,N_4037);
nor U6278 (N_6278,N_5118,N_5709);
nor U6279 (N_6279,N_5441,N_5857);
nor U6280 (N_6280,N_5931,N_5988);
nor U6281 (N_6281,N_5009,N_4882);
nor U6282 (N_6282,N_4044,N_4093);
and U6283 (N_6283,N_4607,N_5846);
nor U6284 (N_6284,N_5782,N_5012);
nand U6285 (N_6285,N_5915,N_4189);
nand U6286 (N_6286,N_4630,N_4179);
nor U6287 (N_6287,N_4123,N_4058);
nor U6288 (N_6288,N_4840,N_5375);
and U6289 (N_6289,N_5875,N_5941);
and U6290 (N_6290,N_5757,N_4916);
and U6291 (N_6291,N_5502,N_5029);
and U6292 (N_6292,N_5736,N_4520);
or U6293 (N_6293,N_5794,N_5105);
nand U6294 (N_6294,N_5828,N_4679);
and U6295 (N_6295,N_5035,N_5237);
nand U6296 (N_6296,N_5874,N_5034);
and U6297 (N_6297,N_5207,N_5044);
nor U6298 (N_6298,N_5365,N_4698);
or U6299 (N_6299,N_5549,N_4152);
nor U6300 (N_6300,N_5590,N_5606);
nand U6301 (N_6301,N_4357,N_5196);
and U6302 (N_6302,N_4834,N_4742);
nand U6303 (N_6303,N_5660,N_5723);
and U6304 (N_6304,N_5714,N_5058);
or U6305 (N_6305,N_5488,N_5197);
nand U6306 (N_6306,N_4976,N_4437);
and U6307 (N_6307,N_4931,N_4480);
or U6308 (N_6308,N_4609,N_4933);
nor U6309 (N_6309,N_4098,N_5323);
or U6310 (N_6310,N_4361,N_4398);
and U6311 (N_6311,N_4688,N_4637);
nand U6312 (N_6312,N_5408,N_5973);
and U6313 (N_6313,N_4167,N_4416);
and U6314 (N_6314,N_5933,N_5056);
and U6315 (N_6315,N_5801,N_4850);
nor U6316 (N_6316,N_5936,N_4248);
and U6317 (N_6317,N_5921,N_5944);
and U6318 (N_6318,N_4781,N_4378);
and U6319 (N_6319,N_4388,N_5045);
or U6320 (N_6320,N_4517,N_5553);
and U6321 (N_6321,N_4013,N_4027);
or U6322 (N_6322,N_5373,N_4644);
or U6323 (N_6323,N_4130,N_5403);
nor U6324 (N_6324,N_5026,N_5540);
and U6325 (N_6325,N_5054,N_5713);
or U6326 (N_6326,N_4553,N_4508);
and U6327 (N_6327,N_5667,N_4586);
nand U6328 (N_6328,N_4481,N_4513);
nand U6329 (N_6329,N_4096,N_5424);
nor U6330 (N_6330,N_4974,N_4278);
and U6331 (N_6331,N_4419,N_4260);
or U6332 (N_6332,N_5582,N_5974);
nand U6333 (N_6333,N_5683,N_4497);
nand U6334 (N_6334,N_4271,N_5825);
nand U6335 (N_6335,N_5703,N_4668);
nand U6336 (N_6336,N_5059,N_4293);
nand U6337 (N_6337,N_5621,N_5011);
and U6338 (N_6338,N_5473,N_5456);
or U6339 (N_6339,N_5597,N_4622);
and U6340 (N_6340,N_4002,N_5354);
nand U6341 (N_6341,N_5389,N_4371);
or U6342 (N_6342,N_5676,N_5599);
nor U6343 (N_6343,N_4190,N_4431);
nor U6344 (N_6344,N_5565,N_4581);
and U6345 (N_6345,N_5759,N_4030);
and U6346 (N_6346,N_5551,N_4842);
or U6347 (N_6347,N_4786,N_4112);
or U6348 (N_6348,N_5372,N_5126);
and U6349 (N_6349,N_4380,N_5524);
nand U6350 (N_6350,N_4064,N_5371);
nor U6351 (N_6351,N_5692,N_4286);
nor U6352 (N_6352,N_5855,N_4969);
nor U6353 (N_6353,N_4204,N_5958);
or U6354 (N_6354,N_4538,N_4909);
and U6355 (N_6355,N_4703,N_4725);
nor U6356 (N_6356,N_4444,N_5724);
or U6357 (N_6357,N_5145,N_5213);
nor U6358 (N_6358,N_4827,N_5755);
nor U6359 (N_6359,N_4100,N_5422);
or U6360 (N_6360,N_5307,N_4589);
or U6361 (N_6361,N_5469,N_5509);
nor U6362 (N_6362,N_4458,N_5761);
and U6363 (N_6363,N_5131,N_5471);
nand U6364 (N_6364,N_5879,N_4904);
nand U6365 (N_6365,N_5345,N_5842);
nand U6366 (N_6366,N_5832,N_5646);
nand U6367 (N_6367,N_4234,N_4899);
xor U6368 (N_6368,N_5843,N_4963);
nor U6369 (N_6369,N_5443,N_4639);
and U6370 (N_6370,N_5448,N_5763);
or U6371 (N_6371,N_4611,N_5939);
nand U6372 (N_6372,N_4479,N_4551);
nand U6373 (N_6373,N_4788,N_4964);
and U6374 (N_6374,N_5972,N_4730);
nand U6375 (N_6375,N_4676,N_4723);
nand U6376 (N_6376,N_5677,N_5867);
nand U6377 (N_6377,N_4347,N_4141);
or U6378 (N_6378,N_5008,N_4244);
or U6379 (N_6379,N_5164,N_4670);
nand U6380 (N_6380,N_4571,N_4979);
or U6381 (N_6381,N_4053,N_5799);
nor U6382 (N_6382,N_5256,N_4085);
and U6383 (N_6383,N_4060,N_5639);
or U6384 (N_6384,N_5525,N_4124);
nand U6385 (N_6385,N_5911,N_4554);
nand U6386 (N_6386,N_5809,N_5302);
nor U6387 (N_6387,N_5598,N_5096);
or U6388 (N_6388,N_5352,N_5554);
nor U6389 (N_6389,N_4087,N_4299);
and U6390 (N_6390,N_5212,N_5762);
or U6391 (N_6391,N_5672,N_5577);
and U6392 (N_6392,N_4405,N_4327);
or U6393 (N_6393,N_4321,N_4134);
and U6394 (N_6394,N_5839,N_5142);
nand U6395 (N_6395,N_5243,N_4986);
and U6396 (N_6396,N_5740,N_4323);
or U6397 (N_6397,N_4031,N_4155);
nor U6398 (N_6398,N_5864,N_4400);
nand U6399 (N_6399,N_5823,N_4747);
nor U6400 (N_6400,N_4116,N_4792);
nor U6401 (N_6401,N_5733,N_5379);
or U6402 (N_6402,N_4268,N_5548);
nand U6403 (N_6403,N_5468,N_4126);
and U6404 (N_6404,N_4075,N_5998);
nand U6405 (N_6405,N_5113,N_4890);
nand U6406 (N_6406,N_4510,N_4634);
and U6407 (N_6407,N_4094,N_5700);
or U6408 (N_6408,N_4540,N_5109);
nor U6409 (N_6409,N_5592,N_4176);
or U6410 (N_6410,N_5148,N_5783);
nand U6411 (N_6411,N_5311,N_4006);
and U6412 (N_6412,N_4157,N_4839);
and U6413 (N_6413,N_5025,N_4181);
and U6414 (N_6414,N_4076,N_5033);
or U6415 (N_6415,N_5750,N_5916);
nor U6416 (N_6416,N_4773,N_4775);
and U6417 (N_6417,N_4292,N_4325);
and U6418 (N_6418,N_4898,N_4242);
and U6419 (N_6419,N_4122,N_4072);
or U6420 (N_6420,N_5306,N_4694);
or U6421 (N_6421,N_5153,N_5078);
nand U6422 (N_6422,N_4426,N_5979);
nand U6423 (N_6423,N_5172,N_4366);
or U6424 (N_6424,N_5234,N_4838);
and U6425 (N_6425,N_5491,N_5064);
or U6426 (N_6426,N_5122,N_4505);
nor U6427 (N_6427,N_4917,N_4722);
nor U6428 (N_6428,N_5517,N_5249);
and U6429 (N_6429,N_4026,N_5264);
and U6430 (N_6430,N_4034,N_4407);
or U6431 (N_6431,N_5503,N_5579);
nand U6432 (N_6432,N_4521,N_4727);
or U6433 (N_6433,N_5115,N_5152);
or U6434 (N_6434,N_5633,N_4082);
nand U6435 (N_6435,N_5173,N_4312);
nor U6436 (N_6436,N_4950,N_5704);
nor U6437 (N_6437,N_5178,N_5957);
nor U6438 (N_6438,N_4414,N_4831);
nor U6439 (N_6439,N_5278,N_5912);
nor U6440 (N_6440,N_4393,N_5028);
or U6441 (N_6441,N_4133,N_4005);
nand U6442 (N_6442,N_5511,N_4140);
nand U6443 (N_6443,N_4620,N_5555);
and U6444 (N_6444,N_4057,N_5370);
or U6445 (N_6445,N_5678,N_4797);
nor U6446 (N_6446,N_5258,N_4762);
and U6447 (N_6447,N_4780,N_5626);
nand U6448 (N_6448,N_4998,N_5948);
and U6449 (N_6449,N_4874,N_4651);
and U6450 (N_6450,N_4922,N_5559);
xor U6451 (N_6451,N_4272,N_4810);
and U6452 (N_6452,N_5039,N_4641);
nor U6453 (N_6453,N_5092,N_5981);
nand U6454 (N_6454,N_4223,N_5315);
nor U6455 (N_6455,N_5060,N_5791);
and U6456 (N_6456,N_5708,N_4217);
nor U6457 (N_6457,N_4601,N_4219);
and U6458 (N_6458,N_5971,N_5760);
or U6459 (N_6459,N_4789,N_4794);
and U6460 (N_6460,N_4744,N_4512);
nand U6461 (N_6461,N_4056,N_4605);
or U6462 (N_6462,N_4343,N_5260);
or U6463 (N_6463,N_4873,N_4091);
nor U6464 (N_6464,N_5863,N_5463);
or U6465 (N_6465,N_5860,N_5720);
or U6466 (N_6466,N_5573,N_5466);
nor U6467 (N_6467,N_4149,N_4577);
nand U6468 (N_6468,N_5866,N_5534);
and U6469 (N_6469,N_4636,N_4073);
and U6470 (N_6470,N_5032,N_5144);
nor U6471 (N_6471,N_4269,N_4049);
and U6472 (N_6472,N_5896,N_5385);
or U6473 (N_6473,N_5568,N_5610);
and U6474 (N_6474,N_4791,N_5426);
nand U6475 (N_6475,N_5747,N_5670);
and U6476 (N_6476,N_5288,N_5363);
or U6477 (N_6477,N_5495,N_4161);
or U6478 (N_6478,N_4117,N_5519);
nand U6479 (N_6479,N_4448,N_4981);
nand U6480 (N_6480,N_5596,N_4151);
and U6481 (N_6481,N_4113,N_5872);
and U6482 (N_6482,N_4295,N_4449);
and U6483 (N_6483,N_4618,N_5569);
and U6484 (N_6484,N_4530,N_4755);
and U6485 (N_6485,N_5952,N_5774);
or U6486 (N_6486,N_5483,N_5880);
or U6487 (N_6487,N_5869,N_5410);
nand U6488 (N_6488,N_4159,N_5820);
or U6489 (N_6489,N_4180,N_5314);
or U6490 (N_6490,N_5557,N_4196);
nor U6491 (N_6491,N_5220,N_4543);
nand U6492 (N_6492,N_4487,N_5150);
or U6493 (N_6493,N_5119,N_4763);
nand U6494 (N_6494,N_4352,N_4710);
nor U6495 (N_6495,N_4089,N_5376);
or U6496 (N_6496,N_5608,N_5072);
nand U6497 (N_6497,N_4364,N_4422);
and U6498 (N_6498,N_5758,N_5068);
nor U6499 (N_6499,N_4615,N_5992);
nand U6500 (N_6500,N_4462,N_5461);
and U6501 (N_6501,N_4348,N_4741);
nand U6502 (N_6502,N_5478,N_4800);
and U6503 (N_6503,N_4531,N_4424);
or U6504 (N_6504,N_5902,N_4045);
or U6505 (N_6505,N_4944,N_4552);
nand U6506 (N_6506,N_4229,N_4750);
nand U6507 (N_6507,N_4466,N_5247);
and U6508 (N_6508,N_5642,N_5831);
nand U6509 (N_6509,N_4102,N_5227);
or U6510 (N_6510,N_5494,N_4956);
or U6511 (N_6511,N_5859,N_4379);
nand U6512 (N_6512,N_5652,N_5206);
or U6513 (N_6513,N_5792,N_5467);
nand U6514 (N_6514,N_4358,N_4569);
or U6515 (N_6515,N_5501,N_4519);
or U6516 (N_6516,N_4493,N_5174);
nand U6517 (N_6517,N_4930,N_5567);
nand U6518 (N_6518,N_5387,N_5193);
nand U6519 (N_6519,N_5342,N_5344);
nor U6520 (N_6520,N_4224,N_4640);
nor U6521 (N_6521,N_4127,N_5405);
nor U6522 (N_6522,N_5308,N_5562);
nand U6523 (N_6523,N_4353,N_5537);
or U6524 (N_6524,N_5838,N_4851);
nor U6525 (N_6525,N_4713,N_4700);
nor U6526 (N_6526,N_4907,N_4685);
nand U6527 (N_6527,N_5452,N_5147);
nor U6528 (N_6528,N_4362,N_4858);
and U6529 (N_6529,N_4438,N_5080);
nand U6530 (N_6530,N_4960,N_5625);
or U6531 (N_6531,N_5816,N_5533);
or U6532 (N_6532,N_5745,N_5442);
and U6533 (N_6533,N_5018,N_4712);
nand U6534 (N_6534,N_4539,N_4804);
nor U6535 (N_6535,N_4820,N_5121);
nand U6536 (N_6536,N_4836,N_4186);
nand U6537 (N_6537,N_4665,N_5788);
nand U6538 (N_6538,N_4172,N_5435);
and U6539 (N_6539,N_5922,N_5886);
or U6540 (N_6540,N_4991,N_4291);
or U6541 (N_6541,N_5103,N_4467);
and U6542 (N_6542,N_5343,N_4790);
nand U6543 (N_6543,N_5914,N_4095);
and U6544 (N_6544,N_4135,N_4250);
and U6545 (N_6545,N_5053,N_5027);
and U6546 (N_6546,N_4383,N_5655);
nor U6547 (N_6547,N_4137,N_5749);
nand U6548 (N_6548,N_4097,N_4170);
nand U6549 (N_6549,N_4844,N_5330);
nand U6550 (N_6550,N_5280,N_5166);
nor U6551 (N_6551,N_4033,N_5881);
or U6552 (N_6552,N_4619,N_5459);
and U6553 (N_6553,N_4659,N_4623);
and U6554 (N_6554,N_5901,N_4621);
nor U6555 (N_6555,N_5870,N_4815);
nor U6556 (N_6556,N_5827,N_5023);
or U6557 (N_6557,N_5717,N_4696);
and U6558 (N_6558,N_5048,N_4435);
nor U6559 (N_6559,N_4128,N_5349);
nor U6560 (N_6560,N_5458,N_5808);
and U6561 (N_6561,N_4826,N_5380);
and U6562 (N_6562,N_4344,N_5604);
or U6563 (N_6563,N_4305,N_5110);
nor U6564 (N_6564,N_5199,N_5438);
nor U6565 (N_6565,N_5942,N_4678);
or U6566 (N_6566,N_4913,N_5665);
or U6567 (N_6567,N_5482,N_5492);
nor U6568 (N_6568,N_4216,N_4961);
and U6569 (N_6569,N_4565,N_4498);
nor U6570 (N_6570,N_5046,N_4937);
nor U6571 (N_6571,N_4495,N_5228);
or U6572 (N_6572,N_4590,N_4483);
or U6573 (N_6573,N_4402,N_4684);
nand U6574 (N_6574,N_5485,N_4328);
and U6575 (N_6575,N_5134,N_5583);
nor U6576 (N_6576,N_4911,N_5619);
nor U6577 (N_6577,N_4816,N_5133);
nor U6578 (N_6578,N_5225,N_5182);
or U6579 (N_6579,N_4499,N_4997);
or U6580 (N_6580,N_4572,N_5416);
nor U6581 (N_6581,N_4885,N_5919);
nor U6582 (N_6582,N_4643,N_5572);
nand U6583 (N_6583,N_4681,N_5613);
or U6584 (N_6584,N_5014,N_4999);
nand U6585 (N_6585,N_5003,N_5789);
xor U6586 (N_6586,N_5997,N_5698);
nor U6587 (N_6587,N_5806,N_5364);
or U6588 (N_6588,N_4276,N_4024);
or U6589 (N_6589,N_4912,N_5836);
and U6590 (N_6590,N_5814,N_5541);
and U6591 (N_6591,N_4069,N_4047);
and U6592 (N_6592,N_5303,N_5187);
nor U6593 (N_6593,N_5591,N_5699);
or U6594 (N_6594,N_5871,N_5418);
nor U6595 (N_6595,N_4003,N_5336);
and U6596 (N_6596,N_4753,N_4772);
xor U6597 (N_6597,N_5593,N_4342);
nor U6598 (N_6598,N_5849,N_5694);
nor U6599 (N_6599,N_5019,N_4923);
and U6600 (N_6600,N_5242,N_5804);
and U6601 (N_6601,N_4339,N_4427);
nor U6602 (N_6602,N_5584,N_4957);
or U6603 (N_6603,N_5850,N_4046);
and U6604 (N_6604,N_5527,N_4274);
nand U6605 (N_6605,N_4896,N_5340);
nor U6606 (N_6606,N_5455,N_5602);
and U6607 (N_6607,N_5211,N_5273);
and U6608 (N_6608,N_4654,N_4454);
or U6609 (N_6609,N_4436,N_5335);
nor U6610 (N_6610,N_5252,N_4993);
or U6611 (N_6611,N_4946,N_4074);
or U6612 (N_6612,N_4166,N_4847);
or U6613 (N_6613,N_4596,N_4258);
nor U6614 (N_6614,N_4592,N_5560);
and U6615 (N_6615,N_4025,N_4376);
nor U6616 (N_6616,N_4142,N_4990);
and U6617 (N_6617,N_5084,N_4211);
nor U6618 (N_6618,N_4954,N_4261);
and U6619 (N_6619,N_5628,N_5177);
and U6620 (N_6620,N_4107,N_5635);
nor U6621 (N_6621,N_5854,N_4215);
or U6622 (N_6622,N_5114,N_5545);
or U6623 (N_6623,N_5159,N_4210);
and U6624 (N_6624,N_5038,N_4707);
nand U6625 (N_6625,N_4953,N_5595);
and U6626 (N_6626,N_4208,N_4285);
or U6627 (N_6627,N_4550,N_5991);
and U6628 (N_6628,N_4334,N_5218);
nor U6629 (N_6629,N_5413,N_4776);
or U6630 (N_6630,N_4232,N_5498);
or U6631 (N_6631,N_5965,N_5155);
and U6632 (N_6632,N_5730,N_4488);
nor U6633 (N_6633,N_4175,N_4724);
or U6634 (N_6634,N_4485,N_4852);
nand U6635 (N_6635,N_5317,N_4169);
and U6636 (N_6636,N_5510,N_5411);
or U6637 (N_6637,N_4450,N_5883);
nand U6638 (N_6638,N_4647,N_4459);
or U6639 (N_6639,N_5061,N_5654);
nand U6640 (N_6640,N_5504,N_5607);
nand U6641 (N_6641,N_5844,N_5384);
nor U6642 (N_6642,N_5520,N_4695);
nand U6643 (N_6643,N_5951,N_5643);
and U6644 (N_6644,N_4735,N_4059);
or U6645 (N_6645,N_4984,N_4532);
nand U6646 (N_6646,N_4529,N_5437);
nor U6647 (N_6647,N_4600,N_4915);
or U6648 (N_6648,N_5157,N_5090);
nor U6649 (N_6649,N_5099,N_4473);
nor U6650 (N_6650,N_4301,N_4967);
and U6651 (N_6651,N_4929,N_5817);
or U6652 (N_6652,N_5219,N_4887);
or U6653 (N_6653,N_5588,N_4555);
nor U6654 (N_6654,N_4927,N_4734);
or U6655 (N_6655,N_4282,N_5318);
nand U6656 (N_6656,N_4680,N_5938);
nand U6657 (N_6657,N_5000,N_5807);
and U6658 (N_6658,N_4423,N_4862);
and U6659 (N_6659,N_5127,N_5955);
and U6660 (N_6660,N_5244,N_5292);
nand U6661 (N_6661,N_5433,N_4115);
nand U6662 (N_6662,N_5480,N_5508);
or U6663 (N_6663,N_5235,N_5744);
or U6664 (N_6664,N_4617,N_5246);
and U6665 (N_6665,N_5924,N_4503);
or U6666 (N_6666,N_4001,N_5050);
and U6667 (N_6667,N_4413,N_5210);
or U6668 (N_6668,N_4941,N_5803);
or U6669 (N_6669,N_5802,N_4021);
nand U6670 (N_6670,N_5521,N_4871);
and U6671 (N_6671,N_5522,N_5930);
or U6672 (N_6672,N_5493,N_5255);
and U6673 (N_6673,N_4653,N_5645);
or U6674 (N_6674,N_4038,N_5325);
or U6675 (N_6675,N_4548,N_5010);
and U6676 (N_6676,N_4996,N_4147);
or U6677 (N_6677,N_5130,N_4042);
nand U6678 (N_6678,N_4926,N_5543);
nor U6679 (N_6679,N_4228,N_4320);
or U6680 (N_6680,N_4959,N_5083);
nor U6681 (N_6681,N_4598,N_4194);
nand U6682 (N_6682,N_4465,N_5776);
nor U6683 (N_6683,N_5263,N_5996);
nand U6684 (N_6684,N_4257,N_5656);
or U6685 (N_6685,N_4469,N_4205);
or U6686 (N_6686,N_4225,N_4970);
nand U6687 (N_6687,N_5322,N_4849);
nand U6688 (N_6688,N_4066,N_4198);
and U6689 (N_6689,N_5767,N_4677);
and U6690 (N_6690,N_4350,N_4631);
and U6691 (N_6691,N_4645,N_5117);
and U6692 (N_6692,N_4368,N_4287);
or U6693 (N_6693,N_4252,N_5350);
nand U6694 (N_6694,N_5279,N_5532);
and U6695 (N_6695,N_4284,N_4404);
nand U6696 (N_6696,N_4642,N_4434);
and U6697 (N_6697,N_5427,N_4410);
nand U6698 (N_6698,N_5331,N_5128);
and U6699 (N_6699,N_4666,N_5269);
nor U6700 (N_6700,N_4154,N_5544);
or U6701 (N_6701,N_4627,N_5085);
xor U6702 (N_6702,N_5299,N_4702);
nand U6703 (N_6703,N_4241,N_4036);
nor U6704 (N_6704,N_5853,N_4943);
or U6705 (N_6705,N_4432,N_5600);
and U6706 (N_6706,N_5769,N_4322);
nor U6707 (N_6707,N_5304,N_5785);
or U6708 (N_6708,N_4977,N_4525);
nor U6709 (N_6709,N_5276,N_4290);
or U6710 (N_6710,N_4359,N_4582);
and U6711 (N_6711,N_4333,N_4331);
nand U6712 (N_6712,N_5188,N_4114);
or U6713 (N_6713,N_4309,N_4471);
or U6714 (N_6714,N_5284,N_4153);
nand U6715 (N_6715,N_4227,N_5216);
or U6716 (N_6716,N_5095,N_4417);
nor U6717 (N_6717,N_5890,N_4240);
or U6718 (N_6718,N_5378,N_4491);
nor U6719 (N_6719,N_5977,N_4080);
or U6720 (N_6720,N_4534,N_5239);
nand U6721 (N_6721,N_4635,N_5696);
or U6722 (N_6722,N_5070,N_5848);
nand U6723 (N_6723,N_5191,N_4384);
nor U6724 (N_6724,N_4235,N_5390);
nor U6725 (N_6725,N_5618,N_5232);
or U6726 (N_6726,N_4403,N_5735);
and U6727 (N_6727,N_4065,N_5753);
or U6728 (N_6728,N_4895,N_5751);
nor U6729 (N_6729,N_4377,N_4752);
nand U6730 (N_6730,N_5470,N_4796);
and U6731 (N_6731,N_4337,N_5691);
nor U6732 (N_6732,N_4955,N_5245);
xor U6733 (N_6733,N_4370,N_4901);
nor U6734 (N_6734,N_5731,N_4691);
nand U6735 (N_6735,N_5404,N_4787);
and U6736 (N_6736,N_5611,N_5891);
nor U6737 (N_6737,N_4962,N_5795);
nand U6738 (N_6738,N_5002,N_4288);
and U6739 (N_6739,N_4893,N_4324);
nor U6740 (N_6740,N_5840,N_5895);
nand U6741 (N_6741,N_5935,N_4004);
nor U6742 (N_6742,N_4511,N_5516);
or U6743 (N_6743,N_5112,N_5140);
nor U6744 (N_6744,N_5986,N_5190);
or U6745 (N_6745,N_5460,N_4132);
nor U6746 (N_6746,N_4878,N_5862);
nand U6747 (N_6747,N_5161,N_5638);
nor U6748 (N_6748,N_5414,N_5309);
and U6749 (N_6749,N_5585,N_5203);
or U6750 (N_6750,N_4938,N_5184);
and U6751 (N_6751,N_4243,N_5423);
or U6752 (N_6752,N_4507,N_5787);
or U6753 (N_6753,N_5800,N_4062);
nor U6754 (N_6754,N_4446,N_5169);
nor U6755 (N_6755,N_4382,N_5253);
nor U6756 (N_6756,N_5746,N_5920);
and U6757 (N_6757,N_5200,N_5586);
or U6758 (N_6758,N_5160,N_5088);
nand U6759 (N_6759,N_5649,N_5984);
nand U6760 (N_6760,N_5648,N_4793);
or U6761 (N_6761,N_5499,N_4411);
nand U6762 (N_6762,N_5903,N_4000);
and U6763 (N_6763,N_5739,N_5063);
nand U6764 (N_6764,N_4297,N_4992);
nor U6765 (N_6765,N_4704,N_4054);
nand U6766 (N_6766,N_5170,N_5711);
and U6767 (N_6767,N_4908,N_5813);
and U6768 (N_6768,N_4795,N_5194);
and U6769 (N_6769,N_5429,N_5824);
and U6770 (N_6770,N_4921,N_4263);
nand U6771 (N_6771,N_5885,N_4010);
or U6772 (N_6772,N_4533,N_4657);
or U6773 (N_6773,N_4206,N_4801);
nor U6774 (N_6774,N_4509,N_5436);
and U6775 (N_6775,N_5420,N_4594);
nor U6776 (N_6776,N_4894,N_5980);
nand U6777 (N_6777,N_5141,N_4546);
nor U6778 (N_6778,N_4433,N_4756);
and U6779 (N_6779,N_5031,N_4360);
and U6780 (N_6780,N_5067,N_5664);
nand U6781 (N_6781,N_5888,N_4706);
and U6782 (N_6782,N_4109,N_4245);
or U6783 (N_6783,N_4903,N_4430);
nand U6784 (N_6784,N_5326,N_4504);
and U6785 (N_6785,N_5929,N_4386);
nor U6786 (N_6786,N_5395,N_5826);
and U6787 (N_6787,N_4673,N_5146);
or U6788 (N_6788,N_4478,N_5796);
or U6789 (N_6789,N_4200,N_5451);
nand U6790 (N_6790,N_5337,N_4008);
nand U6791 (N_6791,N_5055,N_5236);
nor U6792 (N_6792,N_5043,N_5679);
and U6793 (N_6793,N_4855,N_4515);
nand U6794 (N_6794,N_4595,N_5811);
xnor U6795 (N_6795,N_5514,N_5765);
or U6796 (N_6796,N_5017,N_5818);
or U6797 (N_6797,N_5576,N_4182);
or U6798 (N_6798,N_5081,N_4496);
or U6799 (N_6799,N_4314,N_4575);
or U6800 (N_6800,N_4174,N_4121);
or U6801 (N_6801,N_5240,N_5728);
and U6802 (N_6802,N_4583,N_4418);
or U6803 (N_6803,N_5091,N_5274);
or U6804 (N_6804,N_4306,N_5301);
or U6805 (N_6805,N_4629,N_5022);
nand U6806 (N_6806,N_5386,N_5434);
nand U6807 (N_6807,N_5877,N_5754);
or U6808 (N_6808,N_4872,N_4401);
nand U6809 (N_6809,N_5231,N_5074);
or U6810 (N_6810,N_4561,N_5001);
and U6811 (N_6811,N_4474,N_4918);
nand U6812 (N_6812,N_4007,N_4599);
nor U6813 (N_6813,N_4516,N_5321);
nor U6814 (N_6814,N_5894,N_5819);
nand U6815 (N_6815,N_5087,N_5637);
nand U6816 (N_6816,N_4683,N_5407);
nand U6817 (N_6817,N_4891,N_4863);
and U6818 (N_6818,N_4470,N_5398);
or U6819 (N_6819,N_4866,N_4656);
and U6820 (N_6820,N_5185,N_5449);
and U6821 (N_6821,N_4638,N_5089);
or U6822 (N_6822,N_5057,N_5718);
nor U6823 (N_6823,N_5049,N_5702);
nand U6824 (N_6824,N_5208,N_5513);
and U6825 (N_6825,N_4451,N_5620);
and U6826 (N_6826,N_5697,N_4965);
nand U6827 (N_6827,N_4502,N_4051);
nor U6828 (N_6828,N_5179,N_5024);
nor U6829 (N_6829,N_5107,N_4928);
nor U6830 (N_6830,N_5662,N_5741);
nand U6831 (N_6831,N_5640,N_4761);
nand U6832 (N_6832,N_4041,N_5472);
nand U6833 (N_6833,N_4192,N_5201);
nand U6834 (N_6834,N_5316,N_5268);
and U6835 (N_6835,N_5995,N_4751);
or U6836 (N_6836,N_5961,N_4717);
and U6837 (N_6837,N_4460,N_4012);
and U6838 (N_6838,N_5727,N_5756);
nor U6839 (N_6839,N_5108,N_4718);
nor U6840 (N_6840,N_5561,N_5293);
or U6841 (N_6841,N_5512,N_4662);
or U6842 (N_6842,N_4557,N_4067);
and U6843 (N_6843,N_4867,N_5313);
or U6844 (N_6844,N_5428,N_5465);
nor U6845 (N_6845,N_5954,N_5928);
or U6846 (N_6846,N_5296,N_4856);
nor U6847 (N_6847,N_5181,N_5132);
nand U6848 (N_6848,N_4824,N_4745);
nand U6849 (N_6849,N_5574,N_4171);
nand U6850 (N_6850,N_5341,N_4222);
and U6851 (N_6851,N_4549,N_5430);
nor U6852 (N_6852,N_4392,N_4440);
nand U6853 (N_6853,N_4818,N_4484);
nand U6854 (N_6854,N_5793,N_5695);
or U6855 (N_6855,N_5722,N_4319);
and U6856 (N_6856,N_5612,N_5766);
or U6857 (N_6857,N_4011,N_4541);
and U6858 (N_6858,N_5675,N_5189);
nor U6859 (N_6859,N_5120,N_5949);
nand U6860 (N_6860,N_5462,N_5616);
nand U6861 (N_6861,N_4289,N_5778);
nand U6862 (N_6862,N_5346,N_4468);
and U6863 (N_6863,N_4982,N_4560);
nand U6864 (N_6864,N_5892,N_4310);
nand U6865 (N_6865,N_4385,N_5810);
or U6866 (N_6866,N_5630,N_5406);
nand U6867 (N_6867,N_4425,N_4860);
nor U6868 (N_6868,N_5281,N_4052);
nor U6869 (N_6869,N_5779,N_5444);
nand U6870 (N_6870,N_5668,N_5812);
or U6871 (N_6871,N_5865,N_5829);
nand U6872 (N_6872,N_5609,N_4387);
and U6873 (N_6873,N_4111,N_5614);
nor U6874 (N_6874,N_5086,N_4987);
nor U6875 (N_6875,N_5052,N_5605);
nand U6876 (N_6876,N_5013,N_4819);
nand U6877 (N_6877,N_4580,N_4714);
and U6878 (N_6878,N_4177,N_4237);
or U6879 (N_6879,N_5162,N_5453);
xor U6880 (N_6880,N_5893,N_5238);
nor U6881 (N_6881,N_4584,N_4837);
nand U6882 (N_6882,N_4682,N_4018);
and U6883 (N_6883,N_4455,N_5535);
xnor U6884 (N_6884,N_5566,N_5065);
and U6885 (N_6885,N_5969,N_4409);
and U6886 (N_6886,N_4667,N_4726);
and U6887 (N_6887,N_5123,N_5298);
and U6888 (N_6888,N_5721,N_4973);
nor U6889 (N_6889,N_4119,N_5129);
or U6890 (N_6890,N_4669,N_4399);
nor U6891 (N_6891,N_5329,N_4821);
or U6892 (N_6892,N_5388,N_4055);
nand U6893 (N_6893,N_4578,N_5712);
nand U6894 (N_6894,N_4165,N_5450);
or U6895 (N_6895,N_4341,N_4443);
nor U6896 (N_6896,N_4564,N_5042);
nor U6897 (N_6897,N_4686,N_5887);
and U6898 (N_6898,N_4785,N_5272);
nor U6899 (N_6899,N_5382,N_4199);
nand U6900 (N_6900,N_4308,N_5899);
and U6901 (N_6901,N_5047,N_5686);
nor U6902 (N_6902,N_4740,N_4209);
and U6903 (N_6903,N_5421,N_4283);
and U6904 (N_6904,N_5006,N_4749);
or U6905 (N_6905,N_4330,N_5439);
or U6906 (N_6906,N_4743,N_5476);
nor U6907 (N_6907,N_4239,N_5989);
and U6908 (N_6908,N_5082,N_5381);
or U6909 (N_6909,N_5641,N_5136);
and U6910 (N_6910,N_4563,N_4193);
nor U6911 (N_6911,N_4708,N_4129);
or U6912 (N_6912,N_5858,N_5898);
xnor U6913 (N_6913,N_4689,N_4524);
nor U6914 (N_6914,N_5623,N_5217);
nand U6915 (N_6915,N_4759,N_5312);
nand U6916 (N_6916,N_5710,N_5192);
nor U6917 (N_6917,N_4022,N_5947);
and U6918 (N_6918,N_4579,N_4811);
and U6919 (N_6919,N_5094,N_5205);
and U6920 (N_6920,N_4833,N_4231);
nand U6921 (N_6921,N_5156,N_4562);
nand U6922 (N_6922,N_4829,N_4865);
or U6923 (N_6923,N_5546,N_5402);
nand U6924 (N_6924,N_5180,N_4978);
and U6925 (N_6925,N_4160,N_5959);
and U6926 (N_6926,N_4500,N_5397);
and U6927 (N_6927,N_4604,N_5319);
nand U6928 (N_6928,N_4886,N_5822);
nor U6929 (N_6929,N_4275,N_4482);
nand U6930 (N_6930,N_5098,N_4336);
nor U6931 (N_6931,N_4183,N_4251);
or U6932 (N_6932,N_5908,N_4294);
or U6933 (N_6933,N_4613,N_5987);
nor U6934 (N_6934,N_5575,N_4544);
or U6935 (N_6935,N_5570,N_4646);
and U6936 (N_6936,N_4868,N_5603);
nand U6937 (N_6937,N_5530,N_4832);
and U6938 (N_6938,N_5563,N_4514);
nor U6939 (N_6939,N_4900,N_4784);
nand U6940 (N_6940,N_4573,N_4373);
nand U6941 (N_6941,N_4588,N_5993);
and U6942 (N_6942,N_5481,N_5975);
nor U6943 (N_6943,N_4369,N_4077);
and U6944 (N_6944,N_4203,N_5926);
or U6945 (N_6945,N_5151,N_5358);
nand U6946 (N_6946,N_4817,N_4711);
or U6947 (N_6947,N_4768,N_5432);
or U6948 (N_6948,N_5004,N_5230);
nand U6949 (N_6949,N_5671,N_4825);
and U6950 (N_6950,N_5176,N_4958);
nand U6951 (N_6951,N_5834,N_4202);
or U6952 (N_6952,N_4994,N_5497);
nand U6953 (N_6953,N_4587,N_5454);
or U6954 (N_6954,N_4709,N_5681);
nand U6955 (N_6955,N_5016,N_5139);
and U6956 (N_6956,N_5332,N_5701);
nor U6957 (N_6957,N_5328,N_4489);
and U6958 (N_6958,N_4527,N_5149);
or U6959 (N_6959,N_5392,N_5797);
nor U6960 (N_6960,N_4266,N_5835);
nand U6961 (N_6961,N_4084,N_4092);
nor U6962 (N_6962,N_4335,N_4236);
or U6963 (N_6963,N_4086,N_4139);
and U6964 (N_6964,N_4110,N_5594);
and U6965 (N_6965,N_5357,N_4633);
nand U6966 (N_6966,N_4221,N_4523);
or U6967 (N_6967,N_5716,N_5651);
or U6968 (N_6968,N_5275,N_4136);
nor U6969 (N_6969,N_5290,N_5737);
and U6970 (N_6970,N_4869,N_5409);
or U6971 (N_6971,N_4238,N_4158);
or U6972 (N_6972,N_5950,N_5401);
or U6973 (N_6973,N_5644,N_4356);
nor U6974 (N_6974,N_4168,N_5477);
nor U6975 (N_6975,N_4568,N_5571);
nand U6976 (N_6976,N_5168,N_4070);
nor U6977 (N_6977,N_4220,N_5666);
or U6978 (N_6978,N_4395,N_4626);
nand U6979 (N_6979,N_5489,N_4767);
nor U6980 (N_6980,N_5154,N_4146);
or U6981 (N_6981,N_4083,N_5289);
nor U6982 (N_6982,N_4628,N_4345);
and U6983 (N_6983,N_5285,N_5259);
nor U6984 (N_6984,N_4612,N_5658);
or U6985 (N_6985,N_4807,N_5457);
or U6986 (N_6986,N_5135,N_4934);
nand U6987 (N_6987,N_4945,N_5320);
or U6988 (N_6988,N_4902,N_4939);
nor U6989 (N_6989,N_5873,N_5333);
nor U6990 (N_6990,N_5837,N_5531);
or U6991 (N_6991,N_5539,N_4671);
nor U6992 (N_6992,N_5815,N_5529);
nor U6993 (N_6993,N_4848,N_4690);
and U6994 (N_6994,N_4648,N_4870);
nand U6995 (N_6995,N_5339,N_4017);
and U6996 (N_6996,N_4715,N_4148);
nand U6997 (N_6997,N_4910,N_4326);
and U6998 (N_6998,N_5659,N_4476);
and U6999 (N_6999,N_4457,N_4652);
or U7000 (N_7000,N_4646,N_4135);
nor U7001 (N_7001,N_4135,N_4528);
or U7002 (N_7002,N_5840,N_5013);
nand U7003 (N_7003,N_5945,N_4524);
nand U7004 (N_7004,N_4933,N_4323);
nand U7005 (N_7005,N_4340,N_4159);
or U7006 (N_7006,N_4052,N_4809);
and U7007 (N_7007,N_5420,N_4596);
and U7008 (N_7008,N_5376,N_4287);
nand U7009 (N_7009,N_5707,N_5123);
and U7010 (N_7010,N_5313,N_4211);
nand U7011 (N_7011,N_5480,N_4806);
or U7012 (N_7012,N_4679,N_5943);
or U7013 (N_7013,N_5025,N_4210);
and U7014 (N_7014,N_5608,N_5716);
xor U7015 (N_7015,N_4273,N_5308);
and U7016 (N_7016,N_4105,N_5483);
nand U7017 (N_7017,N_5043,N_5239);
and U7018 (N_7018,N_5320,N_5142);
nand U7019 (N_7019,N_4207,N_4206);
or U7020 (N_7020,N_4665,N_4650);
nand U7021 (N_7021,N_4072,N_4054);
nor U7022 (N_7022,N_4234,N_5849);
nor U7023 (N_7023,N_5051,N_5400);
or U7024 (N_7024,N_5406,N_5838);
and U7025 (N_7025,N_5732,N_4203);
nand U7026 (N_7026,N_4137,N_5616);
nand U7027 (N_7027,N_5345,N_4952);
or U7028 (N_7028,N_4192,N_5179);
nor U7029 (N_7029,N_5774,N_5009);
nor U7030 (N_7030,N_4478,N_4775);
nor U7031 (N_7031,N_4295,N_4195);
nand U7032 (N_7032,N_4486,N_5108);
or U7033 (N_7033,N_5162,N_5151);
and U7034 (N_7034,N_5914,N_5976);
or U7035 (N_7035,N_4510,N_4373);
nand U7036 (N_7036,N_5405,N_5491);
nor U7037 (N_7037,N_4506,N_4179);
or U7038 (N_7038,N_4007,N_4195);
or U7039 (N_7039,N_5948,N_4523);
or U7040 (N_7040,N_4577,N_4135);
nor U7041 (N_7041,N_4597,N_5085);
or U7042 (N_7042,N_4190,N_5602);
nor U7043 (N_7043,N_5819,N_5424);
or U7044 (N_7044,N_4438,N_5632);
and U7045 (N_7045,N_5066,N_4583);
and U7046 (N_7046,N_4765,N_4993);
nor U7047 (N_7047,N_4625,N_4853);
or U7048 (N_7048,N_4530,N_5276);
and U7049 (N_7049,N_5321,N_4767);
or U7050 (N_7050,N_5051,N_5980);
or U7051 (N_7051,N_4778,N_4935);
and U7052 (N_7052,N_4591,N_5234);
nor U7053 (N_7053,N_4000,N_4815);
and U7054 (N_7054,N_5104,N_5806);
and U7055 (N_7055,N_4263,N_5369);
and U7056 (N_7056,N_4831,N_4060);
nand U7057 (N_7057,N_4434,N_5970);
nand U7058 (N_7058,N_4972,N_5702);
and U7059 (N_7059,N_4619,N_5407);
nor U7060 (N_7060,N_5821,N_5238);
nand U7061 (N_7061,N_4361,N_5707);
nand U7062 (N_7062,N_5735,N_5033);
or U7063 (N_7063,N_5653,N_5138);
or U7064 (N_7064,N_4754,N_5896);
nand U7065 (N_7065,N_5326,N_4620);
nor U7066 (N_7066,N_5965,N_5340);
and U7067 (N_7067,N_5357,N_5197);
nor U7068 (N_7068,N_4881,N_5756);
nand U7069 (N_7069,N_5849,N_5913);
or U7070 (N_7070,N_4174,N_4062);
and U7071 (N_7071,N_4470,N_5519);
nand U7072 (N_7072,N_5052,N_5855);
nor U7073 (N_7073,N_5475,N_4126);
nand U7074 (N_7074,N_4724,N_4413);
or U7075 (N_7075,N_5422,N_4846);
nor U7076 (N_7076,N_4963,N_5081);
nand U7077 (N_7077,N_4610,N_5185);
or U7078 (N_7078,N_5445,N_5418);
and U7079 (N_7079,N_4716,N_5319);
or U7080 (N_7080,N_5884,N_4590);
nand U7081 (N_7081,N_5133,N_5756);
nor U7082 (N_7082,N_4338,N_4917);
nor U7083 (N_7083,N_4827,N_5357);
or U7084 (N_7084,N_4982,N_4008);
and U7085 (N_7085,N_4316,N_5152);
nor U7086 (N_7086,N_5703,N_4136);
nor U7087 (N_7087,N_5270,N_4018);
and U7088 (N_7088,N_4330,N_4728);
nor U7089 (N_7089,N_5531,N_4391);
nor U7090 (N_7090,N_4498,N_5571);
or U7091 (N_7091,N_5152,N_4134);
nand U7092 (N_7092,N_4415,N_5895);
nor U7093 (N_7093,N_5910,N_5924);
or U7094 (N_7094,N_5173,N_4531);
and U7095 (N_7095,N_5802,N_4427);
nor U7096 (N_7096,N_5706,N_4849);
or U7097 (N_7097,N_5125,N_5119);
nand U7098 (N_7098,N_5455,N_4573);
or U7099 (N_7099,N_4742,N_5533);
or U7100 (N_7100,N_4534,N_5681);
and U7101 (N_7101,N_4187,N_5394);
and U7102 (N_7102,N_5701,N_4877);
nand U7103 (N_7103,N_4994,N_5266);
nand U7104 (N_7104,N_4795,N_4179);
or U7105 (N_7105,N_5340,N_4694);
and U7106 (N_7106,N_5268,N_4166);
or U7107 (N_7107,N_5760,N_5929);
nor U7108 (N_7108,N_4621,N_5553);
nor U7109 (N_7109,N_4651,N_5560);
or U7110 (N_7110,N_4198,N_5338);
and U7111 (N_7111,N_4003,N_5590);
or U7112 (N_7112,N_4946,N_4761);
and U7113 (N_7113,N_4322,N_4755);
nand U7114 (N_7114,N_5163,N_4638);
or U7115 (N_7115,N_4856,N_4234);
and U7116 (N_7116,N_4943,N_5843);
nor U7117 (N_7117,N_5885,N_5643);
nor U7118 (N_7118,N_4808,N_5851);
and U7119 (N_7119,N_5853,N_4452);
nor U7120 (N_7120,N_4021,N_4165);
nand U7121 (N_7121,N_5667,N_5184);
nor U7122 (N_7122,N_5264,N_5449);
or U7123 (N_7123,N_5270,N_4674);
and U7124 (N_7124,N_4974,N_4110);
and U7125 (N_7125,N_5101,N_5988);
nand U7126 (N_7126,N_5638,N_4987);
and U7127 (N_7127,N_4118,N_4000);
and U7128 (N_7128,N_5125,N_4249);
and U7129 (N_7129,N_4733,N_5361);
and U7130 (N_7130,N_5367,N_4791);
nand U7131 (N_7131,N_4880,N_4943);
and U7132 (N_7132,N_4773,N_4143);
nand U7133 (N_7133,N_4510,N_5239);
and U7134 (N_7134,N_5739,N_4214);
or U7135 (N_7135,N_4167,N_5314);
nand U7136 (N_7136,N_5036,N_4885);
and U7137 (N_7137,N_4560,N_5299);
nand U7138 (N_7138,N_5650,N_4270);
and U7139 (N_7139,N_4535,N_4330);
nand U7140 (N_7140,N_4851,N_5601);
and U7141 (N_7141,N_5508,N_5969);
nand U7142 (N_7142,N_5264,N_5724);
nand U7143 (N_7143,N_4958,N_4795);
nor U7144 (N_7144,N_5377,N_5695);
and U7145 (N_7145,N_4120,N_4586);
nor U7146 (N_7146,N_5217,N_4696);
nand U7147 (N_7147,N_4966,N_5583);
and U7148 (N_7148,N_4536,N_5595);
nand U7149 (N_7149,N_4951,N_5282);
nand U7150 (N_7150,N_4712,N_4445);
or U7151 (N_7151,N_4600,N_5041);
nand U7152 (N_7152,N_4573,N_4448);
or U7153 (N_7153,N_5902,N_5617);
nor U7154 (N_7154,N_5502,N_5959);
nor U7155 (N_7155,N_5214,N_4529);
nor U7156 (N_7156,N_5719,N_4007);
nand U7157 (N_7157,N_5394,N_5239);
nand U7158 (N_7158,N_5718,N_5639);
nor U7159 (N_7159,N_5015,N_5877);
and U7160 (N_7160,N_5178,N_4446);
nor U7161 (N_7161,N_4849,N_5931);
and U7162 (N_7162,N_5898,N_4696);
or U7163 (N_7163,N_5486,N_5651);
and U7164 (N_7164,N_5925,N_4761);
and U7165 (N_7165,N_5429,N_4934);
and U7166 (N_7166,N_5077,N_4697);
and U7167 (N_7167,N_4321,N_4904);
or U7168 (N_7168,N_4644,N_4628);
or U7169 (N_7169,N_5168,N_5421);
or U7170 (N_7170,N_4594,N_5515);
or U7171 (N_7171,N_4318,N_4840);
nand U7172 (N_7172,N_5322,N_5157);
and U7173 (N_7173,N_4394,N_5795);
and U7174 (N_7174,N_4932,N_4207);
and U7175 (N_7175,N_4726,N_5379);
or U7176 (N_7176,N_5866,N_5009);
xnor U7177 (N_7177,N_4079,N_5208);
or U7178 (N_7178,N_4868,N_5901);
nand U7179 (N_7179,N_4693,N_5089);
and U7180 (N_7180,N_4168,N_4568);
nand U7181 (N_7181,N_5499,N_4957);
nand U7182 (N_7182,N_4640,N_5255);
and U7183 (N_7183,N_5271,N_4137);
or U7184 (N_7184,N_4385,N_4599);
and U7185 (N_7185,N_5194,N_5238);
or U7186 (N_7186,N_5335,N_5270);
and U7187 (N_7187,N_5453,N_5822);
or U7188 (N_7188,N_5112,N_5460);
nor U7189 (N_7189,N_4340,N_4989);
nand U7190 (N_7190,N_5889,N_5166);
and U7191 (N_7191,N_5335,N_5394);
and U7192 (N_7192,N_5552,N_4329);
or U7193 (N_7193,N_4464,N_4115);
xor U7194 (N_7194,N_4578,N_4102);
and U7195 (N_7195,N_4635,N_4012);
and U7196 (N_7196,N_4935,N_4160);
nor U7197 (N_7197,N_5648,N_4375);
or U7198 (N_7198,N_4940,N_5159);
nand U7199 (N_7199,N_5444,N_5192);
or U7200 (N_7200,N_4835,N_4053);
nor U7201 (N_7201,N_4355,N_4365);
and U7202 (N_7202,N_4491,N_4833);
or U7203 (N_7203,N_4394,N_4329);
nand U7204 (N_7204,N_5358,N_5379);
nand U7205 (N_7205,N_4000,N_5223);
or U7206 (N_7206,N_4775,N_5168);
nor U7207 (N_7207,N_4288,N_4007);
nand U7208 (N_7208,N_5648,N_4211);
nor U7209 (N_7209,N_5544,N_4406);
nor U7210 (N_7210,N_5991,N_4759);
or U7211 (N_7211,N_5655,N_5121);
nor U7212 (N_7212,N_5568,N_4096);
and U7213 (N_7213,N_5662,N_4341);
nand U7214 (N_7214,N_4667,N_5398);
nor U7215 (N_7215,N_5290,N_4324);
nor U7216 (N_7216,N_4121,N_4685);
nand U7217 (N_7217,N_5483,N_4880);
nor U7218 (N_7218,N_4845,N_4755);
or U7219 (N_7219,N_4985,N_5048);
nor U7220 (N_7220,N_5443,N_5382);
nor U7221 (N_7221,N_4380,N_5254);
or U7222 (N_7222,N_4109,N_5195);
and U7223 (N_7223,N_5811,N_4482);
and U7224 (N_7224,N_5712,N_4917);
nor U7225 (N_7225,N_4505,N_4385);
nand U7226 (N_7226,N_5166,N_4882);
nand U7227 (N_7227,N_4261,N_4860);
nor U7228 (N_7228,N_5480,N_5410);
nand U7229 (N_7229,N_4833,N_5979);
nor U7230 (N_7230,N_4183,N_5486);
and U7231 (N_7231,N_4149,N_5552);
nand U7232 (N_7232,N_5721,N_4671);
or U7233 (N_7233,N_4336,N_5704);
nand U7234 (N_7234,N_5821,N_5236);
or U7235 (N_7235,N_5162,N_4937);
or U7236 (N_7236,N_4136,N_4703);
or U7237 (N_7237,N_5672,N_4721);
nor U7238 (N_7238,N_4549,N_4781);
nand U7239 (N_7239,N_4416,N_4033);
or U7240 (N_7240,N_5560,N_5058);
nand U7241 (N_7241,N_5490,N_5080);
nor U7242 (N_7242,N_5719,N_5975);
nand U7243 (N_7243,N_4523,N_5534);
nand U7244 (N_7244,N_5380,N_4480);
nor U7245 (N_7245,N_4171,N_4244);
and U7246 (N_7246,N_5778,N_4464);
nand U7247 (N_7247,N_4619,N_5057);
nand U7248 (N_7248,N_4274,N_4377);
nand U7249 (N_7249,N_5861,N_4602);
nor U7250 (N_7250,N_5535,N_5058);
or U7251 (N_7251,N_4008,N_5407);
and U7252 (N_7252,N_5610,N_5290);
nand U7253 (N_7253,N_5634,N_4194);
or U7254 (N_7254,N_5137,N_5476);
nor U7255 (N_7255,N_5601,N_5214);
nor U7256 (N_7256,N_5959,N_5355);
or U7257 (N_7257,N_4359,N_4834);
or U7258 (N_7258,N_5531,N_4694);
nand U7259 (N_7259,N_5041,N_5449);
nand U7260 (N_7260,N_4932,N_5215);
nand U7261 (N_7261,N_5118,N_5262);
and U7262 (N_7262,N_4087,N_4363);
nand U7263 (N_7263,N_5531,N_5357);
nor U7264 (N_7264,N_5188,N_5765);
or U7265 (N_7265,N_5987,N_5795);
and U7266 (N_7266,N_4611,N_4951);
and U7267 (N_7267,N_5894,N_4740);
nand U7268 (N_7268,N_4156,N_5242);
nor U7269 (N_7269,N_5281,N_4535);
nand U7270 (N_7270,N_4659,N_5639);
or U7271 (N_7271,N_5317,N_5967);
nor U7272 (N_7272,N_5525,N_5067);
and U7273 (N_7273,N_5372,N_4682);
nand U7274 (N_7274,N_4125,N_5117);
nand U7275 (N_7275,N_5120,N_5292);
nand U7276 (N_7276,N_5817,N_5246);
nand U7277 (N_7277,N_5210,N_4699);
and U7278 (N_7278,N_5239,N_5778);
nor U7279 (N_7279,N_4433,N_5591);
nor U7280 (N_7280,N_4117,N_5644);
or U7281 (N_7281,N_4392,N_5801);
and U7282 (N_7282,N_5185,N_5526);
nor U7283 (N_7283,N_5388,N_4923);
nand U7284 (N_7284,N_5911,N_5201);
and U7285 (N_7285,N_4315,N_4950);
or U7286 (N_7286,N_5165,N_4913);
and U7287 (N_7287,N_5449,N_4607);
nand U7288 (N_7288,N_5368,N_5103);
nor U7289 (N_7289,N_5707,N_5919);
nand U7290 (N_7290,N_5560,N_5952);
or U7291 (N_7291,N_5671,N_5289);
nand U7292 (N_7292,N_5640,N_4188);
nand U7293 (N_7293,N_5872,N_5880);
or U7294 (N_7294,N_5342,N_4993);
nand U7295 (N_7295,N_4720,N_4899);
nand U7296 (N_7296,N_4191,N_5759);
and U7297 (N_7297,N_5959,N_4732);
nor U7298 (N_7298,N_4312,N_5546);
nor U7299 (N_7299,N_5523,N_5506);
or U7300 (N_7300,N_4674,N_4644);
and U7301 (N_7301,N_5394,N_5092);
nor U7302 (N_7302,N_5420,N_4668);
or U7303 (N_7303,N_4827,N_4353);
or U7304 (N_7304,N_5565,N_4307);
nand U7305 (N_7305,N_4609,N_4952);
and U7306 (N_7306,N_4954,N_5020);
or U7307 (N_7307,N_5592,N_5153);
or U7308 (N_7308,N_5393,N_5503);
nand U7309 (N_7309,N_4828,N_5177);
or U7310 (N_7310,N_4230,N_4923);
or U7311 (N_7311,N_4725,N_5867);
or U7312 (N_7312,N_5141,N_5351);
nand U7313 (N_7313,N_4576,N_4139);
nand U7314 (N_7314,N_4786,N_5504);
nand U7315 (N_7315,N_4519,N_5978);
or U7316 (N_7316,N_5846,N_5691);
or U7317 (N_7317,N_5237,N_4839);
nand U7318 (N_7318,N_4061,N_5456);
and U7319 (N_7319,N_5752,N_4052);
nor U7320 (N_7320,N_4313,N_5917);
nor U7321 (N_7321,N_4524,N_4559);
nor U7322 (N_7322,N_4075,N_5790);
or U7323 (N_7323,N_5346,N_5605);
or U7324 (N_7324,N_4869,N_5438);
and U7325 (N_7325,N_5372,N_4251);
and U7326 (N_7326,N_5083,N_4551);
nand U7327 (N_7327,N_5453,N_5978);
and U7328 (N_7328,N_5317,N_4535);
and U7329 (N_7329,N_5906,N_5093);
and U7330 (N_7330,N_4797,N_4613);
nor U7331 (N_7331,N_4209,N_4208);
or U7332 (N_7332,N_5116,N_5621);
or U7333 (N_7333,N_4596,N_5380);
or U7334 (N_7334,N_5319,N_5282);
nor U7335 (N_7335,N_4666,N_5227);
nor U7336 (N_7336,N_4156,N_4840);
nand U7337 (N_7337,N_4706,N_4397);
nand U7338 (N_7338,N_5321,N_5830);
and U7339 (N_7339,N_5119,N_4895);
nand U7340 (N_7340,N_4678,N_5631);
or U7341 (N_7341,N_4768,N_4861);
nand U7342 (N_7342,N_4690,N_4746);
and U7343 (N_7343,N_5238,N_4855);
nor U7344 (N_7344,N_5089,N_4155);
nand U7345 (N_7345,N_5836,N_4970);
or U7346 (N_7346,N_4180,N_5194);
and U7347 (N_7347,N_4720,N_5187);
nor U7348 (N_7348,N_4289,N_4704);
nand U7349 (N_7349,N_4906,N_4753);
nor U7350 (N_7350,N_4613,N_5104);
or U7351 (N_7351,N_5215,N_4000);
nand U7352 (N_7352,N_5885,N_4248);
nor U7353 (N_7353,N_5206,N_5419);
or U7354 (N_7354,N_4893,N_5363);
xnor U7355 (N_7355,N_4150,N_4533);
or U7356 (N_7356,N_5180,N_5573);
or U7357 (N_7357,N_5582,N_4149);
nor U7358 (N_7358,N_5608,N_4190);
and U7359 (N_7359,N_5766,N_4383);
and U7360 (N_7360,N_5413,N_5942);
nor U7361 (N_7361,N_4704,N_4251);
nand U7362 (N_7362,N_5076,N_5172);
xor U7363 (N_7363,N_4203,N_5094);
nor U7364 (N_7364,N_5127,N_5565);
and U7365 (N_7365,N_4700,N_4651);
or U7366 (N_7366,N_4002,N_4022);
nand U7367 (N_7367,N_4006,N_4818);
and U7368 (N_7368,N_4124,N_5601);
nor U7369 (N_7369,N_4918,N_4020);
and U7370 (N_7370,N_4920,N_4134);
or U7371 (N_7371,N_5633,N_5079);
nand U7372 (N_7372,N_5426,N_5636);
nor U7373 (N_7373,N_5733,N_4461);
or U7374 (N_7374,N_5832,N_5628);
nand U7375 (N_7375,N_5727,N_5653);
nand U7376 (N_7376,N_5475,N_5613);
nand U7377 (N_7377,N_4551,N_4556);
nand U7378 (N_7378,N_5062,N_5667);
nor U7379 (N_7379,N_5087,N_5559);
nor U7380 (N_7380,N_4080,N_4609);
nor U7381 (N_7381,N_5343,N_5542);
nor U7382 (N_7382,N_5420,N_5696);
and U7383 (N_7383,N_4271,N_4289);
nor U7384 (N_7384,N_4006,N_4473);
or U7385 (N_7385,N_4451,N_5386);
or U7386 (N_7386,N_4635,N_5816);
or U7387 (N_7387,N_5134,N_5313);
or U7388 (N_7388,N_5049,N_4833);
or U7389 (N_7389,N_5615,N_5289);
nand U7390 (N_7390,N_5663,N_4359);
and U7391 (N_7391,N_5271,N_5994);
and U7392 (N_7392,N_4182,N_5195);
nor U7393 (N_7393,N_5668,N_4559);
or U7394 (N_7394,N_5158,N_5997);
nor U7395 (N_7395,N_5657,N_4571);
nor U7396 (N_7396,N_5618,N_5691);
and U7397 (N_7397,N_4414,N_4811);
nor U7398 (N_7398,N_5934,N_5227);
nand U7399 (N_7399,N_4484,N_4470);
nand U7400 (N_7400,N_4145,N_5257);
and U7401 (N_7401,N_4662,N_4114);
or U7402 (N_7402,N_4862,N_4856);
and U7403 (N_7403,N_4741,N_5951);
or U7404 (N_7404,N_5299,N_5532);
or U7405 (N_7405,N_4093,N_5472);
nand U7406 (N_7406,N_5242,N_5934);
nand U7407 (N_7407,N_5383,N_5442);
nor U7408 (N_7408,N_4530,N_4167);
nor U7409 (N_7409,N_4162,N_5024);
nor U7410 (N_7410,N_4670,N_4931);
nand U7411 (N_7411,N_4928,N_5613);
nor U7412 (N_7412,N_4003,N_5192);
or U7413 (N_7413,N_5024,N_4529);
nor U7414 (N_7414,N_5133,N_4835);
nor U7415 (N_7415,N_4585,N_5579);
and U7416 (N_7416,N_4877,N_5795);
nand U7417 (N_7417,N_4352,N_5764);
nand U7418 (N_7418,N_5984,N_4124);
nor U7419 (N_7419,N_4341,N_4977);
and U7420 (N_7420,N_4440,N_4201);
and U7421 (N_7421,N_5989,N_5644);
nor U7422 (N_7422,N_5384,N_4910);
or U7423 (N_7423,N_4385,N_4412);
nor U7424 (N_7424,N_4335,N_4650);
nor U7425 (N_7425,N_5336,N_4096);
nor U7426 (N_7426,N_5677,N_5315);
and U7427 (N_7427,N_4907,N_5319);
and U7428 (N_7428,N_4669,N_5099);
nand U7429 (N_7429,N_4610,N_4002);
nor U7430 (N_7430,N_5487,N_4143);
and U7431 (N_7431,N_4158,N_4569);
and U7432 (N_7432,N_4113,N_5776);
nor U7433 (N_7433,N_5678,N_5487);
or U7434 (N_7434,N_5926,N_4945);
and U7435 (N_7435,N_4505,N_4575);
nor U7436 (N_7436,N_5894,N_5703);
nand U7437 (N_7437,N_5695,N_4887);
and U7438 (N_7438,N_5153,N_4361);
nor U7439 (N_7439,N_5585,N_4727);
and U7440 (N_7440,N_4217,N_4262);
nand U7441 (N_7441,N_4474,N_4796);
nor U7442 (N_7442,N_4079,N_4743);
nor U7443 (N_7443,N_4273,N_5421);
and U7444 (N_7444,N_4862,N_4719);
or U7445 (N_7445,N_4257,N_5627);
or U7446 (N_7446,N_4840,N_5348);
or U7447 (N_7447,N_5867,N_5171);
and U7448 (N_7448,N_4124,N_4168);
and U7449 (N_7449,N_5525,N_5305);
and U7450 (N_7450,N_4067,N_5894);
and U7451 (N_7451,N_4561,N_4366);
nor U7452 (N_7452,N_4372,N_4422);
nand U7453 (N_7453,N_4571,N_5511);
nor U7454 (N_7454,N_4873,N_4341);
nand U7455 (N_7455,N_5517,N_5824);
nor U7456 (N_7456,N_4900,N_5808);
nand U7457 (N_7457,N_4462,N_4534);
nand U7458 (N_7458,N_5347,N_5351);
nor U7459 (N_7459,N_5581,N_4828);
nor U7460 (N_7460,N_5268,N_5948);
or U7461 (N_7461,N_5916,N_5567);
nand U7462 (N_7462,N_4728,N_5500);
nor U7463 (N_7463,N_5158,N_4443);
or U7464 (N_7464,N_5030,N_5091);
nand U7465 (N_7465,N_5301,N_5666);
nand U7466 (N_7466,N_5906,N_4551);
nand U7467 (N_7467,N_4968,N_5006);
nor U7468 (N_7468,N_5422,N_4361);
and U7469 (N_7469,N_4760,N_5214);
or U7470 (N_7470,N_4691,N_5515);
and U7471 (N_7471,N_5683,N_5251);
nor U7472 (N_7472,N_4722,N_4438);
nor U7473 (N_7473,N_5644,N_4336);
nor U7474 (N_7474,N_5557,N_5526);
xor U7475 (N_7475,N_4079,N_5038);
nand U7476 (N_7476,N_4293,N_4234);
xor U7477 (N_7477,N_5449,N_4543);
and U7478 (N_7478,N_5520,N_4699);
and U7479 (N_7479,N_4848,N_4596);
or U7480 (N_7480,N_5386,N_4124);
and U7481 (N_7481,N_4059,N_5029);
nand U7482 (N_7482,N_4582,N_5616);
nor U7483 (N_7483,N_5305,N_4551);
nand U7484 (N_7484,N_5302,N_4742);
or U7485 (N_7485,N_4069,N_4242);
and U7486 (N_7486,N_5814,N_4953);
nor U7487 (N_7487,N_5800,N_5430);
nand U7488 (N_7488,N_4633,N_5009);
and U7489 (N_7489,N_4441,N_5481);
nand U7490 (N_7490,N_4456,N_4708);
or U7491 (N_7491,N_5847,N_4339);
or U7492 (N_7492,N_4246,N_4989);
or U7493 (N_7493,N_4813,N_4558);
nor U7494 (N_7494,N_4534,N_5391);
nand U7495 (N_7495,N_5936,N_4961);
or U7496 (N_7496,N_4696,N_4235);
nor U7497 (N_7497,N_4496,N_5145);
nor U7498 (N_7498,N_4657,N_4035);
or U7499 (N_7499,N_4705,N_4928);
and U7500 (N_7500,N_5105,N_4690);
or U7501 (N_7501,N_4378,N_5497);
or U7502 (N_7502,N_5279,N_4061);
or U7503 (N_7503,N_4532,N_4468);
or U7504 (N_7504,N_4165,N_4871);
nand U7505 (N_7505,N_5431,N_4510);
and U7506 (N_7506,N_5016,N_5764);
nor U7507 (N_7507,N_4577,N_4837);
or U7508 (N_7508,N_4846,N_5348);
nand U7509 (N_7509,N_5443,N_4684);
or U7510 (N_7510,N_4783,N_5983);
and U7511 (N_7511,N_4599,N_5860);
and U7512 (N_7512,N_5013,N_5934);
nor U7513 (N_7513,N_4588,N_5340);
and U7514 (N_7514,N_4616,N_4022);
nand U7515 (N_7515,N_5106,N_5839);
nor U7516 (N_7516,N_5363,N_4920);
and U7517 (N_7517,N_4440,N_4027);
xor U7518 (N_7518,N_4625,N_5917);
or U7519 (N_7519,N_5337,N_5641);
nand U7520 (N_7520,N_4787,N_4637);
or U7521 (N_7521,N_5956,N_5596);
nor U7522 (N_7522,N_5746,N_5906);
nor U7523 (N_7523,N_4905,N_4964);
or U7524 (N_7524,N_4460,N_4437);
or U7525 (N_7525,N_5458,N_5770);
and U7526 (N_7526,N_4661,N_5353);
nor U7527 (N_7527,N_4547,N_5578);
and U7528 (N_7528,N_5094,N_4173);
nor U7529 (N_7529,N_4197,N_4686);
nand U7530 (N_7530,N_4571,N_5128);
and U7531 (N_7531,N_4130,N_5699);
and U7532 (N_7532,N_5610,N_4922);
or U7533 (N_7533,N_5923,N_5262);
and U7534 (N_7534,N_5811,N_4196);
and U7535 (N_7535,N_4128,N_4416);
or U7536 (N_7536,N_4134,N_5120);
nor U7537 (N_7537,N_4849,N_5170);
or U7538 (N_7538,N_4823,N_5304);
and U7539 (N_7539,N_5156,N_4029);
and U7540 (N_7540,N_5977,N_5913);
nand U7541 (N_7541,N_5257,N_4594);
or U7542 (N_7542,N_5389,N_5281);
nor U7543 (N_7543,N_5414,N_5609);
nor U7544 (N_7544,N_5653,N_5227);
and U7545 (N_7545,N_4871,N_5651);
and U7546 (N_7546,N_4048,N_4626);
or U7547 (N_7547,N_5250,N_4020);
or U7548 (N_7548,N_4473,N_4884);
nor U7549 (N_7549,N_5302,N_5621);
nor U7550 (N_7550,N_4860,N_4101);
nor U7551 (N_7551,N_5109,N_4659);
and U7552 (N_7552,N_5802,N_4421);
or U7553 (N_7553,N_5641,N_4440);
or U7554 (N_7554,N_5146,N_4693);
nand U7555 (N_7555,N_5798,N_5678);
and U7556 (N_7556,N_4132,N_5595);
or U7557 (N_7557,N_5522,N_4390);
and U7558 (N_7558,N_4888,N_4846);
nand U7559 (N_7559,N_5367,N_4065);
and U7560 (N_7560,N_5705,N_5319);
or U7561 (N_7561,N_4935,N_4166);
nor U7562 (N_7562,N_4923,N_5040);
or U7563 (N_7563,N_4993,N_5085);
nand U7564 (N_7564,N_4295,N_5944);
and U7565 (N_7565,N_5620,N_4703);
and U7566 (N_7566,N_4568,N_5436);
and U7567 (N_7567,N_4367,N_5635);
nand U7568 (N_7568,N_5128,N_5181);
nor U7569 (N_7569,N_4464,N_4282);
nand U7570 (N_7570,N_4771,N_4077);
nor U7571 (N_7571,N_5483,N_5313);
nand U7572 (N_7572,N_5709,N_4003);
nand U7573 (N_7573,N_4446,N_4251);
nand U7574 (N_7574,N_5270,N_4930);
nor U7575 (N_7575,N_5181,N_5458);
and U7576 (N_7576,N_5391,N_5508);
and U7577 (N_7577,N_4786,N_4550);
nand U7578 (N_7578,N_5408,N_4104);
nor U7579 (N_7579,N_4257,N_5331);
nand U7580 (N_7580,N_4305,N_4088);
nor U7581 (N_7581,N_5808,N_4807);
or U7582 (N_7582,N_5537,N_5365);
nor U7583 (N_7583,N_5829,N_4148);
and U7584 (N_7584,N_4064,N_5300);
nor U7585 (N_7585,N_5248,N_5374);
nor U7586 (N_7586,N_4276,N_5310);
nand U7587 (N_7587,N_5904,N_4270);
and U7588 (N_7588,N_5871,N_4458);
nand U7589 (N_7589,N_5012,N_4190);
and U7590 (N_7590,N_4678,N_5015);
nor U7591 (N_7591,N_5768,N_5167);
nand U7592 (N_7592,N_5538,N_5109);
nand U7593 (N_7593,N_4632,N_4290);
or U7594 (N_7594,N_4561,N_5814);
and U7595 (N_7595,N_5326,N_5676);
and U7596 (N_7596,N_5582,N_5913);
nand U7597 (N_7597,N_5648,N_5548);
nand U7598 (N_7598,N_4125,N_4676);
nand U7599 (N_7599,N_5690,N_4185);
nand U7600 (N_7600,N_5151,N_4360);
nand U7601 (N_7601,N_4538,N_5239);
and U7602 (N_7602,N_5306,N_5512);
or U7603 (N_7603,N_5688,N_4367);
nand U7604 (N_7604,N_5493,N_4929);
or U7605 (N_7605,N_5813,N_4090);
nor U7606 (N_7606,N_4221,N_5693);
and U7607 (N_7607,N_4859,N_4586);
nand U7608 (N_7608,N_4826,N_5926);
or U7609 (N_7609,N_5984,N_4824);
nand U7610 (N_7610,N_4811,N_4524);
nand U7611 (N_7611,N_5081,N_5295);
or U7612 (N_7612,N_4526,N_5090);
and U7613 (N_7613,N_5196,N_4593);
nor U7614 (N_7614,N_5760,N_5071);
nor U7615 (N_7615,N_4203,N_5961);
nor U7616 (N_7616,N_4239,N_5092);
nand U7617 (N_7617,N_4393,N_5660);
nand U7618 (N_7618,N_4001,N_5817);
xor U7619 (N_7619,N_5772,N_5695);
nor U7620 (N_7620,N_4637,N_5341);
nand U7621 (N_7621,N_5710,N_4880);
and U7622 (N_7622,N_5596,N_5592);
and U7623 (N_7623,N_5352,N_4405);
or U7624 (N_7624,N_4165,N_4898);
and U7625 (N_7625,N_4601,N_4370);
or U7626 (N_7626,N_4592,N_4144);
and U7627 (N_7627,N_4785,N_4822);
or U7628 (N_7628,N_5147,N_4348);
or U7629 (N_7629,N_4393,N_4516);
and U7630 (N_7630,N_4204,N_4160);
and U7631 (N_7631,N_5768,N_5503);
and U7632 (N_7632,N_4308,N_5139);
nand U7633 (N_7633,N_4152,N_5846);
nand U7634 (N_7634,N_4224,N_4027);
nand U7635 (N_7635,N_4005,N_4582);
and U7636 (N_7636,N_4136,N_5770);
and U7637 (N_7637,N_4492,N_4866);
and U7638 (N_7638,N_4095,N_5647);
nor U7639 (N_7639,N_5803,N_4737);
nor U7640 (N_7640,N_4537,N_5896);
and U7641 (N_7641,N_4259,N_5512);
nand U7642 (N_7642,N_4771,N_5891);
nand U7643 (N_7643,N_5432,N_4249);
or U7644 (N_7644,N_5485,N_4866);
nor U7645 (N_7645,N_5076,N_4845);
nand U7646 (N_7646,N_4676,N_4545);
or U7647 (N_7647,N_5236,N_4987);
nand U7648 (N_7648,N_5138,N_4946);
nor U7649 (N_7649,N_4086,N_5590);
nor U7650 (N_7650,N_5118,N_4064);
and U7651 (N_7651,N_4546,N_5818);
nor U7652 (N_7652,N_4935,N_5323);
nor U7653 (N_7653,N_5975,N_5744);
nor U7654 (N_7654,N_5009,N_4848);
nand U7655 (N_7655,N_5804,N_4955);
nand U7656 (N_7656,N_4617,N_4072);
nor U7657 (N_7657,N_4401,N_4118);
nor U7658 (N_7658,N_4506,N_5706);
nor U7659 (N_7659,N_4444,N_4663);
nor U7660 (N_7660,N_4265,N_5579);
nor U7661 (N_7661,N_4398,N_5173);
and U7662 (N_7662,N_4021,N_5605);
nand U7663 (N_7663,N_5963,N_4411);
nor U7664 (N_7664,N_5033,N_4099);
or U7665 (N_7665,N_4606,N_4446);
nor U7666 (N_7666,N_5330,N_5937);
nand U7667 (N_7667,N_5927,N_5862);
nand U7668 (N_7668,N_5945,N_4067);
or U7669 (N_7669,N_5701,N_5712);
and U7670 (N_7670,N_4721,N_5841);
nand U7671 (N_7671,N_5905,N_5110);
and U7672 (N_7672,N_4857,N_4041);
nor U7673 (N_7673,N_5716,N_5592);
nand U7674 (N_7674,N_5069,N_5587);
nor U7675 (N_7675,N_4464,N_4971);
nand U7676 (N_7676,N_4245,N_4582);
nand U7677 (N_7677,N_5914,N_4514);
nand U7678 (N_7678,N_4818,N_5809);
and U7679 (N_7679,N_4485,N_4613);
or U7680 (N_7680,N_4751,N_4916);
nand U7681 (N_7681,N_4905,N_5373);
nor U7682 (N_7682,N_4240,N_4776);
and U7683 (N_7683,N_4013,N_5371);
or U7684 (N_7684,N_4146,N_4208);
nand U7685 (N_7685,N_4332,N_4691);
nor U7686 (N_7686,N_4764,N_5248);
nor U7687 (N_7687,N_5488,N_5005);
nand U7688 (N_7688,N_5081,N_4051);
xor U7689 (N_7689,N_4860,N_5236);
nand U7690 (N_7690,N_5983,N_5589);
and U7691 (N_7691,N_5983,N_4219);
nand U7692 (N_7692,N_5753,N_5042);
or U7693 (N_7693,N_4247,N_5533);
and U7694 (N_7694,N_4206,N_5417);
xor U7695 (N_7695,N_5299,N_4178);
xor U7696 (N_7696,N_5007,N_5583);
nand U7697 (N_7697,N_5912,N_4804);
or U7698 (N_7698,N_4069,N_4061);
or U7699 (N_7699,N_4209,N_5368);
and U7700 (N_7700,N_4677,N_5987);
or U7701 (N_7701,N_5324,N_5291);
nor U7702 (N_7702,N_4025,N_5737);
or U7703 (N_7703,N_4264,N_4982);
nor U7704 (N_7704,N_5809,N_4218);
or U7705 (N_7705,N_5024,N_5774);
nand U7706 (N_7706,N_4081,N_5677);
or U7707 (N_7707,N_5068,N_4380);
nand U7708 (N_7708,N_4410,N_5784);
and U7709 (N_7709,N_4524,N_5241);
nor U7710 (N_7710,N_4035,N_5673);
or U7711 (N_7711,N_5439,N_5330);
nor U7712 (N_7712,N_5780,N_4955);
nor U7713 (N_7713,N_4513,N_5765);
or U7714 (N_7714,N_5425,N_4352);
or U7715 (N_7715,N_4206,N_4093);
or U7716 (N_7716,N_5005,N_4457);
nand U7717 (N_7717,N_4711,N_4553);
or U7718 (N_7718,N_5042,N_4722);
nor U7719 (N_7719,N_5921,N_4717);
nor U7720 (N_7720,N_5352,N_5490);
xor U7721 (N_7721,N_5661,N_4680);
nor U7722 (N_7722,N_5272,N_4071);
nor U7723 (N_7723,N_5541,N_4627);
nand U7724 (N_7724,N_5145,N_4666);
nand U7725 (N_7725,N_4503,N_5588);
and U7726 (N_7726,N_4870,N_4887);
nor U7727 (N_7727,N_5235,N_4187);
and U7728 (N_7728,N_5266,N_4802);
nand U7729 (N_7729,N_5941,N_4289);
or U7730 (N_7730,N_5722,N_5259);
nand U7731 (N_7731,N_4588,N_5470);
and U7732 (N_7732,N_4512,N_4630);
or U7733 (N_7733,N_4358,N_4138);
and U7734 (N_7734,N_4136,N_4258);
or U7735 (N_7735,N_4109,N_5181);
nand U7736 (N_7736,N_4265,N_5781);
nor U7737 (N_7737,N_4765,N_4430);
and U7738 (N_7738,N_5577,N_4923);
nand U7739 (N_7739,N_5340,N_4222);
or U7740 (N_7740,N_4297,N_4179);
and U7741 (N_7741,N_5353,N_4075);
nand U7742 (N_7742,N_5276,N_4932);
nor U7743 (N_7743,N_4363,N_4712);
nor U7744 (N_7744,N_4799,N_4264);
and U7745 (N_7745,N_5823,N_5692);
or U7746 (N_7746,N_5732,N_4844);
or U7747 (N_7747,N_4266,N_4940);
nor U7748 (N_7748,N_5334,N_5593);
or U7749 (N_7749,N_4482,N_5323);
nor U7750 (N_7750,N_5213,N_4665);
or U7751 (N_7751,N_5598,N_4795);
or U7752 (N_7752,N_5885,N_4163);
or U7753 (N_7753,N_4276,N_4212);
nor U7754 (N_7754,N_5344,N_4310);
and U7755 (N_7755,N_4301,N_5964);
and U7756 (N_7756,N_4772,N_4295);
or U7757 (N_7757,N_4535,N_4830);
and U7758 (N_7758,N_4046,N_5857);
and U7759 (N_7759,N_5282,N_5277);
or U7760 (N_7760,N_4978,N_4281);
nand U7761 (N_7761,N_5665,N_5844);
nand U7762 (N_7762,N_5928,N_4490);
or U7763 (N_7763,N_5676,N_4608);
or U7764 (N_7764,N_4517,N_4003);
or U7765 (N_7765,N_4419,N_4588);
and U7766 (N_7766,N_4982,N_4587);
nor U7767 (N_7767,N_4947,N_5034);
nand U7768 (N_7768,N_4222,N_5916);
or U7769 (N_7769,N_4108,N_5710);
nand U7770 (N_7770,N_4765,N_5823);
nand U7771 (N_7771,N_4487,N_5317);
nor U7772 (N_7772,N_5309,N_5089);
nand U7773 (N_7773,N_5490,N_4122);
nand U7774 (N_7774,N_5705,N_5575);
nor U7775 (N_7775,N_4915,N_5932);
nor U7776 (N_7776,N_5332,N_4911);
nand U7777 (N_7777,N_4416,N_5237);
or U7778 (N_7778,N_5297,N_5644);
and U7779 (N_7779,N_5987,N_4441);
or U7780 (N_7780,N_4240,N_5194);
or U7781 (N_7781,N_5598,N_4417);
nor U7782 (N_7782,N_4267,N_5977);
xnor U7783 (N_7783,N_5453,N_5882);
nand U7784 (N_7784,N_5229,N_5693);
or U7785 (N_7785,N_5233,N_4064);
and U7786 (N_7786,N_4289,N_5408);
or U7787 (N_7787,N_5160,N_5863);
nor U7788 (N_7788,N_5359,N_4396);
or U7789 (N_7789,N_5049,N_5023);
nand U7790 (N_7790,N_4516,N_5610);
and U7791 (N_7791,N_5039,N_5783);
and U7792 (N_7792,N_5962,N_4585);
nor U7793 (N_7793,N_4198,N_4766);
and U7794 (N_7794,N_4126,N_4989);
and U7795 (N_7795,N_4566,N_5246);
or U7796 (N_7796,N_5884,N_4614);
and U7797 (N_7797,N_5516,N_4228);
or U7798 (N_7798,N_5918,N_5152);
or U7799 (N_7799,N_4843,N_5292);
or U7800 (N_7800,N_4694,N_5731);
nand U7801 (N_7801,N_4185,N_4905);
nor U7802 (N_7802,N_5423,N_4717);
and U7803 (N_7803,N_4196,N_5423);
or U7804 (N_7804,N_5001,N_5171);
or U7805 (N_7805,N_4020,N_5802);
nor U7806 (N_7806,N_5593,N_5381);
nand U7807 (N_7807,N_5294,N_5888);
nand U7808 (N_7808,N_5168,N_4691);
xnor U7809 (N_7809,N_5352,N_5276);
and U7810 (N_7810,N_4893,N_4658);
and U7811 (N_7811,N_4939,N_4343);
xnor U7812 (N_7812,N_4641,N_5952);
or U7813 (N_7813,N_5866,N_5833);
nor U7814 (N_7814,N_5929,N_4710);
or U7815 (N_7815,N_4220,N_4952);
nor U7816 (N_7816,N_4549,N_5647);
and U7817 (N_7817,N_4891,N_4199);
or U7818 (N_7818,N_5512,N_4058);
or U7819 (N_7819,N_5787,N_4024);
nand U7820 (N_7820,N_5312,N_5439);
or U7821 (N_7821,N_5561,N_5500);
or U7822 (N_7822,N_4731,N_4285);
or U7823 (N_7823,N_4364,N_5983);
and U7824 (N_7824,N_4339,N_4951);
or U7825 (N_7825,N_5958,N_4450);
or U7826 (N_7826,N_4443,N_5333);
nor U7827 (N_7827,N_4563,N_5720);
or U7828 (N_7828,N_5761,N_4533);
nor U7829 (N_7829,N_5027,N_5537);
nand U7830 (N_7830,N_5671,N_4063);
or U7831 (N_7831,N_4155,N_5363);
or U7832 (N_7832,N_4133,N_5413);
nor U7833 (N_7833,N_4666,N_4597);
and U7834 (N_7834,N_4868,N_4570);
and U7835 (N_7835,N_4977,N_4751);
nor U7836 (N_7836,N_5923,N_4901);
and U7837 (N_7837,N_4679,N_5805);
or U7838 (N_7838,N_5408,N_4504);
xor U7839 (N_7839,N_4572,N_5964);
and U7840 (N_7840,N_5359,N_4854);
nor U7841 (N_7841,N_5443,N_4477);
or U7842 (N_7842,N_5591,N_4599);
nor U7843 (N_7843,N_4456,N_4976);
and U7844 (N_7844,N_5707,N_4197);
nand U7845 (N_7845,N_4969,N_4086);
nor U7846 (N_7846,N_4673,N_5447);
or U7847 (N_7847,N_4578,N_4258);
and U7848 (N_7848,N_5382,N_5262);
nand U7849 (N_7849,N_5971,N_4664);
and U7850 (N_7850,N_4554,N_4826);
nor U7851 (N_7851,N_5144,N_4165);
or U7852 (N_7852,N_5693,N_4733);
or U7853 (N_7853,N_4997,N_4717);
or U7854 (N_7854,N_4195,N_4740);
xnor U7855 (N_7855,N_4499,N_4799);
nand U7856 (N_7856,N_5499,N_5870);
and U7857 (N_7857,N_4700,N_5688);
nor U7858 (N_7858,N_4250,N_5638);
nand U7859 (N_7859,N_4966,N_4429);
and U7860 (N_7860,N_4423,N_4205);
nor U7861 (N_7861,N_4542,N_4750);
or U7862 (N_7862,N_5629,N_4820);
nor U7863 (N_7863,N_5210,N_5137);
or U7864 (N_7864,N_5205,N_5104);
nand U7865 (N_7865,N_4405,N_4868);
and U7866 (N_7866,N_4888,N_5368);
nand U7867 (N_7867,N_4467,N_5417);
nor U7868 (N_7868,N_5202,N_5927);
and U7869 (N_7869,N_5907,N_5254);
nor U7870 (N_7870,N_4226,N_5027);
nor U7871 (N_7871,N_4988,N_5447);
nor U7872 (N_7872,N_5231,N_4581);
and U7873 (N_7873,N_4109,N_4843);
nand U7874 (N_7874,N_4791,N_5194);
or U7875 (N_7875,N_5018,N_4832);
and U7876 (N_7876,N_4553,N_4582);
nand U7877 (N_7877,N_5619,N_5727);
or U7878 (N_7878,N_5086,N_4608);
nand U7879 (N_7879,N_5352,N_5816);
nand U7880 (N_7880,N_4619,N_4785);
nor U7881 (N_7881,N_5196,N_4842);
nor U7882 (N_7882,N_4480,N_4315);
nor U7883 (N_7883,N_5736,N_5051);
and U7884 (N_7884,N_4082,N_4333);
and U7885 (N_7885,N_5372,N_4630);
and U7886 (N_7886,N_5733,N_5490);
nand U7887 (N_7887,N_4468,N_5566);
nor U7888 (N_7888,N_5688,N_4659);
nand U7889 (N_7889,N_5933,N_4003);
nand U7890 (N_7890,N_5240,N_4737);
and U7891 (N_7891,N_5649,N_4253);
and U7892 (N_7892,N_4205,N_4341);
or U7893 (N_7893,N_4423,N_5943);
nand U7894 (N_7894,N_5269,N_5270);
or U7895 (N_7895,N_5010,N_4507);
and U7896 (N_7896,N_4529,N_5946);
nor U7897 (N_7897,N_5928,N_4701);
nor U7898 (N_7898,N_5426,N_4722);
or U7899 (N_7899,N_5617,N_5832);
and U7900 (N_7900,N_4219,N_5093);
nand U7901 (N_7901,N_4543,N_4313);
or U7902 (N_7902,N_4563,N_5067);
or U7903 (N_7903,N_5651,N_5799);
and U7904 (N_7904,N_5387,N_5097);
or U7905 (N_7905,N_5850,N_5248);
nand U7906 (N_7906,N_4969,N_4475);
and U7907 (N_7907,N_4529,N_5961);
nor U7908 (N_7908,N_5428,N_4554);
nor U7909 (N_7909,N_4266,N_4456);
or U7910 (N_7910,N_5573,N_5841);
nand U7911 (N_7911,N_5898,N_5655);
and U7912 (N_7912,N_4169,N_4370);
nor U7913 (N_7913,N_5281,N_5424);
nand U7914 (N_7914,N_4989,N_5252);
and U7915 (N_7915,N_5144,N_5140);
and U7916 (N_7916,N_4881,N_4166);
or U7917 (N_7917,N_4028,N_5578);
nor U7918 (N_7918,N_5444,N_4370);
nor U7919 (N_7919,N_4237,N_5112);
or U7920 (N_7920,N_5206,N_4386);
or U7921 (N_7921,N_4112,N_5469);
and U7922 (N_7922,N_4460,N_4794);
and U7923 (N_7923,N_5237,N_4384);
and U7924 (N_7924,N_5203,N_4182);
xnor U7925 (N_7925,N_4084,N_5217);
xor U7926 (N_7926,N_4178,N_5425);
or U7927 (N_7927,N_5785,N_5646);
and U7928 (N_7928,N_4243,N_5591);
nor U7929 (N_7929,N_5820,N_5976);
nand U7930 (N_7930,N_5954,N_5285);
nand U7931 (N_7931,N_5307,N_5072);
nand U7932 (N_7932,N_5340,N_5543);
or U7933 (N_7933,N_4483,N_4208);
or U7934 (N_7934,N_5205,N_5444);
and U7935 (N_7935,N_5951,N_5808);
and U7936 (N_7936,N_5313,N_4371);
nand U7937 (N_7937,N_4220,N_5294);
nand U7938 (N_7938,N_5951,N_4893);
nor U7939 (N_7939,N_5902,N_5094);
or U7940 (N_7940,N_4995,N_5924);
nand U7941 (N_7941,N_4257,N_4285);
nor U7942 (N_7942,N_4378,N_5808);
nand U7943 (N_7943,N_4685,N_5846);
nor U7944 (N_7944,N_4818,N_4444);
nand U7945 (N_7945,N_5530,N_4533);
and U7946 (N_7946,N_5115,N_4154);
or U7947 (N_7947,N_5597,N_4592);
or U7948 (N_7948,N_4115,N_5435);
nor U7949 (N_7949,N_4894,N_4451);
nor U7950 (N_7950,N_4435,N_5774);
nand U7951 (N_7951,N_4347,N_4613);
xnor U7952 (N_7952,N_5949,N_5248);
nand U7953 (N_7953,N_4347,N_4670);
and U7954 (N_7954,N_5150,N_4529);
nor U7955 (N_7955,N_4488,N_5876);
nand U7956 (N_7956,N_5298,N_4435);
and U7957 (N_7957,N_5844,N_5792);
and U7958 (N_7958,N_4898,N_4356);
and U7959 (N_7959,N_4971,N_4804);
nor U7960 (N_7960,N_5314,N_4371);
nand U7961 (N_7961,N_5590,N_5996);
and U7962 (N_7962,N_5076,N_5878);
and U7963 (N_7963,N_4988,N_5307);
and U7964 (N_7964,N_5256,N_4384);
nor U7965 (N_7965,N_4896,N_5844);
or U7966 (N_7966,N_5628,N_5436);
or U7967 (N_7967,N_4550,N_5780);
or U7968 (N_7968,N_5204,N_5972);
nor U7969 (N_7969,N_4845,N_5042);
or U7970 (N_7970,N_4894,N_5710);
or U7971 (N_7971,N_5094,N_4196);
and U7972 (N_7972,N_4788,N_5893);
nand U7973 (N_7973,N_5922,N_5392);
nor U7974 (N_7974,N_4590,N_5173);
and U7975 (N_7975,N_4553,N_4466);
nand U7976 (N_7976,N_4695,N_5681);
and U7977 (N_7977,N_5081,N_4016);
nand U7978 (N_7978,N_4644,N_4323);
and U7979 (N_7979,N_4458,N_5330);
nand U7980 (N_7980,N_5768,N_5562);
nand U7981 (N_7981,N_5455,N_4984);
or U7982 (N_7982,N_5572,N_5220);
or U7983 (N_7983,N_5090,N_5427);
nor U7984 (N_7984,N_5461,N_5543);
nor U7985 (N_7985,N_5755,N_4863);
and U7986 (N_7986,N_5845,N_4446);
or U7987 (N_7987,N_4548,N_4496);
and U7988 (N_7988,N_5756,N_4108);
and U7989 (N_7989,N_5476,N_4947);
nor U7990 (N_7990,N_5647,N_4113);
nor U7991 (N_7991,N_4298,N_4327);
nand U7992 (N_7992,N_4073,N_5866);
nand U7993 (N_7993,N_5233,N_4255);
nor U7994 (N_7994,N_4959,N_4414);
nand U7995 (N_7995,N_4020,N_4283);
and U7996 (N_7996,N_4999,N_4979);
or U7997 (N_7997,N_4238,N_5646);
nor U7998 (N_7998,N_4441,N_4865);
and U7999 (N_7999,N_4668,N_5958);
or U8000 (N_8000,N_7831,N_6676);
nor U8001 (N_8001,N_7193,N_6689);
or U8002 (N_8002,N_7672,N_7025);
or U8003 (N_8003,N_7994,N_7230);
or U8004 (N_8004,N_6204,N_7507);
nor U8005 (N_8005,N_6443,N_6209);
or U8006 (N_8006,N_7717,N_7481);
nor U8007 (N_8007,N_7549,N_6810);
and U8008 (N_8008,N_7220,N_6243);
or U8009 (N_8009,N_6920,N_7685);
and U8010 (N_8010,N_6526,N_7370);
nor U8011 (N_8011,N_6165,N_6085);
and U8012 (N_8012,N_6587,N_6698);
nor U8013 (N_8013,N_7542,N_6850);
or U8014 (N_8014,N_7879,N_7848);
nand U8015 (N_8015,N_7505,N_7005);
nand U8016 (N_8016,N_6717,N_6666);
or U8017 (N_8017,N_6685,N_6762);
and U8018 (N_8018,N_7449,N_7476);
nor U8019 (N_8019,N_7828,N_6068);
nand U8020 (N_8020,N_7209,N_6706);
nand U8021 (N_8021,N_7718,N_6994);
xor U8022 (N_8022,N_7534,N_7153);
nand U8023 (N_8023,N_6259,N_6329);
and U8024 (N_8024,N_6694,N_6733);
nor U8025 (N_8025,N_7937,N_7055);
nor U8026 (N_8026,N_7281,N_6188);
nand U8027 (N_8027,N_7561,N_7635);
and U8028 (N_8028,N_6276,N_6976);
nor U8029 (N_8029,N_7019,N_6396);
nand U8030 (N_8030,N_6664,N_6321);
and U8031 (N_8031,N_6064,N_6556);
and U8032 (N_8032,N_7749,N_7160);
nor U8033 (N_8033,N_6568,N_7519);
and U8034 (N_8034,N_6703,N_7002);
nor U8035 (N_8035,N_6506,N_6932);
nor U8036 (N_8036,N_7930,N_6109);
nor U8037 (N_8037,N_6977,N_6967);
and U8038 (N_8038,N_7909,N_7889);
nand U8039 (N_8039,N_7859,N_7675);
nor U8040 (N_8040,N_6848,N_6375);
or U8041 (N_8041,N_6857,N_6711);
nand U8042 (N_8042,N_7078,N_7264);
or U8043 (N_8043,N_7392,N_7663);
and U8044 (N_8044,N_7940,N_7360);
nor U8045 (N_8045,N_7928,N_6988);
and U8046 (N_8046,N_6362,N_6984);
nand U8047 (N_8047,N_7978,N_6467);
or U8048 (N_8048,N_6794,N_6422);
nor U8049 (N_8049,N_6000,N_7676);
nand U8050 (N_8050,N_7790,N_6617);
nand U8051 (N_8051,N_6424,N_7755);
xnor U8052 (N_8052,N_6914,N_6572);
and U8053 (N_8053,N_7910,N_7829);
or U8054 (N_8054,N_6129,N_7254);
and U8055 (N_8055,N_7226,N_6344);
nor U8056 (N_8056,N_7446,N_6287);
nand U8057 (N_8057,N_7354,N_6067);
nand U8058 (N_8058,N_7263,N_6671);
or U8059 (N_8059,N_7939,N_7693);
nor U8060 (N_8060,N_6428,N_7794);
nand U8061 (N_8061,N_6638,N_6753);
nand U8062 (N_8062,N_7275,N_7420);
nor U8063 (N_8063,N_6048,N_7168);
and U8064 (N_8064,N_7678,N_7748);
or U8065 (N_8065,N_7007,N_7863);
nor U8066 (N_8066,N_6594,N_7712);
nand U8067 (N_8067,N_6586,N_6683);
or U8068 (N_8068,N_6414,N_7329);
nor U8069 (N_8069,N_7905,N_7488);
or U8070 (N_8070,N_7458,N_7799);
nor U8071 (N_8071,N_7784,N_7970);
xnor U8072 (N_8072,N_7289,N_6913);
nor U8073 (N_8073,N_7816,N_6839);
nor U8074 (N_8074,N_7362,N_6262);
nand U8075 (N_8075,N_7723,N_6416);
nand U8076 (N_8076,N_7690,N_7942);
and U8077 (N_8077,N_6775,N_7958);
and U8078 (N_8078,N_7069,N_6783);
nand U8079 (N_8079,N_6894,N_6955);
or U8080 (N_8080,N_7839,N_7417);
and U8081 (N_8081,N_6282,N_7067);
and U8082 (N_8082,N_6846,N_7396);
nand U8083 (N_8083,N_7886,N_6249);
and U8084 (N_8084,N_7130,N_7283);
nand U8085 (N_8085,N_7951,N_6611);
or U8086 (N_8086,N_7843,N_6435);
nand U8087 (N_8087,N_7047,N_7441);
or U8088 (N_8088,N_7639,N_6363);
and U8089 (N_8089,N_7623,N_6652);
or U8090 (N_8090,N_7614,N_6041);
nor U8091 (N_8091,N_7604,N_7452);
and U8092 (N_8092,N_6648,N_7398);
nor U8093 (N_8093,N_7222,N_7974);
and U8094 (N_8094,N_7459,N_6633);
xor U8095 (N_8095,N_6620,N_6799);
or U8096 (N_8096,N_6474,N_7897);
and U8097 (N_8097,N_7016,N_6644);
and U8098 (N_8098,N_7785,N_6766);
or U8099 (N_8099,N_7310,N_7625);
nand U8100 (N_8100,N_7238,N_7397);
nand U8101 (N_8101,N_7428,N_6463);
nor U8102 (N_8102,N_6593,N_7662);
and U8103 (N_8103,N_7056,N_7110);
or U8104 (N_8104,N_6286,N_7746);
and U8105 (N_8105,N_6272,N_6090);
nor U8106 (N_8106,N_6551,N_7462);
xor U8107 (N_8107,N_7554,N_7334);
nor U8108 (N_8108,N_7369,N_6953);
nor U8109 (N_8109,N_7709,N_6057);
nand U8110 (N_8110,N_7135,N_6827);
nor U8111 (N_8111,N_6316,N_6401);
and U8112 (N_8112,N_7282,N_7044);
or U8113 (N_8113,N_7483,N_7927);
nor U8114 (N_8114,N_7911,N_6693);
nor U8115 (N_8115,N_7500,N_6771);
or U8116 (N_8116,N_6182,N_7896);
or U8117 (N_8117,N_6636,N_6815);
and U8118 (N_8118,N_6074,N_7553);
nor U8119 (N_8119,N_6060,N_6929);
nand U8120 (N_8120,N_7118,N_7648);
and U8121 (N_8121,N_7477,N_6616);
and U8122 (N_8122,N_7482,N_6024);
and U8123 (N_8123,N_7518,N_7813);
and U8124 (N_8124,N_6842,N_7058);
nand U8125 (N_8125,N_6211,N_6682);
or U8126 (N_8126,N_6145,N_6570);
and U8127 (N_8127,N_7895,N_7570);
and U8128 (N_8128,N_7125,N_7317);
nor U8129 (N_8129,N_6342,N_7624);
or U8130 (N_8130,N_7032,N_6947);
nor U8131 (N_8131,N_6904,N_7001);
nor U8132 (N_8132,N_6626,N_6780);
nand U8133 (N_8133,N_7628,N_6426);
nand U8134 (N_8134,N_6849,N_6115);
nor U8135 (N_8135,N_7277,N_7425);
nor U8136 (N_8136,N_6530,N_6635);
and U8137 (N_8137,N_7929,N_6095);
nor U8138 (N_8138,N_7853,N_6687);
nor U8139 (N_8139,N_7361,N_6531);
nand U8140 (N_8140,N_7729,N_6834);
or U8141 (N_8141,N_7117,N_6924);
and U8142 (N_8142,N_6823,N_6196);
nor U8143 (N_8143,N_6037,N_6198);
nand U8144 (N_8144,N_6816,N_6867);
or U8145 (N_8145,N_6480,N_7004);
nand U8146 (N_8146,N_6229,N_6388);
nor U8147 (N_8147,N_6721,N_7564);
or U8148 (N_8148,N_6575,N_7963);
or U8149 (N_8149,N_6240,N_7860);
or U8150 (N_8150,N_6308,N_7739);
nand U8151 (N_8151,N_7126,N_7116);
nor U8152 (N_8152,N_7212,N_6529);
nand U8153 (N_8153,N_7364,N_6012);
or U8154 (N_8154,N_7260,N_7022);
nor U8155 (N_8155,N_6535,N_7062);
and U8156 (N_8156,N_7342,N_7506);
and U8157 (N_8157,N_7399,N_6772);
nand U8158 (N_8158,N_6997,N_7550);
nor U8159 (N_8159,N_6374,N_6907);
or U8160 (N_8160,N_7495,N_7584);
nand U8161 (N_8161,N_6665,N_6136);
and U8162 (N_8162,N_6452,N_6847);
nor U8163 (N_8163,N_6478,N_7844);
and U8164 (N_8164,N_6039,N_6437);
and U8165 (N_8165,N_6759,N_6716);
and U8166 (N_8166,N_6054,N_7981);
and U8167 (N_8167,N_6710,N_6011);
nand U8168 (N_8168,N_6325,N_7138);
nor U8169 (N_8169,N_7965,N_6122);
or U8170 (N_8170,N_7188,N_6444);
nor U8171 (N_8171,N_6335,N_6887);
and U8172 (N_8172,N_7228,N_7340);
or U8173 (N_8173,N_6553,N_6393);
nand U8174 (N_8174,N_7487,N_7795);
and U8175 (N_8175,N_6172,N_7923);
and U8176 (N_8176,N_6820,N_6059);
nor U8177 (N_8177,N_6538,N_6879);
and U8178 (N_8178,N_6852,N_6659);
or U8179 (N_8179,N_6808,N_6315);
nor U8180 (N_8180,N_6187,N_7450);
and U8181 (N_8181,N_6925,N_6077);
nor U8182 (N_8182,N_7599,N_7652);
nor U8183 (N_8183,N_6173,N_7345);
nor U8184 (N_8184,N_6778,N_6151);
xnor U8185 (N_8185,N_7589,N_7924);
nand U8186 (N_8186,N_7983,N_7586);
and U8187 (N_8187,N_7962,N_6974);
and U8188 (N_8188,N_6893,N_7694);
nand U8189 (N_8189,N_6697,N_6811);
nor U8190 (N_8190,N_6105,N_7592);
or U8191 (N_8191,N_6134,N_7123);
nand U8192 (N_8192,N_7808,N_7665);
or U8193 (N_8193,N_7559,N_7865);
nor U8194 (N_8194,N_7852,N_6514);
nor U8195 (N_8195,N_6571,N_7869);
and U8196 (N_8196,N_7018,N_6297);
and U8197 (N_8197,N_6154,N_7894);
or U8198 (N_8198,N_6641,N_6776);
nand U8199 (N_8199,N_6471,N_7594);
nor U8200 (N_8200,N_6554,N_7390);
and U8201 (N_8201,N_6186,N_6918);
nor U8202 (N_8202,N_6838,N_7498);
nor U8203 (N_8203,N_7421,N_7404);
and U8204 (N_8204,N_6167,N_7697);
nor U8205 (N_8205,N_6114,N_6515);
nor U8206 (N_8206,N_6564,N_7992);
nor U8207 (N_8207,N_7967,N_6273);
nor U8208 (N_8208,N_7840,N_6208);
and U8209 (N_8209,N_7753,N_6911);
nand U8210 (N_8210,N_7292,N_6333);
or U8211 (N_8211,N_7683,N_6391);
nand U8212 (N_8212,N_6817,N_6858);
and U8213 (N_8213,N_7834,N_6327);
and U8214 (N_8214,N_6432,N_6826);
and U8215 (N_8215,N_7847,N_6083);
nor U8216 (N_8216,N_7305,N_7347);
and U8217 (N_8217,N_7257,N_6619);
and U8218 (N_8218,N_7447,N_7637);
or U8219 (N_8219,N_6035,N_6091);
nor U8220 (N_8220,N_6102,N_7177);
or U8221 (N_8221,N_6113,N_6928);
nor U8222 (N_8222,N_7537,N_6562);
nor U8223 (N_8223,N_6739,N_6313);
or U8224 (N_8224,N_6409,N_7268);
nor U8225 (N_8225,N_7621,N_7395);
or U8226 (N_8226,N_7908,N_7657);
nand U8227 (N_8227,N_6675,N_7875);
nor U8228 (N_8228,N_7680,N_7837);
nand U8229 (N_8229,N_6653,N_6770);
nor U8230 (N_8230,N_7405,N_6413);
nand U8231 (N_8231,N_7609,N_7706);
and U8232 (N_8232,N_6518,N_7540);
or U8233 (N_8233,N_6292,N_7862);
and U8234 (N_8234,N_7164,N_7877);
and U8235 (N_8235,N_7687,N_7473);
and U8236 (N_8236,N_7146,N_6298);
or U8237 (N_8237,N_7351,N_7669);
and U8238 (N_8238,N_7195,N_6268);
or U8239 (N_8239,N_6439,N_7162);
nor U8240 (N_8240,N_6940,N_6052);
nand U8241 (N_8241,N_6258,N_7357);
and U8242 (N_8242,N_7095,N_7957);
or U8243 (N_8243,N_7376,N_6504);
nand U8244 (N_8244,N_7603,N_7109);
nor U8245 (N_8245,N_6881,N_7516);
nor U8246 (N_8246,N_6423,N_6120);
nand U8247 (N_8247,N_7976,N_7722);
and U8248 (N_8248,N_7804,N_7131);
or U8249 (N_8249,N_7841,N_6361);
nor U8250 (N_8250,N_6880,N_7655);
nand U8251 (N_8251,N_7855,N_7251);
or U8252 (N_8252,N_6921,N_7899);
or U8253 (N_8253,N_6436,N_7120);
or U8254 (N_8254,N_6053,N_6473);
nor U8255 (N_8255,N_7243,N_7702);
nor U8256 (N_8256,N_7122,N_7239);
nor U8257 (N_8257,N_7322,N_7736);
nand U8258 (N_8258,N_7008,N_7543);
nand U8259 (N_8259,N_6384,N_6031);
and U8260 (N_8260,N_7793,N_7527);
and U8261 (N_8261,N_7033,N_7779);
or U8262 (N_8262,N_6969,N_7596);
or U8263 (N_8263,N_7371,N_7968);
nor U8264 (N_8264,N_7223,N_6336);
nand U8265 (N_8265,N_6560,N_6242);
nor U8266 (N_8266,N_6625,N_6699);
nand U8267 (N_8267,N_6642,N_6740);
or U8268 (N_8268,N_7290,N_6797);
nor U8269 (N_8269,N_7355,N_6156);
nand U8270 (N_8270,N_6294,N_7020);
and U8271 (N_8271,N_7535,N_7832);
nor U8272 (N_8272,N_6946,N_6519);
and U8273 (N_8273,N_6814,N_7196);
nand U8274 (N_8274,N_7526,N_6548);
nand U8275 (N_8275,N_6807,N_6995);
or U8276 (N_8276,N_7469,N_6910);
or U8277 (N_8277,N_6981,N_6343);
and U8278 (N_8278,N_6830,N_6786);
and U8279 (N_8279,N_6590,N_6749);
nor U8280 (N_8280,N_7576,N_7904);
or U8281 (N_8281,N_6107,N_7088);
and U8282 (N_8282,N_7437,N_6614);
or U8283 (N_8283,N_6457,N_6263);
nand U8284 (N_8284,N_6378,N_6868);
or U8285 (N_8285,N_6859,N_7316);
and U8286 (N_8286,N_6222,N_6502);
or U8287 (N_8287,N_6466,N_6900);
and U8288 (N_8288,N_6585,N_7103);
or U8289 (N_8289,N_7378,N_6782);
nand U8290 (N_8290,N_7472,N_7485);
and U8291 (N_8291,N_7703,N_7070);
or U8292 (N_8292,N_6104,N_6791);
nand U8293 (N_8293,N_6305,N_7689);
and U8294 (N_8294,N_7943,N_7618);
nand U8295 (N_8295,N_7312,N_6055);
or U8296 (N_8296,N_7999,N_6366);
nand U8297 (N_8297,N_6591,N_7756);
nor U8298 (N_8298,N_7269,N_6341);
or U8299 (N_8299,N_7271,N_7991);
nor U8300 (N_8300,N_7913,N_6364);
nand U8301 (N_8301,N_6014,N_7780);
nand U8302 (N_8302,N_7023,N_6709);
nor U8303 (N_8303,N_7466,N_6103);
or U8304 (N_8304,N_7011,N_6631);
nor U8305 (N_8305,N_6021,N_7040);
nor U8306 (N_8306,N_7724,N_7806);
or U8307 (N_8307,N_6277,N_7867);
xor U8308 (N_8308,N_6661,N_7097);
or U8309 (N_8309,N_7936,N_6898);
and U8310 (N_8310,N_7424,N_6030);
nor U8311 (N_8311,N_7045,N_6080);
nor U8312 (N_8312,N_7906,N_6891);
nand U8313 (N_8313,N_7169,N_6809);
and U8314 (N_8314,N_7003,N_7511);
nor U8315 (N_8315,N_7769,N_6528);
and U8316 (N_8316,N_7575,N_7165);
nor U8317 (N_8317,N_7871,N_6756);
and U8318 (N_8318,N_7650,N_6882);
or U8319 (N_8319,N_6679,N_7760);
and U8320 (N_8320,N_6195,N_6610);
nor U8321 (N_8321,N_6472,N_6408);
and U8322 (N_8322,N_6726,N_7328);
nor U8323 (N_8323,N_6453,N_7330);
or U8324 (N_8324,N_6563,N_7734);
nand U8325 (N_8325,N_6431,N_7633);
and U8326 (N_8326,N_6257,N_6399);
nor U8327 (N_8327,N_6832,N_6952);
nand U8328 (N_8328,N_6274,N_6523);
or U8329 (N_8329,N_7595,N_6704);
or U8330 (N_8330,N_6744,N_7876);
nand U8331 (N_8331,N_7587,N_6445);
and U8332 (N_8332,N_7985,N_6061);
nor U8333 (N_8333,N_6118,N_6330);
and U8334 (N_8334,N_6128,N_7552);
nor U8335 (N_8335,N_6833,N_7947);
nor U8336 (N_8336,N_7732,N_7253);
and U8337 (N_8337,N_6958,N_7572);
and U8338 (N_8338,N_7366,N_6130);
and U8339 (N_8339,N_6584,N_7274);
and U8340 (N_8340,N_7737,N_7901);
nor U8341 (N_8341,N_7339,N_6433);
nand U8342 (N_8342,N_6792,N_7812);
and U8343 (N_8343,N_7438,N_6957);
or U8344 (N_8344,N_6036,N_6696);
or U8345 (N_8345,N_6695,N_6214);
nand U8346 (N_8346,N_7854,N_6993);
nand U8347 (N_8347,N_6806,N_7076);
and U8348 (N_8348,N_7463,N_7810);
nand U8349 (N_8349,N_6684,N_7142);
nand U8350 (N_8350,N_6835,N_7960);
and U8351 (N_8351,N_7815,N_7479);
nand U8352 (N_8352,N_6171,N_7333);
nand U8353 (N_8353,N_7558,N_6906);
nor U8354 (N_8354,N_7075,N_7027);
nor U8355 (N_8355,N_7645,N_7807);
nand U8356 (N_8356,N_7866,N_7825);
or U8357 (N_8357,N_7764,N_6875);
or U8358 (N_8358,N_6561,N_6322);
and U8359 (N_8359,N_7250,N_6395);
and U8360 (N_8360,N_7338,N_6420);
nand U8361 (N_8361,N_6812,N_7197);
and U8362 (N_8362,N_6752,N_6403);
xnor U8363 (N_8363,N_7982,N_7156);
nor U8364 (N_8364,N_6009,N_7884);
nand U8365 (N_8365,N_6600,N_6549);
or U8366 (N_8366,N_6367,N_6008);
and U8367 (N_8367,N_6318,N_6398);
nand U8368 (N_8368,N_7372,N_6559);
nand U8369 (N_8369,N_6417,N_7814);
or U8370 (N_8370,N_7221,N_7607);
nor U8371 (N_8371,N_6966,N_6200);
or U8372 (N_8372,N_6674,N_7523);
nor U8373 (N_8373,N_7585,N_6650);
nor U8374 (N_8374,N_6701,N_7105);
or U8375 (N_8375,N_6720,N_6734);
and U8376 (N_8376,N_7386,N_6654);
nor U8377 (N_8377,N_7445,N_7050);
and U8378 (N_8378,N_6438,N_7730);
nand U8379 (N_8379,N_7509,N_6233);
and U8380 (N_8380,N_6479,N_7817);
and U8381 (N_8381,N_6542,N_6836);
nand U8382 (N_8382,N_6582,N_6270);
or U8383 (N_8383,N_7335,N_7528);
nand U8384 (N_8384,N_7562,N_7101);
nand U8385 (N_8385,N_7949,N_7115);
and U8386 (N_8386,N_7842,N_7434);
nand U8387 (N_8387,N_7719,N_6784);
nor U8388 (N_8388,N_6864,N_7107);
nand U8389 (N_8389,N_6916,N_6058);
nand U8390 (N_8390,N_7944,N_7577);
nor U8391 (N_8391,N_7063,N_7267);
nand U8392 (N_8392,N_6228,N_6979);
nand U8393 (N_8393,N_6093,N_7430);
nor U8394 (N_8394,N_7163,N_6179);
or U8395 (N_8395,N_6755,N_6482);
or U8396 (N_8396,N_6948,N_7819);
nor U8397 (N_8397,N_6539,N_6429);
nor U8398 (N_8398,N_7072,N_7049);
xor U8399 (N_8399,N_7311,N_6081);
nor U8400 (N_8400,N_7181,N_7419);
nor U8401 (N_8401,N_6392,N_7224);
or U8402 (N_8402,N_7295,N_6764);
or U8403 (N_8403,N_6804,N_7851);
and U8404 (N_8404,N_6760,N_6248);
nand U8405 (N_8405,N_7993,N_7051);
or U8406 (N_8406,N_7489,N_7240);
or U8407 (N_8407,N_7104,N_6691);
or U8408 (N_8408,N_7619,N_7077);
nor U8409 (N_8409,N_6727,N_6862);
nand U8410 (N_8410,N_7931,N_6522);
nor U8411 (N_8411,N_7979,N_6267);
and U8412 (N_8412,N_7214,N_7280);
nor U8413 (N_8413,N_7580,N_7997);
nand U8414 (N_8414,N_7213,N_6998);
nand U8415 (N_8415,N_6731,N_7747);
and U8416 (N_8416,N_6983,N_6124);
nand U8417 (N_8417,N_6581,N_7121);
nor U8418 (N_8418,N_6781,N_6291);
nor U8419 (N_8419,N_7315,N_6493);
or U8420 (N_8420,N_7711,N_7776);
and U8421 (N_8421,N_7173,N_6533);
and U8422 (N_8422,N_7442,N_7898);
nand U8423 (N_8423,N_6745,N_7531);
or U8424 (N_8424,N_7391,N_7757);
nand U8425 (N_8425,N_6069,N_7612);
and U8426 (N_8426,N_7634,N_6527);
and U8427 (N_8427,N_6829,N_6450);
xor U8428 (N_8428,N_7758,N_6131);
or U8429 (N_8429,N_6853,N_7341);
and U8430 (N_8430,N_7917,N_7377);
nand U8431 (N_8431,N_6044,N_7581);
nor U8432 (N_8432,N_6459,N_6877);
or U8433 (N_8433,N_6427,N_7845);
and U8434 (N_8434,N_7891,N_6996);
nor U8435 (N_8435,N_6148,N_6138);
and U8436 (N_8436,N_6337,N_7919);
nor U8437 (N_8437,N_7824,N_6304);
or U8438 (N_8438,N_7620,N_7933);
or U8439 (N_8439,N_6802,N_7856);
or U8440 (N_8440,N_6328,N_6841);
and U8441 (N_8441,N_6369,N_6458);
nand U8442 (N_8442,N_7468,N_6608);
nor U8443 (N_8443,N_7231,N_6796);
or U8444 (N_8444,N_7191,N_6288);
nor U8445 (N_8445,N_6331,N_7414);
or U8446 (N_8446,N_7060,N_6855);
and U8447 (N_8447,N_7089,N_6181);
or U8448 (N_8448,N_7133,N_7359);
nand U8449 (N_8449,N_7200,N_7034);
xnor U8450 (N_8450,N_6219,N_6729);
and U8451 (N_8451,N_6845,N_6098);
or U8452 (N_8452,N_6246,N_7912);
or U8453 (N_8453,N_6798,N_6380);
and U8454 (N_8454,N_7336,N_7486);
and U8455 (N_8455,N_6213,N_7696);
or U8456 (N_8456,N_6987,N_6897);
and U8457 (N_8457,N_6954,N_6492);
or U8458 (N_8458,N_6447,N_6871);
nand U8459 (N_8459,N_6822,N_7323);
or U8460 (N_8460,N_6649,N_6425);
nor U8461 (N_8461,N_6100,N_7520);
nand U8462 (N_8462,N_6464,N_6892);
nand U8463 (N_8463,N_6092,N_6597);
and U8464 (N_8464,N_6777,N_7515);
nand U8465 (N_8465,N_6499,N_7211);
nor U8466 (N_8466,N_6547,N_7504);
nand U8467 (N_8467,N_6884,N_7611);
nor U8468 (N_8468,N_6461,N_6247);
nand U8469 (N_8469,N_6170,N_7954);
or U8470 (N_8470,N_6117,N_7966);
nor U8471 (N_8471,N_6005,N_6303);
and U8472 (N_8472,N_6669,N_6501);
nor U8473 (N_8473,N_7471,N_7140);
nor U8474 (N_8474,N_6174,N_7788);
or U8475 (N_8475,N_7512,N_7881);
nand U8476 (N_8476,N_6446,N_7846);
and U8477 (N_8477,N_6338,N_7206);
nor U8478 (N_8478,N_6986,N_6801);
nor U8479 (N_8479,N_7582,N_6935);
or U8480 (N_8480,N_6462,N_7684);
nand U8481 (N_8481,N_7945,N_6566);
or U8482 (N_8482,N_7084,N_7382);
nand U8483 (N_8483,N_7643,N_6296);
and U8484 (N_8484,N_6544,N_6738);
nor U8485 (N_8485,N_7474,N_7266);
and U8486 (N_8486,N_6899,N_7741);
and U8487 (N_8487,N_7679,N_6099);
or U8488 (N_8488,N_7613,N_6106);
nand U8489 (N_8489,N_7108,N_6576);
and U8490 (N_8490,N_7086,N_6965);
nor U8491 (N_8491,N_7098,N_6536);
and U8492 (N_8492,N_6116,N_6565);
and U8493 (N_8493,N_7176,N_7907);
and U8494 (N_8494,N_6854,N_7134);
and U8495 (N_8495,N_7183,N_7654);
and U8496 (N_8496,N_7774,N_7179);
and U8497 (N_8497,N_7319,N_7522);
and U8498 (N_8498,N_7887,N_7490);
nand U8499 (N_8499,N_7946,N_6767);
and U8500 (N_8500,N_6511,N_6878);
nand U8501 (N_8501,N_6700,N_7367);
and U8502 (N_8502,N_7216,N_7092);
or U8503 (N_8503,N_6629,N_6469);
and U8504 (N_8504,N_6056,N_6137);
or U8505 (N_8505,N_7809,N_7850);
nor U8506 (N_8506,N_6033,N_7157);
nand U8507 (N_8507,N_6750,N_7144);
nor U8508 (N_8508,N_6236,N_7670);
or U8509 (N_8509,N_6567,N_6956);
and U8510 (N_8510,N_6598,N_7080);
nand U8511 (N_8511,N_7128,N_6359);
nor U8512 (N_8512,N_6254,N_7343);
and U8513 (N_8513,N_6803,N_7448);
nand U8514 (N_8514,N_6002,N_6078);
nand U8515 (N_8515,N_6349,N_7667);
nor U8516 (N_8516,N_7496,N_6027);
and U8517 (N_8517,N_7743,N_7557);
nand U8518 (N_8518,N_7219,N_6917);
and U8519 (N_8519,N_7259,N_7754);
and U8520 (N_8520,N_6517,N_7470);
or U8521 (N_8521,N_7174,N_6615);
or U8522 (N_8522,N_7969,N_7262);
nand U8523 (N_8523,N_6460,N_7309);
or U8524 (N_8524,N_6231,N_7041);
or U8525 (N_8525,N_6189,N_7478);
nand U8526 (N_8526,N_7158,N_6264);
and U8527 (N_8527,N_6097,N_7087);
nand U8528 (N_8528,N_6722,N_7781);
or U8529 (N_8529,N_7900,N_6394);
nor U8530 (N_8530,N_6255,N_6084);
or U8531 (N_8531,N_7307,N_7858);
nor U8532 (N_8532,N_6730,N_6640);
and U8533 (N_8533,N_7256,N_7868);
and U8534 (N_8534,N_7597,N_6178);
and U8535 (N_8535,N_6510,N_7726);
xor U8536 (N_8536,N_6415,N_7569);
nor U8537 (N_8537,N_6658,N_7998);
nor U8538 (N_8538,N_7356,N_6164);
or U8539 (N_8539,N_6662,N_7590);
nand U8540 (N_8540,N_6079,N_7751);
nor U8541 (N_8541,N_6051,N_7833);
or U8542 (N_8542,N_6605,N_6550);
and U8543 (N_8543,N_7061,N_6184);
nand U8544 (N_8544,N_6112,N_7503);
nor U8545 (N_8545,N_6483,N_7827);
or U8546 (N_8546,N_6588,N_6221);
or U8547 (N_8547,N_6193,N_6111);
and U8548 (N_8548,N_6951,N_6089);
nor U8549 (N_8549,N_6158,N_6634);
and U8550 (N_8550,N_7300,N_6863);
and U8551 (N_8551,N_6942,N_6937);
or U8552 (N_8552,N_7325,N_7857);
or U8553 (N_8553,N_6681,N_7956);
or U8554 (N_8554,N_7301,N_6500);
or U8555 (N_8555,N_6314,N_6609);
nand U8556 (N_8556,N_7952,N_6162);
nand U8557 (N_8557,N_6520,N_6612);
or U8558 (N_8558,N_7948,N_6793);
or U8559 (N_8559,N_6876,N_6306);
nand U8560 (N_8560,N_7698,N_7205);
or U8561 (N_8561,N_6348,N_6150);
xnor U8562 (N_8562,N_6795,N_6127);
or U8563 (N_8563,N_6225,N_6360);
and U8564 (N_8564,N_7805,N_6140);
or U8565 (N_8565,N_6324,N_6261);
and U8566 (N_8566,N_6319,N_7454);
and U8567 (N_8567,N_6923,N_6788);
and U8568 (N_8568,N_7765,N_7830);
nand U8569 (N_8569,N_6715,N_7984);
nand U8570 (N_8570,N_6774,N_7731);
nor U8571 (N_8571,N_6373,N_6505);
and U8572 (N_8572,N_7529,N_6843);
nor U8573 (N_8573,N_6144,N_7385);
nand U8574 (N_8574,N_7995,N_6350);
and U8575 (N_8575,N_7068,N_7874);
or U8576 (N_8576,N_6234,N_6339);
nor U8577 (N_8577,N_6779,N_6741);
and U8578 (N_8578,N_7166,N_7210);
nor U8579 (N_8579,N_6534,N_7986);
or U8580 (N_8580,N_6326,N_6824);
or U8581 (N_8581,N_6238,N_7826);
and U8582 (N_8582,N_6583,N_6323);
nor U8583 (N_8583,N_7031,N_6023);
nand U8584 (N_8584,N_6390,N_6441);
nor U8585 (N_8585,N_7872,N_7926);
and U8586 (N_8586,N_6279,N_6207);
and U8587 (N_8587,N_7801,N_6627);
nand U8588 (N_8588,N_6702,N_7838);
or U8589 (N_8589,N_7167,N_6110);
and U8590 (N_8590,N_6025,N_7770);
or U8591 (N_8591,N_6412,N_7823);
nand U8592 (N_8592,N_6475,N_6637);
and U8593 (N_8593,N_6216,N_6289);
nor U8594 (N_8594,N_6142,N_6299);
nand U8595 (N_8595,N_7288,N_6604);
and U8596 (N_8596,N_6206,N_7849);
and U8597 (N_8597,N_7431,N_6404);
nor U8598 (N_8598,N_6660,N_6736);
or U8599 (N_8599,N_6503,N_7453);
xnor U8600 (N_8600,N_7201,N_7090);
nor U8601 (N_8601,N_6623,N_7111);
or U8602 (N_8602,N_7773,N_7727);
or U8603 (N_8603,N_7642,N_6411);
or U8604 (N_8604,N_7218,N_7460);
nand U8605 (N_8605,N_7096,N_7400);
and U8606 (N_8606,N_6663,N_7038);
nor U8607 (N_8607,N_7079,N_6552);
nor U8608 (N_8608,N_6132,N_6400);
and U8609 (N_8609,N_7494,N_6028);
nor U8610 (N_8610,N_7880,N_7291);
or U8611 (N_8611,N_7715,N_7627);
nor U8612 (N_8612,N_6334,N_6271);
or U8613 (N_8613,N_7091,N_6241);
nor U8614 (N_8614,N_6844,N_6082);
nand U8615 (N_8615,N_7457,N_6194);
and U8616 (N_8616,N_7902,N_6218);
xnor U8617 (N_8617,N_6320,N_6227);
and U8618 (N_8618,N_6295,N_6494);
or U8619 (N_8619,N_6293,N_6743);
and U8620 (N_8620,N_7740,N_7710);
nand U8621 (N_8621,N_7811,N_7775);
and U8622 (N_8622,N_6197,N_6901);
nor U8623 (N_8623,N_6513,N_6758);
and U8624 (N_8624,N_7321,N_7566);
or U8625 (N_8625,N_7203,N_6013);
nand U8626 (N_8626,N_7975,N_7082);
and U8627 (N_8627,N_7102,N_7065);
or U8628 (N_8628,N_7888,N_6183);
xor U8629 (N_8629,N_6352,N_6332);
nor U8630 (N_8630,N_6905,N_6309);
or U8631 (N_8631,N_6595,N_7346);
nand U8632 (N_8632,N_6963,N_6902);
or U8633 (N_8633,N_7217,N_7890);
nand U8634 (N_8634,N_6224,N_7818);
nand U8635 (N_8635,N_7761,N_7039);
nor U8636 (N_8636,N_6096,N_7410);
and U8637 (N_8637,N_7605,N_7297);
or U8638 (N_8638,N_7681,N_7971);
nand U8639 (N_8639,N_6861,N_7284);
and U8640 (N_8640,N_7759,N_7682);
nor U8641 (N_8641,N_6992,N_7567);
and U8642 (N_8642,N_6789,N_6269);
or U8643 (N_8643,N_6389,N_7556);
nand U8644 (N_8644,N_6888,N_7583);
and U8645 (N_8645,N_7426,N_6018);
nor U8646 (N_8646,N_7416,N_6599);
or U8647 (N_8647,N_7293,N_7057);
or U8648 (N_8648,N_6454,N_7387);
or U8649 (N_8649,N_6205,N_7215);
or U8650 (N_8650,N_6161,N_6147);
nor U8651 (N_8651,N_7934,N_6382);
and U8652 (N_8652,N_7870,N_6558);
nor U8653 (N_8653,N_6930,N_6125);
nor U8654 (N_8654,N_6908,N_6126);
and U8655 (N_8655,N_6386,N_6769);
and U8656 (N_8656,N_6250,N_6883);
and U8657 (N_8657,N_7432,N_7249);
nand U8658 (N_8658,N_7010,N_6284);
or U8659 (N_8659,N_6668,N_7738);
nor U8660 (N_8660,N_7246,N_7252);
or U8661 (N_8661,N_6577,N_7182);
nor U8662 (N_8662,N_6139,N_6050);
nor U8663 (N_8663,N_7074,N_7248);
or U8664 (N_8664,N_7530,N_6713);
nor U8665 (N_8665,N_7408,N_7199);
or U8666 (N_8666,N_6580,N_6714);
or U8667 (N_8667,N_7145,N_7800);
nand U8668 (N_8668,N_7278,N_7407);
or U8669 (N_8669,N_6088,N_6532);
nor U8670 (N_8670,N_7147,N_7972);
xor U8671 (N_8671,N_6985,N_6230);
or U8672 (N_8672,N_6010,N_6541);
nand U8673 (N_8673,N_6746,N_6040);
and U8674 (N_8674,N_7545,N_7402);
nor U8675 (N_8675,N_7279,N_6982);
and U8676 (N_8676,N_7538,N_6280);
nor U8677 (N_8677,N_6639,N_6470);
nand U8678 (N_8678,N_6869,N_7042);
nor U8679 (N_8679,N_6410,N_6964);
or U8680 (N_8680,N_6075,N_7053);
nor U8681 (N_8681,N_7071,N_6889);
or U8682 (N_8682,N_6210,N_7836);
or U8683 (N_8683,N_6705,N_7409);
or U8684 (N_8684,N_7571,N_6909);
nand U8685 (N_8685,N_6163,N_7433);
nor U8686 (N_8686,N_6828,N_6149);
or U8687 (N_8687,N_7568,N_7720);
and U8688 (N_8688,N_7155,N_7054);
nand U8689 (N_8689,N_7422,N_7306);
and U8690 (N_8690,N_7178,N_7046);
nor U8691 (N_8691,N_7803,N_6667);
nor U8692 (N_8692,N_7501,N_7413);
or U8693 (N_8693,N_7318,N_7112);
or U8694 (N_8694,N_7194,N_6354);
or U8695 (N_8695,N_7024,N_7644);
nand U8696 (N_8696,N_6922,N_7427);
and U8697 (N_8697,N_6387,N_7245);
and U8698 (N_8698,N_7412,N_7659);
nor U8699 (N_8699,N_6451,N_7352);
or U8700 (N_8700,N_7822,N_7955);
and U8701 (N_8701,N_7332,N_6317);
or U8702 (N_8702,N_7510,N_7602);
nand U8703 (N_8703,N_7465,N_6175);
nand U8704 (N_8704,N_7789,N_7415);
xor U8705 (N_8705,N_7691,N_6119);
or U8706 (N_8706,N_7270,N_6723);
or U8707 (N_8707,N_7429,N_6724);
and U8708 (N_8708,N_6311,N_7187);
or U8709 (N_8709,N_7508,N_7658);
and U8710 (N_8710,N_6190,N_6961);
nand U8711 (N_8711,N_6978,N_7513);
or U8712 (N_8712,N_7021,N_7656);
and U8713 (N_8713,N_7521,N_6490);
nand U8714 (N_8714,N_6166,N_7517);
nand U8715 (N_8715,N_6256,N_7705);
nor U8716 (N_8716,N_7052,N_7925);
and U8717 (N_8717,N_6212,N_7327);
nor U8718 (N_8718,N_7373,N_6448);
or U8719 (N_8719,N_6959,N_6232);
nand U8720 (N_8720,N_7873,N_6540);
or U8721 (N_8721,N_7265,N_7326);
and U8722 (N_8722,N_6860,N_7186);
or U8723 (N_8723,N_6143,N_7533);
nor U8724 (N_8724,N_7380,N_6307);
and U8725 (N_8725,N_6719,N_7532);
nand U8726 (N_8726,N_7961,N_6485);
nor U8727 (N_8727,N_7258,N_6972);
nand U8728 (N_8728,N_6169,N_6022);
nand U8729 (N_8729,N_7752,N_6927);
or U8730 (N_8730,N_7247,N_6168);
and U8731 (N_8731,N_6926,N_7384);
nand U8732 (N_8732,N_7237,N_7574);
nand U8733 (N_8733,N_6990,N_6047);
and U8734 (N_8734,N_7700,N_7651);
and U8735 (N_8735,N_7579,N_6133);
and U8736 (N_8736,N_7725,N_7921);
nand U8737 (N_8737,N_7006,N_6971);
and U8738 (N_8738,N_6601,N_7353);
xnor U8739 (N_8739,N_6831,N_7236);
and U8740 (N_8740,N_7771,N_6773);
or U8741 (N_8741,N_6896,N_7389);
nand U8742 (N_8742,N_6063,N_6146);
and U8743 (N_8743,N_6545,N_7094);
nand U8744 (N_8744,N_7792,N_7093);
and U8745 (N_8745,N_7916,N_7893);
and U8746 (N_8746,N_7673,N_7615);
and U8747 (N_8747,N_7286,N_7440);
nand U8748 (N_8748,N_7547,N_7802);
or U8749 (N_8749,N_7171,N_7797);
or U8750 (N_8750,N_6606,N_6718);
and U8751 (N_8751,N_6353,N_7677);
nand U8752 (N_8752,N_7744,N_6430);
nor U8753 (N_8753,N_6543,N_6690);
and U8754 (N_8754,N_6819,N_6686);
or U8755 (N_8755,N_7000,N_7475);
nor U8756 (N_8756,N_6488,N_7763);
and U8757 (N_8757,N_7106,N_7443);
nor U8758 (N_8758,N_6874,N_7381);
nor U8759 (N_8759,N_7320,N_6521);
or U8760 (N_8760,N_6655,N_7541);
or U8761 (N_8761,N_7864,N_6498);
and U8762 (N_8762,N_7660,N_7099);
nor U8763 (N_8763,N_6677,N_6643);
nor U8764 (N_8764,N_6573,N_7989);
and U8765 (N_8765,N_7649,N_7914);
nor U8766 (N_8766,N_6751,N_7456);
and U8767 (N_8767,N_6496,N_6943);
nor U8768 (N_8768,N_7996,N_7796);
or U8769 (N_8769,N_6960,N_7148);
nand U8770 (N_8770,N_7546,N_7235);
nor U8771 (N_8771,N_6220,N_6421);
nor U8772 (N_8772,N_7184,N_7699);
nor U8773 (N_8773,N_7403,N_7314);
nand U8774 (N_8774,N_6555,N_6019);
nand U8775 (N_8775,N_6281,N_6152);
or U8776 (N_8776,N_7418,N_7941);
nand U8777 (N_8777,N_6507,N_7578);
or U8778 (N_8778,N_7973,N_7861);
and U8779 (N_8779,N_6670,N_7348);
nand U8780 (N_8780,N_7324,N_7393);
nand U8781 (N_8781,N_6939,N_6856);
nor U8782 (N_8782,N_7745,N_7783);
and U8783 (N_8783,N_7636,N_7638);
nand U8784 (N_8784,N_6121,N_7674);
nor U8785 (N_8785,N_6086,N_6596);
or U8786 (N_8786,N_7451,N_7383);
and U8787 (N_8787,N_6180,N_7551);
nand U8788 (N_8788,N_7692,N_7379);
or U8789 (N_8789,N_7143,N_6252);
and U8790 (N_8790,N_7444,N_6818);
nand U8791 (N_8791,N_6442,N_6840);
and U8792 (N_8792,N_7190,N_7227);
or U8793 (N_8793,N_7151,N_7374);
and U8794 (N_8794,N_6508,N_6226);
or U8795 (N_8795,N_6790,N_7241);
or U8796 (N_8796,N_6991,N_7204);
or U8797 (N_8797,N_6465,N_6578);
and U8798 (N_8798,N_7368,N_6895);
or U8799 (N_8799,N_6931,N_6381);
nor U8800 (N_8800,N_6237,N_7461);
nor U8801 (N_8801,N_6673,N_7641);
or U8802 (N_8802,N_7114,N_6355);
nand U8803 (N_8803,N_7411,N_7064);
nand U8804 (N_8804,N_7647,N_7029);
nand U8805 (N_8805,N_6557,N_7132);
xor U8806 (N_8806,N_6062,N_7035);
and U8807 (N_8807,N_7964,N_7524);
and U8808 (N_8808,N_7539,N_7686);
or U8809 (N_8809,N_6265,N_6785);
and U8810 (N_8810,N_6712,N_7180);
nor U8811 (N_8811,N_6525,N_6688);
or U8812 (N_8812,N_6737,N_7012);
and U8813 (N_8813,N_6886,N_6748);
nor U8814 (N_8814,N_6434,N_7136);
nand U8815 (N_8815,N_7626,N_6630);
nand U8816 (N_8816,N_6516,N_7786);
nand U8817 (N_8817,N_6049,N_6340);
nor U8818 (N_8818,N_6787,N_6312);
nor U8819 (N_8819,N_7388,N_6890);
and U8820 (N_8820,N_6346,N_7152);
nor U8821 (N_8821,N_6251,N_6592);
nand U8822 (N_8822,N_6066,N_7950);
nor U8823 (N_8823,N_6607,N_6477);
nand U8824 (N_8824,N_6042,N_7959);
or U8825 (N_8825,N_7192,N_7401);
nand U8826 (N_8826,N_6933,N_7632);
and U8827 (N_8827,N_7189,N_6487);
nand U8828 (N_8828,N_7514,N_6383);
and U8829 (N_8829,N_6285,N_6397);
or U8830 (N_8830,N_7666,N_7565);
nand U8831 (N_8831,N_6153,N_6017);
xnor U8832 (N_8832,N_7337,N_6624);
nor U8833 (N_8833,N_7721,N_6938);
or U8834 (N_8834,N_6239,N_7349);
or U8835 (N_8835,N_7661,N_7629);
nand U8836 (N_8836,N_6191,N_7059);
nand U8837 (N_8837,N_6372,N_7139);
nand U8838 (N_8838,N_7915,N_6481);
xor U8839 (N_8839,N_6800,N_6356);
or U8840 (N_8840,N_7161,N_7363);
nor U8841 (N_8841,N_6975,N_6509);
nor U8842 (N_8842,N_6283,N_7009);
or U8843 (N_8843,N_7708,N_6537);
or U8844 (N_8844,N_6157,N_6484);
and U8845 (N_8845,N_7882,N_6290);
or U8846 (N_8846,N_6805,N_7977);
nand U8847 (N_8847,N_7081,N_6678);
and U8848 (N_8848,N_7435,N_6376);
and U8849 (N_8849,N_7085,N_7988);
nand U8850 (N_8850,N_6656,N_7015);
nor U8851 (N_8851,N_6377,N_7028);
or U8852 (N_8852,N_7229,N_6569);
and U8853 (N_8853,N_7766,N_6405);
nand U8854 (N_8854,N_7601,N_6821);
or U8855 (N_8855,N_7767,N_6919);
or U8856 (N_8856,N_6177,N_6020);
nand U8857 (N_8857,N_7772,N_7073);
and U8858 (N_8858,N_7119,N_6001);
nor U8859 (N_8859,N_6029,N_6449);
xor U8860 (N_8860,N_7591,N_6949);
xor U8861 (N_8861,N_6260,N_7821);
nand U8862 (N_8862,N_7630,N_7100);
nor U8863 (N_8863,N_7714,N_7640);
and U8864 (N_8864,N_7303,N_7671);
and U8865 (N_8865,N_6708,N_7272);
or U8866 (N_8866,N_7716,N_6851);
or U8867 (N_8867,N_6873,N_7480);
nand U8868 (N_8868,N_6275,N_6945);
nor U8869 (N_8869,N_7980,N_7892);
nand U8870 (N_8870,N_7791,N_7232);
or U8871 (N_8871,N_7185,N_6813);
nand U8872 (N_8872,N_7273,N_6347);
xor U8873 (N_8873,N_6941,N_6108);
xnor U8874 (N_8874,N_7548,N_6546);
and U8875 (N_8875,N_6870,N_6094);
nor U8876 (N_8876,N_6371,N_7113);
and U8877 (N_8877,N_7617,N_6915);
and U8878 (N_8878,N_6968,N_6368);
nor U8879 (N_8879,N_6135,N_6007);
nor U8880 (N_8880,N_6757,N_7713);
or U8881 (N_8881,N_6936,N_7608);
and U8882 (N_8882,N_6015,N_6345);
nor U8883 (N_8883,N_6365,N_7616);
and U8884 (N_8884,N_6223,N_7066);
and U8885 (N_8885,N_7598,N_6070);
or U8886 (N_8886,N_7903,N_6621);
and U8887 (N_8887,N_7883,N_7885);
nand U8888 (N_8888,N_6491,N_7653);
nor U8889 (N_8889,N_7285,N_6999);
nand U8890 (N_8890,N_6486,N_6692);
and U8891 (N_8891,N_6646,N_6735);
and U8892 (N_8892,N_6087,N_6155);
nor U8893 (N_8893,N_7436,N_7365);
and U8894 (N_8894,N_6245,N_7688);
and U8895 (N_8895,N_7296,N_7208);
nand U8896 (N_8896,N_7610,N_7787);
or U8897 (N_8897,N_7704,N_6004);
nand U8898 (N_8898,N_6603,N_7464);
and U8899 (N_8899,N_6765,N_6407);
nand U8900 (N_8900,N_7394,N_7304);
or U8901 (N_8901,N_7026,N_6072);
nand U8902 (N_8902,N_6351,N_6201);
or U8903 (N_8903,N_6026,N_6934);
nor U8904 (N_8904,N_6006,N_6176);
and U8905 (N_8905,N_6725,N_7344);
nor U8906 (N_8906,N_6885,N_6192);
nor U8907 (N_8907,N_6622,N_7762);
nor U8908 (N_8908,N_6495,N_6073);
and U8909 (N_8909,N_7573,N_7777);
nand U8910 (N_8910,N_6618,N_6003);
nand U8911 (N_8911,N_7175,N_6742);
nand U8912 (N_8912,N_6761,N_6980);
or U8913 (N_8913,N_6468,N_7242);
and U8914 (N_8914,N_7695,N_6406);
nand U8915 (N_8915,N_7932,N_6456);
nor U8916 (N_8916,N_6419,N_7668);
and U8917 (N_8917,N_7294,N_7493);
nand U8918 (N_8918,N_7234,N_6912);
or U8919 (N_8919,N_6278,N_7560);
nand U8920 (N_8920,N_6613,N_6645);
or U8921 (N_8921,N_7313,N_7622);
and U8922 (N_8922,N_7137,N_7502);
or U8923 (N_8923,N_7127,N_6370);
nand U8924 (N_8924,N_6301,N_6235);
nand U8925 (N_8925,N_7124,N_7198);
nand U8926 (N_8926,N_7331,N_7499);
or U8927 (N_8927,N_6141,N_6199);
and U8928 (N_8928,N_7497,N_7358);
nand U8929 (N_8929,N_7491,N_7820);
and U8930 (N_8930,N_6440,N_7350);
nand U8931 (N_8931,N_7276,N_7798);
and U8932 (N_8932,N_7037,N_7735);
and U8933 (N_8933,N_6628,N_7631);
or U8934 (N_8934,N_6489,N_7172);
nand U8935 (N_8935,N_7244,N_6524);
or U8936 (N_8936,N_7439,N_7036);
or U8937 (N_8937,N_6476,N_7588);
nor U8938 (N_8938,N_7742,N_7308);
nor U8939 (N_8939,N_6512,N_6038);
xnor U8940 (N_8940,N_6065,N_7141);
nor U8941 (N_8941,N_6159,N_7298);
and U8942 (N_8942,N_7918,N_7129);
nor U8943 (N_8943,N_6300,N_6302);
nand U8944 (N_8944,N_7233,N_6266);
or U8945 (N_8945,N_7606,N_7646);
or U8946 (N_8946,N_6707,N_7835);
nand U8947 (N_8947,N_7536,N_6989);
or U8948 (N_8948,N_7406,N_6632);
or U8949 (N_8949,N_6962,N_6903);
nor U8950 (N_8950,N_6357,N_6763);
or U8951 (N_8951,N_6754,N_7782);
nor U8952 (N_8952,N_6768,N_7707);
or U8953 (N_8953,N_6379,N_7170);
or U8954 (N_8954,N_7593,N_7484);
and U8955 (N_8955,N_7750,N_7149);
and U8956 (N_8956,N_7375,N_7544);
and U8957 (N_8957,N_6402,N_6657);
or U8958 (N_8958,N_6747,N_7600);
or U8959 (N_8959,N_7048,N_7953);
nor U8960 (N_8960,N_6602,N_6310);
nor U8961 (N_8961,N_6497,N_6045);
and U8962 (N_8962,N_6185,N_6647);
xor U8963 (N_8963,N_7492,N_7728);
nand U8964 (N_8964,N_6651,N_6728);
nor U8965 (N_8965,N_6101,N_6160);
or U8966 (N_8966,N_7423,N_7261);
nand U8967 (N_8967,N_7083,N_6872);
and U8968 (N_8968,N_7555,N_7525);
and U8969 (N_8969,N_6825,N_6076);
nand U8970 (N_8970,N_7990,N_6043);
nor U8971 (N_8971,N_7150,N_7014);
nor U8972 (N_8972,N_6202,N_7922);
or U8973 (N_8973,N_7043,N_6970);
nand U8974 (N_8974,N_7299,N_7287);
nor U8975 (N_8975,N_7778,N_6203);
nor U8976 (N_8976,N_7255,N_7768);
and U8977 (N_8977,N_7701,N_7935);
and U8978 (N_8978,N_6973,N_7938);
and U8979 (N_8979,N_6865,N_6244);
nor U8980 (N_8980,N_6866,N_6837);
or U8981 (N_8981,N_7017,N_6680);
or U8982 (N_8982,N_6253,N_6455);
and U8983 (N_8983,N_7987,N_6418);
nor U8984 (N_8984,N_7920,N_6574);
nor U8985 (N_8985,N_7030,N_7154);
or U8986 (N_8986,N_6016,N_6944);
or U8987 (N_8987,N_6034,N_6579);
or U8988 (N_8988,N_6032,N_6358);
nand U8989 (N_8989,N_6589,N_7664);
and U8990 (N_8990,N_7563,N_7159);
nor U8991 (N_8991,N_6215,N_7207);
and U8992 (N_8992,N_7733,N_6046);
nand U8993 (N_8993,N_6732,N_7878);
or U8994 (N_8994,N_7455,N_6950);
or U8995 (N_8995,N_6385,N_7202);
and U8996 (N_8996,N_6071,N_7302);
nor U8997 (N_8997,N_7225,N_6123);
or U8998 (N_8998,N_7013,N_6672);
nand U8999 (N_8999,N_6217,N_7467);
and U9000 (N_9000,N_6151,N_6543);
nand U9001 (N_9001,N_6499,N_7893);
nor U9002 (N_9002,N_6075,N_6475);
or U9003 (N_9003,N_7999,N_7823);
nor U9004 (N_9004,N_7091,N_6159);
or U9005 (N_9005,N_7356,N_6388);
nand U9006 (N_9006,N_7553,N_6767);
or U9007 (N_9007,N_6320,N_7142);
nand U9008 (N_9008,N_6136,N_7649);
nand U9009 (N_9009,N_6805,N_7352);
and U9010 (N_9010,N_6495,N_6687);
nor U9011 (N_9011,N_7592,N_7035);
nor U9012 (N_9012,N_7377,N_6961);
or U9013 (N_9013,N_6609,N_6358);
nand U9014 (N_9014,N_7133,N_6800);
nor U9015 (N_9015,N_7035,N_7728);
and U9016 (N_9016,N_7256,N_7558);
and U9017 (N_9017,N_6780,N_6638);
and U9018 (N_9018,N_6036,N_7264);
and U9019 (N_9019,N_6946,N_7846);
and U9020 (N_9020,N_7212,N_7298);
nand U9021 (N_9021,N_7868,N_7074);
nand U9022 (N_9022,N_7724,N_7021);
nand U9023 (N_9023,N_7803,N_7686);
nor U9024 (N_9024,N_6146,N_6690);
and U9025 (N_9025,N_6132,N_6756);
nor U9026 (N_9026,N_7585,N_7944);
nand U9027 (N_9027,N_7467,N_6609);
and U9028 (N_9028,N_7500,N_6586);
nand U9029 (N_9029,N_7332,N_6426);
nand U9030 (N_9030,N_7503,N_7590);
and U9031 (N_9031,N_6376,N_7109);
nand U9032 (N_9032,N_7924,N_7250);
or U9033 (N_9033,N_6931,N_7479);
and U9034 (N_9034,N_7961,N_7201);
nor U9035 (N_9035,N_7515,N_7106);
nand U9036 (N_9036,N_6290,N_7537);
or U9037 (N_9037,N_7085,N_6224);
nand U9038 (N_9038,N_7799,N_7627);
nor U9039 (N_9039,N_6795,N_6983);
nand U9040 (N_9040,N_6755,N_6610);
or U9041 (N_9041,N_6888,N_7201);
or U9042 (N_9042,N_7039,N_7057);
or U9043 (N_9043,N_7610,N_6196);
nor U9044 (N_9044,N_7490,N_6030);
nor U9045 (N_9045,N_6709,N_6076);
or U9046 (N_9046,N_7393,N_7837);
nor U9047 (N_9047,N_6415,N_7393);
or U9048 (N_9048,N_7312,N_6181);
nor U9049 (N_9049,N_7789,N_7579);
and U9050 (N_9050,N_7036,N_7086);
nand U9051 (N_9051,N_6914,N_6076);
nor U9052 (N_9052,N_7975,N_6312);
nand U9053 (N_9053,N_6926,N_7609);
nand U9054 (N_9054,N_6872,N_6502);
nand U9055 (N_9055,N_6356,N_6475);
or U9056 (N_9056,N_6498,N_6708);
nor U9057 (N_9057,N_7143,N_6884);
nand U9058 (N_9058,N_7807,N_6836);
nand U9059 (N_9059,N_7696,N_7964);
nor U9060 (N_9060,N_7552,N_6899);
or U9061 (N_9061,N_7991,N_7384);
nand U9062 (N_9062,N_6405,N_6338);
or U9063 (N_9063,N_6024,N_7742);
or U9064 (N_9064,N_6922,N_7294);
and U9065 (N_9065,N_6862,N_7482);
nand U9066 (N_9066,N_6666,N_7528);
nor U9067 (N_9067,N_7674,N_6616);
or U9068 (N_9068,N_7908,N_7656);
or U9069 (N_9069,N_6537,N_7582);
nor U9070 (N_9070,N_7402,N_6755);
and U9071 (N_9071,N_6367,N_7845);
or U9072 (N_9072,N_6223,N_6705);
nor U9073 (N_9073,N_7157,N_6943);
nor U9074 (N_9074,N_6470,N_7754);
or U9075 (N_9075,N_7239,N_7682);
and U9076 (N_9076,N_6972,N_6416);
nor U9077 (N_9077,N_6595,N_6059);
nor U9078 (N_9078,N_7458,N_6712);
and U9079 (N_9079,N_6022,N_6227);
or U9080 (N_9080,N_6329,N_6266);
nor U9081 (N_9081,N_6008,N_7905);
nand U9082 (N_9082,N_6227,N_6970);
and U9083 (N_9083,N_7011,N_6650);
nand U9084 (N_9084,N_6026,N_7766);
nand U9085 (N_9085,N_6715,N_7126);
nor U9086 (N_9086,N_7491,N_7637);
nor U9087 (N_9087,N_6315,N_7256);
nor U9088 (N_9088,N_7087,N_7529);
nand U9089 (N_9089,N_7592,N_6525);
nor U9090 (N_9090,N_7610,N_6368);
and U9091 (N_9091,N_7782,N_6127);
nor U9092 (N_9092,N_6913,N_6355);
nand U9093 (N_9093,N_7000,N_6456);
and U9094 (N_9094,N_7386,N_7697);
nor U9095 (N_9095,N_7429,N_7801);
and U9096 (N_9096,N_7005,N_6007);
nor U9097 (N_9097,N_7941,N_7105);
nand U9098 (N_9098,N_7513,N_7094);
and U9099 (N_9099,N_7478,N_7616);
nand U9100 (N_9100,N_6562,N_6484);
and U9101 (N_9101,N_7200,N_7032);
nand U9102 (N_9102,N_7528,N_7400);
or U9103 (N_9103,N_6800,N_6159);
nor U9104 (N_9104,N_6971,N_6667);
or U9105 (N_9105,N_6942,N_7505);
or U9106 (N_9106,N_6223,N_7534);
and U9107 (N_9107,N_6653,N_7284);
nand U9108 (N_9108,N_6026,N_7078);
and U9109 (N_9109,N_6558,N_7229);
nor U9110 (N_9110,N_7815,N_6853);
nor U9111 (N_9111,N_7682,N_7313);
nand U9112 (N_9112,N_7322,N_6094);
nand U9113 (N_9113,N_6178,N_7848);
and U9114 (N_9114,N_7005,N_7594);
nor U9115 (N_9115,N_6972,N_7179);
nor U9116 (N_9116,N_7969,N_6121);
or U9117 (N_9117,N_7647,N_7155);
or U9118 (N_9118,N_7710,N_7869);
nand U9119 (N_9119,N_6486,N_6264);
and U9120 (N_9120,N_7777,N_6394);
and U9121 (N_9121,N_7185,N_7158);
nand U9122 (N_9122,N_6807,N_6177);
and U9123 (N_9123,N_7636,N_7712);
and U9124 (N_9124,N_6982,N_7826);
or U9125 (N_9125,N_6389,N_7830);
nor U9126 (N_9126,N_7906,N_7835);
nand U9127 (N_9127,N_6509,N_6868);
and U9128 (N_9128,N_6449,N_6377);
and U9129 (N_9129,N_7100,N_6645);
nor U9130 (N_9130,N_7575,N_6222);
nor U9131 (N_9131,N_7811,N_7081);
nand U9132 (N_9132,N_6274,N_7017);
nor U9133 (N_9133,N_7029,N_7485);
or U9134 (N_9134,N_6378,N_6472);
and U9135 (N_9135,N_7157,N_6492);
and U9136 (N_9136,N_7468,N_7219);
or U9137 (N_9137,N_7208,N_7024);
nand U9138 (N_9138,N_7852,N_6671);
nand U9139 (N_9139,N_7255,N_6097);
or U9140 (N_9140,N_6377,N_6386);
and U9141 (N_9141,N_6581,N_7033);
or U9142 (N_9142,N_7174,N_7022);
and U9143 (N_9143,N_6316,N_7217);
nand U9144 (N_9144,N_6700,N_6842);
nand U9145 (N_9145,N_7248,N_6265);
nor U9146 (N_9146,N_6643,N_7568);
nand U9147 (N_9147,N_6960,N_6061);
nand U9148 (N_9148,N_6306,N_6364);
nand U9149 (N_9149,N_6435,N_7156);
nand U9150 (N_9150,N_7439,N_6676);
and U9151 (N_9151,N_7147,N_6750);
nor U9152 (N_9152,N_6704,N_7129);
nor U9153 (N_9153,N_7860,N_7672);
and U9154 (N_9154,N_7181,N_6909);
xor U9155 (N_9155,N_6187,N_6405);
and U9156 (N_9156,N_7404,N_6459);
or U9157 (N_9157,N_6316,N_7980);
nand U9158 (N_9158,N_6145,N_6321);
and U9159 (N_9159,N_6679,N_7011);
and U9160 (N_9160,N_7346,N_6694);
nand U9161 (N_9161,N_6125,N_7431);
or U9162 (N_9162,N_6149,N_7139);
or U9163 (N_9163,N_7675,N_7811);
nand U9164 (N_9164,N_6910,N_7250);
or U9165 (N_9165,N_6197,N_7660);
or U9166 (N_9166,N_6733,N_6549);
or U9167 (N_9167,N_6296,N_7352);
xor U9168 (N_9168,N_7878,N_7043);
nand U9169 (N_9169,N_7285,N_7314);
xnor U9170 (N_9170,N_7561,N_7534);
nor U9171 (N_9171,N_6373,N_6016);
and U9172 (N_9172,N_6498,N_7851);
nand U9173 (N_9173,N_6655,N_7644);
nand U9174 (N_9174,N_7326,N_6001);
nor U9175 (N_9175,N_6616,N_7699);
nor U9176 (N_9176,N_6208,N_7192);
nand U9177 (N_9177,N_6403,N_6968);
or U9178 (N_9178,N_7157,N_6018);
nor U9179 (N_9179,N_6516,N_7014);
nand U9180 (N_9180,N_6239,N_6763);
nor U9181 (N_9181,N_6814,N_6098);
nand U9182 (N_9182,N_6152,N_6917);
or U9183 (N_9183,N_7031,N_7066);
or U9184 (N_9184,N_7588,N_7341);
or U9185 (N_9185,N_6290,N_7504);
nor U9186 (N_9186,N_6506,N_7791);
and U9187 (N_9187,N_6253,N_7938);
nor U9188 (N_9188,N_6650,N_7008);
and U9189 (N_9189,N_7716,N_6906);
nor U9190 (N_9190,N_6276,N_7990);
nand U9191 (N_9191,N_6853,N_6146);
nand U9192 (N_9192,N_6450,N_7584);
and U9193 (N_9193,N_6129,N_6310);
or U9194 (N_9194,N_6409,N_6219);
xor U9195 (N_9195,N_7314,N_6594);
or U9196 (N_9196,N_7362,N_7829);
or U9197 (N_9197,N_6206,N_6485);
and U9198 (N_9198,N_6409,N_7983);
and U9199 (N_9199,N_6581,N_6913);
xor U9200 (N_9200,N_7167,N_6613);
nand U9201 (N_9201,N_6954,N_6462);
or U9202 (N_9202,N_7256,N_6866);
nor U9203 (N_9203,N_7917,N_6571);
or U9204 (N_9204,N_6780,N_7887);
nand U9205 (N_9205,N_6142,N_6812);
and U9206 (N_9206,N_7155,N_6254);
and U9207 (N_9207,N_7070,N_6400);
or U9208 (N_9208,N_7467,N_6954);
or U9209 (N_9209,N_6998,N_7595);
nor U9210 (N_9210,N_6833,N_6032);
nand U9211 (N_9211,N_7447,N_7620);
nor U9212 (N_9212,N_6654,N_7662);
or U9213 (N_9213,N_7579,N_7843);
and U9214 (N_9214,N_6934,N_6896);
nand U9215 (N_9215,N_7187,N_7131);
nor U9216 (N_9216,N_6988,N_6841);
nand U9217 (N_9217,N_6265,N_6139);
or U9218 (N_9218,N_7467,N_7676);
and U9219 (N_9219,N_7037,N_6890);
and U9220 (N_9220,N_7756,N_6418);
or U9221 (N_9221,N_7751,N_7722);
xnor U9222 (N_9222,N_6350,N_6118);
nand U9223 (N_9223,N_6630,N_6938);
nor U9224 (N_9224,N_6531,N_6423);
or U9225 (N_9225,N_6308,N_6665);
nor U9226 (N_9226,N_7118,N_7676);
or U9227 (N_9227,N_6763,N_6378);
nor U9228 (N_9228,N_6551,N_6633);
and U9229 (N_9229,N_6992,N_7969);
nand U9230 (N_9230,N_6850,N_7138);
or U9231 (N_9231,N_6765,N_7406);
nand U9232 (N_9232,N_6158,N_6829);
nor U9233 (N_9233,N_6926,N_6718);
nor U9234 (N_9234,N_7191,N_7235);
and U9235 (N_9235,N_6314,N_7341);
nor U9236 (N_9236,N_6326,N_7786);
and U9237 (N_9237,N_7160,N_7970);
and U9238 (N_9238,N_7614,N_7791);
and U9239 (N_9239,N_7432,N_7732);
and U9240 (N_9240,N_6163,N_6580);
nor U9241 (N_9241,N_6113,N_6142);
and U9242 (N_9242,N_7209,N_7229);
nand U9243 (N_9243,N_7024,N_6329);
nand U9244 (N_9244,N_6117,N_6297);
nand U9245 (N_9245,N_7160,N_7619);
and U9246 (N_9246,N_7811,N_7369);
nor U9247 (N_9247,N_6273,N_6908);
nand U9248 (N_9248,N_6564,N_7035);
nor U9249 (N_9249,N_6282,N_6648);
nor U9250 (N_9250,N_6588,N_6755);
nand U9251 (N_9251,N_7229,N_6811);
and U9252 (N_9252,N_6977,N_7307);
nor U9253 (N_9253,N_7432,N_6548);
or U9254 (N_9254,N_6364,N_7953);
and U9255 (N_9255,N_7346,N_7164);
nand U9256 (N_9256,N_6595,N_6739);
nor U9257 (N_9257,N_6007,N_6829);
and U9258 (N_9258,N_6292,N_6833);
nor U9259 (N_9259,N_6087,N_6411);
nor U9260 (N_9260,N_6038,N_6228);
nor U9261 (N_9261,N_7536,N_6574);
and U9262 (N_9262,N_7749,N_6770);
and U9263 (N_9263,N_7381,N_7095);
nor U9264 (N_9264,N_6930,N_6183);
or U9265 (N_9265,N_7493,N_6175);
nor U9266 (N_9266,N_6875,N_7843);
or U9267 (N_9267,N_6886,N_6538);
and U9268 (N_9268,N_6050,N_6580);
or U9269 (N_9269,N_7049,N_6986);
nor U9270 (N_9270,N_7449,N_6875);
nor U9271 (N_9271,N_6852,N_6974);
or U9272 (N_9272,N_7260,N_6891);
nor U9273 (N_9273,N_7358,N_7633);
and U9274 (N_9274,N_7803,N_7867);
nand U9275 (N_9275,N_7850,N_7531);
nand U9276 (N_9276,N_7570,N_7006);
nand U9277 (N_9277,N_6062,N_7599);
nor U9278 (N_9278,N_6123,N_7298);
nor U9279 (N_9279,N_6436,N_7895);
nor U9280 (N_9280,N_7084,N_7797);
nand U9281 (N_9281,N_7945,N_7642);
or U9282 (N_9282,N_7494,N_6068);
nor U9283 (N_9283,N_6985,N_7683);
nand U9284 (N_9284,N_7005,N_7657);
and U9285 (N_9285,N_6186,N_6697);
nor U9286 (N_9286,N_7493,N_6414);
nor U9287 (N_9287,N_6505,N_6341);
nand U9288 (N_9288,N_6156,N_6125);
nor U9289 (N_9289,N_7958,N_6941);
or U9290 (N_9290,N_6055,N_6670);
nand U9291 (N_9291,N_6992,N_6462);
or U9292 (N_9292,N_7188,N_7754);
nor U9293 (N_9293,N_6985,N_6903);
nand U9294 (N_9294,N_6355,N_7850);
or U9295 (N_9295,N_7022,N_7613);
and U9296 (N_9296,N_6100,N_7601);
and U9297 (N_9297,N_7129,N_6816);
or U9298 (N_9298,N_6970,N_6441);
or U9299 (N_9299,N_6893,N_6002);
nor U9300 (N_9300,N_6981,N_6141);
xor U9301 (N_9301,N_7681,N_7731);
or U9302 (N_9302,N_7831,N_6591);
and U9303 (N_9303,N_7420,N_7570);
and U9304 (N_9304,N_7379,N_7466);
nand U9305 (N_9305,N_7611,N_6028);
or U9306 (N_9306,N_7543,N_6272);
or U9307 (N_9307,N_6524,N_7177);
or U9308 (N_9308,N_6184,N_7629);
nor U9309 (N_9309,N_6161,N_6969);
or U9310 (N_9310,N_7152,N_7836);
nor U9311 (N_9311,N_7909,N_6559);
xnor U9312 (N_9312,N_7729,N_6904);
and U9313 (N_9313,N_7280,N_6300);
xnor U9314 (N_9314,N_6238,N_7943);
nor U9315 (N_9315,N_6907,N_7579);
nor U9316 (N_9316,N_6003,N_6801);
and U9317 (N_9317,N_6167,N_6664);
or U9318 (N_9318,N_6515,N_6562);
nor U9319 (N_9319,N_6943,N_7446);
nand U9320 (N_9320,N_6903,N_7356);
nand U9321 (N_9321,N_6735,N_6828);
nor U9322 (N_9322,N_7583,N_7261);
and U9323 (N_9323,N_7215,N_6132);
and U9324 (N_9324,N_6880,N_7720);
nor U9325 (N_9325,N_7011,N_6046);
or U9326 (N_9326,N_6501,N_7672);
and U9327 (N_9327,N_6046,N_7665);
nor U9328 (N_9328,N_6815,N_7394);
nor U9329 (N_9329,N_6816,N_7883);
nor U9330 (N_9330,N_6704,N_6074);
nor U9331 (N_9331,N_6638,N_6801);
nand U9332 (N_9332,N_7087,N_6452);
or U9333 (N_9333,N_7381,N_6610);
nor U9334 (N_9334,N_7563,N_7674);
or U9335 (N_9335,N_7777,N_6914);
or U9336 (N_9336,N_6252,N_6844);
or U9337 (N_9337,N_7325,N_6215);
or U9338 (N_9338,N_7974,N_7447);
xnor U9339 (N_9339,N_6065,N_6502);
and U9340 (N_9340,N_7234,N_6097);
and U9341 (N_9341,N_7766,N_6011);
or U9342 (N_9342,N_7651,N_6297);
nor U9343 (N_9343,N_7424,N_7742);
nor U9344 (N_9344,N_7609,N_6620);
or U9345 (N_9345,N_7204,N_6919);
nand U9346 (N_9346,N_7834,N_7390);
and U9347 (N_9347,N_6761,N_6301);
nor U9348 (N_9348,N_7805,N_6478);
nand U9349 (N_9349,N_6090,N_7090);
or U9350 (N_9350,N_7217,N_7027);
nand U9351 (N_9351,N_7799,N_6499);
nand U9352 (N_9352,N_7926,N_6817);
nor U9353 (N_9353,N_7489,N_7568);
nand U9354 (N_9354,N_6595,N_7720);
nand U9355 (N_9355,N_6027,N_7685);
nand U9356 (N_9356,N_6223,N_6243);
or U9357 (N_9357,N_7997,N_6543);
or U9358 (N_9358,N_6227,N_6873);
and U9359 (N_9359,N_6747,N_7399);
or U9360 (N_9360,N_6120,N_7714);
or U9361 (N_9361,N_6167,N_7729);
nor U9362 (N_9362,N_6766,N_7334);
and U9363 (N_9363,N_7578,N_6629);
and U9364 (N_9364,N_7747,N_6410);
nand U9365 (N_9365,N_7979,N_6810);
nand U9366 (N_9366,N_6882,N_7206);
nand U9367 (N_9367,N_6526,N_7871);
or U9368 (N_9368,N_6010,N_6396);
or U9369 (N_9369,N_6587,N_6609);
or U9370 (N_9370,N_7246,N_6162);
xor U9371 (N_9371,N_6701,N_7686);
or U9372 (N_9372,N_6072,N_7835);
and U9373 (N_9373,N_6723,N_6295);
nand U9374 (N_9374,N_6007,N_6056);
or U9375 (N_9375,N_6868,N_7062);
and U9376 (N_9376,N_6755,N_7174);
and U9377 (N_9377,N_6376,N_6106);
and U9378 (N_9378,N_7946,N_7936);
or U9379 (N_9379,N_6149,N_6794);
nor U9380 (N_9380,N_6996,N_6779);
and U9381 (N_9381,N_7317,N_7771);
and U9382 (N_9382,N_6419,N_7231);
and U9383 (N_9383,N_7629,N_6821);
xor U9384 (N_9384,N_6782,N_6317);
or U9385 (N_9385,N_7216,N_7309);
or U9386 (N_9386,N_7067,N_7700);
or U9387 (N_9387,N_7182,N_7432);
or U9388 (N_9388,N_6101,N_6768);
and U9389 (N_9389,N_6214,N_6540);
or U9390 (N_9390,N_7427,N_6113);
or U9391 (N_9391,N_7656,N_7911);
and U9392 (N_9392,N_7874,N_7152);
and U9393 (N_9393,N_7068,N_6421);
nand U9394 (N_9394,N_6670,N_7809);
nand U9395 (N_9395,N_6913,N_6386);
and U9396 (N_9396,N_6029,N_6846);
and U9397 (N_9397,N_6413,N_6092);
nor U9398 (N_9398,N_7261,N_7794);
or U9399 (N_9399,N_7548,N_6363);
and U9400 (N_9400,N_6062,N_6224);
or U9401 (N_9401,N_6414,N_6031);
nand U9402 (N_9402,N_7849,N_7218);
and U9403 (N_9403,N_6298,N_7929);
nor U9404 (N_9404,N_7460,N_7693);
nor U9405 (N_9405,N_7181,N_7506);
or U9406 (N_9406,N_6773,N_6921);
and U9407 (N_9407,N_6142,N_6403);
and U9408 (N_9408,N_6751,N_6459);
and U9409 (N_9409,N_7468,N_6866);
xnor U9410 (N_9410,N_7854,N_7440);
nand U9411 (N_9411,N_7015,N_6727);
and U9412 (N_9412,N_7147,N_6689);
and U9413 (N_9413,N_6341,N_7584);
nand U9414 (N_9414,N_7289,N_7170);
nor U9415 (N_9415,N_7796,N_6501);
or U9416 (N_9416,N_6799,N_7386);
nand U9417 (N_9417,N_7970,N_7908);
or U9418 (N_9418,N_6603,N_6121);
or U9419 (N_9419,N_6512,N_7939);
nor U9420 (N_9420,N_7835,N_7403);
nor U9421 (N_9421,N_6713,N_7819);
and U9422 (N_9422,N_6958,N_7542);
or U9423 (N_9423,N_7079,N_7346);
nor U9424 (N_9424,N_6236,N_6171);
or U9425 (N_9425,N_6648,N_6640);
nor U9426 (N_9426,N_7841,N_7744);
and U9427 (N_9427,N_6205,N_6781);
and U9428 (N_9428,N_6657,N_7733);
nor U9429 (N_9429,N_7346,N_6611);
nor U9430 (N_9430,N_7037,N_6927);
nand U9431 (N_9431,N_6876,N_7484);
or U9432 (N_9432,N_7861,N_7369);
nor U9433 (N_9433,N_6817,N_7190);
nor U9434 (N_9434,N_7982,N_6663);
and U9435 (N_9435,N_7538,N_7361);
or U9436 (N_9436,N_7297,N_7223);
nor U9437 (N_9437,N_7583,N_7830);
and U9438 (N_9438,N_6410,N_6207);
and U9439 (N_9439,N_6883,N_6869);
nor U9440 (N_9440,N_7114,N_6678);
or U9441 (N_9441,N_6119,N_7467);
nor U9442 (N_9442,N_7434,N_7123);
and U9443 (N_9443,N_7745,N_7832);
or U9444 (N_9444,N_7851,N_7534);
or U9445 (N_9445,N_6153,N_7956);
nor U9446 (N_9446,N_6093,N_7211);
nand U9447 (N_9447,N_6866,N_7650);
nor U9448 (N_9448,N_6514,N_7730);
nand U9449 (N_9449,N_7943,N_6740);
or U9450 (N_9450,N_7212,N_6123);
or U9451 (N_9451,N_7523,N_7197);
or U9452 (N_9452,N_6078,N_7846);
or U9453 (N_9453,N_6414,N_6302);
nand U9454 (N_9454,N_6045,N_7424);
nor U9455 (N_9455,N_7882,N_6815);
nor U9456 (N_9456,N_6510,N_6401);
and U9457 (N_9457,N_7182,N_6562);
nor U9458 (N_9458,N_7738,N_7377);
nand U9459 (N_9459,N_6633,N_7385);
nand U9460 (N_9460,N_6717,N_7207);
nor U9461 (N_9461,N_6731,N_7874);
nor U9462 (N_9462,N_6907,N_7895);
nor U9463 (N_9463,N_6669,N_7288);
or U9464 (N_9464,N_7610,N_6403);
and U9465 (N_9465,N_6451,N_7335);
nand U9466 (N_9466,N_7606,N_7594);
nor U9467 (N_9467,N_6849,N_6931);
or U9468 (N_9468,N_7739,N_6348);
and U9469 (N_9469,N_6967,N_6508);
or U9470 (N_9470,N_6002,N_6384);
nor U9471 (N_9471,N_6357,N_7037);
or U9472 (N_9472,N_7989,N_7750);
nor U9473 (N_9473,N_6561,N_6012);
and U9474 (N_9474,N_7832,N_7916);
nand U9475 (N_9475,N_6213,N_7112);
and U9476 (N_9476,N_6104,N_7190);
or U9477 (N_9477,N_7020,N_6007);
or U9478 (N_9478,N_6813,N_7967);
and U9479 (N_9479,N_6991,N_7672);
nor U9480 (N_9480,N_6871,N_6218);
nor U9481 (N_9481,N_7353,N_7831);
and U9482 (N_9482,N_7739,N_6419);
nand U9483 (N_9483,N_6283,N_6282);
or U9484 (N_9484,N_6054,N_6170);
nor U9485 (N_9485,N_6117,N_6788);
nor U9486 (N_9486,N_7978,N_6312);
nor U9487 (N_9487,N_6177,N_6227);
and U9488 (N_9488,N_7941,N_6486);
nor U9489 (N_9489,N_6744,N_6012);
and U9490 (N_9490,N_7764,N_7399);
nand U9491 (N_9491,N_7170,N_6517);
nand U9492 (N_9492,N_7714,N_6056);
or U9493 (N_9493,N_6227,N_7863);
nor U9494 (N_9494,N_6238,N_6325);
or U9495 (N_9495,N_7841,N_7683);
nor U9496 (N_9496,N_7481,N_6445);
nor U9497 (N_9497,N_6274,N_7332);
nor U9498 (N_9498,N_6349,N_6270);
nand U9499 (N_9499,N_7458,N_6403);
nor U9500 (N_9500,N_7077,N_7623);
or U9501 (N_9501,N_6042,N_6897);
or U9502 (N_9502,N_7214,N_7058);
nor U9503 (N_9503,N_6142,N_6081);
or U9504 (N_9504,N_6698,N_6726);
or U9505 (N_9505,N_7672,N_6169);
or U9506 (N_9506,N_7298,N_7674);
nor U9507 (N_9507,N_6817,N_6019);
nand U9508 (N_9508,N_7282,N_7832);
or U9509 (N_9509,N_7436,N_6204);
nor U9510 (N_9510,N_7797,N_7663);
nand U9511 (N_9511,N_6035,N_6994);
and U9512 (N_9512,N_7158,N_6975);
nor U9513 (N_9513,N_7727,N_6498);
and U9514 (N_9514,N_7787,N_7737);
nor U9515 (N_9515,N_6142,N_7850);
and U9516 (N_9516,N_7502,N_6767);
xnor U9517 (N_9517,N_7505,N_6429);
or U9518 (N_9518,N_6615,N_6316);
nand U9519 (N_9519,N_7399,N_7408);
or U9520 (N_9520,N_7321,N_7562);
and U9521 (N_9521,N_6767,N_7555);
nand U9522 (N_9522,N_6065,N_7757);
or U9523 (N_9523,N_6865,N_6579);
or U9524 (N_9524,N_6580,N_7938);
nor U9525 (N_9525,N_6843,N_6010);
or U9526 (N_9526,N_7878,N_7292);
nand U9527 (N_9527,N_7761,N_7138);
and U9528 (N_9528,N_6677,N_6283);
nor U9529 (N_9529,N_6150,N_7549);
and U9530 (N_9530,N_7225,N_6760);
nor U9531 (N_9531,N_6976,N_7760);
nand U9532 (N_9532,N_6156,N_7230);
or U9533 (N_9533,N_6781,N_6068);
nor U9534 (N_9534,N_6773,N_7861);
and U9535 (N_9535,N_7472,N_6842);
or U9536 (N_9536,N_7131,N_7548);
and U9537 (N_9537,N_7632,N_6366);
nor U9538 (N_9538,N_6934,N_7109);
nor U9539 (N_9539,N_6668,N_7410);
and U9540 (N_9540,N_7132,N_7332);
xor U9541 (N_9541,N_6322,N_6420);
and U9542 (N_9542,N_6835,N_6521);
nand U9543 (N_9543,N_7336,N_7668);
nor U9544 (N_9544,N_6920,N_7099);
nor U9545 (N_9545,N_7024,N_7400);
nand U9546 (N_9546,N_6461,N_7980);
nand U9547 (N_9547,N_7277,N_7812);
or U9548 (N_9548,N_6004,N_7164);
or U9549 (N_9549,N_6971,N_6731);
or U9550 (N_9550,N_7624,N_7439);
nor U9551 (N_9551,N_7578,N_7617);
and U9552 (N_9552,N_6922,N_6609);
and U9553 (N_9553,N_6911,N_7566);
and U9554 (N_9554,N_7154,N_6001);
or U9555 (N_9555,N_7466,N_6612);
and U9556 (N_9556,N_6153,N_6362);
or U9557 (N_9557,N_7556,N_6598);
nand U9558 (N_9558,N_7684,N_6629);
xnor U9559 (N_9559,N_6363,N_6610);
nand U9560 (N_9560,N_7912,N_7550);
or U9561 (N_9561,N_7610,N_7530);
xnor U9562 (N_9562,N_7780,N_7841);
and U9563 (N_9563,N_7966,N_6419);
or U9564 (N_9564,N_7324,N_7836);
and U9565 (N_9565,N_7914,N_6935);
or U9566 (N_9566,N_6282,N_6610);
and U9567 (N_9567,N_7218,N_6723);
nor U9568 (N_9568,N_7643,N_6517);
nor U9569 (N_9569,N_6948,N_6606);
nand U9570 (N_9570,N_6355,N_7407);
and U9571 (N_9571,N_7885,N_6348);
nor U9572 (N_9572,N_6794,N_6530);
nand U9573 (N_9573,N_7246,N_6053);
nor U9574 (N_9574,N_6078,N_7417);
and U9575 (N_9575,N_7250,N_7060);
nor U9576 (N_9576,N_7254,N_7003);
nand U9577 (N_9577,N_7764,N_6923);
nor U9578 (N_9578,N_7800,N_6933);
or U9579 (N_9579,N_7219,N_6974);
nand U9580 (N_9580,N_6932,N_6860);
or U9581 (N_9581,N_6681,N_7401);
nor U9582 (N_9582,N_7132,N_6014);
nor U9583 (N_9583,N_6577,N_6735);
or U9584 (N_9584,N_6740,N_6416);
or U9585 (N_9585,N_6131,N_6880);
nand U9586 (N_9586,N_7753,N_7822);
nor U9587 (N_9587,N_7528,N_7604);
nor U9588 (N_9588,N_7629,N_6472);
nand U9589 (N_9589,N_7342,N_6912);
or U9590 (N_9590,N_7261,N_6102);
nand U9591 (N_9591,N_7851,N_6662);
or U9592 (N_9592,N_6487,N_6091);
nor U9593 (N_9593,N_7358,N_6098);
or U9594 (N_9594,N_7706,N_7257);
nand U9595 (N_9595,N_7150,N_7300);
or U9596 (N_9596,N_7812,N_7749);
and U9597 (N_9597,N_6504,N_7340);
or U9598 (N_9598,N_7967,N_6160);
nand U9599 (N_9599,N_6671,N_6598);
nor U9600 (N_9600,N_6489,N_6720);
and U9601 (N_9601,N_6334,N_7706);
nand U9602 (N_9602,N_6493,N_6727);
and U9603 (N_9603,N_7884,N_7636);
or U9604 (N_9604,N_6104,N_7281);
or U9605 (N_9605,N_7020,N_7281);
or U9606 (N_9606,N_6601,N_6463);
nand U9607 (N_9607,N_6161,N_7278);
or U9608 (N_9608,N_6099,N_7952);
nand U9609 (N_9609,N_6696,N_6633);
nand U9610 (N_9610,N_6775,N_6439);
nor U9611 (N_9611,N_6666,N_7366);
nand U9612 (N_9612,N_7912,N_7338);
and U9613 (N_9613,N_6196,N_7283);
nand U9614 (N_9614,N_7418,N_6933);
nand U9615 (N_9615,N_6989,N_6087);
or U9616 (N_9616,N_6852,N_6527);
or U9617 (N_9617,N_6837,N_6670);
or U9618 (N_9618,N_7266,N_7323);
and U9619 (N_9619,N_6971,N_7022);
nand U9620 (N_9620,N_7661,N_7367);
nor U9621 (N_9621,N_6883,N_7718);
nand U9622 (N_9622,N_6247,N_6704);
nand U9623 (N_9623,N_6288,N_7641);
nand U9624 (N_9624,N_6638,N_7151);
nand U9625 (N_9625,N_7803,N_6116);
and U9626 (N_9626,N_7521,N_7991);
nor U9627 (N_9627,N_6918,N_7991);
nor U9628 (N_9628,N_7696,N_7993);
or U9629 (N_9629,N_7703,N_7756);
and U9630 (N_9630,N_7403,N_6144);
and U9631 (N_9631,N_7106,N_7731);
nand U9632 (N_9632,N_6369,N_6330);
nand U9633 (N_9633,N_6187,N_6241);
nor U9634 (N_9634,N_6576,N_7818);
nand U9635 (N_9635,N_6918,N_6395);
and U9636 (N_9636,N_7446,N_7103);
nand U9637 (N_9637,N_6350,N_7224);
nand U9638 (N_9638,N_6062,N_6591);
nand U9639 (N_9639,N_7458,N_6633);
or U9640 (N_9640,N_7044,N_6301);
or U9641 (N_9641,N_7950,N_7185);
nand U9642 (N_9642,N_6691,N_7301);
and U9643 (N_9643,N_6322,N_7221);
nor U9644 (N_9644,N_7913,N_7486);
nand U9645 (N_9645,N_7153,N_7816);
or U9646 (N_9646,N_7027,N_7507);
or U9647 (N_9647,N_7594,N_7766);
nand U9648 (N_9648,N_7812,N_7445);
or U9649 (N_9649,N_7399,N_7137);
nand U9650 (N_9650,N_7330,N_7318);
nand U9651 (N_9651,N_7689,N_6806);
xor U9652 (N_9652,N_6162,N_7003);
and U9653 (N_9653,N_7171,N_7871);
and U9654 (N_9654,N_7658,N_7131);
nand U9655 (N_9655,N_6767,N_6472);
nand U9656 (N_9656,N_7721,N_6439);
or U9657 (N_9657,N_7605,N_6753);
nand U9658 (N_9658,N_6957,N_7981);
nor U9659 (N_9659,N_6064,N_7551);
nor U9660 (N_9660,N_7454,N_6556);
nor U9661 (N_9661,N_6261,N_6110);
nor U9662 (N_9662,N_7029,N_6846);
nand U9663 (N_9663,N_6640,N_6613);
nand U9664 (N_9664,N_6520,N_7780);
and U9665 (N_9665,N_7018,N_6697);
nor U9666 (N_9666,N_6512,N_6067);
or U9667 (N_9667,N_6725,N_6637);
nor U9668 (N_9668,N_6335,N_7911);
or U9669 (N_9669,N_7710,N_6964);
and U9670 (N_9670,N_7354,N_6221);
or U9671 (N_9671,N_6875,N_6445);
nand U9672 (N_9672,N_7911,N_7517);
nand U9673 (N_9673,N_7331,N_6667);
and U9674 (N_9674,N_6345,N_6298);
and U9675 (N_9675,N_7935,N_6927);
or U9676 (N_9676,N_7602,N_6407);
or U9677 (N_9677,N_7746,N_7496);
or U9678 (N_9678,N_6662,N_6642);
or U9679 (N_9679,N_7160,N_6811);
or U9680 (N_9680,N_6555,N_6708);
nand U9681 (N_9681,N_7686,N_7324);
nor U9682 (N_9682,N_6333,N_7564);
or U9683 (N_9683,N_7527,N_6028);
nand U9684 (N_9684,N_6456,N_6762);
nand U9685 (N_9685,N_7437,N_7780);
nand U9686 (N_9686,N_6464,N_6788);
and U9687 (N_9687,N_7493,N_7823);
or U9688 (N_9688,N_6363,N_6614);
or U9689 (N_9689,N_6363,N_7651);
or U9690 (N_9690,N_7052,N_6743);
nor U9691 (N_9691,N_6594,N_7402);
nor U9692 (N_9692,N_6128,N_6638);
nand U9693 (N_9693,N_7182,N_6617);
or U9694 (N_9694,N_6962,N_6314);
and U9695 (N_9695,N_6792,N_6205);
nand U9696 (N_9696,N_6738,N_7456);
nand U9697 (N_9697,N_7895,N_6011);
or U9698 (N_9698,N_6523,N_6860);
or U9699 (N_9699,N_7399,N_6569);
and U9700 (N_9700,N_6168,N_7936);
or U9701 (N_9701,N_7127,N_7326);
nand U9702 (N_9702,N_7205,N_6683);
nor U9703 (N_9703,N_6984,N_6802);
nor U9704 (N_9704,N_7384,N_6137);
nor U9705 (N_9705,N_7931,N_6959);
and U9706 (N_9706,N_7678,N_7274);
nand U9707 (N_9707,N_6198,N_7061);
and U9708 (N_9708,N_6875,N_6843);
and U9709 (N_9709,N_7131,N_6584);
and U9710 (N_9710,N_6641,N_6262);
and U9711 (N_9711,N_6950,N_6960);
nor U9712 (N_9712,N_7369,N_6544);
and U9713 (N_9713,N_6874,N_7409);
and U9714 (N_9714,N_7323,N_6653);
and U9715 (N_9715,N_7845,N_6262);
and U9716 (N_9716,N_6187,N_7201);
nand U9717 (N_9717,N_7900,N_6953);
and U9718 (N_9718,N_6476,N_6763);
nand U9719 (N_9719,N_6444,N_7029);
xnor U9720 (N_9720,N_7298,N_6082);
or U9721 (N_9721,N_6938,N_6133);
and U9722 (N_9722,N_6101,N_6290);
nor U9723 (N_9723,N_7889,N_6595);
or U9724 (N_9724,N_6297,N_6229);
or U9725 (N_9725,N_6482,N_6967);
nor U9726 (N_9726,N_7891,N_6359);
nor U9727 (N_9727,N_6289,N_6125);
and U9728 (N_9728,N_7010,N_6681);
nand U9729 (N_9729,N_7240,N_6331);
nand U9730 (N_9730,N_7372,N_6084);
nand U9731 (N_9731,N_7421,N_7406);
or U9732 (N_9732,N_7032,N_6154);
nand U9733 (N_9733,N_7573,N_7865);
nor U9734 (N_9734,N_7192,N_6911);
nor U9735 (N_9735,N_7584,N_7471);
and U9736 (N_9736,N_6362,N_7761);
and U9737 (N_9737,N_7179,N_7658);
nor U9738 (N_9738,N_6817,N_7527);
or U9739 (N_9739,N_7097,N_7455);
and U9740 (N_9740,N_6436,N_7707);
nor U9741 (N_9741,N_6292,N_6741);
nor U9742 (N_9742,N_6661,N_6760);
nand U9743 (N_9743,N_7296,N_7131);
xor U9744 (N_9744,N_6459,N_6135);
or U9745 (N_9745,N_7111,N_6330);
and U9746 (N_9746,N_7407,N_7524);
and U9747 (N_9747,N_6314,N_7758);
nand U9748 (N_9748,N_7529,N_6617);
and U9749 (N_9749,N_7679,N_6723);
nor U9750 (N_9750,N_7046,N_7787);
or U9751 (N_9751,N_7319,N_6894);
nor U9752 (N_9752,N_7536,N_7660);
and U9753 (N_9753,N_7214,N_6723);
nand U9754 (N_9754,N_6304,N_6700);
nor U9755 (N_9755,N_6513,N_7764);
nor U9756 (N_9756,N_7723,N_7207);
or U9757 (N_9757,N_7723,N_6593);
or U9758 (N_9758,N_6311,N_6572);
xor U9759 (N_9759,N_6859,N_6668);
nand U9760 (N_9760,N_7744,N_7338);
and U9761 (N_9761,N_7270,N_7360);
and U9762 (N_9762,N_7506,N_7442);
nand U9763 (N_9763,N_7556,N_7964);
nand U9764 (N_9764,N_7404,N_6561);
nand U9765 (N_9765,N_6959,N_7363);
or U9766 (N_9766,N_7064,N_7253);
and U9767 (N_9767,N_6903,N_6987);
nor U9768 (N_9768,N_7077,N_6851);
and U9769 (N_9769,N_6506,N_6316);
nand U9770 (N_9770,N_6613,N_6680);
nor U9771 (N_9771,N_6392,N_6212);
or U9772 (N_9772,N_7706,N_6329);
nor U9773 (N_9773,N_7148,N_6529);
nor U9774 (N_9774,N_7764,N_6164);
and U9775 (N_9775,N_6340,N_6904);
or U9776 (N_9776,N_6178,N_7288);
or U9777 (N_9777,N_6109,N_6021);
and U9778 (N_9778,N_6879,N_7969);
or U9779 (N_9779,N_7033,N_7859);
and U9780 (N_9780,N_6420,N_7962);
nor U9781 (N_9781,N_6813,N_7885);
and U9782 (N_9782,N_7749,N_7212);
or U9783 (N_9783,N_7266,N_6722);
nand U9784 (N_9784,N_7175,N_7197);
nor U9785 (N_9785,N_6307,N_7761);
nor U9786 (N_9786,N_6821,N_6601);
or U9787 (N_9787,N_6670,N_6377);
nand U9788 (N_9788,N_7610,N_6168);
xnor U9789 (N_9789,N_7317,N_7371);
nor U9790 (N_9790,N_7095,N_7338);
nand U9791 (N_9791,N_6415,N_6382);
nor U9792 (N_9792,N_6982,N_7444);
nand U9793 (N_9793,N_6366,N_7902);
and U9794 (N_9794,N_6927,N_7860);
or U9795 (N_9795,N_7805,N_7227);
nor U9796 (N_9796,N_6340,N_6162);
nor U9797 (N_9797,N_6865,N_7163);
nor U9798 (N_9798,N_7965,N_6545);
nor U9799 (N_9799,N_7650,N_6946);
or U9800 (N_9800,N_7654,N_7196);
nor U9801 (N_9801,N_6578,N_6512);
nand U9802 (N_9802,N_6036,N_7637);
or U9803 (N_9803,N_7655,N_6476);
nand U9804 (N_9804,N_6112,N_6120);
or U9805 (N_9805,N_6803,N_7423);
and U9806 (N_9806,N_7503,N_7882);
nand U9807 (N_9807,N_6213,N_7753);
nor U9808 (N_9808,N_6847,N_7961);
nand U9809 (N_9809,N_6985,N_6479);
and U9810 (N_9810,N_6959,N_6722);
nand U9811 (N_9811,N_7738,N_6844);
nand U9812 (N_9812,N_7606,N_7130);
nor U9813 (N_9813,N_6344,N_7343);
nand U9814 (N_9814,N_6963,N_7937);
nor U9815 (N_9815,N_7234,N_6074);
nand U9816 (N_9816,N_7412,N_7674);
nor U9817 (N_9817,N_6743,N_7215);
nand U9818 (N_9818,N_6366,N_7780);
and U9819 (N_9819,N_6108,N_7408);
or U9820 (N_9820,N_7325,N_6542);
and U9821 (N_9821,N_7256,N_7065);
nor U9822 (N_9822,N_7989,N_7341);
nor U9823 (N_9823,N_7900,N_7309);
and U9824 (N_9824,N_6595,N_7508);
and U9825 (N_9825,N_6596,N_6122);
and U9826 (N_9826,N_7224,N_7042);
or U9827 (N_9827,N_6723,N_6939);
or U9828 (N_9828,N_6386,N_6146);
and U9829 (N_9829,N_7896,N_6559);
nor U9830 (N_9830,N_6924,N_6853);
nor U9831 (N_9831,N_6806,N_6433);
or U9832 (N_9832,N_7967,N_6300);
or U9833 (N_9833,N_7353,N_7484);
or U9834 (N_9834,N_6434,N_7476);
nand U9835 (N_9835,N_6244,N_7153);
nand U9836 (N_9836,N_7704,N_6432);
or U9837 (N_9837,N_7996,N_7274);
nor U9838 (N_9838,N_6041,N_7654);
nand U9839 (N_9839,N_6341,N_6031);
nor U9840 (N_9840,N_7238,N_7279);
nor U9841 (N_9841,N_7380,N_6750);
or U9842 (N_9842,N_6285,N_7642);
nor U9843 (N_9843,N_7976,N_6673);
and U9844 (N_9844,N_7600,N_7598);
nor U9845 (N_9845,N_6074,N_6218);
nor U9846 (N_9846,N_7029,N_6776);
xnor U9847 (N_9847,N_7742,N_6659);
and U9848 (N_9848,N_7544,N_6273);
nand U9849 (N_9849,N_6073,N_6338);
nor U9850 (N_9850,N_6434,N_7300);
nor U9851 (N_9851,N_7172,N_6414);
nand U9852 (N_9852,N_7875,N_6703);
nand U9853 (N_9853,N_6519,N_7572);
and U9854 (N_9854,N_7968,N_6870);
or U9855 (N_9855,N_7774,N_7609);
nand U9856 (N_9856,N_6044,N_6437);
or U9857 (N_9857,N_6755,N_7323);
nor U9858 (N_9858,N_7926,N_7328);
nand U9859 (N_9859,N_6417,N_7911);
or U9860 (N_9860,N_7116,N_7784);
or U9861 (N_9861,N_7916,N_6252);
or U9862 (N_9862,N_7344,N_6592);
or U9863 (N_9863,N_6267,N_6101);
nor U9864 (N_9864,N_6166,N_6663);
nor U9865 (N_9865,N_6572,N_7900);
and U9866 (N_9866,N_6512,N_6640);
or U9867 (N_9867,N_7652,N_7664);
nor U9868 (N_9868,N_6867,N_7582);
nand U9869 (N_9869,N_6775,N_6920);
nor U9870 (N_9870,N_6934,N_7863);
nor U9871 (N_9871,N_6261,N_7588);
and U9872 (N_9872,N_6248,N_7925);
or U9873 (N_9873,N_7026,N_6579);
nor U9874 (N_9874,N_7626,N_6110);
nor U9875 (N_9875,N_6809,N_6290);
nand U9876 (N_9876,N_6243,N_7041);
and U9877 (N_9877,N_7310,N_7142);
nor U9878 (N_9878,N_6283,N_7947);
and U9879 (N_9879,N_7046,N_7615);
nand U9880 (N_9880,N_7069,N_6621);
or U9881 (N_9881,N_7142,N_7320);
or U9882 (N_9882,N_7307,N_7250);
and U9883 (N_9883,N_6376,N_7980);
or U9884 (N_9884,N_7664,N_7057);
or U9885 (N_9885,N_7779,N_7189);
nor U9886 (N_9886,N_7089,N_7979);
nand U9887 (N_9887,N_6502,N_7884);
or U9888 (N_9888,N_6442,N_6162);
nor U9889 (N_9889,N_7258,N_7339);
nor U9890 (N_9890,N_6989,N_7657);
and U9891 (N_9891,N_7187,N_7191);
nand U9892 (N_9892,N_7950,N_7033);
or U9893 (N_9893,N_6984,N_6512);
nand U9894 (N_9894,N_7240,N_6485);
nand U9895 (N_9895,N_6841,N_7536);
nor U9896 (N_9896,N_7246,N_7679);
nand U9897 (N_9897,N_6999,N_6640);
nor U9898 (N_9898,N_7387,N_6361);
nor U9899 (N_9899,N_6712,N_7926);
and U9900 (N_9900,N_6705,N_7136);
or U9901 (N_9901,N_6723,N_7336);
and U9902 (N_9902,N_6150,N_6105);
and U9903 (N_9903,N_6622,N_7575);
or U9904 (N_9904,N_7181,N_6589);
and U9905 (N_9905,N_7250,N_6149);
or U9906 (N_9906,N_6003,N_6709);
or U9907 (N_9907,N_6278,N_6046);
or U9908 (N_9908,N_7381,N_6753);
nand U9909 (N_9909,N_6526,N_6386);
or U9910 (N_9910,N_6728,N_7713);
nor U9911 (N_9911,N_6590,N_7930);
and U9912 (N_9912,N_6015,N_7513);
nor U9913 (N_9913,N_6213,N_6157);
or U9914 (N_9914,N_7732,N_7452);
and U9915 (N_9915,N_6385,N_7417);
and U9916 (N_9916,N_7286,N_6091);
or U9917 (N_9917,N_6270,N_7010);
nor U9918 (N_9918,N_7619,N_6194);
nand U9919 (N_9919,N_7497,N_7999);
and U9920 (N_9920,N_6398,N_7513);
and U9921 (N_9921,N_6761,N_6555);
and U9922 (N_9922,N_6602,N_7989);
or U9923 (N_9923,N_6120,N_7085);
nand U9924 (N_9924,N_6246,N_7790);
and U9925 (N_9925,N_7255,N_7853);
and U9926 (N_9926,N_6397,N_7682);
and U9927 (N_9927,N_6276,N_7719);
nand U9928 (N_9928,N_6995,N_7099);
and U9929 (N_9929,N_6384,N_6489);
and U9930 (N_9930,N_7876,N_6199);
nand U9931 (N_9931,N_7061,N_7336);
nand U9932 (N_9932,N_7337,N_7454);
nand U9933 (N_9933,N_6716,N_7095);
or U9934 (N_9934,N_7539,N_7502);
nor U9935 (N_9935,N_6951,N_7484);
nand U9936 (N_9936,N_6100,N_7504);
nor U9937 (N_9937,N_6461,N_7628);
nand U9938 (N_9938,N_7752,N_6308);
or U9939 (N_9939,N_7313,N_6201);
or U9940 (N_9940,N_6490,N_6939);
nor U9941 (N_9941,N_6760,N_7364);
or U9942 (N_9942,N_7166,N_6277);
nor U9943 (N_9943,N_6264,N_6672);
or U9944 (N_9944,N_6817,N_7337);
nand U9945 (N_9945,N_7616,N_7079);
and U9946 (N_9946,N_6070,N_7239);
or U9947 (N_9947,N_6949,N_7322);
and U9948 (N_9948,N_7198,N_7061);
nand U9949 (N_9949,N_7946,N_6479);
nand U9950 (N_9950,N_6868,N_6857);
nor U9951 (N_9951,N_6172,N_7776);
or U9952 (N_9952,N_7562,N_6058);
and U9953 (N_9953,N_7640,N_7599);
nor U9954 (N_9954,N_7332,N_6236);
or U9955 (N_9955,N_7964,N_6257);
or U9956 (N_9956,N_6757,N_7536);
or U9957 (N_9957,N_7038,N_6143);
nor U9958 (N_9958,N_7046,N_6634);
nor U9959 (N_9959,N_7208,N_6375);
and U9960 (N_9960,N_6481,N_7809);
nand U9961 (N_9961,N_7820,N_7750);
nor U9962 (N_9962,N_7604,N_7062);
and U9963 (N_9963,N_7395,N_6183);
nor U9964 (N_9964,N_7170,N_7884);
nor U9965 (N_9965,N_7791,N_6925);
or U9966 (N_9966,N_6170,N_6952);
or U9967 (N_9967,N_6200,N_7516);
or U9968 (N_9968,N_7195,N_6727);
nor U9969 (N_9969,N_7760,N_7657);
nor U9970 (N_9970,N_7519,N_6618);
nand U9971 (N_9971,N_6695,N_6315);
nand U9972 (N_9972,N_7133,N_6967);
or U9973 (N_9973,N_7718,N_6045);
or U9974 (N_9974,N_6636,N_6712);
nand U9975 (N_9975,N_6475,N_6372);
nand U9976 (N_9976,N_6793,N_6879);
nor U9977 (N_9977,N_7423,N_7943);
nand U9978 (N_9978,N_6468,N_6808);
or U9979 (N_9979,N_6594,N_7713);
or U9980 (N_9980,N_7751,N_6518);
nand U9981 (N_9981,N_7643,N_7599);
nor U9982 (N_9982,N_6102,N_6475);
nand U9983 (N_9983,N_7039,N_6645);
or U9984 (N_9984,N_6732,N_6048);
or U9985 (N_9985,N_6935,N_7124);
nand U9986 (N_9986,N_7573,N_7737);
nand U9987 (N_9987,N_7999,N_7707);
or U9988 (N_9988,N_7480,N_7034);
or U9989 (N_9989,N_7407,N_6714);
nand U9990 (N_9990,N_6196,N_7790);
nand U9991 (N_9991,N_6883,N_6633);
or U9992 (N_9992,N_7104,N_7067);
and U9993 (N_9993,N_7910,N_6716);
nor U9994 (N_9994,N_7285,N_7549);
nor U9995 (N_9995,N_6270,N_6243);
nor U9996 (N_9996,N_6186,N_7673);
and U9997 (N_9997,N_6570,N_6051);
nor U9998 (N_9998,N_7009,N_7662);
or U9999 (N_9999,N_6902,N_6145);
nand UO_0 (O_0,N_9765,N_9877);
nand UO_1 (O_1,N_9682,N_9132);
nor UO_2 (O_2,N_9689,N_8671);
and UO_3 (O_3,N_9910,N_8675);
nand UO_4 (O_4,N_9511,N_9961);
and UO_5 (O_5,N_8480,N_8944);
nor UO_6 (O_6,N_9169,N_8875);
or UO_7 (O_7,N_8287,N_9977);
or UO_8 (O_8,N_8752,N_8054);
or UO_9 (O_9,N_8840,N_8750);
and UO_10 (O_10,N_8585,N_9659);
nand UO_11 (O_11,N_9879,N_8443);
nand UO_12 (O_12,N_9767,N_9321);
nand UO_13 (O_13,N_8324,N_9971);
or UO_14 (O_14,N_9542,N_9563);
and UO_15 (O_15,N_8793,N_8362);
or UO_16 (O_16,N_8406,N_9479);
and UO_17 (O_17,N_8327,N_8146);
nand UO_18 (O_18,N_9848,N_9196);
or UO_19 (O_19,N_8125,N_8274);
nor UO_20 (O_20,N_9964,N_8968);
or UO_21 (O_21,N_8971,N_8728);
nand UO_22 (O_22,N_9868,N_9601);
and UO_23 (O_23,N_8666,N_9438);
nor UO_24 (O_24,N_9535,N_8042);
and UO_25 (O_25,N_8495,N_9711);
nand UO_26 (O_26,N_8885,N_8498);
and UO_27 (O_27,N_8828,N_8296);
nand UO_28 (O_28,N_8580,N_8520);
nand UO_29 (O_29,N_8444,N_9249);
or UO_30 (O_30,N_9584,N_8800);
or UO_31 (O_31,N_8445,N_8414);
nand UO_32 (O_32,N_8733,N_9561);
or UO_33 (O_33,N_8094,N_8158);
nor UO_34 (O_34,N_8899,N_9189);
nand UO_35 (O_35,N_8252,N_9182);
or UO_36 (O_36,N_9137,N_8115);
nor UO_37 (O_37,N_8514,N_8240);
nor UO_38 (O_38,N_8391,N_9119);
and UO_39 (O_39,N_8487,N_8594);
or UO_40 (O_40,N_9636,N_9557);
nand UO_41 (O_41,N_9081,N_9047);
nand UO_42 (O_42,N_8477,N_9115);
xnor UO_43 (O_43,N_8832,N_9322);
or UO_44 (O_44,N_8893,N_9002);
or UO_45 (O_45,N_9443,N_9568);
or UO_46 (O_46,N_9324,N_8931);
or UO_47 (O_47,N_9477,N_8188);
nand UO_48 (O_48,N_8434,N_8182);
and UO_49 (O_49,N_8415,N_8166);
nor UO_50 (O_50,N_9257,N_8669);
or UO_51 (O_51,N_8954,N_9161);
nor UO_52 (O_52,N_8446,N_9095);
nor UO_53 (O_53,N_8597,N_9501);
nand UO_54 (O_54,N_8868,N_9459);
and UO_55 (O_55,N_9234,N_9295);
and UO_56 (O_56,N_9899,N_9688);
nor UO_57 (O_57,N_8276,N_9282);
or UO_58 (O_58,N_8651,N_8055);
nor UO_59 (O_59,N_8212,N_9394);
and UO_60 (O_60,N_8260,N_8199);
and UO_61 (O_61,N_8630,N_9934);
nor UO_62 (O_62,N_8482,N_8454);
or UO_63 (O_63,N_8400,N_9787);
nand UO_64 (O_64,N_8687,N_9344);
or UO_65 (O_65,N_9622,N_9198);
nor UO_66 (O_66,N_8164,N_8297);
nand UO_67 (O_67,N_8235,N_9147);
nand UO_68 (O_68,N_8229,N_8242);
or UO_69 (O_69,N_9401,N_9045);
and UO_70 (O_70,N_9068,N_9224);
nand UO_71 (O_71,N_9063,N_8243);
nor UO_72 (O_72,N_9426,N_9651);
or UO_73 (O_73,N_8626,N_9184);
nor UO_74 (O_74,N_8784,N_8790);
or UO_75 (O_75,N_9120,N_8973);
nand UO_76 (O_76,N_9398,N_8349);
nand UO_77 (O_77,N_9629,N_8140);
nor UO_78 (O_78,N_8535,N_9312);
nand UO_79 (O_79,N_8596,N_8171);
and UO_80 (O_80,N_9795,N_9415);
nor UO_81 (O_81,N_8371,N_9986);
nor UO_82 (O_82,N_8003,N_8841);
nand UO_83 (O_83,N_8088,N_8927);
nor UO_84 (O_84,N_9212,N_8262);
and UO_85 (O_85,N_8845,N_8325);
or UO_86 (O_86,N_9356,N_8447);
or UO_87 (O_87,N_8467,N_9240);
nor UO_88 (O_88,N_8072,N_8989);
nand UO_89 (O_89,N_9508,N_9607);
nor UO_90 (O_90,N_9476,N_8956);
nand UO_91 (O_91,N_8478,N_9875);
xnor UO_92 (O_92,N_9248,N_8746);
nor UO_93 (O_93,N_8364,N_8073);
nor UO_94 (O_94,N_9284,N_9980);
and UO_95 (O_95,N_9025,N_8223);
nand UO_96 (O_96,N_9325,N_9136);
and UO_97 (O_97,N_9761,N_9378);
and UO_98 (O_98,N_8079,N_8619);
nand UO_99 (O_99,N_9255,N_9128);
nand UO_100 (O_100,N_8078,N_8867);
nand UO_101 (O_101,N_8633,N_9088);
and UO_102 (O_102,N_8493,N_8040);
nor UO_103 (O_103,N_8184,N_8536);
nand UO_104 (O_104,N_9367,N_9959);
nand UO_105 (O_105,N_8465,N_9805);
nand UO_106 (O_106,N_9730,N_9044);
nor UO_107 (O_107,N_9118,N_9159);
or UO_108 (O_108,N_9849,N_8644);
nand UO_109 (O_109,N_8063,N_8114);
and UO_110 (O_110,N_9000,N_9071);
nand UO_111 (O_111,N_8431,N_9303);
nor UO_112 (O_112,N_8314,N_8494);
and UO_113 (O_113,N_8095,N_9702);
nand UO_114 (O_114,N_9363,N_9059);
nor UO_115 (O_115,N_8366,N_9171);
and UO_116 (O_116,N_9089,N_8322);
and UO_117 (O_117,N_8416,N_9432);
nand UO_118 (O_118,N_9251,N_8939);
and UO_119 (O_119,N_9751,N_9539);
and UO_120 (O_120,N_8578,N_9313);
or UO_121 (O_121,N_9353,N_9298);
nor UO_122 (O_122,N_8479,N_8216);
and UO_123 (O_123,N_8462,N_8375);
nor UO_124 (O_124,N_8238,N_9345);
nand UO_125 (O_125,N_8987,N_9262);
nand UO_126 (O_126,N_8312,N_8439);
and UO_127 (O_127,N_9509,N_9102);
and UO_128 (O_128,N_9012,N_8060);
nor UO_129 (O_129,N_9220,N_9552);
and UO_130 (O_130,N_9522,N_8550);
nand UO_131 (O_131,N_9897,N_9468);
nand UO_132 (O_132,N_9770,N_8113);
nand UO_133 (O_133,N_9085,N_8685);
and UO_134 (O_134,N_8678,N_9610);
nor UO_135 (O_135,N_9870,N_9299);
nor UO_136 (O_136,N_8858,N_9675);
or UO_137 (O_137,N_8138,N_9722);
and UO_138 (O_138,N_8882,N_9158);
and UO_139 (O_139,N_9117,N_9517);
nor UO_140 (O_140,N_8869,N_8802);
nor UO_141 (O_141,N_8378,N_8815);
nor UO_142 (O_142,N_9125,N_8118);
xnor UO_143 (O_143,N_8429,N_9811);
nor UO_144 (O_144,N_9888,N_9982);
nand UO_145 (O_145,N_9750,N_8782);
nor UO_146 (O_146,N_9287,N_9529);
nand UO_147 (O_147,N_8136,N_8048);
nor UO_148 (O_148,N_9828,N_9151);
nand UO_149 (O_149,N_9757,N_9792);
or UO_150 (O_150,N_9348,N_8700);
or UO_151 (O_151,N_8698,N_9619);
nor UO_152 (O_152,N_8451,N_8656);
and UO_153 (O_153,N_9652,N_9766);
nand UO_154 (O_154,N_9486,N_8665);
nand UO_155 (O_155,N_8284,N_8731);
nand UO_156 (O_156,N_9819,N_9233);
nor UO_157 (O_157,N_8455,N_8635);
or UO_158 (O_158,N_9153,N_8348);
and UO_159 (O_159,N_9188,N_9978);
and UO_160 (O_160,N_8066,N_9732);
and UO_161 (O_161,N_8211,N_8852);
and UO_162 (O_162,N_8387,N_8174);
nand UO_163 (O_163,N_9924,N_9241);
nand UO_164 (O_164,N_8350,N_9994);
nor UO_165 (O_165,N_9191,N_9365);
nor UO_166 (O_166,N_8604,N_8181);
and UO_167 (O_167,N_8299,N_8220);
nor UO_168 (O_168,N_8667,N_8126);
and UO_169 (O_169,N_9373,N_8689);
or UO_170 (O_170,N_9989,N_9519);
or UO_171 (O_171,N_8173,N_8137);
and UO_172 (O_172,N_9109,N_9166);
nand UO_173 (O_173,N_9793,N_9461);
or UO_174 (O_174,N_8425,N_9887);
nor UO_175 (O_175,N_9215,N_9167);
nor UO_176 (O_176,N_8374,N_9360);
nand UO_177 (O_177,N_8565,N_8310);
nand UO_178 (O_178,N_8770,N_9555);
or UO_179 (O_179,N_8949,N_9116);
nand UO_180 (O_180,N_9901,N_9134);
nor UO_181 (O_181,N_8153,N_8900);
nor UO_182 (O_182,N_9847,N_9510);
nand UO_183 (O_183,N_9328,N_8881);
nand UO_184 (O_184,N_9384,N_9856);
nand UO_185 (O_185,N_8552,N_9537);
and UO_186 (O_186,N_9335,N_8621);
nand UO_187 (O_187,N_9268,N_8386);
or UO_188 (O_188,N_9950,N_8873);
nand UO_189 (O_189,N_9747,N_8797);
nor UO_190 (O_190,N_9646,N_9800);
and UO_191 (O_191,N_8165,N_9574);
nand UO_192 (O_192,N_8313,N_9038);
and UO_193 (O_193,N_9326,N_9616);
nand UO_194 (O_194,N_9441,N_8693);
nand UO_195 (O_195,N_9009,N_9912);
and UO_196 (O_196,N_9445,N_9375);
and UO_197 (O_197,N_8600,N_8803);
nor UO_198 (O_198,N_8475,N_9370);
nor UO_199 (O_199,N_9114,N_8345);
nor UO_200 (O_200,N_9798,N_9826);
nor UO_201 (O_201,N_8877,N_9804);
or UO_202 (O_202,N_9381,N_8704);
or UO_203 (O_203,N_9049,N_9319);
nand UO_204 (O_204,N_8768,N_9187);
nand UO_205 (O_205,N_8527,N_8030);
or UO_206 (O_206,N_9281,N_8903);
nor UO_207 (O_207,N_8982,N_8518);
nor UO_208 (O_208,N_9157,N_8210);
or UO_209 (O_209,N_8609,N_8278);
or UO_210 (O_210,N_9180,N_8926);
nand UO_211 (O_211,N_9687,N_8582);
or UO_212 (O_212,N_8771,N_8807);
nor UO_213 (O_213,N_8833,N_9753);
and UO_214 (O_214,N_8021,N_8584);
and UO_215 (O_215,N_8266,N_8677);
or UO_216 (O_216,N_9504,N_8896);
nand UO_217 (O_217,N_9270,N_9968);
nor UO_218 (O_218,N_8329,N_8117);
nor UO_219 (O_219,N_9124,N_8718);
nor UO_220 (O_220,N_8449,N_8005);
and UO_221 (O_221,N_8418,N_9396);
and UO_222 (O_222,N_9222,N_9430);
nor UO_223 (O_223,N_9067,N_8464);
xor UO_224 (O_224,N_8910,N_9070);
and UO_225 (O_225,N_8397,N_9194);
and UO_226 (O_226,N_8344,N_8537);
nor UO_227 (O_227,N_9593,N_8340);
or UO_228 (O_228,N_9790,N_8224);
nor UO_229 (O_229,N_8791,N_9165);
and UO_230 (O_230,N_9640,N_8683);
nor UO_231 (O_231,N_9228,N_8037);
and UO_232 (O_232,N_8025,N_8301);
nor UO_233 (O_233,N_9039,N_8657);
nor UO_234 (O_234,N_8905,N_8300);
or UO_235 (O_235,N_8589,N_8742);
nand UO_236 (O_236,N_8501,N_9855);
or UO_237 (O_237,N_9949,N_9237);
and UO_238 (O_238,N_8682,N_9471);
or UO_239 (O_239,N_9015,N_8513);
nand UO_240 (O_240,N_9979,N_8196);
or UO_241 (O_241,N_9776,N_8909);
or UO_242 (O_242,N_8438,N_9421);
nand UO_243 (O_243,N_9832,N_8365);
or UO_244 (O_244,N_8059,N_9569);
xnor UO_245 (O_245,N_8028,N_8152);
and UO_246 (O_246,N_8214,N_8969);
nand UO_247 (O_247,N_9181,N_9974);
nor UO_248 (O_248,N_8461,N_8541);
nor UO_249 (O_249,N_9786,N_8844);
nor UO_250 (O_250,N_9531,N_9211);
or UO_251 (O_251,N_8197,N_8638);
nand UO_252 (O_252,N_8389,N_8050);
and UO_253 (O_253,N_8819,N_9668);
nand UO_254 (O_254,N_8856,N_8990);
nand UO_255 (O_255,N_8891,N_9200);
nor UO_256 (O_256,N_8504,N_8557);
nand UO_257 (O_257,N_8123,N_9083);
nand UO_258 (O_258,N_9410,N_9036);
nor UO_259 (O_259,N_9869,N_9528);
nand UO_260 (O_260,N_8920,N_9449);
and UO_261 (O_261,N_9480,N_8735);
and UO_262 (O_262,N_8979,N_9138);
nand UO_263 (O_263,N_9988,N_9331);
nor UO_264 (O_264,N_9041,N_9946);
and UO_265 (O_265,N_8044,N_8194);
or UO_266 (O_266,N_8039,N_8709);
or UO_267 (O_267,N_8328,N_9058);
nand UO_268 (O_268,N_8653,N_9976);
or UO_269 (O_269,N_9017,N_8924);
nor UO_270 (O_270,N_8147,N_9617);
nor UO_271 (O_271,N_8241,N_8823);
nor UO_272 (O_272,N_9097,N_9797);
nand UO_273 (O_273,N_8895,N_8601);
xnor UO_274 (O_274,N_9694,N_8654);
nand UO_275 (O_275,N_8918,N_8405);
and UO_276 (O_276,N_9156,N_8338);
and UO_277 (O_277,N_8069,N_9470);
or UO_278 (O_278,N_9473,N_9951);
nor UO_279 (O_279,N_9873,N_8865);
nand UO_280 (O_280,N_9272,N_8420);
nand UO_281 (O_281,N_8627,N_9882);
nand UO_282 (O_282,N_8821,N_8838);
and UO_283 (O_283,N_8859,N_9500);
nor UO_284 (O_284,N_8998,N_9148);
nor UO_285 (O_285,N_9462,N_9420);
or UO_286 (O_286,N_8440,N_9442);
xor UO_287 (O_287,N_9444,N_9639);
and UO_288 (O_288,N_9520,N_8046);
nor UO_289 (O_289,N_8052,N_8526);
nand UO_290 (O_290,N_9716,N_8563);
nor UO_291 (O_291,N_9301,N_9559);
and UO_292 (O_292,N_9999,N_9554);
or UO_293 (O_293,N_9698,N_8889);
nand UO_294 (O_294,N_8696,N_9496);
or UO_295 (O_295,N_8703,N_8019);
and UO_296 (O_296,N_8264,N_9371);
nand UO_297 (O_297,N_9472,N_8530);
nor UO_298 (O_298,N_8690,N_8294);
nor UO_299 (O_299,N_8629,N_8977);
nor UO_300 (O_300,N_8974,N_9595);
or UO_301 (O_301,N_9567,N_9507);
or UO_302 (O_302,N_9553,N_9831);
nor UO_303 (O_303,N_9708,N_8205);
and UO_304 (O_304,N_9290,N_9709);
nor UO_305 (O_305,N_8806,N_9772);
or UO_306 (O_306,N_9721,N_9960);
nand UO_307 (O_307,N_8936,N_8825);
nor UO_308 (O_308,N_9707,N_8670);
and UO_309 (O_309,N_9207,N_9860);
xor UO_310 (O_310,N_8599,N_9830);
or UO_311 (O_311,N_8236,N_9857);
nand UO_312 (O_312,N_9300,N_8180);
or UO_313 (O_313,N_9972,N_9635);
or UO_314 (O_314,N_9822,N_8641);
nand UO_315 (O_315,N_8051,N_8155);
or UO_316 (O_316,N_8065,N_9416);
and UO_317 (O_317,N_9582,N_9448);
and UO_318 (O_318,N_8228,N_8381);
nand UO_319 (O_319,N_9925,N_9874);
and UO_320 (O_320,N_9631,N_8437);
or UO_321 (O_321,N_9302,N_9674);
nor UO_322 (O_322,N_9955,N_8000);
or UO_323 (O_323,N_8623,N_9078);
nand UO_324 (O_324,N_8127,N_9076);
nand UO_325 (O_325,N_8539,N_9774);
nand UO_326 (O_326,N_8710,N_9431);
nor UO_327 (O_327,N_9992,N_8160);
nand UO_328 (O_328,N_9458,N_8128);
nor UO_329 (O_329,N_8170,N_8286);
nand UO_330 (O_330,N_8788,N_9122);
nor UO_331 (O_331,N_8333,N_8441);
nor UO_332 (O_332,N_9407,N_9763);
and UO_333 (O_333,N_9178,N_8290);
nor UO_334 (O_334,N_9852,N_9643);
and UO_335 (O_335,N_9838,N_8570);
nor UO_336 (O_336,N_9532,N_9842);
or UO_337 (O_337,N_9297,N_8795);
nand UO_338 (O_338,N_9176,N_8412);
xnor UO_339 (O_339,N_8524,N_9238);
nor UO_340 (O_340,N_9389,N_8660);
nor UO_341 (O_341,N_8029,N_8777);
and UO_342 (O_342,N_9032,N_8227);
or UO_343 (O_343,N_8749,N_8016);
nand UO_344 (O_344,N_8734,N_9362);
nand UO_345 (O_345,N_9417,N_9916);
or UO_346 (O_346,N_8435,N_9043);
nand UO_347 (O_347,N_8458,N_9706);
and UO_348 (O_348,N_8532,N_9627);
or UO_349 (O_349,N_8473,N_8688);
nand UO_350 (O_350,N_8648,N_8183);
nor UO_351 (O_351,N_8500,N_8679);
nand UO_352 (O_352,N_8195,N_9278);
or UO_353 (O_353,N_9625,N_8237);
nand UO_354 (O_354,N_9346,N_9231);
nor UO_355 (O_355,N_9928,N_8659);
and UO_356 (O_356,N_8760,N_8393);
nand UO_357 (O_357,N_9379,N_8036);
or UO_358 (O_358,N_8808,N_8942);
nand UO_359 (O_359,N_8448,N_8215);
nand UO_360 (O_360,N_9332,N_8139);
nand UO_361 (O_361,N_8714,N_8586);
or UO_362 (O_362,N_9727,N_9294);
or UO_363 (O_363,N_9383,N_9073);
nand UO_364 (O_364,N_8279,N_9466);
and UO_365 (O_365,N_8799,N_8606);
or UO_366 (O_366,N_9170,N_9991);
or UO_367 (O_367,N_9502,N_8367);
and UO_368 (O_368,N_8640,N_8298);
nand UO_369 (O_369,N_8817,N_8486);
nor UO_370 (O_370,N_9086,N_8853);
nand UO_371 (O_371,N_9611,N_8934);
or UO_372 (O_372,N_8064,N_9933);
nand UO_373 (O_373,N_9467,N_8551);
and UO_374 (O_374,N_9634,N_8528);
nor UO_375 (O_375,N_8038,N_8246);
nor UO_376 (O_376,N_8758,N_8135);
nor UO_377 (O_377,N_8874,N_9827);
nand UO_378 (O_378,N_8860,N_9696);
and UO_379 (O_379,N_8093,N_9139);
or UO_380 (O_380,N_9304,N_8639);
and UO_381 (O_381,N_8534,N_9638);
nand UO_382 (O_382,N_9921,N_9174);
and UO_383 (O_383,N_8729,N_9033);
nand UO_384 (O_384,N_9062,N_9141);
nor UO_385 (O_385,N_8617,N_8045);
or UO_386 (O_386,N_9666,N_8091);
nor UO_387 (O_387,N_9150,N_9057);
or UO_388 (O_388,N_9918,N_8245);
and UO_389 (O_389,N_9760,N_8732);
nand UO_390 (O_390,N_8457,N_9492);
nand UO_391 (O_391,N_9973,N_8142);
or UO_392 (O_392,N_8553,N_8024);
nor UO_393 (O_393,N_9010,N_8192);
and UO_394 (O_394,N_9351,N_8658);
or UO_395 (O_395,N_8144,N_9749);
or UO_396 (O_396,N_8169,N_8813);
or UO_397 (O_397,N_8506,N_8380);
nand UO_398 (O_398,N_8603,N_9720);
nand UO_399 (O_399,N_8738,N_9724);
nand UO_400 (O_400,N_8101,N_8232);
and UO_401 (O_401,N_9376,N_8295);
and UO_402 (O_402,N_9164,N_8363);
nand UO_403 (O_403,N_8980,N_9390);
nand UO_404 (O_404,N_8318,N_8883);
and UO_405 (O_405,N_8921,N_8319);
nand UO_406 (O_406,N_8549,N_9547);
and UO_407 (O_407,N_8943,N_9691);
nor UO_408 (O_408,N_8084,N_8254);
nor UO_409 (O_409,N_8577,N_8177);
nor UO_410 (O_410,N_9320,N_9665);
nor UO_411 (O_411,N_9144,N_8684);
nor UO_412 (O_412,N_9387,N_8104);
nand UO_413 (O_413,N_8612,N_8058);
or UO_414 (O_414,N_8624,N_9541);
nand UO_415 (O_415,N_9475,N_9409);
and UO_416 (O_416,N_9895,N_9745);
nor UO_417 (O_417,N_9437,N_8303);
and UO_418 (O_418,N_8453,N_8592);
nor UO_419 (O_419,N_9112,N_8157);
nand UO_420 (O_420,N_8542,N_8966);
nand UO_421 (O_421,N_8265,N_9662);
and UO_422 (O_422,N_9587,N_9173);
nor UO_423 (O_423,N_9658,N_8335);
or UO_424 (O_424,N_9906,N_9591);
nand UO_425 (O_425,N_8615,N_9392);
and UO_426 (O_426,N_9664,N_8130);
or UO_427 (O_427,N_8202,N_9019);
and UO_428 (O_428,N_9850,N_9050);
or UO_429 (O_429,N_9514,N_8090);
or UO_430 (O_430,N_9266,N_8581);
nand UO_431 (O_431,N_8470,N_9752);
or UO_432 (O_432,N_8976,N_9741);
and UO_433 (O_433,N_8331,N_8730);
and UO_434 (O_434,N_9337,N_9111);
and UO_435 (O_435,N_9549,N_8792);
and UO_436 (O_436,N_9368,N_9931);
nand UO_437 (O_437,N_8890,N_9903);
xnor UO_438 (O_438,N_9618,N_9311);
and UO_439 (O_439,N_8663,N_8781);
and UO_440 (O_440,N_8983,N_9523);
xnor UO_441 (O_441,N_8077,N_9100);
nand UO_442 (O_442,N_8106,N_8922);
xor UO_443 (O_443,N_9965,N_8080);
and UO_444 (O_444,N_9482,N_9740);
nand UO_445 (O_445,N_8953,N_9993);
or UO_446 (O_446,N_9149,N_8716);
and UO_447 (O_447,N_8964,N_9048);
nand UO_448 (O_448,N_9876,N_8020);
and UO_449 (O_449,N_9003,N_9079);
nand UO_450 (O_450,N_8250,N_9229);
nand UO_451 (O_451,N_8395,N_8200);
nor UO_452 (O_452,N_8488,N_9835);
nand UO_453 (O_453,N_8505,N_9686);
and UO_454 (O_454,N_8459,N_9104);
and UO_455 (O_455,N_8801,N_8306);
or UO_456 (O_456,N_9123,N_8089);
nand UO_457 (O_457,N_8851,N_8317);
nor UO_458 (O_458,N_8923,N_8826);
and UO_459 (O_459,N_9578,N_9883);
nand UO_460 (O_460,N_9656,N_9785);
nand UO_461 (O_461,N_8778,N_8672);
and UO_462 (O_462,N_9024,N_8219);
or UO_463 (O_463,N_9168,N_9613);
nor UO_464 (O_464,N_9710,N_8647);
nor UO_465 (O_465,N_9526,N_8929);
or UO_466 (O_466,N_8161,N_9521);
or UO_467 (O_467,N_9859,N_8272);
or UO_468 (O_468,N_9604,N_9435);
and UO_469 (O_469,N_9397,N_8512);
or UO_470 (O_470,N_9288,N_9594);
nor UO_471 (O_471,N_9013,N_9544);
nor UO_472 (O_472,N_9781,N_9440);
nor UO_473 (O_473,N_8886,N_8835);
or UO_474 (O_474,N_9515,N_8997);
or UO_475 (O_475,N_9612,N_8309);
nor UO_476 (O_476,N_8715,N_8277);
and UO_477 (O_477,N_8822,N_9155);
nand UO_478 (O_478,N_8359,N_8004);
and UO_479 (O_479,N_8256,N_9891);
or UO_480 (O_480,N_8593,N_8699);
nand UO_481 (O_481,N_9609,N_9323);
and UO_482 (O_482,N_9277,N_9446);
and UO_483 (O_483,N_8613,N_9391);
nand UO_484 (O_484,N_9645,N_8740);
nand UO_485 (O_485,N_9499,N_8846);
and UO_486 (O_486,N_9424,N_8010);
nor UO_487 (O_487,N_9624,N_8492);
or UO_488 (O_488,N_8775,N_9280);
nand UO_489 (O_489,N_8411,N_8408);
nor UO_490 (O_490,N_9935,N_9372);
nor UO_491 (O_491,N_8047,N_8385);
nor UO_492 (O_492,N_9518,N_9984);
nor UO_493 (O_493,N_9232,N_8427);
and UO_494 (O_494,N_8566,N_9427);
nor UO_495 (O_495,N_8756,N_8515);
and UO_496 (O_496,N_9914,N_9031);
and UO_497 (O_497,N_9179,N_8251);
or UO_498 (O_498,N_8209,N_9592);
nand UO_499 (O_499,N_9087,N_9863);
nand UO_500 (O_500,N_9400,N_8848);
or UO_501 (O_501,N_9690,N_8820);
or UO_502 (O_502,N_8785,N_8898);
nor UO_503 (O_503,N_8727,N_9271);
nor UO_504 (O_504,N_8062,N_8002);
nor UO_505 (O_505,N_9654,N_8884);
or UO_506 (O_506,N_8426,N_9395);
nor UO_507 (O_507,N_8743,N_8955);
nor UO_508 (O_508,N_8339,N_9536);
or UO_509 (O_509,N_9937,N_8794);
nor UO_510 (O_510,N_9004,N_8008);
and UO_511 (O_511,N_9789,N_9641);
or UO_512 (O_512,N_9065,N_8769);
nand UO_513 (O_513,N_8694,N_8267);
nor UO_514 (O_514,N_8945,N_9411);
and UO_515 (O_515,N_8424,N_8725);
nand UO_516 (O_516,N_8722,N_8620);
or UO_517 (O_517,N_9551,N_9713);
nor UO_518 (O_518,N_8087,N_8132);
or UO_519 (O_519,N_9399,N_9227);
or UO_520 (O_520,N_8022,N_8347);
or UO_521 (O_521,N_9650,N_8805);
or UO_522 (O_522,N_9769,N_8507);
nor UO_523 (O_523,N_9598,N_8928);
xor UO_524 (O_524,N_9602,N_9864);
nor UO_525 (O_525,N_8558,N_9199);
and UO_526 (O_526,N_9975,N_8863);
or UO_527 (O_527,N_8061,N_9020);
nand UO_528 (O_528,N_9943,N_8757);
xnor UO_529 (O_529,N_8765,N_8567);
nor UO_530 (O_530,N_8713,N_9731);
nor UO_531 (O_531,N_8814,N_8485);
nand UO_532 (O_532,N_8384,N_8637);
or UO_533 (O_533,N_9334,N_8293);
nand UO_534 (O_534,N_9885,N_8304);
and UO_535 (O_535,N_8097,N_9648);
or UO_536 (O_536,N_9318,N_9452);
or UO_537 (O_537,N_8396,N_8871);
nor UO_538 (O_538,N_9160,N_9712);
nand UO_539 (O_539,N_9803,N_9620);
or UO_540 (O_540,N_9201,N_9755);
or UO_541 (O_541,N_9764,N_9309);
and UO_542 (O_542,N_8233,N_8509);
and UO_543 (O_543,N_9226,N_9821);
or UO_544 (O_544,N_8914,N_9052);
nor UO_545 (O_545,N_8616,N_8311);
nor UO_546 (O_546,N_9001,N_8258);
nand UO_547 (O_547,N_9962,N_8655);
and UO_548 (O_548,N_8281,N_9908);
nand UO_549 (O_549,N_9970,N_8409);
and UO_550 (O_550,N_9154,N_9192);
nor UO_551 (O_551,N_9783,N_8156);
or UO_552 (O_552,N_9402,N_8354);
and UO_553 (O_553,N_8531,N_8291);
and UO_554 (O_554,N_9341,N_8984);
or UO_555 (O_555,N_9512,N_8519);
nor UO_556 (O_556,N_8489,N_9818);
nand UO_557 (O_557,N_8204,N_9824);
and UO_558 (O_558,N_9491,N_9223);
nand UO_559 (O_559,N_9213,N_8031);
nand UO_560 (O_560,N_9889,N_8259);
nor UO_561 (O_561,N_8239,N_9382);
and UO_562 (O_562,N_9243,N_8041);
nand UO_563 (O_563,N_9451,N_9843);
or UO_564 (O_564,N_8282,N_9205);
nand UO_565 (O_565,N_8452,N_8013);
and UO_566 (O_566,N_8661,N_8032);
and UO_567 (O_567,N_8320,N_9195);
nand UO_568 (O_568,N_9990,N_9600);
nand UO_569 (O_569,N_9524,N_9872);
or UO_570 (O_570,N_8402,N_9487);
and UO_571 (O_571,N_9902,N_9106);
or UO_572 (O_572,N_9190,N_8831);
or UO_573 (O_573,N_8428,N_9193);
nor UO_574 (O_574,N_9904,N_8755);
nand UO_575 (O_575,N_9737,N_9846);
and UO_576 (O_576,N_8056,N_8967);
or UO_577 (O_577,N_9366,N_8681);
nor UO_578 (O_578,N_8522,N_8148);
and UO_579 (O_579,N_8234,N_9743);
or UO_580 (O_580,N_9162,N_8351);
nor UO_581 (O_581,N_9796,N_8786);
or UO_582 (O_582,N_8105,N_9028);
and UO_583 (O_583,N_9131,N_9947);
nor UO_584 (O_584,N_9865,N_8285);
nand UO_585 (O_585,N_8421,N_9945);
and UO_586 (O_586,N_8634,N_9630);
or UO_587 (O_587,N_8568,N_8472);
and UO_588 (O_588,N_9746,N_9098);
nor UO_589 (O_589,N_8745,N_9406);
nand UO_590 (O_590,N_8560,N_8816);
and UO_591 (O_591,N_8739,N_8432);
nor UO_592 (O_592,N_8878,N_8787);
or UO_593 (O_593,N_8579,N_9715);
nand UO_594 (O_594,N_9208,N_9560);
and UO_595 (O_595,N_9014,N_9583);
and UO_596 (O_596,N_9540,N_8925);
or UO_597 (O_597,N_8076,N_9516);
nor UO_598 (O_598,N_8026,N_9726);
nor UO_599 (O_599,N_9940,N_9909);
and UO_600 (O_600,N_9703,N_8463);
nor UO_601 (O_601,N_9829,N_8422);
and UO_602 (O_602,N_9866,N_8717);
nor UO_603 (O_603,N_9314,N_9428);
nor UO_604 (O_604,N_8834,N_8403);
and UO_605 (O_605,N_9728,N_8902);
nand UO_606 (O_606,N_8680,N_9204);
and UO_607 (O_607,N_9505,N_8880);
nor UO_608 (O_608,N_8796,N_8218);
nor UO_609 (O_609,N_9525,N_8009);
or UO_610 (O_610,N_9930,N_9177);
and UO_611 (O_611,N_9253,N_8697);
and UO_612 (O_612,N_9754,N_9605);
xor UO_613 (O_613,N_9893,N_9285);
and UO_614 (O_614,N_8941,N_9210);
nor UO_615 (O_615,N_8830,N_9900);
nand UO_616 (O_616,N_8401,N_8720);
or UO_617 (O_617,N_8358,N_9506);
or UO_618 (O_618,N_8876,N_9305);
nor UO_619 (O_619,N_9572,N_8993);
nand UO_620 (O_620,N_9364,N_9684);
nor UO_621 (O_621,N_9573,N_8779);
nand UO_622 (O_622,N_8018,N_8643);
nand UO_623 (O_623,N_8145,N_8074);
and UO_624 (O_624,N_9632,N_9784);
nand UO_625 (O_625,N_9642,N_9758);
or UO_626 (O_626,N_9967,N_8747);
nor UO_627 (O_627,N_8767,N_8843);
nor UO_628 (O_628,N_8124,N_9806);
or UO_629 (O_629,N_9245,N_8748);
nand UO_630 (O_630,N_9898,N_9725);
nor UO_631 (O_631,N_8222,N_8836);
and UO_632 (O_632,N_9836,N_9172);
nand UO_633 (O_633,N_9361,N_8917);
nor UO_634 (O_634,N_8308,N_9729);
or UO_635 (O_635,N_9649,N_9562);
and UO_636 (O_636,N_9672,N_8861);
nand UO_637 (O_637,N_9538,N_8662);
or UO_638 (O_638,N_9355,N_9545);
and UO_639 (O_639,N_8608,N_9018);
nand UO_640 (O_640,N_9920,N_9927);
nor UO_641 (O_641,N_9692,N_8271);
or UO_642 (O_642,N_9660,N_8190);
nand UO_643 (O_643,N_9099,N_9216);
nor UO_644 (O_644,N_8083,N_8394);
or UO_645 (O_645,N_9008,N_8368);
and UO_646 (O_646,N_8706,N_8992);
or UO_647 (O_647,N_8517,N_8413);
or UO_648 (O_648,N_9289,N_8049);
nor UO_649 (O_649,N_9881,N_8372);
nand UO_650 (O_650,N_8912,N_9939);
nand UO_651 (O_651,N_9633,N_8499);
nand UO_652 (O_652,N_8510,N_8175);
or UO_653 (O_653,N_9621,N_8474);
nand UO_654 (O_654,N_8849,N_8963);
nand UO_655 (O_655,N_9336,N_8316);
xor UO_656 (O_656,N_9952,N_9225);
and UO_657 (O_657,N_9352,N_8419);
nand UO_658 (O_658,N_8189,N_9077);
nand UO_659 (O_659,N_8598,N_8764);
and UO_660 (O_660,N_8556,N_9209);
nand UO_661 (O_661,N_9006,N_8185);
and UO_662 (O_662,N_9113,N_9439);
nor UO_663 (O_663,N_9615,N_8538);
or UO_664 (O_664,N_9966,N_9723);
nand UO_665 (O_665,N_8086,N_8894);
and UO_666 (O_666,N_8602,N_9839);
or UO_667 (O_667,N_9279,N_9074);
and UO_668 (O_668,N_9941,N_8650);
nand UO_669 (O_669,N_9546,N_9082);
nor UO_670 (O_670,N_8270,N_8761);
nor UO_671 (O_671,N_8576,N_9543);
and UO_672 (O_672,N_9329,N_9606);
nand UO_673 (O_673,N_8525,N_9236);
nor UO_674 (O_674,N_9714,N_8695);
nand UO_675 (O_675,N_9217,N_9588);
or UO_676 (O_676,N_8547,N_9586);
or UO_677 (O_677,N_9046,N_9056);
nand UO_678 (O_678,N_9425,N_8085);
nor UO_679 (O_679,N_8323,N_8053);
or UO_680 (O_680,N_9474,N_8573);
nor UO_681 (O_681,N_9359,N_9135);
nand UO_682 (O_682,N_9533,N_8466);
nand UO_683 (O_683,N_8569,N_9867);
nor UO_684 (O_684,N_9093,N_9307);
nor UO_685 (O_685,N_9069,N_9779);
and UO_686 (O_686,N_9197,N_9944);
and UO_687 (O_687,N_9369,N_8543);
or UO_688 (O_688,N_8850,N_8471);
and UO_689 (O_689,N_8460,N_9388);
nand UO_690 (O_690,N_8332,N_8149);
nor UO_691 (O_691,N_9274,N_8523);
or UO_692 (O_692,N_9628,N_8203);
nor UO_693 (O_693,N_9956,N_8150);
and UO_694 (O_694,N_8737,N_9465);
nand UO_695 (O_695,N_9485,N_8972);
or UO_696 (O_696,N_8879,N_9825);
nor UO_697 (O_697,N_9414,N_8015);
or UO_698 (O_698,N_9550,N_9423);
nand UO_699 (O_699,N_8162,N_8159);
nor UO_700 (O_700,N_8719,N_8870);
nor UO_701 (O_701,N_9090,N_9896);
nor UO_702 (O_702,N_8373,N_9239);
or UO_703 (O_703,N_9385,N_8911);
nor UO_704 (O_704,N_8111,N_9996);
nor UO_705 (O_705,N_9075,N_8996);
nor UO_706 (O_706,N_9484,N_9963);
or UO_707 (O_707,N_9953,N_8529);
nor UO_708 (O_708,N_8533,N_9697);
and UO_709 (O_709,N_9347,N_8932);
nand UO_710 (O_710,N_9503,N_8108);
nand UO_711 (O_711,N_8935,N_8605);
or UO_712 (O_712,N_9556,N_9673);
or UO_713 (O_713,N_8321,N_8390);
nor UO_714 (O_714,N_9969,N_9023);
or UO_715 (O_715,N_8201,N_9405);
or UO_716 (O_716,N_8417,N_9527);
or UO_717 (O_717,N_9403,N_8186);
or UO_718 (O_718,N_8986,N_8330);
nand UO_719 (O_719,N_8433,N_8337);
and UO_720 (O_720,N_9663,N_9878);
or UO_721 (O_721,N_9814,N_9815);
nor UO_722 (O_722,N_9676,N_8490);
nand UO_723 (O_723,N_8904,N_9308);
or UO_724 (O_724,N_8107,N_9837);
nor UO_725 (O_725,N_8774,N_9478);
or UO_726 (O_726,N_8810,N_9599);
nor UO_727 (O_727,N_9339,N_8591);
nor UO_728 (O_728,N_9130,N_9218);
or UO_729 (O_729,N_8555,N_8023);
nand UO_730 (O_730,N_8948,N_8721);
nor UO_731 (O_731,N_9699,N_9580);
and UO_732 (O_732,N_8178,N_8864);
or UO_733 (O_733,N_9267,N_9291);
nor UO_734 (O_734,N_8965,N_9490);
and UO_735 (O_735,N_9072,N_9744);
or UO_736 (O_736,N_8554,N_9489);
or UO_737 (O_737,N_9954,N_9330);
nor UO_738 (O_738,N_8244,N_9434);
nand UO_739 (O_739,N_9488,N_9037);
or UO_740 (O_740,N_8208,N_9575);
and UO_741 (O_741,N_9778,N_8940);
nor UO_742 (O_742,N_9146,N_9812);
nand UO_743 (O_743,N_8842,N_9777);
nor UO_744 (O_744,N_8789,N_9739);
nor UO_745 (O_745,N_8957,N_8221);
nor UO_746 (O_746,N_8268,N_9080);
nor UO_747 (O_747,N_8154,N_9061);
nand UO_748 (O_748,N_9809,N_9005);
or UO_749 (O_749,N_9817,N_8590);
and UO_750 (O_750,N_8958,N_9719);
or UO_751 (O_751,N_9589,N_8508);
and UO_752 (O_752,N_8292,N_8574);
or UO_753 (O_753,N_9260,N_8827);
and UO_754 (O_754,N_9327,N_8172);
nand UO_755 (O_755,N_8120,N_9316);
nor UO_756 (O_756,N_8360,N_9317);
xor UO_757 (O_757,N_9734,N_8248);
nor UO_758 (O_758,N_8017,N_9021);
nor UO_759 (O_759,N_9890,N_8151);
and UO_760 (O_760,N_8082,N_9498);
nor UO_761 (O_761,N_9263,N_9221);
and UO_762 (O_762,N_9614,N_9055);
nand UO_763 (O_763,N_9565,N_8872);
nand UO_764 (O_764,N_9923,N_9064);
nand UO_765 (O_765,N_9293,N_9027);
and UO_766 (O_766,N_9655,N_8253);
nor UO_767 (O_767,N_8999,N_9029);
nand UO_768 (O_768,N_9775,N_8571);
nand UO_769 (O_769,N_9011,N_9823);
nor UO_770 (O_770,N_8377,N_9564);
nor UO_771 (O_771,N_8960,N_9374);
nand UO_772 (O_772,N_8342,N_8686);
nand UO_773 (O_773,N_8110,N_8607);
or UO_774 (O_774,N_8798,N_9608);
nor UO_775 (O_775,N_8930,N_9469);
nand UO_776 (O_776,N_9998,N_8692);
nand UO_777 (O_777,N_8649,N_9603);
nor UO_778 (O_778,N_9026,N_9661);
or UO_779 (O_779,N_8652,N_8341);
or UO_780 (O_780,N_8230,N_8847);
or UO_781 (O_781,N_9700,N_9084);
nor UO_782 (O_782,N_9840,N_8947);
nand UO_783 (O_783,N_9040,N_8288);
nand UO_784 (O_784,N_9762,N_9338);
nand UO_785 (O_785,N_9259,N_9246);
nor UO_786 (O_786,N_8033,N_8356);
or UO_787 (O_787,N_8206,N_8625);
and UO_788 (O_788,N_9590,N_9788);
nor UO_789 (O_789,N_9143,N_9858);
or UO_790 (O_790,N_9597,N_8357);
nor UO_791 (O_791,N_8766,N_8610);
or UO_792 (O_792,N_9261,N_9463);
nor UO_793 (O_793,N_8561,N_8007);
nand UO_794 (O_794,N_9186,N_8668);
nand UO_795 (O_795,N_9094,N_8001);
nand UO_796 (O_796,N_8207,N_8773);
or UO_797 (O_797,N_8071,N_8636);
and UO_798 (O_798,N_9342,N_8937);
and UO_799 (O_799,N_8481,N_9315);
nand UO_800 (O_800,N_9418,N_8632);
or UO_801 (O_801,N_9570,N_8548);
and UO_802 (O_802,N_8887,N_9653);
nand UO_803 (O_803,N_9513,N_8430);
and UO_804 (O_804,N_8255,N_8991);
nor UO_805 (O_805,N_9756,N_9042);
xor UO_806 (O_806,N_9497,N_8131);
nor UO_807 (O_807,N_8352,N_9091);
and UO_808 (O_808,N_8133,N_8736);
or UO_809 (O_809,N_9693,N_9886);
nand UO_810 (O_810,N_8141,N_9913);
or UO_811 (O_811,N_9942,N_8067);
nand UO_812 (O_812,N_9626,N_9717);
and UO_813 (O_813,N_9296,N_9704);
or UO_814 (O_814,N_8575,N_9358);
and UO_815 (O_815,N_8263,N_9422);
nor UO_816 (O_816,N_8398,N_8545);
nor UO_817 (O_817,N_8198,N_9258);
nor UO_818 (O_818,N_8121,N_9493);
nor UO_819 (O_819,N_8343,N_9412);
nor UO_820 (O_820,N_8564,N_8981);
and UO_821 (O_821,N_9349,N_8119);
nor UO_822 (O_822,N_9457,N_8933);
or UO_823 (O_823,N_8383,N_9671);
or UO_824 (O_824,N_8754,N_8167);
nand UO_825 (O_825,N_9264,N_9292);
and UO_826 (O_826,N_8622,N_8961);
and UO_827 (O_827,N_8355,N_9183);
and UO_828 (O_828,N_8283,N_8780);
or UO_829 (O_829,N_8497,N_9738);
nand UO_830 (O_830,N_9230,N_9834);
and UO_831 (O_831,N_9140,N_9911);
nand UO_832 (O_832,N_8280,N_9007);
and UO_833 (O_833,N_9782,N_9733);
nor UO_834 (O_834,N_8404,N_9035);
or UO_835 (O_835,N_8450,N_8857);
and UO_836 (O_836,N_8096,N_8913);
and UO_837 (O_837,N_9286,N_9558);
or UO_838 (O_838,N_9380,N_9917);
and UO_839 (O_839,N_9810,N_8273);
nand UO_840 (O_840,N_8901,N_9343);
nand UO_841 (O_841,N_8915,N_9142);
and UO_842 (O_842,N_9310,N_8103);
and UO_843 (O_843,N_9107,N_8673);
nor UO_844 (O_844,N_8511,N_8908);
or UO_845 (O_845,N_9129,N_8257);
nor UO_846 (O_846,N_8631,N_8759);
nor UO_847 (O_847,N_9748,N_9735);
nand UO_848 (O_848,N_8226,N_8962);
and UO_849 (O_849,N_9016,N_8469);
nand UO_850 (O_850,N_9453,N_8741);
nor UO_851 (O_851,N_8916,N_9103);
and UO_852 (O_852,N_9919,N_8100);
nand UO_853 (O_853,N_8163,N_9202);
and UO_854 (O_854,N_9780,N_8225);
nand UO_855 (O_855,N_8057,N_9455);
nor UO_856 (O_856,N_9948,N_9844);
and UO_857 (O_857,N_8572,N_8975);
nand UO_858 (O_858,N_8583,N_9736);
nor UO_859 (O_859,N_8027,N_8382);
and UO_860 (O_860,N_8483,N_8664);
nor UO_861 (O_861,N_8702,N_9685);
nand UO_862 (O_862,N_9022,N_8407);
or UO_863 (O_863,N_9571,N_8034);
or UO_864 (O_864,N_8540,N_9801);
nor UO_865 (O_865,N_9121,N_9851);
or UO_866 (O_866,N_9377,N_8109);
and UO_867 (O_867,N_9861,N_8112);
nand UO_868 (O_868,N_9596,N_9929);
or UO_869 (O_869,N_9853,N_8410);
nor UO_870 (O_870,N_8011,N_9957);
and UO_871 (O_871,N_9742,N_9256);
or UO_872 (O_872,N_9680,N_9585);
and UO_873 (O_873,N_8217,N_9481);
or UO_874 (O_874,N_8484,N_9333);
nand UO_875 (O_875,N_9254,N_8370);
and UO_876 (O_876,N_9841,N_8809);
or UO_877 (O_877,N_9915,N_8676);
nor UO_878 (O_878,N_8906,N_9203);
and UO_879 (O_879,N_8456,N_9030);
nand UO_880 (O_880,N_8723,N_8092);
nand UO_881 (O_881,N_8919,N_8744);
nand UO_882 (O_882,N_9433,N_9581);
nor UO_883 (O_883,N_9816,N_8866);
nor UO_884 (O_884,N_8907,N_9454);
nand UO_885 (O_885,N_8829,N_9637);
or UO_886 (O_886,N_9219,N_8191);
or UO_887 (O_887,N_8099,N_8353);
nand UO_888 (O_888,N_9791,N_8701);
nand UO_889 (O_889,N_9242,N_9252);
nand UO_890 (O_890,N_8705,N_8985);
nand UO_891 (O_891,N_8753,N_9958);
and UO_892 (O_892,N_8334,N_9436);
nand UO_893 (O_893,N_9429,N_9579);
nand UO_894 (O_894,N_9244,N_8892);
or UO_895 (O_895,N_8888,N_8116);
nor UO_896 (O_896,N_8854,N_9456);
nor UO_897 (O_897,N_9350,N_8336);
nand UO_898 (O_898,N_8812,N_9820);
or UO_899 (O_899,N_8897,N_9133);
or UO_900 (O_900,N_8946,N_8307);
or UO_901 (O_901,N_9404,N_9413);
or UO_902 (O_902,N_8952,N_9548);
and UO_903 (O_903,N_9995,N_9932);
and UO_904 (O_904,N_9283,N_9105);
and UO_905 (O_905,N_9054,N_9110);
and UO_906 (O_906,N_9667,N_8959);
or UO_907 (O_907,N_8707,N_9214);
or UO_908 (O_908,N_9306,N_8502);
or UO_909 (O_909,N_8436,N_8562);
nand UO_910 (O_910,N_8818,N_9926);
nand UO_911 (O_911,N_8376,N_8559);
nor UO_912 (O_912,N_8994,N_9677);
and UO_913 (O_913,N_8711,N_8995);
nand UO_914 (O_914,N_9670,N_9534);
nand UO_915 (O_915,N_9759,N_8168);
or UO_916 (O_916,N_8176,N_9705);
nand UO_917 (O_917,N_8326,N_8804);
or UO_918 (O_918,N_8708,N_8122);
nor UO_919 (O_919,N_8645,N_9386);
nand UO_920 (O_920,N_8193,N_9108);
or UO_921 (O_921,N_9495,N_9247);
nand UO_922 (O_922,N_8302,N_8491);
nand UO_923 (O_923,N_8305,N_8614);
or UO_924 (O_924,N_9892,N_9393);
nand UO_925 (O_925,N_9845,N_9718);
nor UO_926 (O_926,N_8503,N_8179);
nor UO_927 (O_927,N_9060,N_8261);
and UO_928 (O_928,N_8346,N_8275);
nor UO_929 (O_929,N_9768,N_9794);
and UO_930 (O_930,N_9152,N_8776);
and UO_931 (O_931,N_9905,N_9269);
nand UO_932 (O_932,N_9894,N_9530);
and UO_933 (O_933,N_9808,N_9408);
and UO_934 (O_934,N_8043,N_8712);
and UO_935 (O_935,N_9447,N_8361);
or UO_936 (O_936,N_8674,N_9273);
nand UO_937 (O_937,N_8068,N_8269);
nand UO_938 (O_938,N_9871,N_9034);
nor UO_939 (O_939,N_8951,N_8938);
nor UO_940 (O_940,N_8772,N_9175);
nor UO_941 (O_941,N_8388,N_9576);
nand UO_942 (O_942,N_9802,N_8496);
nand UO_943 (O_943,N_9206,N_8521);
and UO_944 (O_944,N_9679,N_9450);
or UO_945 (O_945,N_9127,N_9833);
or UO_946 (O_946,N_9126,N_9185);
nand UO_947 (O_947,N_9862,N_9265);
nor UO_948 (O_948,N_9657,N_9145);
nand UO_949 (O_949,N_9813,N_9096);
nor UO_950 (O_950,N_9235,N_9681);
nor UO_951 (O_951,N_8081,N_9695);
and UO_952 (O_952,N_8315,N_9678);
or UO_953 (O_953,N_9983,N_9647);
or UO_954 (O_954,N_9771,N_8006);
nand UO_955 (O_955,N_8399,N_9483);
or UO_956 (O_956,N_8247,N_8442);
nor UO_957 (O_957,N_8546,N_9340);
nor UO_958 (O_958,N_9922,N_9807);
nand UO_959 (O_959,N_9101,N_8950);
xnor UO_960 (O_960,N_8611,N_9460);
and UO_961 (O_961,N_8249,N_8628);
and UO_962 (O_962,N_8143,N_9669);
nand UO_963 (O_963,N_8783,N_8102);
and UO_964 (O_964,N_8129,N_8855);
nor UO_965 (O_965,N_8726,N_8595);
or UO_966 (O_966,N_8379,N_8014);
and UO_967 (O_967,N_8646,N_8392);
xor UO_968 (O_968,N_8231,N_9354);
nand UO_969 (O_969,N_9985,N_8618);
nand UO_970 (O_970,N_8369,N_8811);
and UO_971 (O_971,N_9250,N_8751);
and UO_972 (O_972,N_9419,N_9683);
and UO_973 (O_973,N_9880,N_9577);
or UO_974 (O_974,N_8423,N_9907);
nand UO_975 (O_975,N_8516,N_9644);
or UO_976 (O_976,N_8691,N_8213);
and UO_977 (O_977,N_8724,N_9799);
or UO_978 (O_978,N_8587,N_9701);
or UO_979 (O_979,N_8837,N_9053);
or UO_980 (O_980,N_9936,N_9163);
nand UO_981 (O_981,N_9092,N_8289);
nand UO_982 (O_982,N_9981,N_8012);
nand UO_983 (O_983,N_8075,N_9854);
or UO_984 (O_984,N_9773,N_9884);
nand UO_985 (O_985,N_8187,N_8544);
nor UO_986 (O_986,N_9938,N_8839);
and UO_987 (O_987,N_9623,N_9051);
or UO_988 (O_988,N_8978,N_8588);
nand UO_989 (O_989,N_9997,N_9987);
xnor UO_990 (O_990,N_8970,N_8476);
or UO_991 (O_991,N_9276,N_9566);
nor UO_992 (O_992,N_8098,N_8824);
nand UO_993 (O_993,N_9066,N_8134);
nand UO_994 (O_994,N_8988,N_8468);
or UO_995 (O_995,N_9357,N_8763);
and UO_996 (O_996,N_8035,N_8070);
nor UO_997 (O_997,N_8862,N_9275);
nor UO_998 (O_998,N_9464,N_8762);
or UO_999 (O_999,N_9494,N_8642);
nor UO_1000 (O_1000,N_8769,N_8248);
and UO_1001 (O_1001,N_8017,N_8011);
nor UO_1002 (O_1002,N_8594,N_9825);
nor UO_1003 (O_1003,N_8873,N_8827);
nor UO_1004 (O_1004,N_8468,N_8433);
nor UO_1005 (O_1005,N_9053,N_9994);
nor UO_1006 (O_1006,N_8961,N_9072);
nor UO_1007 (O_1007,N_8227,N_8916);
nand UO_1008 (O_1008,N_8948,N_9477);
nor UO_1009 (O_1009,N_8383,N_8563);
or UO_1010 (O_1010,N_9046,N_9725);
or UO_1011 (O_1011,N_8290,N_9702);
nor UO_1012 (O_1012,N_9266,N_8211);
nand UO_1013 (O_1013,N_8259,N_9253);
or UO_1014 (O_1014,N_9547,N_9762);
or UO_1015 (O_1015,N_8776,N_9192);
nor UO_1016 (O_1016,N_8862,N_9658);
or UO_1017 (O_1017,N_9359,N_8113);
nand UO_1018 (O_1018,N_8626,N_8789);
and UO_1019 (O_1019,N_8491,N_9589);
nand UO_1020 (O_1020,N_9220,N_9710);
nand UO_1021 (O_1021,N_9196,N_8015);
nor UO_1022 (O_1022,N_9313,N_9563);
or UO_1023 (O_1023,N_8707,N_8234);
nand UO_1024 (O_1024,N_8833,N_9354);
nand UO_1025 (O_1025,N_9211,N_9537);
nand UO_1026 (O_1026,N_8711,N_9982);
or UO_1027 (O_1027,N_9199,N_8098);
or UO_1028 (O_1028,N_9720,N_8467);
nand UO_1029 (O_1029,N_9016,N_8254);
nor UO_1030 (O_1030,N_9698,N_9744);
or UO_1031 (O_1031,N_9734,N_8097);
nor UO_1032 (O_1032,N_9841,N_8030);
nand UO_1033 (O_1033,N_9672,N_9927);
or UO_1034 (O_1034,N_8806,N_9739);
or UO_1035 (O_1035,N_8992,N_9463);
nor UO_1036 (O_1036,N_9862,N_9794);
nand UO_1037 (O_1037,N_8197,N_8118);
or UO_1038 (O_1038,N_9689,N_8109);
or UO_1039 (O_1039,N_9010,N_8588);
nand UO_1040 (O_1040,N_8725,N_8896);
nand UO_1041 (O_1041,N_8048,N_9915);
or UO_1042 (O_1042,N_9526,N_9947);
nand UO_1043 (O_1043,N_9119,N_9312);
and UO_1044 (O_1044,N_9318,N_8573);
and UO_1045 (O_1045,N_8110,N_9578);
and UO_1046 (O_1046,N_8541,N_9216);
and UO_1047 (O_1047,N_9990,N_9510);
nor UO_1048 (O_1048,N_9989,N_8088);
nor UO_1049 (O_1049,N_8539,N_8369);
and UO_1050 (O_1050,N_8560,N_9040);
nand UO_1051 (O_1051,N_9756,N_9018);
nand UO_1052 (O_1052,N_9055,N_8021);
nor UO_1053 (O_1053,N_8692,N_9049);
or UO_1054 (O_1054,N_8697,N_9640);
nor UO_1055 (O_1055,N_8481,N_9353);
and UO_1056 (O_1056,N_8856,N_8775);
or UO_1057 (O_1057,N_8762,N_9895);
or UO_1058 (O_1058,N_9547,N_8910);
nor UO_1059 (O_1059,N_8555,N_8483);
nand UO_1060 (O_1060,N_9877,N_8810);
or UO_1061 (O_1061,N_9478,N_8169);
nor UO_1062 (O_1062,N_9092,N_9645);
or UO_1063 (O_1063,N_8614,N_9668);
and UO_1064 (O_1064,N_9743,N_8312);
nor UO_1065 (O_1065,N_8737,N_9490);
nand UO_1066 (O_1066,N_8122,N_8421);
and UO_1067 (O_1067,N_8813,N_8677);
and UO_1068 (O_1068,N_8489,N_9296);
nand UO_1069 (O_1069,N_9336,N_8403);
nand UO_1070 (O_1070,N_9027,N_8145);
nor UO_1071 (O_1071,N_8488,N_8793);
and UO_1072 (O_1072,N_9955,N_8463);
or UO_1073 (O_1073,N_8955,N_8954);
nand UO_1074 (O_1074,N_9554,N_9432);
nand UO_1075 (O_1075,N_8231,N_9005);
or UO_1076 (O_1076,N_9506,N_8565);
nand UO_1077 (O_1077,N_8342,N_8076);
or UO_1078 (O_1078,N_9837,N_8556);
nand UO_1079 (O_1079,N_8212,N_8510);
nor UO_1080 (O_1080,N_8286,N_9133);
and UO_1081 (O_1081,N_9890,N_8696);
and UO_1082 (O_1082,N_9142,N_8265);
and UO_1083 (O_1083,N_9204,N_9647);
nor UO_1084 (O_1084,N_9435,N_9201);
or UO_1085 (O_1085,N_8482,N_9112);
or UO_1086 (O_1086,N_9596,N_9498);
nand UO_1087 (O_1087,N_9536,N_9548);
and UO_1088 (O_1088,N_8254,N_8235);
nand UO_1089 (O_1089,N_8943,N_8319);
nor UO_1090 (O_1090,N_9283,N_9583);
nor UO_1091 (O_1091,N_9774,N_8486);
nand UO_1092 (O_1092,N_9427,N_8183);
or UO_1093 (O_1093,N_9995,N_8541);
and UO_1094 (O_1094,N_8559,N_9011);
nand UO_1095 (O_1095,N_8804,N_8458);
or UO_1096 (O_1096,N_8807,N_8125);
nor UO_1097 (O_1097,N_9918,N_8887);
or UO_1098 (O_1098,N_8265,N_8432);
or UO_1099 (O_1099,N_9362,N_9474);
or UO_1100 (O_1100,N_8721,N_8797);
or UO_1101 (O_1101,N_8484,N_9055);
or UO_1102 (O_1102,N_8041,N_9628);
nor UO_1103 (O_1103,N_8923,N_8655);
and UO_1104 (O_1104,N_8751,N_8262);
nand UO_1105 (O_1105,N_8544,N_9479);
and UO_1106 (O_1106,N_8594,N_8681);
or UO_1107 (O_1107,N_9927,N_9730);
and UO_1108 (O_1108,N_9534,N_8156);
or UO_1109 (O_1109,N_9024,N_9669);
nand UO_1110 (O_1110,N_8953,N_9395);
nor UO_1111 (O_1111,N_9148,N_8321);
nor UO_1112 (O_1112,N_8831,N_8371);
or UO_1113 (O_1113,N_9874,N_8457);
nor UO_1114 (O_1114,N_9945,N_9601);
or UO_1115 (O_1115,N_8045,N_8623);
nand UO_1116 (O_1116,N_8401,N_9720);
nor UO_1117 (O_1117,N_8765,N_8520);
and UO_1118 (O_1118,N_9904,N_8870);
or UO_1119 (O_1119,N_8433,N_8827);
nor UO_1120 (O_1120,N_8237,N_9009);
or UO_1121 (O_1121,N_9338,N_9560);
nor UO_1122 (O_1122,N_8085,N_8271);
and UO_1123 (O_1123,N_8123,N_8625);
nor UO_1124 (O_1124,N_9772,N_8485);
and UO_1125 (O_1125,N_9312,N_9728);
nor UO_1126 (O_1126,N_9981,N_9052);
and UO_1127 (O_1127,N_8415,N_8741);
nor UO_1128 (O_1128,N_9554,N_9957);
nand UO_1129 (O_1129,N_8855,N_9964);
or UO_1130 (O_1130,N_8977,N_9819);
and UO_1131 (O_1131,N_8357,N_8977);
and UO_1132 (O_1132,N_8565,N_9260);
nor UO_1133 (O_1133,N_9662,N_8538);
or UO_1134 (O_1134,N_8216,N_8510);
nor UO_1135 (O_1135,N_9513,N_8425);
nand UO_1136 (O_1136,N_8159,N_9649);
and UO_1137 (O_1137,N_8579,N_9888);
nor UO_1138 (O_1138,N_9821,N_8332);
nor UO_1139 (O_1139,N_9254,N_9016);
nand UO_1140 (O_1140,N_8028,N_8673);
nor UO_1141 (O_1141,N_9457,N_9932);
or UO_1142 (O_1142,N_9022,N_9562);
nand UO_1143 (O_1143,N_8713,N_9156);
nand UO_1144 (O_1144,N_8633,N_9489);
and UO_1145 (O_1145,N_8573,N_9052);
and UO_1146 (O_1146,N_9277,N_8138);
xor UO_1147 (O_1147,N_8108,N_9937);
or UO_1148 (O_1148,N_8628,N_9588);
and UO_1149 (O_1149,N_8197,N_9195);
and UO_1150 (O_1150,N_9510,N_8743);
nor UO_1151 (O_1151,N_9587,N_9664);
and UO_1152 (O_1152,N_9487,N_9447);
and UO_1153 (O_1153,N_9932,N_9212);
and UO_1154 (O_1154,N_8408,N_8481);
and UO_1155 (O_1155,N_8095,N_8712);
nor UO_1156 (O_1156,N_8766,N_9106);
nor UO_1157 (O_1157,N_9602,N_9535);
nand UO_1158 (O_1158,N_9699,N_8947);
or UO_1159 (O_1159,N_8434,N_9839);
nand UO_1160 (O_1160,N_8369,N_8043);
and UO_1161 (O_1161,N_9034,N_8148);
nor UO_1162 (O_1162,N_9257,N_9430);
nand UO_1163 (O_1163,N_8782,N_9839);
nor UO_1164 (O_1164,N_8819,N_8735);
xor UO_1165 (O_1165,N_9939,N_8560);
nor UO_1166 (O_1166,N_8004,N_9701);
and UO_1167 (O_1167,N_9245,N_9282);
nor UO_1168 (O_1168,N_8872,N_8231);
and UO_1169 (O_1169,N_8373,N_9394);
or UO_1170 (O_1170,N_8971,N_9443);
nor UO_1171 (O_1171,N_9027,N_8692);
nand UO_1172 (O_1172,N_8764,N_9440);
and UO_1173 (O_1173,N_8485,N_9270);
or UO_1174 (O_1174,N_9842,N_9920);
nor UO_1175 (O_1175,N_9512,N_8020);
nand UO_1176 (O_1176,N_8670,N_9577);
nor UO_1177 (O_1177,N_8485,N_9956);
nor UO_1178 (O_1178,N_8362,N_8152);
nand UO_1179 (O_1179,N_9019,N_9696);
nand UO_1180 (O_1180,N_8711,N_9411);
and UO_1181 (O_1181,N_9092,N_8234);
or UO_1182 (O_1182,N_8947,N_8901);
nand UO_1183 (O_1183,N_9333,N_9461);
nand UO_1184 (O_1184,N_8469,N_9905);
nor UO_1185 (O_1185,N_8270,N_8476);
or UO_1186 (O_1186,N_8677,N_8422);
nor UO_1187 (O_1187,N_8726,N_8229);
nor UO_1188 (O_1188,N_8718,N_9986);
nor UO_1189 (O_1189,N_9091,N_9655);
or UO_1190 (O_1190,N_8638,N_9970);
nand UO_1191 (O_1191,N_9465,N_8050);
nand UO_1192 (O_1192,N_8790,N_8599);
or UO_1193 (O_1193,N_9410,N_9507);
or UO_1194 (O_1194,N_9203,N_8469);
nand UO_1195 (O_1195,N_8879,N_9657);
nor UO_1196 (O_1196,N_9531,N_9937);
nand UO_1197 (O_1197,N_9856,N_8537);
nor UO_1198 (O_1198,N_9271,N_8447);
or UO_1199 (O_1199,N_8377,N_8067);
or UO_1200 (O_1200,N_9658,N_9804);
nor UO_1201 (O_1201,N_8336,N_9938);
or UO_1202 (O_1202,N_9072,N_8147);
or UO_1203 (O_1203,N_8619,N_8283);
nor UO_1204 (O_1204,N_8295,N_9022);
and UO_1205 (O_1205,N_9422,N_8172);
nand UO_1206 (O_1206,N_9280,N_9547);
or UO_1207 (O_1207,N_8983,N_8019);
or UO_1208 (O_1208,N_8340,N_9524);
nand UO_1209 (O_1209,N_8888,N_9642);
nor UO_1210 (O_1210,N_8537,N_8586);
or UO_1211 (O_1211,N_9819,N_8370);
nor UO_1212 (O_1212,N_8893,N_8871);
nand UO_1213 (O_1213,N_9971,N_8777);
and UO_1214 (O_1214,N_9844,N_9159);
nand UO_1215 (O_1215,N_8447,N_8259);
or UO_1216 (O_1216,N_8871,N_9651);
nor UO_1217 (O_1217,N_9858,N_8917);
or UO_1218 (O_1218,N_8515,N_8826);
and UO_1219 (O_1219,N_8248,N_9375);
and UO_1220 (O_1220,N_8074,N_9737);
nand UO_1221 (O_1221,N_8059,N_8238);
or UO_1222 (O_1222,N_8044,N_8586);
nor UO_1223 (O_1223,N_8121,N_9835);
nor UO_1224 (O_1224,N_8147,N_9028);
or UO_1225 (O_1225,N_8121,N_8696);
or UO_1226 (O_1226,N_8909,N_9145);
nor UO_1227 (O_1227,N_8605,N_8547);
nor UO_1228 (O_1228,N_9757,N_8539);
or UO_1229 (O_1229,N_9454,N_8263);
and UO_1230 (O_1230,N_9188,N_9179);
nand UO_1231 (O_1231,N_8512,N_8469);
or UO_1232 (O_1232,N_9656,N_9767);
and UO_1233 (O_1233,N_8419,N_8938);
nor UO_1234 (O_1234,N_8830,N_8607);
and UO_1235 (O_1235,N_9611,N_8444);
nor UO_1236 (O_1236,N_8185,N_8506);
or UO_1237 (O_1237,N_8087,N_8733);
nand UO_1238 (O_1238,N_9259,N_9562);
and UO_1239 (O_1239,N_9409,N_8545);
or UO_1240 (O_1240,N_9005,N_9879);
and UO_1241 (O_1241,N_9564,N_8512);
and UO_1242 (O_1242,N_9882,N_8346);
and UO_1243 (O_1243,N_8776,N_8351);
and UO_1244 (O_1244,N_9546,N_9092);
nor UO_1245 (O_1245,N_8705,N_8741);
nor UO_1246 (O_1246,N_8511,N_8937);
or UO_1247 (O_1247,N_8679,N_8715);
and UO_1248 (O_1248,N_8053,N_8288);
nor UO_1249 (O_1249,N_8847,N_9178);
nor UO_1250 (O_1250,N_9640,N_8036);
nor UO_1251 (O_1251,N_9193,N_8690);
nand UO_1252 (O_1252,N_8546,N_8650);
nand UO_1253 (O_1253,N_9044,N_9370);
or UO_1254 (O_1254,N_8856,N_8415);
nor UO_1255 (O_1255,N_9988,N_8016);
and UO_1256 (O_1256,N_8064,N_8088);
or UO_1257 (O_1257,N_9341,N_8871);
or UO_1258 (O_1258,N_9163,N_8275);
or UO_1259 (O_1259,N_8578,N_8439);
nor UO_1260 (O_1260,N_8630,N_8105);
nor UO_1261 (O_1261,N_8144,N_8686);
nor UO_1262 (O_1262,N_9819,N_8760);
or UO_1263 (O_1263,N_8745,N_8986);
or UO_1264 (O_1264,N_9488,N_8304);
or UO_1265 (O_1265,N_8708,N_8661);
nor UO_1266 (O_1266,N_8849,N_9760);
nor UO_1267 (O_1267,N_9752,N_8914);
nor UO_1268 (O_1268,N_9363,N_9811);
and UO_1269 (O_1269,N_8662,N_9098);
nor UO_1270 (O_1270,N_9223,N_8953);
nand UO_1271 (O_1271,N_8492,N_8477);
or UO_1272 (O_1272,N_8415,N_8008);
nand UO_1273 (O_1273,N_8303,N_9901);
and UO_1274 (O_1274,N_8589,N_9276);
nand UO_1275 (O_1275,N_8621,N_9445);
nand UO_1276 (O_1276,N_9856,N_8827);
nor UO_1277 (O_1277,N_8250,N_8468);
and UO_1278 (O_1278,N_9153,N_9161);
or UO_1279 (O_1279,N_9024,N_9941);
nand UO_1280 (O_1280,N_9077,N_8828);
nor UO_1281 (O_1281,N_9063,N_8773);
nor UO_1282 (O_1282,N_8879,N_8464);
nand UO_1283 (O_1283,N_8748,N_8573);
or UO_1284 (O_1284,N_9225,N_8381);
nand UO_1285 (O_1285,N_9766,N_8640);
nor UO_1286 (O_1286,N_9462,N_8691);
and UO_1287 (O_1287,N_8961,N_8387);
or UO_1288 (O_1288,N_9121,N_8843);
nor UO_1289 (O_1289,N_8968,N_8501);
and UO_1290 (O_1290,N_9966,N_9913);
nor UO_1291 (O_1291,N_9672,N_9284);
nand UO_1292 (O_1292,N_9726,N_8887);
and UO_1293 (O_1293,N_9562,N_8887);
nand UO_1294 (O_1294,N_9162,N_9822);
and UO_1295 (O_1295,N_8565,N_9125);
nor UO_1296 (O_1296,N_9085,N_8857);
nand UO_1297 (O_1297,N_9001,N_8837);
nand UO_1298 (O_1298,N_8507,N_8946);
nand UO_1299 (O_1299,N_9211,N_8933);
or UO_1300 (O_1300,N_9245,N_8320);
nor UO_1301 (O_1301,N_9858,N_9865);
nand UO_1302 (O_1302,N_9340,N_9676);
and UO_1303 (O_1303,N_8471,N_8495);
nand UO_1304 (O_1304,N_9843,N_8558);
nand UO_1305 (O_1305,N_9013,N_8955);
and UO_1306 (O_1306,N_8037,N_9219);
or UO_1307 (O_1307,N_9842,N_9757);
or UO_1308 (O_1308,N_8208,N_8398);
or UO_1309 (O_1309,N_8371,N_8761);
and UO_1310 (O_1310,N_8387,N_8653);
nor UO_1311 (O_1311,N_9218,N_9648);
and UO_1312 (O_1312,N_8193,N_8869);
nand UO_1313 (O_1313,N_8994,N_9443);
nand UO_1314 (O_1314,N_9898,N_9981);
nor UO_1315 (O_1315,N_9335,N_9631);
or UO_1316 (O_1316,N_9850,N_8195);
nand UO_1317 (O_1317,N_8000,N_9873);
nand UO_1318 (O_1318,N_8216,N_8006);
nand UO_1319 (O_1319,N_9246,N_8452);
nor UO_1320 (O_1320,N_8218,N_9028);
nor UO_1321 (O_1321,N_9389,N_8633);
nand UO_1322 (O_1322,N_8803,N_9988);
and UO_1323 (O_1323,N_8057,N_9287);
or UO_1324 (O_1324,N_8329,N_9799);
nand UO_1325 (O_1325,N_8399,N_9934);
nor UO_1326 (O_1326,N_9440,N_8734);
and UO_1327 (O_1327,N_9801,N_8088);
and UO_1328 (O_1328,N_9976,N_8492);
or UO_1329 (O_1329,N_8554,N_9744);
or UO_1330 (O_1330,N_9497,N_8671);
and UO_1331 (O_1331,N_8649,N_9155);
nand UO_1332 (O_1332,N_9592,N_8221);
or UO_1333 (O_1333,N_9287,N_9514);
and UO_1334 (O_1334,N_8990,N_8686);
nand UO_1335 (O_1335,N_8152,N_8132);
and UO_1336 (O_1336,N_8296,N_8196);
and UO_1337 (O_1337,N_8170,N_9653);
and UO_1338 (O_1338,N_8829,N_8456);
or UO_1339 (O_1339,N_9625,N_9916);
nor UO_1340 (O_1340,N_8635,N_8383);
nand UO_1341 (O_1341,N_9543,N_9269);
and UO_1342 (O_1342,N_8959,N_9018);
and UO_1343 (O_1343,N_8802,N_8260);
or UO_1344 (O_1344,N_8074,N_8832);
or UO_1345 (O_1345,N_9279,N_8286);
nor UO_1346 (O_1346,N_9980,N_8415);
nor UO_1347 (O_1347,N_8656,N_9768);
nor UO_1348 (O_1348,N_9253,N_9604);
and UO_1349 (O_1349,N_8394,N_8709);
nor UO_1350 (O_1350,N_8670,N_9097);
nand UO_1351 (O_1351,N_8714,N_9859);
nand UO_1352 (O_1352,N_8767,N_8043);
or UO_1353 (O_1353,N_9185,N_9187);
nor UO_1354 (O_1354,N_9337,N_9134);
nor UO_1355 (O_1355,N_9701,N_9525);
nand UO_1356 (O_1356,N_9532,N_8403);
and UO_1357 (O_1357,N_9834,N_8469);
or UO_1358 (O_1358,N_9289,N_9935);
and UO_1359 (O_1359,N_9182,N_9389);
xnor UO_1360 (O_1360,N_8403,N_8660);
nor UO_1361 (O_1361,N_9598,N_9774);
nor UO_1362 (O_1362,N_9024,N_9398);
and UO_1363 (O_1363,N_8417,N_8360);
nor UO_1364 (O_1364,N_9847,N_8329);
or UO_1365 (O_1365,N_8382,N_9872);
nand UO_1366 (O_1366,N_9761,N_9023);
nand UO_1367 (O_1367,N_9324,N_9339);
nor UO_1368 (O_1368,N_8449,N_8465);
and UO_1369 (O_1369,N_9592,N_9492);
nand UO_1370 (O_1370,N_9771,N_8294);
or UO_1371 (O_1371,N_8048,N_8689);
or UO_1372 (O_1372,N_9657,N_8631);
and UO_1373 (O_1373,N_8227,N_8313);
or UO_1374 (O_1374,N_9009,N_8629);
nand UO_1375 (O_1375,N_9174,N_9594);
or UO_1376 (O_1376,N_9627,N_9284);
and UO_1377 (O_1377,N_9136,N_9284);
and UO_1378 (O_1378,N_8091,N_8444);
or UO_1379 (O_1379,N_9887,N_8510);
nand UO_1380 (O_1380,N_8721,N_9527);
or UO_1381 (O_1381,N_8311,N_8655);
nand UO_1382 (O_1382,N_8998,N_9291);
and UO_1383 (O_1383,N_8173,N_8805);
or UO_1384 (O_1384,N_8369,N_9989);
nor UO_1385 (O_1385,N_8173,N_9614);
or UO_1386 (O_1386,N_8058,N_9963);
or UO_1387 (O_1387,N_9960,N_9617);
and UO_1388 (O_1388,N_9259,N_8472);
nand UO_1389 (O_1389,N_8890,N_8909);
and UO_1390 (O_1390,N_9448,N_9953);
or UO_1391 (O_1391,N_8580,N_9142);
nand UO_1392 (O_1392,N_8272,N_8454);
and UO_1393 (O_1393,N_9276,N_8164);
nand UO_1394 (O_1394,N_9270,N_8444);
nand UO_1395 (O_1395,N_9164,N_8487);
nor UO_1396 (O_1396,N_8196,N_9810);
nor UO_1397 (O_1397,N_8686,N_8403);
and UO_1398 (O_1398,N_9419,N_9813);
or UO_1399 (O_1399,N_8898,N_9713);
or UO_1400 (O_1400,N_8635,N_8909);
and UO_1401 (O_1401,N_9257,N_8174);
nand UO_1402 (O_1402,N_9511,N_9479);
nand UO_1403 (O_1403,N_8488,N_8412);
or UO_1404 (O_1404,N_8011,N_8863);
and UO_1405 (O_1405,N_9842,N_8438);
nand UO_1406 (O_1406,N_9354,N_9110);
nand UO_1407 (O_1407,N_9652,N_8991);
nand UO_1408 (O_1408,N_9344,N_8641);
nand UO_1409 (O_1409,N_9747,N_9667);
and UO_1410 (O_1410,N_8777,N_8383);
nand UO_1411 (O_1411,N_8460,N_9019);
or UO_1412 (O_1412,N_8119,N_9143);
or UO_1413 (O_1413,N_9623,N_8522);
or UO_1414 (O_1414,N_8446,N_8668);
nand UO_1415 (O_1415,N_8479,N_9006);
nand UO_1416 (O_1416,N_8759,N_8703);
nor UO_1417 (O_1417,N_8215,N_9936);
or UO_1418 (O_1418,N_9968,N_8835);
nor UO_1419 (O_1419,N_8003,N_9098);
nor UO_1420 (O_1420,N_8761,N_9740);
and UO_1421 (O_1421,N_9882,N_9978);
nor UO_1422 (O_1422,N_9039,N_9640);
nand UO_1423 (O_1423,N_8200,N_9683);
nand UO_1424 (O_1424,N_9415,N_8142);
or UO_1425 (O_1425,N_8125,N_9359);
nand UO_1426 (O_1426,N_8514,N_9184);
or UO_1427 (O_1427,N_8080,N_8347);
nor UO_1428 (O_1428,N_8855,N_9121);
or UO_1429 (O_1429,N_8971,N_8229);
or UO_1430 (O_1430,N_9520,N_9597);
nor UO_1431 (O_1431,N_9789,N_8051);
nand UO_1432 (O_1432,N_8662,N_8493);
or UO_1433 (O_1433,N_8875,N_9229);
nor UO_1434 (O_1434,N_9768,N_8930);
nor UO_1435 (O_1435,N_9288,N_9714);
nor UO_1436 (O_1436,N_8850,N_9502);
and UO_1437 (O_1437,N_8222,N_8757);
nand UO_1438 (O_1438,N_8085,N_9106);
and UO_1439 (O_1439,N_9535,N_8570);
or UO_1440 (O_1440,N_8179,N_8637);
and UO_1441 (O_1441,N_8377,N_8931);
nand UO_1442 (O_1442,N_9988,N_9170);
nand UO_1443 (O_1443,N_9047,N_8447);
and UO_1444 (O_1444,N_9077,N_8789);
and UO_1445 (O_1445,N_8573,N_8420);
nor UO_1446 (O_1446,N_8025,N_9047);
or UO_1447 (O_1447,N_8137,N_9126);
nand UO_1448 (O_1448,N_9395,N_8210);
nor UO_1449 (O_1449,N_9001,N_8031);
nor UO_1450 (O_1450,N_8499,N_8515);
and UO_1451 (O_1451,N_9998,N_9685);
xor UO_1452 (O_1452,N_9769,N_8226);
and UO_1453 (O_1453,N_9799,N_9779);
nor UO_1454 (O_1454,N_9192,N_8593);
nor UO_1455 (O_1455,N_8105,N_8872);
or UO_1456 (O_1456,N_8908,N_9136);
nand UO_1457 (O_1457,N_8816,N_9513);
or UO_1458 (O_1458,N_8715,N_9128);
nand UO_1459 (O_1459,N_9837,N_9396);
nand UO_1460 (O_1460,N_8860,N_8293);
nor UO_1461 (O_1461,N_9205,N_9160);
nand UO_1462 (O_1462,N_9535,N_8189);
and UO_1463 (O_1463,N_9593,N_8269);
xnor UO_1464 (O_1464,N_9653,N_9189);
or UO_1465 (O_1465,N_8181,N_9068);
nor UO_1466 (O_1466,N_9342,N_9897);
nand UO_1467 (O_1467,N_9720,N_8667);
or UO_1468 (O_1468,N_8660,N_8406);
nand UO_1469 (O_1469,N_8570,N_8643);
or UO_1470 (O_1470,N_9697,N_8146);
xnor UO_1471 (O_1471,N_9468,N_8299);
nand UO_1472 (O_1472,N_8755,N_9645);
and UO_1473 (O_1473,N_9360,N_8540);
nand UO_1474 (O_1474,N_8520,N_8647);
or UO_1475 (O_1475,N_8698,N_9207);
nand UO_1476 (O_1476,N_9647,N_8418);
nor UO_1477 (O_1477,N_9790,N_8386);
nor UO_1478 (O_1478,N_9222,N_9418);
or UO_1479 (O_1479,N_8531,N_8987);
nand UO_1480 (O_1480,N_8812,N_8490);
nand UO_1481 (O_1481,N_9454,N_9488);
and UO_1482 (O_1482,N_8938,N_8105);
or UO_1483 (O_1483,N_9414,N_9178);
nor UO_1484 (O_1484,N_8797,N_9773);
or UO_1485 (O_1485,N_9206,N_8350);
nand UO_1486 (O_1486,N_8821,N_8692);
and UO_1487 (O_1487,N_9554,N_9423);
and UO_1488 (O_1488,N_8666,N_8244);
nand UO_1489 (O_1489,N_9236,N_8103);
and UO_1490 (O_1490,N_9546,N_8477);
or UO_1491 (O_1491,N_9687,N_9311);
nor UO_1492 (O_1492,N_9408,N_9584);
or UO_1493 (O_1493,N_8571,N_9623);
nor UO_1494 (O_1494,N_9176,N_9604);
and UO_1495 (O_1495,N_9631,N_8574);
or UO_1496 (O_1496,N_9697,N_8046);
nor UO_1497 (O_1497,N_8420,N_8803);
nand UO_1498 (O_1498,N_8832,N_8892);
nand UO_1499 (O_1499,N_8366,N_9279);
endmodule