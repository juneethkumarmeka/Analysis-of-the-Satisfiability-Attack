module basic_1000_10000_1500_2_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5004,N_5005,N_5007,N_5010,N_5011,N_5014,N_5015,N_5018,N_5019,N_5020,N_5025,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5038,N_5043,N_5044,N_5045,N_5046,N_5050,N_5051,N_5054,N_5055,N_5057,N_5058,N_5059,N_5060,N_5061,N_5067,N_5069,N_5070,N_5073,N_5074,N_5075,N_5076,N_5077,N_5080,N_5081,N_5082,N_5088,N_5089,N_5090,N_5092,N_5093,N_5094,N_5095,N_5096,N_5098,N_5099,N_5101,N_5102,N_5103,N_5104,N_5105,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5114,N_5116,N_5117,N_5121,N_5122,N_5123,N_5125,N_5126,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5139,N_5140,N_5141,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5152,N_5156,N_5159,N_5160,N_5162,N_5163,N_5164,N_5168,N_5169,N_5171,N_5172,N_5175,N_5176,N_5177,N_5178,N_5180,N_5181,N_5184,N_5186,N_5188,N_5189,N_5190,N_5191,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5202,N_5203,N_5204,N_5206,N_5208,N_5209,N_5213,N_5215,N_5216,N_5219,N_5220,N_5222,N_5224,N_5227,N_5229,N_5231,N_5232,N_5233,N_5234,N_5236,N_5237,N_5239,N_5240,N_5248,N_5249,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5260,N_5262,N_5264,N_5265,N_5266,N_5267,N_5269,N_5270,N_5274,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5283,N_5286,N_5289,N_5290,N_5291,N_5292,N_5294,N_5296,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5310,N_5311,N_5312,N_5313,N_5314,N_5316,N_5317,N_5319,N_5323,N_5326,N_5329,N_5330,N_5331,N_5332,N_5335,N_5336,N_5337,N_5339,N_5342,N_5343,N_5344,N_5346,N_5347,N_5348,N_5349,N_5351,N_5352,N_5353,N_5354,N_5355,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5366,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5375,N_5377,N_5379,N_5380,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5392,N_5393,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5404,N_5405,N_5406,N_5409,N_5410,N_5413,N_5414,N_5415,N_5417,N_5419,N_5420,N_5421,N_5422,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5435,N_5436,N_5437,N_5438,N_5440,N_5442,N_5443,N_5445,N_5447,N_5450,N_5452,N_5454,N_5456,N_5458,N_5459,N_5461,N_5462,N_5463,N_5465,N_5467,N_5468,N_5469,N_5472,N_5474,N_5475,N_5476,N_5478,N_5479,N_5480,N_5481,N_5482,N_5484,N_5487,N_5488,N_5490,N_5494,N_5496,N_5499,N_5500,N_5504,N_5506,N_5507,N_5508,N_5509,N_5511,N_5512,N_5513,N_5514,N_5516,N_5519,N_5520,N_5521,N_5522,N_5524,N_5525,N_5526,N_5528,N_5529,N_5530,N_5534,N_5536,N_5537,N_5538,N_5541,N_5542,N_5546,N_5548,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5561,N_5562,N_5564,N_5565,N_5566,N_5567,N_5569,N_5570,N_5571,N_5574,N_5579,N_5580,N_5581,N_5583,N_5584,N_5586,N_5587,N_5589,N_5590,N_5592,N_5603,N_5605,N_5606,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5615,N_5617,N_5618,N_5619,N_5621,N_5623,N_5624,N_5625,N_5626,N_5628,N_5629,N_5631,N_5634,N_5635,N_5637,N_5638,N_5639,N_5641,N_5642,N_5644,N_5645,N_5646,N_5647,N_5651,N_5652,N_5658,N_5659,N_5661,N_5662,N_5663,N_5664,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5677,N_5678,N_5681,N_5682,N_5686,N_5687,N_5688,N_5691,N_5693,N_5694,N_5695,N_5696,N_5699,N_5701,N_5704,N_5705,N_5706,N_5709,N_5710,N_5712,N_5713,N_5715,N_5716,N_5717,N_5718,N_5719,N_5721,N_5722,N_5723,N_5725,N_5726,N_5728,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5740,N_5741,N_5744,N_5746,N_5747,N_5748,N_5751,N_5752,N_5753,N_5755,N_5757,N_5758,N_5762,N_5763,N_5764,N_5768,N_5771,N_5772,N_5773,N_5774,N_5775,N_5780,N_5784,N_5785,N_5787,N_5788,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5800,N_5801,N_5803,N_5805,N_5808,N_5811,N_5812,N_5815,N_5818,N_5819,N_5821,N_5823,N_5825,N_5826,N_5827,N_5829,N_5830,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5840,N_5841,N_5842,N_5843,N_5846,N_5847,N_5850,N_5851,N_5853,N_5854,N_5855,N_5857,N_5859,N_5860,N_5864,N_5865,N_5866,N_5867,N_5874,N_5877,N_5878,N_5883,N_5884,N_5885,N_5887,N_5889,N_5891,N_5892,N_5894,N_5896,N_5897,N_5898,N_5902,N_5903,N_5905,N_5907,N_5908,N_5909,N_5911,N_5912,N_5916,N_5918,N_5923,N_5925,N_5926,N_5927,N_5929,N_5930,N_5932,N_5933,N_5934,N_5935,N_5938,N_5943,N_5945,N_5947,N_5949,N_5950,N_5951,N_5952,N_5954,N_5955,N_5956,N_5958,N_5960,N_5962,N_5965,N_5968,N_5970,N_5971,N_5974,N_5975,N_5977,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5994,N_5995,N_5996,N_5997,N_5999,N_6000,N_6001,N_6002,N_6003,N_6005,N_6006,N_6008,N_6009,N_6010,N_6012,N_6014,N_6015,N_6017,N_6018,N_6019,N_6021,N_6022,N_6024,N_6025,N_6026,N_6028,N_6032,N_6036,N_6037,N_6038,N_6039,N_6042,N_6043,N_6044,N_6047,N_6048,N_6050,N_6051,N_6052,N_6055,N_6057,N_6058,N_6066,N_6067,N_6068,N_6069,N_6070,N_6073,N_6074,N_6076,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6095,N_6096,N_6097,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6108,N_6111,N_6115,N_6117,N_6118,N_6119,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6131,N_6132,N_6133,N_6137,N_6138,N_6139,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6150,N_6151,N_6152,N_6153,N_6157,N_6159,N_6161,N_6163,N_6166,N_6167,N_6169,N_6172,N_6174,N_6175,N_6176,N_6180,N_6181,N_6183,N_6184,N_6187,N_6189,N_6190,N_6191,N_6194,N_6195,N_6196,N_6197,N_6198,N_6202,N_6204,N_6205,N_6206,N_6208,N_6209,N_6210,N_6213,N_6215,N_6216,N_6222,N_6223,N_6226,N_6227,N_6230,N_6232,N_6235,N_6236,N_6238,N_6239,N_6240,N_6241,N_6242,N_6245,N_6246,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6256,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6272,N_6276,N_6278,N_6279,N_6284,N_6286,N_6287,N_6289,N_6290,N_6292,N_6293,N_6294,N_6295,N_6297,N_6298,N_6299,N_6300,N_6301,N_6304,N_6305,N_6306,N_6313,N_6314,N_6316,N_6317,N_6320,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6330,N_6333,N_6336,N_6340,N_6341,N_6346,N_6348,N_6349,N_6351,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6366,N_6367,N_6368,N_6370,N_6372,N_6375,N_6376,N_6380,N_6381,N_6384,N_6385,N_6390,N_6394,N_6395,N_6397,N_6398,N_6399,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6412,N_6414,N_6416,N_6418,N_6419,N_6420,N_6422,N_6423,N_6424,N_6425,N_6430,N_6433,N_6434,N_6435,N_6436,N_6439,N_6443,N_6444,N_6446,N_6449,N_6452,N_6454,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6465,N_6466,N_6470,N_6472,N_6473,N_6475,N_6480,N_6481,N_6482,N_6483,N_6484,N_6487,N_6488,N_6489,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6499,N_6500,N_6502,N_6503,N_6504,N_6506,N_6507,N_6508,N_6509,N_6510,N_6512,N_6513,N_6514,N_6516,N_6518,N_6520,N_6522,N_6523,N_6527,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6538,N_6541,N_6542,N_6543,N_6546,N_6547,N_6549,N_6551,N_6553,N_6554,N_6556,N_6558,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6571,N_6577,N_6578,N_6585,N_6588,N_6589,N_6592,N_6594,N_6595,N_6596,N_6597,N_6598,N_6600,N_6601,N_6602,N_6603,N_6606,N_6607,N_6608,N_6609,N_6610,N_6612,N_6616,N_6617,N_6618,N_6620,N_6621,N_6623,N_6624,N_6626,N_6629,N_6630,N_6632,N_6634,N_6635,N_6636,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6646,N_6647,N_6648,N_6649,N_6651,N_6652,N_6653,N_6655,N_6656,N_6658,N_6659,N_6660,N_6661,N_6663,N_6664,N_6665,N_6667,N_6670,N_6671,N_6672,N_6675,N_6676,N_6678,N_6679,N_6684,N_6685,N_6689,N_6691,N_6692,N_6693,N_6694,N_6696,N_6697,N_6698,N_6699,N_6700,N_6702,N_6704,N_6705,N_6706,N_6707,N_6712,N_6717,N_6718,N_6719,N_6720,N_6725,N_6726,N_6727,N_6730,N_6733,N_6734,N_6736,N_6737,N_6739,N_6742,N_6743,N_6744,N_6746,N_6747,N_6748,N_6750,N_6754,N_6756,N_6757,N_6759,N_6760,N_6762,N_6764,N_6765,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6778,N_6779,N_6780,N_6781,N_6783,N_6785,N_6786,N_6787,N_6788,N_6790,N_6791,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6802,N_6803,N_6804,N_6806,N_6808,N_6809,N_6810,N_6813,N_6814,N_6815,N_6816,N_6818,N_6824,N_6826,N_6828,N_6829,N_6830,N_6832,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6843,N_6844,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6853,N_6855,N_6859,N_6860,N_6861,N_6862,N_6863,N_6865,N_6866,N_6867,N_6870,N_6871,N_6873,N_6874,N_6875,N_6877,N_6879,N_6883,N_6885,N_6886,N_6887,N_6888,N_6890,N_6893,N_6895,N_6899,N_6900,N_6901,N_6902,N_6904,N_6905,N_6907,N_6908,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6917,N_6918,N_6919,N_6920,N_6923,N_6924,N_6925,N_6927,N_6929,N_6930,N_6934,N_6935,N_6939,N_6940,N_6941,N_6942,N_6944,N_6948,N_6949,N_6953,N_6954,N_6957,N_6959,N_6960,N_6961,N_6963,N_6966,N_6968,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6978,N_6979,N_6981,N_6982,N_6983,N_6986,N_6987,N_6988,N_6989,N_6991,N_6992,N_6993,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7002,N_7003,N_7006,N_7008,N_7010,N_7011,N_7012,N_7014,N_7015,N_7017,N_7018,N_7021,N_7022,N_7024,N_7025,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7038,N_7042,N_7043,N_7044,N_7045,N_7047,N_7048,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7057,N_7058,N_7059,N_7062,N_7063,N_7064,N_7066,N_7068,N_7070,N_7073,N_7074,N_7076,N_7077,N_7080,N_7083,N_7084,N_7086,N_7087,N_7090,N_7091,N_7092,N_7094,N_7095,N_7096,N_7098,N_7100,N_7103,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7117,N_7118,N_7119,N_7122,N_7124,N_7125,N_7126,N_7127,N_7128,N_7130,N_7131,N_7132,N_7134,N_7135,N_7136,N_7142,N_7144,N_7146,N_7147,N_7148,N_7149,N_7150,N_7153,N_7154,N_7155,N_7156,N_7159,N_7160,N_7162,N_7165,N_7168,N_7171,N_7175,N_7177,N_7178,N_7180,N_7181,N_7182,N_7183,N_7185,N_7187,N_7188,N_7192,N_7193,N_7195,N_7196,N_7201,N_7203,N_7205,N_7206,N_7207,N_7209,N_7210,N_7213,N_7216,N_7217,N_7220,N_7225,N_7226,N_7227,N_7229,N_7230,N_7231,N_7233,N_7235,N_7236,N_7237,N_7238,N_7239,N_7241,N_7242,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7255,N_7256,N_7257,N_7259,N_7260,N_7261,N_7263,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7272,N_7274,N_7276,N_7277,N_7278,N_7282,N_7283,N_7284,N_7287,N_7290,N_7291,N_7292,N_7295,N_7296,N_7299,N_7303,N_7308,N_7312,N_7314,N_7315,N_7316,N_7317,N_7319,N_7320,N_7321,N_7322,N_7324,N_7325,N_7326,N_7327,N_7329,N_7331,N_7334,N_7335,N_7340,N_7342,N_7343,N_7349,N_7351,N_7353,N_7354,N_7355,N_7358,N_7361,N_7362,N_7363,N_7364,N_7366,N_7367,N_7368,N_7369,N_7371,N_7372,N_7373,N_7374,N_7376,N_7377,N_7378,N_7379,N_7381,N_7383,N_7384,N_7385,N_7387,N_7391,N_7392,N_7394,N_7396,N_7398,N_7399,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7408,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7435,N_7438,N_7439,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7448,N_7450,N_7451,N_7453,N_7454,N_7456,N_7457,N_7459,N_7460,N_7462,N_7463,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7476,N_7478,N_7483,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7492,N_7493,N_7494,N_7495,N_7499,N_7502,N_7503,N_7504,N_7505,N_7506,N_7508,N_7509,N_7510,N_7511,N_7514,N_7515,N_7516,N_7518,N_7521,N_7522,N_7525,N_7526,N_7527,N_7531,N_7532,N_7533,N_7534,N_7536,N_7538,N_7540,N_7541,N_7542,N_7543,N_7544,N_7546,N_7548,N_7551,N_7552,N_7554,N_7556,N_7559,N_7560,N_7561,N_7562,N_7564,N_7565,N_7566,N_7568,N_7569,N_7572,N_7573,N_7576,N_7577,N_7580,N_7582,N_7588,N_7589,N_7590,N_7592,N_7596,N_7598,N_7599,N_7600,N_7601,N_7602,N_7605,N_7607,N_7610,N_7612,N_7613,N_7614,N_7616,N_7618,N_7619,N_7622,N_7623,N_7624,N_7625,N_7626,N_7628,N_7629,N_7630,N_7631,N_7634,N_7636,N_7640,N_7641,N_7644,N_7645,N_7646,N_7647,N_7648,N_7650,N_7653,N_7654,N_7655,N_7657,N_7659,N_7667,N_7668,N_7672,N_7673,N_7674,N_7682,N_7683,N_7684,N_7685,N_7687,N_7692,N_7694,N_7697,N_7698,N_7700,N_7701,N_7707,N_7709,N_7710,N_7711,N_7713,N_7714,N_7715,N_7716,N_7718,N_7719,N_7724,N_7725,N_7726,N_7727,N_7729,N_7731,N_7732,N_7734,N_7737,N_7738,N_7740,N_7741,N_7742,N_7743,N_7744,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7758,N_7759,N_7761,N_7763,N_7764,N_7765,N_7769,N_7771,N_7772,N_7773,N_7774,N_7776,N_7777,N_7779,N_7781,N_7783,N_7785,N_7786,N_7787,N_7788,N_7790,N_7794,N_7795,N_7797,N_7799,N_7800,N_7801,N_7803,N_7804,N_7805,N_7807,N_7809,N_7810,N_7811,N_7815,N_7816,N_7817,N_7818,N_7822,N_7825,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7840,N_7844,N_7845,N_7846,N_7847,N_7850,N_7853,N_7854,N_7855,N_7856,N_7857,N_7859,N_7860,N_7861,N_7863,N_7865,N_7867,N_7868,N_7869,N_7871,N_7872,N_7875,N_7876,N_7877,N_7879,N_7880,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7891,N_7892,N_7896,N_7897,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7909,N_7910,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7924,N_7926,N_7928,N_7933,N_7934,N_7935,N_7937,N_7939,N_7940,N_7945,N_7946,N_7947,N_7948,N_7949,N_7952,N_7953,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7964,N_7966,N_7971,N_7976,N_7980,N_7981,N_7984,N_7985,N_7986,N_7987,N_7989,N_7991,N_7992,N_7994,N_7995,N_7996,N_7997,N_7998,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8007,N_8008,N_8011,N_8013,N_8014,N_8017,N_8019,N_8020,N_8023,N_8026,N_8031,N_8033,N_8036,N_8037,N_8038,N_8039,N_8040,N_8042,N_8043,N_8044,N_8047,N_8049,N_8050,N_8054,N_8055,N_8056,N_8057,N_8059,N_8060,N_8061,N_8062,N_8063,N_8066,N_8067,N_8068,N_8069,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8080,N_8081,N_8084,N_8085,N_8086,N_8087,N_8088,N_8090,N_8096,N_8097,N_8101,N_8104,N_8105,N_8107,N_8108,N_8110,N_8113,N_8114,N_8115,N_8116,N_8117,N_8120,N_8123,N_8126,N_8130,N_8131,N_8133,N_8134,N_8135,N_8137,N_8138,N_8140,N_8141,N_8142,N_8143,N_8145,N_8146,N_8149,N_8150,N_8151,N_8152,N_8153,N_8155,N_8157,N_8159,N_8161,N_8162,N_8164,N_8165,N_8166,N_8168,N_8169,N_8171,N_8172,N_8177,N_8179,N_8180,N_8182,N_8183,N_8184,N_8185,N_8189,N_8190,N_8191,N_8194,N_8198,N_8199,N_8200,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8211,N_8213,N_8214,N_8215,N_8223,N_8224,N_8226,N_8227,N_8228,N_8229,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8242,N_8243,N_8244,N_8247,N_8248,N_8249,N_8250,N_8251,N_8254,N_8255,N_8258,N_8260,N_8261,N_8263,N_8264,N_8266,N_8267,N_8269,N_8271,N_8273,N_8275,N_8278,N_8279,N_8280,N_8281,N_8284,N_8286,N_8289,N_8290,N_8291,N_8293,N_8294,N_8295,N_8296,N_8297,N_8301,N_8302,N_8303,N_8305,N_8308,N_8309,N_8310,N_8311,N_8313,N_8316,N_8317,N_8318,N_8319,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8336,N_8337,N_8338,N_8342,N_8343,N_8344,N_8345,N_8346,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8368,N_8370,N_8371,N_8373,N_8374,N_8376,N_8377,N_8379,N_8382,N_8384,N_8385,N_8386,N_8388,N_8389,N_8390,N_8391,N_8394,N_8395,N_8396,N_8397,N_8398,N_8403,N_8404,N_8405,N_8406,N_8407,N_8409,N_8410,N_8413,N_8417,N_8418,N_8419,N_8422,N_8423,N_8424,N_8426,N_8427,N_8430,N_8431,N_8432,N_8433,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8443,N_8444,N_8447,N_8448,N_8449,N_8450,N_8452,N_8453,N_8454,N_8456,N_8457,N_8458,N_8461,N_8462,N_8464,N_8466,N_8467,N_8468,N_8470,N_8471,N_8472,N_8473,N_8476,N_8478,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8489,N_8491,N_8492,N_8494,N_8497,N_8499,N_8501,N_8502,N_8504,N_8505,N_8506,N_8507,N_8510,N_8514,N_8517,N_8519,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8531,N_8533,N_8535,N_8536,N_8537,N_8538,N_8539,N_8542,N_8544,N_8545,N_8546,N_8547,N_8549,N_8551,N_8552,N_8553,N_8556,N_8557,N_8558,N_8561,N_8562,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8571,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8595,N_8598,N_8599,N_8600,N_8604,N_8606,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8618,N_8619,N_8621,N_8622,N_8623,N_8627,N_8629,N_8633,N_8634,N_8635,N_8640,N_8641,N_8642,N_8645,N_8649,N_8651,N_8654,N_8657,N_8658,N_8660,N_8661,N_8664,N_8665,N_8666,N_8670,N_8671,N_8680,N_8683,N_8684,N_8685,N_8687,N_8688,N_8689,N_8690,N_8691,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8709,N_8710,N_8712,N_8714,N_8715,N_8716,N_8718,N_8719,N_8720,N_8722,N_8723,N_8725,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8737,N_8738,N_8740,N_8742,N_8743,N_8744,N_8746,N_8749,N_8751,N_8752,N_8753,N_8754,N_8757,N_8758,N_8761,N_8763,N_8764,N_8765,N_8768,N_8769,N_8771,N_8772,N_8773,N_8774,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8783,N_8786,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8799,N_8800,N_8802,N_8803,N_8804,N_8805,N_8806,N_8808,N_8809,N_8810,N_8811,N_8814,N_8817,N_8818,N_8819,N_8821,N_8823,N_8824,N_8827,N_8828,N_8830,N_8831,N_8833,N_8834,N_8836,N_8837,N_8838,N_8839,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8859,N_8860,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8872,N_8873,N_8875,N_8876,N_8877,N_8878,N_8880,N_8882,N_8883,N_8884,N_8886,N_8887,N_8889,N_8890,N_8893,N_8894,N_8896,N_8897,N_8898,N_8900,N_8902,N_8903,N_8904,N_8905,N_8907,N_8910,N_8911,N_8912,N_8913,N_8914,N_8916,N_8918,N_8919,N_8920,N_8921,N_8922,N_8927,N_8929,N_8930,N_8931,N_8933,N_8934,N_8935,N_8936,N_8938,N_8940,N_8942,N_8943,N_8944,N_8947,N_8948,N_8949,N_8950,N_8952,N_8954,N_8956,N_8957,N_8960,N_8962,N_8964,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8974,N_8976,N_8977,N_8978,N_8979,N_8981,N_8983,N_8984,N_8988,N_8990,N_8991,N_8992,N_8993,N_8994,N_8996,N_8997,N_8998,N_8999,N_9003,N_9006,N_9010,N_9011,N_9013,N_9014,N_9015,N_9016,N_9017,N_9020,N_9022,N_9023,N_9026,N_9028,N_9029,N_9030,N_9032,N_9033,N_9034,N_9035,N_9036,N_9039,N_9040,N_9042,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9055,N_9056,N_9059,N_9062,N_9064,N_9066,N_9069,N_9071,N_9072,N_9073,N_9074,N_9075,N_9078,N_9080,N_9082,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9096,N_9097,N_9099,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9116,N_9117,N_9118,N_9119,N_9121,N_9123,N_9125,N_9129,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9138,N_9143,N_9144,N_9145,N_9147,N_9148,N_9151,N_9153,N_9156,N_9157,N_9159,N_9160,N_9161,N_9162,N_9165,N_9167,N_9169,N_9170,N_9172,N_9173,N_9175,N_9176,N_9177,N_9178,N_9180,N_9181,N_9184,N_9187,N_9189,N_9191,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9213,N_9214,N_9215,N_9216,N_9220,N_9222,N_9223,N_9225,N_9226,N_9228,N_9229,N_9232,N_9233,N_9235,N_9237,N_9238,N_9239,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9250,N_9251,N_9252,N_9254,N_9255,N_9258,N_9259,N_9262,N_9263,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9273,N_9275,N_9277,N_9278,N_9279,N_9280,N_9283,N_9285,N_9286,N_9288,N_9289,N_9290,N_9292,N_9293,N_9297,N_9298,N_9299,N_9300,N_9301,N_9304,N_9305,N_9306,N_9308,N_9309,N_9310,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9322,N_9323,N_9324,N_9326,N_9328,N_9329,N_9333,N_9334,N_9335,N_9337,N_9338,N_9340,N_9341,N_9342,N_9344,N_9346,N_9347,N_9349,N_9351,N_9353,N_9355,N_9356,N_9358,N_9359,N_9361,N_9363,N_9364,N_9365,N_9368,N_9369,N_9371,N_9373,N_9374,N_9375,N_9377,N_9380,N_9381,N_9382,N_9384,N_9385,N_9387,N_9388,N_9390,N_9391,N_9394,N_9395,N_9397,N_9399,N_9400,N_9402,N_9411,N_9412,N_9413,N_9414,N_9415,N_9417,N_9421,N_9423,N_9425,N_9429,N_9430,N_9431,N_9438,N_9439,N_9440,N_9441,N_9443,N_9444,N_9447,N_9448,N_9449,N_9450,N_9451,N_9454,N_9456,N_9457,N_9461,N_9462,N_9464,N_9465,N_9466,N_9473,N_9474,N_9475,N_9478,N_9479,N_9480,N_9484,N_9485,N_9486,N_9492,N_9494,N_9495,N_9500,N_9501,N_9502,N_9504,N_9506,N_9507,N_9508,N_9509,N_9512,N_9513,N_9514,N_9515,N_9517,N_9518,N_9520,N_9521,N_9525,N_9526,N_9527,N_9528,N_9530,N_9531,N_9533,N_9534,N_9535,N_9536,N_9537,N_9540,N_9541,N_9542,N_9543,N_9544,N_9546,N_9547,N_9549,N_9553,N_9554,N_9557,N_9559,N_9562,N_9563,N_9564,N_9566,N_9568,N_9569,N_9571,N_9572,N_9573,N_9576,N_9578,N_9579,N_9580,N_9581,N_9585,N_9588,N_9590,N_9591,N_9592,N_9594,N_9597,N_9599,N_9600,N_9602,N_9605,N_9613,N_9614,N_9616,N_9618,N_9623,N_9624,N_9625,N_9627,N_9630,N_9631,N_9632,N_9635,N_9638,N_9639,N_9640,N_9642,N_9647,N_9648,N_9649,N_9651,N_9653,N_9656,N_9657,N_9659,N_9660,N_9661,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9675,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9689,N_9692,N_9696,N_9699,N_9701,N_9704,N_9705,N_9708,N_9710,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9722,N_9723,N_9724,N_9725,N_9726,N_9728,N_9729,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9742,N_9744,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9754,N_9755,N_9756,N_9758,N_9759,N_9760,N_9761,N_9763,N_9764,N_9767,N_9769,N_9770,N_9772,N_9773,N_9776,N_9777,N_9779,N_9780,N_9782,N_9783,N_9785,N_9786,N_9788,N_9790,N_9791,N_9793,N_9794,N_9795,N_9796,N_9798,N_9800,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9809,N_9810,N_9813,N_9814,N_9816,N_9820,N_9823,N_9824,N_9827,N_9828,N_9829,N_9830,N_9832,N_9833,N_9834,N_9840,N_9847,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9856,N_9857,N_9858,N_9859,N_9860,N_9864,N_9865,N_9866,N_9867,N_9873,N_9874,N_9875,N_9876,N_9879,N_9881,N_9884,N_9888,N_9891,N_9894,N_9895,N_9900,N_9903,N_9904,N_9905,N_9907,N_9909,N_9910,N_9912,N_9913,N_9914,N_9915,N_9916,N_9918,N_9919,N_9920,N_9921,N_9922,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9932,N_9933,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9950,N_9951,N_9952,N_9953,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9965,N_9967,N_9969,N_9970,N_9971,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9995,N_9996,N_9997,N_9998;
nand U0 (N_0,In_327,In_430);
or U1 (N_1,In_410,In_291);
or U2 (N_2,In_446,In_648);
nand U3 (N_3,In_477,In_520);
or U4 (N_4,In_270,In_783);
nand U5 (N_5,In_338,In_813);
nand U6 (N_6,In_998,In_57);
and U7 (N_7,In_618,In_473);
nor U8 (N_8,In_498,In_468);
or U9 (N_9,In_116,In_319);
nand U10 (N_10,In_527,In_476);
or U11 (N_11,In_518,In_119);
and U12 (N_12,In_471,In_662);
nand U13 (N_13,In_21,In_534);
nand U14 (N_14,In_918,In_912);
xor U15 (N_15,In_891,In_395);
nor U16 (N_16,In_986,In_16);
nand U17 (N_17,In_735,In_553);
nor U18 (N_18,In_80,In_386);
nor U19 (N_19,In_834,In_859);
and U20 (N_20,In_968,In_145);
xor U21 (N_21,In_526,In_8);
or U22 (N_22,In_335,In_387);
and U23 (N_23,In_582,In_823);
nor U24 (N_24,In_762,In_447);
or U25 (N_25,In_302,In_159);
or U26 (N_26,In_426,In_257);
nand U27 (N_27,In_598,In_601);
and U28 (N_28,In_744,In_128);
nand U29 (N_29,In_536,In_339);
or U30 (N_30,In_467,In_710);
nand U31 (N_31,In_631,In_826);
nand U32 (N_32,In_723,In_732);
or U33 (N_33,In_658,In_693);
or U34 (N_34,In_221,In_401);
and U35 (N_35,In_572,In_89);
nand U36 (N_36,In_209,In_427);
xnor U37 (N_37,In_558,In_851);
or U38 (N_38,In_576,In_665);
nor U39 (N_39,In_853,In_925);
or U40 (N_40,In_874,In_803);
xor U41 (N_41,In_362,In_179);
or U42 (N_42,In_481,In_231);
nand U43 (N_43,In_168,In_671);
nor U44 (N_44,In_367,In_494);
or U45 (N_45,In_736,In_69);
nand U46 (N_46,In_350,In_624);
nor U47 (N_47,In_899,In_800);
nor U48 (N_48,In_474,In_84);
or U49 (N_49,In_163,In_909);
nand U50 (N_50,In_642,In_81);
nand U51 (N_51,In_269,In_821);
nor U52 (N_52,In_645,In_53);
or U53 (N_53,In_333,In_566);
xor U54 (N_54,In_996,In_40);
xor U55 (N_55,In_931,In_927);
and U56 (N_56,In_411,In_470);
xnor U57 (N_57,In_244,In_465);
or U58 (N_58,In_840,In_997);
and U59 (N_59,In_832,In_186);
or U60 (N_60,In_730,In_196);
nand U61 (N_61,In_118,In_19);
nor U62 (N_62,In_589,In_784);
and U63 (N_63,In_304,In_63);
and U64 (N_64,In_42,In_725);
and U65 (N_65,In_268,In_442);
nand U66 (N_66,In_121,In_6);
nor U67 (N_67,In_884,In_796);
and U68 (N_68,In_361,In_100);
or U69 (N_69,In_58,In_830);
xor U70 (N_70,In_299,In_177);
nor U71 (N_71,In_849,In_46);
xnor U72 (N_72,In_495,In_464);
and U73 (N_73,In_529,In_524);
and U74 (N_74,In_174,In_510);
nor U75 (N_75,In_863,In_633);
or U76 (N_76,In_959,In_842);
nand U77 (N_77,In_415,In_202);
nor U78 (N_78,In_105,In_885);
and U79 (N_79,In_607,In_525);
nor U80 (N_80,In_341,In_551);
xnor U81 (N_81,In_158,In_767);
xor U82 (N_82,In_737,In_413);
nand U83 (N_83,In_363,In_945);
and U84 (N_84,In_808,In_513);
nand U85 (N_85,In_505,In_436);
xnor U86 (N_86,In_332,In_301);
nor U87 (N_87,In_970,In_812);
or U88 (N_88,In_846,In_161);
nor U89 (N_89,In_535,In_691);
xnor U90 (N_90,In_616,In_150);
nor U91 (N_91,In_810,In_560);
xor U92 (N_92,In_903,In_508);
nor U93 (N_93,In_747,In_532);
and U94 (N_94,In_381,In_881);
nor U95 (N_95,In_455,In_711);
nor U96 (N_96,In_342,In_902);
nand U97 (N_97,In_388,In_789);
nor U98 (N_98,In_488,In_435);
or U99 (N_99,In_441,In_194);
or U100 (N_100,In_377,In_462);
and U101 (N_101,In_422,In_277);
xnor U102 (N_102,In_734,In_348);
or U103 (N_103,In_841,In_318);
or U104 (N_104,In_253,In_975);
nor U105 (N_105,In_490,In_234);
nand U106 (N_106,In_233,In_833);
nor U107 (N_107,In_433,In_611);
or U108 (N_108,In_690,In_214);
and U109 (N_109,In_20,In_901);
or U110 (N_110,In_379,In_557);
or U111 (N_111,In_65,In_483);
nand U112 (N_112,In_394,In_236);
nand U113 (N_113,In_983,In_432);
nor U114 (N_114,In_380,In_802);
nand U115 (N_115,In_207,In_317);
xnor U116 (N_116,In_647,In_602);
or U117 (N_117,In_574,In_370);
or U118 (N_118,In_403,In_932);
or U119 (N_119,In_792,In_402);
nor U120 (N_120,In_754,In_795);
nand U121 (N_121,In_870,In_722);
nand U122 (N_122,In_199,In_809);
or U123 (N_123,In_533,In_314);
nand U124 (N_124,In_372,In_219);
nand U125 (N_125,In_967,In_506);
and U126 (N_126,In_858,In_680);
nand U127 (N_127,In_115,In_652);
and U128 (N_128,In_716,In_756);
or U129 (N_129,In_814,In_260);
xor U130 (N_130,In_791,In_59);
and U131 (N_131,In_935,In_964);
nor U132 (N_132,In_130,In_905);
and U133 (N_133,In_603,In_27);
and U134 (N_134,In_7,In_805);
nand U135 (N_135,In_92,In_47);
nor U136 (N_136,In_99,In_570);
or U137 (N_137,In_175,In_843);
xnor U138 (N_138,In_764,In_669);
nand U139 (N_139,In_801,In_522);
xor U140 (N_140,In_530,In_579);
nand U141 (N_141,In_171,In_770);
or U142 (N_142,In_106,In_449);
and U143 (N_143,In_499,In_563);
or U144 (N_144,In_153,In_938);
xor U145 (N_145,In_963,In_571);
xor U146 (N_146,In_897,In_396);
nor U147 (N_147,In_85,In_187);
xnor U148 (N_148,In_608,In_284);
xor U149 (N_149,In_210,In_406);
xor U150 (N_150,In_285,In_896);
nand U151 (N_151,In_156,In_31);
and U152 (N_152,In_599,In_604);
nand U153 (N_153,In_282,In_203);
or U154 (N_154,In_12,In_829);
or U155 (N_155,In_472,In_384);
nor U156 (N_156,In_928,In_879);
nor U157 (N_157,In_475,In_418);
or U158 (N_158,In_686,In_428);
nor U159 (N_159,In_414,In_949);
nand U160 (N_160,In_757,In_519);
and U161 (N_161,In_324,In_714);
or U162 (N_162,In_705,In_531);
and U163 (N_163,In_517,In_160);
nor U164 (N_164,In_248,In_182);
and U165 (N_165,In_399,In_751);
and U166 (N_166,In_544,In_738);
xor U167 (N_167,In_101,In_954);
or U168 (N_168,In_828,In_591);
and U169 (N_169,In_588,In_126);
or U170 (N_170,In_135,In_294);
xor U171 (N_171,In_143,In_555);
nor U172 (N_172,In_868,In_696);
nor U173 (N_173,In_977,In_637);
or U174 (N_174,In_201,In_347);
nand U175 (N_175,In_322,In_698);
nand U176 (N_176,In_96,In_354);
and U177 (N_177,In_771,In_672);
or U178 (N_178,In_674,In_875);
xor U179 (N_179,In_343,In_117);
xnor U180 (N_180,In_35,In_664);
xnor U181 (N_181,In_659,In_458);
nand U182 (N_182,In_729,In_124);
nand U183 (N_183,In_898,In_559);
nand U184 (N_184,In_644,In_369);
nand U185 (N_185,In_971,In_980);
or U186 (N_186,In_981,In_288);
xnor U187 (N_187,In_906,In_818);
nand U188 (N_188,In_144,In_854);
nor U189 (N_189,In_670,In_451);
xnor U190 (N_190,In_457,In_404);
or U191 (N_191,In_765,In_515);
and U192 (N_192,In_62,In_721);
nand U193 (N_193,In_915,In_157);
and U194 (N_194,In_742,In_831);
nor U195 (N_195,In_992,In_249);
nor U196 (N_196,In_61,In_577);
or U197 (N_197,In_390,In_501);
and U198 (N_198,In_929,In_251);
nand U199 (N_199,In_545,In_491);
or U200 (N_200,In_88,In_774);
nand U201 (N_201,In_316,In_781);
nor U202 (N_202,In_438,In_628);
nor U203 (N_203,In_569,In_609);
nand U204 (N_204,In_727,In_425);
nor U205 (N_205,In_523,In_972);
xor U206 (N_206,In_578,In_417);
and U207 (N_207,In_787,In_798);
or U208 (N_208,In_264,In_923);
xor U209 (N_209,In_180,In_646);
nand U210 (N_210,In_140,In_643);
or U211 (N_211,In_552,In_635);
nor U212 (N_212,In_496,In_750);
or U213 (N_213,In_817,In_668);
xnor U214 (N_214,In_336,In_775);
xnor U215 (N_215,In_70,In_663);
nor U216 (N_216,In_108,In_454);
xor U217 (N_217,In_307,In_890);
or U218 (N_218,In_15,In_592);
nand U219 (N_219,In_497,In_739);
xnor U220 (N_220,In_208,In_123);
and U221 (N_221,In_34,In_797);
xor U222 (N_222,In_407,In_786);
xnor U223 (N_223,In_993,In_947);
or U224 (N_224,In_596,In_328);
nor U225 (N_225,In_655,In_590);
or U226 (N_226,In_753,In_25);
and U227 (N_227,In_79,In_340);
and U228 (N_228,In_974,In_279);
nor U229 (N_229,In_91,In_778);
nor U230 (N_230,In_943,In_271);
or U231 (N_231,In_819,In_478);
nand U232 (N_232,In_516,In_661);
and U233 (N_233,In_13,In_703);
or U234 (N_234,In_820,In_865);
xnor U235 (N_235,In_955,In_702);
and U236 (N_236,In_583,In_83);
or U237 (N_237,In_788,In_429);
nor U238 (N_238,In_989,In_305);
and U239 (N_239,In_26,In_749);
or U240 (N_240,In_676,In_373);
nor U241 (N_241,In_740,In_888);
or U242 (N_242,In_839,In_225);
nor U243 (N_243,In_298,In_122);
xor U244 (N_244,In_882,In_112);
nand U245 (N_245,In_987,In_951);
and U246 (N_246,In_872,In_541);
and U247 (N_247,In_585,In_717);
nand U248 (N_248,In_685,In_358);
nor U249 (N_249,In_994,In_678);
or U250 (N_250,In_456,In_266);
nor U251 (N_251,In_877,In_445);
xnor U252 (N_252,In_252,In_807);
nand U253 (N_253,In_707,In_164);
and U254 (N_254,In_60,In_697);
and U255 (N_255,In_237,In_151);
and U256 (N_256,In_656,In_258);
nor U257 (N_257,In_66,In_741);
and U258 (N_258,In_622,In_192);
or U259 (N_259,In_779,In_939);
or U260 (N_260,In_619,In_917);
or U261 (N_261,In_193,In_86);
or U262 (N_262,In_593,In_908);
nand U263 (N_263,In_11,In_82);
nand U264 (N_264,In_554,In_393);
and U265 (N_265,In_567,In_999);
xor U266 (N_266,In_303,In_946);
nand U267 (N_267,In_638,In_170);
nor U268 (N_268,In_706,In_97);
xnor U269 (N_269,In_357,In_485);
or U270 (N_270,In_165,In_836);
nand U271 (N_271,In_982,In_469);
or U272 (N_272,In_930,In_245);
or U273 (N_273,In_45,In_51);
nor U274 (N_274,In_215,In_824);
xor U275 (N_275,In_713,In_924);
nor U276 (N_276,In_374,In_238);
and U277 (N_277,In_804,In_246);
or U278 (N_278,In_408,In_550);
nand U279 (N_279,In_976,In_565);
nand U280 (N_280,In_922,In_920);
or U281 (N_281,In_371,In_845);
and U282 (N_282,In_3,In_136);
xnor U283 (N_283,In_262,In_183);
or U284 (N_284,In_587,In_629);
and U285 (N_285,In_220,In_308);
nor U286 (N_286,In_625,In_376);
nor U287 (N_287,In_883,In_620);
and U288 (N_288,In_806,In_424);
nor U289 (N_289,In_312,In_71);
and U290 (N_290,In_461,In_382);
nand U291 (N_291,In_247,In_852);
nand U292 (N_292,In_235,In_166);
nand U293 (N_293,In_259,In_850);
xor U294 (N_294,In_154,In_597);
nand U295 (N_295,In_724,In_239);
and U296 (N_296,In_562,In_634);
and U297 (N_297,In_914,In_176);
nor U298 (N_298,In_953,In_198);
or U299 (N_299,In_990,In_273);
nand U300 (N_300,In_985,In_759);
nand U301 (N_301,In_934,In_4);
xnor U302 (N_302,In_857,In_32);
and U303 (N_303,In_492,In_521);
xor U304 (N_304,In_397,In_421);
nor U305 (N_305,In_537,In_5);
or U306 (N_306,In_613,In_173);
nor U307 (N_307,In_825,In_866);
and U308 (N_308,In_346,In_17);
xnor U309 (N_309,In_688,In_793);
nand U310 (N_310,In_952,In_37);
nor U311 (N_311,In_300,In_763);
xor U312 (N_312,In_267,In_412);
xor U313 (N_313,In_287,In_848);
and U314 (N_314,In_169,In_480);
or U315 (N_315,In_229,In_1);
and U316 (N_316,In_405,In_600);
and U317 (N_317,In_694,In_704);
nand U318 (N_318,In_549,In_365);
nor U319 (N_319,In_443,In_692);
or U320 (N_320,In_114,In_768);
and U321 (N_321,In_961,In_561);
and U322 (N_322,In_10,In_864);
xnor U323 (N_323,In_984,In_969);
nor U324 (N_324,In_855,In_835);
xor U325 (N_325,In_326,In_761);
xor U326 (N_326,In_958,In_514);
and U327 (N_327,In_211,In_323);
or U328 (N_328,In_460,In_43);
nor U329 (N_329,In_799,In_98);
nor U330 (N_330,In_605,In_580);
nand U331 (N_331,In_223,In_263);
xor U332 (N_332,In_48,In_584);
and U333 (N_333,In_29,In_329);
xor U334 (N_334,In_907,In_904);
xnor U335 (N_335,In_206,In_261);
and U336 (N_336,In_745,In_389);
xnor U337 (N_337,In_218,In_385);
and U338 (N_338,In_683,In_139);
xnor U339 (N_339,In_699,In_679);
nor U340 (N_340,In_448,In_184);
nor U341 (N_341,In_926,In_111);
nor U342 (N_342,In_224,In_213);
xnor U343 (N_343,In_681,In_636);
xnor U344 (N_344,In_73,In_546);
and U345 (N_345,In_639,In_30);
and U346 (N_346,In_102,In_331);
and U347 (N_347,In_718,In_538);
nand U348 (N_348,In_878,In_615);
or U349 (N_349,In_614,In_650);
or U350 (N_350,In_90,In_640);
xnor U351 (N_351,In_419,In_191);
nand U352 (N_352,In_933,In_641);
nor U353 (N_353,In_360,In_701);
xnor U354 (N_354,In_14,In_493);
nor U355 (N_355,In_420,In_568);
nand U356 (N_356,In_889,In_973);
nand U357 (N_357,In_230,In_540);
or U358 (N_358,In_265,In_228);
and U359 (N_359,In_594,In_212);
nand U360 (N_360,In_39,In_507);
nand U361 (N_361,In_275,In_109);
or U362 (N_362,In_965,In_137);
or U363 (N_363,In_423,In_960);
nand U364 (N_364,In_649,In_222);
and U365 (N_365,In_0,In_489);
nor U366 (N_366,In_712,In_28);
xnor U367 (N_367,In_320,In_575);
xnor U368 (N_368,In_666,In_867);
and U369 (N_369,In_673,In_667);
and U370 (N_370,In_979,In_197);
or U371 (N_371,In_780,In_728);
or U372 (N_372,In_232,In_325);
or U373 (N_373,In_172,In_988);
nand U374 (N_374,In_632,In_293);
nor U375 (N_375,In_148,In_450);
xor U376 (N_376,In_147,In_330);
or U377 (N_377,In_309,In_746);
or U378 (N_378,In_398,In_677);
nor U379 (N_379,In_466,In_368);
nor U380 (N_380,In_777,In_966);
and U381 (N_381,In_785,In_916);
xor U382 (N_382,In_827,In_772);
or U383 (N_383,In_189,In_627);
or U384 (N_384,In_311,In_138);
and U385 (N_385,In_621,In_94);
xor U386 (N_386,In_657,In_205);
xor U387 (N_387,In_487,In_286);
nor U388 (N_388,In_543,In_254);
or U389 (N_389,In_142,In_295);
and U390 (N_390,In_416,In_400);
or U391 (N_391,In_995,In_276);
or U392 (N_392,In_250,In_95);
nand U393 (N_393,In_617,In_769);
or U394 (N_394,In_38,In_292);
nor U395 (N_395,In_77,In_104);
nor U396 (N_396,In_272,In_383);
nand U397 (N_397,In_682,In_847);
xnor U398 (N_398,In_913,In_444);
or U399 (N_399,In_861,In_256);
xor U400 (N_400,In_226,In_782);
xnor U401 (N_401,In_2,In_752);
or U402 (N_402,In_586,In_359);
or U403 (N_403,In_900,In_178);
xor U404 (N_404,In_280,In_353);
or U405 (N_405,In_528,In_72);
xnor U406 (N_406,In_152,In_895);
xnor U407 (N_407,In_141,In_107);
xor U408 (N_408,In_131,In_274);
and U409 (N_409,In_310,In_440);
or U410 (N_410,In_651,In_74);
and U411 (N_411,In_500,In_675);
xor U412 (N_412,In_479,In_610);
nand U413 (N_413,In_195,In_950);
and U414 (N_414,In_816,In_719);
or U415 (N_415,In_911,In_313);
and U416 (N_416,In_134,In_720);
or U417 (N_417,In_366,In_281);
nand U418 (N_418,In_630,In_297);
xnor U419 (N_419,In_880,In_794);
nand U420 (N_420,In_146,In_700);
nor U421 (N_421,In_941,In_893);
xnor U422 (N_422,In_9,In_41);
or U423 (N_423,In_217,In_919);
nand U424 (N_424,In_894,In_776);
xor U425 (N_425,In_185,In_944);
nor U426 (N_426,In_283,In_103);
nand U427 (N_427,In_542,In_811);
xor U428 (N_428,In_556,In_684);
nor U429 (N_429,In_155,In_860);
nor U430 (N_430,In_289,In_790);
nand U431 (N_431,In_862,In_871);
nor U432 (N_432,In_547,In_623);
xnor U433 (N_433,In_936,In_942);
xor U434 (N_434,In_509,In_437);
and U435 (N_435,In_743,In_484);
xnor U436 (N_436,In_511,In_937);
xnor U437 (N_437,In_758,In_459);
nor U438 (N_438,In_337,In_708);
nand U439 (N_439,In_75,In_352);
or U440 (N_440,In_50,In_654);
xnor U441 (N_441,In_216,In_23);
and U442 (N_442,In_837,In_344);
and U443 (N_443,In_887,In_760);
or U444 (N_444,In_24,In_54);
nand U445 (N_445,In_453,In_120);
and U446 (N_446,In_87,In_626);
xnor U447 (N_447,In_181,In_773);
nor U448 (N_448,In_242,In_76);
or U449 (N_449,In_876,In_687);
and U450 (N_450,In_956,In_255);
nand U451 (N_451,In_22,In_243);
nand U452 (N_452,In_127,In_240);
and U453 (N_453,In_539,In_67);
xnor U454 (N_454,In_129,In_978);
xor U455 (N_455,In_482,In_355);
nand U456 (N_456,In_110,In_595);
nor U457 (N_457,In_378,In_56);
xor U458 (N_458,In_33,In_715);
xor U459 (N_459,In_726,In_227);
and U460 (N_460,In_113,In_948);
nor U461 (N_461,In_838,In_334);
xnor U462 (N_462,In_606,In_321);
nor U463 (N_463,In_748,In_132);
nor U464 (N_464,In_162,In_52);
or U465 (N_465,In_910,In_815);
nand U466 (N_466,In_125,In_431);
xnor U467 (N_467,In_822,In_660);
nand U468 (N_468,In_349,In_957);
xnor U469 (N_469,In_564,In_204);
and U470 (N_470,In_49,In_869);
xor U471 (N_471,In_731,In_439);
and U472 (N_472,In_612,In_290);
or U473 (N_473,In_296,In_892);
nand U474 (N_474,In_315,In_133);
or U475 (N_475,In_200,In_149);
nor U476 (N_476,In_409,In_962);
nand U477 (N_477,In_503,In_55);
nand U478 (N_478,In_392,In_573);
and U479 (N_479,In_940,In_856);
nand U480 (N_480,In_502,In_653);
and U481 (N_481,In_463,In_512);
and U482 (N_482,In_36,In_64);
and U483 (N_483,In_695,In_921);
nor U484 (N_484,In_733,In_689);
or U485 (N_485,In_356,In_844);
nand U486 (N_486,In_766,In_755);
xor U487 (N_487,In_364,In_504);
nor U488 (N_488,In_44,In_68);
or U489 (N_489,In_78,In_709);
nand U490 (N_490,In_886,In_278);
nand U491 (N_491,In_991,In_375);
xor U492 (N_492,In_452,In_434);
nand U493 (N_493,In_306,In_18);
or U494 (N_494,In_190,In_93);
nand U495 (N_495,In_391,In_188);
xor U496 (N_496,In_351,In_873);
nor U497 (N_497,In_548,In_241);
or U498 (N_498,In_581,In_486);
or U499 (N_499,In_345,In_167);
or U500 (N_500,In_759,In_928);
xnor U501 (N_501,In_222,In_281);
xnor U502 (N_502,In_224,In_193);
xnor U503 (N_503,In_308,In_989);
nor U504 (N_504,In_329,In_939);
and U505 (N_505,In_906,In_980);
xor U506 (N_506,In_459,In_590);
nor U507 (N_507,In_107,In_585);
nor U508 (N_508,In_841,In_245);
xor U509 (N_509,In_120,In_734);
nor U510 (N_510,In_869,In_895);
nand U511 (N_511,In_383,In_616);
nand U512 (N_512,In_868,In_438);
xor U513 (N_513,In_456,In_137);
nor U514 (N_514,In_649,In_850);
nor U515 (N_515,In_827,In_426);
and U516 (N_516,In_109,In_344);
nor U517 (N_517,In_72,In_306);
xnor U518 (N_518,In_274,In_993);
or U519 (N_519,In_241,In_814);
nor U520 (N_520,In_711,In_12);
nor U521 (N_521,In_817,In_868);
xnor U522 (N_522,In_777,In_327);
nor U523 (N_523,In_905,In_532);
xor U524 (N_524,In_370,In_724);
nor U525 (N_525,In_725,In_862);
nand U526 (N_526,In_61,In_124);
xor U527 (N_527,In_97,In_780);
and U528 (N_528,In_618,In_314);
or U529 (N_529,In_406,In_821);
nor U530 (N_530,In_376,In_936);
nand U531 (N_531,In_654,In_734);
nand U532 (N_532,In_711,In_375);
nor U533 (N_533,In_900,In_813);
nor U534 (N_534,In_562,In_584);
nor U535 (N_535,In_469,In_465);
or U536 (N_536,In_935,In_149);
nor U537 (N_537,In_335,In_115);
xor U538 (N_538,In_555,In_33);
or U539 (N_539,In_108,In_994);
and U540 (N_540,In_725,In_496);
nand U541 (N_541,In_206,In_319);
nor U542 (N_542,In_158,In_512);
nand U543 (N_543,In_423,In_415);
nand U544 (N_544,In_680,In_419);
and U545 (N_545,In_798,In_753);
nand U546 (N_546,In_335,In_978);
nand U547 (N_547,In_437,In_841);
nand U548 (N_548,In_352,In_778);
or U549 (N_549,In_711,In_179);
xor U550 (N_550,In_11,In_401);
nand U551 (N_551,In_872,In_212);
and U552 (N_552,In_543,In_36);
or U553 (N_553,In_466,In_415);
nand U554 (N_554,In_597,In_192);
nand U555 (N_555,In_261,In_21);
xor U556 (N_556,In_476,In_669);
and U557 (N_557,In_382,In_190);
or U558 (N_558,In_582,In_829);
nor U559 (N_559,In_488,In_548);
xor U560 (N_560,In_480,In_323);
nand U561 (N_561,In_57,In_368);
or U562 (N_562,In_318,In_503);
or U563 (N_563,In_576,In_736);
and U564 (N_564,In_89,In_946);
nand U565 (N_565,In_308,In_384);
or U566 (N_566,In_860,In_528);
xnor U567 (N_567,In_883,In_69);
and U568 (N_568,In_675,In_55);
nand U569 (N_569,In_281,In_110);
nand U570 (N_570,In_730,In_671);
xor U571 (N_571,In_742,In_116);
nor U572 (N_572,In_953,In_157);
nand U573 (N_573,In_871,In_664);
or U574 (N_574,In_26,In_85);
xor U575 (N_575,In_679,In_437);
or U576 (N_576,In_157,In_556);
or U577 (N_577,In_476,In_491);
or U578 (N_578,In_941,In_105);
or U579 (N_579,In_162,In_425);
or U580 (N_580,In_6,In_73);
nor U581 (N_581,In_84,In_408);
or U582 (N_582,In_972,In_487);
nor U583 (N_583,In_149,In_164);
nand U584 (N_584,In_27,In_826);
nor U585 (N_585,In_601,In_33);
nor U586 (N_586,In_826,In_909);
or U587 (N_587,In_349,In_455);
xnor U588 (N_588,In_947,In_49);
nand U589 (N_589,In_695,In_486);
and U590 (N_590,In_434,In_886);
and U591 (N_591,In_835,In_592);
or U592 (N_592,In_689,In_811);
nand U593 (N_593,In_860,In_38);
xor U594 (N_594,In_259,In_31);
nand U595 (N_595,In_329,In_575);
nand U596 (N_596,In_372,In_300);
or U597 (N_597,In_287,In_595);
xnor U598 (N_598,In_741,In_667);
and U599 (N_599,In_291,In_405);
nor U600 (N_600,In_431,In_561);
nand U601 (N_601,In_275,In_84);
or U602 (N_602,In_100,In_327);
or U603 (N_603,In_573,In_393);
nor U604 (N_604,In_662,In_180);
nand U605 (N_605,In_881,In_7);
xnor U606 (N_606,In_902,In_234);
nand U607 (N_607,In_733,In_434);
nor U608 (N_608,In_478,In_161);
nand U609 (N_609,In_352,In_832);
nor U610 (N_610,In_841,In_303);
nand U611 (N_611,In_365,In_884);
xor U612 (N_612,In_341,In_364);
nand U613 (N_613,In_878,In_18);
and U614 (N_614,In_310,In_869);
nand U615 (N_615,In_774,In_21);
or U616 (N_616,In_31,In_643);
or U617 (N_617,In_155,In_585);
nand U618 (N_618,In_472,In_191);
nor U619 (N_619,In_747,In_902);
and U620 (N_620,In_665,In_447);
and U621 (N_621,In_139,In_137);
nor U622 (N_622,In_39,In_569);
nor U623 (N_623,In_36,In_196);
or U624 (N_624,In_258,In_416);
or U625 (N_625,In_538,In_280);
xnor U626 (N_626,In_47,In_36);
nand U627 (N_627,In_398,In_909);
nand U628 (N_628,In_214,In_592);
or U629 (N_629,In_404,In_367);
or U630 (N_630,In_50,In_230);
nand U631 (N_631,In_65,In_366);
xnor U632 (N_632,In_362,In_402);
and U633 (N_633,In_873,In_960);
xnor U634 (N_634,In_878,In_971);
and U635 (N_635,In_972,In_129);
xnor U636 (N_636,In_571,In_412);
nor U637 (N_637,In_237,In_312);
and U638 (N_638,In_470,In_419);
xnor U639 (N_639,In_826,In_532);
or U640 (N_640,In_396,In_885);
and U641 (N_641,In_965,In_633);
nand U642 (N_642,In_643,In_666);
xor U643 (N_643,In_605,In_802);
or U644 (N_644,In_512,In_452);
xnor U645 (N_645,In_684,In_793);
nor U646 (N_646,In_103,In_753);
nand U647 (N_647,In_961,In_254);
and U648 (N_648,In_320,In_300);
nand U649 (N_649,In_916,In_183);
nor U650 (N_650,In_693,In_447);
nand U651 (N_651,In_691,In_646);
nand U652 (N_652,In_176,In_976);
nand U653 (N_653,In_120,In_381);
xor U654 (N_654,In_236,In_496);
xor U655 (N_655,In_664,In_236);
xnor U656 (N_656,In_95,In_159);
or U657 (N_657,In_85,In_29);
nor U658 (N_658,In_31,In_688);
xnor U659 (N_659,In_527,In_58);
and U660 (N_660,In_668,In_927);
nand U661 (N_661,In_952,In_194);
xor U662 (N_662,In_341,In_282);
nand U663 (N_663,In_546,In_854);
nor U664 (N_664,In_796,In_635);
or U665 (N_665,In_366,In_865);
and U666 (N_666,In_325,In_936);
nand U667 (N_667,In_947,In_432);
and U668 (N_668,In_930,In_975);
nand U669 (N_669,In_106,In_300);
and U670 (N_670,In_585,In_389);
nor U671 (N_671,In_712,In_431);
xnor U672 (N_672,In_979,In_895);
nor U673 (N_673,In_549,In_380);
xnor U674 (N_674,In_393,In_563);
or U675 (N_675,In_920,In_667);
nand U676 (N_676,In_231,In_556);
xor U677 (N_677,In_200,In_379);
xor U678 (N_678,In_541,In_406);
xor U679 (N_679,In_675,In_239);
xor U680 (N_680,In_10,In_495);
nor U681 (N_681,In_160,In_351);
and U682 (N_682,In_241,In_437);
and U683 (N_683,In_630,In_759);
or U684 (N_684,In_569,In_948);
nand U685 (N_685,In_397,In_56);
or U686 (N_686,In_418,In_852);
xor U687 (N_687,In_665,In_800);
or U688 (N_688,In_637,In_125);
nand U689 (N_689,In_650,In_920);
nand U690 (N_690,In_213,In_356);
or U691 (N_691,In_819,In_38);
nand U692 (N_692,In_872,In_684);
and U693 (N_693,In_220,In_876);
and U694 (N_694,In_507,In_416);
nand U695 (N_695,In_695,In_30);
or U696 (N_696,In_901,In_599);
xnor U697 (N_697,In_549,In_201);
nand U698 (N_698,In_995,In_505);
xor U699 (N_699,In_908,In_725);
or U700 (N_700,In_111,In_529);
nor U701 (N_701,In_213,In_148);
xnor U702 (N_702,In_981,In_267);
and U703 (N_703,In_381,In_927);
nor U704 (N_704,In_244,In_983);
or U705 (N_705,In_384,In_893);
and U706 (N_706,In_43,In_486);
xnor U707 (N_707,In_293,In_65);
and U708 (N_708,In_478,In_92);
xnor U709 (N_709,In_318,In_436);
xnor U710 (N_710,In_539,In_385);
xor U711 (N_711,In_765,In_290);
or U712 (N_712,In_71,In_367);
nand U713 (N_713,In_662,In_316);
nand U714 (N_714,In_454,In_56);
and U715 (N_715,In_905,In_164);
or U716 (N_716,In_866,In_649);
xnor U717 (N_717,In_577,In_73);
or U718 (N_718,In_56,In_985);
or U719 (N_719,In_752,In_291);
and U720 (N_720,In_273,In_367);
nand U721 (N_721,In_573,In_300);
and U722 (N_722,In_579,In_932);
nor U723 (N_723,In_733,In_98);
xor U724 (N_724,In_109,In_269);
xnor U725 (N_725,In_259,In_196);
or U726 (N_726,In_308,In_959);
and U727 (N_727,In_651,In_797);
nor U728 (N_728,In_72,In_359);
and U729 (N_729,In_691,In_378);
nor U730 (N_730,In_452,In_94);
nor U731 (N_731,In_255,In_218);
and U732 (N_732,In_85,In_281);
and U733 (N_733,In_63,In_349);
xor U734 (N_734,In_81,In_612);
and U735 (N_735,In_189,In_789);
xnor U736 (N_736,In_820,In_741);
or U737 (N_737,In_865,In_478);
or U738 (N_738,In_933,In_268);
nand U739 (N_739,In_882,In_6);
nand U740 (N_740,In_803,In_839);
and U741 (N_741,In_690,In_753);
or U742 (N_742,In_373,In_767);
or U743 (N_743,In_910,In_445);
xnor U744 (N_744,In_120,In_352);
nor U745 (N_745,In_836,In_691);
nor U746 (N_746,In_916,In_879);
nand U747 (N_747,In_484,In_711);
nor U748 (N_748,In_783,In_17);
nor U749 (N_749,In_434,In_177);
nor U750 (N_750,In_686,In_519);
and U751 (N_751,In_569,In_464);
and U752 (N_752,In_275,In_972);
and U753 (N_753,In_577,In_500);
or U754 (N_754,In_765,In_786);
xor U755 (N_755,In_43,In_541);
nor U756 (N_756,In_767,In_284);
or U757 (N_757,In_520,In_388);
xnor U758 (N_758,In_78,In_388);
nand U759 (N_759,In_4,In_952);
or U760 (N_760,In_300,In_717);
nand U761 (N_761,In_782,In_904);
and U762 (N_762,In_391,In_604);
nand U763 (N_763,In_93,In_551);
and U764 (N_764,In_823,In_975);
nand U765 (N_765,In_986,In_417);
nand U766 (N_766,In_873,In_542);
xor U767 (N_767,In_556,In_51);
or U768 (N_768,In_433,In_159);
and U769 (N_769,In_314,In_792);
and U770 (N_770,In_362,In_164);
and U771 (N_771,In_402,In_319);
and U772 (N_772,In_810,In_222);
nand U773 (N_773,In_797,In_91);
or U774 (N_774,In_338,In_51);
and U775 (N_775,In_386,In_391);
and U776 (N_776,In_349,In_284);
or U777 (N_777,In_523,In_736);
xnor U778 (N_778,In_839,In_899);
xor U779 (N_779,In_298,In_28);
nor U780 (N_780,In_451,In_911);
and U781 (N_781,In_244,In_215);
xor U782 (N_782,In_798,In_519);
nand U783 (N_783,In_511,In_565);
or U784 (N_784,In_218,In_313);
xnor U785 (N_785,In_998,In_202);
and U786 (N_786,In_692,In_169);
or U787 (N_787,In_103,In_536);
nand U788 (N_788,In_22,In_787);
nand U789 (N_789,In_421,In_159);
and U790 (N_790,In_407,In_272);
and U791 (N_791,In_689,In_561);
or U792 (N_792,In_52,In_117);
and U793 (N_793,In_608,In_860);
nand U794 (N_794,In_614,In_768);
xnor U795 (N_795,In_983,In_197);
or U796 (N_796,In_54,In_804);
or U797 (N_797,In_593,In_967);
nor U798 (N_798,In_839,In_811);
and U799 (N_799,In_643,In_337);
and U800 (N_800,In_644,In_68);
nor U801 (N_801,In_363,In_769);
nand U802 (N_802,In_183,In_491);
nor U803 (N_803,In_38,In_326);
xnor U804 (N_804,In_413,In_118);
xnor U805 (N_805,In_404,In_819);
nand U806 (N_806,In_847,In_609);
nor U807 (N_807,In_829,In_486);
xor U808 (N_808,In_701,In_70);
nand U809 (N_809,In_603,In_418);
and U810 (N_810,In_397,In_791);
or U811 (N_811,In_944,In_586);
nand U812 (N_812,In_122,In_763);
xnor U813 (N_813,In_905,In_562);
nand U814 (N_814,In_983,In_913);
nand U815 (N_815,In_203,In_22);
nor U816 (N_816,In_887,In_989);
nor U817 (N_817,In_288,In_274);
and U818 (N_818,In_820,In_963);
nand U819 (N_819,In_519,In_425);
and U820 (N_820,In_108,In_822);
or U821 (N_821,In_549,In_947);
xor U822 (N_822,In_892,In_456);
or U823 (N_823,In_51,In_329);
or U824 (N_824,In_873,In_167);
or U825 (N_825,In_241,In_880);
or U826 (N_826,In_444,In_548);
nand U827 (N_827,In_674,In_266);
nor U828 (N_828,In_887,In_153);
nand U829 (N_829,In_496,In_787);
xor U830 (N_830,In_602,In_486);
and U831 (N_831,In_963,In_565);
nand U832 (N_832,In_433,In_702);
nor U833 (N_833,In_754,In_946);
xor U834 (N_834,In_977,In_168);
nand U835 (N_835,In_14,In_461);
xnor U836 (N_836,In_25,In_15);
nand U837 (N_837,In_427,In_587);
xor U838 (N_838,In_276,In_609);
nor U839 (N_839,In_377,In_214);
and U840 (N_840,In_938,In_166);
and U841 (N_841,In_929,In_41);
nand U842 (N_842,In_419,In_130);
and U843 (N_843,In_1,In_414);
and U844 (N_844,In_484,In_948);
or U845 (N_845,In_943,In_848);
nor U846 (N_846,In_206,In_28);
nand U847 (N_847,In_931,In_855);
nor U848 (N_848,In_196,In_721);
nor U849 (N_849,In_827,In_390);
or U850 (N_850,In_398,In_456);
nand U851 (N_851,In_110,In_698);
xor U852 (N_852,In_543,In_829);
and U853 (N_853,In_54,In_339);
and U854 (N_854,In_78,In_277);
or U855 (N_855,In_439,In_554);
or U856 (N_856,In_438,In_537);
nand U857 (N_857,In_614,In_796);
xor U858 (N_858,In_249,In_863);
or U859 (N_859,In_230,In_256);
nor U860 (N_860,In_398,In_241);
or U861 (N_861,In_5,In_790);
and U862 (N_862,In_410,In_940);
xor U863 (N_863,In_412,In_555);
xor U864 (N_864,In_774,In_229);
xnor U865 (N_865,In_646,In_526);
nor U866 (N_866,In_358,In_939);
xor U867 (N_867,In_127,In_431);
xor U868 (N_868,In_37,In_786);
nor U869 (N_869,In_647,In_469);
xnor U870 (N_870,In_83,In_444);
xor U871 (N_871,In_884,In_594);
nor U872 (N_872,In_689,In_51);
or U873 (N_873,In_828,In_948);
xor U874 (N_874,In_453,In_388);
xnor U875 (N_875,In_442,In_701);
xor U876 (N_876,In_988,In_711);
and U877 (N_877,In_486,In_837);
or U878 (N_878,In_454,In_244);
nor U879 (N_879,In_168,In_492);
xnor U880 (N_880,In_720,In_188);
nor U881 (N_881,In_323,In_580);
or U882 (N_882,In_218,In_181);
xnor U883 (N_883,In_307,In_339);
or U884 (N_884,In_959,In_799);
xnor U885 (N_885,In_281,In_409);
and U886 (N_886,In_557,In_396);
and U887 (N_887,In_304,In_817);
nor U888 (N_888,In_20,In_125);
xor U889 (N_889,In_436,In_736);
nand U890 (N_890,In_766,In_366);
nand U891 (N_891,In_306,In_600);
and U892 (N_892,In_969,In_289);
nor U893 (N_893,In_689,In_910);
nor U894 (N_894,In_147,In_295);
xnor U895 (N_895,In_937,In_494);
xor U896 (N_896,In_886,In_973);
xor U897 (N_897,In_964,In_789);
nor U898 (N_898,In_603,In_376);
xnor U899 (N_899,In_320,In_927);
xor U900 (N_900,In_671,In_95);
or U901 (N_901,In_722,In_573);
xnor U902 (N_902,In_870,In_438);
or U903 (N_903,In_539,In_607);
nand U904 (N_904,In_677,In_984);
xor U905 (N_905,In_708,In_450);
nor U906 (N_906,In_871,In_875);
and U907 (N_907,In_70,In_830);
xor U908 (N_908,In_840,In_363);
and U909 (N_909,In_286,In_485);
or U910 (N_910,In_603,In_266);
and U911 (N_911,In_843,In_209);
xor U912 (N_912,In_770,In_75);
and U913 (N_913,In_461,In_355);
xor U914 (N_914,In_772,In_521);
nand U915 (N_915,In_515,In_128);
nor U916 (N_916,In_130,In_488);
or U917 (N_917,In_837,In_977);
xnor U918 (N_918,In_59,In_700);
nand U919 (N_919,In_958,In_302);
or U920 (N_920,In_845,In_295);
xnor U921 (N_921,In_123,In_352);
nor U922 (N_922,In_365,In_493);
xnor U923 (N_923,In_821,In_884);
xnor U924 (N_924,In_316,In_134);
nand U925 (N_925,In_947,In_510);
xor U926 (N_926,In_542,In_724);
xnor U927 (N_927,In_766,In_58);
and U928 (N_928,In_943,In_739);
xor U929 (N_929,In_324,In_567);
nand U930 (N_930,In_908,In_105);
or U931 (N_931,In_465,In_679);
nor U932 (N_932,In_413,In_249);
nand U933 (N_933,In_537,In_715);
nor U934 (N_934,In_845,In_278);
or U935 (N_935,In_654,In_140);
or U936 (N_936,In_685,In_620);
nand U937 (N_937,In_970,In_798);
or U938 (N_938,In_288,In_324);
nor U939 (N_939,In_630,In_855);
nand U940 (N_940,In_864,In_684);
xnor U941 (N_941,In_456,In_180);
nand U942 (N_942,In_538,In_49);
nor U943 (N_943,In_411,In_194);
xnor U944 (N_944,In_115,In_164);
and U945 (N_945,In_821,In_30);
or U946 (N_946,In_235,In_438);
nor U947 (N_947,In_866,In_501);
nand U948 (N_948,In_353,In_407);
and U949 (N_949,In_547,In_315);
and U950 (N_950,In_817,In_326);
nor U951 (N_951,In_344,In_896);
and U952 (N_952,In_786,In_810);
nor U953 (N_953,In_33,In_589);
nand U954 (N_954,In_617,In_330);
nor U955 (N_955,In_932,In_934);
xor U956 (N_956,In_228,In_430);
nor U957 (N_957,In_252,In_711);
xnor U958 (N_958,In_916,In_896);
nand U959 (N_959,In_774,In_145);
nand U960 (N_960,In_669,In_636);
and U961 (N_961,In_487,In_174);
and U962 (N_962,In_980,In_211);
xnor U963 (N_963,In_89,In_260);
nand U964 (N_964,In_262,In_224);
xnor U965 (N_965,In_523,In_779);
xor U966 (N_966,In_372,In_439);
or U967 (N_967,In_92,In_965);
nor U968 (N_968,In_772,In_717);
xor U969 (N_969,In_87,In_275);
nor U970 (N_970,In_262,In_189);
xnor U971 (N_971,In_119,In_365);
nand U972 (N_972,In_218,In_846);
and U973 (N_973,In_243,In_882);
xor U974 (N_974,In_581,In_323);
xor U975 (N_975,In_43,In_894);
nand U976 (N_976,In_84,In_492);
xnor U977 (N_977,In_937,In_859);
nand U978 (N_978,In_749,In_43);
nor U979 (N_979,In_626,In_63);
xnor U980 (N_980,In_500,In_713);
nand U981 (N_981,In_883,In_520);
or U982 (N_982,In_430,In_748);
or U983 (N_983,In_400,In_456);
nor U984 (N_984,In_96,In_681);
and U985 (N_985,In_950,In_542);
or U986 (N_986,In_667,In_14);
or U987 (N_987,In_875,In_418);
nor U988 (N_988,In_337,In_132);
xor U989 (N_989,In_51,In_629);
or U990 (N_990,In_870,In_96);
xnor U991 (N_991,In_72,In_254);
xnor U992 (N_992,In_745,In_708);
xor U993 (N_993,In_189,In_867);
nand U994 (N_994,In_787,In_87);
nor U995 (N_995,In_430,In_191);
xnor U996 (N_996,In_505,In_401);
xor U997 (N_997,In_748,In_718);
and U998 (N_998,In_135,In_982);
or U999 (N_999,In_78,In_81);
nand U1000 (N_1000,In_862,In_909);
nor U1001 (N_1001,In_945,In_536);
nand U1002 (N_1002,In_515,In_632);
nor U1003 (N_1003,In_782,In_327);
and U1004 (N_1004,In_944,In_758);
nand U1005 (N_1005,In_980,In_593);
xnor U1006 (N_1006,In_111,In_569);
nor U1007 (N_1007,In_913,In_131);
nand U1008 (N_1008,In_788,In_822);
nand U1009 (N_1009,In_59,In_913);
xnor U1010 (N_1010,In_239,In_714);
or U1011 (N_1011,In_474,In_764);
and U1012 (N_1012,In_877,In_742);
xor U1013 (N_1013,In_113,In_463);
or U1014 (N_1014,In_586,In_495);
nand U1015 (N_1015,In_512,In_570);
nand U1016 (N_1016,In_135,In_493);
and U1017 (N_1017,In_487,In_780);
nand U1018 (N_1018,In_841,In_777);
xnor U1019 (N_1019,In_72,In_36);
and U1020 (N_1020,In_640,In_592);
nor U1021 (N_1021,In_449,In_558);
and U1022 (N_1022,In_858,In_640);
and U1023 (N_1023,In_865,In_928);
and U1024 (N_1024,In_721,In_848);
nor U1025 (N_1025,In_174,In_864);
and U1026 (N_1026,In_45,In_581);
and U1027 (N_1027,In_532,In_553);
nor U1028 (N_1028,In_79,In_48);
nand U1029 (N_1029,In_998,In_487);
nand U1030 (N_1030,In_986,In_62);
xnor U1031 (N_1031,In_719,In_84);
and U1032 (N_1032,In_429,In_458);
and U1033 (N_1033,In_407,In_197);
nor U1034 (N_1034,In_499,In_2);
and U1035 (N_1035,In_345,In_993);
and U1036 (N_1036,In_335,In_432);
nand U1037 (N_1037,In_531,In_689);
or U1038 (N_1038,In_703,In_280);
nand U1039 (N_1039,In_56,In_739);
nand U1040 (N_1040,In_536,In_214);
xnor U1041 (N_1041,In_791,In_950);
or U1042 (N_1042,In_960,In_179);
nand U1043 (N_1043,In_592,In_78);
nand U1044 (N_1044,In_27,In_521);
or U1045 (N_1045,In_954,In_294);
or U1046 (N_1046,In_255,In_411);
xor U1047 (N_1047,In_647,In_972);
nor U1048 (N_1048,In_545,In_966);
and U1049 (N_1049,In_200,In_608);
xor U1050 (N_1050,In_11,In_451);
and U1051 (N_1051,In_793,In_891);
nand U1052 (N_1052,In_761,In_247);
and U1053 (N_1053,In_931,In_374);
or U1054 (N_1054,In_434,In_363);
xor U1055 (N_1055,In_950,In_701);
and U1056 (N_1056,In_978,In_536);
nand U1057 (N_1057,In_905,In_689);
and U1058 (N_1058,In_529,In_500);
xnor U1059 (N_1059,In_253,In_795);
nor U1060 (N_1060,In_138,In_871);
xor U1061 (N_1061,In_394,In_175);
or U1062 (N_1062,In_62,In_553);
xnor U1063 (N_1063,In_80,In_65);
or U1064 (N_1064,In_910,In_857);
and U1065 (N_1065,In_767,In_683);
and U1066 (N_1066,In_189,In_830);
nor U1067 (N_1067,In_120,In_973);
and U1068 (N_1068,In_351,In_977);
nor U1069 (N_1069,In_131,In_721);
or U1070 (N_1070,In_819,In_527);
or U1071 (N_1071,In_566,In_697);
nor U1072 (N_1072,In_90,In_25);
xnor U1073 (N_1073,In_407,In_670);
nor U1074 (N_1074,In_689,In_508);
nor U1075 (N_1075,In_762,In_114);
or U1076 (N_1076,In_656,In_999);
or U1077 (N_1077,In_208,In_469);
nand U1078 (N_1078,In_40,In_798);
or U1079 (N_1079,In_419,In_271);
or U1080 (N_1080,In_97,In_215);
nor U1081 (N_1081,In_894,In_189);
nand U1082 (N_1082,In_234,In_127);
nor U1083 (N_1083,In_368,In_292);
xor U1084 (N_1084,In_88,In_259);
and U1085 (N_1085,In_617,In_972);
and U1086 (N_1086,In_606,In_84);
and U1087 (N_1087,In_722,In_709);
xor U1088 (N_1088,In_334,In_857);
or U1089 (N_1089,In_833,In_968);
and U1090 (N_1090,In_954,In_624);
or U1091 (N_1091,In_669,In_814);
nor U1092 (N_1092,In_334,In_289);
nand U1093 (N_1093,In_318,In_240);
nor U1094 (N_1094,In_71,In_256);
nand U1095 (N_1095,In_122,In_511);
or U1096 (N_1096,In_433,In_263);
nor U1097 (N_1097,In_837,In_922);
and U1098 (N_1098,In_190,In_599);
nor U1099 (N_1099,In_122,In_71);
nand U1100 (N_1100,In_847,In_904);
xor U1101 (N_1101,In_720,In_647);
nand U1102 (N_1102,In_524,In_996);
or U1103 (N_1103,In_16,In_848);
nand U1104 (N_1104,In_87,In_991);
xor U1105 (N_1105,In_67,In_413);
nand U1106 (N_1106,In_713,In_157);
nand U1107 (N_1107,In_802,In_303);
nor U1108 (N_1108,In_129,In_232);
or U1109 (N_1109,In_527,In_555);
or U1110 (N_1110,In_947,In_987);
nand U1111 (N_1111,In_613,In_725);
nor U1112 (N_1112,In_648,In_561);
or U1113 (N_1113,In_484,In_399);
nor U1114 (N_1114,In_604,In_551);
nand U1115 (N_1115,In_794,In_434);
nor U1116 (N_1116,In_411,In_189);
or U1117 (N_1117,In_560,In_563);
or U1118 (N_1118,In_409,In_527);
nor U1119 (N_1119,In_219,In_893);
nand U1120 (N_1120,In_915,In_225);
nand U1121 (N_1121,In_486,In_327);
nand U1122 (N_1122,In_809,In_776);
or U1123 (N_1123,In_7,In_204);
xor U1124 (N_1124,In_929,In_850);
nor U1125 (N_1125,In_958,In_641);
nor U1126 (N_1126,In_582,In_662);
and U1127 (N_1127,In_348,In_639);
and U1128 (N_1128,In_771,In_772);
nand U1129 (N_1129,In_287,In_705);
nand U1130 (N_1130,In_83,In_78);
nand U1131 (N_1131,In_63,In_390);
or U1132 (N_1132,In_683,In_695);
or U1133 (N_1133,In_825,In_253);
or U1134 (N_1134,In_282,In_991);
xor U1135 (N_1135,In_100,In_106);
xnor U1136 (N_1136,In_57,In_260);
nor U1137 (N_1137,In_465,In_830);
or U1138 (N_1138,In_514,In_468);
nand U1139 (N_1139,In_440,In_959);
nand U1140 (N_1140,In_627,In_604);
nor U1141 (N_1141,In_467,In_507);
nand U1142 (N_1142,In_591,In_275);
nand U1143 (N_1143,In_278,In_254);
and U1144 (N_1144,In_151,In_766);
and U1145 (N_1145,In_774,In_191);
xor U1146 (N_1146,In_467,In_459);
nand U1147 (N_1147,In_375,In_753);
xor U1148 (N_1148,In_491,In_33);
xor U1149 (N_1149,In_625,In_865);
nand U1150 (N_1150,In_223,In_825);
xnor U1151 (N_1151,In_357,In_159);
and U1152 (N_1152,In_331,In_581);
nand U1153 (N_1153,In_749,In_583);
nand U1154 (N_1154,In_523,In_308);
nor U1155 (N_1155,In_947,In_127);
or U1156 (N_1156,In_334,In_173);
nor U1157 (N_1157,In_781,In_281);
nor U1158 (N_1158,In_331,In_631);
xor U1159 (N_1159,In_564,In_336);
and U1160 (N_1160,In_859,In_719);
and U1161 (N_1161,In_722,In_238);
or U1162 (N_1162,In_819,In_253);
nand U1163 (N_1163,In_972,In_839);
or U1164 (N_1164,In_432,In_7);
and U1165 (N_1165,In_973,In_603);
nand U1166 (N_1166,In_565,In_585);
nand U1167 (N_1167,In_53,In_549);
xnor U1168 (N_1168,In_53,In_715);
nor U1169 (N_1169,In_94,In_169);
and U1170 (N_1170,In_844,In_102);
nor U1171 (N_1171,In_662,In_411);
nand U1172 (N_1172,In_653,In_145);
or U1173 (N_1173,In_757,In_371);
or U1174 (N_1174,In_716,In_58);
nand U1175 (N_1175,In_46,In_213);
and U1176 (N_1176,In_77,In_587);
or U1177 (N_1177,In_647,In_723);
or U1178 (N_1178,In_60,In_354);
nor U1179 (N_1179,In_594,In_3);
nor U1180 (N_1180,In_626,In_886);
xnor U1181 (N_1181,In_752,In_208);
xor U1182 (N_1182,In_587,In_107);
xnor U1183 (N_1183,In_374,In_489);
and U1184 (N_1184,In_392,In_384);
or U1185 (N_1185,In_501,In_74);
and U1186 (N_1186,In_4,In_275);
or U1187 (N_1187,In_645,In_905);
xor U1188 (N_1188,In_396,In_816);
nand U1189 (N_1189,In_132,In_328);
or U1190 (N_1190,In_316,In_216);
xnor U1191 (N_1191,In_628,In_28);
nand U1192 (N_1192,In_227,In_49);
xor U1193 (N_1193,In_816,In_463);
or U1194 (N_1194,In_237,In_38);
or U1195 (N_1195,In_707,In_71);
nor U1196 (N_1196,In_811,In_41);
nand U1197 (N_1197,In_445,In_698);
nor U1198 (N_1198,In_649,In_307);
xor U1199 (N_1199,In_675,In_213);
or U1200 (N_1200,In_737,In_260);
or U1201 (N_1201,In_381,In_580);
xnor U1202 (N_1202,In_926,In_872);
nand U1203 (N_1203,In_724,In_804);
and U1204 (N_1204,In_942,In_120);
nand U1205 (N_1205,In_541,In_635);
nand U1206 (N_1206,In_413,In_583);
or U1207 (N_1207,In_959,In_333);
and U1208 (N_1208,In_390,In_761);
and U1209 (N_1209,In_25,In_732);
xor U1210 (N_1210,In_47,In_538);
nand U1211 (N_1211,In_104,In_817);
nor U1212 (N_1212,In_725,In_729);
nand U1213 (N_1213,In_850,In_50);
nand U1214 (N_1214,In_622,In_120);
xnor U1215 (N_1215,In_809,In_185);
xnor U1216 (N_1216,In_564,In_934);
or U1217 (N_1217,In_587,In_242);
nor U1218 (N_1218,In_301,In_863);
nand U1219 (N_1219,In_489,In_389);
xnor U1220 (N_1220,In_821,In_850);
and U1221 (N_1221,In_139,In_715);
and U1222 (N_1222,In_946,In_387);
nor U1223 (N_1223,In_464,In_769);
xor U1224 (N_1224,In_275,In_631);
xnor U1225 (N_1225,In_907,In_633);
and U1226 (N_1226,In_377,In_491);
nor U1227 (N_1227,In_901,In_400);
xor U1228 (N_1228,In_987,In_591);
nand U1229 (N_1229,In_565,In_66);
xor U1230 (N_1230,In_313,In_30);
nor U1231 (N_1231,In_118,In_916);
nor U1232 (N_1232,In_129,In_254);
nor U1233 (N_1233,In_896,In_15);
xor U1234 (N_1234,In_865,In_164);
or U1235 (N_1235,In_118,In_996);
xnor U1236 (N_1236,In_84,In_637);
xnor U1237 (N_1237,In_492,In_615);
and U1238 (N_1238,In_245,In_98);
nor U1239 (N_1239,In_61,In_482);
or U1240 (N_1240,In_600,In_117);
nand U1241 (N_1241,In_669,In_190);
or U1242 (N_1242,In_818,In_941);
or U1243 (N_1243,In_99,In_154);
nor U1244 (N_1244,In_303,In_220);
nor U1245 (N_1245,In_448,In_406);
nor U1246 (N_1246,In_773,In_880);
and U1247 (N_1247,In_304,In_354);
xnor U1248 (N_1248,In_886,In_112);
xnor U1249 (N_1249,In_224,In_183);
nor U1250 (N_1250,In_684,In_994);
or U1251 (N_1251,In_766,In_32);
and U1252 (N_1252,In_312,In_25);
and U1253 (N_1253,In_202,In_984);
nor U1254 (N_1254,In_211,In_883);
nand U1255 (N_1255,In_252,In_294);
xnor U1256 (N_1256,In_262,In_355);
xor U1257 (N_1257,In_865,In_354);
nor U1258 (N_1258,In_3,In_305);
nand U1259 (N_1259,In_541,In_854);
or U1260 (N_1260,In_90,In_766);
nand U1261 (N_1261,In_166,In_229);
nand U1262 (N_1262,In_779,In_872);
and U1263 (N_1263,In_976,In_428);
nand U1264 (N_1264,In_665,In_560);
or U1265 (N_1265,In_257,In_831);
xor U1266 (N_1266,In_456,In_720);
nor U1267 (N_1267,In_170,In_3);
and U1268 (N_1268,In_680,In_628);
nand U1269 (N_1269,In_133,In_311);
xnor U1270 (N_1270,In_789,In_49);
or U1271 (N_1271,In_277,In_65);
xor U1272 (N_1272,In_251,In_572);
nand U1273 (N_1273,In_516,In_884);
nor U1274 (N_1274,In_481,In_898);
nand U1275 (N_1275,In_931,In_470);
and U1276 (N_1276,In_709,In_822);
nand U1277 (N_1277,In_669,In_467);
nand U1278 (N_1278,In_690,In_383);
xnor U1279 (N_1279,In_129,In_831);
nor U1280 (N_1280,In_198,In_676);
xnor U1281 (N_1281,In_821,In_760);
and U1282 (N_1282,In_107,In_618);
xor U1283 (N_1283,In_591,In_291);
or U1284 (N_1284,In_739,In_721);
and U1285 (N_1285,In_882,In_577);
nand U1286 (N_1286,In_789,In_126);
nor U1287 (N_1287,In_931,In_553);
or U1288 (N_1288,In_871,In_618);
or U1289 (N_1289,In_125,In_445);
xnor U1290 (N_1290,In_326,In_821);
nor U1291 (N_1291,In_643,In_305);
and U1292 (N_1292,In_578,In_997);
xnor U1293 (N_1293,In_491,In_239);
and U1294 (N_1294,In_90,In_308);
or U1295 (N_1295,In_867,In_365);
nand U1296 (N_1296,In_542,In_189);
or U1297 (N_1297,In_666,In_206);
or U1298 (N_1298,In_635,In_857);
nor U1299 (N_1299,In_654,In_361);
or U1300 (N_1300,In_460,In_687);
xnor U1301 (N_1301,In_600,In_110);
and U1302 (N_1302,In_620,In_175);
nor U1303 (N_1303,In_241,In_652);
nand U1304 (N_1304,In_625,In_836);
nor U1305 (N_1305,In_127,In_926);
or U1306 (N_1306,In_237,In_183);
nand U1307 (N_1307,In_31,In_94);
or U1308 (N_1308,In_787,In_676);
nor U1309 (N_1309,In_32,In_416);
xnor U1310 (N_1310,In_406,In_751);
and U1311 (N_1311,In_149,In_904);
and U1312 (N_1312,In_747,In_195);
nand U1313 (N_1313,In_473,In_271);
nand U1314 (N_1314,In_420,In_345);
xnor U1315 (N_1315,In_582,In_583);
or U1316 (N_1316,In_476,In_56);
nor U1317 (N_1317,In_885,In_493);
xor U1318 (N_1318,In_102,In_897);
nand U1319 (N_1319,In_211,In_187);
nand U1320 (N_1320,In_132,In_30);
or U1321 (N_1321,In_337,In_838);
or U1322 (N_1322,In_958,In_207);
or U1323 (N_1323,In_226,In_272);
and U1324 (N_1324,In_284,In_617);
xnor U1325 (N_1325,In_646,In_461);
nor U1326 (N_1326,In_255,In_173);
nor U1327 (N_1327,In_669,In_896);
xnor U1328 (N_1328,In_156,In_804);
nand U1329 (N_1329,In_884,In_236);
nor U1330 (N_1330,In_577,In_890);
xnor U1331 (N_1331,In_344,In_150);
xor U1332 (N_1332,In_162,In_127);
xor U1333 (N_1333,In_833,In_688);
xnor U1334 (N_1334,In_761,In_47);
or U1335 (N_1335,In_146,In_792);
or U1336 (N_1336,In_387,In_369);
or U1337 (N_1337,In_931,In_746);
nor U1338 (N_1338,In_203,In_957);
or U1339 (N_1339,In_860,In_656);
and U1340 (N_1340,In_534,In_540);
xor U1341 (N_1341,In_729,In_971);
nor U1342 (N_1342,In_706,In_269);
nand U1343 (N_1343,In_422,In_36);
nand U1344 (N_1344,In_500,In_755);
or U1345 (N_1345,In_329,In_630);
and U1346 (N_1346,In_619,In_809);
xor U1347 (N_1347,In_499,In_444);
xor U1348 (N_1348,In_884,In_430);
and U1349 (N_1349,In_116,In_461);
nor U1350 (N_1350,In_540,In_111);
and U1351 (N_1351,In_385,In_220);
nand U1352 (N_1352,In_102,In_909);
xor U1353 (N_1353,In_140,In_230);
nand U1354 (N_1354,In_268,In_274);
nor U1355 (N_1355,In_321,In_431);
nor U1356 (N_1356,In_116,In_450);
nor U1357 (N_1357,In_14,In_914);
or U1358 (N_1358,In_805,In_826);
or U1359 (N_1359,In_666,In_58);
nand U1360 (N_1360,In_229,In_183);
xor U1361 (N_1361,In_930,In_721);
and U1362 (N_1362,In_431,In_639);
nand U1363 (N_1363,In_472,In_617);
and U1364 (N_1364,In_324,In_419);
nand U1365 (N_1365,In_122,In_911);
nor U1366 (N_1366,In_483,In_232);
and U1367 (N_1367,In_314,In_896);
and U1368 (N_1368,In_285,In_902);
nor U1369 (N_1369,In_312,In_764);
nand U1370 (N_1370,In_280,In_450);
xor U1371 (N_1371,In_42,In_958);
or U1372 (N_1372,In_369,In_162);
xnor U1373 (N_1373,In_662,In_20);
nand U1374 (N_1374,In_438,In_45);
and U1375 (N_1375,In_553,In_195);
nor U1376 (N_1376,In_153,In_719);
and U1377 (N_1377,In_974,In_1);
xnor U1378 (N_1378,In_658,In_171);
or U1379 (N_1379,In_493,In_195);
nor U1380 (N_1380,In_254,In_299);
nand U1381 (N_1381,In_715,In_330);
and U1382 (N_1382,In_987,In_70);
xor U1383 (N_1383,In_881,In_854);
or U1384 (N_1384,In_612,In_706);
or U1385 (N_1385,In_888,In_996);
nor U1386 (N_1386,In_519,In_308);
xnor U1387 (N_1387,In_623,In_517);
nand U1388 (N_1388,In_767,In_193);
xnor U1389 (N_1389,In_3,In_267);
xnor U1390 (N_1390,In_931,In_852);
xor U1391 (N_1391,In_68,In_543);
and U1392 (N_1392,In_497,In_604);
xnor U1393 (N_1393,In_632,In_603);
or U1394 (N_1394,In_819,In_428);
nor U1395 (N_1395,In_806,In_532);
or U1396 (N_1396,In_178,In_826);
or U1397 (N_1397,In_586,In_499);
or U1398 (N_1398,In_656,In_288);
or U1399 (N_1399,In_614,In_656);
or U1400 (N_1400,In_910,In_863);
xor U1401 (N_1401,In_336,In_921);
and U1402 (N_1402,In_724,In_668);
nand U1403 (N_1403,In_598,In_614);
xnor U1404 (N_1404,In_141,In_275);
nor U1405 (N_1405,In_211,In_421);
or U1406 (N_1406,In_957,In_863);
or U1407 (N_1407,In_526,In_220);
and U1408 (N_1408,In_951,In_625);
or U1409 (N_1409,In_226,In_536);
nor U1410 (N_1410,In_822,In_484);
nand U1411 (N_1411,In_350,In_560);
nand U1412 (N_1412,In_551,In_155);
nor U1413 (N_1413,In_181,In_224);
nor U1414 (N_1414,In_190,In_75);
xnor U1415 (N_1415,In_667,In_838);
or U1416 (N_1416,In_970,In_672);
and U1417 (N_1417,In_507,In_713);
nand U1418 (N_1418,In_152,In_278);
nor U1419 (N_1419,In_483,In_533);
and U1420 (N_1420,In_601,In_814);
or U1421 (N_1421,In_593,In_902);
nor U1422 (N_1422,In_375,In_488);
xnor U1423 (N_1423,In_468,In_563);
nand U1424 (N_1424,In_257,In_439);
and U1425 (N_1425,In_573,In_521);
nor U1426 (N_1426,In_873,In_474);
and U1427 (N_1427,In_540,In_826);
nand U1428 (N_1428,In_614,In_128);
nor U1429 (N_1429,In_258,In_933);
xnor U1430 (N_1430,In_227,In_633);
xor U1431 (N_1431,In_858,In_788);
and U1432 (N_1432,In_969,In_550);
and U1433 (N_1433,In_144,In_515);
nand U1434 (N_1434,In_534,In_564);
and U1435 (N_1435,In_986,In_896);
nor U1436 (N_1436,In_9,In_20);
nor U1437 (N_1437,In_735,In_377);
and U1438 (N_1438,In_201,In_752);
and U1439 (N_1439,In_218,In_947);
and U1440 (N_1440,In_108,In_503);
and U1441 (N_1441,In_705,In_414);
and U1442 (N_1442,In_649,In_445);
or U1443 (N_1443,In_733,In_549);
xnor U1444 (N_1444,In_52,In_6);
and U1445 (N_1445,In_796,In_896);
nand U1446 (N_1446,In_108,In_976);
or U1447 (N_1447,In_832,In_826);
nand U1448 (N_1448,In_202,In_373);
and U1449 (N_1449,In_993,In_691);
nand U1450 (N_1450,In_354,In_444);
and U1451 (N_1451,In_762,In_954);
nor U1452 (N_1452,In_335,In_779);
nor U1453 (N_1453,In_667,In_585);
and U1454 (N_1454,In_410,In_777);
and U1455 (N_1455,In_459,In_765);
or U1456 (N_1456,In_608,In_147);
or U1457 (N_1457,In_5,In_295);
and U1458 (N_1458,In_338,In_86);
nand U1459 (N_1459,In_462,In_906);
nor U1460 (N_1460,In_114,In_726);
nor U1461 (N_1461,In_170,In_332);
nor U1462 (N_1462,In_49,In_75);
or U1463 (N_1463,In_513,In_166);
or U1464 (N_1464,In_995,In_601);
and U1465 (N_1465,In_63,In_498);
or U1466 (N_1466,In_405,In_821);
nand U1467 (N_1467,In_561,In_626);
xor U1468 (N_1468,In_952,In_146);
nor U1469 (N_1469,In_275,In_669);
xor U1470 (N_1470,In_515,In_656);
xor U1471 (N_1471,In_804,In_492);
or U1472 (N_1472,In_829,In_256);
and U1473 (N_1473,In_50,In_342);
nor U1474 (N_1474,In_339,In_738);
xnor U1475 (N_1475,In_128,In_396);
nor U1476 (N_1476,In_553,In_243);
nor U1477 (N_1477,In_642,In_874);
or U1478 (N_1478,In_349,In_10);
and U1479 (N_1479,In_223,In_967);
nor U1480 (N_1480,In_785,In_235);
nor U1481 (N_1481,In_621,In_719);
nor U1482 (N_1482,In_569,In_608);
or U1483 (N_1483,In_11,In_798);
nor U1484 (N_1484,In_620,In_262);
xor U1485 (N_1485,In_590,In_185);
xor U1486 (N_1486,In_598,In_474);
or U1487 (N_1487,In_876,In_784);
nand U1488 (N_1488,In_551,In_780);
or U1489 (N_1489,In_263,In_793);
nor U1490 (N_1490,In_781,In_398);
xnor U1491 (N_1491,In_97,In_447);
xnor U1492 (N_1492,In_303,In_309);
and U1493 (N_1493,In_981,In_332);
nand U1494 (N_1494,In_0,In_693);
nor U1495 (N_1495,In_476,In_925);
or U1496 (N_1496,In_768,In_69);
nand U1497 (N_1497,In_597,In_753);
nand U1498 (N_1498,In_229,In_263);
nor U1499 (N_1499,In_785,In_795);
nor U1500 (N_1500,In_732,In_754);
nand U1501 (N_1501,In_314,In_508);
nor U1502 (N_1502,In_297,In_488);
and U1503 (N_1503,In_643,In_623);
nand U1504 (N_1504,In_668,In_482);
nor U1505 (N_1505,In_311,In_458);
and U1506 (N_1506,In_777,In_535);
and U1507 (N_1507,In_996,In_224);
or U1508 (N_1508,In_515,In_233);
nor U1509 (N_1509,In_656,In_204);
and U1510 (N_1510,In_917,In_218);
and U1511 (N_1511,In_279,In_897);
nor U1512 (N_1512,In_202,In_189);
or U1513 (N_1513,In_452,In_870);
or U1514 (N_1514,In_720,In_859);
or U1515 (N_1515,In_836,In_313);
or U1516 (N_1516,In_17,In_709);
or U1517 (N_1517,In_914,In_4);
and U1518 (N_1518,In_226,In_457);
or U1519 (N_1519,In_885,In_817);
xnor U1520 (N_1520,In_199,In_624);
and U1521 (N_1521,In_647,In_281);
nor U1522 (N_1522,In_889,In_701);
xor U1523 (N_1523,In_505,In_581);
nor U1524 (N_1524,In_461,In_961);
and U1525 (N_1525,In_8,In_882);
and U1526 (N_1526,In_20,In_658);
nand U1527 (N_1527,In_815,In_299);
nand U1528 (N_1528,In_520,In_991);
or U1529 (N_1529,In_709,In_476);
and U1530 (N_1530,In_184,In_20);
and U1531 (N_1531,In_969,In_556);
or U1532 (N_1532,In_663,In_63);
and U1533 (N_1533,In_850,In_968);
xor U1534 (N_1534,In_387,In_114);
nor U1535 (N_1535,In_476,In_887);
or U1536 (N_1536,In_895,In_435);
or U1537 (N_1537,In_584,In_478);
nand U1538 (N_1538,In_198,In_414);
nor U1539 (N_1539,In_687,In_668);
nor U1540 (N_1540,In_723,In_629);
nor U1541 (N_1541,In_609,In_595);
and U1542 (N_1542,In_289,In_443);
or U1543 (N_1543,In_598,In_571);
nor U1544 (N_1544,In_948,In_114);
or U1545 (N_1545,In_850,In_121);
nor U1546 (N_1546,In_167,In_459);
xnor U1547 (N_1547,In_447,In_748);
nand U1548 (N_1548,In_722,In_172);
and U1549 (N_1549,In_587,In_907);
xor U1550 (N_1550,In_362,In_481);
nand U1551 (N_1551,In_824,In_131);
nand U1552 (N_1552,In_46,In_135);
xnor U1553 (N_1553,In_886,In_896);
or U1554 (N_1554,In_224,In_887);
or U1555 (N_1555,In_829,In_391);
nand U1556 (N_1556,In_155,In_755);
nor U1557 (N_1557,In_896,In_87);
or U1558 (N_1558,In_642,In_928);
nor U1559 (N_1559,In_303,In_706);
or U1560 (N_1560,In_517,In_419);
nand U1561 (N_1561,In_743,In_845);
or U1562 (N_1562,In_655,In_653);
and U1563 (N_1563,In_192,In_863);
nor U1564 (N_1564,In_131,In_176);
nand U1565 (N_1565,In_220,In_380);
xor U1566 (N_1566,In_267,In_967);
and U1567 (N_1567,In_374,In_16);
nor U1568 (N_1568,In_609,In_529);
and U1569 (N_1569,In_253,In_719);
nand U1570 (N_1570,In_526,In_376);
or U1571 (N_1571,In_240,In_656);
nand U1572 (N_1572,In_982,In_398);
nor U1573 (N_1573,In_652,In_428);
nand U1574 (N_1574,In_412,In_729);
and U1575 (N_1575,In_309,In_193);
nor U1576 (N_1576,In_190,In_894);
or U1577 (N_1577,In_415,In_599);
xnor U1578 (N_1578,In_292,In_669);
and U1579 (N_1579,In_165,In_895);
or U1580 (N_1580,In_42,In_281);
nor U1581 (N_1581,In_393,In_301);
nand U1582 (N_1582,In_509,In_274);
and U1583 (N_1583,In_959,In_378);
xor U1584 (N_1584,In_722,In_741);
nor U1585 (N_1585,In_810,In_141);
or U1586 (N_1586,In_312,In_408);
and U1587 (N_1587,In_717,In_971);
and U1588 (N_1588,In_534,In_589);
nand U1589 (N_1589,In_602,In_148);
xnor U1590 (N_1590,In_872,In_694);
nand U1591 (N_1591,In_131,In_51);
and U1592 (N_1592,In_659,In_176);
or U1593 (N_1593,In_938,In_980);
xor U1594 (N_1594,In_451,In_255);
nand U1595 (N_1595,In_537,In_400);
and U1596 (N_1596,In_240,In_267);
and U1597 (N_1597,In_733,In_235);
or U1598 (N_1598,In_156,In_883);
nor U1599 (N_1599,In_647,In_930);
nand U1600 (N_1600,In_551,In_540);
xnor U1601 (N_1601,In_929,In_920);
or U1602 (N_1602,In_791,In_618);
nand U1603 (N_1603,In_923,In_212);
or U1604 (N_1604,In_461,In_15);
nor U1605 (N_1605,In_325,In_885);
or U1606 (N_1606,In_522,In_579);
or U1607 (N_1607,In_589,In_962);
xor U1608 (N_1608,In_544,In_550);
or U1609 (N_1609,In_480,In_381);
nand U1610 (N_1610,In_202,In_454);
xnor U1611 (N_1611,In_355,In_709);
or U1612 (N_1612,In_97,In_841);
or U1613 (N_1613,In_972,In_0);
nand U1614 (N_1614,In_937,In_640);
and U1615 (N_1615,In_318,In_76);
nor U1616 (N_1616,In_719,In_873);
and U1617 (N_1617,In_106,In_878);
nand U1618 (N_1618,In_98,In_741);
nor U1619 (N_1619,In_250,In_597);
nor U1620 (N_1620,In_644,In_632);
and U1621 (N_1621,In_475,In_501);
or U1622 (N_1622,In_474,In_453);
nand U1623 (N_1623,In_551,In_765);
nand U1624 (N_1624,In_56,In_444);
nor U1625 (N_1625,In_463,In_674);
nor U1626 (N_1626,In_697,In_436);
and U1627 (N_1627,In_513,In_441);
nand U1628 (N_1628,In_565,In_142);
or U1629 (N_1629,In_207,In_425);
nand U1630 (N_1630,In_835,In_932);
nor U1631 (N_1631,In_980,In_198);
nand U1632 (N_1632,In_988,In_739);
nor U1633 (N_1633,In_477,In_704);
or U1634 (N_1634,In_532,In_984);
and U1635 (N_1635,In_859,In_108);
nor U1636 (N_1636,In_348,In_94);
and U1637 (N_1637,In_665,In_501);
or U1638 (N_1638,In_43,In_129);
and U1639 (N_1639,In_697,In_647);
or U1640 (N_1640,In_452,In_960);
nor U1641 (N_1641,In_286,In_629);
or U1642 (N_1642,In_586,In_839);
and U1643 (N_1643,In_403,In_347);
xnor U1644 (N_1644,In_917,In_434);
nand U1645 (N_1645,In_359,In_583);
or U1646 (N_1646,In_430,In_198);
nand U1647 (N_1647,In_460,In_214);
or U1648 (N_1648,In_286,In_217);
and U1649 (N_1649,In_813,In_828);
and U1650 (N_1650,In_871,In_909);
and U1651 (N_1651,In_302,In_875);
nor U1652 (N_1652,In_809,In_405);
or U1653 (N_1653,In_753,In_430);
nand U1654 (N_1654,In_625,In_13);
xnor U1655 (N_1655,In_719,In_902);
or U1656 (N_1656,In_549,In_821);
xnor U1657 (N_1657,In_595,In_606);
xnor U1658 (N_1658,In_454,In_468);
nor U1659 (N_1659,In_115,In_159);
nor U1660 (N_1660,In_932,In_386);
and U1661 (N_1661,In_426,In_856);
xnor U1662 (N_1662,In_955,In_464);
nor U1663 (N_1663,In_425,In_864);
and U1664 (N_1664,In_309,In_196);
nand U1665 (N_1665,In_590,In_739);
xor U1666 (N_1666,In_999,In_768);
nand U1667 (N_1667,In_794,In_197);
or U1668 (N_1668,In_729,In_998);
and U1669 (N_1669,In_184,In_705);
or U1670 (N_1670,In_952,In_830);
and U1671 (N_1671,In_362,In_897);
and U1672 (N_1672,In_722,In_541);
nor U1673 (N_1673,In_302,In_700);
or U1674 (N_1674,In_30,In_599);
and U1675 (N_1675,In_393,In_827);
or U1676 (N_1676,In_652,In_916);
or U1677 (N_1677,In_230,In_657);
nor U1678 (N_1678,In_231,In_260);
nand U1679 (N_1679,In_543,In_835);
and U1680 (N_1680,In_357,In_785);
nand U1681 (N_1681,In_559,In_128);
nand U1682 (N_1682,In_397,In_364);
or U1683 (N_1683,In_170,In_370);
nor U1684 (N_1684,In_842,In_987);
nand U1685 (N_1685,In_387,In_842);
or U1686 (N_1686,In_741,In_176);
nor U1687 (N_1687,In_427,In_127);
or U1688 (N_1688,In_870,In_113);
and U1689 (N_1689,In_52,In_541);
nor U1690 (N_1690,In_134,In_935);
and U1691 (N_1691,In_836,In_279);
xnor U1692 (N_1692,In_629,In_110);
xor U1693 (N_1693,In_842,In_184);
or U1694 (N_1694,In_909,In_108);
nand U1695 (N_1695,In_895,In_612);
xor U1696 (N_1696,In_774,In_660);
xor U1697 (N_1697,In_965,In_962);
nor U1698 (N_1698,In_703,In_270);
nor U1699 (N_1699,In_255,In_23);
nor U1700 (N_1700,In_853,In_751);
nor U1701 (N_1701,In_491,In_267);
xnor U1702 (N_1702,In_586,In_834);
nor U1703 (N_1703,In_986,In_968);
nor U1704 (N_1704,In_547,In_724);
nand U1705 (N_1705,In_602,In_960);
nand U1706 (N_1706,In_966,In_39);
and U1707 (N_1707,In_170,In_682);
or U1708 (N_1708,In_358,In_42);
nor U1709 (N_1709,In_339,In_961);
and U1710 (N_1710,In_292,In_477);
and U1711 (N_1711,In_23,In_904);
or U1712 (N_1712,In_9,In_601);
nor U1713 (N_1713,In_749,In_619);
nand U1714 (N_1714,In_844,In_967);
and U1715 (N_1715,In_842,In_543);
or U1716 (N_1716,In_527,In_624);
and U1717 (N_1717,In_470,In_413);
and U1718 (N_1718,In_521,In_577);
and U1719 (N_1719,In_95,In_619);
nand U1720 (N_1720,In_503,In_538);
nand U1721 (N_1721,In_629,In_756);
or U1722 (N_1722,In_916,In_159);
and U1723 (N_1723,In_597,In_224);
nor U1724 (N_1724,In_851,In_358);
nand U1725 (N_1725,In_229,In_572);
and U1726 (N_1726,In_272,In_26);
xor U1727 (N_1727,In_110,In_364);
or U1728 (N_1728,In_437,In_755);
and U1729 (N_1729,In_375,In_381);
and U1730 (N_1730,In_635,In_51);
nor U1731 (N_1731,In_666,In_455);
or U1732 (N_1732,In_717,In_819);
nand U1733 (N_1733,In_222,In_384);
nand U1734 (N_1734,In_486,In_678);
and U1735 (N_1735,In_710,In_110);
or U1736 (N_1736,In_543,In_101);
and U1737 (N_1737,In_974,In_566);
and U1738 (N_1738,In_3,In_349);
nand U1739 (N_1739,In_57,In_813);
xnor U1740 (N_1740,In_304,In_525);
nor U1741 (N_1741,In_748,In_696);
nor U1742 (N_1742,In_88,In_776);
and U1743 (N_1743,In_130,In_793);
nor U1744 (N_1744,In_301,In_206);
nor U1745 (N_1745,In_829,In_126);
xnor U1746 (N_1746,In_956,In_340);
nand U1747 (N_1747,In_736,In_942);
nand U1748 (N_1748,In_760,In_731);
and U1749 (N_1749,In_287,In_701);
and U1750 (N_1750,In_485,In_807);
and U1751 (N_1751,In_773,In_240);
nor U1752 (N_1752,In_329,In_861);
and U1753 (N_1753,In_266,In_308);
nor U1754 (N_1754,In_126,In_733);
or U1755 (N_1755,In_306,In_504);
xor U1756 (N_1756,In_252,In_472);
xor U1757 (N_1757,In_64,In_769);
and U1758 (N_1758,In_688,In_786);
nand U1759 (N_1759,In_649,In_995);
nand U1760 (N_1760,In_218,In_42);
nor U1761 (N_1761,In_969,In_548);
or U1762 (N_1762,In_793,In_281);
xor U1763 (N_1763,In_578,In_783);
nand U1764 (N_1764,In_682,In_445);
or U1765 (N_1765,In_831,In_823);
nor U1766 (N_1766,In_136,In_543);
xnor U1767 (N_1767,In_194,In_18);
xor U1768 (N_1768,In_178,In_353);
nand U1769 (N_1769,In_131,In_241);
xor U1770 (N_1770,In_457,In_396);
nor U1771 (N_1771,In_271,In_122);
nor U1772 (N_1772,In_306,In_353);
or U1773 (N_1773,In_493,In_6);
nand U1774 (N_1774,In_269,In_997);
xor U1775 (N_1775,In_264,In_874);
nand U1776 (N_1776,In_307,In_421);
nor U1777 (N_1777,In_196,In_323);
xnor U1778 (N_1778,In_43,In_842);
nor U1779 (N_1779,In_727,In_580);
nor U1780 (N_1780,In_959,In_524);
nor U1781 (N_1781,In_109,In_933);
xor U1782 (N_1782,In_916,In_412);
and U1783 (N_1783,In_804,In_480);
nor U1784 (N_1784,In_945,In_782);
or U1785 (N_1785,In_867,In_868);
and U1786 (N_1786,In_502,In_335);
nor U1787 (N_1787,In_522,In_503);
or U1788 (N_1788,In_991,In_836);
and U1789 (N_1789,In_257,In_214);
nand U1790 (N_1790,In_158,In_918);
nor U1791 (N_1791,In_882,In_284);
nor U1792 (N_1792,In_921,In_168);
or U1793 (N_1793,In_681,In_115);
or U1794 (N_1794,In_788,In_434);
nor U1795 (N_1795,In_412,In_454);
or U1796 (N_1796,In_501,In_278);
nor U1797 (N_1797,In_935,In_73);
and U1798 (N_1798,In_888,In_812);
and U1799 (N_1799,In_398,In_534);
or U1800 (N_1800,In_92,In_269);
nand U1801 (N_1801,In_715,In_55);
or U1802 (N_1802,In_970,In_924);
nand U1803 (N_1803,In_924,In_507);
nor U1804 (N_1804,In_926,In_387);
xnor U1805 (N_1805,In_40,In_573);
nand U1806 (N_1806,In_223,In_443);
or U1807 (N_1807,In_989,In_500);
nor U1808 (N_1808,In_875,In_330);
or U1809 (N_1809,In_851,In_526);
nor U1810 (N_1810,In_641,In_53);
xor U1811 (N_1811,In_151,In_722);
xnor U1812 (N_1812,In_487,In_875);
nand U1813 (N_1813,In_811,In_622);
xnor U1814 (N_1814,In_317,In_76);
nand U1815 (N_1815,In_30,In_906);
or U1816 (N_1816,In_814,In_67);
xnor U1817 (N_1817,In_734,In_279);
xor U1818 (N_1818,In_293,In_117);
xor U1819 (N_1819,In_704,In_457);
and U1820 (N_1820,In_804,In_22);
or U1821 (N_1821,In_379,In_329);
or U1822 (N_1822,In_504,In_125);
and U1823 (N_1823,In_331,In_4);
nand U1824 (N_1824,In_653,In_576);
or U1825 (N_1825,In_577,In_401);
xor U1826 (N_1826,In_284,In_254);
nand U1827 (N_1827,In_112,In_440);
nor U1828 (N_1828,In_87,In_369);
and U1829 (N_1829,In_930,In_863);
nand U1830 (N_1830,In_101,In_776);
xor U1831 (N_1831,In_831,In_606);
xnor U1832 (N_1832,In_527,In_451);
or U1833 (N_1833,In_503,In_238);
xor U1834 (N_1834,In_7,In_596);
xor U1835 (N_1835,In_96,In_728);
nor U1836 (N_1836,In_73,In_418);
xnor U1837 (N_1837,In_212,In_361);
or U1838 (N_1838,In_949,In_13);
xnor U1839 (N_1839,In_412,In_813);
and U1840 (N_1840,In_410,In_709);
or U1841 (N_1841,In_722,In_210);
and U1842 (N_1842,In_435,In_370);
or U1843 (N_1843,In_533,In_894);
and U1844 (N_1844,In_858,In_20);
nor U1845 (N_1845,In_84,In_284);
nand U1846 (N_1846,In_549,In_720);
and U1847 (N_1847,In_685,In_825);
nor U1848 (N_1848,In_508,In_628);
nor U1849 (N_1849,In_895,In_172);
xnor U1850 (N_1850,In_531,In_373);
and U1851 (N_1851,In_143,In_614);
and U1852 (N_1852,In_199,In_399);
xor U1853 (N_1853,In_850,In_770);
xor U1854 (N_1854,In_645,In_126);
or U1855 (N_1855,In_91,In_115);
nor U1856 (N_1856,In_736,In_887);
nor U1857 (N_1857,In_425,In_252);
nand U1858 (N_1858,In_8,In_465);
xnor U1859 (N_1859,In_502,In_997);
nand U1860 (N_1860,In_498,In_379);
and U1861 (N_1861,In_945,In_568);
and U1862 (N_1862,In_605,In_723);
xnor U1863 (N_1863,In_459,In_768);
or U1864 (N_1864,In_575,In_138);
nor U1865 (N_1865,In_394,In_485);
nor U1866 (N_1866,In_38,In_142);
xnor U1867 (N_1867,In_474,In_502);
and U1868 (N_1868,In_108,In_224);
nor U1869 (N_1869,In_324,In_54);
xor U1870 (N_1870,In_699,In_110);
xor U1871 (N_1871,In_916,In_235);
nand U1872 (N_1872,In_495,In_137);
xnor U1873 (N_1873,In_592,In_186);
and U1874 (N_1874,In_396,In_279);
or U1875 (N_1875,In_846,In_815);
xnor U1876 (N_1876,In_886,In_636);
or U1877 (N_1877,In_703,In_146);
or U1878 (N_1878,In_796,In_165);
and U1879 (N_1879,In_596,In_158);
or U1880 (N_1880,In_980,In_74);
xor U1881 (N_1881,In_389,In_144);
nand U1882 (N_1882,In_376,In_26);
or U1883 (N_1883,In_981,In_615);
and U1884 (N_1884,In_771,In_134);
and U1885 (N_1885,In_749,In_590);
nor U1886 (N_1886,In_135,In_265);
nand U1887 (N_1887,In_137,In_630);
nand U1888 (N_1888,In_984,In_115);
and U1889 (N_1889,In_298,In_738);
or U1890 (N_1890,In_2,In_459);
nor U1891 (N_1891,In_906,In_672);
or U1892 (N_1892,In_842,In_119);
nand U1893 (N_1893,In_4,In_889);
or U1894 (N_1894,In_758,In_48);
or U1895 (N_1895,In_514,In_333);
nor U1896 (N_1896,In_86,In_323);
nor U1897 (N_1897,In_261,In_867);
nand U1898 (N_1898,In_313,In_910);
or U1899 (N_1899,In_948,In_9);
nor U1900 (N_1900,In_724,In_428);
and U1901 (N_1901,In_494,In_185);
nand U1902 (N_1902,In_21,In_699);
xnor U1903 (N_1903,In_705,In_516);
xor U1904 (N_1904,In_125,In_978);
nor U1905 (N_1905,In_832,In_484);
xnor U1906 (N_1906,In_860,In_1);
nor U1907 (N_1907,In_553,In_229);
nand U1908 (N_1908,In_729,In_651);
nor U1909 (N_1909,In_910,In_554);
nand U1910 (N_1910,In_319,In_489);
nand U1911 (N_1911,In_483,In_326);
or U1912 (N_1912,In_917,In_606);
or U1913 (N_1913,In_857,In_407);
nor U1914 (N_1914,In_48,In_194);
nor U1915 (N_1915,In_992,In_830);
xor U1916 (N_1916,In_835,In_68);
nor U1917 (N_1917,In_128,In_720);
nand U1918 (N_1918,In_114,In_966);
and U1919 (N_1919,In_41,In_604);
or U1920 (N_1920,In_972,In_311);
nor U1921 (N_1921,In_595,In_126);
nor U1922 (N_1922,In_887,In_213);
and U1923 (N_1923,In_386,In_242);
xor U1924 (N_1924,In_733,In_780);
xor U1925 (N_1925,In_546,In_423);
or U1926 (N_1926,In_268,In_588);
or U1927 (N_1927,In_165,In_481);
xnor U1928 (N_1928,In_363,In_872);
or U1929 (N_1929,In_852,In_953);
or U1930 (N_1930,In_770,In_302);
nor U1931 (N_1931,In_245,In_761);
xnor U1932 (N_1932,In_551,In_363);
nor U1933 (N_1933,In_656,In_82);
or U1934 (N_1934,In_33,In_644);
and U1935 (N_1935,In_161,In_307);
xnor U1936 (N_1936,In_446,In_417);
xnor U1937 (N_1937,In_543,In_669);
xor U1938 (N_1938,In_302,In_988);
nand U1939 (N_1939,In_395,In_422);
or U1940 (N_1940,In_698,In_669);
xor U1941 (N_1941,In_935,In_524);
or U1942 (N_1942,In_177,In_565);
nand U1943 (N_1943,In_811,In_560);
xor U1944 (N_1944,In_722,In_967);
or U1945 (N_1945,In_436,In_577);
nor U1946 (N_1946,In_849,In_133);
nand U1947 (N_1947,In_8,In_741);
and U1948 (N_1948,In_934,In_692);
xor U1949 (N_1949,In_256,In_171);
nand U1950 (N_1950,In_794,In_571);
nor U1951 (N_1951,In_576,In_283);
or U1952 (N_1952,In_113,In_738);
or U1953 (N_1953,In_94,In_966);
nand U1954 (N_1954,In_609,In_745);
and U1955 (N_1955,In_685,In_775);
xor U1956 (N_1956,In_365,In_777);
xor U1957 (N_1957,In_125,In_360);
nand U1958 (N_1958,In_65,In_397);
nor U1959 (N_1959,In_15,In_63);
or U1960 (N_1960,In_785,In_883);
and U1961 (N_1961,In_266,In_332);
xnor U1962 (N_1962,In_79,In_19);
xnor U1963 (N_1963,In_411,In_46);
or U1964 (N_1964,In_421,In_738);
and U1965 (N_1965,In_613,In_218);
nor U1966 (N_1966,In_551,In_231);
nor U1967 (N_1967,In_715,In_283);
nor U1968 (N_1968,In_684,In_10);
and U1969 (N_1969,In_543,In_4);
nand U1970 (N_1970,In_818,In_920);
nor U1971 (N_1971,In_101,In_902);
nand U1972 (N_1972,In_307,In_432);
nand U1973 (N_1973,In_328,In_721);
nor U1974 (N_1974,In_432,In_594);
and U1975 (N_1975,In_459,In_710);
or U1976 (N_1976,In_279,In_543);
or U1977 (N_1977,In_287,In_388);
and U1978 (N_1978,In_678,In_864);
and U1979 (N_1979,In_817,In_840);
nor U1980 (N_1980,In_225,In_701);
nand U1981 (N_1981,In_50,In_955);
nand U1982 (N_1982,In_904,In_679);
and U1983 (N_1983,In_617,In_2);
nand U1984 (N_1984,In_969,In_9);
nor U1985 (N_1985,In_855,In_711);
nor U1986 (N_1986,In_231,In_622);
nor U1987 (N_1987,In_48,In_56);
or U1988 (N_1988,In_825,In_211);
and U1989 (N_1989,In_550,In_915);
xor U1990 (N_1990,In_367,In_188);
nor U1991 (N_1991,In_8,In_187);
xnor U1992 (N_1992,In_427,In_281);
and U1993 (N_1993,In_276,In_568);
and U1994 (N_1994,In_550,In_486);
and U1995 (N_1995,In_847,In_309);
and U1996 (N_1996,In_893,In_610);
and U1997 (N_1997,In_366,In_901);
nor U1998 (N_1998,In_855,In_475);
or U1999 (N_1999,In_586,In_293);
or U2000 (N_2000,In_984,In_497);
or U2001 (N_2001,In_224,In_713);
nor U2002 (N_2002,In_969,In_46);
xnor U2003 (N_2003,In_296,In_663);
and U2004 (N_2004,In_67,In_959);
nor U2005 (N_2005,In_397,In_592);
nor U2006 (N_2006,In_12,In_146);
nor U2007 (N_2007,In_570,In_579);
and U2008 (N_2008,In_667,In_595);
nand U2009 (N_2009,In_131,In_822);
xnor U2010 (N_2010,In_15,In_980);
xor U2011 (N_2011,In_862,In_534);
xor U2012 (N_2012,In_760,In_78);
nor U2013 (N_2013,In_112,In_156);
nor U2014 (N_2014,In_849,In_9);
or U2015 (N_2015,In_527,In_962);
and U2016 (N_2016,In_670,In_825);
or U2017 (N_2017,In_645,In_725);
nor U2018 (N_2018,In_960,In_878);
nor U2019 (N_2019,In_684,In_903);
or U2020 (N_2020,In_191,In_63);
or U2021 (N_2021,In_401,In_78);
and U2022 (N_2022,In_449,In_251);
and U2023 (N_2023,In_175,In_600);
nor U2024 (N_2024,In_534,In_979);
nand U2025 (N_2025,In_241,In_40);
and U2026 (N_2026,In_3,In_392);
or U2027 (N_2027,In_555,In_559);
xnor U2028 (N_2028,In_849,In_991);
and U2029 (N_2029,In_287,In_269);
nor U2030 (N_2030,In_503,In_791);
xor U2031 (N_2031,In_357,In_676);
nand U2032 (N_2032,In_806,In_357);
nand U2033 (N_2033,In_799,In_953);
nand U2034 (N_2034,In_377,In_465);
nand U2035 (N_2035,In_377,In_640);
and U2036 (N_2036,In_957,In_838);
nand U2037 (N_2037,In_0,In_257);
nand U2038 (N_2038,In_495,In_412);
nand U2039 (N_2039,In_289,In_132);
and U2040 (N_2040,In_86,In_208);
nor U2041 (N_2041,In_435,In_780);
nand U2042 (N_2042,In_189,In_846);
and U2043 (N_2043,In_678,In_400);
and U2044 (N_2044,In_704,In_282);
nor U2045 (N_2045,In_860,In_297);
and U2046 (N_2046,In_819,In_353);
and U2047 (N_2047,In_429,In_373);
nand U2048 (N_2048,In_698,In_990);
xor U2049 (N_2049,In_46,In_842);
or U2050 (N_2050,In_939,In_707);
nand U2051 (N_2051,In_149,In_899);
and U2052 (N_2052,In_660,In_654);
nand U2053 (N_2053,In_455,In_248);
nor U2054 (N_2054,In_591,In_166);
nand U2055 (N_2055,In_730,In_153);
or U2056 (N_2056,In_516,In_183);
or U2057 (N_2057,In_849,In_233);
or U2058 (N_2058,In_579,In_576);
or U2059 (N_2059,In_281,In_333);
nor U2060 (N_2060,In_860,In_365);
nand U2061 (N_2061,In_272,In_640);
xnor U2062 (N_2062,In_772,In_445);
xor U2063 (N_2063,In_674,In_905);
and U2064 (N_2064,In_672,In_8);
and U2065 (N_2065,In_782,In_990);
and U2066 (N_2066,In_576,In_718);
and U2067 (N_2067,In_69,In_510);
and U2068 (N_2068,In_866,In_218);
xnor U2069 (N_2069,In_205,In_80);
or U2070 (N_2070,In_211,In_802);
xnor U2071 (N_2071,In_773,In_96);
and U2072 (N_2072,In_992,In_94);
xor U2073 (N_2073,In_580,In_131);
nand U2074 (N_2074,In_619,In_461);
and U2075 (N_2075,In_999,In_791);
xor U2076 (N_2076,In_122,In_120);
and U2077 (N_2077,In_390,In_920);
and U2078 (N_2078,In_723,In_345);
and U2079 (N_2079,In_272,In_715);
or U2080 (N_2080,In_327,In_845);
nand U2081 (N_2081,In_42,In_834);
and U2082 (N_2082,In_379,In_829);
and U2083 (N_2083,In_119,In_678);
or U2084 (N_2084,In_214,In_986);
xor U2085 (N_2085,In_347,In_513);
nand U2086 (N_2086,In_912,In_615);
nand U2087 (N_2087,In_783,In_524);
nor U2088 (N_2088,In_353,In_36);
nand U2089 (N_2089,In_501,In_573);
nor U2090 (N_2090,In_802,In_487);
or U2091 (N_2091,In_866,In_968);
xor U2092 (N_2092,In_142,In_190);
xnor U2093 (N_2093,In_425,In_972);
nor U2094 (N_2094,In_525,In_388);
nor U2095 (N_2095,In_735,In_677);
nor U2096 (N_2096,In_235,In_82);
xnor U2097 (N_2097,In_961,In_374);
and U2098 (N_2098,In_136,In_497);
xnor U2099 (N_2099,In_271,In_160);
nor U2100 (N_2100,In_740,In_471);
or U2101 (N_2101,In_254,In_443);
nand U2102 (N_2102,In_306,In_738);
nor U2103 (N_2103,In_627,In_82);
nand U2104 (N_2104,In_652,In_668);
and U2105 (N_2105,In_164,In_957);
xnor U2106 (N_2106,In_901,In_389);
nand U2107 (N_2107,In_883,In_549);
nor U2108 (N_2108,In_299,In_247);
nor U2109 (N_2109,In_232,In_12);
and U2110 (N_2110,In_293,In_330);
xnor U2111 (N_2111,In_275,In_129);
xor U2112 (N_2112,In_431,In_545);
or U2113 (N_2113,In_845,In_99);
and U2114 (N_2114,In_757,In_826);
xor U2115 (N_2115,In_862,In_793);
nor U2116 (N_2116,In_983,In_240);
nand U2117 (N_2117,In_612,In_352);
or U2118 (N_2118,In_345,In_826);
xnor U2119 (N_2119,In_460,In_239);
nor U2120 (N_2120,In_176,In_195);
xor U2121 (N_2121,In_169,In_828);
xnor U2122 (N_2122,In_661,In_215);
nor U2123 (N_2123,In_699,In_662);
xnor U2124 (N_2124,In_382,In_587);
or U2125 (N_2125,In_859,In_396);
and U2126 (N_2126,In_287,In_183);
nand U2127 (N_2127,In_156,In_159);
nand U2128 (N_2128,In_410,In_773);
or U2129 (N_2129,In_469,In_652);
or U2130 (N_2130,In_912,In_863);
nand U2131 (N_2131,In_431,In_103);
nand U2132 (N_2132,In_676,In_69);
and U2133 (N_2133,In_270,In_941);
or U2134 (N_2134,In_619,In_46);
and U2135 (N_2135,In_683,In_418);
xnor U2136 (N_2136,In_429,In_410);
nand U2137 (N_2137,In_383,In_681);
xor U2138 (N_2138,In_976,In_153);
nand U2139 (N_2139,In_389,In_302);
or U2140 (N_2140,In_35,In_567);
xnor U2141 (N_2141,In_996,In_267);
nand U2142 (N_2142,In_597,In_239);
or U2143 (N_2143,In_760,In_384);
and U2144 (N_2144,In_306,In_552);
nor U2145 (N_2145,In_793,In_43);
and U2146 (N_2146,In_843,In_135);
nand U2147 (N_2147,In_33,In_779);
nand U2148 (N_2148,In_907,In_148);
nor U2149 (N_2149,In_21,In_236);
or U2150 (N_2150,In_288,In_105);
nand U2151 (N_2151,In_662,In_465);
nand U2152 (N_2152,In_633,In_989);
and U2153 (N_2153,In_337,In_718);
nor U2154 (N_2154,In_773,In_351);
nor U2155 (N_2155,In_884,In_785);
or U2156 (N_2156,In_722,In_963);
or U2157 (N_2157,In_17,In_547);
nand U2158 (N_2158,In_170,In_60);
nand U2159 (N_2159,In_393,In_77);
and U2160 (N_2160,In_540,In_797);
xnor U2161 (N_2161,In_601,In_790);
or U2162 (N_2162,In_257,In_509);
or U2163 (N_2163,In_517,In_876);
or U2164 (N_2164,In_66,In_249);
xnor U2165 (N_2165,In_175,In_9);
nor U2166 (N_2166,In_424,In_745);
xnor U2167 (N_2167,In_416,In_434);
nand U2168 (N_2168,In_288,In_658);
or U2169 (N_2169,In_14,In_197);
or U2170 (N_2170,In_845,In_777);
nand U2171 (N_2171,In_782,In_350);
nand U2172 (N_2172,In_902,In_569);
or U2173 (N_2173,In_674,In_954);
and U2174 (N_2174,In_185,In_802);
xnor U2175 (N_2175,In_271,In_87);
xor U2176 (N_2176,In_536,In_670);
nor U2177 (N_2177,In_125,In_687);
or U2178 (N_2178,In_307,In_549);
or U2179 (N_2179,In_883,In_981);
nor U2180 (N_2180,In_630,In_825);
or U2181 (N_2181,In_206,In_603);
xor U2182 (N_2182,In_290,In_299);
or U2183 (N_2183,In_531,In_739);
nor U2184 (N_2184,In_697,In_185);
or U2185 (N_2185,In_950,In_112);
and U2186 (N_2186,In_336,In_175);
and U2187 (N_2187,In_562,In_891);
and U2188 (N_2188,In_883,In_52);
and U2189 (N_2189,In_36,In_502);
nor U2190 (N_2190,In_131,In_469);
and U2191 (N_2191,In_10,In_671);
and U2192 (N_2192,In_686,In_738);
nor U2193 (N_2193,In_487,In_722);
or U2194 (N_2194,In_978,In_912);
nor U2195 (N_2195,In_677,In_872);
nor U2196 (N_2196,In_444,In_512);
or U2197 (N_2197,In_2,In_434);
or U2198 (N_2198,In_581,In_306);
and U2199 (N_2199,In_690,In_995);
xor U2200 (N_2200,In_489,In_746);
nor U2201 (N_2201,In_94,In_61);
nor U2202 (N_2202,In_857,In_92);
nand U2203 (N_2203,In_88,In_135);
nor U2204 (N_2204,In_899,In_823);
nand U2205 (N_2205,In_793,In_267);
or U2206 (N_2206,In_716,In_737);
or U2207 (N_2207,In_231,In_905);
and U2208 (N_2208,In_400,In_185);
xor U2209 (N_2209,In_937,In_479);
or U2210 (N_2210,In_362,In_41);
nand U2211 (N_2211,In_352,In_687);
nand U2212 (N_2212,In_705,In_295);
xnor U2213 (N_2213,In_107,In_687);
and U2214 (N_2214,In_381,In_522);
or U2215 (N_2215,In_295,In_107);
nand U2216 (N_2216,In_754,In_998);
and U2217 (N_2217,In_520,In_15);
or U2218 (N_2218,In_988,In_190);
or U2219 (N_2219,In_738,In_793);
xnor U2220 (N_2220,In_830,In_711);
and U2221 (N_2221,In_607,In_247);
nand U2222 (N_2222,In_693,In_840);
or U2223 (N_2223,In_926,In_280);
and U2224 (N_2224,In_739,In_270);
or U2225 (N_2225,In_475,In_480);
nor U2226 (N_2226,In_913,In_354);
and U2227 (N_2227,In_145,In_629);
nand U2228 (N_2228,In_0,In_663);
nor U2229 (N_2229,In_118,In_376);
nor U2230 (N_2230,In_538,In_941);
and U2231 (N_2231,In_212,In_603);
nor U2232 (N_2232,In_769,In_475);
xnor U2233 (N_2233,In_26,In_802);
xnor U2234 (N_2234,In_364,In_947);
nor U2235 (N_2235,In_308,In_578);
nor U2236 (N_2236,In_107,In_481);
xnor U2237 (N_2237,In_452,In_951);
or U2238 (N_2238,In_423,In_775);
xnor U2239 (N_2239,In_325,In_753);
nand U2240 (N_2240,In_491,In_727);
nand U2241 (N_2241,In_325,In_968);
or U2242 (N_2242,In_30,In_108);
and U2243 (N_2243,In_588,In_934);
nand U2244 (N_2244,In_354,In_489);
nor U2245 (N_2245,In_90,In_726);
or U2246 (N_2246,In_456,In_644);
and U2247 (N_2247,In_541,In_893);
or U2248 (N_2248,In_679,In_315);
or U2249 (N_2249,In_87,In_297);
nor U2250 (N_2250,In_232,In_912);
or U2251 (N_2251,In_878,In_678);
nand U2252 (N_2252,In_846,In_717);
or U2253 (N_2253,In_866,In_306);
and U2254 (N_2254,In_544,In_210);
nor U2255 (N_2255,In_451,In_749);
nor U2256 (N_2256,In_123,In_374);
or U2257 (N_2257,In_55,In_745);
or U2258 (N_2258,In_443,In_643);
or U2259 (N_2259,In_973,In_156);
nand U2260 (N_2260,In_506,In_202);
nand U2261 (N_2261,In_73,In_972);
and U2262 (N_2262,In_327,In_960);
xnor U2263 (N_2263,In_320,In_3);
nor U2264 (N_2264,In_753,In_675);
nor U2265 (N_2265,In_979,In_357);
or U2266 (N_2266,In_405,In_968);
or U2267 (N_2267,In_769,In_753);
nor U2268 (N_2268,In_891,In_170);
nand U2269 (N_2269,In_442,In_740);
nor U2270 (N_2270,In_233,In_386);
or U2271 (N_2271,In_545,In_236);
nor U2272 (N_2272,In_220,In_674);
and U2273 (N_2273,In_921,In_309);
xor U2274 (N_2274,In_363,In_86);
or U2275 (N_2275,In_818,In_597);
xnor U2276 (N_2276,In_117,In_570);
nand U2277 (N_2277,In_858,In_551);
or U2278 (N_2278,In_555,In_128);
nor U2279 (N_2279,In_639,In_326);
xor U2280 (N_2280,In_62,In_875);
xnor U2281 (N_2281,In_483,In_404);
and U2282 (N_2282,In_862,In_42);
or U2283 (N_2283,In_452,In_983);
and U2284 (N_2284,In_789,In_359);
and U2285 (N_2285,In_961,In_716);
or U2286 (N_2286,In_956,In_853);
nand U2287 (N_2287,In_921,In_402);
and U2288 (N_2288,In_206,In_324);
nand U2289 (N_2289,In_426,In_544);
nor U2290 (N_2290,In_175,In_178);
xnor U2291 (N_2291,In_592,In_72);
nand U2292 (N_2292,In_610,In_152);
and U2293 (N_2293,In_989,In_506);
and U2294 (N_2294,In_313,In_29);
nor U2295 (N_2295,In_579,In_238);
xor U2296 (N_2296,In_127,In_458);
nor U2297 (N_2297,In_896,In_422);
xnor U2298 (N_2298,In_911,In_960);
nand U2299 (N_2299,In_555,In_872);
nor U2300 (N_2300,In_635,In_163);
xnor U2301 (N_2301,In_621,In_658);
and U2302 (N_2302,In_482,In_161);
or U2303 (N_2303,In_458,In_391);
xnor U2304 (N_2304,In_327,In_970);
nor U2305 (N_2305,In_192,In_594);
or U2306 (N_2306,In_267,In_589);
nand U2307 (N_2307,In_257,In_22);
or U2308 (N_2308,In_784,In_921);
and U2309 (N_2309,In_606,In_704);
nor U2310 (N_2310,In_38,In_782);
or U2311 (N_2311,In_386,In_238);
xor U2312 (N_2312,In_869,In_297);
or U2313 (N_2313,In_536,In_156);
xor U2314 (N_2314,In_370,In_636);
xnor U2315 (N_2315,In_873,In_624);
or U2316 (N_2316,In_292,In_413);
nand U2317 (N_2317,In_631,In_65);
and U2318 (N_2318,In_879,In_880);
xnor U2319 (N_2319,In_845,In_879);
or U2320 (N_2320,In_542,In_805);
nor U2321 (N_2321,In_222,In_496);
and U2322 (N_2322,In_170,In_339);
nand U2323 (N_2323,In_124,In_230);
and U2324 (N_2324,In_568,In_679);
nor U2325 (N_2325,In_557,In_51);
nand U2326 (N_2326,In_352,In_322);
nor U2327 (N_2327,In_844,In_124);
and U2328 (N_2328,In_107,In_541);
or U2329 (N_2329,In_206,In_106);
and U2330 (N_2330,In_50,In_455);
and U2331 (N_2331,In_167,In_935);
nor U2332 (N_2332,In_415,In_642);
nand U2333 (N_2333,In_780,In_89);
xnor U2334 (N_2334,In_778,In_20);
xnor U2335 (N_2335,In_515,In_733);
nand U2336 (N_2336,In_222,In_236);
and U2337 (N_2337,In_194,In_99);
or U2338 (N_2338,In_218,In_137);
and U2339 (N_2339,In_310,In_56);
or U2340 (N_2340,In_581,In_124);
nor U2341 (N_2341,In_218,In_685);
and U2342 (N_2342,In_220,In_173);
or U2343 (N_2343,In_549,In_93);
xor U2344 (N_2344,In_341,In_308);
xor U2345 (N_2345,In_402,In_316);
nand U2346 (N_2346,In_378,In_112);
and U2347 (N_2347,In_408,In_169);
or U2348 (N_2348,In_571,In_163);
or U2349 (N_2349,In_794,In_942);
nor U2350 (N_2350,In_866,In_822);
nor U2351 (N_2351,In_506,In_645);
nand U2352 (N_2352,In_565,In_567);
nand U2353 (N_2353,In_381,In_354);
nand U2354 (N_2354,In_224,In_783);
xor U2355 (N_2355,In_202,In_220);
or U2356 (N_2356,In_230,In_263);
nand U2357 (N_2357,In_770,In_707);
xnor U2358 (N_2358,In_474,In_492);
and U2359 (N_2359,In_308,In_712);
nand U2360 (N_2360,In_92,In_691);
and U2361 (N_2361,In_260,In_735);
and U2362 (N_2362,In_370,In_946);
nand U2363 (N_2363,In_341,In_337);
or U2364 (N_2364,In_780,In_620);
xnor U2365 (N_2365,In_570,In_414);
nand U2366 (N_2366,In_506,In_791);
nor U2367 (N_2367,In_863,In_856);
nor U2368 (N_2368,In_642,In_913);
nor U2369 (N_2369,In_504,In_235);
nand U2370 (N_2370,In_496,In_202);
or U2371 (N_2371,In_541,In_987);
or U2372 (N_2372,In_513,In_211);
nand U2373 (N_2373,In_383,In_124);
and U2374 (N_2374,In_805,In_929);
nor U2375 (N_2375,In_764,In_595);
and U2376 (N_2376,In_610,In_796);
nand U2377 (N_2377,In_563,In_24);
xnor U2378 (N_2378,In_649,In_50);
or U2379 (N_2379,In_663,In_920);
nor U2380 (N_2380,In_15,In_985);
and U2381 (N_2381,In_846,In_954);
nand U2382 (N_2382,In_596,In_792);
and U2383 (N_2383,In_460,In_536);
nor U2384 (N_2384,In_217,In_727);
and U2385 (N_2385,In_496,In_979);
and U2386 (N_2386,In_675,In_179);
or U2387 (N_2387,In_20,In_354);
and U2388 (N_2388,In_998,In_40);
nor U2389 (N_2389,In_101,In_601);
nand U2390 (N_2390,In_950,In_910);
nor U2391 (N_2391,In_260,In_93);
and U2392 (N_2392,In_790,In_451);
nor U2393 (N_2393,In_456,In_824);
nand U2394 (N_2394,In_472,In_207);
xnor U2395 (N_2395,In_989,In_39);
or U2396 (N_2396,In_677,In_631);
xnor U2397 (N_2397,In_869,In_562);
nor U2398 (N_2398,In_512,In_244);
nor U2399 (N_2399,In_686,In_110);
nor U2400 (N_2400,In_540,In_295);
nand U2401 (N_2401,In_778,In_390);
nor U2402 (N_2402,In_965,In_706);
and U2403 (N_2403,In_965,In_33);
or U2404 (N_2404,In_57,In_710);
nor U2405 (N_2405,In_587,In_128);
nor U2406 (N_2406,In_498,In_473);
nor U2407 (N_2407,In_854,In_684);
nor U2408 (N_2408,In_167,In_171);
xnor U2409 (N_2409,In_221,In_641);
and U2410 (N_2410,In_140,In_803);
and U2411 (N_2411,In_163,In_449);
or U2412 (N_2412,In_312,In_2);
nand U2413 (N_2413,In_104,In_652);
nor U2414 (N_2414,In_616,In_584);
xor U2415 (N_2415,In_18,In_286);
or U2416 (N_2416,In_579,In_738);
nor U2417 (N_2417,In_302,In_263);
xor U2418 (N_2418,In_236,In_74);
or U2419 (N_2419,In_686,In_908);
and U2420 (N_2420,In_30,In_863);
or U2421 (N_2421,In_323,In_264);
xnor U2422 (N_2422,In_984,In_226);
nor U2423 (N_2423,In_250,In_344);
nor U2424 (N_2424,In_986,In_21);
or U2425 (N_2425,In_562,In_699);
nor U2426 (N_2426,In_490,In_526);
nand U2427 (N_2427,In_312,In_908);
or U2428 (N_2428,In_737,In_26);
and U2429 (N_2429,In_941,In_439);
and U2430 (N_2430,In_15,In_87);
xnor U2431 (N_2431,In_951,In_158);
nor U2432 (N_2432,In_190,In_754);
xor U2433 (N_2433,In_100,In_326);
and U2434 (N_2434,In_33,In_828);
nor U2435 (N_2435,In_421,In_334);
nand U2436 (N_2436,In_945,In_178);
nor U2437 (N_2437,In_594,In_816);
xnor U2438 (N_2438,In_619,In_351);
and U2439 (N_2439,In_411,In_38);
and U2440 (N_2440,In_655,In_119);
xor U2441 (N_2441,In_407,In_409);
xor U2442 (N_2442,In_783,In_172);
xor U2443 (N_2443,In_367,In_103);
and U2444 (N_2444,In_79,In_18);
and U2445 (N_2445,In_413,In_643);
nand U2446 (N_2446,In_73,In_466);
nor U2447 (N_2447,In_210,In_87);
xnor U2448 (N_2448,In_593,In_616);
xor U2449 (N_2449,In_65,In_690);
or U2450 (N_2450,In_438,In_492);
and U2451 (N_2451,In_374,In_692);
nor U2452 (N_2452,In_455,In_326);
nor U2453 (N_2453,In_466,In_573);
or U2454 (N_2454,In_792,In_147);
or U2455 (N_2455,In_797,In_850);
and U2456 (N_2456,In_316,In_263);
and U2457 (N_2457,In_848,In_213);
xnor U2458 (N_2458,In_884,In_81);
nor U2459 (N_2459,In_82,In_588);
nand U2460 (N_2460,In_907,In_220);
xor U2461 (N_2461,In_588,In_830);
nand U2462 (N_2462,In_671,In_504);
nand U2463 (N_2463,In_460,In_25);
nand U2464 (N_2464,In_453,In_563);
and U2465 (N_2465,In_534,In_687);
xnor U2466 (N_2466,In_507,In_811);
xnor U2467 (N_2467,In_822,In_626);
nor U2468 (N_2468,In_29,In_115);
and U2469 (N_2469,In_592,In_82);
and U2470 (N_2470,In_506,In_218);
and U2471 (N_2471,In_417,In_375);
xor U2472 (N_2472,In_412,In_541);
nand U2473 (N_2473,In_685,In_557);
nor U2474 (N_2474,In_217,In_99);
xnor U2475 (N_2475,In_978,In_117);
and U2476 (N_2476,In_3,In_988);
and U2477 (N_2477,In_111,In_133);
or U2478 (N_2478,In_156,In_504);
nand U2479 (N_2479,In_488,In_526);
and U2480 (N_2480,In_984,In_423);
nor U2481 (N_2481,In_154,In_500);
and U2482 (N_2482,In_405,In_635);
nand U2483 (N_2483,In_917,In_865);
nand U2484 (N_2484,In_374,In_601);
nand U2485 (N_2485,In_11,In_306);
xor U2486 (N_2486,In_311,In_341);
and U2487 (N_2487,In_613,In_707);
or U2488 (N_2488,In_915,In_613);
or U2489 (N_2489,In_944,In_549);
and U2490 (N_2490,In_799,In_139);
nor U2491 (N_2491,In_972,In_599);
and U2492 (N_2492,In_660,In_497);
nor U2493 (N_2493,In_141,In_352);
xor U2494 (N_2494,In_364,In_614);
nand U2495 (N_2495,In_2,In_349);
nor U2496 (N_2496,In_939,In_308);
nand U2497 (N_2497,In_610,In_428);
xor U2498 (N_2498,In_257,In_414);
or U2499 (N_2499,In_808,In_32);
nand U2500 (N_2500,In_897,In_785);
xor U2501 (N_2501,In_961,In_77);
nand U2502 (N_2502,In_42,In_258);
nand U2503 (N_2503,In_105,In_99);
or U2504 (N_2504,In_136,In_713);
nor U2505 (N_2505,In_574,In_506);
xnor U2506 (N_2506,In_369,In_728);
nor U2507 (N_2507,In_347,In_975);
and U2508 (N_2508,In_880,In_134);
and U2509 (N_2509,In_223,In_754);
or U2510 (N_2510,In_41,In_522);
nand U2511 (N_2511,In_777,In_163);
and U2512 (N_2512,In_608,In_179);
or U2513 (N_2513,In_348,In_442);
xnor U2514 (N_2514,In_616,In_53);
nand U2515 (N_2515,In_306,In_750);
nor U2516 (N_2516,In_732,In_718);
nor U2517 (N_2517,In_209,In_256);
xnor U2518 (N_2518,In_362,In_378);
and U2519 (N_2519,In_774,In_582);
nand U2520 (N_2520,In_443,In_834);
nor U2521 (N_2521,In_130,In_93);
xor U2522 (N_2522,In_873,In_922);
xor U2523 (N_2523,In_392,In_25);
xnor U2524 (N_2524,In_370,In_883);
xnor U2525 (N_2525,In_992,In_258);
or U2526 (N_2526,In_166,In_744);
and U2527 (N_2527,In_716,In_418);
nand U2528 (N_2528,In_632,In_947);
nor U2529 (N_2529,In_133,In_956);
or U2530 (N_2530,In_648,In_317);
xnor U2531 (N_2531,In_359,In_607);
nor U2532 (N_2532,In_935,In_47);
xnor U2533 (N_2533,In_23,In_517);
or U2534 (N_2534,In_97,In_631);
or U2535 (N_2535,In_522,In_30);
or U2536 (N_2536,In_725,In_324);
and U2537 (N_2537,In_265,In_238);
and U2538 (N_2538,In_245,In_488);
nor U2539 (N_2539,In_259,In_950);
and U2540 (N_2540,In_565,In_806);
xor U2541 (N_2541,In_917,In_741);
xnor U2542 (N_2542,In_549,In_862);
and U2543 (N_2543,In_217,In_619);
xnor U2544 (N_2544,In_749,In_674);
nor U2545 (N_2545,In_942,In_572);
nor U2546 (N_2546,In_340,In_489);
nand U2547 (N_2547,In_609,In_224);
nand U2548 (N_2548,In_414,In_29);
and U2549 (N_2549,In_68,In_398);
nand U2550 (N_2550,In_251,In_988);
and U2551 (N_2551,In_241,In_823);
or U2552 (N_2552,In_755,In_438);
and U2553 (N_2553,In_726,In_94);
or U2554 (N_2554,In_265,In_534);
and U2555 (N_2555,In_824,In_361);
or U2556 (N_2556,In_458,In_543);
nor U2557 (N_2557,In_655,In_270);
and U2558 (N_2558,In_928,In_572);
or U2559 (N_2559,In_731,In_499);
nor U2560 (N_2560,In_324,In_100);
nor U2561 (N_2561,In_27,In_731);
and U2562 (N_2562,In_173,In_536);
or U2563 (N_2563,In_891,In_339);
or U2564 (N_2564,In_624,In_654);
and U2565 (N_2565,In_787,In_382);
nor U2566 (N_2566,In_246,In_266);
and U2567 (N_2567,In_843,In_104);
or U2568 (N_2568,In_322,In_816);
nand U2569 (N_2569,In_632,In_979);
xnor U2570 (N_2570,In_711,In_178);
or U2571 (N_2571,In_545,In_235);
or U2572 (N_2572,In_652,In_129);
nor U2573 (N_2573,In_659,In_876);
nand U2574 (N_2574,In_70,In_423);
and U2575 (N_2575,In_792,In_503);
nand U2576 (N_2576,In_915,In_358);
nand U2577 (N_2577,In_78,In_421);
xnor U2578 (N_2578,In_921,In_293);
or U2579 (N_2579,In_862,In_834);
nand U2580 (N_2580,In_957,In_846);
and U2581 (N_2581,In_755,In_310);
and U2582 (N_2582,In_700,In_81);
nand U2583 (N_2583,In_125,In_740);
or U2584 (N_2584,In_748,In_778);
or U2585 (N_2585,In_350,In_640);
nand U2586 (N_2586,In_743,In_619);
nand U2587 (N_2587,In_645,In_816);
nor U2588 (N_2588,In_171,In_731);
and U2589 (N_2589,In_563,In_376);
nor U2590 (N_2590,In_219,In_325);
and U2591 (N_2591,In_501,In_120);
nand U2592 (N_2592,In_198,In_931);
and U2593 (N_2593,In_36,In_21);
nor U2594 (N_2594,In_484,In_630);
nand U2595 (N_2595,In_173,In_682);
xor U2596 (N_2596,In_163,In_408);
xor U2597 (N_2597,In_954,In_521);
or U2598 (N_2598,In_857,In_380);
or U2599 (N_2599,In_796,In_61);
nor U2600 (N_2600,In_725,In_871);
and U2601 (N_2601,In_887,In_714);
and U2602 (N_2602,In_517,In_591);
nand U2603 (N_2603,In_340,In_140);
xor U2604 (N_2604,In_395,In_271);
and U2605 (N_2605,In_596,In_369);
or U2606 (N_2606,In_453,In_998);
xor U2607 (N_2607,In_198,In_249);
nor U2608 (N_2608,In_406,In_594);
and U2609 (N_2609,In_636,In_11);
nand U2610 (N_2610,In_550,In_120);
xor U2611 (N_2611,In_101,In_577);
nand U2612 (N_2612,In_449,In_763);
and U2613 (N_2613,In_559,In_204);
xnor U2614 (N_2614,In_335,In_866);
and U2615 (N_2615,In_446,In_82);
or U2616 (N_2616,In_263,In_443);
nor U2617 (N_2617,In_218,In_55);
and U2618 (N_2618,In_995,In_98);
xnor U2619 (N_2619,In_652,In_90);
nor U2620 (N_2620,In_831,In_929);
xor U2621 (N_2621,In_92,In_103);
and U2622 (N_2622,In_571,In_578);
or U2623 (N_2623,In_156,In_405);
or U2624 (N_2624,In_792,In_305);
and U2625 (N_2625,In_73,In_547);
nor U2626 (N_2626,In_568,In_163);
xnor U2627 (N_2627,In_870,In_211);
and U2628 (N_2628,In_565,In_339);
xor U2629 (N_2629,In_868,In_5);
nor U2630 (N_2630,In_446,In_23);
nor U2631 (N_2631,In_147,In_827);
nand U2632 (N_2632,In_624,In_819);
and U2633 (N_2633,In_771,In_20);
and U2634 (N_2634,In_53,In_378);
nor U2635 (N_2635,In_139,In_324);
xor U2636 (N_2636,In_58,In_499);
and U2637 (N_2637,In_254,In_938);
nor U2638 (N_2638,In_967,In_144);
nand U2639 (N_2639,In_278,In_888);
and U2640 (N_2640,In_155,In_183);
or U2641 (N_2641,In_375,In_403);
nand U2642 (N_2642,In_714,In_896);
nand U2643 (N_2643,In_297,In_548);
xor U2644 (N_2644,In_779,In_828);
nor U2645 (N_2645,In_685,In_766);
nor U2646 (N_2646,In_197,In_732);
or U2647 (N_2647,In_110,In_525);
or U2648 (N_2648,In_626,In_547);
nand U2649 (N_2649,In_969,In_828);
nand U2650 (N_2650,In_567,In_467);
or U2651 (N_2651,In_995,In_148);
or U2652 (N_2652,In_672,In_511);
and U2653 (N_2653,In_724,In_527);
nand U2654 (N_2654,In_464,In_651);
xnor U2655 (N_2655,In_401,In_617);
nand U2656 (N_2656,In_476,In_426);
nand U2657 (N_2657,In_949,In_482);
nor U2658 (N_2658,In_448,In_307);
nand U2659 (N_2659,In_193,In_644);
xor U2660 (N_2660,In_232,In_977);
nand U2661 (N_2661,In_969,In_955);
xnor U2662 (N_2662,In_773,In_16);
and U2663 (N_2663,In_826,In_674);
or U2664 (N_2664,In_588,In_516);
or U2665 (N_2665,In_911,In_567);
xor U2666 (N_2666,In_411,In_797);
nand U2667 (N_2667,In_142,In_973);
or U2668 (N_2668,In_965,In_283);
nor U2669 (N_2669,In_326,In_325);
nor U2670 (N_2670,In_788,In_258);
or U2671 (N_2671,In_406,In_925);
nor U2672 (N_2672,In_394,In_435);
and U2673 (N_2673,In_174,In_87);
nor U2674 (N_2674,In_661,In_66);
or U2675 (N_2675,In_632,In_98);
xor U2676 (N_2676,In_836,In_171);
nor U2677 (N_2677,In_723,In_141);
or U2678 (N_2678,In_355,In_183);
and U2679 (N_2679,In_573,In_161);
or U2680 (N_2680,In_855,In_996);
xor U2681 (N_2681,In_687,In_36);
nand U2682 (N_2682,In_228,In_360);
and U2683 (N_2683,In_242,In_93);
or U2684 (N_2684,In_744,In_569);
and U2685 (N_2685,In_607,In_886);
nor U2686 (N_2686,In_383,In_936);
and U2687 (N_2687,In_895,In_734);
and U2688 (N_2688,In_490,In_282);
or U2689 (N_2689,In_122,In_266);
xnor U2690 (N_2690,In_38,In_494);
and U2691 (N_2691,In_442,In_924);
and U2692 (N_2692,In_687,In_992);
or U2693 (N_2693,In_636,In_238);
nor U2694 (N_2694,In_709,In_629);
nor U2695 (N_2695,In_370,In_711);
nor U2696 (N_2696,In_168,In_270);
and U2697 (N_2697,In_637,In_88);
nor U2698 (N_2698,In_429,In_157);
nand U2699 (N_2699,In_731,In_850);
nor U2700 (N_2700,In_86,In_965);
nor U2701 (N_2701,In_311,In_466);
nand U2702 (N_2702,In_64,In_239);
xnor U2703 (N_2703,In_888,In_435);
and U2704 (N_2704,In_605,In_166);
and U2705 (N_2705,In_305,In_275);
or U2706 (N_2706,In_788,In_274);
nor U2707 (N_2707,In_705,In_235);
nor U2708 (N_2708,In_410,In_572);
nor U2709 (N_2709,In_460,In_163);
nor U2710 (N_2710,In_260,In_372);
and U2711 (N_2711,In_363,In_568);
xnor U2712 (N_2712,In_542,In_420);
xnor U2713 (N_2713,In_238,In_800);
nand U2714 (N_2714,In_429,In_786);
nand U2715 (N_2715,In_439,In_450);
nor U2716 (N_2716,In_983,In_775);
and U2717 (N_2717,In_806,In_47);
or U2718 (N_2718,In_15,In_554);
or U2719 (N_2719,In_257,In_486);
xnor U2720 (N_2720,In_780,In_809);
nand U2721 (N_2721,In_113,In_277);
and U2722 (N_2722,In_801,In_844);
xnor U2723 (N_2723,In_349,In_953);
nor U2724 (N_2724,In_523,In_695);
nor U2725 (N_2725,In_658,In_834);
or U2726 (N_2726,In_954,In_121);
nor U2727 (N_2727,In_588,In_987);
and U2728 (N_2728,In_893,In_685);
nand U2729 (N_2729,In_112,In_95);
xor U2730 (N_2730,In_580,In_775);
xor U2731 (N_2731,In_7,In_93);
nand U2732 (N_2732,In_654,In_566);
nor U2733 (N_2733,In_877,In_205);
xnor U2734 (N_2734,In_716,In_408);
nand U2735 (N_2735,In_83,In_413);
nand U2736 (N_2736,In_521,In_359);
xnor U2737 (N_2737,In_819,In_968);
nor U2738 (N_2738,In_989,In_670);
and U2739 (N_2739,In_245,In_838);
and U2740 (N_2740,In_349,In_428);
xor U2741 (N_2741,In_940,In_685);
and U2742 (N_2742,In_887,In_89);
xor U2743 (N_2743,In_905,In_572);
or U2744 (N_2744,In_937,In_228);
and U2745 (N_2745,In_271,In_699);
and U2746 (N_2746,In_717,In_140);
and U2747 (N_2747,In_369,In_144);
nand U2748 (N_2748,In_850,In_894);
xnor U2749 (N_2749,In_722,In_229);
or U2750 (N_2750,In_49,In_201);
and U2751 (N_2751,In_81,In_701);
or U2752 (N_2752,In_409,In_86);
nor U2753 (N_2753,In_132,In_126);
xor U2754 (N_2754,In_4,In_193);
and U2755 (N_2755,In_887,In_83);
and U2756 (N_2756,In_665,In_729);
and U2757 (N_2757,In_944,In_155);
and U2758 (N_2758,In_544,In_255);
xor U2759 (N_2759,In_151,In_779);
or U2760 (N_2760,In_926,In_358);
nand U2761 (N_2761,In_433,In_109);
and U2762 (N_2762,In_952,In_185);
nor U2763 (N_2763,In_85,In_805);
nand U2764 (N_2764,In_121,In_760);
and U2765 (N_2765,In_376,In_73);
xnor U2766 (N_2766,In_602,In_781);
nand U2767 (N_2767,In_333,In_273);
or U2768 (N_2768,In_93,In_811);
xor U2769 (N_2769,In_23,In_156);
nand U2770 (N_2770,In_776,In_552);
nor U2771 (N_2771,In_18,In_295);
nor U2772 (N_2772,In_701,In_542);
xnor U2773 (N_2773,In_671,In_390);
nor U2774 (N_2774,In_322,In_646);
and U2775 (N_2775,In_554,In_456);
and U2776 (N_2776,In_364,In_990);
xor U2777 (N_2777,In_377,In_424);
nand U2778 (N_2778,In_918,In_292);
nand U2779 (N_2779,In_835,In_333);
nand U2780 (N_2780,In_910,In_449);
nand U2781 (N_2781,In_723,In_703);
nor U2782 (N_2782,In_645,In_672);
nor U2783 (N_2783,In_968,In_999);
or U2784 (N_2784,In_903,In_162);
or U2785 (N_2785,In_521,In_916);
nor U2786 (N_2786,In_164,In_147);
nand U2787 (N_2787,In_786,In_545);
and U2788 (N_2788,In_636,In_649);
nand U2789 (N_2789,In_293,In_594);
nor U2790 (N_2790,In_630,In_381);
and U2791 (N_2791,In_12,In_628);
nor U2792 (N_2792,In_626,In_481);
or U2793 (N_2793,In_992,In_95);
nor U2794 (N_2794,In_114,In_701);
xor U2795 (N_2795,In_477,In_245);
xnor U2796 (N_2796,In_88,In_108);
xnor U2797 (N_2797,In_873,In_827);
xor U2798 (N_2798,In_607,In_352);
or U2799 (N_2799,In_445,In_84);
nand U2800 (N_2800,In_1,In_568);
nor U2801 (N_2801,In_860,In_344);
nor U2802 (N_2802,In_660,In_526);
or U2803 (N_2803,In_123,In_679);
or U2804 (N_2804,In_532,In_518);
nand U2805 (N_2805,In_679,In_907);
and U2806 (N_2806,In_434,In_163);
or U2807 (N_2807,In_154,In_641);
nand U2808 (N_2808,In_53,In_854);
and U2809 (N_2809,In_546,In_830);
xnor U2810 (N_2810,In_245,In_194);
xor U2811 (N_2811,In_262,In_702);
nor U2812 (N_2812,In_402,In_642);
and U2813 (N_2813,In_479,In_332);
or U2814 (N_2814,In_742,In_281);
nor U2815 (N_2815,In_80,In_204);
and U2816 (N_2816,In_354,In_92);
xor U2817 (N_2817,In_417,In_682);
nand U2818 (N_2818,In_924,In_658);
or U2819 (N_2819,In_751,In_741);
and U2820 (N_2820,In_420,In_165);
nor U2821 (N_2821,In_108,In_495);
or U2822 (N_2822,In_652,In_332);
xor U2823 (N_2823,In_237,In_579);
xnor U2824 (N_2824,In_426,In_341);
xnor U2825 (N_2825,In_280,In_609);
and U2826 (N_2826,In_197,In_100);
nor U2827 (N_2827,In_149,In_387);
nand U2828 (N_2828,In_344,In_100);
or U2829 (N_2829,In_482,In_849);
nand U2830 (N_2830,In_632,In_449);
xor U2831 (N_2831,In_204,In_59);
nand U2832 (N_2832,In_134,In_616);
and U2833 (N_2833,In_150,In_531);
xor U2834 (N_2834,In_367,In_369);
or U2835 (N_2835,In_947,In_140);
nand U2836 (N_2836,In_691,In_532);
or U2837 (N_2837,In_937,In_496);
and U2838 (N_2838,In_926,In_183);
nor U2839 (N_2839,In_62,In_807);
nor U2840 (N_2840,In_95,In_625);
nand U2841 (N_2841,In_592,In_613);
and U2842 (N_2842,In_682,In_197);
and U2843 (N_2843,In_559,In_784);
nor U2844 (N_2844,In_693,In_687);
and U2845 (N_2845,In_847,In_89);
or U2846 (N_2846,In_922,In_604);
or U2847 (N_2847,In_451,In_267);
or U2848 (N_2848,In_117,In_621);
or U2849 (N_2849,In_483,In_19);
nand U2850 (N_2850,In_929,In_663);
xnor U2851 (N_2851,In_551,In_866);
xor U2852 (N_2852,In_721,In_682);
xor U2853 (N_2853,In_710,In_11);
xor U2854 (N_2854,In_730,In_526);
nand U2855 (N_2855,In_675,In_392);
xor U2856 (N_2856,In_52,In_792);
nor U2857 (N_2857,In_177,In_227);
nor U2858 (N_2858,In_199,In_709);
and U2859 (N_2859,In_40,In_523);
nor U2860 (N_2860,In_482,In_998);
and U2861 (N_2861,In_241,In_902);
or U2862 (N_2862,In_993,In_398);
and U2863 (N_2863,In_445,In_880);
xor U2864 (N_2864,In_40,In_582);
or U2865 (N_2865,In_945,In_686);
xor U2866 (N_2866,In_860,In_257);
nor U2867 (N_2867,In_984,In_492);
or U2868 (N_2868,In_985,In_488);
or U2869 (N_2869,In_140,In_157);
or U2870 (N_2870,In_532,In_668);
or U2871 (N_2871,In_1,In_266);
nor U2872 (N_2872,In_738,In_252);
or U2873 (N_2873,In_109,In_533);
or U2874 (N_2874,In_493,In_759);
nand U2875 (N_2875,In_200,In_932);
or U2876 (N_2876,In_81,In_424);
nor U2877 (N_2877,In_568,In_753);
xor U2878 (N_2878,In_486,In_862);
or U2879 (N_2879,In_836,In_485);
and U2880 (N_2880,In_913,In_229);
nand U2881 (N_2881,In_363,In_567);
nand U2882 (N_2882,In_770,In_620);
xor U2883 (N_2883,In_296,In_5);
xnor U2884 (N_2884,In_824,In_559);
xnor U2885 (N_2885,In_945,In_678);
or U2886 (N_2886,In_216,In_480);
nor U2887 (N_2887,In_905,In_809);
or U2888 (N_2888,In_125,In_280);
nor U2889 (N_2889,In_795,In_261);
and U2890 (N_2890,In_150,In_216);
nor U2891 (N_2891,In_832,In_979);
and U2892 (N_2892,In_438,In_140);
nor U2893 (N_2893,In_462,In_766);
nor U2894 (N_2894,In_613,In_591);
and U2895 (N_2895,In_33,In_395);
xor U2896 (N_2896,In_66,In_74);
or U2897 (N_2897,In_524,In_917);
xor U2898 (N_2898,In_419,In_76);
xnor U2899 (N_2899,In_362,In_20);
xnor U2900 (N_2900,In_662,In_603);
nand U2901 (N_2901,In_946,In_995);
nand U2902 (N_2902,In_348,In_410);
xnor U2903 (N_2903,In_975,In_192);
nand U2904 (N_2904,In_906,In_103);
nor U2905 (N_2905,In_883,In_59);
nand U2906 (N_2906,In_372,In_972);
or U2907 (N_2907,In_575,In_232);
nand U2908 (N_2908,In_544,In_182);
and U2909 (N_2909,In_962,In_267);
xor U2910 (N_2910,In_759,In_358);
xor U2911 (N_2911,In_364,In_586);
nand U2912 (N_2912,In_494,In_800);
or U2913 (N_2913,In_801,In_898);
nand U2914 (N_2914,In_65,In_582);
and U2915 (N_2915,In_863,In_121);
or U2916 (N_2916,In_521,In_847);
xor U2917 (N_2917,In_265,In_782);
xnor U2918 (N_2918,In_295,In_221);
and U2919 (N_2919,In_678,In_601);
nor U2920 (N_2920,In_869,In_546);
nor U2921 (N_2921,In_762,In_223);
and U2922 (N_2922,In_624,In_540);
nand U2923 (N_2923,In_533,In_571);
and U2924 (N_2924,In_629,In_2);
nand U2925 (N_2925,In_830,In_563);
and U2926 (N_2926,In_565,In_280);
or U2927 (N_2927,In_523,In_60);
and U2928 (N_2928,In_636,In_257);
nand U2929 (N_2929,In_322,In_69);
nor U2930 (N_2930,In_101,In_947);
nor U2931 (N_2931,In_593,In_961);
nand U2932 (N_2932,In_824,In_188);
nand U2933 (N_2933,In_351,In_354);
nor U2934 (N_2934,In_713,In_736);
nand U2935 (N_2935,In_671,In_182);
nand U2936 (N_2936,In_429,In_259);
and U2937 (N_2937,In_156,In_510);
or U2938 (N_2938,In_256,In_691);
nor U2939 (N_2939,In_709,In_487);
nor U2940 (N_2940,In_29,In_228);
and U2941 (N_2941,In_671,In_533);
xnor U2942 (N_2942,In_120,In_428);
or U2943 (N_2943,In_847,In_749);
nor U2944 (N_2944,In_935,In_604);
nand U2945 (N_2945,In_102,In_227);
and U2946 (N_2946,In_892,In_278);
xnor U2947 (N_2947,In_97,In_886);
or U2948 (N_2948,In_272,In_650);
and U2949 (N_2949,In_55,In_495);
or U2950 (N_2950,In_991,In_940);
or U2951 (N_2951,In_710,In_656);
nor U2952 (N_2952,In_529,In_214);
or U2953 (N_2953,In_404,In_417);
xnor U2954 (N_2954,In_403,In_333);
or U2955 (N_2955,In_422,In_383);
and U2956 (N_2956,In_166,In_756);
nor U2957 (N_2957,In_424,In_43);
or U2958 (N_2958,In_652,In_542);
xor U2959 (N_2959,In_355,In_342);
and U2960 (N_2960,In_737,In_141);
nor U2961 (N_2961,In_908,In_903);
and U2962 (N_2962,In_802,In_875);
nand U2963 (N_2963,In_143,In_222);
nand U2964 (N_2964,In_951,In_505);
nor U2965 (N_2965,In_358,In_224);
nand U2966 (N_2966,In_970,In_512);
xnor U2967 (N_2967,In_573,In_348);
and U2968 (N_2968,In_310,In_398);
nor U2969 (N_2969,In_114,In_240);
xnor U2970 (N_2970,In_569,In_852);
xnor U2971 (N_2971,In_473,In_802);
and U2972 (N_2972,In_994,In_388);
or U2973 (N_2973,In_133,In_590);
nor U2974 (N_2974,In_298,In_413);
and U2975 (N_2975,In_333,In_851);
and U2976 (N_2976,In_576,In_20);
xor U2977 (N_2977,In_832,In_887);
or U2978 (N_2978,In_785,In_514);
and U2979 (N_2979,In_320,In_416);
nand U2980 (N_2980,In_104,In_483);
nor U2981 (N_2981,In_651,In_788);
nand U2982 (N_2982,In_846,In_993);
nor U2983 (N_2983,In_436,In_939);
xnor U2984 (N_2984,In_999,In_179);
or U2985 (N_2985,In_563,In_241);
nor U2986 (N_2986,In_837,In_255);
xor U2987 (N_2987,In_72,In_858);
nand U2988 (N_2988,In_201,In_21);
or U2989 (N_2989,In_209,In_900);
or U2990 (N_2990,In_726,In_715);
nor U2991 (N_2991,In_990,In_444);
nand U2992 (N_2992,In_183,In_689);
nor U2993 (N_2993,In_225,In_10);
and U2994 (N_2994,In_200,In_432);
nor U2995 (N_2995,In_577,In_653);
xor U2996 (N_2996,In_735,In_844);
and U2997 (N_2997,In_408,In_260);
and U2998 (N_2998,In_685,In_293);
nor U2999 (N_2999,In_51,In_137);
nor U3000 (N_3000,In_647,In_518);
and U3001 (N_3001,In_170,In_488);
nand U3002 (N_3002,In_969,In_124);
nor U3003 (N_3003,In_922,In_711);
nand U3004 (N_3004,In_804,In_60);
nand U3005 (N_3005,In_553,In_954);
nor U3006 (N_3006,In_717,In_970);
nor U3007 (N_3007,In_533,In_270);
nor U3008 (N_3008,In_795,In_347);
xor U3009 (N_3009,In_418,In_270);
or U3010 (N_3010,In_102,In_379);
and U3011 (N_3011,In_510,In_513);
nor U3012 (N_3012,In_150,In_199);
and U3013 (N_3013,In_127,In_741);
nor U3014 (N_3014,In_867,In_791);
nand U3015 (N_3015,In_437,In_454);
and U3016 (N_3016,In_867,In_142);
nand U3017 (N_3017,In_701,In_123);
xor U3018 (N_3018,In_507,In_178);
nor U3019 (N_3019,In_362,In_805);
or U3020 (N_3020,In_346,In_437);
xor U3021 (N_3021,In_111,In_713);
xnor U3022 (N_3022,In_539,In_267);
and U3023 (N_3023,In_880,In_365);
or U3024 (N_3024,In_688,In_121);
or U3025 (N_3025,In_464,In_69);
nor U3026 (N_3026,In_210,In_879);
and U3027 (N_3027,In_16,In_406);
xor U3028 (N_3028,In_956,In_880);
xnor U3029 (N_3029,In_197,In_948);
and U3030 (N_3030,In_277,In_609);
or U3031 (N_3031,In_408,In_458);
nand U3032 (N_3032,In_259,In_807);
nand U3033 (N_3033,In_332,In_612);
xor U3034 (N_3034,In_930,In_47);
xnor U3035 (N_3035,In_813,In_632);
xnor U3036 (N_3036,In_608,In_532);
or U3037 (N_3037,In_396,In_475);
nand U3038 (N_3038,In_154,In_325);
and U3039 (N_3039,In_60,In_532);
and U3040 (N_3040,In_321,In_278);
and U3041 (N_3041,In_23,In_576);
and U3042 (N_3042,In_866,In_752);
and U3043 (N_3043,In_376,In_1);
or U3044 (N_3044,In_898,In_593);
nor U3045 (N_3045,In_679,In_713);
and U3046 (N_3046,In_177,In_452);
xor U3047 (N_3047,In_493,In_998);
nor U3048 (N_3048,In_94,In_647);
nor U3049 (N_3049,In_607,In_902);
and U3050 (N_3050,In_968,In_565);
xnor U3051 (N_3051,In_487,In_960);
nor U3052 (N_3052,In_934,In_331);
nor U3053 (N_3053,In_413,In_191);
nand U3054 (N_3054,In_341,In_409);
xnor U3055 (N_3055,In_589,In_474);
xnor U3056 (N_3056,In_174,In_896);
nand U3057 (N_3057,In_200,In_557);
xor U3058 (N_3058,In_225,In_763);
xor U3059 (N_3059,In_427,In_226);
nor U3060 (N_3060,In_430,In_549);
and U3061 (N_3061,In_210,In_320);
and U3062 (N_3062,In_355,In_85);
xnor U3063 (N_3063,In_243,In_597);
nand U3064 (N_3064,In_519,In_692);
xnor U3065 (N_3065,In_341,In_588);
nor U3066 (N_3066,In_976,In_421);
nor U3067 (N_3067,In_804,In_189);
xnor U3068 (N_3068,In_213,In_312);
or U3069 (N_3069,In_851,In_168);
nor U3070 (N_3070,In_343,In_714);
and U3071 (N_3071,In_469,In_196);
and U3072 (N_3072,In_912,In_468);
or U3073 (N_3073,In_277,In_711);
or U3074 (N_3074,In_684,In_318);
xor U3075 (N_3075,In_764,In_376);
nand U3076 (N_3076,In_934,In_551);
and U3077 (N_3077,In_137,In_777);
nand U3078 (N_3078,In_837,In_638);
or U3079 (N_3079,In_463,In_175);
nor U3080 (N_3080,In_212,In_563);
nor U3081 (N_3081,In_553,In_711);
and U3082 (N_3082,In_737,In_281);
and U3083 (N_3083,In_943,In_477);
xor U3084 (N_3084,In_493,In_930);
and U3085 (N_3085,In_837,In_623);
or U3086 (N_3086,In_518,In_394);
nor U3087 (N_3087,In_607,In_453);
nand U3088 (N_3088,In_625,In_954);
and U3089 (N_3089,In_18,In_881);
and U3090 (N_3090,In_919,In_607);
xnor U3091 (N_3091,In_883,In_479);
xor U3092 (N_3092,In_105,In_40);
nand U3093 (N_3093,In_40,In_205);
or U3094 (N_3094,In_313,In_193);
or U3095 (N_3095,In_434,In_638);
nor U3096 (N_3096,In_512,In_439);
and U3097 (N_3097,In_185,In_276);
nand U3098 (N_3098,In_829,In_389);
or U3099 (N_3099,In_350,In_414);
and U3100 (N_3100,In_832,In_624);
and U3101 (N_3101,In_516,In_171);
nor U3102 (N_3102,In_6,In_799);
nor U3103 (N_3103,In_281,In_836);
and U3104 (N_3104,In_602,In_363);
or U3105 (N_3105,In_563,In_405);
and U3106 (N_3106,In_283,In_903);
or U3107 (N_3107,In_483,In_529);
nor U3108 (N_3108,In_61,In_993);
xnor U3109 (N_3109,In_826,In_440);
xor U3110 (N_3110,In_996,In_776);
nor U3111 (N_3111,In_943,In_230);
xnor U3112 (N_3112,In_456,In_164);
xor U3113 (N_3113,In_747,In_518);
nor U3114 (N_3114,In_522,In_825);
and U3115 (N_3115,In_264,In_590);
xor U3116 (N_3116,In_328,In_766);
xnor U3117 (N_3117,In_477,In_818);
nor U3118 (N_3118,In_718,In_226);
nand U3119 (N_3119,In_265,In_482);
nand U3120 (N_3120,In_65,In_773);
nand U3121 (N_3121,In_120,In_777);
xnor U3122 (N_3122,In_384,In_108);
or U3123 (N_3123,In_515,In_244);
nand U3124 (N_3124,In_239,In_856);
and U3125 (N_3125,In_23,In_41);
and U3126 (N_3126,In_192,In_196);
or U3127 (N_3127,In_297,In_478);
and U3128 (N_3128,In_522,In_191);
xnor U3129 (N_3129,In_537,In_500);
and U3130 (N_3130,In_516,In_241);
nand U3131 (N_3131,In_318,In_160);
nor U3132 (N_3132,In_442,In_279);
or U3133 (N_3133,In_697,In_689);
or U3134 (N_3134,In_208,In_485);
xnor U3135 (N_3135,In_495,In_852);
nand U3136 (N_3136,In_917,In_757);
and U3137 (N_3137,In_132,In_539);
and U3138 (N_3138,In_103,In_143);
or U3139 (N_3139,In_950,In_328);
nor U3140 (N_3140,In_204,In_39);
xor U3141 (N_3141,In_586,In_662);
and U3142 (N_3142,In_954,In_336);
nand U3143 (N_3143,In_762,In_900);
xor U3144 (N_3144,In_654,In_364);
or U3145 (N_3145,In_5,In_513);
and U3146 (N_3146,In_348,In_977);
xnor U3147 (N_3147,In_161,In_520);
xor U3148 (N_3148,In_859,In_496);
nand U3149 (N_3149,In_627,In_640);
xor U3150 (N_3150,In_287,In_647);
nand U3151 (N_3151,In_59,In_546);
nand U3152 (N_3152,In_703,In_255);
and U3153 (N_3153,In_109,In_409);
nand U3154 (N_3154,In_733,In_17);
and U3155 (N_3155,In_393,In_763);
nand U3156 (N_3156,In_524,In_640);
nor U3157 (N_3157,In_582,In_45);
and U3158 (N_3158,In_620,In_127);
or U3159 (N_3159,In_985,In_573);
xor U3160 (N_3160,In_371,In_150);
or U3161 (N_3161,In_163,In_731);
nand U3162 (N_3162,In_369,In_901);
or U3163 (N_3163,In_582,In_328);
nor U3164 (N_3164,In_931,In_541);
and U3165 (N_3165,In_150,In_970);
and U3166 (N_3166,In_89,In_524);
or U3167 (N_3167,In_676,In_458);
or U3168 (N_3168,In_519,In_525);
nor U3169 (N_3169,In_973,In_731);
xnor U3170 (N_3170,In_97,In_981);
nand U3171 (N_3171,In_564,In_412);
xnor U3172 (N_3172,In_237,In_724);
xor U3173 (N_3173,In_271,In_626);
nor U3174 (N_3174,In_973,In_195);
nand U3175 (N_3175,In_915,In_300);
nor U3176 (N_3176,In_125,In_298);
or U3177 (N_3177,In_5,In_786);
and U3178 (N_3178,In_579,In_13);
xnor U3179 (N_3179,In_152,In_877);
nor U3180 (N_3180,In_488,In_960);
or U3181 (N_3181,In_217,In_944);
or U3182 (N_3182,In_655,In_630);
nor U3183 (N_3183,In_240,In_434);
and U3184 (N_3184,In_109,In_247);
nor U3185 (N_3185,In_450,In_493);
nand U3186 (N_3186,In_957,In_585);
nand U3187 (N_3187,In_95,In_235);
xor U3188 (N_3188,In_201,In_335);
or U3189 (N_3189,In_64,In_997);
or U3190 (N_3190,In_814,In_765);
and U3191 (N_3191,In_261,In_696);
xnor U3192 (N_3192,In_368,In_691);
nor U3193 (N_3193,In_615,In_494);
nand U3194 (N_3194,In_945,In_987);
and U3195 (N_3195,In_942,In_436);
nor U3196 (N_3196,In_783,In_475);
and U3197 (N_3197,In_667,In_989);
and U3198 (N_3198,In_405,In_999);
or U3199 (N_3199,In_738,In_969);
nor U3200 (N_3200,In_3,In_13);
or U3201 (N_3201,In_359,In_803);
nor U3202 (N_3202,In_793,In_794);
or U3203 (N_3203,In_403,In_925);
or U3204 (N_3204,In_368,In_478);
and U3205 (N_3205,In_503,In_862);
and U3206 (N_3206,In_83,In_546);
xor U3207 (N_3207,In_510,In_604);
nand U3208 (N_3208,In_924,In_565);
nand U3209 (N_3209,In_777,In_5);
xor U3210 (N_3210,In_243,In_361);
and U3211 (N_3211,In_720,In_94);
and U3212 (N_3212,In_394,In_922);
nand U3213 (N_3213,In_53,In_956);
or U3214 (N_3214,In_432,In_622);
and U3215 (N_3215,In_169,In_54);
nand U3216 (N_3216,In_433,In_662);
nand U3217 (N_3217,In_369,In_879);
nand U3218 (N_3218,In_364,In_701);
or U3219 (N_3219,In_903,In_854);
xnor U3220 (N_3220,In_684,In_686);
xnor U3221 (N_3221,In_117,In_523);
and U3222 (N_3222,In_913,In_416);
nand U3223 (N_3223,In_161,In_920);
and U3224 (N_3224,In_303,In_19);
nand U3225 (N_3225,In_483,In_532);
nand U3226 (N_3226,In_258,In_799);
nor U3227 (N_3227,In_694,In_886);
nand U3228 (N_3228,In_371,In_934);
nor U3229 (N_3229,In_323,In_201);
or U3230 (N_3230,In_718,In_937);
nand U3231 (N_3231,In_523,In_990);
and U3232 (N_3232,In_837,In_717);
nor U3233 (N_3233,In_331,In_192);
nand U3234 (N_3234,In_120,In_190);
and U3235 (N_3235,In_832,In_694);
xnor U3236 (N_3236,In_511,In_829);
or U3237 (N_3237,In_884,In_433);
and U3238 (N_3238,In_740,In_49);
or U3239 (N_3239,In_662,In_716);
and U3240 (N_3240,In_224,In_238);
xor U3241 (N_3241,In_182,In_494);
nor U3242 (N_3242,In_121,In_735);
nand U3243 (N_3243,In_803,In_654);
nor U3244 (N_3244,In_317,In_337);
nand U3245 (N_3245,In_339,In_919);
or U3246 (N_3246,In_674,In_524);
or U3247 (N_3247,In_442,In_440);
nand U3248 (N_3248,In_307,In_722);
nor U3249 (N_3249,In_860,In_959);
nor U3250 (N_3250,In_393,In_877);
and U3251 (N_3251,In_515,In_935);
nor U3252 (N_3252,In_466,In_377);
nand U3253 (N_3253,In_867,In_409);
nor U3254 (N_3254,In_211,In_561);
nor U3255 (N_3255,In_616,In_225);
xor U3256 (N_3256,In_367,In_24);
nand U3257 (N_3257,In_978,In_554);
nand U3258 (N_3258,In_500,In_461);
xor U3259 (N_3259,In_293,In_678);
xor U3260 (N_3260,In_222,In_362);
or U3261 (N_3261,In_558,In_82);
xor U3262 (N_3262,In_767,In_299);
and U3263 (N_3263,In_737,In_681);
nor U3264 (N_3264,In_877,In_457);
nand U3265 (N_3265,In_734,In_5);
nor U3266 (N_3266,In_748,In_765);
xor U3267 (N_3267,In_132,In_803);
nor U3268 (N_3268,In_444,In_677);
and U3269 (N_3269,In_394,In_86);
nor U3270 (N_3270,In_728,In_79);
xnor U3271 (N_3271,In_949,In_645);
nor U3272 (N_3272,In_673,In_386);
and U3273 (N_3273,In_915,In_708);
nand U3274 (N_3274,In_201,In_8);
xor U3275 (N_3275,In_32,In_571);
and U3276 (N_3276,In_373,In_905);
nand U3277 (N_3277,In_960,In_579);
or U3278 (N_3278,In_39,In_206);
xor U3279 (N_3279,In_810,In_517);
xor U3280 (N_3280,In_829,In_771);
and U3281 (N_3281,In_6,In_998);
nand U3282 (N_3282,In_489,In_406);
or U3283 (N_3283,In_230,In_65);
xnor U3284 (N_3284,In_487,In_92);
or U3285 (N_3285,In_685,In_983);
or U3286 (N_3286,In_886,In_379);
nor U3287 (N_3287,In_298,In_533);
xor U3288 (N_3288,In_363,In_90);
or U3289 (N_3289,In_490,In_641);
or U3290 (N_3290,In_39,In_366);
xor U3291 (N_3291,In_937,In_780);
nor U3292 (N_3292,In_393,In_898);
xor U3293 (N_3293,In_877,In_214);
nand U3294 (N_3294,In_171,In_443);
xor U3295 (N_3295,In_239,In_551);
nor U3296 (N_3296,In_448,In_923);
nand U3297 (N_3297,In_341,In_312);
and U3298 (N_3298,In_467,In_961);
nor U3299 (N_3299,In_266,In_441);
nor U3300 (N_3300,In_551,In_884);
and U3301 (N_3301,In_505,In_636);
xor U3302 (N_3302,In_131,In_620);
or U3303 (N_3303,In_286,In_656);
xnor U3304 (N_3304,In_704,In_990);
and U3305 (N_3305,In_915,In_692);
nand U3306 (N_3306,In_901,In_689);
nand U3307 (N_3307,In_23,In_790);
and U3308 (N_3308,In_54,In_1);
xnor U3309 (N_3309,In_516,In_879);
or U3310 (N_3310,In_56,In_62);
or U3311 (N_3311,In_360,In_623);
nand U3312 (N_3312,In_652,In_491);
nor U3313 (N_3313,In_266,In_907);
xnor U3314 (N_3314,In_303,In_379);
xnor U3315 (N_3315,In_166,In_416);
nor U3316 (N_3316,In_176,In_893);
nand U3317 (N_3317,In_214,In_223);
nand U3318 (N_3318,In_130,In_853);
and U3319 (N_3319,In_539,In_297);
or U3320 (N_3320,In_376,In_520);
and U3321 (N_3321,In_645,In_812);
or U3322 (N_3322,In_502,In_935);
nor U3323 (N_3323,In_77,In_634);
xor U3324 (N_3324,In_517,In_460);
nor U3325 (N_3325,In_730,In_770);
and U3326 (N_3326,In_681,In_220);
nand U3327 (N_3327,In_197,In_877);
and U3328 (N_3328,In_422,In_601);
and U3329 (N_3329,In_956,In_461);
nor U3330 (N_3330,In_614,In_229);
nor U3331 (N_3331,In_42,In_865);
or U3332 (N_3332,In_614,In_820);
nand U3333 (N_3333,In_868,In_854);
and U3334 (N_3334,In_803,In_787);
and U3335 (N_3335,In_599,In_357);
and U3336 (N_3336,In_644,In_424);
nand U3337 (N_3337,In_341,In_929);
xnor U3338 (N_3338,In_544,In_713);
nor U3339 (N_3339,In_941,In_273);
nor U3340 (N_3340,In_768,In_247);
nor U3341 (N_3341,In_990,In_828);
nand U3342 (N_3342,In_73,In_730);
and U3343 (N_3343,In_96,In_14);
xor U3344 (N_3344,In_261,In_145);
or U3345 (N_3345,In_288,In_688);
and U3346 (N_3346,In_742,In_829);
and U3347 (N_3347,In_887,In_531);
or U3348 (N_3348,In_260,In_232);
or U3349 (N_3349,In_501,In_526);
nor U3350 (N_3350,In_3,In_504);
nand U3351 (N_3351,In_818,In_544);
or U3352 (N_3352,In_794,In_738);
nand U3353 (N_3353,In_677,In_16);
or U3354 (N_3354,In_580,In_215);
xnor U3355 (N_3355,In_419,In_772);
and U3356 (N_3356,In_615,In_324);
nand U3357 (N_3357,In_365,In_782);
and U3358 (N_3358,In_539,In_957);
or U3359 (N_3359,In_533,In_1);
nor U3360 (N_3360,In_860,In_791);
or U3361 (N_3361,In_868,In_607);
or U3362 (N_3362,In_330,In_97);
xnor U3363 (N_3363,In_928,In_588);
xnor U3364 (N_3364,In_181,In_622);
xor U3365 (N_3365,In_688,In_509);
or U3366 (N_3366,In_165,In_992);
and U3367 (N_3367,In_54,In_993);
xor U3368 (N_3368,In_247,In_759);
xnor U3369 (N_3369,In_873,In_139);
and U3370 (N_3370,In_944,In_935);
xnor U3371 (N_3371,In_743,In_315);
nand U3372 (N_3372,In_929,In_881);
nor U3373 (N_3373,In_596,In_431);
or U3374 (N_3374,In_991,In_879);
nand U3375 (N_3375,In_969,In_623);
nor U3376 (N_3376,In_321,In_935);
xnor U3377 (N_3377,In_398,In_38);
and U3378 (N_3378,In_543,In_801);
nor U3379 (N_3379,In_818,In_995);
nand U3380 (N_3380,In_232,In_16);
nor U3381 (N_3381,In_614,In_728);
xor U3382 (N_3382,In_709,In_68);
nand U3383 (N_3383,In_122,In_781);
or U3384 (N_3384,In_529,In_487);
nor U3385 (N_3385,In_708,In_711);
or U3386 (N_3386,In_864,In_220);
and U3387 (N_3387,In_722,In_919);
or U3388 (N_3388,In_348,In_587);
xor U3389 (N_3389,In_313,In_688);
nor U3390 (N_3390,In_722,In_765);
nor U3391 (N_3391,In_247,In_64);
nand U3392 (N_3392,In_130,In_892);
and U3393 (N_3393,In_371,In_568);
or U3394 (N_3394,In_946,In_731);
or U3395 (N_3395,In_698,In_194);
xor U3396 (N_3396,In_737,In_961);
nand U3397 (N_3397,In_8,In_681);
or U3398 (N_3398,In_200,In_533);
or U3399 (N_3399,In_358,In_860);
nand U3400 (N_3400,In_416,In_235);
or U3401 (N_3401,In_817,In_440);
nor U3402 (N_3402,In_433,In_791);
nor U3403 (N_3403,In_558,In_465);
and U3404 (N_3404,In_407,In_889);
and U3405 (N_3405,In_726,In_785);
nor U3406 (N_3406,In_779,In_457);
or U3407 (N_3407,In_611,In_569);
nor U3408 (N_3408,In_667,In_692);
xor U3409 (N_3409,In_304,In_186);
nand U3410 (N_3410,In_555,In_108);
or U3411 (N_3411,In_661,In_866);
nor U3412 (N_3412,In_811,In_392);
nor U3413 (N_3413,In_772,In_776);
xor U3414 (N_3414,In_192,In_267);
and U3415 (N_3415,In_415,In_18);
and U3416 (N_3416,In_557,In_171);
nand U3417 (N_3417,In_388,In_631);
nor U3418 (N_3418,In_731,In_963);
and U3419 (N_3419,In_953,In_625);
xnor U3420 (N_3420,In_624,In_625);
or U3421 (N_3421,In_176,In_726);
and U3422 (N_3422,In_194,In_966);
xor U3423 (N_3423,In_41,In_705);
nor U3424 (N_3424,In_917,In_514);
and U3425 (N_3425,In_621,In_959);
xnor U3426 (N_3426,In_857,In_628);
nand U3427 (N_3427,In_146,In_748);
nand U3428 (N_3428,In_353,In_570);
xnor U3429 (N_3429,In_187,In_667);
and U3430 (N_3430,In_821,In_16);
xor U3431 (N_3431,In_304,In_778);
xor U3432 (N_3432,In_540,In_227);
and U3433 (N_3433,In_80,In_479);
or U3434 (N_3434,In_180,In_562);
or U3435 (N_3435,In_62,In_215);
nand U3436 (N_3436,In_63,In_611);
or U3437 (N_3437,In_983,In_151);
nor U3438 (N_3438,In_841,In_814);
and U3439 (N_3439,In_917,In_47);
xor U3440 (N_3440,In_366,In_747);
or U3441 (N_3441,In_30,In_657);
nor U3442 (N_3442,In_544,In_306);
nor U3443 (N_3443,In_382,In_794);
or U3444 (N_3444,In_445,In_334);
or U3445 (N_3445,In_884,In_390);
xor U3446 (N_3446,In_599,In_565);
and U3447 (N_3447,In_950,In_256);
or U3448 (N_3448,In_605,In_94);
nor U3449 (N_3449,In_782,In_153);
nor U3450 (N_3450,In_938,In_916);
or U3451 (N_3451,In_84,In_679);
and U3452 (N_3452,In_685,In_212);
nor U3453 (N_3453,In_51,In_191);
nand U3454 (N_3454,In_219,In_840);
nor U3455 (N_3455,In_657,In_176);
nand U3456 (N_3456,In_66,In_558);
nand U3457 (N_3457,In_256,In_969);
nor U3458 (N_3458,In_779,In_128);
nand U3459 (N_3459,In_218,In_959);
and U3460 (N_3460,In_930,In_405);
xor U3461 (N_3461,In_767,In_812);
or U3462 (N_3462,In_201,In_412);
nand U3463 (N_3463,In_845,In_780);
and U3464 (N_3464,In_95,In_716);
and U3465 (N_3465,In_386,In_732);
xor U3466 (N_3466,In_584,In_283);
nor U3467 (N_3467,In_82,In_447);
or U3468 (N_3468,In_49,In_373);
or U3469 (N_3469,In_456,In_742);
and U3470 (N_3470,In_902,In_596);
and U3471 (N_3471,In_260,In_519);
nor U3472 (N_3472,In_683,In_742);
and U3473 (N_3473,In_480,In_347);
and U3474 (N_3474,In_770,In_68);
xor U3475 (N_3475,In_638,In_641);
nand U3476 (N_3476,In_544,In_998);
nor U3477 (N_3477,In_175,In_381);
or U3478 (N_3478,In_770,In_741);
nor U3479 (N_3479,In_282,In_900);
nor U3480 (N_3480,In_405,In_455);
or U3481 (N_3481,In_378,In_381);
xnor U3482 (N_3482,In_712,In_792);
nand U3483 (N_3483,In_506,In_577);
xnor U3484 (N_3484,In_199,In_431);
or U3485 (N_3485,In_633,In_367);
nand U3486 (N_3486,In_281,In_678);
or U3487 (N_3487,In_619,In_289);
nand U3488 (N_3488,In_858,In_441);
or U3489 (N_3489,In_994,In_644);
nand U3490 (N_3490,In_682,In_897);
nor U3491 (N_3491,In_387,In_799);
or U3492 (N_3492,In_847,In_615);
nand U3493 (N_3493,In_263,In_98);
and U3494 (N_3494,In_770,In_609);
nor U3495 (N_3495,In_838,In_566);
xor U3496 (N_3496,In_675,In_816);
nand U3497 (N_3497,In_212,In_294);
nand U3498 (N_3498,In_933,In_341);
and U3499 (N_3499,In_671,In_273);
and U3500 (N_3500,In_853,In_330);
nand U3501 (N_3501,In_333,In_736);
or U3502 (N_3502,In_278,In_19);
xnor U3503 (N_3503,In_803,In_201);
or U3504 (N_3504,In_355,In_923);
nand U3505 (N_3505,In_177,In_224);
xor U3506 (N_3506,In_417,In_315);
or U3507 (N_3507,In_475,In_96);
or U3508 (N_3508,In_330,In_433);
or U3509 (N_3509,In_250,In_986);
or U3510 (N_3510,In_670,In_109);
nor U3511 (N_3511,In_62,In_242);
and U3512 (N_3512,In_222,In_241);
xnor U3513 (N_3513,In_967,In_264);
nor U3514 (N_3514,In_131,In_165);
and U3515 (N_3515,In_107,In_337);
xor U3516 (N_3516,In_175,In_140);
and U3517 (N_3517,In_80,In_801);
and U3518 (N_3518,In_792,In_105);
nand U3519 (N_3519,In_549,In_410);
and U3520 (N_3520,In_884,In_836);
xor U3521 (N_3521,In_896,In_555);
nand U3522 (N_3522,In_277,In_117);
xor U3523 (N_3523,In_800,In_704);
or U3524 (N_3524,In_738,In_156);
or U3525 (N_3525,In_642,In_948);
xor U3526 (N_3526,In_160,In_217);
and U3527 (N_3527,In_101,In_471);
nand U3528 (N_3528,In_83,In_990);
and U3529 (N_3529,In_365,In_952);
nand U3530 (N_3530,In_920,In_923);
nand U3531 (N_3531,In_109,In_327);
and U3532 (N_3532,In_545,In_238);
nand U3533 (N_3533,In_350,In_478);
and U3534 (N_3534,In_766,In_560);
nor U3535 (N_3535,In_19,In_288);
and U3536 (N_3536,In_594,In_500);
or U3537 (N_3537,In_36,In_7);
or U3538 (N_3538,In_523,In_859);
nand U3539 (N_3539,In_491,In_388);
nand U3540 (N_3540,In_72,In_743);
or U3541 (N_3541,In_894,In_426);
nor U3542 (N_3542,In_123,In_651);
or U3543 (N_3543,In_419,In_867);
nor U3544 (N_3544,In_112,In_274);
and U3545 (N_3545,In_939,In_544);
xnor U3546 (N_3546,In_563,In_556);
or U3547 (N_3547,In_689,In_169);
or U3548 (N_3548,In_907,In_961);
and U3549 (N_3549,In_305,In_214);
xor U3550 (N_3550,In_643,In_55);
nor U3551 (N_3551,In_990,In_15);
or U3552 (N_3552,In_167,In_87);
nand U3553 (N_3553,In_59,In_348);
or U3554 (N_3554,In_314,In_860);
and U3555 (N_3555,In_813,In_588);
or U3556 (N_3556,In_732,In_819);
nand U3557 (N_3557,In_755,In_820);
or U3558 (N_3558,In_999,In_613);
and U3559 (N_3559,In_470,In_504);
or U3560 (N_3560,In_251,In_558);
nor U3561 (N_3561,In_610,In_997);
and U3562 (N_3562,In_301,In_524);
nor U3563 (N_3563,In_818,In_46);
and U3564 (N_3564,In_914,In_296);
nor U3565 (N_3565,In_546,In_942);
nor U3566 (N_3566,In_648,In_315);
nand U3567 (N_3567,In_315,In_886);
nor U3568 (N_3568,In_560,In_203);
and U3569 (N_3569,In_790,In_732);
nand U3570 (N_3570,In_134,In_673);
or U3571 (N_3571,In_276,In_558);
or U3572 (N_3572,In_806,In_759);
and U3573 (N_3573,In_755,In_325);
or U3574 (N_3574,In_366,In_356);
or U3575 (N_3575,In_5,In_504);
and U3576 (N_3576,In_343,In_99);
nor U3577 (N_3577,In_370,In_451);
and U3578 (N_3578,In_89,In_85);
or U3579 (N_3579,In_86,In_780);
nor U3580 (N_3580,In_591,In_557);
and U3581 (N_3581,In_791,In_555);
and U3582 (N_3582,In_307,In_302);
and U3583 (N_3583,In_151,In_978);
xor U3584 (N_3584,In_66,In_255);
nor U3585 (N_3585,In_572,In_395);
nand U3586 (N_3586,In_897,In_666);
nor U3587 (N_3587,In_871,In_591);
nand U3588 (N_3588,In_906,In_59);
nand U3589 (N_3589,In_793,In_575);
nor U3590 (N_3590,In_246,In_79);
or U3591 (N_3591,In_176,In_142);
xor U3592 (N_3592,In_93,In_756);
nand U3593 (N_3593,In_666,In_636);
nor U3594 (N_3594,In_603,In_876);
nand U3595 (N_3595,In_650,In_741);
nor U3596 (N_3596,In_113,In_316);
nor U3597 (N_3597,In_69,In_231);
or U3598 (N_3598,In_266,In_361);
or U3599 (N_3599,In_737,In_35);
and U3600 (N_3600,In_492,In_871);
xnor U3601 (N_3601,In_391,In_845);
xor U3602 (N_3602,In_925,In_603);
xnor U3603 (N_3603,In_782,In_835);
and U3604 (N_3604,In_285,In_57);
or U3605 (N_3605,In_623,In_249);
xnor U3606 (N_3606,In_865,In_264);
xnor U3607 (N_3607,In_689,In_933);
nor U3608 (N_3608,In_558,In_997);
nand U3609 (N_3609,In_367,In_171);
and U3610 (N_3610,In_251,In_123);
nand U3611 (N_3611,In_787,In_189);
xnor U3612 (N_3612,In_754,In_659);
and U3613 (N_3613,In_461,In_241);
nor U3614 (N_3614,In_615,In_657);
or U3615 (N_3615,In_800,In_394);
and U3616 (N_3616,In_406,In_911);
or U3617 (N_3617,In_145,In_687);
nor U3618 (N_3618,In_774,In_767);
xor U3619 (N_3619,In_565,In_294);
or U3620 (N_3620,In_356,In_411);
nand U3621 (N_3621,In_508,In_763);
nand U3622 (N_3622,In_882,In_985);
or U3623 (N_3623,In_899,In_599);
nand U3624 (N_3624,In_770,In_645);
nand U3625 (N_3625,In_131,In_261);
or U3626 (N_3626,In_412,In_597);
xor U3627 (N_3627,In_334,In_854);
and U3628 (N_3628,In_970,In_520);
or U3629 (N_3629,In_798,In_767);
or U3630 (N_3630,In_404,In_4);
nor U3631 (N_3631,In_30,In_635);
and U3632 (N_3632,In_829,In_807);
nor U3633 (N_3633,In_431,In_52);
and U3634 (N_3634,In_129,In_553);
nand U3635 (N_3635,In_451,In_968);
nor U3636 (N_3636,In_241,In_796);
nor U3637 (N_3637,In_346,In_118);
and U3638 (N_3638,In_380,In_934);
and U3639 (N_3639,In_357,In_342);
and U3640 (N_3640,In_814,In_798);
or U3641 (N_3641,In_213,In_769);
nand U3642 (N_3642,In_121,In_285);
nor U3643 (N_3643,In_842,In_367);
xor U3644 (N_3644,In_837,In_217);
and U3645 (N_3645,In_838,In_845);
or U3646 (N_3646,In_592,In_363);
or U3647 (N_3647,In_757,In_376);
and U3648 (N_3648,In_328,In_488);
or U3649 (N_3649,In_266,In_474);
xnor U3650 (N_3650,In_264,In_4);
xnor U3651 (N_3651,In_729,In_800);
or U3652 (N_3652,In_626,In_304);
and U3653 (N_3653,In_600,In_371);
xor U3654 (N_3654,In_996,In_22);
and U3655 (N_3655,In_802,In_691);
nand U3656 (N_3656,In_252,In_393);
nand U3657 (N_3657,In_931,In_938);
and U3658 (N_3658,In_158,In_19);
nor U3659 (N_3659,In_440,In_461);
nor U3660 (N_3660,In_148,In_379);
nand U3661 (N_3661,In_348,In_40);
and U3662 (N_3662,In_181,In_179);
nor U3663 (N_3663,In_338,In_311);
nand U3664 (N_3664,In_888,In_347);
and U3665 (N_3665,In_306,In_338);
nand U3666 (N_3666,In_120,In_705);
xor U3667 (N_3667,In_776,In_467);
xnor U3668 (N_3668,In_75,In_866);
xnor U3669 (N_3669,In_788,In_805);
xnor U3670 (N_3670,In_428,In_87);
xor U3671 (N_3671,In_679,In_495);
xor U3672 (N_3672,In_603,In_567);
xnor U3673 (N_3673,In_789,In_379);
nand U3674 (N_3674,In_731,In_809);
xor U3675 (N_3675,In_430,In_387);
nand U3676 (N_3676,In_668,In_870);
nor U3677 (N_3677,In_981,In_531);
or U3678 (N_3678,In_872,In_189);
or U3679 (N_3679,In_374,In_181);
and U3680 (N_3680,In_982,In_606);
or U3681 (N_3681,In_730,In_991);
nor U3682 (N_3682,In_379,In_483);
nand U3683 (N_3683,In_501,In_616);
nor U3684 (N_3684,In_114,In_462);
or U3685 (N_3685,In_46,In_807);
and U3686 (N_3686,In_203,In_490);
nor U3687 (N_3687,In_808,In_969);
nor U3688 (N_3688,In_941,In_352);
nand U3689 (N_3689,In_869,In_32);
or U3690 (N_3690,In_682,In_622);
xor U3691 (N_3691,In_21,In_413);
and U3692 (N_3692,In_125,In_406);
or U3693 (N_3693,In_709,In_172);
nand U3694 (N_3694,In_122,In_977);
nand U3695 (N_3695,In_590,In_326);
nand U3696 (N_3696,In_407,In_629);
and U3697 (N_3697,In_927,In_92);
nor U3698 (N_3698,In_68,In_899);
or U3699 (N_3699,In_187,In_597);
nand U3700 (N_3700,In_320,In_274);
nor U3701 (N_3701,In_259,In_978);
and U3702 (N_3702,In_994,In_88);
nand U3703 (N_3703,In_409,In_934);
nand U3704 (N_3704,In_468,In_260);
or U3705 (N_3705,In_794,In_212);
and U3706 (N_3706,In_774,In_201);
or U3707 (N_3707,In_496,In_277);
xor U3708 (N_3708,In_327,In_665);
xnor U3709 (N_3709,In_801,In_496);
nand U3710 (N_3710,In_651,In_682);
and U3711 (N_3711,In_778,In_386);
and U3712 (N_3712,In_596,In_315);
nand U3713 (N_3713,In_326,In_400);
or U3714 (N_3714,In_510,In_788);
xnor U3715 (N_3715,In_744,In_449);
or U3716 (N_3716,In_811,In_574);
nand U3717 (N_3717,In_515,In_13);
xnor U3718 (N_3718,In_948,In_633);
nand U3719 (N_3719,In_150,In_172);
xnor U3720 (N_3720,In_859,In_656);
or U3721 (N_3721,In_158,In_380);
and U3722 (N_3722,In_867,In_191);
or U3723 (N_3723,In_575,In_847);
nand U3724 (N_3724,In_921,In_660);
nor U3725 (N_3725,In_917,In_760);
xor U3726 (N_3726,In_223,In_198);
or U3727 (N_3727,In_179,In_396);
and U3728 (N_3728,In_54,In_699);
and U3729 (N_3729,In_111,In_257);
nand U3730 (N_3730,In_57,In_257);
and U3731 (N_3731,In_556,In_252);
nor U3732 (N_3732,In_200,In_315);
nand U3733 (N_3733,In_602,In_183);
nor U3734 (N_3734,In_327,In_0);
xnor U3735 (N_3735,In_866,In_400);
nand U3736 (N_3736,In_958,In_983);
and U3737 (N_3737,In_301,In_669);
nand U3738 (N_3738,In_880,In_473);
nand U3739 (N_3739,In_282,In_828);
xnor U3740 (N_3740,In_63,In_898);
or U3741 (N_3741,In_727,In_757);
or U3742 (N_3742,In_768,In_181);
and U3743 (N_3743,In_414,In_937);
nand U3744 (N_3744,In_731,In_60);
nor U3745 (N_3745,In_782,In_359);
nor U3746 (N_3746,In_665,In_407);
and U3747 (N_3747,In_926,In_94);
and U3748 (N_3748,In_44,In_301);
or U3749 (N_3749,In_369,In_802);
and U3750 (N_3750,In_870,In_288);
xor U3751 (N_3751,In_14,In_842);
and U3752 (N_3752,In_56,In_832);
nor U3753 (N_3753,In_879,In_380);
or U3754 (N_3754,In_784,In_139);
or U3755 (N_3755,In_341,In_566);
and U3756 (N_3756,In_601,In_613);
or U3757 (N_3757,In_552,In_932);
xor U3758 (N_3758,In_893,In_25);
xor U3759 (N_3759,In_294,In_211);
nand U3760 (N_3760,In_141,In_846);
nand U3761 (N_3761,In_482,In_993);
nor U3762 (N_3762,In_51,In_61);
nand U3763 (N_3763,In_817,In_799);
nor U3764 (N_3764,In_29,In_40);
nor U3765 (N_3765,In_691,In_911);
nand U3766 (N_3766,In_168,In_209);
and U3767 (N_3767,In_4,In_119);
or U3768 (N_3768,In_316,In_495);
nand U3769 (N_3769,In_515,In_343);
xnor U3770 (N_3770,In_596,In_556);
xor U3771 (N_3771,In_759,In_176);
or U3772 (N_3772,In_147,In_559);
xor U3773 (N_3773,In_646,In_171);
or U3774 (N_3774,In_377,In_307);
or U3775 (N_3775,In_515,In_143);
and U3776 (N_3776,In_901,In_872);
nor U3777 (N_3777,In_753,In_299);
or U3778 (N_3778,In_26,In_275);
or U3779 (N_3779,In_166,In_900);
nand U3780 (N_3780,In_577,In_771);
and U3781 (N_3781,In_245,In_68);
and U3782 (N_3782,In_881,In_594);
or U3783 (N_3783,In_394,In_677);
nand U3784 (N_3784,In_522,In_508);
and U3785 (N_3785,In_146,In_22);
nand U3786 (N_3786,In_781,In_280);
or U3787 (N_3787,In_487,In_853);
nor U3788 (N_3788,In_524,In_259);
or U3789 (N_3789,In_741,In_940);
nor U3790 (N_3790,In_952,In_711);
nand U3791 (N_3791,In_700,In_346);
or U3792 (N_3792,In_21,In_271);
xor U3793 (N_3793,In_570,In_904);
or U3794 (N_3794,In_443,In_262);
nand U3795 (N_3795,In_941,In_308);
and U3796 (N_3796,In_399,In_724);
or U3797 (N_3797,In_183,In_811);
nand U3798 (N_3798,In_177,In_244);
and U3799 (N_3799,In_156,In_729);
and U3800 (N_3800,In_614,In_693);
nor U3801 (N_3801,In_645,In_721);
nand U3802 (N_3802,In_265,In_305);
nor U3803 (N_3803,In_314,In_330);
nor U3804 (N_3804,In_514,In_893);
nand U3805 (N_3805,In_474,In_962);
or U3806 (N_3806,In_4,In_191);
nor U3807 (N_3807,In_863,In_42);
or U3808 (N_3808,In_203,In_976);
or U3809 (N_3809,In_713,In_317);
or U3810 (N_3810,In_221,In_947);
and U3811 (N_3811,In_880,In_238);
or U3812 (N_3812,In_122,In_295);
nand U3813 (N_3813,In_178,In_224);
xor U3814 (N_3814,In_172,In_749);
nor U3815 (N_3815,In_408,In_691);
nor U3816 (N_3816,In_825,In_11);
xor U3817 (N_3817,In_120,In_243);
nand U3818 (N_3818,In_516,In_51);
and U3819 (N_3819,In_446,In_238);
and U3820 (N_3820,In_472,In_490);
and U3821 (N_3821,In_617,In_388);
nand U3822 (N_3822,In_366,In_768);
nand U3823 (N_3823,In_429,In_585);
and U3824 (N_3824,In_422,In_870);
or U3825 (N_3825,In_432,In_943);
or U3826 (N_3826,In_665,In_251);
xor U3827 (N_3827,In_48,In_178);
xnor U3828 (N_3828,In_386,In_882);
xnor U3829 (N_3829,In_122,In_333);
xnor U3830 (N_3830,In_121,In_146);
and U3831 (N_3831,In_921,In_78);
and U3832 (N_3832,In_918,In_911);
xnor U3833 (N_3833,In_443,In_744);
or U3834 (N_3834,In_575,In_739);
or U3835 (N_3835,In_669,In_595);
xnor U3836 (N_3836,In_453,In_150);
nand U3837 (N_3837,In_882,In_446);
nand U3838 (N_3838,In_369,In_274);
xor U3839 (N_3839,In_982,In_198);
nor U3840 (N_3840,In_181,In_947);
nand U3841 (N_3841,In_436,In_258);
xor U3842 (N_3842,In_536,In_502);
xor U3843 (N_3843,In_136,In_845);
or U3844 (N_3844,In_93,In_278);
and U3845 (N_3845,In_401,In_275);
xnor U3846 (N_3846,In_42,In_578);
and U3847 (N_3847,In_538,In_943);
nor U3848 (N_3848,In_439,In_86);
nand U3849 (N_3849,In_764,In_377);
nand U3850 (N_3850,In_9,In_677);
nor U3851 (N_3851,In_326,In_423);
or U3852 (N_3852,In_941,In_133);
xnor U3853 (N_3853,In_981,In_698);
nor U3854 (N_3854,In_667,In_574);
and U3855 (N_3855,In_902,In_622);
and U3856 (N_3856,In_55,In_479);
and U3857 (N_3857,In_622,In_767);
nand U3858 (N_3858,In_574,In_317);
and U3859 (N_3859,In_549,In_869);
nor U3860 (N_3860,In_498,In_635);
or U3861 (N_3861,In_757,In_665);
nor U3862 (N_3862,In_312,In_564);
nor U3863 (N_3863,In_896,In_519);
and U3864 (N_3864,In_499,In_926);
or U3865 (N_3865,In_159,In_227);
xor U3866 (N_3866,In_553,In_755);
or U3867 (N_3867,In_781,In_782);
nand U3868 (N_3868,In_788,In_438);
and U3869 (N_3869,In_322,In_369);
or U3870 (N_3870,In_793,In_376);
and U3871 (N_3871,In_154,In_950);
and U3872 (N_3872,In_463,In_653);
nor U3873 (N_3873,In_4,In_999);
nand U3874 (N_3874,In_687,In_268);
xor U3875 (N_3875,In_918,In_184);
and U3876 (N_3876,In_64,In_464);
xor U3877 (N_3877,In_480,In_351);
and U3878 (N_3878,In_212,In_710);
nor U3879 (N_3879,In_683,In_460);
nand U3880 (N_3880,In_207,In_38);
or U3881 (N_3881,In_130,In_970);
nand U3882 (N_3882,In_410,In_618);
or U3883 (N_3883,In_276,In_357);
or U3884 (N_3884,In_960,In_745);
and U3885 (N_3885,In_373,In_509);
xor U3886 (N_3886,In_847,In_114);
or U3887 (N_3887,In_489,In_327);
nor U3888 (N_3888,In_954,In_461);
and U3889 (N_3889,In_549,In_625);
xor U3890 (N_3890,In_457,In_914);
or U3891 (N_3891,In_364,In_503);
nor U3892 (N_3892,In_14,In_683);
nor U3893 (N_3893,In_807,In_102);
nand U3894 (N_3894,In_63,In_551);
xor U3895 (N_3895,In_581,In_974);
nor U3896 (N_3896,In_414,In_938);
or U3897 (N_3897,In_768,In_554);
nand U3898 (N_3898,In_989,In_337);
and U3899 (N_3899,In_553,In_867);
nand U3900 (N_3900,In_400,In_622);
nor U3901 (N_3901,In_566,In_674);
or U3902 (N_3902,In_150,In_477);
or U3903 (N_3903,In_520,In_781);
and U3904 (N_3904,In_313,In_182);
xor U3905 (N_3905,In_417,In_791);
nor U3906 (N_3906,In_751,In_378);
xnor U3907 (N_3907,In_353,In_310);
xnor U3908 (N_3908,In_386,In_396);
or U3909 (N_3909,In_657,In_567);
nor U3910 (N_3910,In_193,In_91);
or U3911 (N_3911,In_442,In_56);
or U3912 (N_3912,In_630,In_16);
nand U3913 (N_3913,In_557,In_56);
nor U3914 (N_3914,In_819,In_98);
nand U3915 (N_3915,In_337,In_937);
nor U3916 (N_3916,In_650,In_744);
nand U3917 (N_3917,In_521,In_655);
nand U3918 (N_3918,In_952,In_469);
xnor U3919 (N_3919,In_840,In_545);
nand U3920 (N_3920,In_81,In_983);
xor U3921 (N_3921,In_449,In_319);
nand U3922 (N_3922,In_887,In_674);
nand U3923 (N_3923,In_482,In_713);
or U3924 (N_3924,In_739,In_918);
and U3925 (N_3925,In_764,In_498);
nand U3926 (N_3926,In_350,In_702);
nand U3927 (N_3927,In_503,In_273);
xnor U3928 (N_3928,In_64,In_905);
nand U3929 (N_3929,In_799,In_681);
nand U3930 (N_3930,In_425,In_797);
nor U3931 (N_3931,In_953,In_433);
and U3932 (N_3932,In_311,In_613);
and U3933 (N_3933,In_521,In_215);
xnor U3934 (N_3934,In_112,In_101);
nor U3935 (N_3935,In_753,In_332);
and U3936 (N_3936,In_853,In_72);
nor U3937 (N_3937,In_111,In_900);
nor U3938 (N_3938,In_677,In_304);
nor U3939 (N_3939,In_399,In_809);
or U3940 (N_3940,In_901,In_60);
nor U3941 (N_3941,In_853,In_437);
or U3942 (N_3942,In_997,In_371);
and U3943 (N_3943,In_574,In_304);
and U3944 (N_3944,In_933,In_471);
xor U3945 (N_3945,In_219,In_920);
nor U3946 (N_3946,In_8,In_834);
or U3947 (N_3947,In_193,In_69);
nand U3948 (N_3948,In_826,In_194);
nor U3949 (N_3949,In_511,In_84);
nand U3950 (N_3950,In_625,In_880);
or U3951 (N_3951,In_57,In_591);
xor U3952 (N_3952,In_401,In_878);
and U3953 (N_3953,In_533,In_517);
xor U3954 (N_3954,In_128,In_450);
nand U3955 (N_3955,In_526,In_785);
nand U3956 (N_3956,In_578,In_186);
xnor U3957 (N_3957,In_920,In_517);
xor U3958 (N_3958,In_530,In_238);
nand U3959 (N_3959,In_929,In_555);
nor U3960 (N_3960,In_885,In_198);
xnor U3961 (N_3961,In_134,In_383);
and U3962 (N_3962,In_66,In_382);
or U3963 (N_3963,In_325,In_126);
nand U3964 (N_3964,In_407,In_199);
xnor U3965 (N_3965,In_95,In_768);
xor U3966 (N_3966,In_908,In_13);
or U3967 (N_3967,In_466,In_785);
xor U3968 (N_3968,In_396,In_588);
and U3969 (N_3969,In_630,In_164);
nor U3970 (N_3970,In_722,In_276);
or U3971 (N_3971,In_966,In_145);
nor U3972 (N_3972,In_555,In_42);
and U3973 (N_3973,In_381,In_240);
xnor U3974 (N_3974,In_497,In_882);
nand U3975 (N_3975,In_352,In_627);
and U3976 (N_3976,In_682,In_116);
and U3977 (N_3977,In_701,In_19);
nor U3978 (N_3978,In_685,In_315);
nor U3979 (N_3979,In_859,In_89);
nand U3980 (N_3980,In_243,In_719);
and U3981 (N_3981,In_891,In_916);
nand U3982 (N_3982,In_483,In_167);
and U3983 (N_3983,In_280,In_475);
nand U3984 (N_3984,In_167,In_554);
nand U3985 (N_3985,In_486,In_509);
nor U3986 (N_3986,In_272,In_13);
nand U3987 (N_3987,In_363,In_580);
nor U3988 (N_3988,In_123,In_803);
xor U3989 (N_3989,In_657,In_241);
nor U3990 (N_3990,In_321,In_559);
and U3991 (N_3991,In_497,In_481);
nor U3992 (N_3992,In_261,In_433);
and U3993 (N_3993,In_993,In_377);
or U3994 (N_3994,In_457,In_79);
or U3995 (N_3995,In_842,In_668);
nor U3996 (N_3996,In_976,In_118);
and U3997 (N_3997,In_642,In_646);
or U3998 (N_3998,In_451,In_221);
xor U3999 (N_3999,In_385,In_86);
and U4000 (N_4000,In_434,In_747);
or U4001 (N_4001,In_531,In_608);
and U4002 (N_4002,In_914,In_977);
or U4003 (N_4003,In_288,In_996);
nor U4004 (N_4004,In_956,In_578);
nand U4005 (N_4005,In_275,In_908);
xnor U4006 (N_4006,In_4,In_663);
nand U4007 (N_4007,In_599,In_6);
and U4008 (N_4008,In_677,In_395);
nand U4009 (N_4009,In_55,In_490);
or U4010 (N_4010,In_721,In_693);
nand U4011 (N_4011,In_273,In_119);
and U4012 (N_4012,In_464,In_732);
nor U4013 (N_4013,In_378,In_675);
and U4014 (N_4014,In_911,In_306);
and U4015 (N_4015,In_49,In_470);
or U4016 (N_4016,In_446,In_579);
and U4017 (N_4017,In_8,In_84);
nand U4018 (N_4018,In_802,In_552);
nor U4019 (N_4019,In_596,In_472);
xnor U4020 (N_4020,In_21,In_971);
and U4021 (N_4021,In_88,In_344);
nand U4022 (N_4022,In_612,In_995);
xnor U4023 (N_4023,In_931,In_776);
or U4024 (N_4024,In_141,In_930);
or U4025 (N_4025,In_696,In_913);
xnor U4026 (N_4026,In_797,In_871);
xor U4027 (N_4027,In_162,In_100);
nor U4028 (N_4028,In_344,In_392);
and U4029 (N_4029,In_949,In_739);
nand U4030 (N_4030,In_432,In_385);
xnor U4031 (N_4031,In_558,In_418);
or U4032 (N_4032,In_255,In_30);
xor U4033 (N_4033,In_511,In_938);
or U4034 (N_4034,In_966,In_527);
xnor U4035 (N_4035,In_948,In_978);
nor U4036 (N_4036,In_536,In_54);
and U4037 (N_4037,In_882,In_372);
or U4038 (N_4038,In_270,In_378);
or U4039 (N_4039,In_276,In_730);
or U4040 (N_4040,In_306,In_330);
nor U4041 (N_4041,In_821,In_578);
or U4042 (N_4042,In_178,In_209);
or U4043 (N_4043,In_947,In_239);
nor U4044 (N_4044,In_604,In_533);
nor U4045 (N_4045,In_937,In_510);
and U4046 (N_4046,In_635,In_713);
nor U4047 (N_4047,In_113,In_493);
nor U4048 (N_4048,In_285,In_501);
and U4049 (N_4049,In_410,In_178);
xor U4050 (N_4050,In_198,In_486);
or U4051 (N_4051,In_625,In_157);
and U4052 (N_4052,In_972,In_452);
and U4053 (N_4053,In_994,In_10);
nor U4054 (N_4054,In_539,In_918);
nand U4055 (N_4055,In_605,In_551);
and U4056 (N_4056,In_538,In_787);
nand U4057 (N_4057,In_35,In_312);
xnor U4058 (N_4058,In_206,In_687);
xnor U4059 (N_4059,In_697,In_435);
and U4060 (N_4060,In_172,In_180);
nand U4061 (N_4061,In_496,In_334);
or U4062 (N_4062,In_572,In_378);
or U4063 (N_4063,In_622,In_890);
and U4064 (N_4064,In_385,In_161);
or U4065 (N_4065,In_932,In_858);
and U4066 (N_4066,In_800,In_360);
nand U4067 (N_4067,In_779,In_541);
nor U4068 (N_4068,In_580,In_913);
xnor U4069 (N_4069,In_588,In_721);
nand U4070 (N_4070,In_918,In_257);
nor U4071 (N_4071,In_324,In_874);
xor U4072 (N_4072,In_128,In_660);
nand U4073 (N_4073,In_995,In_497);
or U4074 (N_4074,In_167,In_916);
xnor U4075 (N_4075,In_918,In_105);
or U4076 (N_4076,In_570,In_789);
and U4077 (N_4077,In_185,In_104);
or U4078 (N_4078,In_613,In_990);
nor U4079 (N_4079,In_53,In_156);
xor U4080 (N_4080,In_975,In_517);
xnor U4081 (N_4081,In_696,In_942);
nor U4082 (N_4082,In_931,In_179);
nor U4083 (N_4083,In_911,In_153);
and U4084 (N_4084,In_265,In_78);
nand U4085 (N_4085,In_995,In_255);
nor U4086 (N_4086,In_316,In_463);
nor U4087 (N_4087,In_183,In_643);
xnor U4088 (N_4088,In_103,In_579);
nand U4089 (N_4089,In_23,In_870);
or U4090 (N_4090,In_860,In_527);
xor U4091 (N_4091,In_992,In_79);
or U4092 (N_4092,In_168,In_912);
nor U4093 (N_4093,In_396,In_275);
xnor U4094 (N_4094,In_240,In_452);
nor U4095 (N_4095,In_203,In_698);
xnor U4096 (N_4096,In_103,In_422);
and U4097 (N_4097,In_939,In_18);
or U4098 (N_4098,In_573,In_13);
nor U4099 (N_4099,In_276,In_5);
and U4100 (N_4100,In_32,In_545);
xnor U4101 (N_4101,In_657,In_254);
or U4102 (N_4102,In_404,In_835);
and U4103 (N_4103,In_639,In_626);
xor U4104 (N_4104,In_134,In_853);
or U4105 (N_4105,In_806,In_237);
xor U4106 (N_4106,In_327,In_92);
and U4107 (N_4107,In_359,In_848);
nor U4108 (N_4108,In_820,In_433);
and U4109 (N_4109,In_124,In_615);
xor U4110 (N_4110,In_864,In_91);
or U4111 (N_4111,In_858,In_874);
nor U4112 (N_4112,In_338,In_604);
xor U4113 (N_4113,In_814,In_55);
and U4114 (N_4114,In_236,In_87);
xor U4115 (N_4115,In_348,In_521);
and U4116 (N_4116,In_841,In_624);
nand U4117 (N_4117,In_235,In_440);
and U4118 (N_4118,In_297,In_26);
nor U4119 (N_4119,In_858,In_584);
xor U4120 (N_4120,In_199,In_276);
xor U4121 (N_4121,In_329,In_898);
nand U4122 (N_4122,In_104,In_915);
and U4123 (N_4123,In_554,In_106);
xnor U4124 (N_4124,In_207,In_43);
or U4125 (N_4125,In_119,In_55);
and U4126 (N_4126,In_905,In_337);
nor U4127 (N_4127,In_201,In_272);
xor U4128 (N_4128,In_826,In_587);
nor U4129 (N_4129,In_194,In_714);
or U4130 (N_4130,In_989,In_55);
nor U4131 (N_4131,In_885,In_866);
nor U4132 (N_4132,In_507,In_593);
nand U4133 (N_4133,In_362,In_806);
nor U4134 (N_4134,In_294,In_576);
nand U4135 (N_4135,In_684,In_153);
and U4136 (N_4136,In_902,In_537);
and U4137 (N_4137,In_198,In_300);
and U4138 (N_4138,In_827,In_711);
or U4139 (N_4139,In_584,In_30);
nand U4140 (N_4140,In_781,In_43);
and U4141 (N_4141,In_905,In_195);
or U4142 (N_4142,In_614,In_935);
and U4143 (N_4143,In_350,In_754);
and U4144 (N_4144,In_632,In_26);
xnor U4145 (N_4145,In_550,In_759);
and U4146 (N_4146,In_887,In_467);
and U4147 (N_4147,In_336,In_29);
xor U4148 (N_4148,In_930,In_658);
and U4149 (N_4149,In_148,In_37);
nand U4150 (N_4150,In_183,In_530);
xnor U4151 (N_4151,In_441,In_811);
or U4152 (N_4152,In_119,In_555);
xor U4153 (N_4153,In_313,In_321);
or U4154 (N_4154,In_61,In_823);
nand U4155 (N_4155,In_884,In_413);
or U4156 (N_4156,In_196,In_215);
and U4157 (N_4157,In_588,In_214);
nor U4158 (N_4158,In_433,In_316);
or U4159 (N_4159,In_181,In_410);
nand U4160 (N_4160,In_822,In_234);
and U4161 (N_4161,In_52,In_62);
nand U4162 (N_4162,In_227,In_747);
or U4163 (N_4163,In_96,In_874);
or U4164 (N_4164,In_693,In_477);
nand U4165 (N_4165,In_97,In_824);
xor U4166 (N_4166,In_59,In_36);
nand U4167 (N_4167,In_436,In_455);
xor U4168 (N_4168,In_123,In_846);
xnor U4169 (N_4169,In_614,In_983);
xor U4170 (N_4170,In_395,In_869);
nand U4171 (N_4171,In_353,In_731);
nor U4172 (N_4172,In_950,In_526);
or U4173 (N_4173,In_328,In_415);
or U4174 (N_4174,In_467,In_343);
or U4175 (N_4175,In_359,In_517);
nand U4176 (N_4176,In_698,In_773);
xor U4177 (N_4177,In_265,In_909);
nand U4178 (N_4178,In_122,In_507);
nand U4179 (N_4179,In_807,In_212);
xor U4180 (N_4180,In_353,In_683);
xor U4181 (N_4181,In_312,In_826);
xnor U4182 (N_4182,In_889,In_199);
nor U4183 (N_4183,In_810,In_706);
and U4184 (N_4184,In_455,In_527);
xor U4185 (N_4185,In_214,In_46);
or U4186 (N_4186,In_295,In_928);
nor U4187 (N_4187,In_859,In_866);
or U4188 (N_4188,In_381,In_483);
and U4189 (N_4189,In_946,In_81);
nand U4190 (N_4190,In_728,In_659);
nor U4191 (N_4191,In_67,In_771);
nand U4192 (N_4192,In_345,In_133);
xor U4193 (N_4193,In_490,In_252);
xor U4194 (N_4194,In_389,In_19);
or U4195 (N_4195,In_27,In_774);
xnor U4196 (N_4196,In_399,In_668);
xnor U4197 (N_4197,In_365,In_629);
xor U4198 (N_4198,In_823,In_488);
nand U4199 (N_4199,In_457,In_182);
nor U4200 (N_4200,In_15,In_570);
and U4201 (N_4201,In_188,In_301);
xor U4202 (N_4202,In_129,In_616);
nand U4203 (N_4203,In_586,In_282);
nand U4204 (N_4204,In_176,In_795);
nand U4205 (N_4205,In_771,In_256);
nor U4206 (N_4206,In_301,In_194);
or U4207 (N_4207,In_129,In_896);
or U4208 (N_4208,In_320,In_185);
xor U4209 (N_4209,In_749,In_729);
nor U4210 (N_4210,In_683,In_892);
and U4211 (N_4211,In_697,In_34);
xor U4212 (N_4212,In_490,In_823);
nand U4213 (N_4213,In_560,In_844);
xor U4214 (N_4214,In_462,In_420);
or U4215 (N_4215,In_596,In_355);
xor U4216 (N_4216,In_332,In_353);
xor U4217 (N_4217,In_57,In_981);
or U4218 (N_4218,In_138,In_30);
xor U4219 (N_4219,In_474,In_605);
nand U4220 (N_4220,In_330,In_528);
nor U4221 (N_4221,In_510,In_252);
nand U4222 (N_4222,In_818,In_27);
nand U4223 (N_4223,In_343,In_21);
xnor U4224 (N_4224,In_883,In_291);
or U4225 (N_4225,In_18,In_500);
and U4226 (N_4226,In_352,In_556);
and U4227 (N_4227,In_28,In_642);
and U4228 (N_4228,In_237,In_378);
or U4229 (N_4229,In_681,In_516);
or U4230 (N_4230,In_738,In_401);
or U4231 (N_4231,In_667,In_770);
or U4232 (N_4232,In_289,In_445);
nor U4233 (N_4233,In_599,In_77);
nor U4234 (N_4234,In_593,In_644);
and U4235 (N_4235,In_132,In_698);
xor U4236 (N_4236,In_87,In_410);
nor U4237 (N_4237,In_512,In_797);
and U4238 (N_4238,In_243,In_639);
or U4239 (N_4239,In_109,In_937);
xnor U4240 (N_4240,In_27,In_880);
or U4241 (N_4241,In_475,In_105);
nor U4242 (N_4242,In_109,In_236);
nand U4243 (N_4243,In_455,In_397);
and U4244 (N_4244,In_287,In_804);
nand U4245 (N_4245,In_247,In_419);
nand U4246 (N_4246,In_130,In_414);
or U4247 (N_4247,In_266,In_113);
nor U4248 (N_4248,In_446,In_732);
nor U4249 (N_4249,In_114,In_973);
and U4250 (N_4250,In_233,In_744);
xnor U4251 (N_4251,In_379,In_346);
xor U4252 (N_4252,In_227,In_262);
nand U4253 (N_4253,In_79,In_175);
nand U4254 (N_4254,In_906,In_189);
and U4255 (N_4255,In_235,In_91);
nand U4256 (N_4256,In_334,In_137);
nand U4257 (N_4257,In_335,In_161);
xor U4258 (N_4258,In_901,In_966);
or U4259 (N_4259,In_507,In_802);
or U4260 (N_4260,In_635,In_993);
nor U4261 (N_4261,In_460,In_932);
nand U4262 (N_4262,In_195,In_799);
nand U4263 (N_4263,In_593,In_903);
xor U4264 (N_4264,In_728,In_72);
or U4265 (N_4265,In_930,In_728);
and U4266 (N_4266,In_878,In_97);
and U4267 (N_4267,In_104,In_357);
nand U4268 (N_4268,In_5,In_838);
and U4269 (N_4269,In_686,In_206);
or U4270 (N_4270,In_29,In_277);
nand U4271 (N_4271,In_98,In_692);
nand U4272 (N_4272,In_534,In_581);
nor U4273 (N_4273,In_494,In_788);
xor U4274 (N_4274,In_495,In_810);
xnor U4275 (N_4275,In_849,In_141);
xnor U4276 (N_4276,In_689,In_416);
nand U4277 (N_4277,In_672,In_578);
nand U4278 (N_4278,In_682,In_301);
nand U4279 (N_4279,In_324,In_679);
nor U4280 (N_4280,In_588,In_862);
xnor U4281 (N_4281,In_414,In_115);
nor U4282 (N_4282,In_315,In_355);
or U4283 (N_4283,In_207,In_130);
xor U4284 (N_4284,In_486,In_106);
nor U4285 (N_4285,In_885,In_841);
nand U4286 (N_4286,In_121,In_65);
or U4287 (N_4287,In_726,In_493);
nand U4288 (N_4288,In_265,In_181);
nor U4289 (N_4289,In_966,In_59);
and U4290 (N_4290,In_923,In_251);
nor U4291 (N_4291,In_224,In_158);
xnor U4292 (N_4292,In_251,In_934);
or U4293 (N_4293,In_801,In_201);
nor U4294 (N_4294,In_146,In_130);
nand U4295 (N_4295,In_737,In_947);
or U4296 (N_4296,In_311,In_371);
and U4297 (N_4297,In_718,In_692);
xnor U4298 (N_4298,In_208,In_274);
xnor U4299 (N_4299,In_438,In_903);
xnor U4300 (N_4300,In_181,In_282);
nor U4301 (N_4301,In_371,In_297);
and U4302 (N_4302,In_583,In_933);
nor U4303 (N_4303,In_919,In_542);
nor U4304 (N_4304,In_4,In_120);
and U4305 (N_4305,In_522,In_813);
nor U4306 (N_4306,In_936,In_468);
xnor U4307 (N_4307,In_207,In_905);
or U4308 (N_4308,In_995,In_950);
and U4309 (N_4309,In_506,In_620);
or U4310 (N_4310,In_107,In_208);
nand U4311 (N_4311,In_340,In_177);
xnor U4312 (N_4312,In_218,In_750);
xor U4313 (N_4313,In_878,In_933);
and U4314 (N_4314,In_988,In_710);
xnor U4315 (N_4315,In_742,In_389);
xnor U4316 (N_4316,In_429,In_145);
xor U4317 (N_4317,In_910,In_685);
and U4318 (N_4318,In_129,In_951);
xnor U4319 (N_4319,In_688,In_599);
and U4320 (N_4320,In_780,In_858);
xor U4321 (N_4321,In_618,In_420);
xnor U4322 (N_4322,In_14,In_522);
nand U4323 (N_4323,In_162,In_253);
xnor U4324 (N_4324,In_440,In_971);
nand U4325 (N_4325,In_287,In_656);
nand U4326 (N_4326,In_31,In_935);
nor U4327 (N_4327,In_831,In_9);
and U4328 (N_4328,In_321,In_259);
and U4329 (N_4329,In_960,In_640);
nor U4330 (N_4330,In_357,In_91);
xnor U4331 (N_4331,In_273,In_264);
nor U4332 (N_4332,In_537,In_545);
nand U4333 (N_4333,In_221,In_204);
or U4334 (N_4334,In_66,In_104);
and U4335 (N_4335,In_42,In_425);
nor U4336 (N_4336,In_919,In_546);
xor U4337 (N_4337,In_458,In_63);
xnor U4338 (N_4338,In_191,In_508);
or U4339 (N_4339,In_441,In_718);
nor U4340 (N_4340,In_541,In_758);
and U4341 (N_4341,In_4,In_414);
nor U4342 (N_4342,In_197,In_319);
and U4343 (N_4343,In_331,In_760);
or U4344 (N_4344,In_544,In_936);
xnor U4345 (N_4345,In_836,In_629);
xnor U4346 (N_4346,In_949,In_524);
and U4347 (N_4347,In_470,In_410);
or U4348 (N_4348,In_428,In_56);
xor U4349 (N_4349,In_497,In_306);
xnor U4350 (N_4350,In_306,In_991);
xor U4351 (N_4351,In_520,In_346);
or U4352 (N_4352,In_858,In_894);
and U4353 (N_4353,In_416,In_291);
and U4354 (N_4354,In_375,In_909);
nor U4355 (N_4355,In_144,In_440);
xnor U4356 (N_4356,In_465,In_846);
xor U4357 (N_4357,In_845,In_138);
and U4358 (N_4358,In_57,In_382);
xnor U4359 (N_4359,In_246,In_75);
and U4360 (N_4360,In_703,In_367);
or U4361 (N_4361,In_117,In_44);
nand U4362 (N_4362,In_868,In_835);
nor U4363 (N_4363,In_268,In_12);
or U4364 (N_4364,In_914,In_845);
nand U4365 (N_4365,In_564,In_348);
and U4366 (N_4366,In_540,In_386);
and U4367 (N_4367,In_433,In_677);
nor U4368 (N_4368,In_160,In_943);
or U4369 (N_4369,In_22,In_139);
or U4370 (N_4370,In_438,In_396);
xor U4371 (N_4371,In_892,In_170);
nor U4372 (N_4372,In_362,In_874);
xor U4373 (N_4373,In_31,In_41);
or U4374 (N_4374,In_689,In_355);
nor U4375 (N_4375,In_770,In_46);
nand U4376 (N_4376,In_427,In_989);
and U4377 (N_4377,In_947,In_228);
and U4378 (N_4378,In_722,In_473);
or U4379 (N_4379,In_780,In_646);
nand U4380 (N_4380,In_135,In_386);
nand U4381 (N_4381,In_531,In_784);
nor U4382 (N_4382,In_320,In_222);
xnor U4383 (N_4383,In_12,In_487);
or U4384 (N_4384,In_796,In_132);
or U4385 (N_4385,In_832,In_366);
nor U4386 (N_4386,In_229,In_531);
xnor U4387 (N_4387,In_667,In_897);
nand U4388 (N_4388,In_132,In_885);
nand U4389 (N_4389,In_102,In_700);
or U4390 (N_4390,In_585,In_589);
and U4391 (N_4391,In_98,In_160);
nor U4392 (N_4392,In_519,In_275);
xnor U4393 (N_4393,In_849,In_977);
xor U4394 (N_4394,In_864,In_480);
nand U4395 (N_4395,In_503,In_169);
or U4396 (N_4396,In_990,In_36);
or U4397 (N_4397,In_452,In_444);
or U4398 (N_4398,In_79,In_898);
or U4399 (N_4399,In_274,In_418);
nand U4400 (N_4400,In_27,In_407);
or U4401 (N_4401,In_995,In_226);
and U4402 (N_4402,In_32,In_13);
or U4403 (N_4403,In_750,In_905);
nand U4404 (N_4404,In_445,In_40);
nor U4405 (N_4405,In_722,In_534);
xor U4406 (N_4406,In_837,In_256);
and U4407 (N_4407,In_495,In_808);
and U4408 (N_4408,In_438,In_257);
or U4409 (N_4409,In_416,In_897);
or U4410 (N_4410,In_303,In_163);
nand U4411 (N_4411,In_479,In_531);
and U4412 (N_4412,In_909,In_922);
nor U4413 (N_4413,In_736,In_579);
nand U4414 (N_4414,In_580,In_610);
or U4415 (N_4415,In_46,In_461);
nor U4416 (N_4416,In_573,In_264);
nor U4417 (N_4417,In_430,In_823);
or U4418 (N_4418,In_376,In_538);
nand U4419 (N_4419,In_659,In_138);
nand U4420 (N_4420,In_161,In_814);
nand U4421 (N_4421,In_159,In_44);
nand U4422 (N_4422,In_340,In_584);
nor U4423 (N_4423,In_648,In_728);
nand U4424 (N_4424,In_402,In_193);
xnor U4425 (N_4425,In_893,In_951);
xnor U4426 (N_4426,In_831,In_803);
or U4427 (N_4427,In_869,In_587);
nor U4428 (N_4428,In_782,In_487);
and U4429 (N_4429,In_361,In_730);
xor U4430 (N_4430,In_152,In_571);
xor U4431 (N_4431,In_270,In_809);
nor U4432 (N_4432,In_899,In_521);
and U4433 (N_4433,In_775,In_547);
xor U4434 (N_4434,In_912,In_315);
xor U4435 (N_4435,In_140,In_376);
nor U4436 (N_4436,In_590,In_561);
or U4437 (N_4437,In_153,In_73);
and U4438 (N_4438,In_927,In_620);
xor U4439 (N_4439,In_494,In_208);
and U4440 (N_4440,In_809,In_779);
xnor U4441 (N_4441,In_438,In_828);
nand U4442 (N_4442,In_178,In_630);
and U4443 (N_4443,In_704,In_588);
nand U4444 (N_4444,In_268,In_97);
or U4445 (N_4445,In_295,In_17);
or U4446 (N_4446,In_572,In_939);
xnor U4447 (N_4447,In_342,In_609);
and U4448 (N_4448,In_402,In_544);
xor U4449 (N_4449,In_771,In_473);
and U4450 (N_4450,In_354,In_831);
or U4451 (N_4451,In_621,In_771);
or U4452 (N_4452,In_156,In_382);
and U4453 (N_4453,In_903,In_976);
or U4454 (N_4454,In_224,In_528);
nor U4455 (N_4455,In_956,In_635);
or U4456 (N_4456,In_792,In_653);
nor U4457 (N_4457,In_764,In_531);
nand U4458 (N_4458,In_548,In_39);
and U4459 (N_4459,In_413,In_578);
nor U4460 (N_4460,In_993,In_27);
xnor U4461 (N_4461,In_456,In_459);
nand U4462 (N_4462,In_97,In_560);
and U4463 (N_4463,In_65,In_551);
xor U4464 (N_4464,In_685,In_699);
nor U4465 (N_4465,In_559,In_671);
nor U4466 (N_4466,In_617,In_913);
xor U4467 (N_4467,In_947,In_602);
nand U4468 (N_4468,In_459,In_109);
xnor U4469 (N_4469,In_888,In_66);
and U4470 (N_4470,In_516,In_820);
xnor U4471 (N_4471,In_402,In_600);
nor U4472 (N_4472,In_59,In_234);
or U4473 (N_4473,In_529,In_537);
xnor U4474 (N_4474,In_525,In_505);
xnor U4475 (N_4475,In_515,In_95);
nand U4476 (N_4476,In_176,In_738);
xnor U4477 (N_4477,In_410,In_287);
nor U4478 (N_4478,In_619,In_567);
and U4479 (N_4479,In_516,In_965);
nand U4480 (N_4480,In_363,In_226);
or U4481 (N_4481,In_57,In_118);
and U4482 (N_4482,In_224,In_446);
nor U4483 (N_4483,In_320,In_515);
and U4484 (N_4484,In_72,In_547);
nor U4485 (N_4485,In_738,In_849);
and U4486 (N_4486,In_97,In_850);
nand U4487 (N_4487,In_571,In_704);
and U4488 (N_4488,In_897,In_735);
nor U4489 (N_4489,In_343,In_494);
nand U4490 (N_4490,In_781,In_0);
and U4491 (N_4491,In_829,In_659);
xor U4492 (N_4492,In_680,In_112);
nand U4493 (N_4493,In_796,In_496);
xor U4494 (N_4494,In_488,In_926);
or U4495 (N_4495,In_187,In_514);
xnor U4496 (N_4496,In_171,In_664);
xnor U4497 (N_4497,In_7,In_85);
nor U4498 (N_4498,In_443,In_358);
nor U4499 (N_4499,In_522,In_713);
nor U4500 (N_4500,In_749,In_760);
xnor U4501 (N_4501,In_659,In_189);
nor U4502 (N_4502,In_896,In_381);
or U4503 (N_4503,In_772,In_223);
and U4504 (N_4504,In_47,In_57);
and U4505 (N_4505,In_937,In_607);
xnor U4506 (N_4506,In_243,In_991);
or U4507 (N_4507,In_475,In_614);
xor U4508 (N_4508,In_691,In_99);
nand U4509 (N_4509,In_73,In_655);
and U4510 (N_4510,In_479,In_475);
nor U4511 (N_4511,In_572,In_111);
nor U4512 (N_4512,In_625,In_823);
and U4513 (N_4513,In_479,In_999);
xor U4514 (N_4514,In_148,In_211);
nor U4515 (N_4515,In_267,In_697);
and U4516 (N_4516,In_925,In_191);
and U4517 (N_4517,In_1,In_818);
or U4518 (N_4518,In_485,In_162);
nand U4519 (N_4519,In_499,In_30);
nor U4520 (N_4520,In_313,In_76);
nor U4521 (N_4521,In_480,In_483);
nor U4522 (N_4522,In_428,In_669);
nand U4523 (N_4523,In_245,In_834);
xor U4524 (N_4524,In_63,In_826);
nor U4525 (N_4525,In_103,In_368);
or U4526 (N_4526,In_790,In_504);
nand U4527 (N_4527,In_104,In_712);
xnor U4528 (N_4528,In_291,In_919);
nand U4529 (N_4529,In_279,In_313);
or U4530 (N_4530,In_377,In_927);
or U4531 (N_4531,In_730,In_715);
nor U4532 (N_4532,In_992,In_724);
xor U4533 (N_4533,In_255,In_440);
and U4534 (N_4534,In_915,In_433);
xnor U4535 (N_4535,In_537,In_895);
or U4536 (N_4536,In_195,In_217);
nor U4537 (N_4537,In_17,In_113);
or U4538 (N_4538,In_879,In_247);
xnor U4539 (N_4539,In_595,In_435);
and U4540 (N_4540,In_393,In_355);
nor U4541 (N_4541,In_585,In_493);
nor U4542 (N_4542,In_284,In_847);
nor U4543 (N_4543,In_85,In_890);
nor U4544 (N_4544,In_934,In_782);
or U4545 (N_4545,In_754,In_836);
nor U4546 (N_4546,In_273,In_470);
nor U4547 (N_4547,In_29,In_208);
nand U4548 (N_4548,In_855,In_634);
or U4549 (N_4549,In_949,In_797);
xor U4550 (N_4550,In_461,In_255);
or U4551 (N_4551,In_942,In_47);
and U4552 (N_4552,In_841,In_436);
xor U4553 (N_4553,In_845,In_306);
xor U4554 (N_4554,In_508,In_379);
or U4555 (N_4555,In_816,In_472);
nor U4556 (N_4556,In_51,In_664);
xnor U4557 (N_4557,In_58,In_631);
xor U4558 (N_4558,In_799,In_920);
or U4559 (N_4559,In_371,In_12);
xnor U4560 (N_4560,In_300,In_81);
xnor U4561 (N_4561,In_218,In_216);
nor U4562 (N_4562,In_312,In_464);
nor U4563 (N_4563,In_428,In_66);
and U4564 (N_4564,In_121,In_31);
or U4565 (N_4565,In_827,In_965);
and U4566 (N_4566,In_540,In_581);
and U4567 (N_4567,In_162,In_302);
or U4568 (N_4568,In_803,In_953);
nor U4569 (N_4569,In_349,In_510);
nor U4570 (N_4570,In_443,In_716);
nor U4571 (N_4571,In_694,In_306);
or U4572 (N_4572,In_916,In_431);
xor U4573 (N_4573,In_511,In_910);
or U4574 (N_4574,In_917,In_785);
nand U4575 (N_4575,In_623,In_760);
nand U4576 (N_4576,In_192,In_427);
nand U4577 (N_4577,In_824,In_727);
and U4578 (N_4578,In_642,In_914);
or U4579 (N_4579,In_503,In_150);
or U4580 (N_4580,In_659,In_586);
nor U4581 (N_4581,In_964,In_120);
xnor U4582 (N_4582,In_901,In_559);
xnor U4583 (N_4583,In_544,In_353);
nand U4584 (N_4584,In_512,In_101);
nand U4585 (N_4585,In_673,In_968);
or U4586 (N_4586,In_743,In_330);
xor U4587 (N_4587,In_227,In_550);
nor U4588 (N_4588,In_754,In_637);
nand U4589 (N_4589,In_910,In_305);
or U4590 (N_4590,In_364,In_273);
nor U4591 (N_4591,In_109,In_510);
nor U4592 (N_4592,In_904,In_939);
nand U4593 (N_4593,In_643,In_145);
nand U4594 (N_4594,In_557,In_45);
or U4595 (N_4595,In_494,In_508);
nand U4596 (N_4596,In_460,In_969);
nor U4597 (N_4597,In_521,In_13);
xnor U4598 (N_4598,In_461,In_684);
nand U4599 (N_4599,In_764,In_83);
and U4600 (N_4600,In_340,In_50);
nor U4601 (N_4601,In_892,In_574);
nand U4602 (N_4602,In_265,In_451);
and U4603 (N_4603,In_535,In_674);
or U4604 (N_4604,In_920,In_262);
nor U4605 (N_4605,In_920,In_470);
or U4606 (N_4606,In_8,In_424);
and U4607 (N_4607,In_655,In_631);
xor U4608 (N_4608,In_913,In_841);
and U4609 (N_4609,In_893,In_672);
nor U4610 (N_4610,In_924,In_794);
xnor U4611 (N_4611,In_794,In_353);
nor U4612 (N_4612,In_58,In_898);
xnor U4613 (N_4613,In_804,In_102);
nand U4614 (N_4614,In_615,In_431);
nor U4615 (N_4615,In_60,In_153);
nand U4616 (N_4616,In_701,In_822);
and U4617 (N_4617,In_444,In_21);
nand U4618 (N_4618,In_772,In_110);
nand U4619 (N_4619,In_144,In_705);
nor U4620 (N_4620,In_352,In_50);
and U4621 (N_4621,In_323,In_726);
and U4622 (N_4622,In_685,In_106);
or U4623 (N_4623,In_295,In_219);
nor U4624 (N_4624,In_427,In_289);
nor U4625 (N_4625,In_894,In_94);
xnor U4626 (N_4626,In_193,In_476);
and U4627 (N_4627,In_244,In_727);
or U4628 (N_4628,In_428,In_887);
xor U4629 (N_4629,In_404,In_295);
nor U4630 (N_4630,In_508,In_966);
nand U4631 (N_4631,In_254,In_290);
nand U4632 (N_4632,In_183,In_795);
xnor U4633 (N_4633,In_961,In_288);
and U4634 (N_4634,In_390,In_205);
nand U4635 (N_4635,In_44,In_842);
and U4636 (N_4636,In_276,In_631);
nand U4637 (N_4637,In_950,In_888);
nand U4638 (N_4638,In_246,In_59);
or U4639 (N_4639,In_219,In_63);
or U4640 (N_4640,In_442,In_610);
nand U4641 (N_4641,In_406,In_131);
nor U4642 (N_4642,In_646,In_174);
xnor U4643 (N_4643,In_240,In_170);
xor U4644 (N_4644,In_598,In_829);
xor U4645 (N_4645,In_94,In_500);
xor U4646 (N_4646,In_426,In_107);
and U4647 (N_4647,In_336,In_524);
nor U4648 (N_4648,In_189,In_473);
or U4649 (N_4649,In_609,In_165);
and U4650 (N_4650,In_770,In_961);
nand U4651 (N_4651,In_788,In_473);
nand U4652 (N_4652,In_665,In_797);
or U4653 (N_4653,In_927,In_471);
nor U4654 (N_4654,In_248,In_747);
nor U4655 (N_4655,In_564,In_124);
nand U4656 (N_4656,In_528,In_397);
and U4657 (N_4657,In_206,In_552);
and U4658 (N_4658,In_595,In_467);
and U4659 (N_4659,In_962,In_358);
xor U4660 (N_4660,In_818,In_250);
nor U4661 (N_4661,In_538,In_792);
nor U4662 (N_4662,In_519,In_462);
or U4663 (N_4663,In_984,In_68);
nor U4664 (N_4664,In_854,In_618);
or U4665 (N_4665,In_258,In_40);
and U4666 (N_4666,In_279,In_222);
nor U4667 (N_4667,In_472,In_825);
nor U4668 (N_4668,In_854,In_301);
xnor U4669 (N_4669,In_312,In_745);
nand U4670 (N_4670,In_264,In_940);
or U4671 (N_4671,In_267,In_788);
or U4672 (N_4672,In_395,In_620);
xor U4673 (N_4673,In_929,In_486);
xor U4674 (N_4674,In_141,In_862);
xor U4675 (N_4675,In_669,In_303);
or U4676 (N_4676,In_267,In_343);
or U4677 (N_4677,In_637,In_680);
and U4678 (N_4678,In_351,In_592);
or U4679 (N_4679,In_601,In_382);
or U4680 (N_4680,In_129,In_982);
nor U4681 (N_4681,In_806,In_36);
xor U4682 (N_4682,In_73,In_105);
xor U4683 (N_4683,In_612,In_660);
xor U4684 (N_4684,In_492,In_533);
or U4685 (N_4685,In_102,In_750);
nor U4686 (N_4686,In_557,In_496);
xnor U4687 (N_4687,In_799,In_516);
xor U4688 (N_4688,In_420,In_797);
and U4689 (N_4689,In_887,In_134);
and U4690 (N_4690,In_781,In_466);
xnor U4691 (N_4691,In_402,In_363);
and U4692 (N_4692,In_860,In_414);
or U4693 (N_4693,In_922,In_8);
nand U4694 (N_4694,In_383,In_910);
or U4695 (N_4695,In_103,In_865);
nand U4696 (N_4696,In_837,In_592);
xnor U4697 (N_4697,In_224,In_144);
or U4698 (N_4698,In_551,In_728);
and U4699 (N_4699,In_409,In_988);
xnor U4700 (N_4700,In_946,In_581);
or U4701 (N_4701,In_109,In_336);
xor U4702 (N_4702,In_889,In_625);
nand U4703 (N_4703,In_699,In_257);
nand U4704 (N_4704,In_908,In_855);
or U4705 (N_4705,In_601,In_782);
nor U4706 (N_4706,In_898,In_879);
and U4707 (N_4707,In_281,In_850);
or U4708 (N_4708,In_386,In_823);
nand U4709 (N_4709,In_214,In_760);
nor U4710 (N_4710,In_473,In_676);
or U4711 (N_4711,In_415,In_625);
or U4712 (N_4712,In_524,In_431);
nor U4713 (N_4713,In_939,In_240);
nand U4714 (N_4714,In_33,In_516);
or U4715 (N_4715,In_150,In_953);
xnor U4716 (N_4716,In_962,In_297);
and U4717 (N_4717,In_288,In_767);
nand U4718 (N_4718,In_226,In_822);
or U4719 (N_4719,In_166,In_320);
or U4720 (N_4720,In_925,In_61);
and U4721 (N_4721,In_450,In_456);
nand U4722 (N_4722,In_317,In_205);
nor U4723 (N_4723,In_412,In_82);
nor U4724 (N_4724,In_66,In_763);
nor U4725 (N_4725,In_183,In_15);
or U4726 (N_4726,In_695,In_745);
or U4727 (N_4727,In_420,In_653);
and U4728 (N_4728,In_791,In_464);
nor U4729 (N_4729,In_140,In_992);
or U4730 (N_4730,In_450,In_554);
and U4731 (N_4731,In_529,In_653);
and U4732 (N_4732,In_203,In_561);
nand U4733 (N_4733,In_627,In_104);
or U4734 (N_4734,In_74,In_909);
nor U4735 (N_4735,In_980,In_525);
or U4736 (N_4736,In_406,In_986);
nand U4737 (N_4737,In_626,In_101);
xnor U4738 (N_4738,In_949,In_558);
and U4739 (N_4739,In_907,In_270);
nand U4740 (N_4740,In_480,In_636);
nand U4741 (N_4741,In_184,In_554);
xor U4742 (N_4742,In_176,In_524);
nand U4743 (N_4743,In_401,In_996);
xnor U4744 (N_4744,In_392,In_741);
nor U4745 (N_4745,In_362,In_792);
or U4746 (N_4746,In_539,In_678);
or U4747 (N_4747,In_127,In_133);
or U4748 (N_4748,In_999,In_685);
nor U4749 (N_4749,In_905,In_793);
or U4750 (N_4750,In_313,In_583);
nor U4751 (N_4751,In_632,In_371);
and U4752 (N_4752,In_683,In_858);
or U4753 (N_4753,In_180,In_994);
nor U4754 (N_4754,In_534,In_579);
nor U4755 (N_4755,In_122,In_816);
or U4756 (N_4756,In_691,In_789);
and U4757 (N_4757,In_603,In_993);
nand U4758 (N_4758,In_161,In_26);
or U4759 (N_4759,In_179,In_963);
xnor U4760 (N_4760,In_989,In_690);
nor U4761 (N_4761,In_854,In_210);
xor U4762 (N_4762,In_607,In_481);
and U4763 (N_4763,In_790,In_131);
and U4764 (N_4764,In_711,In_263);
nand U4765 (N_4765,In_704,In_313);
or U4766 (N_4766,In_834,In_623);
xor U4767 (N_4767,In_494,In_768);
nor U4768 (N_4768,In_993,In_626);
and U4769 (N_4769,In_503,In_881);
or U4770 (N_4770,In_895,In_885);
or U4771 (N_4771,In_475,In_504);
and U4772 (N_4772,In_497,In_127);
or U4773 (N_4773,In_672,In_754);
nor U4774 (N_4774,In_261,In_542);
nand U4775 (N_4775,In_838,In_628);
or U4776 (N_4776,In_974,In_106);
or U4777 (N_4777,In_554,In_206);
or U4778 (N_4778,In_549,In_558);
xnor U4779 (N_4779,In_84,In_178);
nand U4780 (N_4780,In_416,In_410);
xnor U4781 (N_4781,In_709,In_265);
nand U4782 (N_4782,In_596,In_106);
or U4783 (N_4783,In_473,In_643);
nor U4784 (N_4784,In_827,In_228);
xnor U4785 (N_4785,In_880,In_464);
xor U4786 (N_4786,In_846,In_120);
or U4787 (N_4787,In_921,In_214);
xnor U4788 (N_4788,In_689,In_182);
nor U4789 (N_4789,In_260,In_792);
or U4790 (N_4790,In_352,In_294);
nor U4791 (N_4791,In_489,In_208);
or U4792 (N_4792,In_71,In_331);
or U4793 (N_4793,In_864,In_275);
and U4794 (N_4794,In_391,In_329);
or U4795 (N_4795,In_911,In_846);
xor U4796 (N_4796,In_128,In_71);
nand U4797 (N_4797,In_439,In_553);
nand U4798 (N_4798,In_865,In_170);
and U4799 (N_4799,In_745,In_72);
and U4800 (N_4800,In_654,In_178);
xnor U4801 (N_4801,In_480,In_257);
nand U4802 (N_4802,In_61,In_298);
nand U4803 (N_4803,In_564,In_299);
xor U4804 (N_4804,In_254,In_593);
nor U4805 (N_4805,In_137,In_860);
and U4806 (N_4806,In_870,In_980);
nor U4807 (N_4807,In_472,In_389);
and U4808 (N_4808,In_157,In_672);
nand U4809 (N_4809,In_951,In_281);
or U4810 (N_4810,In_288,In_515);
xor U4811 (N_4811,In_739,In_599);
or U4812 (N_4812,In_822,In_441);
nor U4813 (N_4813,In_559,In_865);
and U4814 (N_4814,In_406,In_132);
nand U4815 (N_4815,In_121,In_290);
nand U4816 (N_4816,In_254,In_353);
xor U4817 (N_4817,In_691,In_761);
nand U4818 (N_4818,In_359,In_620);
and U4819 (N_4819,In_31,In_109);
nand U4820 (N_4820,In_20,In_315);
or U4821 (N_4821,In_634,In_710);
nand U4822 (N_4822,In_542,In_110);
nand U4823 (N_4823,In_665,In_890);
nor U4824 (N_4824,In_288,In_65);
or U4825 (N_4825,In_772,In_628);
nand U4826 (N_4826,In_913,In_332);
or U4827 (N_4827,In_223,In_549);
xnor U4828 (N_4828,In_480,In_242);
or U4829 (N_4829,In_41,In_553);
nor U4830 (N_4830,In_113,In_102);
xnor U4831 (N_4831,In_966,In_985);
nor U4832 (N_4832,In_789,In_991);
or U4833 (N_4833,In_226,In_920);
nor U4834 (N_4834,In_600,In_898);
xnor U4835 (N_4835,In_208,In_643);
xor U4836 (N_4836,In_751,In_896);
or U4837 (N_4837,In_99,In_444);
xnor U4838 (N_4838,In_465,In_999);
and U4839 (N_4839,In_936,In_550);
nor U4840 (N_4840,In_22,In_907);
or U4841 (N_4841,In_629,In_445);
xnor U4842 (N_4842,In_12,In_611);
nor U4843 (N_4843,In_694,In_612);
nand U4844 (N_4844,In_441,In_10);
xnor U4845 (N_4845,In_433,In_664);
or U4846 (N_4846,In_872,In_646);
xor U4847 (N_4847,In_850,In_6);
and U4848 (N_4848,In_826,In_624);
and U4849 (N_4849,In_724,In_512);
and U4850 (N_4850,In_654,In_871);
nand U4851 (N_4851,In_762,In_639);
and U4852 (N_4852,In_478,In_564);
or U4853 (N_4853,In_155,In_588);
or U4854 (N_4854,In_198,In_950);
and U4855 (N_4855,In_867,In_305);
xor U4856 (N_4856,In_314,In_657);
nand U4857 (N_4857,In_699,In_57);
xor U4858 (N_4858,In_332,In_852);
or U4859 (N_4859,In_868,In_248);
or U4860 (N_4860,In_731,In_218);
or U4861 (N_4861,In_503,In_511);
or U4862 (N_4862,In_594,In_176);
nor U4863 (N_4863,In_513,In_537);
nor U4864 (N_4864,In_623,In_542);
or U4865 (N_4865,In_608,In_169);
and U4866 (N_4866,In_787,In_903);
nand U4867 (N_4867,In_814,In_344);
nand U4868 (N_4868,In_858,In_958);
xor U4869 (N_4869,In_599,In_687);
or U4870 (N_4870,In_862,In_741);
or U4871 (N_4871,In_301,In_154);
xor U4872 (N_4872,In_64,In_912);
nand U4873 (N_4873,In_938,In_444);
xor U4874 (N_4874,In_47,In_720);
and U4875 (N_4875,In_953,In_956);
and U4876 (N_4876,In_434,In_574);
or U4877 (N_4877,In_556,In_523);
xnor U4878 (N_4878,In_406,In_714);
nor U4879 (N_4879,In_257,In_924);
nor U4880 (N_4880,In_446,In_439);
nor U4881 (N_4881,In_260,In_529);
or U4882 (N_4882,In_343,In_25);
xnor U4883 (N_4883,In_447,In_187);
or U4884 (N_4884,In_479,In_922);
nand U4885 (N_4885,In_843,In_178);
and U4886 (N_4886,In_701,In_841);
nand U4887 (N_4887,In_676,In_789);
and U4888 (N_4888,In_765,In_395);
nor U4889 (N_4889,In_606,In_428);
and U4890 (N_4890,In_140,In_417);
and U4891 (N_4891,In_228,In_985);
or U4892 (N_4892,In_173,In_698);
nand U4893 (N_4893,In_637,In_970);
nand U4894 (N_4894,In_74,In_757);
or U4895 (N_4895,In_318,In_615);
nor U4896 (N_4896,In_24,In_603);
nor U4897 (N_4897,In_943,In_976);
nand U4898 (N_4898,In_697,In_494);
nor U4899 (N_4899,In_111,In_495);
nand U4900 (N_4900,In_770,In_210);
nor U4901 (N_4901,In_914,In_590);
xor U4902 (N_4902,In_109,In_501);
nor U4903 (N_4903,In_219,In_528);
nor U4904 (N_4904,In_547,In_442);
and U4905 (N_4905,In_40,In_365);
and U4906 (N_4906,In_987,In_519);
or U4907 (N_4907,In_16,In_300);
nand U4908 (N_4908,In_344,In_184);
and U4909 (N_4909,In_358,In_917);
or U4910 (N_4910,In_428,In_889);
nor U4911 (N_4911,In_422,In_506);
nand U4912 (N_4912,In_309,In_492);
and U4913 (N_4913,In_656,In_7);
nand U4914 (N_4914,In_254,In_583);
xor U4915 (N_4915,In_615,In_990);
and U4916 (N_4916,In_800,In_382);
and U4917 (N_4917,In_231,In_763);
or U4918 (N_4918,In_663,In_56);
nor U4919 (N_4919,In_668,In_500);
nand U4920 (N_4920,In_970,In_378);
or U4921 (N_4921,In_433,In_696);
and U4922 (N_4922,In_585,In_65);
nor U4923 (N_4923,In_268,In_540);
xnor U4924 (N_4924,In_791,In_601);
nand U4925 (N_4925,In_8,In_256);
and U4926 (N_4926,In_66,In_384);
and U4927 (N_4927,In_59,In_695);
or U4928 (N_4928,In_605,In_183);
and U4929 (N_4929,In_902,In_15);
nor U4930 (N_4930,In_824,In_116);
xor U4931 (N_4931,In_336,In_511);
xor U4932 (N_4932,In_521,In_985);
or U4933 (N_4933,In_82,In_361);
nor U4934 (N_4934,In_333,In_867);
nand U4935 (N_4935,In_98,In_587);
or U4936 (N_4936,In_112,In_161);
nor U4937 (N_4937,In_696,In_443);
nand U4938 (N_4938,In_747,In_545);
and U4939 (N_4939,In_282,In_791);
and U4940 (N_4940,In_278,In_704);
xnor U4941 (N_4941,In_489,In_369);
xor U4942 (N_4942,In_253,In_957);
or U4943 (N_4943,In_205,In_513);
or U4944 (N_4944,In_929,In_553);
nand U4945 (N_4945,In_732,In_119);
or U4946 (N_4946,In_411,In_762);
xor U4947 (N_4947,In_146,In_357);
xnor U4948 (N_4948,In_810,In_251);
or U4949 (N_4949,In_916,In_566);
xnor U4950 (N_4950,In_834,In_844);
and U4951 (N_4951,In_335,In_17);
xnor U4952 (N_4952,In_446,In_964);
nand U4953 (N_4953,In_159,In_694);
and U4954 (N_4954,In_931,In_583);
and U4955 (N_4955,In_862,In_44);
or U4956 (N_4956,In_211,In_437);
nor U4957 (N_4957,In_571,In_429);
and U4958 (N_4958,In_818,In_90);
xnor U4959 (N_4959,In_77,In_831);
nand U4960 (N_4960,In_4,In_575);
and U4961 (N_4961,In_92,In_577);
xor U4962 (N_4962,In_546,In_484);
or U4963 (N_4963,In_629,In_78);
nor U4964 (N_4964,In_327,In_294);
nand U4965 (N_4965,In_684,In_314);
or U4966 (N_4966,In_172,In_935);
or U4967 (N_4967,In_702,In_296);
and U4968 (N_4968,In_191,In_710);
nand U4969 (N_4969,In_212,In_886);
and U4970 (N_4970,In_561,In_28);
or U4971 (N_4971,In_814,In_992);
nor U4972 (N_4972,In_90,In_124);
or U4973 (N_4973,In_422,In_521);
xnor U4974 (N_4974,In_599,In_443);
or U4975 (N_4975,In_830,In_405);
or U4976 (N_4976,In_874,In_551);
xor U4977 (N_4977,In_806,In_248);
nand U4978 (N_4978,In_81,In_315);
or U4979 (N_4979,In_392,In_688);
xnor U4980 (N_4980,In_412,In_439);
nor U4981 (N_4981,In_50,In_213);
and U4982 (N_4982,In_399,In_719);
and U4983 (N_4983,In_480,In_409);
nor U4984 (N_4984,In_194,In_125);
nor U4985 (N_4985,In_450,In_486);
nor U4986 (N_4986,In_662,In_538);
or U4987 (N_4987,In_721,In_906);
or U4988 (N_4988,In_436,In_427);
nor U4989 (N_4989,In_108,In_159);
xor U4990 (N_4990,In_430,In_236);
nand U4991 (N_4991,In_416,In_764);
or U4992 (N_4992,In_277,In_530);
nor U4993 (N_4993,In_779,In_645);
or U4994 (N_4994,In_309,In_498);
xor U4995 (N_4995,In_485,In_991);
and U4996 (N_4996,In_787,In_254);
and U4997 (N_4997,In_964,In_880);
nand U4998 (N_4998,In_145,In_418);
nor U4999 (N_4999,In_851,In_387);
xor U5000 (N_5000,N_2244,N_1024);
and U5001 (N_5001,N_956,N_2687);
or U5002 (N_5002,N_4955,N_4619);
nand U5003 (N_5003,N_1657,N_2147);
and U5004 (N_5004,N_1032,N_3026);
nor U5005 (N_5005,N_2018,N_4943);
and U5006 (N_5006,N_3776,N_3916);
xnor U5007 (N_5007,N_2052,N_2630);
xnor U5008 (N_5008,N_486,N_725);
or U5009 (N_5009,N_1403,N_3389);
or U5010 (N_5010,N_2726,N_3312);
nor U5011 (N_5011,N_1683,N_322);
and U5012 (N_5012,N_227,N_1590);
nor U5013 (N_5013,N_3096,N_4048);
nand U5014 (N_5014,N_4659,N_4354);
and U5015 (N_5015,N_1706,N_4568);
nand U5016 (N_5016,N_3476,N_39);
xor U5017 (N_5017,N_1029,N_4382);
and U5018 (N_5018,N_2287,N_642);
and U5019 (N_5019,N_4475,N_3162);
and U5020 (N_5020,N_1294,N_367);
nor U5021 (N_5021,N_1651,N_2870);
or U5022 (N_5022,N_29,N_4690);
xnor U5023 (N_5023,N_2465,N_4487);
and U5024 (N_5024,N_4915,N_801);
nor U5025 (N_5025,N_3236,N_4812);
and U5026 (N_5026,N_2108,N_677);
nor U5027 (N_5027,N_3483,N_2528);
xor U5028 (N_5028,N_1568,N_3251);
nor U5029 (N_5029,N_2134,N_804);
or U5030 (N_5030,N_3185,N_4790);
nand U5031 (N_5031,N_2047,N_3024);
and U5032 (N_5032,N_1866,N_2948);
or U5033 (N_5033,N_4167,N_1756);
nor U5034 (N_5034,N_4011,N_1816);
and U5035 (N_5035,N_2526,N_3214);
xnor U5036 (N_5036,N_307,N_2040);
xnor U5037 (N_5037,N_3689,N_3232);
and U5038 (N_5038,N_4855,N_1238);
nor U5039 (N_5039,N_1536,N_1502);
nor U5040 (N_5040,N_1445,N_640);
xnor U5041 (N_5041,N_258,N_3374);
or U5042 (N_5042,N_4424,N_2203);
nand U5043 (N_5043,N_4071,N_21);
or U5044 (N_5044,N_4570,N_4821);
xnor U5045 (N_5045,N_3675,N_4119);
xnor U5046 (N_5046,N_3976,N_1615);
and U5047 (N_5047,N_4963,N_829);
or U5048 (N_5048,N_4617,N_2413);
nor U5049 (N_5049,N_1336,N_4344);
and U5050 (N_5050,N_3881,N_1687);
nand U5051 (N_5051,N_4488,N_3158);
or U5052 (N_5052,N_900,N_3225);
and U5053 (N_5053,N_4244,N_933);
xor U5054 (N_5054,N_106,N_1088);
nand U5055 (N_5055,N_3526,N_4358);
and U5056 (N_5056,N_4432,N_2605);
xor U5057 (N_5057,N_810,N_3194);
nor U5058 (N_5058,N_2124,N_3625);
nand U5059 (N_5059,N_4585,N_3636);
or U5060 (N_5060,N_4910,N_2250);
and U5061 (N_5061,N_4852,N_2639);
or U5062 (N_5062,N_910,N_1533);
nor U5063 (N_5063,N_4947,N_2997);
or U5064 (N_5064,N_2770,N_842);
xnor U5065 (N_5065,N_503,N_1196);
or U5066 (N_5066,N_4390,N_4190);
and U5067 (N_5067,N_2354,N_1211);
or U5068 (N_5068,N_2103,N_3501);
xor U5069 (N_5069,N_2114,N_3275);
nor U5070 (N_5070,N_1569,N_1558);
xor U5071 (N_5071,N_1762,N_415);
or U5072 (N_5072,N_319,N_2030);
or U5073 (N_5073,N_114,N_468);
xnor U5074 (N_5074,N_669,N_1296);
or U5075 (N_5075,N_701,N_2711);
xor U5076 (N_5076,N_2425,N_4666);
or U5077 (N_5077,N_2824,N_2332);
xnor U5078 (N_5078,N_492,N_1595);
and U5079 (N_5079,N_1636,N_5);
nor U5080 (N_5080,N_3363,N_2903);
nor U5081 (N_5081,N_1660,N_10);
and U5082 (N_5082,N_353,N_68);
and U5083 (N_5083,N_331,N_3553);
xor U5084 (N_5084,N_1970,N_4802);
or U5085 (N_5085,N_2340,N_1551);
or U5086 (N_5086,N_937,N_4891);
xor U5087 (N_5087,N_2923,N_2335);
or U5088 (N_5088,N_2640,N_1061);
or U5089 (N_5089,N_3375,N_3603);
and U5090 (N_5090,N_2441,N_2145);
and U5091 (N_5091,N_2602,N_3186);
xor U5092 (N_5092,N_3392,N_2373);
xnor U5093 (N_5093,N_1072,N_2468);
xnor U5094 (N_5094,N_3727,N_970);
or U5095 (N_5095,N_4439,N_4776);
nand U5096 (N_5096,N_3690,N_1310);
and U5097 (N_5097,N_621,N_1912);
or U5098 (N_5098,N_233,N_365);
nand U5099 (N_5099,N_2178,N_4663);
nor U5100 (N_5100,N_4333,N_789);
nor U5101 (N_5101,N_619,N_4902);
or U5102 (N_5102,N_2628,N_1812);
and U5103 (N_5103,N_1725,N_1875);
nor U5104 (N_5104,N_2182,N_2080);
and U5105 (N_5105,N_3958,N_4597);
or U5106 (N_5106,N_1357,N_1891);
xor U5107 (N_5107,N_4974,N_3330);
xor U5108 (N_5108,N_722,N_3406);
nand U5109 (N_5109,N_2918,N_3567);
and U5110 (N_5110,N_2621,N_1934);
xor U5111 (N_5111,N_3370,N_1402);
nor U5112 (N_5112,N_4882,N_3493);
or U5113 (N_5113,N_3545,N_388);
and U5114 (N_5114,N_2159,N_4691);
or U5115 (N_5115,N_4170,N_4589);
nor U5116 (N_5116,N_4272,N_3432);
nor U5117 (N_5117,N_1216,N_4627);
or U5118 (N_5118,N_2459,N_3914);
xnor U5119 (N_5119,N_2837,N_2345);
nor U5120 (N_5120,N_4669,N_4117);
nand U5121 (N_5121,N_924,N_3372);
or U5122 (N_5122,N_4559,N_2754);
and U5123 (N_5123,N_766,N_4295);
xnor U5124 (N_5124,N_4697,N_3937);
and U5125 (N_5125,N_4962,N_895);
or U5126 (N_5126,N_2977,N_2228);
or U5127 (N_5127,N_1579,N_4115);
or U5128 (N_5128,N_3620,N_1822);
nand U5129 (N_5129,N_4430,N_3997);
nand U5130 (N_5130,N_663,N_3640);
nand U5131 (N_5131,N_1534,N_1721);
xor U5132 (N_5132,N_514,N_3068);
nor U5133 (N_5133,N_4534,N_3775);
nand U5134 (N_5134,N_3456,N_4046);
xor U5135 (N_5135,N_4287,N_682);
nand U5136 (N_5136,N_3939,N_1442);
or U5137 (N_5137,N_3490,N_2667);
xor U5138 (N_5138,N_382,N_694);
or U5139 (N_5139,N_2790,N_3845);
and U5140 (N_5140,N_1757,N_2949);
xor U5141 (N_5141,N_3717,N_285);
xnor U5142 (N_5142,N_36,N_1666);
or U5143 (N_5143,N_195,N_750);
nand U5144 (N_5144,N_294,N_4880);
nor U5145 (N_5145,N_3030,N_2294);
xnor U5146 (N_5146,N_2663,N_3504);
and U5147 (N_5147,N_324,N_1532);
and U5148 (N_5148,N_1159,N_2282);
nor U5149 (N_5149,N_2449,N_1184);
and U5150 (N_5150,N_3742,N_1952);
nor U5151 (N_5151,N_4015,N_4448);
nor U5152 (N_5152,N_1035,N_3781);
xor U5153 (N_5153,N_2657,N_3266);
and U5154 (N_5154,N_1472,N_4041);
and U5155 (N_5155,N_3136,N_1859);
nand U5156 (N_5156,N_184,N_1105);
xnor U5157 (N_5157,N_4942,N_460);
nor U5158 (N_5158,N_4131,N_988);
xnor U5159 (N_5159,N_2198,N_3050);
xnor U5160 (N_5160,N_2987,N_2435);
or U5161 (N_5161,N_4851,N_2753);
nor U5162 (N_5162,N_2729,N_256);
nand U5163 (N_5163,N_614,N_3261);
or U5164 (N_5164,N_3182,N_1741);
nand U5165 (N_5165,N_2169,N_2473);
or U5166 (N_5166,N_275,N_728);
or U5167 (N_5167,N_2012,N_1152);
or U5168 (N_5168,N_1412,N_1627);
nand U5169 (N_5169,N_414,N_3435);
and U5170 (N_5170,N_2772,N_1398);
or U5171 (N_5171,N_3272,N_2877);
xor U5172 (N_5172,N_643,N_3103);
xnor U5173 (N_5173,N_1702,N_18);
or U5174 (N_5174,N_1526,N_885);
or U5175 (N_5175,N_1538,N_4370);
nand U5176 (N_5176,N_2410,N_4785);
xor U5177 (N_5177,N_1454,N_4874);
or U5178 (N_5178,N_3972,N_2185);
nor U5179 (N_5179,N_2941,N_869);
xor U5180 (N_5180,N_3129,N_4065);
nand U5181 (N_5181,N_2454,N_884);
and U5182 (N_5182,N_1796,N_3498);
and U5183 (N_5183,N_4049,N_202);
nor U5184 (N_5184,N_1933,N_2204);
and U5185 (N_5185,N_1194,N_16);
nor U5186 (N_5186,N_3209,N_4379);
nand U5187 (N_5187,N_3405,N_3280);
or U5188 (N_5188,N_550,N_3863);
nor U5189 (N_5189,N_3040,N_3323);
or U5190 (N_5190,N_205,N_4141);
nand U5191 (N_5191,N_4747,N_4936);
and U5192 (N_5192,N_2716,N_4361);
and U5193 (N_5193,N_4805,N_2810);
nand U5194 (N_5194,N_781,N_1737);
and U5195 (N_5195,N_2847,N_4335);
or U5196 (N_5196,N_1893,N_3536);
nand U5197 (N_5197,N_1118,N_939);
nand U5198 (N_5198,N_4086,N_4620);
and U5199 (N_5199,N_1574,N_4331);
nor U5200 (N_5200,N_4284,N_3941);
nor U5201 (N_5201,N_2952,N_4426);
nor U5202 (N_5202,N_786,N_2533);
and U5203 (N_5203,N_4464,N_4098);
or U5204 (N_5204,N_2635,N_662);
xor U5205 (N_5205,N_2170,N_2158);
xnor U5206 (N_5206,N_2298,N_855);
and U5207 (N_5207,N_4780,N_4401);
nor U5208 (N_5208,N_4770,N_390);
nand U5209 (N_5209,N_1860,N_208);
or U5210 (N_5210,N_4712,N_4843);
nand U5211 (N_5211,N_3509,N_4093);
or U5212 (N_5212,N_1305,N_4266);
or U5213 (N_5213,N_2218,N_312);
nand U5214 (N_5214,N_4879,N_209);
and U5215 (N_5215,N_1342,N_4723);
xnor U5216 (N_5216,N_1940,N_2906);
nor U5217 (N_5217,N_4923,N_3685);
nand U5218 (N_5218,N_1544,N_4908);
nand U5219 (N_5219,N_429,N_2327);
and U5220 (N_5220,N_975,N_3758);
or U5221 (N_5221,N_4083,N_3656);
xor U5222 (N_5222,N_2365,N_3173);
xnor U5223 (N_5223,N_2448,N_4479);
and U5224 (N_5224,N_1186,N_182);
nand U5225 (N_5225,N_3960,N_433);
nand U5226 (N_5226,N_1167,N_549);
nand U5227 (N_5227,N_2236,N_4105);
nor U5228 (N_5228,N_1504,N_3098);
nand U5229 (N_5229,N_4553,N_2069);
or U5230 (N_5230,N_217,N_4765);
xor U5231 (N_5231,N_3956,N_2302);
xnor U5232 (N_5232,N_2755,N_447);
and U5233 (N_5233,N_3286,N_4660);
xnor U5234 (N_5234,N_2890,N_3329);
nand U5235 (N_5235,N_3653,N_2280);
xor U5236 (N_5236,N_1197,N_2437);
nand U5237 (N_5237,N_3179,N_3320);
xnor U5238 (N_5238,N_1381,N_3168);
or U5239 (N_5239,N_4219,N_1783);
or U5240 (N_5240,N_1518,N_866);
and U5241 (N_5241,N_2190,N_4547);
nor U5242 (N_5242,N_3293,N_1347);
nand U5243 (N_5243,N_2133,N_3304);
and U5244 (N_5244,N_2874,N_968);
nand U5245 (N_5245,N_4248,N_3694);
xor U5246 (N_5246,N_878,N_4494);
xor U5247 (N_5247,N_1591,N_3593);
or U5248 (N_5248,N_1281,N_531);
and U5249 (N_5249,N_3904,N_4321);
nor U5250 (N_5250,N_4311,N_3786);
or U5251 (N_5251,N_1332,N_2943);
xnor U5252 (N_5252,N_3449,N_4473);
and U5253 (N_5253,N_3169,N_3757);
nor U5254 (N_5254,N_3979,N_389);
or U5255 (N_5255,N_1172,N_1503);
and U5256 (N_5256,N_1144,N_3227);
xnor U5257 (N_5257,N_902,N_4308);
xor U5258 (N_5258,N_120,N_4214);
xnor U5259 (N_5259,N_360,N_4252);
and U5260 (N_5260,N_3079,N_299);
and U5261 (N_5261,N_363,N_309);
and U5262 (N_5262,N_3877,N_2125);
or U5263 (N_5263,N_807,N_2054);
or U5264 (N_5264,N_4057,N_3166);
or U5265 (N_5265,N_3475,N_4667);
nand U5266 (N_5266,N_301,N_3990);
and U5267 (N_5267,N_890,N_1941);
nor U5268 (N_5268,N_1069,N_1451);
nor U5269 (N_5269,N_2234,N_3884);
or U5270 (N_5270,N_3478,N_4341);
nand U5271 (N_5271,N_4823,N_830);
or U5272 (N_5272,N_4841,N_2764);
nor U5273 (N_5273,N_80,N_164);
and U5274 (N_5274,N_478,N_3768);
nand U5275 (N_5275,N_3451,N_2721);
or U5276 (N_5276,N_3535,N_2458);
nand U5277 (N_5277,N_2434,N_4262);
nor U5278 (N_5278,N_3299,N_2175);
nand U5279 (N_5279,N_4745,N_989);
nand U5280 (N_5280,N_2208,N_831);
xor U5281 (N_5281,N_3302,N_770);
nor U5282 (N_5282,N_1290,N_3891);
and U5283 (N_5283,N_4800,N_169);
nor U5284 (N_5284,N_718,N_2537);
or U5285 (N_5285,N_3199,N_4540);
and U5286 (N_5286,N_3740,N_1292);
or U5287 (N_5287,N_4625,N_73);
nor U5288 (N_5288,N_1039,N_3908);
nor U5289 (N_5289,N_4183,N_4175);
and U5290 (N_5290,N_723,N_77);
and U5291 (N_5291,N_4508,N_441);
or U5292 (N_5292,N_4134,N_3797);
and U5293 (N_5293,N_282,N_4005);
or U5294 (N_5294,N_4414,N_3659);
nor U5295 (N_5295,N_849,N_610);
xnor U5296 (N_5296,N_624,N_576);
nand U5297 (N_5297,N_1215,N_1539);
nand U5298 (N_5298,N_2757,N_4708);
and U5299 (N_5299,N_3719,N_4522);
and U5300 (N_5300,N_2507,N_1549);
nor U5301 (N_5301,N_1208,N_4655);
nor U5302 (N_5302,N_1164,N_1314);
or U5303 (N_5303,N_384,N_1075);
xnor U5304 (N_5304,N_1852,N_4767);
nor U5305 (N_5305,N_1902,N_2007);
or U5306 (N_5306,N_2440,N_1733);
and U5307 (N_5307,N_86,N_4147);
nor U5308 (N_5308,N_4312,N_735);
nand U5309 (N_5309,N_876,N_3357);
nor U5310 (N_5310,N_3539,N_3629);
nand U5311 (N_5311,N_4634,N_923);
nor U5312 (N_5312,N_3421,N_224);
nand U5313 (N_5313,N_3083,N_3837);
nor U5314 (N_5314,N_4340,N_1861);
xor U5315 (N_5315,N_2738,N_2181);
xor U5316 (N_5316,N_3041,N_4729);
or U5317 (N_5317,N_2596,N_2419);
nand U5318 (N_5318,N_4072,N_3245);
xnor U5319 (N_5319,N_3815,N_438);
or U5320 (N_5320,N_304,N_730);
and U5321 (N_5321,N_2820,N_1643);
and U5322 (N_5322,N_4433,N_1594);
and U5323 (N_5323,N_3813,N_4595);
nand U5324 (N_5324,N_4192,N_3167);
xnor U5325 (N_5325,N_4037,N_2712);
xor U5326 (N_5326,N_2362,N_4246);
xnor U5327 (N_5327,N_374,N_269);
or U5328 (N_5328,N_4647,N_4889);
nor U5329 (N_5329,N_1236,N_4378);
nand U5330 (N_5330,N_4656,N_613);
and U5331 (N_5331,N_3969,N_4773);
or U5332 (N_5332,N_4109,N_1014);
nand U5333 (N_5333,N_496,N_3454);
and U5334 (N_5334,N_3601,N_3574);
xnor U5335 (N_5335,N_1221,N_2442);
and U5336 (N_5336,N_3126,N_4);
or U5337 (N_5337,N_2768,N_3326);
and U5338 (N_5338,N_4689,N_1896);
and U5339 (N_5339,N_2295,N_630);
and U5340 (N_5340,N_4478,N_2380);
nor U5341 (N_5341,N_4803,N_4089);
and U5342 (N_5342,N_1045,N_3565);
nor U5343 (N_5343,N_356,N_1647);
and U5344 (N_5344,N_1570,N_2759);
or U5345 (N_5345,N_2981,N_3922);
xor U5346 (N_5346,N_1301,N_2659);
xnor U5347 (N_5347,N_2004,N_2252);
xor U5348 (N_5348,N_124,N_2128);
nand U5349 (N_5349,N_2676,N_1366);
nand U5350 (N_5350,N_3200,N_2389);
and U5351 (N_5351,N_3384,N_1958);
or U5352 (N_5352,N_3089,N_705);
xnor U5353 (N_5353,N_4829,N_605);
nand U5354 (N_5354,N_4436,N_3390);
nor U5355 (N_5355,N_2618,N_4504);
and U5356 (N_5356,N_3839,N_1942);
and U5357 (N_5357,N_584,N_4929);
and U5358 (N_5358,N_3784,N_1331);
or U5359 (N_5359,N_4493,N_4750);
and U5360 (N_5360,N_2557,N_2819);
or U5361 (N_5361,N_2213,N_2115);
nand U5362 (N_5362,N_2205,N_4067);
nor U5363 (N_5363,N_2829,N_1419);
and U5364 (N_5364,N_736,N_3688);
or U5365 (N_5365,N_3521,N_4772);
nor U5366 (N_5366,N_1821,N_2786);
or U5367 (N_5367,N_4536,N_4913);
nand U5368 (N_5368,N_3844,N_2140);
xor U5369 (N_5369,N_4886,N_4637);
or U5370 (N_5370,N_4768,N_4241);
nand U5371 (N_5371,N_1592,N_1112);
nand U5372 (N_5372,N_402,N_1936);
nor U5373 (N_5373,N_1777,N_3743);
and U5374 (N_5374,N_4292,N_4918);
or U5375 (N_5375,N_3646,N_3613);
or U5376 (N_5376,N_4665,N_4171);
nor U5377 (N_5377,N_2075,N_783);
nand U5378 (N_5378,N_1593,N_51);
or U5379 (N_5379,N_2576,N_434);
xor U5380 (N_5380,N_2223,N_2868);
nor U5381 (N_5381,N_2098,N_1603);
xnor U5382 (N_5382,N_1397,N_4063);
and U5383 (N_5383,N_3788,N_727);
xnor U5384 (N_5384,N_4416,N_2805);
nor U5385 (N_5385,N_1935,N_2342);
xor U5386 (N_5386,N_3745,N_4813);
and U5387 (N_5387,N_343,N_4845);
nand U5388 (N_5388,N_3680,N_2900);
xnor U5389 (N_5389,N_4693,N_4054);
and U5390 (N_5390,N_4546,N_1448);
xor U5391 (N_5391,N_901,N_552);
nor U5392 (N_5392,N_3107,N_1277);
xnor U5393 (N_5393,N_4236,N_2050);
nor U5394 (N_5394,N_4164,N_1011);
and U5395 (N_5395,N_2778,N_3631);
nand U5396 (N_5396,N_2015,N_3519);
nor U5397 (N_5397,N_355,N_1956);
xnor U5398 (N_5398,N_4956,N_741);
and U5399 (N_5399,N_3269,N_2256);
and U5400 (N_5400,N_4728,N_1051);
xnor U5401 (N_5401,N_2443,N_874);
or U5402 (N_5402,N_1851,N_1825);
or U5403 (N_5403,N_2727,N_4569);
or U5404 (N_5404,N_2680,N_4298);
nand U5405 (N_5405,N_2623,N_3623);
and U5406 (N_5406,N_2285,N_3159);
xnor U5407 (N_5407,N_1694,N_2130);
or U5408 (N_5408,N_3181,N_2366);
xor U5409 (N_5409,N_1966,N_1258);
nand U5410 (N_5410,N_2136,N_3996);
and U5411 (N_5411,N_4463,N_957);
nand U5412 (N_5412,N_2227,N_3282);
or U5413 (N_5413,N_1855,N_1103);
nand U5414 (N_5414,N_3912,N_3953);
and U5415 (N_5415,N_2081,N_1265);
or U5416 (N_5416,N_444,N_1053);
or U5417 (N_5417,N_911,N_877);
nand U5418 (N_5418,N_1110,N_2322);
xnor U5419 (N_5419,N_2144,N_1303);
nand U5420 (N_5420,N_4349,N_2245);
or U5421 (N_5421,N_3691,N_2148);
nor U5422 (N_5422,N_1079,N_2622);
nor U5423 (N_5423,N_1548,N_2049);
nand U5424 (N_5424,N_2154,N_4445);
and U5425 (N_5425,N_2494,N_2344);
and U5426 (N_5426,N_3606,N_527);
nand U5427 (N_5427,N_2897,N_1607);
and U5428 (N_5428,N_1139,N_4253);
or U5429 (N_5429,N_3720,N_2731);
xor U5430 (N_5430,N_2211,N_4636);
and U5431 (N_5431,N_3621,N_4680);
nor U5432 (N_5432,N_4481,N_4462);
xnor U5433 (N_5433,N_655,N_2966);
xnor U5434 (N_5434,N_2643,N_1134);
and U5435 (N_5435,N_4169,N_2246);
nand U5436 (N_5436,N_3446,N_4431);
or U5437 (N_5437,N_1559,N_3645);
nand U5438 (N_5438,N_1023,N_4418);
nand U5439 (N_5439,N_1994,N_3981);
nor U5440 (N_5440,N_1531,N_346);
nor U5441 (N_5441,N_4056,N_4384);
nand U5442 (N_5442,N_3038,N_4921);
and U5443 (N_5443,N_3670,N_1596);
xor U5444 (N_5444,N_1753,N_1865);
or U5445 (N_5445,N_3533,N_4003);
nor U5446 (N_5446,N_2469,N_1619);
and U5447 (N_5447,N_4116,N_4450);
and U5448 (N_5448,N_2356,N_2780);
or U5449 (N_5449,N_1080,N_2595);
xor U5450 (N_5450,N_4927,N_145);
nor U5451 (N_5451,N_4014,N_964);
nor U5452 (N_5452,N_259,N_243);
and U5453 (N_5453,N_3624,N_2936);
or U5454 (N_5454,N_2480,N_926);
or U5455 (N_5455,N_1001,N_3065);
nand U5456 (N_5456,N_1691,N_3045);
nor U5457 (N_5457,N_1766,N_2039);
xor U5458 (N_5458,N_3436,N_1241);
and U5459 (N_5459,N_2929,N_101);
nor U5460 (N_5460,N_4458,N_3084);
nand U5461 (N_5461,N_386,N_2281);
or U5462 (N_5462,N_1537,N_4389);
xnor U5463 (N_5463,N_4944,N_2464);
or U5464 (N_5464,N_2193,N_4683);
and U5465 (N_5465,N_788,N_1947);
xor U5466 (N_5466,N_4700,N_2965);
xor U5467 (N_5467,N_1372,N_4123);
xor U5468 (N_5468,N_4888,N_2543);
nand U5469 (N_5469,N_1316,N_2463);
nor U5470 (N_5470,N_4410,N_4027);
xor U5471 (N_5471,N_3499,N_3555);
xnor U5472 (N_5472,N_2773,N_3542);
or U5473 (N_5473,N_908,N_3368);
nand U5474 (N_5474,N_2902,N_3101);
nand U5475 (N_5475,N_2947,N_1155);
xor U5476 (N_5476,N_2121,N_1337);
or U5477 (N_5477,N_3032,N_2179);
or U5478 (N_5478,N_3128,N_85);
nand U5479 (N_5479,N_1715,N_1877);
xor U5480 (N_5480,N_3464,N_3132);
or U5481 (N_5481,N_134,N_2627);
and U5482 (N_5482,N_4489,N_3318);
nor U5483 (N_5483,N_2857,N_4074);
and U5484 (N_5484,N_4761,N_1471);
nand U5485 (N_5485,N_540,N_1352);
nand U5486 (N_5486,N_4814,N_1844);
xor U5487 (N_5487,N_1529,N_489);
xnor U5488 (N_5488,N_1249,N_1652);
nand U5489 (N_5489,N_1688,N_4221);
or U5490 (N_5490,N_23,N_242);
and U5491 (N_5491,N_803,N_1245);
nand U5492 (N_5492,N_4434,N_1100);
xnor U5493 (N_5493,N_834,N_3397);
and U5494 (N_5494,N_1466,N_2268);
nor U5495 (N_5495,N_3147,N_2411);
or U5496 (N_5496,N_241,N_2581);
nand U5497 (N_5497,N_206,N_1257);
nand U5498 (N_5498,N_3989,N_2112);
or U5499 (N_5499,N_2499,N_2745);
xor U5500 (N_5500,N_4541,N_2131);
nor U5501 (N_5501,N_483,N_194);
and U5502 (N_5502,N_3944,N_4720);
or U5503 (N_5503,N_3241,N_4124);
and U5504 (N_5504,N_3595,N_4185);
xnor U5505 (N_5505,N_4087,N_1982);
xnor U5506 (N_5506,N_2690,N_2014);
or U5507 (N_5507,N_4088,N_476);
or U5508 (N_5508,N_3906,N_1578);
nor U5509 (N_5509,N_2424,N_2311);
nand U5510 (N_5510,N_2359,N_3457);
or U5511 (N_5511,N_2296,N_2209);
nand U5512 (N_5512,N_3809,N_3751);
or U5513 (N_5513,N_1223,N_2860);
or U5514 (N_5514,N_2284,N_2762);
xnor U5515 (N_5515,N_3651,N_1312);
or U5516 (N_5516,N_2397,N_4607);
xnor U5517 (N_5517,N_2318,N_1870);
xnor U5518 (N_5518,N_526,N_3827);
and U5519 (N_5519,N_4887,N_953);
xor U5520 (N_5520,N_2430,N_589);
nor U5521 (N_5521,N_4859,N_4338);
or U5522 (N_5522,N_4143,N_3202);
or U5523 (N_5523,N_2735,N_1732);
nor U5524 (N_5524,N_2645,N_533);
nand U5525 (N_5525,N_1987,N_4515);
or U5526 (N_5526,N_146,N_1611);
nand U5527 (N_5527,N_3648,N_1055);
nor U5528 (N_5528,N_3422,N_2930);
or U5529 (N_5529,N_1931,N_2585);
nor U5530 (N_5530,N_54,N_2348);
xnor U5531 (N_5531,N_295,N_2748);
xnor U5532 (N_5532,N_4999,N_3790);
nor U5533 (N_5533,N_808,N_4133);
or U5534 (N_5534,N_2850,N_3025);
and U5535 (N_5535,N_2455,N_3559);
nand U5536 (N_5536,N_3544,N_4080);
nor U5537 (N_5537,N_4702,N_3712);
nor U5538 (N_5538,N_4939,N_850);
nor U5539 (N_5539,N_2504,N_329);
or U5540 (N_5540,N_475,N_1132);
or U5541 (N_5541,N_171,N_4423);
and U5542 (N_5542,N_615,N_4223);
nand U5543 (N_5543,N_2323,N_1685);
nor U5544 (N_5544,N_2299,N_1776);
or U5545 (N_5545,N_2350,N_1107);
xor U5546 (N_5546,N_1073,N_3063);
and U5547 (N_5547,N_3120,N_1698);
and U5548 (N_5548,N_813,N_1597);
nand U5549 (N_5549,N_985,N_3331);
nor U5550 (N_5550,N_1008,N_1665);
nor U5551 (N_5551,N_3134,N_4628);
xor U5552 (N_5552,N_2058,N_2698);
nor U5553 (N_5553,N_1116,N_3111);
and U5554 (N_5554,N_156,N_2855);
and U5555 (N_5555,N_1787,N_3267);
nand U5556 (N_5556,N_4586,N_2325);
or U5557 (N_5557,N_4545,N_420);
nor U5558 (N_5558,N_1566,N_4686);
and U5559 (N_5559,N_1018,N_4245);
nand U5560 (N_5560,N_3349,N_4084);
and U5561 (N_5561,N_4930,N_2995);
or U5562 (N_5562,N_3371,N_1327);
xnor U5563 (N_5563,N_4739,N_3865);
xor U5564 (N_5564,N_424,N_1233);
xnor U5565 (N_5565,N_1017,N_695);
xor U5566 (N_5566,N_327,N_3962);
and U5567 (N_5567,N_3873,N_2967);
or U5568 (N_5568,N_1348,N_3667);
nor U5569 (N_5569,N_3508,N_354);
nor U5570 (N_5570,N_1420,N_967);
and U5571 (N_5571,N_148,N_4664);
or U5572 (N_5572,N_2102,N_1511);
nand U5573 (N_5573,N_3106,N_2549);
xnor U5574 (N_5574,N_1985,N_1156);
or U5575 (N_5575,N_1843,N_4503);
nor U5576 (N_5576,N_4870,N_3889);
nand U5577 (N_5577,N_336,N_1711);
and U5578 (N_5578,N_4774,N_71);
and U5579 (N_5579,N_3860,N_272);
nor U5580 (N_5580,N_1409,N_421);
nand U5581 (N_5581,N_4551,N_1645);
nor U5582 (N_5582,N_2852,N_3016);
nand U5583 (N_5583,N_2577,N_375);
nand U5584 (N_5584,N_1433,N_262);
or U5585 (N_5585,N_4705,N_2994);
or U5586 (N_5586,N_254,N_4937);
nor U5587 (N_5587,N_3332,N_381);
xnor U5588 (N_5588,N_1175,N_556);
or U5589 (N_5589,N_4500,N_1703);
nand U5590 (N_5590,N_4283,N_4009);
xor U5591 (N_5591,N_163,N_4658);
xor U5592 (N_5592,N_1514,N_3787);
and U5593 (N_5593,N_4687,N_3488);
and U5594 (N_5594,N_2910,N_3678);
nor U5595 (N_5595,N_2321,N_4314);
or U5596 (N_5596,N_3192,N_3522);
nor U5597 (N_5597,N_4976,N_4611);
nor U5598 (N_5598,N_4217,N_4588);
nor U5599 (N_5599,N_4854,N_4359);
nand U5600 (N_5600,N_3759,N_882);
nand U5601 (N_5601,N_1746,N_1587);
nand U5602 (N_5602,N_495,N_181);
nand U5603 (N_5603,N_592,N_3414);
or U5604 (N_5604,N_4961,N_1369);
xor U5605 (N_5605,N_4091,N_3804);
or U5606 (N_5606,N_1562,N_4600);
nand U5607 (N_5607,N_248,N_2412);
xnor U5608 (N_5608,N_648,N_960);
and U5609 (N_5609,N_3339,N_3394);
nand U5610 (N_5610,N_4988,N_1148);
xnor U5611 (N_5611,N_3761,N_4916);
nand U5612 (N_5612,N_4255,N_2489);
xor U5613 (N_5613,N_2882,N_3709);
nand U5614 (N_5614,N_3949,N_1999);
nand U5615 (N_5615,N_3036,N_567);
xnor U5616 (N_5616,N_2887,N_3971);
nand U5617 (N_5617,N_314,N_469);
or U5618 (N_5618,N_3572,N_1499);
and U5619 (N_5619,N_3849,N_2044);
nand U5620 (N_5620,N_2224,N_3538);
nand U5621 (N_5621,N_1335,N_4216);
nor U5622 (N_5622,N_2445,N_1131);
and U5623 (N_5623,N_2393,N_2895);
xor U5624 (N_5624,N_2085,N_880);
xnor U5625 (N_5625,N_2351,N_3882);
and U5626 (N_5626,N_3105,N_1176);
or U5627 (N_5627,N_1580,N_3291);
xor U5628 (N_5628,N_2517,N_894);
xor U5629 (N_5629,N_1811,N_4422);
nor U5630 (N_5630,N_2779,N_4706);
and U5631 (N_5631,N_2016,N_4791);
nand U5632 (N_5632,N_1641,N_500);
nor U5633 (N_5633,N_1183,N_493);
xor U5634 (N_5634,N_250,N_3954);
nand U5635 (N_5635,N_3829,N_2370);
or U5636 (N_5636,N_3704,N_523);
nand U5637 (N_5637,N_3915,N_3736);
nand U5638 (N_5638,N_2675,N_3468);
nor U5639 (N_5639,N_1616,N_3190);
xnor U5640 (N_5640,N_1085,N_1261);
xnor U5641 (N_5641,N_1842,N_2650);
nor U5642 (N_5642,N_2928,N_659);
nand U5643 (N_5643,N_3654,N_4764);
nand U5644 (N_5644,N_1806,N_1624);
xnor U5645 (N_5645,N_1628,N_4521);
nand U5646 (N_5646,N_1457,N_980);
or U5647 (N_5647,N_1047,N_1203);
xnor U5648 (N_5648,N_2070,N_562);
xnor U5649 (N_5649,N_4052,N_4492);
nor U5650 (N_5650,N_4097,N_3671);
xnor U5651 (N_5651,N_186,N_1522);
or U5652 (N_5652,N_2417,N_76);
nor U5653 (N_5653,N_2767,N_1308);
xnor U5654 (N_5654,N_2242,N_3838);
nor U5655 (N_5655,N_2041,N_4971);
or U5656 (N_5656,N_3239,N_3085);
or U5657 (N_5657,N_4161,N_2803);
and U5658 (N_5658,N_3428,N_4034);
xor U5659 (N_5659,N_1883,N_1092);
and U5660 (N_5660,N_3911,N_4442);
or U5661 (N_5661,N_4452,N_3327);
and U5662 (N_5662,N_4387,N_2665);
nand U5663 (N_5663,N_733,N_959);
nand U5664 (N_5664,N_4180,N_1400);
nor U5665 (N_5665,N_3229,N_4815);
xnor U5666 (N_5666,N_1748,N_2324);
and U5667 (N_5667,N_2403,N_3502);
or U5668 (N_5668,N_4953,N_1356);
nand U5669 (N_5669,N_1498,N_2769);
and U5670 (N_5670,N_4873,N_2099);
and U5671 (N_5671,N_3387,N_3119);
nor U5672 (N_5672,N_2619,N_833);
and U5673 (N_5673,N_3300,N_2956);
nor U5674 (N_5674,N_809,N_751);
nor U5675 (N_5675,N_3276,N_3695);
xnor U5676 (N_5676,N_918,N_1654);
xor U5677 (N_5677,N_4012,N_2958);
nand U5678 (N_5678,N_734,N_4238);
nand U5679 (N_5679,N_1007,N_1363);
and U5680 (N_5680,N_2317,N_3340);
and U5681 (N_5681,N_3415,N_3723);
and U5682 (N_5682,N_2582,N_1486);
or U5683 (N_5683,N_4850,N_4635);
xor U5684 (N_5684,N_2186,N_3864);
xnor U5685 (N_5685,N_2617,N_2301);
and U5686 (N_5686,N_4329,N_481);
nor U5687 (N_5687,N_2082,N_1041);
or U5688 (N_5688,N_4081,N_991);
nand U5689 (N_5689,N_2497,N_2919);
xor U5690 (N_5690,N_3638,N_3256);
or U5691 (N_5691,N_674,N_2705);
or U5692 (N_5692,N_969,N_161);
xor U5693 (N_5693,N_137,N_3474);
nand U5694 (N_5694,N_64,N_4797);
nand U5695 (N_5695,N_4965,N_3600);
and U5696 (N_5696,N_1282,N_3910);
or U5697 (N_5697,N_667,N_3224);
and U5698 (N_5698,N_1128,N_470);
or U5699 (N_5699,N_4995,N_3328);
or U5700 (N_5700,N_2053,N_1117);
and U5701 (N_5701,N_1867,N_1309);
and U5702 (N_5702,N_2800,N_1997);
nor U5703 (N_5703,N_4397,N_3023);
nor U5704 (N_5704,N_1943,N_4237);
and U5705 (N_5705,N_4612,N_3296);
xor U5706 (N_5706,N_2388,N_292);
xor U5707 (N_5707,N_4563,N_3099);
xnor U5708 (N_5708,N_4578,N_2615);
nand U5709 (N_5709,N_2993,N_4355);
nor U5710 (N_5710,N_697,N_1199);
nor U5711 (N_5711,N_3630,N_1874);
and U5712 (N_5712,N_2511,N_3706);
xor U5713 (N_5713,N_4137,N_2452);
nor U5714 (N_5714,N_1975,N_2835);
nand U5715 (N_5715,N_4032,N_2239);
nor U5716 (N_5716,N_2583,N_3520);
and U5717 (N_5717,N_1791,N_198);
or U5718 (N_5718,N_8,N_2878);
nor U5719 (N_5719,N_3943,N_3322);
nand U5720 (N_5720,N_325,N_4250);
xnor U5721 (N_5721,N_393,N_4381);
xnor U5722 (N_5722,N_450,N_913);
nor U5723 (N_5723,N_223,N_1151);
xnor U5724 (N_5724,N_2374,N_3721);
or U5725 (N_5725,N_2957,N_3672);
and U5726 (N_5726,N_501,N_397);
xnor U5727 (N_5727,N_1315,N_2920);
xor U5728 (N_5728,N_2414,N_543);
xnor U5729 (N_5729,N_33,N_3348);
nor U5730 (N_5730,N_2747,N_3398);
or U5731 (N_5731,N_4787,N_4145);
nand U5732 (N_5732,N_1953,N_811);
xor U5733 (N_5733,N_986,N_1247);
nand U5734 (N_5734,N_162,N_744);
xnor U5735 (N_5735,N_3489,N_474);
and U5736 (N_5736,N_585,N_2334);
nand U5737 (N_5737,N_4825,N_321);
or U5738 (N_5738,N_3263,N_1334);
or U5739 (N_5739,N_1602,N_771);
and U5740 (N_5740,N_97,N_4662);
nand U5741 (N_5741,N_4610,N_2149);
xnor U5742 (N_5742,N_660,N_3077);
and U5743 (N_5743,N_966,N_359);
nor U5744 (N_5744,N_951,N_94);
or U5745 (N_5745,N_2253,N_3246);
xnor U5746 (N_5746,N_3696,N_4827);
xnor U5747 (N_5747,N_792,N_2552);
nor U5748 (N_5748,N_1563,N_3247);
xor U5749 (N_5749,N_2962,N_4510);
and U5750 (N_5750,N_2990,N_3427);
and U5751 (N_5751,N_1415,N_3257);
and U5752 (N_5752,N_535,N_215);
and U5753 (N_5753,N_4777,N_1157);
or U5754 (N_5754,N_138,N_2737);
and U5755 (N_5755,N_4215,N_2498);
xor U5756 (N_5756,N_3615,N_4499);
nor U5757 (N_5757,N_2177,N_4451);
and U5758 (N_5758,N_3124,N_2522);
nand U5759 (N_5759,N_4028,N_2091);
nor U5760 (N_5760,N_3846,N_1496);
or U5761 (N_5761,N_4839,N_4150);
and U5762 (N_5762,N_3716,N_1364);
xnor U5763 (N_5763,N_758,N_637);
and U5764 (N_5764,N_4309,N_2604);
nor U5765 (N_5765,N_1109,N_2553);
nor U5766 (N_5766,N_561,N_4760);
nand U5767 (N_5767,N_342,N_4045);
and U5768 (N_5768,N_4419,N_1392);
nand U5769 (N_5769,N_3178,N_4296);
xnor U5770 (N_5770,N_4230,N_3378);
nand U5771 (N_5771,N_3616,N_3530);
or U5772 (N_5772,N_2539,N_3424);
nor U5773 (N_5773,N_2834,N_3123);
nand U5774 (N_5774,N_3027,N_1338);
xor U5775 (N_5775,N_853,N_1976);
and U5776 (N_5776,N_4471,N_2787);
and U5777 (N_5777,N_2853,N_1220);
xor U5778 (N_5778,N_20,N_2176);
nand U5779 (N_5779,N_3311,N_4848);
or U5780 (N_5780,N_2861,N_3021);
or U5781 (N_5781,N_4638,N_289);
nor U5782 (N_5782,N_1384,N_2173);
nand U5783 (N_5783,N_4290,N_3983);
nand U5784 (N_5784,N_4368,N_3218);
or U5785 (N_5785,N_2263,N_2598);
or U5786 (N_5786,N_2568,N_3744);
and U5787 (N_5787,N_3554,N_3108);
and U5788 (N_5788,N_340,N_1873);
and U5789 (N_5789,N_797,N_1009);
nor U5790 (N_5790,N_816,N_2341);
nand U5791 (N_5791,N_1136,N_4738);
or U5792 (N_5792,N_437,N_4544);
xnor U5793 (N_5793,N_1273,N_2901);
nand U5794 (N_5794,N_3702,N_2110);
and U5795 (N_5795,N_4609,N_4762);
nor U5796 (N_5796,N_3399,N_3747);
nand U5797 (N_5797,N_1229,N_1640);
xor U5798 (N_5798,N_4757,N_4249);
and U5799 (N_5799,N_3566,N_3380);
or U5800 (N_5800,N_2883,N_639);
or U5801 (N_5801,N_2843,N_3614);
or U5802 (N_5802,N_3794,N_4631);
and U5803 (N_5803,N_1095,N_3164);
and U5804 (N_5804,N_1304,N_2188);
nand U5805 (N_5805,N_4792,N_2614);
xnor U5806 (N_5806,N_4574,N_4435);
and U5807 (N_5807,N_1495,N_3807);
xor U5808 (N_5808,N_2978,N_1786);
nand U5809 (N_5809,N_2593,N_840);
and U5810 (N_5810,N_949,N_2875);
and U5811 (N_5811,N_1320,N_680);
xnor U5812 (N_5812,N_2095,N_832);
and U5813 (N_5813,N_2163,N_2566);
xnor U5814 (N_5814,N_4872,N_729);
nand U5815 (N_5815,N_623,N_4518);
and U5816 (N_5816,N_3798,N_3381);
and U5817 (N_5817,N_4304,N_1621);
nor U5818 (N_5818,N_3552,N_4591);
and U5819 (N_5819,N_2912,N_96);
xnor U5820 (N_5820,N_4403,N_2431);
xnor U5821 (N_5821,N_4409,N_4204);
nand U5822 (N_5822,N_1345,N_1423);
and U5823 (N_5823,N_672,N_2446);
xnor U5824 (N_5824,N_1179,N_2603);
or U5825 (N_5825,N_3799,N_544);
or U5826 (N_5826,N_3673,N_3002);
nand U5827 (N_5827,N_2573,N_63);
or U5828 (N_5828,N_1195,N_3367);
xnor U5829 (N_5829,N_4197,N_4062);
or U5830 (N_5830,N_4079,N_1460);
or U5831 (N_5831,N_1218,N_4548);
nor U5832 (N_5832,N_4914,N_1803);
xor U5833 (N_5833,N_3057,N_2338);
and U5834 (N_5834,N_4948,N_4293);
nor U5835 (N_5835,N_3626,N_4516);
nor U5836 (N_5836,N_1251,N_794);
or U5837 (N_5837,N_1407,N_1713);
xor U5838 (N_5838,N_2283,N_157);
nand U5839 (N_5839,N_745,N_2666);
nand U5840 (N_5840,N_3472,N_3198);
nor U5841 (N_5841,N_3551,N_4385);
or U5842 (N_5842,N_160,N_925);
and U5843 (N_5843,N_4260,N_2168);
nor U5844 (N_5844,N_661,N_1759);
or U5845 (N_5845,N_763,N_3726);
or U5846 (N_5846,N_4661,N_3466);
nand U5847 (N_5847,N_3770,N_4302);
or U5848 (N_5848,N_2034,N_2275);
nor U5849 (N_5849,N_1191,N_378);
nand U5850 (N_5850,N_4191,N_4831);
nand U5851 (N_5851,N_260,N_3880);
and U5852 (N_5852,N_541,N_3919);
xor U5853 (N_5853,N_4526,N_4822);
and U5854 (N_5854,N_1673,N_4505);
or U5855 (N_5855,N_4579,N_140);
or U5856 (N_5856,N_551,N_1299);
nand U5857 (N_5857,N_3393,N_2954);
or U5858 (N_5858,N_4783,N_881);
nor U5859 (N_5859,N_4077,N_398);
xor U5860 (N_5860,N_973,N_1482);
and U5861 (N_5861,N_1917,N_317);
nand U5862 (N_5862,N_724,N_1070);
xor U5863 (N_5863,N_4520,N_3642);
and U5864 (N_5864,N_2785,N_4393);
or U5865 (N_5865,N_4694,N_310);
nor U5866 (N_5866,N_2542,N_4182);
or U5867 (N_5867,N_4590,N_4649);
nor U5868 (N_5868,N_2988,N_2109);
or U5869 (N_5869,N_4596,N_35);
nand U5870 (N_5870,N_125,N_3156);
nand U5871 (N_5871,N_4793,N_3548);
xnor U5872 (N_5872,N_4334,N_4132);
nand U5873 (N_5873,N_377,N_4396);
or U5874 (N_5874,N_436,N_581);
or U5875 (N_5875,N_4429,N_738);
xor U5876 (N_5876,N_2806,N_1474);
or U5877 (N_5877,N_936,N_1063);
and U5878 (N_5878,N_462,N_2229);
and U5879 (N_5879,N_3418,N_3984);
xnor U5880 (N_5880,N_767,N_3580);
nand U5881 (N_5881,N_3968,N_681);
nor U5882 (N_5882,N_3701,N_3594);
nand U5883 (N_5883,N_4094,N_2409);
or U5884 (N_5884,N_4905,N_3518);
nand U5885 (N_5885,N_4907,N_690);
nor U5886 (N_5886,N_4593,N_3531);
xor U5887 (N_5887,N_3495,N_4834);
and U5888 (N_5888,N_200,N_4682);
xor U5889 (N_5889,N_1287,N_3728);
nand U5890 (N_5890,N_706,N_1924);
and U5891 (N_5891,N_2530,N_4731);
nand U5892 (N_5892,N_456,N_1509);
and U5893 (N_5893,N_1764,N_1771);
nor U5894 (N_5894,N_4583,N_4629);
nor U5895 (N_5895,N_2924,N_3760);
nand U5896 (N_5896,N_2845,N_3234);
xor U5897 (N_5897,N_4343,N_1298);
and U5898 (N_5898,N_4374,N_135);
nor U5899 (N_5899,N_2231,N_4112);
or U5900 (N_5900,N_1797,N_822);
nand U5901 (N_5901,N_296,N_3017);
nor U5902 (N_5902,N_3683,N_3301);
xnor U5903 (N_5903,N_2415,N_2678);
or U5904 (N_5904,N_4806,N_3416);
nor U5905 (N_5905,N_2485,N_3376);
nor U5906 (N_5906,N_2288,N_820);
xor U5907 (N_5907,N_4817,N_1248);
nor U5908 (N_5908,N_4188,N_439);
xnor U5909 (N_5909,N_487,N_1840);
or U5910 (N_5910,N_1333,N_3344);
nor U5911 (N_5911,N_546,N_2802);
and U5912 (N_5912,N_3754,N_1808);
nor U5913 (N_5913,N_4200,N_3986);
nor U5914 (N_5914,N_3306,N_263);
xnor U5915 (N_5915,N_4744,N_2739);
nor U5916 (N_5916,N_3133,N_3800);
xnor U5917 (N_5917,N_2451,N_588);
xnor U5918 (N_5918,N_1667,N_4816);
nor U5919 (N_5919,N_4350,N_2001);
nor U5920 (N_5920,N_2732,N_2031);
or U5921 (N_5921,N_2563,N_4996);
or U5922 (N_5922,N_3752,N_1154);
or U5923 (N_5923,N_1456,N_2858);
or U5924 (N_5924,N_2817,N_405);
nand U5925 (N_5925,N_4153,N_1986);
nor U5926 (N_5926,N_3127,N_1648);
or U5927 (N_5927,N_1093,N_1984);
nand U5928 (N_5928,N_1722,N_3307);
or U5929 (N_5929,N_779,N_2814);
nand U5930 (N_5930,N_3092,N_1037);
nand U5931 (N_5931,N_4826,N_4243);
nor U5932 (N_5932,N_2221,N_1065);
nor U5933 (N_5933,N_1847,N_128);
xnor U5934 (N_5934,N_539,N_4871);
or U5935 (N_5935,N_2807,N_4159);
xor U5936 (N_5936,N_4327,N_3005);
and U5937 (N_5937,N_998,N_4240);
xor U5938 (N_5938,N_371,N_2886);
nand U5939 (N_5939,N_1573,N_4022);
or U5940 (N_5940,N_2505,N_3627);
or U5941 (N_5941,N_3724,N_3762);
nor U5942 (N_5942,N_4924,N_416);
nor U5943 (N_5943,N_297,N_1649);
nand U5944 (N_5944,N_3894,N_4877);
nor U5945 (N_5945,N_4051,N_2071);
xnor U5946 (N_5946,N_3697,N_3513);
and U5947 (N_5947,N_2395,N_2885);
and U5948 (N_5948,N_2601,N_891);
xor U5949 (N_5949,N_1916,N_511);
xor U5950 (N_5950,N_2482,N_2975);
or U5951 (N_5951,N_935,N_471);
and U5952 (N_5952,N_1422,N_3022);
nand U5953 (N_5953,N_2697,N_1650);
or U5954 (N_5954,N_1057,N_4258);
nor U5955 (N_5955,N_4633,N_428);
or U5956 (N_5956,N_2478,N_1021);
and U5957 (N_5957,N_2220,N_4470);
xor U5958 (N_5958,N_3610,N_1869);
and U5959 (N_5959,N_3975,N_4966);
or U5960 (N_5960,N_1491,N_805);
nor U5961 (N_5961,N_2942,N_1693);
and U5962 (N_5962,N_506,N_707);
or U5963 (N_5963,N_574,N_944);
nor U5964 (N_5964,N_1192,N_2695);
and U5965 (N_5965,N_1885,N_2600);
nor U5966 (N_5966,N_4869,N_1505);
nor U5967 (N_5967,N_3961,N_3605);
or U5968 (N_5968,N_1494,N_4351);
or U5969 (N_5969,N_3938,N_2792);
and U5970 (N_5970,N_4979,N_664);
xor U5971 (N_5971,N_2662,N_3966);
nand U5972 (N_5972,N_4402,N_2945);
nor U5973 (N_5973,N_3977,N_2564);
nor U5974 (N_5974,N_4865,N_1492);
nand U5975 (N_5975,N_896,N_2073);
nand U5976 (N_5976,N_1528,N_1427);
nand U5977 (N_5977,N_4212,N_898);
nand U5978 (N_5978,N_825,N_2022);
xnor U5979 (N_5979,N_2713,N_4242);
xor U5980 (N_5980,N_4324,N_3135);
nand U5981 (N_5981,N_2045,N_704);
and U5982 (N_5982,N_4174,N_3191);
or U5983 (N_5983,N_1142,N_1146);
nand U5984 (N_5984,N_2825,N_400);
and U5985 (N_5985,N_2893,N_2933);
xor U5986 (N_5986,N_3774,N_1052);
nor U5987 (N_5987,N_1577,N_2143);
or U5988 (N_5988,N_302,N_2523);
nor U5989 (N_5989,N_2258,N_2155);
nand U5990 (N_5990,N_2556,N_4670);
or U5991 (N_5991,N_2426,N_1871);
and U5992 (N_5992,N_3013,N_395);
or U5993 (N_5993,N_4168,N_852);
nor U5994 (N_5994,N_3856,N_404);
nand U5995 (N_5995,N_1668,N_2743);
xnor U5996 (N_5996,N_2774,N_4582);
nand U5997 (N_5997,N_1516,N_3260);
nor U5998 (N_5998,N_987,N_3549);
or U5999 (N_5999,N_4987,N_3965);
or U6000 (N_6000,N_3396,N_2259);
or U6001 (N_6001,N_370,N_2398);
and U6002 (N_6002,N_2703,N_3130);
and U6003 (N_6003,N_2219,N_3738);
nor U6004 (N_6004,N_4122,N_2863);
or U6005 (N_6005,N_1926,N_4986);
xor U6006 (N_6006,N_4514,N_1535);
xor U6007 (N_6007,N_3767,N_4007);
and U6008 (N_6008,N_3125,N_3563);
or U6009 (N_6009,N_121,N_4685);
xor U6010 (N_6010,N_2391,N_1056);
nor U6011 (N_6011,N_652,N_4799);
xnor U6012 (N_6012,N_4156,N_4157);
nand U6013 (N_6013,N_452,N_3801);
and U6014 (N_6014,N_1690,N_4560);
nor U6015 (N_6015,N_1613,N_4721);
xnor U6016 (N_6016,N_2776,N_4820);
and U6017 (N_6017,N_3693,N_1913);
nand U6018 (N_6018,N_4428,N_742);
xnor U6019 (N_6019,N_1378,N_1684);
nor U6020 (N_6020,N_3578,N_1710);
and U6021 (N_6021,N_281,N_3604);
nor U6022 (N_6022,N_1326,N_3888);
and U6023 (N_6023,N_4140,N_423);
xor U6024 (N_6024,N_2265,N_3854);
nand U6025 (N_6025,N_2162,N_683);
or U6026 (N_6026,N_2013,N_2438);
nor U6027 (N_6027,N_2710,N_4038);
or U6028 (N_6028,N_339,N_1446);
and U6029 (N_6029,N_2382,N_105);
xor U6030 (N_6030,N_2881,N_1872);
nand U6031 (N_6031,N_2744,N_3281);
xor U6032 (N_6032,N_3635,N_3206);
nand U6033 (N_6033,N_4251,N_2420);
or U6034 (N_6034,N_597,N_3803);
xnor U6035 (N_6035,N_4322,N_2346);
nand U6036 (N_6036,N_2856,N_2740);
nor U6037 (N_6037,N_3641,N_861);
or U6038 (N_6038,N_3404,N_570);
and U6039 (N_6039,N_905,N_1523);
xor U6040 (N_6040,N_4372,N_940);
xnor U6041 (N_6041,N_4142,N_2383);
or U6042 (N_6042,N_4964,N_1098);
xor U6043 (N_6043,N_3802,N_4798);
nand U6044 (N_6044,N_2632,N_3874);
or U6045 (N_6045,N_499,N_1908);
xor U6046 (N_6046,N_1781,N_362);
or U6047 (N_6047,N_172,N_1360);
nor U6048 (N_6048,N_401,N_1246);
and U6049 (N_6049,N_1225,N_1507);
or U6050 (N_6050,N_2319,N_1839);
or U6051 (N_6051,N_2037,N_2508);
nand U6052 (N_6052,N_4749,N_1387);
xnor U6053 (N_6053,N_4862,N_3003);
or U6054 (N_6054,N_802,N_2475);
nand U6055 (N_6055,N_1089,N_2226);
xnor U6056 (N_6056,N_601,N_1359);
or U6057 (N_6057,N_4490,N_4151);
nor U6058 (N_6058,N_298,N_3413);
nor U6059 (N_6059,N_2907,N_3060);
xor U6060 (N_6060,N_1027,N_364);
and U6061 (N_6061,N_2869,N_2347);
and U6062 (N_6062,N_3121,N_4053);
and U6063 (N_6063,N_3755,N_774);
or U6064 (N_6064,N_1476,N_3066);
or U6065 (N_6065,N_4575,N_4277);
nor U6066 (N_6066,N_920,N_3313);
nor U6067 (N_6067,N_4042,N_3951);
nand U6068 (N_6068,N_2976,N_4121);
nor U6069 (N_6069,N_3902,N_17);
and U6070 (N_6070,N_3942,N_3012);
and U6071 (N_6071,N_3150,N_3243);
xnor U6072 (N_6072,N_2,N_2064);
nand U6073 (N_6073,N_566,N_647);
xnor U6074 (N_6074,N_2946,N_629);
nand U6075 (N_6075,N_2914,N_3681);
and U6076 (N_6076,N_3851,N_2569);
and U6077 (N_6077,N_856,N_617);
xnor U6078 (N_6078,N_3715,N_83);
or U6079 (N_6079,N_4425,N_4106);
and U6080 (N_6080,N_142,N_15);
or U6081 (N_6081,N_517,N_1439);
nand U6082 (N_6082,N_3317,N_2527);
or U6083 (N_6083,N_1863,N_2891);
or U6084 (N_6084,N_484,N_1140);
and U6085 (N_6085,N_4824,N_1899);
nand U6086 (N_6086,N_2927,N_1174);
nor U6087 (N_6087,N_230,N_2590);
nand U6088 (N_6088,N_4994,N_3353);
nand U6089 (N_6089,N_1404,N_3785);
nand U6090 (N_6090,N_4303,N_748);
nor U6091 (N_6091,N_2888,N_3059);
and U6092 (N_6092,N_2700,N_3819);
and U6093 (N_6093,N_2725,N_4671);
and U6094 (N_6094,N_4892,N_4833);
xor U6095 (N_6095,N_2000,N_3325);
or U6096 (N_6096,N_686,N_399);
or U6097 (N_6097,N_512,N_777);
or U6098 (N_6098,N_3561,N_3237);
nand U6099 (N_6099,N_3825,N_465);
nor U6100 (N_6100,N_1637,N_3834);
nand U6101 (N_6101,N_1658,N_41);
nand U6102 (N_6102,N_1133,N_4725);
xor U6103 (N_6103,N_2333,N_387);
or U6104 (N_6104,N_996,N_709);
and U6105 (N_6105,N_4165,N_2846);
nor U6106 (N_6106,N_2272,N_306);
xnor U6107 (N_6107,N_2503,N_1171);
and U6108 (N_6108,N_1894,N_3835);
xor U6109 (N_6109,N_3292,N_2089);
nor U6110 (N_6110,N_4830,N_187);
xnor U6111 (N_6111,N_981,N_3596);
xor U6112 (N_6112,N_545,N_4525);
xor U6113 (N_6113,N_607,N_3591);
and U6114 (N_6114,N_1903,N_618);
and U6115 (N_6115,N_3297,N_3534);
nor U6116 (N_6116,N_245,N_2599);
nor U6117 (N_6117,N_1121,N_3342);
xor U6118 (N_6118,N_3249,N_2594);
nor U6119 (N_6119,N_2559,N_1291);
or U6120 (N_6120,N_2658,N_2741);
nor U6121 (N_6121,N_2092,N_3138);
and U6122 (N_6122,N_1664,N_1802);
xor U6123 (N_6123,N_721,N_2119);
xnor U6124 (N_6124,N_1465,N_4281);
nor U6125 (N_6125,N_907,N_1389);
nand U6126 (N_6126,N_2638,N_757);
nor U6127 (N_6127,N_4856,N_3308);
and U6128 (N_6128,N_2840,N_4406);
or U6129 (N_6129,N_4289,N_4972);
xnor U6130 (N_6130,N_1091,N_4718);
nor U6131 (N_6131,N_859,N_2160);
xnor U6132 (N_6132,N_1122,N_2360);
or U6133 (N_6133,N_2672,N_2490);
nor U6134 (N_6134,N_1600,N_3999);
or U6135 (N_6135,N_4020,N_962);
nand U6136 (N_6136,N_43,N_858);
xnor U6137 (N_6137,N_692,N_4102);
xnor U6138 (N_6138,N_4206,N_1910);
nor U6139 (N_6139,N_3046,N_1770);
and U6140 (N_6140,N_4152,N_4674);
xnor U6141 (N_6141,N_2751,N_488);
nor U6142 (N_6142,N_1838,N_2724);
nor U6143 (N_6143,N_2830,N_1709);
nor U6144 (N_6144,N_394,N_4675);
or U6145 (N_6145,N_1677,N_4517);
nand U6146 (N_6146,N_4073,N_4868);
and U6147 (N_6147,N_764,N_2547);
and U6148 (N_6148,N_1809,N_326);
or U6149 (N_6149,N_3258,N_2405);
nor U6150 (N_6150,N_4998,N_4846);
xor U6151 (N_6151,N_2165,N_2266);
nand U6152 (N_6152,N_3354,N_4208);
or U6153 (N_6153,N_1583,N_754);
and U6154 (N_6154,N_4940,N_69);
nor U6155 (N_6155,N_782,N_3568);
or U6156 (N_6156,N_4139,N_2580);
nor U6157 (N_6157,N_293,N_4684);
and U6158 (N_6158,N_2028,N_3453);
xnor U6159 (N_6159,N_3477,N_2561);
nand U6160 (N_6160,N_4394,N_1394);
nand U6161 (N_6161,N_2240,N_1681);
xnor U6162 (N_6162,N_775,N_90);
or U6163 (N_6163,N_1901,N_4533);
nand U6164 (N_6164,N_3895,N_2023);
nor U6165 (N_6165,N_341,N_688);
nor U6166 (N_6166,N_3343,N_1096);
xor U6167 (N_6167,N_1878,N_3400);
nand U6168 (N_6168,N_3351,N_1201);
or U6169 (N_6169,N_2093,N_2349);
xor U6170 (N_6170,N_3222,N_3197);
or U6171 (N_6171,N_2558,N_1589);
nor U6172 (N_6172,N_1949,N_524);
xor U6173 (N_6173,N_1267,N_1062);
nand U6174 (N_6174,N_3529,N_3609);
xnor U6175 (N_6175,N_1608,N_3305);
xor U6176 (N_6176,N_1517,N_1662);
or U6177 (N_6177,N_644,N_2811);
nor U6178 (N_6178,N_3756,N_3571);
nand U6179 (N_6179,N_2894,N_3955);
or U6180 (N_6180,N_2309,N_4413);
nor U6181 (N_6181,N_1857,N_979);
nor U6182 (N_6182,N_466,N_3153);
xnor U6183 (N_6183,N_904,N_843);
or U6184 (N_6184,N_1129,N_1835);
nor U6185 (N_6185,N_4513,N_927);
or U6186 (N_6186,N_3588,N_1102);
nand U6187 (N_6187,N_4362,N_1630);
nand U6188 (N_6188,N_1497,N_565);
nor U6189 (N_6189,N_1747,N_3402);
xor U6190 (N_6190,N_4875,N_2156);
or U6191 (N_6191,N_3377,N_2025);
nand U6192 (N_6192,N_4064,N_3618);
xnor U6193 (N_6193,N_4024,N_133);
nand U6194 (N_6194,N_841,N_274);
nor U6195 (N_6195,N_3294,N_3469);
and U6196 (N_6196,N_3497,N_4992);
or U6197 (N_6197,N_3872,N_4746);
xor U6198 (N_6198,N_1487,N_2444);
or U6199 (N_6199,N_84,N_2717);
or U6200 (N_6200,N_2003,N_3204);
nand U6201 (N_6201,N_1330,N_3973);
nor U6202 (N_6202,N_4033,N_2286);
nor U6203 (N_6203,N_3952,N_4193);
nor U6204 (N_6204,N_2688,N_4411);
nor U6205 (N_6205,N_1237,N_4285);
xor U6206 (N_6206,N_3141,N_3663);
nand U6207 (N_6207,N_3442,N_3898);
or U6208 (N_6208,N_3061,N_1669);
xor U6209 (N_6209,N_1350,N_1149);
and U6210 (N_6210,N_1981,N_608);
and U6211 (N_6211,N_4177,N_1087);
nor U6212 (N_6212,N_2989,N_407);
and U6213 (N_6213,N_714,N_3242);
nand U6214 (N_6214,N_1019,N_1324);
or U6215 (N_6215,N_2300,N_1274);
nor U6216 (N_6216,N_1767,N_2167);
or U6217 (N_6217,N_4187,N_2126);
nand U6218 (N_6218,N_4885,N_1388);
and U6219 (N_6219,N_4040,N_2487);
nand U6220 (N_6220,N_3315,N_4207);
or U6221 (N_6221,N_4960,N_978);
or U6222 (N_6222,N_4838,N_3496);
nand U6223 (N_6223,N_719,N_2106);
xor U6224 (N_6224,N_2079,N_2531);
or U6225 (N_6225,N_679,N_396);
and U6226 (N_6226,N_313,N_1605);
nor U6227 (N_6227,N_1905,N_636);
nand U6228 (N_6228,N_479,N_264);
and U6229 (N_6229,N_3634,N_3705);
nor U6230 (N_6230,N_4532,N_239);
nand U6231 (N_6231,N_2329,N_4496);
and U6232 (N_6232,N_1204,N_1228);
and U6233 (N_6233,N_2174,N_74);
or U6234 (N_6234,N_3073,N_3607);
nand U6235 (N_6235,N_4605,N_1461);
xor U6236 (N_6236,N_4580,N_1054);
nor U6237 (N_6237,N_30,N_1002);
nand U6238 (N_6238,N_4810,N_627);
xnor U6239 (N_6239,N_1629,N_1922);
nor U6240 (N_6240,N_4265,N_3324);
or U6241 (N_6241,N_658,N_4681);
or U6242 (N_6242,N_3826,N_4602);
nor U6243 (N_6243,N_1410,N_2982);
nor U6244 (N_6244,N_1582,N_2746);
nor U6245 (N_6245,N_2664,N_3365);
and U6246 (N_6246,N_99,N_1006);
nand U6247 (N_6247,N_3467,N_1553);
nor U6248 (N_6248,N_1745,N_1181);
nand U6249 (N_6249,N_1483,N_207);
or U6250 (N_6250,N_3924,N_1479);
nand U6251 (N_6251,N_2797,N_100);
nor U6252 (N_6252,N_1742,N_609);
or U6253 (N_6253,N_67,N_760);
or U6254 (N_6254,N_3172,N_159);
and U6255 (N_6255,N_409,N_2466);
nand U6256 (N_6256,N_2536,N_2616);
and U6257 (N_6257,N_4307,N_702);
or U6258 (N_6258,N_1846,N_72);
nand U6259 (N_6259,N_573,N_938);
nor U6260 (N_6260,N_3733,N_2934);
xnor U6261 (N_6261,N_3160,N_2951);
nand U6262 (N_6262,N_3171,N_3700);
nor U6263 (N_6263,N_4775,N_787);
and U6264 (N_6264,N_1468,N_4345);
nand U6265 (N_6265,N_1854,N_711);
and U6266 (N_6266,N_3139,N_1353);
and U6267 (N_6267,N_3816,N_578);
nand U6268 (N_6268,N_2540,N_1655);
nor U6269 (N_6269,N_2937,N_2429);
or U6270 (N_6270,N_2107,N_879);
and U6271 (N_6271,N_2871,N_2247);
nand U6272 (N_6272,N_366,N_3221);
nor U6273 (N_6273,N_3622,N_78);
nand U6274 (N_6274,N_3921,N_3259);
nand U6275 (N_6275,N_3450,N_4336);
nor U6276 (N_6276,N_2704,N_1269);
nor U6277 (N_6277,N_3982,N_12);
and U6278 (N_6278,N_4696,N_2122);
nor U6279 (N_6279,N_4247,N_3543);
and U6280 (N_6280,N_1515,N_4407);
nand U6281 (N_6281,N_2120,N_762);
or U6282 (N_6282,N_2376,N_2336);
or U6283 (N_6283,N_1882,N_2842);
nor U6284 (N_6284,N_265,N_4002);
xnor U6285 (N_6285,N_4181,N_2270);
xnor U6286 (N_6286,N_3131,N_4058);
nor U6287 (N_6287,N_1469,N_2801);
xor U6288 (N_6288,N_3284,N_4501);
nand U6289 (N_6289,N_612,N_3855);
nand U6290 (N_6290,N_4184,N_2534);
or U6291 (N_6291,N_3114,N_1609);
nand U6292 (N_6292,N_3570,N_2088);
xnor U6293 (N_6293,N_4421,N_2996);
and U6294 (N_6294,N_3335,N_1554);
xnor U6295 (N_6295,N_3379,N_945);
xor U6296 (N_6296,N_3532,N_817);
xnor U6297 (N_6297,N_4288,N_2456);
nand U6298 (N_6298,N_3753,N_221);
and U6299 (N_6299,N_2516,N_3528);
and U6300 (N_6300,N_4727,N_2551);
nand U6301 (N_6301,N_1374,N_2502);
or U6302 (N_6302,N_82,N_3766);
and U6303 (N_6303,N_1361,N_3086);
or U6304 (N_6304,N_2648,N_236);
nand U6305 (N_6305,N_532,N_1042);
nand U6306 (N_6306,N_1230,N_3852);
xor U6307 (N_6307,N_1805,N_2673);
xor U6308 (N_6308,N_1815,N_3219);
nor U6309 (N_6309,N_1289,N_2898);
nor U6310 (N_6310,N_2418,N_3611);
xnor U6311 (N_6311,N_4618,N_3963);
or U6312 (N_6312,N_3262,N_2613);
xnor U6313 (N_6313,N_1500,N_4530);
xnor U6314 (N_6314,N_3011,N_3226);
or U6315 (N_6315,N_4225,N_2823);
and U6316 (N_6316,N_776,N_1571);
xor U6317 (N_6317,N_2416,N_1283);
and U6318 (N_6318,N_3892,N_1108);
nor U6319 (N_6319,N_963,N_999);
and U6320 (N_6320,N_1810,N_183);
and U6321 (N_6321,N_946,N_1915);
or U6322 (N_6322,N_3602,N_4558);
nand U6323 (N_6323,N_4008,N_3154);
xor U6324 (N_6324,N_3930,N_255);
or U6325 (N_6325,N_1207,N_3163);
nand U6326 (N_6326,N_3228,N_3004);
nor U6327 (N_6327,N_4581,N_3830);
nor U6328 (N_6328,N_4264,N_2192);
nor U6329 (N_6329,N_3437,N_1617);
nand U6330 (N_6330,N_1567,N_671);
xnor U6331 (N_6331,N_1319,N_696);
xnor U6332 (N_6332,N_2750,N_177);
xnor U6333 (N_6333,N_3116,N_1260);
and U6334 (N_6334,N_3769,N_1814);
or U6335 (N_6335,N_2277,N_3048);
nand U6336 (N_6336,N_502,N_130);
and U6337 (N_6337,N_2010,N_3289);
xnor U6338 (N_6338,N_2261,N_1145);
or U6339 (N_6339,N_3088,N_28);
nand U6340 (N_6340,N_2849,N_3564);
nor U6341 (N_6341,N_2313,N_2521);
or U6342 (N_6342,N_4163,N_2986);
nor U6343 (N_6343,N_3558,N_1428);
nor U6344 (N_6344,N_3806,N_4342);
or U6345 (N_6345,N_595,N_167);
or U6346 (N_6346,N_2524,N_1076);
xor U6347 (N_6347,N_22,N_4599);
or U6348 (N_6348,N_4945,N_4722);
xnor U6349 (N_6349,N_1321,N_1111);
nand U6350 (N_6350,N_2859,N_2427);
or U6351 (N_6351,N_1720,N_2251);
xor U6352 (N_6352,N_4369,N_4453);
nand U6353 (N_6353,N_3516,N_1779);
xor U6354 (N_6354,N_1386,N_1719);
nand U6355 (N_6355,N_2212,N_283);
nand U6356 (N_6356,N_3511,N_2320);
nor U6357 (N_6357,N_2390,N_4771);
nor U6358 (N_6358,N_1401,N_4616);
nand U6359 (N_6359,N_4155,N_3679);
and U6360 (N_6360,N_1754,N_4055);
xor U6361 (N_6361,N_3248,N_1086);
or U6362 (N_6362,N_1973,N_3043);
nor U6363 (N_6363,N_622,N_4699);
nand U6364 (N_6364,N_1368,N_2117);
or U6365 (N_6365,N_914,N_3265);
xor U6366 (N_6366,N_1841,N_3735);
nand U6367 (N_6367,N_3665,N_947);
nor U6368 (N_6368,N_110,N_2784);
nor U6369 (N_6369,N_2926,N_2378);
or U6370 (N_6370,N_3009,N_1104);
xnor U6371 (N_6371,N_1012,N_2094);
xnor U6372 (N_6372,N_3805,N_3639);
nand U6373 (N_6373,N_376,N_4754);
xor U6374 (N_6374,N_4678,N_4922);
and U6375 (N_6375,N_152,N_4138);
nand U6376 (N_6376,N_1998,N_3444);
nor U6377 (N_6377,N_3866,N_4047);
and U6378 (N_6378,N_1480,N_528);
or U6379 (N_6379,N_1022,N_534);
nand U6380 (N_6380,N_3780,N_2439);
or U6381 (N_6381,N_2683,N_2063);
and U6382 (N_6382,N_2477,N_2371);
nor U6383 (N_6383,N_836,N_2059);
nor U6384 (N_6384,N_3360,N_4160);
and U6385 (N_6385,N_2074,N_3748);
or U6386 (N_6386,N_1761,N_2386);
xor U6387 (N_6387,N_2636,N_3587);
xnor U6388 (N_6388,N_2765,N_3525);
nand U6389 (N_6389,N_865,N_1644);
nor U6390 (N_6390,N_4935,N_587);
and U6391 (N_6391,N_1506,N_2214);
xor U6392 (N_6392,N_2608,N_330);
and U6393 (N_6393,N_2671,N_1383);
or U6394 (N_6394,N_3395,N_703);
or U6395 (N_6395,N_112,N_2483);
nand U6396 (N_6396,N_3479,N_4118);
nand U6397 (N_6397,N_4482,N_237);
nor U6398 (N_6398,N_2305,N_1960);
nor U6399 (N_6399,N_443,N_1379);
nand U6400 (N_6400,N_4735,N_1438);
xnor U6401 (N_6401,N_2355,N_4614);
and U6402 (N_6402,N_2520,N_4626);
or U6403 (N_6403,N_392,N_4229);
and U6404 (N_6404,N_1964,N_1937);
or U6405 (N_6405,N_2709,N_871);
or U6406 (N_6406,N_2113,N_726);
nand U6407 (N_6407,N_1288,N_3778);
xor U6408 (N_6408,N_4491,N_2461);
or U6409 (N_6409,N_3383,N_3576);
and U6410 (N_6410,N_4412,N_620);
nor U6411 (N_6411,N_3599,N_170);
xor U6412 (N_6412,N_2404,N_1158);
nor U6413 (N_6413,N_349,N_1264);
nor U6414 (N_6414,N_1130,N_56);
nor U6415 (N_6415,N_1377,N_575);
or U6416 (N_6416,N_568,N_2609);
nand U6417 (N_6417,N_2153,N_1586);
nor U6418 (N_6418,N_3917,N_2062);
or U6419 (N_6419,N_3546,N_3840);
or U6420 (N_6420,N_4043,N_1785);
or U6421 (N_6421,N_252,N_3933);
nor U6422 (N_6422,N_4061,N_2771);
nor U6423 (N_6423,N_3789,N_828);
or U6424 (N_6424,N_2462,N_3137);
xnor U6425 (N_6425,N_4353,N_1724);
and U6426 (N_6426,N_3931,N_2314);
nand U6427 (N_6427,N_1425,N_3677);
xor U6428 (N_6428,N_1058,N_253);
and U6429 (N_6429,N_4990,N_0);
nand U6430 (N_6430,N_4031,N_784);
xnor U6431 (N_6431,N_4103,N_1700);
nand U6432 (N_6432,N_2385,N_139);
nand U6433 (N_6433,N_1707,N_4603);
xor U6434 (N_6434,N_2450,N_4279);
and U6435 (N_6435,N_4339,N_685);
nand U6436 (N_6436,N_823,N_1773);
and U6437 (N_6437,N_4405,N_2980);
and U6438 (N_6438,N_1043,N_4993);
or U6439 (N_6439,N_1198,N_4901);
nor U6440 (N_6440,N_3964,N_1727);
nand U6441 (N_6441,N_2904,N_4021);
nor U6442 (N_6442,N_2048,N_2422);
nand U6443 (N_6443,N_3909,N_3993);
nor U6444 (N_6444,N_3037,N_1784);
and U6445 (N_6445,N_3244,N_4601);
xnor U6446 (N_6446,N_1991,N_1399);
xnor U6447 (N_6447,N_1177,N_1272);
or U6448 (N_6448,N_1254,N_1718);
or U6449 (N_6449,N_154,N_3514);
nor U6450 (N_6450,N_778,N_3175);
and U6451 (N_6451,N_3019,N_1697);
nor U6452 (N_6452,N_4539,N_3686);
and U6453 (N_6453,N_3146,N_2838);
or U6454 (N_6454,N_3669,N_2491);
nor U6455 (N_6455,N_886,N_1067);
and U6456 (N_6456,N_4592,N_218);
nor U6457 (N_6457,N_4779,N_1674);
and U6458 (N_6458,N_1735,N_635);
nand U6459 (N_6459,N_1828,N_42);
and U6460 (N_6460,N_4932,N_2067);
nor U6461 (N_6461,N_3081,N_3842);
nand U6462 (N_6462,N_4857,N_3401);
and U6463 (N_6463,N_201,N_1373);
and U6464 (N_6464,N_244,N_3071);
xor U6465 (N_6465,N_4672,N_1351);
or U6466 (N_6466,N_2194,N_3818);
nor U6467 (N_6467,N_1488,N_3907);
xor U6468 (N_6468,N_1790,N_3796);
nand U6469 (N_6469,N_3279,N_547);
xor U6470 (N_6470,N_3858,N_107);
xnor U6471 (N_6471,N_4866,N_4840);
nor U6472 (N_6472,N_3658,N_127);
and U6473 (N_6473,N_1887,N_3230);
and U6474 (N_6474,N_4509,N_848);
nand U6475 (N_6475,N_2588,N_2734);
xor U6476 (N_6476,N_1729,N_4917);
xnor U6477 (N_6477,N_3505,N_4438);
or U6478 (N_6478,N_4668,N_1380);
xnor U6479 (N_6479,N_3459,N_2908);
or U6480 (N_6480,N_203,N_1656);
or U6481 (N_6481,N_646,N_2718);
nor U6482 (N_6482,N_3151,N_2880);
and U6483 (N_6483,N_800,N_3500);
or U6484 (N_6484,N_1788,N_2715);
nand U6485 (N_6485,N_2567,N_4640);
nor U6486 (N_6486,N_4220,N_2821);
xor U6487 (N_6487,N_4529,N_4300);
and U6488 (N_6488,N_3927,N_1639);
or U6489 (N_6489,N_2401,N_2985);
xnor U6490 (N_6490,N_698,N_3853);
nor U6491 (N_6491,N_3283,N_1813);
and U6492 (N_6492,N_4213,N_32);
nand U6493 (N_6493,N_3749,N_132);
and U6494 (N_6494,N_403,N_1546);
nand U6495 (N_6495,N_1313,N_52);
and U6496 (N_6496,N_4162,N_4380);
and U6497 (N_6497,N_2137,N_3612);
nor U6498 (N_6498,N_2554,N_4280);
and U6499 (N_6499,N_4714,N_180);
and U6500 (N_6500,N_1731,N_2172);
nor U6501 (N_6501,N_257,N_3828);
xor U6502 (N_6502,N_591,N_2358);
or U6503 (N_6503,N_3054,N_4468);
or U6504 (N_6504,N_2501,N_2101);
and U6505 (N_6505,N_4893,N_1923);
nor U6506 (N_6506,N_4711,N_982);
xnor U6507 (N_6507,N_3537,N_2387);
and U6508 (N_6508,N_3883,N_2164);
nor U6509 (N_6509,N_4941,N_625);
xnor U6510 (N_6510,N_3649,N_482);
and U6511 (N_6511,N_4968,N_755);
and U6512 (N_6512,N_2065,N_4325);
nand U6513 (N_6513,N_1795,N_4376);
nor U6514 (N_6514,N_1836,N_2804);
nor U6515 (N_6515,N_1911,N_2789);
and U6516 (N_6516,N_2587,N_4567);
and U6517 (N_6517,N_2292,N_191);
nand U6518 (N_6518,N_3991,N_4465);
nor U6519 (N_6519,N_4849,N_4984);
or U6520 (N_6520,N_1200,N_4519);
nand U6521 (N_6521,N_4415,N_2199);
xnor U6522 (N_6522,N_505,N_2652);
nor U6523 (N_6523,N_3113,N_3220);
nor U6524 (N_6524,N_928,N_3708);
or U6525 (N_6525,N_98,N_507);
nand U6526 (N_6526,N_2472,N_922);
nand U6527 (N_6527,N_3426,N_3000);
nor U6528 (N_6528,N_93,N_1266);
or U6529 (N_6529,N_3934,N_3913);
nand U6530 (N_6530,N_4808,N_284);
or U6531 (N_6531,N_1576,N_3441);
xor U6532 (N_6532,N_3582,N_4853);
or U6533 (N_6533,N_2097,N_1699);
nand U6534 (N_6534,N_231,N_4970);
xnor U6535 (N_6535,N_2249,N_2544);
xnor U6536 (N_6536,N_246,N_515);
nor U6537 (N_6537,N_440,N_2720);
nand U6538 (N_6538,N_4271,N_1622);
and U6539 (N_6539,N_596,N_2915);
nand U6540 (N_6540,N_2955,N_3196);
or U6541 (N_6541,N_2624,N_2991);
xnor U6542 (N_6542,N_477,N_3586);
nor U6543 (N_6543,N_3140,N_3878);
nand U6544 (N_6544,N_4000,N_143);
and U6545 (N_6545,N_2471,N_4273);
and U6546 (N_6546,N_4639,N_3661);
or U6547 (N_6547,N_2111,N_3076);
and U6548 (N_6548,N_225,N_3831);
nand U6549 (N_6549,N_261,N_4900);
and U6550 (N_6550,N_626,N_3337);
or U6551 (N_6551,N_1180,N_55);
or U6552 (N_6552,N_2692,N_192);
xor U6553 (N_6553,N_44,N_4890);
and U6554 (N_6554,N_2911,N_2532);
nor U6555 (N_6555,N_2291,N_1979);
or U6556 (N_6556,N_2984,N_1726);
or U6557 (N_6557,N_504,N_656);
nor U6558 (N_6558,N_769,N_4594);
nor U6559 (N_6559,N_9,N_1362);
and U6560 (N_6560,N_2072,N_2685);
xnor U6561 (N_6561,N_2243,N_826);
and U6562 (N_6562,N_3811,N_3506);
or U6563 (N_6563,N_1900,N_3205);
nand U6564 (N_6564,N_4319,N_712);
and U6565 (N_6565,N_3347,N_1355);
nor U6566 (N_6566,N_4707,N_4769);
nand U6567 (N_6567,N_1696,N_1547);
or U6568 (N_6568,N_3080,N_2467);
and U6569 (N_6569,N_2867,N_2862);
xnor U6570 (N_6570,N_1493,N_361);
or U6571 (N_6571,N_3034,N_1099);
xnor U6572 (N_6572,N_1163,N_4095);
nor U6573 (N_6573,N_1862,N_3463);
nor U6574 (N_6574,N_4099,N_903);
nand U6575 (N_6575,N_1868,N_1123);
xnor U6576 (N_6576,N_2646,N_691);
nand U6577 (N_6577,N_1376,N_687);
nand U6578 (N_6578,N_1671,N_3033);
and U6579 (N_6579,N_1162,N_4114);
xor U6580 (N_6580,N_1736,N_4446);
nand U6581 (N_6581,N_1610,N_821);
nand U6582 (N_6582,N_4035,N_3583);
and U6583 (N_6583,N_1417,N_1890);
nand U6584 (N_6584,N_4502,N_1584);
nand U6585 (N_6585,N_2879,N_4256);
nor U6586 (N_6586,N_4904,N_136);
nor U6587 (N_6587,N_994,N_288);
xor U6588 (N_6588,N_1473,N_3932);
and U6589 (N_6589,N_1450,N_2548);
xnor U6590 (N_6590,N_1187,N_995);
or U6591 (N_6591,N_602,N_2248);
or U6592 (N_6592,N_153,N_2644);
nor U6593 (N_6593,N_2963,N_4317);
and U6594 (N_6594,N_4554,N_4758);
xnor U6595 (N_6595,N_1190,N_4466);
xnor U6596 (N_6596,N_291,N_24);
or U6597 (N_6597,N_2447,N_4794);
and U6598 (N_6598,N_122,N_3345);
or U6599 (N_6599,N_1418,N_2303);
xor U6600 (N_6600,N_4650,N_2562);
nor U6601 (N_6601,N_1339,N_1275);
and U6602 (N_6602,N_2055,N_2171);
nor U6603 (N_6603,N_328,N_793);
or U6604 (N_6604,N_3896,N_4323);
or U6605 (N_6605,N_2679,N_4778);
nand U6606 (N_6606,N_941,N_631);
nand U6607 (N_6607,N_4507,N_1778);
nor U6608 (N_6608,N_2649,N_3319);
or U6609 (N_6609,N_2104,N_1792);
or U6610 (N_6610,N_2476,N_654);
nand U6611 (N_6611,N_2017,N_536);
nor U6612 (N_6612,N_3346,N_2210);
nor U6613 (N_6613,N_4320,N_1680);
or U6614 (N_6614,N_3725,N_1831);
and U6615 (N_6615,N_875,N_4957);
or U6616 (N_6616,N_752,N_3445);
or U6617 (N_6617,N_2032,N_1243);
nand U6618 (N_6618,N_2983,N_4371);
nand U6619 (N_6619,N_1114,N_1030);
xnor U6620 (N_6620,N_665,N_2597);
or U6621 (N_6621,N_1470,N_1138);
nor U6622 (N_6622,N_4282,N_102);
and U6623 (N_6623,N_2361,N_872);
and U6624 (N_6624,N_2330,N_3042);
and U6625 (N_6625,N_3980,N_3254);
and U6626 (N_6626,N_412,N_3362);
nor U6627 (N_6627,N_3869,N_1988);
nand U6628 (N_6628,N_2090,N_676);
or U6629 (N_6629,N_650,N_3303);
nand U6630 (N_6630,N_4347,N_4950);
nor U6631 (N_6631,N_1557,N_3440);
nor U6632 (N_6632,N_3429,N_3170);
xnor U6633 (N_6633,N_1921,N_2078);
nand U6634 (N_6634,N_1550,N_4557);
nand U6635 (N_6635,N_13,N_220);
nor U6636 (N_6636,N_1125,N_240);
or U6637 (N_6637,N_1490,N_454);
nor U6638 (N_6638,N_2222,N_2123);
nor U6639 (N_6639,N_2931,N_4392);
xnor U6640 (N_6640,N_641,N_2056);
nand U6641 (N_6641,N_2304,N_4196);
and U6642 (N_6642,N_1938,N_318);
nor U6643 (N_6643,N_1467,N_457);
and U6644 (N_6644,N_2043,N_3959);
or U6645 (N_6645,N_4931,N_1775);
nand U6646 (N_6646,N_1705,N_4294);
or U6647 (N_6647,N_498,N_2940);
xor U6648 (N_6648,N_4565,N_860);
nor U6649 (N_6649,N_2815,N_3056);
and U6650 (N_6650,N_385,N_4523);
nor U6651 (N_6651,N_3201,N_2257);
or U6652 (N_6652,N_2761,N_2375);
or U6653 (N_6653,N_4881,N_280);
xor U6654 (N_6654,N_4195,N_3718);
and U6655 (N_6655,N_3750,N_2312);
and U6656 (N_6656,N_4449,N_81);
or U6657 (N_6657,N_1390,N_2216);
nand U6658 (N_6658,N_684,N_799);
nor U6659 (N_6659,N_4766,N_2254);
and U6660 (N_6660,N_516,N_2591);
xnor U6661 (N_6661,N_2828,N_3644);
and U6662 (N_6662,N_2555,N_4807);
xnor U6663 (N_6663,N_3235,N_3887);
xnor U6664 (N_6664,N_442,N_104);
nor U6665 (N_6665,N_4835,N_3270);
and U6666 (N_6666,N_4259,N_213);
and U6667 (N_6667,N_352,N_4313);
xnor U6668 (N_6668,N_3647,N_863);
nand U6669 (N_6669,N_179,N_3808);
nor U6670 (N_6670,N_2791,N_4044);
and U6671 (N_6671,N_3144,N_3664);
xnor U6672 (N_6672,N_1452,N_57);
nor U6673 (N_6673,N_4828,N_117);
nor U6674 (N_6674,N_188,N_3608);
nor U6675 (N_6675,N_4179,N_4346);
and U6676 (N_6676,N_480,N_419);
and U6677 (N_6677,N_837,N_3945);
nor U6678 (N_6678,N_558,N_305);
xnor U6679 (N_6679,N_1137,N_1064);
nand U6680 (N_6680,N_1884,N_1793);
xnor U6681 (N_6681,N_2139,N_4447);
nor U6682 (N_6682,N_4701,N_1909);
and U6683 (N_6683,N_4467,N_383);
nand U6684 (N_6684,N_38,N_1074);
nor U6685 (N_6685,N_1235,N_932);
xor U6686 (N_6686,N_1382,N_2841);
or U6687 (N_6687,N_780,N_2077);
or U6688 (N_6688,N_3783,N_65);
nor U6689 (N_6689,N_713,N_542);
nor U6690 (N_6690,N_2364,N_251);
and U6691 (N_6691,N_2775,N_3118);
nand U6692 (N_6692,N_1307,N_3207);
xnor U6693 (N_6693,N_3391,N_3833);
nand U6694 (N_6694,N_1206,N_553);
nor U6695 (N_6695,N_594,N_1585);
xor U6696 (N_6696,N_915,N_2694);
nand U6697 (N_6697,N_411,N_3487);
nor U6698 (N_6698,N_158,N_1653);
nand U6699 (N_6699,N_1601,N_4991);
or U6700 (N_6700,N_2310,N_4980);
xor U6701 (N_6701,N_2944,N_2152);
or U6702 (N_6702,N_4030,N_2379);
nand U6703 (N_6703,N_3897,N_494);
and U6704 (N_6704,N_1226,N_66);
nor U6705 (N_6705,N_3947,N_1962);
nor U6706 (N_6706,N_3890,N_2670);
nor U6707 (N_6707,N_2992,N_2872);
and U6708 (N_6708,N_4982,N_45);
and U6709 (N_6709,N_1455,N_4176);
nor U6710 (N_6710,N_1817,N_34);
xor U6711 (N_6711,N_2150,N_2005);
and U6712 (N_6712,N_2808,N_380);
and U6713 (N_6713,N_4441,N_1827);
nand U6714 (N_6714,N_1370,N_2899);
or U6715 (N_6715,N_1153,N_1965);
and U6716 (N_6716,N_4573,N_1025);
or U6717 (N_6717,N_818,N_765);
nor U6718 (N_6718,N_4363,N_529);
xor U6719 (N_6719,N_4026,N_1853);
nand U6720 (N_6720,N_4348,N_3900);
or U6721 (N_6721,N_3795,N_3812);
and U6722 (N_6722,N_4013,N_3090);
nand U6723 (N_6723,N_4512,N_4110);
xnor U6724 (N_6724,N_168,N_1918);
nand U6725 (N_6725,N_3662,N_2560);
and U6726 (N_6726,N_1408,N_1083);
xor U6727 (N_6727,N_2035,N_4836);
nand U6728 (N_6728,N_368,N_3419);
nand U6729 (N_6729,N_2068,N_1214);
or U6730 (N_6730,N_4068,N_929);
and U6731 (N_6731,N_6,N_3562);
nor U6732 (N_6732,N_1919,N_4844);
and U6733 (N_6733,N_2674,N_586);
nor U6734 (N_6734,N_4136,N_1329);
xor U6735 (N_6735,N_3155,N_4459);
nand U6736 (N_6736,N_2276,N_4677);
or U6737 (N_6737,N_2020,N_1);
nor U6738 (N_6738,N_1262,N_1066);
xor U6739 (N_6739,N_3703,N_4108);
xor U6740 (N_6740,N_1686,N_3231);
and U6741 (N_6741,N_4125,N_4703);
or U6742 (N_6742,N_4218,N_1033);
nand U6743 (N_6743,N_3029,N_115);
and U6744 (N_6744,N_4555,N_1302);
or U6745 (N_6745,N_3867,N_2631);
nor U6746 (N_6746,N_3212,N_1325);
xnor U6747 (N_6747,N_1663,N_3547);
nor U6748 (N_6748,N_2876,N_3886);
nor U6749 (N_6749,N_1961,N_3994);
or U6750 (N_6750,N_4096,N_1485);
nand U6751 (N_6751,N_3211,N_1716);
or U6752 (N_6752,N_3698,N_2157);
nor U6753 (N_6753,N_228,N_2315);
nand U6754 (N_6754,N_2428,N_1268);
nor U6755 (N_6755,N_4713,N_4969);
and U6756 (N_6756,N_1545,N_2578);
and U6757 (N_6757,N_1317,N_1371);
nor U6758 (N_6758,N_379,N_4019);
nor U6759 (N_6759,N_3652,N_2189);
or U6760 (N_6760,N_3369,N_417);
or U6761 (N_6761,N_2307,N_1459);
or U6762 (N_6762,N_4795,N_2496);
nor U6763 (N_6763,N_2372,N_2799);
nand U6764 (N_6764,N_4016,N_983);
or U6765 (N_6765,N_1679,N_3470);
and U6766 (N_6766,N_3929,N_189);
and U6767 (N_6767,N_508,N_1751);
or U6768 (N_6768,N_2905,N_611);
or U6769 (N_6769,N_2076,N_2197);
or U6770 (N_6770,N_4832,N_1426);
nand U6771 (N_6771,N_2488,N_1978);
nor U6772 (N_6772,N_2161,N_4199);
and U6773 (N_6773,N_1995,N_1794);
and U6774 (N_6774,N_2046,N_4928);
nor U6775 (N_6775,N_2207,N_2579);
xnor U6776 (N_6776,N_893,N_1437);
nor U6777 (N_6777,N_1135,N_3174);
or U6778 (N_6778,N_1481,N_2184);
nor U6779 (N_6779,N_972,N_4809);
nor U6780 (N_6780,N_583,N_3364);
nand U6781 (N_6781,N_1222,N_1081);
and U6782 (N_6782,N_3482,N_4894);
xnor U6783 (N_6783,N_4861,N_2669);
and U6784 (N_6784,N_2782,N_279);
nor U6785 (N_6785,N_1106,N_2026);
xor U6786 (N_6786,N_4895,N_1046);
nor U6787 (N_6787,N_190,N_678);
xnor U6788 (N_6788,N_3006,N_3739);
and U6789 (N_6789,N_2708,N_1830);
and U6790 (N_6790,N_1678,N_4864);
nand U6791 (N_6791,N_4896,N_2620);
nand U6792 (N_6792,N_2328,N_1543);
nand U6793 (N_6793,N_4782,N_791);
xor U6794 (N_6794,N_1028,N_1646);
xor U6795 (N_6795,N_3095,N_4740);
xor U6796 (N_6796,N_3407,N_2961);
nor U6797 (N_6797,N_2396,N_4301);
or U6798 (N_6798,N_4542,N_838);
or U6799 (N_6799,N_4006,N_2971);
nand U6800 (N_6800,N_4883,N_1127);
nand U6801 (N_6801,N_4228,N_2235);
nand U6802 (N_6802,N_4983,N_1829);
and U6803 (N_6803,N_1632,N_1178);
nand U6804 (N_6804,N_873,N_3274);
or U6805 (N_6805,N_4967,N_867);
nand U6806 (N_6806,N_89,N_149);
nand U6807 (N_6807,N_693,N_4954);
and U6808 (N_6808,N_2241,N_3692);
and U6809 (N_6809,N_4860,N_1749);
nor U6810 (N_6810,N_1623,N_3058);
or U6811 (N_6811,N_273,N_2633);
and U6812 (N_6812,N_2423,N_1285);
nand U6813 (N_6813,N_2781,N_3843);
nand U6814 (N_6814,N_4643,N_916);
xnor U6815 (N_6815,N_4291,N_1115);
xor U6816 (N_6816,N_1031,N_1036);
nand U6817 (N_6817,N_1876,N_4538);
and U6818 (N_6818,N_1429,N_4818);
xor U6819 (N_6819,N_315,N_1013);
nand U6820 (N_6820,N_2684,N_4925);
and U6821 (N_6821,N_2777,N_887);
and U6822 (N_6822,N_4364,N_27);
nor U6823 (N_6823,N_2206,N_4113);
nor U6824 (N_6824,N_773,N_3321);
xnor U6825 (N_6825,N_2402,N_4506);
nand U6826 (N_6826,N_1101,N_2306);
nor U6827 (N_6827,N_4621,N_4408);
or U6828 (N_6828,N_560,N_1633);
nor U6829 (N_6829,N_3920,N_1612);
and U6830 (N_6830,N_3903,N_4646);
nor U6831 (N_6831,N_3946,N_426);
nor U6832 (N_6832,N_4025,N_3049);
xor U6833 (N_6833,N_3352,N_1682);
xor U6834 (N_6834,N_214,N_4622);
and U6835 (N_6835,N_749,N_1478);
and U6836 (N_6836,N_2822,N_3879);
xnor U6837 (N_6837,N_2610,N_513);
nand U6838 (N_6838,N_4561,N_2686);
nor U6839 (N_6839,N_2042,N_267);
and U6840 (N_6840,N_287,N_710);
nor U6841 (N_6841,N_3722,N_451);
xor U6842 (N_6842,N_3824,N_756);
nand U6843 (N_6843,N_4154,N_1160);
nand U6844 (N_6844,N_3666,N_2512);
nor U6845 (N_6845,N_917,N_1227);
or U6846 (N_6846,N_3420,N_1038);
and U6847 (N_6847,N_413,N_934);
nor U6848 (N_6848,N_4564,N_2060);
nand U6849 (N_6849,N_2917,N_4920);
nor U6850 (N_6850,N_1967,N_3699);
nor U6851 (N_6851,N_60,N_2166);
xor U6852 (N_6852,N_2788,N_3836);
or U6853 (N_6853,N_3216,N_3373);
nand U6854 (N_6854,N_3465,N_2682);
xnor U6855 (N_6855,N_2589,N_4386);
or U6856 (N_6856,N_1413,N_2572);
and U6857 (N_6857,N_1581,N_2653);
nand U6858 (N_6858,N_4373,N_651);
and U6859 (N_6859,N_2611,N_2217);
or U6860 (N_6860,N_129,N_3072);
nor U6861 (N_6861,N_4985,N_3655);
or U6862 (N_6862,N_4733,N_1598);
and U6863 (N_6863,N_1026,N_4710);
nor U6864 (N_6864,N_2884,N_1444);
xor U6865 (N_6865,N_431,N_3791);
or U6866 (N_6866,N_796,N_522);
or U6867 (N_6867,N_212,N_1049);
or U6868 (N_6868,N_3208,N_2570);
and U6869 (N_6869,N_3104,N_1971);
xnor U6870 (N_6870,N_2457,N_3070);
xor U6871 (N_6871,N_3355,N_598);
xnor U6872 (N_6872,N_2689,N_3524);
or U6873 (N_6873,N_4788,N_3338);
and U6874 (N_6874,N_4624,N_150);
nor U6875 (N_6875,N_2029,N_1832);
nand U6876 (N_6876,N_266,N_1618);
nor U6877 (N_6877,N_1120,N_2545);
and U6878 (N_6878,N_4576,N_2964);
nor U6879 (N_6879,N_1242,N_2864);
nor U6880 (N_6880,N_3316,N_1185);
and U6881 (N_6881,N_2742,N_3820);
nor U6882 (N_6882,N_1774,N_37);
nand U6883 (N_6883,N_1143,N_942);
and U6884 (N_6884,N_4934,N_1082);
xnor U6885 (N_6885,N_4946,N_977);
or U6886 (N_6886,N_4198,N_3250);
xor U6887 (N_6887,N_87,N_461);
or U6888 (N_6888,N_1974,N_1561);
and U6889 (N_6889,N_204,N_3967);
xor U6890 (N_6890,N_2758,N_338);
and U6891 (N_6891,N_373,N_2656);
nand U6892 (N_6892,N_4460,N_4842);
xor U6893 (N_6893,N_3573,N_2500);
xor U6894 (N_6894,N_4485,N_1341);
nor U6895 (N_6895,N_4060,N_4726);
and U6896 (N_6896,N_3729,N_4201);
and U6897 (N_6897,N_572,N_753);
xnor U6898 (N_6898,N_768,N_2818);
xor U6899 (N_6899,N_26,N_2518);
or U6900 (N_6900,N_3055,N_1914);
or U6901 (N_6901,N_1424,N_518);
nand U6902 (N_6902,N_1094,N_4897);
or U6903 (N_6903,N_1820,N_1239);
xnor U6904 (N_6904,N_761,N_2629);
xor U6905 (N_6905,N_4642,N_1734);
nor U6906 (N_6906,N_3062,N_785);
nand U6907 (N_6907,N_2833,N_3309);
or U6908 (N_6908,N_4365,N_3861);
or U6909 (N_6909,N_812,N_1489);
nand U6910 (N_6910,N_1730,N_4975);
xnor U6911 (N_6911,N_1989,N_1250);
xnor U6912 (N_6912,N_320,N_548);
nand U6913 (N_6913,N_4400,N_1513);
nand U6914 (N_6914,N_4577,N_226);
nor U6915 (N_6915,N_3868,N_819);
and U6916 (N_6916,N_2730,N_847);
xnor U6917 (N_6917,N_1524,N_1231);
and U6918 (N_6918,N_3253,N_2255);
nand U6919 (N_6919,N_14,N_699);
nand U6920 (N_6920,N_2515,N_1972);
or U6921 (N_6921,N_4330,N_2353);
nor U6922 (N_6922,N_1395,N_4328);
and U6923 (N_6923,N_2998,N_2021);
nor U6924 (N_6924,N_4127,N_2262);
or U6925 (N_6925,N_3238,N_3848);
nand U6926 (N_6926,N_4715,N_1599);
nand U6927 (N_6927,N_844,N_2407);
or U6928 (N_6928,N_4743,N_3510);
xnor U6929 (N_6929,N_3203,N_4884);
nand U6930 (N_6930,N_835,N_3082);
nand U6931 (N_6931,N_1256,N_4235);
or U6932 (N_6932,N_2051,N_3713);
and U6933 (N_6933,N_4337,N_3278);
xor U6934 (N_6934,N_4632,N_4004);
xor U6935 (N_6935,N_3925,N_897);
and U6936 (N_6936,N_952,N_2972);
or U6937 (N_6937,N_2019,N_1824);
and U6938 (N_6938,N_1638,N_2827);
and U6939 (N_6939,N_3584,N_593);
or U6940 (N_6940,N_4211,N_1789);
xor U6941 (N_6941,N_3714,N_1525);
or U6942 (N_6942,N_599,N_351);
nor U6943 (N_6943,N_2839,N_851);
or U6944 (N_6944,N_2538,N_2763);
nor U6945 (N_6945,N_3628,N_1951);
nand U6946 (N_6946,N_2696,N_806);
xnor U6947 (N_6947,N_1635,N_1375);
nor U6948 (N_6948,N_2535,N_2191);
and U6949 (N_6949,N_1449,N_247);
xnor U6950 (N_6950,N_1798,N_3481);
nor U6951 (N_6951,N_4239,N_1801);
nand U6952 (N_6952,N_3905,N_3741);
nor U6953 (N_6953,N_2038,N_1845);
nor U6954 (N_6954,N_277,N_4443);
or U6955 (N_6955,N_1435,N_3995);
xnor U6956 (N_6956,N_2519,N_1278);
and U6957 (N_6957,N_1689,N_47);
or U6958 (N_6958,N_3832,N_2486);
xnor U6959 (N_6959,N_3223,N_1692);
xor U6960 (N_6960,N_1219,N_1217);
and U6961 (N_6961,N_2916,N_4562);
nor U6962 (N_6962,N_4717,N_2008);
and U6963 (N_6963,N_798,N_165);
or U6964 (N_6964,N_1161,N_2061);
or U6965 (N_6965,N_4299,N_1892);
nand U6966 (N_6966,N_3014,N_3100);
nand U6967 (N_6967,N_3893,N_1436);
nor U6968 (N_6968,N_2264,N_2230);
nor U6969 (N_6969,N_1659,N_2681);
or U6970 (N_6970,N_278,N_2479);
xnor U6971 (N_6971,N_4804,N_4101);
xor U6972 (N_6972,N_2959,N_3935);
or U6973 (N_6973,N_1300,N_290);
or U6974 (N_6974,N_2637,N_3987);
nor U6975 (N_6975,N_3001,N_2279);
nand U6976 (N_6976,N_3268,N_4444);
nor U6977 (N_6977,N_3431,N_1717);
xor U6978 (N_6978,N_1996,N_3109);
and U6979 (N_6979,N_286,N_3295);
nand U6980 (N_6980,N_178,N_4653);
nor U6981 (N_6981,N_4752,N_3660);
xor U6982 (N_6982,N_4566,N_1889);
or U6983 (N_6983,N_4587,N_2922);
and U6984 (N_6984,N_4356,N_2866);
nand U6985 (N_6985,N_1772,N_892);
or U6986 (N_6986,N_1888,N_3217);
nor U6987 (N_6987,N_3180,N_1969);
and U6988 (N_6988,N_59,N_827);
nor U6989 (N_6989,N_1521,N_2592);
xnor U6990 (N_6990,N_3492,N_4698);
nand U6991 (N_6991,N_3417,N_4497);
nand U6992 (N_6992,N_1453,N_1768);
nand U6993 (N_6993,N_1119,N_4226);
xnor U6994 (N_6994,N_219,N_839);
or U6995 (N_6995,N_2006,N_4286);
or U6996 (N_6996,N_467,N_4796);
nand U6997 (N_6997,N_3409,N_2506);
xnor U6998 (N_6998,N_4903,N_4878);
and U6999 (N_6999,N_4527,N_2105);
xnor U7000 (N_7000,N_3255,N_2851);
xnor U7001 (N_7001,N_1925,N_717);
nor U7002 (N_7002,N_1209,N_4318);
and U7003 (N_7003,N_2460,N_3928);
nand U7004 (N_7004,N_1886,N_193);
xor U7005 (N_7005,N_1367,N_4357);
nand U7006 (N_7006,N_906,N_2470);
nand U7007 (N_7007,N_3298,N_3035);
xor U7008 (N_7008,N_4608,N_2584);
or U7009 (N_7009,N_4695,N_3643);
nor U7010 (N_7010,N_3491,N_958);
nor U7011 (N_7011,N_632,N_1565);
and U7012 (N_7012,N_3018,N_1765);
and U7013 (N_7013,N_2795,N_3408);
or U7014 (N_7014,N_126,N_530);
or U7015 (N_7015,N_1328,N_4210);
nor U7016 (N_7016,N_1286,N_2546);
xnor U7017 (N_7017,N_4454,N_2693);
nand U7018 (N_7018,N_1769,N_1414);
nand U7019 (N_7019,N_3157,N_3423);
or U7020 (N_7020,N_633,N_50);
and U7021 (N_7021,N_2343,N_689);
nor U7022 (N_7022,N_3515,N_316);
xor U7023 (N_7023,N_62,N_3746);
or U7024 (N_7024,N_4938,N_391);
nor U7025 (N_7025,N_1169,N_563);
nand U7026 (N_7026,N_604,N_3579);
nand U7027 (N_7027,N_2331,N_4654);
xnor U7028 (N_7028,N_2009,N_4001);
or U7029 (N_7029,N_1818,N_3657);
and U7030 (N_7030,N_2135,N_2647);
xnor U7031 (N_7031,N_600,N_1005);
and U7032 (N_7032,N_1240,N_369);
xnor U7033 (N_7033,N_868,N_3577);
xnor U7034 (N_7034,N_846,N_4129);
nor U7035 (N_7035,N_2541,N_1068);
or U7036 (N_7036,N_3730,N_634);
or U7037 (N_7037,N_645,N_3948);
nand U7038 (N_7038,N_2100,N_1040);
or U7039 (N_7039,N_4741,N_4604);
nor U7040 (N_7040,N_3841,N_4734);
or U7041 (N_7041,N_889,N_4876);
xor U7042 (N_7042,N_3341,N_2433);
or U7043 (N_7043,N_1928,N_418);
nor U7044 (N_7044,N_1168,N_606);
nor U7045 (N_7045,N_4730,N_4148);
nand U7046 (N_7046,N_334,N_580);
and U7047 (N_7047,N_11,N_3737);
nand U7048 (N_7048,N_1959,N_2481);
nor U7049 (N_7049,N_19,N_653);
xor U7050 (N_7050,N_2142,N_997);
nor U7051 (N_7051,N_4919,N_2196);
and U7052 (N_7052,N_3271,N_3443);
or U7053 (N_7053,N_3857,N_144);
or U7054 (N_7054,N_210,N_4531);
xor U7055 (N_7055,N_2889,N_708);
xnor U7056 (N_7056,N_4233,N_2651);
and U7057 (N_7057,N_3462,N_2453);
or U7058 (N_7058,N_491,N_1519);
xnor U7059 (N_7059,N_3710,N_116);
nor U7060 (N_7060,N_2127,N_3590);
xnor U7061 (N_7061,N_3176,N_3792);
xor U7062 (N_7062,N_4495,N_2024);
xor U7063 (N_7063,N_525,N_3285);
nor U7064 (N_7064,N_1740,N_3213);
or U7065 (N_7065,N_1323,N_2607);
nand U7066 (N_7066,N_993,N_3410);
or U7067 (N_7067,N_1676,N_3682);
nor U7068 (N_7068,N_3075,N_2699);
xnor U7069 (N_7069,N_1463,N_4556);
nand U7070 (N_7070,N_3195,N_3439);
nor U7071 (N_7071,N_1293,N_123);
nor U7072 (N_7072,N_3102,N_649);
nor U7073 (N_7073,N_950,N_348);
or U7074 (N_7074,N_931,N_1799);
nor U7075 (N_7075,N_2400,N_3359);
nand U7076 (N_7076,N_1927,N_3403);
nor U7077 (N_7077,N_3233,N_2529);
nand U7078 (N_7078,N_3277,N_48);
xnor U7079 (N_7079,N_555,N_3926);
xnor U7080 (N_7080,N_4644,N_3970);
or U7081 (N_7081,N_3110,N_3676);
nand U7082 (N_7082,N_537,N_4819);
nor U7083 (N_7083,N_1000,N_2432);
nor U7084 (N_7084,N_2368,N_427);
or U7085 (N_7085,N_1349,N_333);
nand U7086 (N_7086,N_1271,N_3184);
and U7087 (N_7087,N_1510,N_4912);
xor U7088 (N_7088,N_616,N_1897);
and U7089 (N_7089,N_1188,N_1807);
and U7090 (N_7090,N_4297,N_61);
nor U7091 (N_7091,N_1050,N_2367);
or U7092 (N_7092,N_1430,N_3575);
nor U7093 (N_7093,N_432,N_3069);
nand U7094 (N_7094,N_4399,N_1385);
xnor U7095 (N_7095,N_1263,N_4484);
xnor U7096 (N_7096,N_1708,N_7);
and U7097 (N_7097,N_2626,N_1992);
and U7098 (N_7098,N_2399,N_131);
or U7099 (N_7099,N_345,N_1322);
nand U7100 (N_7100,N_271,N_1728);
and U7101 (N_7101,N_3447,N_921);
or U7102 (N_7102,N_2513,N_3143);
and U7103 (N_7103,N_4146,N_4679);
xor U7104 (N_7104,N_1968,N_4050);
nor U7105 (N_7105,N_732,N_1858);
and U7106 (N_7106,N_497,N_308);
nor U7107 (N_7107,N_2271,N_4997);
nand U7108 (N_7108,N_4427,N_464);
nor U7109 (N_7109,N_3350,N_1800);
and U7110 (N_7110,N_772,N_1344);
nor U7111 (N_7111,N_3507,N_2574);
or U7112 (N_7112,N_408,N_3777);
nand U7113 (N_7113,N_1743,N_4724);
xor U7114 (N_7114,N_554,N_1744);
nor U7115 (N_7115,N_3687,N_3461);
nor U7116 (N_7116,N_4571,N_919);
and U7117 (N_7117,N_3597,N_3067);
xor U7118 (N_7118,N_4476,N_2702);
and U7119 (N_7119,N_2677,N_25);
nor U7120 (N_7120,N_4978,N_4552);
and U7121 (N_7121,N_4613,N_2033);
nor U7122 (N_7122,N_2909,N_2514);
or U7123 (N_7123,N_3177,N_1670);
or U7124 (N_7124,N_3480,N_3569);
or U7125 (N_7125,N_3044,N_3015);
nor U7126 (N_7126,N_2269,N_3486);
and U7127 (N_7127,N_350,N_4395);
xor U7128 (N_7128,N_335,N_747);
and U7129 (N_7129,N_4172,N_2668);
nor U7130 (N_7130,N_571,N_3115);
nand U7131 (N_7131,N_4111,N_2141);
xnor U7132 (N_7132,N_4010,N_4268);
or U7133 (N_7133,N_1071,N_2796);
nand U7134 (N_7134,N_176,N_4486);
nor U7135 (N_7135,N_590,N_4732);
and U7136 (N_7136,N_4461,N_3684);
xnor U7137 (N_7137,N_1864,N_520);
xnor U7138 (N_7138,N_4651,N_1346);
and U7139 (N_7139,N_743,N_4440);
nor U7140 (N_7140,N_1780,N_638);
xnor U7141 (N_7141,N_3094,N_4391);
or U7142 (N_7142,N_759,N_4352);
or U7143 (N_7143,N_2352,N_4090);
or U7144 (N_7144,N_4039,N_3);
or U7145 (N_7145,N_1034,N_3455);
and U7146 (N_7146,N_1343,N_3382);
and U7147 (N_7147,N_3165,N_4645);
or U7148 (N_7148,N_2129,N_4480);
and U7149 (N_7149,N_1950,N_943);
and U7150 (N_7150,N_46,N_2969);
nand U7151 (N_7151,N_3438,N_3215);
and U7152 (N_7152,N_4535,N_4837);
and U7153 (N_7153,N_1165,N_1244);
nor U7154 (N_7154,N_4149,N_3122);
nand U7155 (N_7155,N_270,N_3517);
xnor U7156 (N_7156,N_3674,N_1932);
xor U7157 (N_7157,N_232,N_4736);
or U7158 (N_7158,N_3556,N_141);
nor U7159 (N_7159,N_3310,N_2484);
xor U7160 (N_7160,N_2183,N_2812);
and U7161 (N_7161,N_3087,N_2606);
nor U7162 (N_7162,N_3773,N_3503);
nor U7163 (N_7163,N_4537,N_4360);
or U7164 (N_7164,N_4078,N_453);
nand U7165 (N_7165,N_3007,N_1113);
xor U7166 (N_7166,N_4036,N_1189);
and U7167 (N_7167,N_4898,N_3632);
nand U7168 (N_7168,N_3273,N_4477);
nor U7169 (N_7169,N_1193,N_1929);
and U7170 (N_7170,N_4158,N_3010);
and U7171 (N_7171,N_1588,N_4417);
xnor U7172 (N_7172,N_118,N_1750);
and U7173 (N_7173,N_2575,N_4973);
and U7174 (N_7174,N_862,N_3732);
and U7175 (N_7175,N_4615,N_3541);
xnor U7176 (N_7176,N_4135,N_103);
and U7177 (N_7177,N_2816,N_410);
or U7178 (N_7178,N_2436,N_4332);
nand U7179 (N_7179,N_3950,N_3875);
nor U7180 (N_7180,N_3814,N_2195);
or U7181 (N_7181,N_4759,N_731);
xnor U7182 (N_7182,N_628,N_2691);
nor U7183 (N_7183,N_2201,N_425);
and U7184 (N_7184,N_4763,N_2225);
and U7185 (N_7185,N_4933,N_2384);
nand U7186 (N_7186,N_1848,N_1672);
nand U7187 (N_7187,N_2289,N_4066);
nand U7188 (N_7188,N_3617,N_2151);
nor U7189 (N_7189,N_4719,N_4692);
or U7190 (N_7190,N_173,N_3183);
nor U7191 (N_7191,N_2086,N_3940);
nand U7192 (N_7192,N_4498,N_4144);
xor U7193 (N_7193,N_458,N_519);
xnor U7194 (N_7194,N_4688,N_2509);
nand U7195 (N_7195,N_4657,N_2293);
or U7196 (N_7196,N_564,N_3091);
nand U7197 (N_7197,N_1895,N_1512);
nor U7198 (N_7198,N_4209,N_174);
xor U7199 (N_7199,N_4383,N_1954);
nand U7200 (N_7200,N_1253,N_3385);
nor U7201 (N_7201,N_3093,N_3145);
nor U7202 (N_7202,N_4549,N_657);
nand U7203 (N_7203,N_955,N_3821);
nor U7204 (N_7204,N_2813,N_4404);
xnor U7205 (N_7205,N_485,N_2752);
or U7206 (N_7206,N_3334,N_2002);
nand U7207 (N_7207,N_1173,N_899);
and U7208 (N_7208,N_2510,N_4858);
nor U7209 (N_7209,N_1631,N_372);
nor U7210 (N_7210,N_1782,N_1234);
nor U7211 (N_7211,N_4784,N_1147);
xor U7212 (N_7212,N_1416,N_1431);
and U7213 (N_7213,N_1850,N_1124);
nor U7214 (N_7214,N_151,N_4847);
and U7215 (N_7215,N_2935,N_2096);
nand U7216 (N_7216,N_4076,N_4227);
nand U7217 (N_7217,N_3064,N_4305);
and U7218 (N_7218,N_1555,N_4173);
or U7219 (N_7219,N_912,N_3047);
nor U7220 (N_7220,N_1078,N_1015);
nor U7221 (N_7221,N_4085,N_2290);
xor U7222 (N_7222,N_2273,N_2661);
and U7223 (N_7223,N_1255,N_1990);
or U7224 (N_7224,N_4911,N_1642);
xnor U7225 (N_7225,N_3901,N_3361);
or U7226 (N_7226,N_1150,N_1939);
and U7227 (N_7227,N_3598,N_3772);
nor U7228 (N_7228,N_1704,N_1758);
nor U7229 (N_7229,N_2267,N_2913);
or U7230 (N_7230,N_2495,N_984);
or U7231 (N_7231,N_2363,N_4704);
nand U7232 (N_7232,N_2794,N_1856);
xnor U7233 (N_7233,N_1977,N_4909);
xor U7234 (N_7234,N_2831,N_4455);
and U7235 (N_7235,N_815,N_4524);
and U7236 (N_7236,N_357,N_2896);
nand U7237 (N_7237,N_1520,N_2979);
xnor U7238 (N_7238,N_2180,N_4457);
nand U7239 (N_7239,N_4202,N_1477);
or U7240 (N_7240,N_3210,N_3494);
nand U7241 (N_7241,N_300,N_666);
nor U7242 (N_7242,N_716,N_2339);
or U7243 (N_7243,N_3471,N_3193);
xor U7244 (N_7244,N_3885,N_1306);
xnor U7245 (N_7245,N_3899,N_234);
nor U7246 (N_7246,N_1004,N_4316);
or U7247 (N_7247,N_4186,N_2783);
nor U7248 (N_7248,N_2950,N_3314);
nor U7249 (N_7249,N_1205,N_1661);
nand U7250 (N_7250,N_4755,N_1530);
nand U7251 (N_7251,N_3765,N_1202);
nor U7252 (N_7252,N_1311,N_4676);
nand U7253 (N_7253,N_3707,N_1752);
xor U7254 (N_7254,N_1295,N_1755);
xnor U7255 (N_7255,N_4388,N_4572);
nor U7256 (N_7256,N_1620,N_992);
nor U7257 (N_7257,N_1458,N_2011);
or U7258 (N_7258,N_2736,N_4528);
nand U7259 (N_7259,N_1880,N_2260);
xnor U7260 (N_7260,N_1930,N_4989);
nand U7261 (N_7261,N_4906,N_1763);
and U7262 (N_7262,N_577,N_3633);
nand U7263 (N_7263,N_4278,N_4606);
nor U7264 (N_7264,N_1804,N_579);
and U7265 (N_7265,N_1508,N_3448);
nor U7266 (N_7266,N_1280,N_4899);
xor U7267 (N_7267,N_1182,N_4598);
xnor U7268 (N_7268,N_1606,N_2337);
or U7269 (N_7269,N_1760,N_3779);
nor U7270 (N_7270,N_814,N_1955);
nand U7271 (N_7271,N_1572,N_4205);
nor U7272 (N_7272,N_4018,N_3112);
xor U7273 (N_7273,N_961,N_4263);
xor U7274 (N_7274,N_1396,N_4178);
nand U7275 (N_7275,N_2215,N_4070);
xnor U7276 (N_7276,N_990,N_4781);
and U7277 (N_7277,N_4069,N_4751);
nor U7278 (N_7278,N_1542,N_1365);
nor U7279 (N_7279,N_235,N_1224);
and U7280 (N_7280,N_974,N_1048);
and U7281 (N_7281,N_344,N_2707);
xnor U7282 (N_7282,N_2793,N_603);
or U7283 (N_7283,N_2525,N_3988);
and U7284 (N_7284,N_455,N_2394);
nor U7285 (N_7285,N_4483,N_449);
nor U7286 (N_7286,N_1881,N_3039);
and U7287 (N_7287,N_1484,N_1945);
nor U7288 (N_7288,N_715,N_406);
or U7289 (N_7289,N_3117,N_670);
or U7290 (N_7290,N_3998,N_3051);
nor U7291 (N_7291,N_1259,N_185);
nor U7292 (N_7292,N_3460,N_1421);
or U7293 (N_7293,N_2844,N_1540);
and U7294 (N_7294,N_4269,N_2084);
xor U7295 (N_7295,N_332,N_2970);
nand U7296 (N_7296,N_1411,N_1358);
nor U7297 (N_7297,N_3771,N_1712);
or U7298 (N_7298,N_323,N_2392);
and U7299 (N_7299,N_1948,N_1738);
nand U7300 (N_7300,N_3650,N_1834);
or U7301 (N_7301,N_229,N_4231);
xor U7302 (N_7302,N_75,N_4543);
or U7303 (N_7303,N_557,N_4274);
or U7304 (N_7304,N_4377,N_422);
or U7305 (N_7305,N_2973,N_4075);
nor U7306 (N_7306,N_1166,N_3527);
nor U7307 (N_7307,N_2116,N_2938);
or U7308 (N_7308,N_155,N_965);
and U7309 (N_7309,N_1837,N_4267);
nor U7310 (N_7310,N_1625,N_2921);
nand U7311 (N_7311,N_2932,N_1440);
and U7312 (N_7312,N_845,N_1980);
or U7313 (N_7313,N_3388,N_3430);
xor U7314 (N_7314,N_3581,N_1614);
nor U7315 (N_7315,N_3589,N_3592);
or U7316 (N_7316,N_1826,N_3810);
and U7317 (N_7317,N_4789,N_3560);
or U7318 (N_7318,N_3028,N_58);
nor U7319 (N_7319,N_1552,N_2719);
nor U7320 (N_7320,N_1210,N_3434);
and U7321 (N_7321,N_2999,N_1447);
and U7322 (N_7322,N_472,N_675);
or U7323 (N_7323,N_795,N_2571);
nor U7324 (N_7324,N_857,N_2406);
nor U7325 (N_7325,N_4366,N_3366);
xnor U7326 (N_7326,N_448,N_3793);
and U7327 (N_7327,N_3031,N_3974);
nand U7328 (N_7328,N_53,N_175);
xnor U7329 (N_7329,N_3850,N_268);
or U7330 (N_7330,N_2701,N_1141);
xor U7331 (N_7331,N_1907,N_337);
or U7332 (N_7332,N_3484,N_4128);
and U7333 (N_7333,N_166,N_147);
and U7334 (N_7334,N_948,N_3918);
nor U7335 (N_7335,N_2654,N_1475);
or U7336 (N_7336,N_2706,N_79);
xnor U7337 (N_7337,N_3585,N_2586);
and U7338 (N_7338,N_2733,N_3008);
or U7339 (N_7339,N_4469,N_119);
xor U7340 (N_7340,N_2200,N_4958);
nor U7341 (N_7341,N_569,N_4275);
and U7342 (N_7342,N_3187,N_2421);
nor U7343 (N_7343,N_435,N_1441);
nand U7344 (N_7344,N_4104,N_473);
xnor U7345 (N_7345,N_111,N_3356);
nor U7346 (N_7346,N_1879,N_2474);
nor U7347 (N_7347,N_4959,N_1443);
xor U7348 (N_7348,N_1126,N_95);
or U7349 (N_7349,N_909,N_2854);
nand U7350 (N_7350,N_3923,N_1279);
nand U7351 (N_7351,N_790,N_3336);
nor U7352 (N_7352,N_1626,N_4673);
nor U7353 (N_7353,N_521,N_2612);
and U7354 (N_7354,N_954,N_1527);
xnor U7355 (N_7355,N_4398,N_4059);
and U7356 (N_7356,N_1462,N_1318);
and U7357 (N_7357,N_1276,N_4952);
nand U7358 (N_7358,N_4203,N_2326);
nor U7359 (N_7359,N_971,N_1432);
and U7360 (N_7360,N_3764,N_49);
nand U7361 (N_7361,N_3823,N_2118);
and U7362 (N_7362,N_3862,N_4254);
nor U7363 (N_7363,N_3540,N_4811);
and U7364 (N_7364,N_3161,N_509);
nand U7365 (N_7365,N_1020,N_2138);
nand U7366 (N_7366,N_4276,N_1501);
nand U7367 (N_7367,N_2953,N_2083);
or U7368 (N_7368,N_1010,N_3985);
xnor U7369 (N_7369,N_4641,N_1604);
nor U7370 (N_7370,N_1077,N_3290);
or U7371 (N_7371,N_4261,N_4126);
nand U7372 (N_7372,N_3782,N_3433);
xor U7373 (N_7373,N_2892,N_3711);
xor U7374 (N_7374,N_3358,N_2377);
nor U7375 (N_7375,N_673,N_4456);
and U7376 (N_7376,N_3252,N_1090);
and U7377 (N_7377,N_2939,N_4949);
and U7378 (N_7378,N_4511,N_510);
nand U7379 (N_7379,N_3763,N_197);
or U7380 (N_7380,N_4716,N_4742);
xnor U7381 (N_7381,N_668,N_2974);
or U7382 (N_7382,N_3870,N_1084);
xor U7383 (N_7383,N_559,N_2660);
nand U7384 (N_7384,N_740,N_196);
or U7385 (N_7385,N_4306,N_930);
xor U7386 (N_7386,N_3876,N_737);
and U7387 (N_7387,N_4756,N_463);
or U7388 (N_7388,N_347,N_4257);
xnor U7389 (N_7389,N_4437,N_4420);
or U7390 (N_7390,N_3452,N_824);
or U7391 (N_7391,N_222,N_4310);
xnor U7392 (N_7392,N_4375,N_2297);
nor U7393 (N_7393,N_3859,N_4709);
nand U7394 (N_7394,N_3412,N_2960);
and U7395 (N_7395,N_1739,N_4867);
xor U7396 (N_7396,N_4863,N_976);
nor U7397 (N_7397,N_1354,N_3053);
and U7398 (N_7398,N_2237,N_2493);
or U7399 (N_7399,N_2714,N_276);
xnor U7400 (N_7400,N_2655,N_4189);
or U7401 (N_7401,N_2723,N_1060);
or U7402 (N_7402,N_1833,N_249);
or U7403 (N_7403,N_31,N_88);
and U7404 (N_7404,N_1170,N_4166);
xor U7405 (N_7405,N_2749,N_4029);
or U7406 (N_7406,N_70,N_1920);
nor U7407 (N_7407,N_3288,N_1849);
and U7408 (N_7408,N_3992,N_883);
or U7409 (N_7409,N_3512,N_739);
and U7410 (N_7410,N_2625,N_3523);
nand U7411 (N_7411,N_2187,N_4222);
xnor U7412 (N_7412,N_1232,N_1393);
xnor U7413 (N_7413,N_3668,N_3333);
and U7414 (N_7414,N_4315,N_311);
nand U7415 (N_7415,N_4107,N_4270);
and U7416 (N_7416,N_2202,N_4786);
and U7417 (N_7417,N_4224,N_2766);
and U7418 (N_7418,N_1016,N_3473);
and U7419 (N_7419,N_3734,N_3822);
nand U7420 (N_7420,N_459,N_3142);
nor U7421 (N_7421,N_4550,N_2832);
nand U7422 (N_7422,N_1434,N_109);
nor U7423 (N_7423,N_1212,N_2865);
and U7424 (N_7424,N_1464,N_4092);
and U7425 (N_7425,N_3458,N_3957);
nand U7426 (N_7426,N_1701,N_1564);
xnor U7427 (N_7427,N_1059,N_2492);
or U7428 (N_7428,N_113,N_864);
nand U7429 (N_7429,N_3619,N_3148);
nor U7430 (N_7430,N_4977,N_1270);
and U7431 (N_7431,N_4367,N_1819);
nor U7432 (N_7432,N_3978,N_2316);
or U7433 (N_7433,N_3052,N_430);
nand U7434 (N_7434,N_2809,N_3074);
nand U7435 (N_7435,N_4474,N_1963);
nor U7436 (N_7436,N_1898,N_445);
xor U7437 (N_7437,N_2146,N_4082);
xor U7438 (N_7438,N_2756,N_490);
or U7439 (N_7439,N_4748,N_1003);
nor U7440 (N_7440,N_4232,N_1097);
xor U7441 (N_7441,N_3188,N_1405);
and U7442 (N_7442,N_2278,N_746);
nor U7443 (N_7443,N_2565,N_1723);
nor U7444 (N_7444,N_3287,N_3425);
or U7445 (N_7445,N_582,N_3097);
nor U7446 (N_7446,N_1284,N_1904);
xnor U7447 (N_7447,N_3152,N_2722);
or U7448 (N_7448,N_446,N_2836);
nor U7449 (N_7449,N_2873,N_2381);
xnor U7450 (N_7450,N_1213,N_3020);
or U7451 (N_7451,N_3871,N_4737);
and U7452 (N_7452,N_2408,N_870);
and U7453 (N_7453,N_2369,N_1556);
xor U7454 (N_7454,N_4326,N_4951);
nand U7455 (N_7455,N_1675,N_4120);
or U7456 (N_7456,N_2232,N_720);
or U7457 (N_7457,N_3817,N_358);
nor U7458 (N_7458,N_4981,N_2274);
nand U7459 (N_7459,N_1946,N_1575);
and U7460 (N_7460,N_1993,N_216);
nand U7461 (N_7461,N_4472,N_4648);
or U7462 (N_7462,N_211,N_3149);
or U7463 (N_7463,N_2087,N_1044);
xor U7464 (N_7464,N_4623,N_2634);
xnor U7465 (N_7465,N_3550,N_1252);
or U7466 (N_7466,N_1695,N_3386);
and U7467 (N_7467,N_1983,N_3411);
and U7468 (N_7468,N_3240,N_4630);
nand U7469 (N_7469,N_854,N_2760);
nor U7470 (N_7470,N_303,N_4753);
nand U7471 (N_7471,N_4194,N_2233);
xor U7472 (N_7472,N_3637,N_4801);
xnor U7473 (N_7473,N_1406,N_40);
and U7474 (N_7474,N_1906,N_538);
nor U7475 (N_7475,N_2798,N_2027);
and U7476 (N_7476,N_1823,N_4017);
nand U7477 (N_7477,N_4926,N_91);
nand U7478 (N_7478,N_238,N_4130);
or U7479 (N_7479,N_888,N_92);
nand U7480 (N_7480,N_1634,N_2132);
and U7481 (N_7481,N_1714,N_1541);
nand U7482 (N_7482,N_3936,N_2641);
xor U7483 (N_7483,N_2308,N_3731);
xor U7484 (N_7484,N_2238,N_4023);
or U7485 (N_7485,N_1340,N_2036);
or U7486 (N_7486,N_4100,N_1944);
or U7487 (N_7487,N_2642,N_1297);
and U7488 (N_7488,N_2848,N_2057);
nand U7489 (N_7489,N_3189,N_4234);
xor U7490 (N_7490,N_2550,N_2066);
xnor U7491 (N_7491,N_3847,N_2357);
or U7492 (N_7492,N_2728,N_2826);
nand U7493 (N_7493,N_108,N_1391);
nor U7494 (N_7494,N_1957,N_2968);
nor U7495 (N_7495,N_2925,N_199);
or U7496 (N_7496,N_4652,N_3485);
xnor U7497 (N_7497,N_3557,N_4584);
and U7498 (N_7498,N_3264,N_3078);
nor U7499 (N_7499,N_1560,N_700);
nor U7500 (N_7500,N_1232,N_478);
and U7501 (N_7501,N_661,N_1128);
nor U7502 (N_7502,N_149,N_4935);
nand U7503 (N_7503,N_3862,N_1735);
nand U7504 (N_7504,N_1875,N_1027);
nor U7505 (N_7505,N_2125,N_1600);
nand U7506 (N_7506,N_2010,N_2470);
or U7507 (N_7507,N_454,N_569);
xnor U7508 (N_7508,N_4629,N_402);
nand U7509 (N_7509,N_4288,N_1990);
or U7510 (N_7510,N_4590,N_2621);
or U7511 (N_7511,N_4633,N_2186);
or U7512 (N_7512,N_2954,N_4447);
and U7513 (N_7513,N_1485,N_1500);
nand U7514 (N_7514,N_531,N_4228);
xor U7515 (N_7515,N_17,N_654);
nor U7516 (N_7516,N_4281,N_2371);
nor U7517 (N_7517,N_632,N_980);
and U7518 (N_7518,N_3023,N_4761);
xnor U7519 (N_7519,N_924,N_2972);
nand U7520 (N_7520,N_1097,N_2650);
or U7521 (N_7521,N_1027,N_318);
xnor U7522 (N_7522,N_3683,N_4524);
nor U7523 (N_7523,N_473,N_3939);
nand U7524 (N_7524,N_13,N_354);
or U7525 (N_7525,N_3978,N_2292);
nand U7526 (N_7526,N_2375,N_382);
and U7527 (N_7527,N_4516,N_3774);
and U7528 (N_7528,N_3846,N_2563);
and U7529 (N_7529,N_2184,N_3463);
nand U7530 (N_7530,N_2543,N_1807);
nor U7531 (N_7531,N_143,N_4945);
xnor U7532 (N_7532,N_336,N_4993);
xnor U7533 (N_7533,N_3748,N_1339);
or U7534 (N_7534,N_1454,N_3001);
or U7535 (N_7535,N_1427,N_4350);
and U7536 (N_7536,N_4594,N_1555);
nand U7537 (N_7537,N_3960,N_4496);
xnor U7538 (N_7538,N_4481,N_2549);
nand U7539 (N_7539,N_4074,N_305);
xor U7540 (N_7540,N_4285,N_3497);
or U7541 (N_7541,N_4402,N_3962);
or U7542 (N_7542,N_4589,N_4615);
and U7543 (N_7543,N_1900,N_1327);
or U7544 (N_7544,N_1863,N_3861);
nand U7545 (N_7545,N_3068,N_3822);
and U7546 (N_7546,N_2951,N_1516);
nand U7547 (N_7547,N_2256,N_1887);
nor U7548 (N_7548,N_4271,N_2054);
xor U7549 (N_7549,N_3910,N_100);
nand U7550 (N_7550,N_3987,N_4412);
xnor U7551 (N_7551,N_3952,N_339);
or U7552 (N_7552,N_3644,N_3134);
and U7553 (N_7553,N_4040,N_997);
and U7554 (N_7554,N_3868,N_3634);
or U7555 (N_7555,N_3672,N_4766);
and U7556 (N_7556,N_876,N_3485);
xor U7557 (N_7557,N_3955,N_3839);
and U7558 (N_7558,N_4665,N_1470);
or U7559 (N_7559,N_2073,N_898);
or U7560 (N_7560,N_3322,N_1576);
nand U7561 (N_7561,N_4562,N_1748);
and U7562 (N_7562,N_3690,N_2647);
nor U7563 (N_7563,N_567,N_1751);
and U7564 (N_7564,N_781,N_2688);
xnor U7565 (N_7565,N_4153,N_327);
nand U7566 (N_7566,N_1617,N_4057);
and U7567 (N_7567,N_4631,N_993);
and U7568 (N_7568,N_2586,N_3753);
nor U7569 (N_7569,N_137,N_402);
or U7570 (N_7570,N_2125,N_527);
nand U7571 (N_7571,N_2933,N_3761);
xnor U7572 (N_7572,N_875,N_1218);
nor U7573 (N_7573,N_4513,N_1773);
or U7574 (N_7574,N_1231,N_59);
and U7575 (N_7575,N_1504,N_1030);
and U7576 (N_7576,N_4804,N_2736);
or U7577 (N_7577,N_216,N_914);
nand U7578 (N_7578,N_2938,N_3167);
and U7579 (N_7579,N_3960,N_3133);
xnor U7580 (N_7580,N_3637,N_2955);
or U7581 (N_7581,N_170,N_767);
xor U7582 (N_7582,N_3378,N_1619);
nand U7583 (N_7583,N_2598,N_4436);
xor U7584 (N_7584,N_137,N_1650);
or U7585 (N_7585,N_3478,N_400);
nand U7586 (N_7586,N_2040,N_2112);
nand U7587 (N_7587,N_4706,N_828);
nand U7588 (N_7588,N_4630,N_2432);
and U7589 (N_7589,N_648,N_1622);
and U7590 (N_7590,N_4361,N_94);
and U7591 (N_7591,N_3995,N_3353);
nor U7592 (N_7592,N_3547,N_411);
nand U7593 (N_7593,N_608,N_3351);
xnor U7594 (N_7594,N_3139,N_1214);
xor U7595 (N_7595,N_1088,N_1663);
nor U7596 (N_7596,N_4113,N_100);
or U7597 (N_7597,N_1923,N_2352);
nor U7598 (N_7598,N_4745,N_1704);
nor U7599 (N_7599,N_2283,N_4615);
or U7600 (N_7600,N_450,N_1847);
nand U7601 (N_7601,N_3472,N_210);
nand U7602 (N_7602,N_2541,N_2928);
or U7603 (N_7603,N_528,N_2708);
or U7604 (N_7604,N_4130,N_309);
and U7605 (N_7605,N_2670,N_1896);
nand U7606 (N_7606,N_3558,N_1104);
and U7607 (N_7607,N_2655,N_3796);
or U7608 (N_7608,N_4692,N_4010);
or U7609 (N_7609,N_237,N_4980);
and U7610 (N_7610,N_1072,N_3892);
xnor U7611 (N_7611,N_3998,N_657);
and U7612 (N_7612,N_2833,N_3656);
xor U7613 (N_7613,N_4045,N_1891);
nor U7614 (N_7614,N_3786,N_4735);
nor U7615 (N_7615,N_3273,N_998);
xor U7616 (N_7616,N_3248,N_4297);
nor U7617 (N_7617,N_108,N_4384);
or U7618 (N_7618,N_4207,N_3382);
nor U7619 (N_7619,N_2695,N_93);
nor U7620 (N_7620,N_4972,N_4647);
and U7621 (N_7621,N_4969,N_309);
nand U7622 (N_7622,N_2250,N_2797);
or U7623 (N_7623,N_2071,N_2070);
nor U7624 (N_7624,N_2253,N_1014);
xor U7625 (N_7625,N_4428,N_2448);
or U7626 (N_7626,N_569,N_1727);
and U7627 (N_7627,N_3198,N_3169);
nor U7628 (N_7628,N_2603,N_3627);
or U7629 (N_7629,N_3913,N_1561);
nand U7630 (N_7630,N_2597,N_2808);
nand U7631 (N_7631,N_2468,N_865);
xor U7632 (N_7632,N_4786,N_509);
or U7633 (N_7633,N_2026,N_3829);
nand U7634 (N_7634,N_4576,N_3982);
xnor U7635 (N_7635,N_3951,N_4881);
or U7636 (N_7636,N_4646,N_1337);
xnor U7637 (N_7637,N_27,N_2115);
and U7638 (N_7638,N_3421,N_451);
and U7639 (N_7639,N_26,N_1191);
or U7640 (N_7640,N_1354,N_2594);
and U7641 (N_7641,N_4513,N_4568);
or U7642 (N_7642,N_1651,N_2605);
nand U7643 (N_7643,N_3876,N_2030);
and U7644 (N_7644,N_840,N_4843);
and U7645 (N_7645,N_3409,N_2592);
and U7646 (N_7646,N_4324,N_923);
or U7647 (N_7647,N_4776,N_1977);
xor U7648 (N_7648,N_3811,N_3355);
nor U7649 (N_7649,N_2450,N_1689);
xor U7650 (N_7650,N_1628,N_1683);
and U7651 (N_7651,N_2232,N_4073);
or U7652 (N_7652,N_1872,N_4227);
or U7653 (N_7653,N_1472,N_4751);
xor U7654 (N_7654,N_1140,N_4564);
or U7655 (N_7655,N_1432,N_2593);
or U7656 (N_7656,N_659,N_4938);
or U7657 (N_7657,N_4876,N_3802);
or U7658 (N_7658,N_1247,N_611);
nor U7659 (N_7659,N_3586,N_3170);
xnor U7660 (N_7660,N_2643,N_1436);
xnor U7661 (N_7661,N_1973,N_2963);
or U7662 (N_7662,N_1209,N_3279);
xor U7663 (N_7663,N_669,N_1703);
nor U7664 (N_7664,N_4993,N_3366);
xor U7665 (N_7665,N_4325,N_1109);
and U7666 (N_7666,N_3888,N_4274);
or U7667 (N_7667,N_2072,N_2531);
nor U7668 (N_7668,N_4654,N_3943);
and U7669 (N_7669,N_967,N_1102);
xnor U7670 (N_7670,N_1526,N_4015);
and U7671 (N_7671,N_2373,N_2039);
and U7672 (N_7672,N_3105,N_3872);
xor U7673 (N_7673,N_4277,N_3625);
nand U7674 (N_7674,N_3533,N_3328);
and U7675 (N_7675,N_3084,N_3387);
nand U7676 (N_7676,N_401,N_2223);
and U7677 (N_7677,N_2886,N_1856);
or U7678 (N_7678,N_1309,N_4112);
nand U7679 (N_7679,N_1729,N_3197);
or U7680 (N_7680,N_4373,N_253);
nor U7681 (N_7681,N_425,N_4306);
xor U7682 (N_7682,N_4255,N_305);
nor U7683 (N_7683,N_4548,N_785);
xnor U7684 (N_7684,N_1466,N_1574);
xnor U7685 (N_7685,N_3562,N_3373);
nor U7686 (N_7686,N_4174,N_4979);
or U7687 (N_7687,N_3424,N_4696);
or U7688 (N_7688,N_4594,N_40);
or U7689 (N_7689,N_3853,N_2239);
nand U7690 (N_7690,N_2773,N_4477);
nor U7691 (N_7691,N_497,N_3231);
and U7692 (N_7692,N_4190,N_292);
and U7693 (N_7693,N_1842,N_4028);
nor U7694 (N_7694,N_3126,N_390);
and U7695 (N_7695,N_427,N_4325);
nor U7696 (N_7696,N_4787,N_1366);
or U7697 (N_7697,N_4909,N_4671);
xor U7698 (N_7698,N_4567,N_3606);
nor U7699 (N_7699,N_4195,N_2082);
or U7700 (N_7700,N_1691,N_418);
or U7701 (N_7701,N_2479,N_768);
nand U7702 (N_7702,N_4942,N_92);
or U7703 (N_7703,N_2765,N_255);
nand U7704 (N_7704,N_3414,N_1395);
nor U7705 (N_7705,N_127,N_1793);
xor U7706 (N_7706,N_107,N_4742);
nor U7707 (N_7707,N_289,N_3650);
nor U7708 (N_7708,N_4738,N_2029);
nand U7709 (N_7709,N_3437,N_1304);
or U7710 (N_7710,N_4066,N_3238);
xor U7711 (N_7711,N_1589,N_4389);
nor U7712 (N_7712,N_1975,N_2034);
nor U7713 (N_7713,N_1904,N_4080);
or U7714 (N_7714,N_3630,N_457);
and U7715 (N_7715,N_954,N_3760);
xnor U7716 (N_7716,N_2383,N_4873);
xor U7717 (N_7717,N_3408,N_1630);
xnor U7718 (N_7718,N_1335,N_3548);
xor U7719 (N_7719,N_1738,N_577);
nand U7720 (N_7720,N_1505,N_4497);
and U7721 (N_7721,N_2697,N_4309);
nor U7722 (N_7722,N_3723,N_2610);
and U7723 (N_7723,N_4275,N_4013);
and U7724 (N_7724,N_1337,N_599);
nor U7725 (N_7725,N_2712,N_4472);
nor U7726 (N_7726,N_1496,N_3345);
nand U7727 (N_7727,N_3409,N_4688);
nand U7728 (N_7728,N_713,N_1821);
nor U7729 (N_7729,N_2453,N_3706);
nand U7730 (N_7730,N_808,N_1724);
xnor U7731 (N_7731,N_70,N_830);
xnor U7732 (N_7732,N_3631,N_4864);
nor U7733 (N_7733,N_3619,N_4981);
or U7734 (N_7734,N_1700,N_1512);
or U7735 (N_7735,N_1368,N_4430);
and U7736 (N_7736,N_1155,N_2200);
nand U7737 (N_7737,N_4245,N_376);
nand U7738 (N_7738,N_1753,N_2650);
and U7739 (N_7739,N_3334,N_3659);
xnor U7740 (N_7740,N_2726,N_3811);
nor U7741 (N_7741,N_2968,N_4782);
nor U7742 (N_7742,N_4068,N_3966);
nand U7743 (N_7743,N_269,N_2231);
nor U7744 (N_7744,N_1783,N_3616);
or U7745 (N_7745,N_1373,N_340);
nand U7746 (N_7746,N_2870,N_1357);
xor U7747 (N_7747,N_336,N_604);
xnor U7748 (N_7748,N_1021,N_4818);
nor U7749 (N_7749,N_4021,N_3510);
nor U7750 (N_7750,N_3340,N_218);
nor U7751 (N_7751,N_3600,N_3520);
nor U7752 (N_7752,N_3793,N_4136);
or U7753 (N_7753,N_2269,N_781);
nand U7754 (N_7754,N_4127,N_2778);
nand U7755 (N_7755,N_3815,N_3047);
or U7756 (N_7756,N_4482,N_668);
xnor U7757 (N_7757,N_4203,N_1159);
nor U7758 (N_7758,N_1200,N_4669);
and U7759 (N_7759,N_15,N_1248);
and U7760 (N_7760,N_1630,N_4325);
xnor U7761 (N_7761,N_2218,N_3074);
or U7762 (N_7762,N_2422,N_4615);
and U7763 (N_7763,N_3341,N_2666);
or U7764 (N_7764,N_2992,N_296);
and U7765 (N_7765,N_3342,N_1018);
or U7766 (N_7766,N_4354,N_3035);
nor U7767 (N_7767,N_2282,N_2387);
and U7768 (N_7768,N_3786,N_2755);
nor U7769 (N_7769,N_912,N_4370);
xor U7770 (N_7770,N_2263,N_3118);
xor U7771 (N_7771,N_4022,N_2054);
and U7772 (N_7772,N_4069,N_681);
and U7773 (N_7773,N_3852,N_1642);
xor U7774 (N_7774,N_111,N_340);
or U7775 (N_7775,N_3814,N_2089);
nand U7776 (N_7776,N_973,N_4739);
or U7777 (N_7777,N_907,N_1714);
nand U7778 (N_7778,N_4270,N_2562);
nor U7779 (N_7779,N_2359,N_1775);
nand U7780 (N_7780,N_4158,N_18);
nor U7781 (N_7781,N_2422,N_3615);
nand U7782 (N_7782,N_1921,N_4953);
xnor U7783 (N_7783,N_3727,N_4982);
nor U7784 (N_7784,N_2553,N_3563);
nor U7785 (N_7785,N_313,N_4560);
xnor U7786 (N_7786,N_3463,N_2977);
and U7787 (N_7787,N_3114,N_195);
nand U7788 (N_7788,N_158,N_4311);
and U7789 (N_7789,N_1711,N_4350);
nand U7790 (N_7790,N_1621,N_4993);
or U7791 (N_7791,N_313,N_1256);
nand U7792 (N_7792,N_4534,N_294);
nand U7793 (N_7793,N_3489,N_4571);
or U7794 (N_7794,N_956,N_2197);
or U7795 (N_7795,N_793,N_3986);
nor U7796 (N_7796,N_2843,N_2736);
nor U7797 (N_7797,N_4348,N_2034);
xor U7798 (N_7798,N_4461,N_2192);
or U7799 (N_7799,N_4241,N_3179);
and U7800 (N_7800,N_2728,N_3632);
and U7801 (N_7801,N_3072,N_2318);
and U7802 (N_7802,N_2487,N_4988);
nor U7803 (N_7803,N_2808,N_2327);
xnor U7804 (N_7804,N_1480,N_4360);
nor U7805 (N_7805,N_1755,N_360);
xnor U7806 (N_7806,N_4779,N_3281);
and U7807 (N_7807,N_1768,N_2139);
nor U7808 (N_7808,N_577,N_1931);
and U7809 (N_7809,N_1703,N_4062);
xnor U7810 (N_7810,N_2479,N_276);
nor U7811 (N_7811,N_3914,N_2582);
nor U7812 (N_7812,N_192,N_4210);
nor U7813 (N_7813,N_4099,N_1649);
nor U7814 (N_7814,N_1835,N_2529);
and U7815 (N_7815,N_3209,N_1641);
or U7816 (N_7816,N_2510,N_1290);
xnor U7817 (N_7817,N_583,N_4838);
xnor U7818 (N_7818,N_2900,N_2222);
and U7819 (N_7819,N_324,N_3521);
nand U7820 (N_7820,N_2733,N_494);
nor U7821 (N_7821,N_3882,N_1656);
nor U7822 (N_7822,N_359,N_4676);
nor U7823 (N_7823,N_1897,N_3871);
nor U7824 (N_7824,N_833,N_3489);
and U7825 (N_7825,N_866,N_3659);
nor U7826 (N_7826,N_2666,N_2898);
xor U7827 (N_7827,N_4748,N_2634);
xnor U7828 (N_7828,N_4282,N_4488);
nor U7829 (N_7829,N_2953,N_3590);
nor U7830 (N_7830,N_4913,N_54);
and U7831 (N_7831,N_3224,N_831);
xor U7832 (N_7832,N_44,N_2413);
nor U7833 (N_7833,N_4443,N_13);
nand U7834 (N_7834,N_3697,N_4891);
xor U7835 (N_7835,N_3435,N_4304);
nand U7836 (N_7836,N_2236,N_4951);
or U7837 (N_7837,N_2801,N_105);
nor U7838 (N_7838,N_1669,N_4200);
nor U7839 (N_7839,N_688,N_1760);
xnor U7840 (N_7840,N_2366,N_1780);
or U7841 (N_7841,N_434,N_3274);
nand U7842 (N_7842,N_1936,N_929);
or U7843 (N_7843,N_4633,N_4321);
nor U7844 (N_7844,N_934,N_846);
nand U7845 (N_7845,N_159,N_3788);
and U7846 (N_7846,N_2648,N_989);
and U7847 (N_7847,N_2164,N_109);
xnor U7848 (N_7848,N_1776,N_1051);
nand U7849 (N_7849,N_1215,N_1427);
nand U7850 (N_7850,N_1912,N_836);
nand U7851 (N_7851,N_1120,N_1192);
nor U7852 (N_7852,N_602,N_3724);
nor U7853 (N_7853,N_1190,N_1617);
nand U7854 (N_7854,N_1976,N_3506);
or U7855 (N_7855,N_3888,N_3294);
and U7856 (N_7856,N_2136,N_1717);
or U7857 (N_7857,N_1202,N_484);
xnor U7858 (N_7858,N_1491,N_4407);
or U7859 (N_7859,N_3019,N_4528);
and U7860 (N_7860,N_1633,N_3914);
xor U7861 (N_7861,N_149,N_4494);
nor U7862 (N_7862,N_1798,N_1315);
nand U7863 (N_7863,N_758,N_4567);
xnor U7864 (N_7864,N_190,N_3368);
nor U7865 (N_7865,N_2194,N_1081);
nand U7866 (N_7866,N_3933,N_2106);
and U7867 (N_7867,N_2162,N_1142);
and U7868 (N_7868,N_3237,N_806);
nor U7869 (N_7869,N_3070,N_3807);
xnor U7870 (N_7870,N_4511,N_1372);
or U7871 (N_7871,N_4031,N_4523);
or U7872 (N_7872,N_147,N_1805);
and U7873 (N_7873,N_4665,N_908);
or U7874 (N_7874,N_1946,N_4361);
and U7875 (N_7875,N_4832,N_2740);
nand U7876 (N_7876,N_1972,N_3591);
or U7877 (N_7877,N_1668,N_4173);
or U7878 (N_7878,N_1165,N_713);
xor U7879 (N_7879,N_4034,N_3164);
or U7880 (N_7880,N_2050,N_2038);
nand U7881 (N_7881,N_3084,N_4880);
nand U7882 (N_7882,N_2725,N_1027);
or U7883 (N_7883,N_341,N_4707);
nor U7884 (N_7884,N_3511,N_2391);
or U7885 (N_7885,N_4427,N_4991);
xor U7886 (N_7886,N_969,N_2965);
nor U7887 (N_7887,N_2703,N_4708);
and U7888 (N_7888,N_2121,N_4427);
nand U7889 (N_7889,N_1103,N_1584);
xor U7890 (N_7890,N_4638,N_4390);
nor U7891 (N_7891,N_2518,N_2913);
and U7892 (N_7892,N_1574,N_184);
or U7893 (N_7893,N_2623,N_3028);
and U7894 (N_7894,N_1600,N_653);
nand U7895 (N_7895,N_1653,N_1963);
or U7896 (N_7896,N_2091,N_4071);
nand U7897 (N_7897,N_337,N_942);
or U7898 (N_7898,N_3784,N_1398);
xor U7899 (N_7899,N_4898,N_558);
nor U7900 (N_7900,N_2233,N_3015);
or U7901 (N_7901,N_1012,N_1888);
xor U7902 (N_7902,N_4761,N_1929);
xnor U7903 (N_7903,N_455,N_1645);
xor U7904 (N_7904,N_3559,N_4244);
nand U7905 (N_7905,N_1020,N_1807);
or U7906 (N_7906,N_3323,N_960);
nor U7907 (N_7907,N_1110,N_4312);
nand U7908 (N_7908,N_1745,N_2920);
xor U7909 (N_7909,N_1344,N_4903);
nand U7910 (N_7910,N_3050,N_4444);
nand U7911 (N_7911,N_3334,N_2284);
nor U7912 (N_7912,N_4250,N_3463);
xnor U7913 (N_7913,N_1737,N_4297);
or U7914 (N_7914,N_1737,N_3343);
or U7915 (N_7915,N_743,N_1046);
nor U7916 (N_7916,N_4762,N_3333);
xor U7917 (N_7917,N_4101,N_311);
xor U7918 (N_7918,N_3755,N_2474);
xor U7919 (N_7919,N_1175,N_2067);
or U7920 (N_7920,N_3146,N_1361);
nor U7921 (N_7921,N_730,N_684);
nor U7922 (N_7922,N_4867,N_210);
nor U7923 (N_7923,N_4978,N_2847);
nor U7924 (N_7924,N_3491,N_132);
and U7925 (N_7925,N_3460,N_4429);
xor U7926 (N_7926,N_1592,N_3557);
or U7927 (N_7927,N_2251,N_475);
xor U7928 (N_7928,N_3484,N_4939);
nor U7929 (N_7929,N_2658,N_3572);
xnor U7930 (N_7930,N_907,N_2753);
nor U7931 (N_7931,N_4752,N_797);
xor U7932 (N_7932,N_4095,N_4220);
or U7933 (N_7933,N_1302,N_3660);
xor U7934 (N_7934,N_3295,N_2705);
xor U7935 (N_7935,N_351,N_2003);
nand U7936 (N_7936,N_3405,N_96);
or U7937 (N_7937,N_2391,N_1177);
or U7938 (N_7938,N_3714,N_869);
nand U7939 (N_7939,N_697,N_2657);
nand U7940 (N_7940,N_3325,N_571);
xnor U7941 (N_7941,N_83,N_4494);
or U7942 (N_7942,N_1460,N_2440);
or U7943 (N_7943,N_1992,N_16);
or U7944 (N_7944,N_3061,N_3127);
nand U7945 (N_7945,N_4048,N_870);
nor U7946 (N_7946,N_2524,N_4674);
nand U7947 (N_7947,N_2135,N_984);
xnor U7948 (N_7948,N_319,N_191);
or U7949 (N_7949,N_3946,N_530);
nor U7950 (N_7950,N_2587,N_2872);
nor U7951 (N_7951,N_823,N_2026);
or U7952 (N_7952,N_660,N_3267);
xnor U7953 (N_7953,N_3848,N_2160);
nor U7954 (N_7954,N_4365,N_1012);
nand U7955 (N_7955,N_1831,N_4663);
or U7956 (N_7956,N_4103,N_3364);
or U7957 (N_7957,N_2196,N_3476);
nor U7958 (N_7958,N_3982,N_3189);
nor U7959 (N_7959,N_2035,N_4142);
and U7960 (N_7960,N_2621,N_4264);
or U7961 (N_7961,N_1005,N_1249);
and U7962 (N_7962,N_261,N_3987);
nand U7963 (N_7963,N_3053,N_1975);
nand U7964 (N_7964,N_4202,N_2954);
or U7965 (N_7965,N_2692,N_2473);
xnor U7966 (N_7966,N_2455,N_1567);
nand U7967 (N_7967,N_4263,N_2773);
nor U7968 (N_7968,N_2435,N_595);
nor U7969 (N_7969,N_471,N_3611);
nor U7970 (N_7970,N_3704,N_2054);
nor U7971 (N_7971,N_3697,N_2938);
nand U7972 (N_7972,N_1392,N_2606);
xor U7973 (N_7973,N_449,N_4517);
or U7974 (N_7974,N_504,N_574);
nand U7975 (N_7975,N_2461,N_911);
xnor U7976 (N_7976,N_1321,N_891);
or U7977 (N_7977,N_1729,N_3314);
or U7978 (N_7978,N_3717,N_3627);
or U7979 (N_7979,N_1768,N_1195);
nand U7980 (N_7980,N_3787,N_2262);
xnor U7981 (N_7981,N_1674,N_2460);
xnor U7982 (N_7982,N_1568,N_4781);
or U7983 (N_7983,N_199,N_351);
nand U7984 (N_7984,N_482,N_533);
nand U7985 (N_7985,N_2093,N_1530);
nor U7986 (N_7986,N_881,N_3114);
or U7987 (N_7987,N_1754,N_3457);
xnor U7988 (N_7988,N_2689,N_4998);
and U7989 (N_7989,N_493,N_3896);
and U7990 (N_7990,N_3852,N_1391);
xnor U7991 (N_7991,N_55,N_4401);
xnor U7992 (N_7992,N_1544,N_2541);
or U7993 (N_7993,N_3612,N_2909);
xnor U7994 (N_7994,N_1226,N_433);
xnor U7995 (N_7995,N_1184,N_670);
xnor U7996 (N_7996,N_187,N_3942);
or U7997 (N_7997,N_4797,N_2411);
and U7998 (N_7998,N_4560,N_891);
or U7999 (N_7999,N_4920,N_111);
and U8000 (N_8000,N_2917,N_1100);
nand U8001 (N_8001,N_1659,N_750);
nand U8002 (N_8002,N_2826,N_3785);
xnor U8003 (N_8003,N_4478,N_1253);
nor U8004 (N_8004,N_916,N_291);
nand U8005 (N_8005,N_4325,N_2043);
or U8006 (N_8006,N_4154,N_4194);
nor U8007 (N_8007,N_269,N_4067);
and U8008 (N_8008,N_2843,N_3773);
nand U8009 (N_8009,N_3226,N_2653);
xnor U8010 (N_8010,N_3328,N_4156);
and U8011 (N_8011,N_1502,N_2947);
and U8012 (N_8012,N_2607,N_4565);
nand U8013 (N_8013,N_2072,N_2387);
nor U8014 (N_8014,N_3161,N_1841);
nor U8015 (N_8015,N_3199,N_1884);
xnor U8016 (N_8016,N_2067,N_2277);
or U8017 (N_8017,N_2929,N_1018);
xor U8018 (N_8018,N_2954,N_4427);
xor U8019 (N_8019,N_4964,N_398);
and U8020 (N_8020,N_3385,N_4484);
nand U8021 (N_8021,N_1860,N_2249);
nor U8022 (N_8022,N_2434,N_3657);
nor U8023 (N_8023,N_389,N_2790);
or U8024 (N_8024,N_1822,N_4880);
or U8025 (N_8025,N_2945,N_700);
nor U8026 (N_8026,N_3445,N_3651);
nand U8027 (N_8027,N_4940,N_486);
and U8028 (N_8028,N_1846,N_4107);
xor U8029 (N_8029,N_3733,N_4646);
or U8030 (N_8030,N_929,N_3105);
and U8031 (N_8031,N_4424,N_1466);
and U8032 (N_8032,N_2303,N_1456);
xor U8033 (N_8033,N_3009,N_3077);
nand U8034 (N_8034,N_1540,N_3521);
xor U8035 (N_8035,N_2146,N_1522);
nand U8036 (N_8036,N_4546,N_125);
nand U8037 (N_8037,N_1252,N_340);
nor U8038 (N_8038,N_472,N_1976);
and U8039 (N_8039,N_1050,N_1042);
or U8040 (N_8040,N_4845,N_205);
and U8041 (N_8041,N_2471,N_2990);
xnor U8042 (N_8042,N_3902,N_3655);
or U8043 (N_8043,N_1013,N_3134);
and U8044 (N_8044,N_3185,N_372);
xnor U8045 (N_8045,N_1611,N_4);
nor U8046 (N_8046,N_1847,N_478);
or U8047 (N_8047,N_3636,N_4166);
and U8048 (N_8048,N_602,N_3982);
or U8049 (N_8049,N_3054,N_3424);
nand U8050 (N_8050,N_2388,N_335);
nor U8051 (N_8051,N_4220,N_2723);
nor U8052 (N_8052,N_1804,N_3438);
or U8053 (N_8053,N_3400,N_2759);
nand U8054 (N_8054,N_2710,N_3932);
or U8055 (N_8055,N_4894,N_3344);
xor U8056 (N_8056,N_121,N_2074);
xnor U8057 (N_8057,N_4573,N_2966);
and U8058 (N_8058,N_3210,N_3);
nand U8059 (N_8059,N_1465,N_4166);
or U8060 (N_8060,N_1482,N_4756);
nor U8061 (N_8061,N_1131,N_3569);
nor U8062 (N_8062,N_3044,N_2098);
or U8063 (N_8063,N_2140,N_2136);
nand U8064 (N_8064,N_3854,N_1823);
and U8065 (N_8065,N_1025,N_594);
xor U8066 (N_8066,N_2736,N_4412);
or U8067 (N_8067,N_801,N_1706);
nand U8068 (N_8068,N_747,N_695);
nor U8069 (N_8069,N_2007,N_1510);
nand U8070 (N_8070,N_435,N_4946);
or U8071 (N_8071,N_2921,N_3104);
and U8072 (N_8072,N_3954,N_1390);
and U8073 (N_8073,N_1212,N_1244);
xor U8074 (N_8074,N_3977,N_3753);
or U8075 (N_8075,N_2200,N_4299);
nor U8076 (N_8076,N_1263,N_855);
xor U8077 (N_8077,N_1905,N_2020);
or U8078 (N_8078,N_1047,N_1853);
or U8079 (N_8079,N_1248,N_4456);
and U8080 (N_8080,N_3755,N_3334);
or U8081 (N_8081,N_1796,N_4521);
xor U8082 (N_8082,N_4320,N_1827);
xnor U8083 (N_8083,N_2854,N_4024);
xor U8084 (N_8084,N_3460,N_625);
nand U8085 (N_8085,N_1576,N_3671);
nor U8086 (N_8086,N_1616,N_1845);
xnor U8087 (N_8087,N_80,N_242);
nand U8088 (N_8088,N_2423,N_673);
nand U8089 (N_8089,N_3546,N_1946);
nor U8090 (N_8090,N_3074,N_2642);
xor U8091 (N_8091,N_1896,N_3218);
or U8092 (N_8092,N_3841,N_1449);
and U8093 (N_8093,N_3908,N_1959);
nor U8094 (N_8094,N_775,N_1916);
xor U8095 (N_8095,N_111,N_3888);
and U8096 (N_8096,N_4188,N_553);
or U8097 (N_8097,N_2162,N_3013);
or U8098 (N_8098,N_212,N_2282);
nor U8099 (N_8099,N_4035,N_3891);
and U8100 (N_8100,N_3762,N_3800);
xor U8101 (N_8101,N_2794,N_3900);
and U8102 (N_8102,N_562,N_4576);
nor U8103 (N_8103,N_3414,N_954);
nor U8104 (N_8104,N_1760,N_2167);
and U8105 (N_8105,N_2670,N_1947);
xor U8106 (N_8106,N_969,N_3507);
nor U8107 (N_8107,N_4534,N_11);
and U8108 (N_8108,N_4042,N_981);
xnor U8109 (N_8109,N_3794,N_4566);
nand U8110 (N_8110,N_4675,N_675);
or U8111 (N_8111,N_4513,N_1599);
or U8112 (N_8112,N_3307,N_1040);
nand U8113 (N_8113,N_863,N_607);
nor U8114 (N_8114,N_2786,N_2407);
nand U8115 (N_8115,N_2793,N_4014);
nor U8116 (N_8116,N_3832,N_499);
nand U8117 (N_8117,N_3906,N_1354);
or U8118 (N_8118,N_4606,N_3910);
nand U8119 (N_8119,N_3510,N_1223);
nand U8120 (N_8120,N_4088,N_4744);
nand U8121 (N_8121,N_1790,N_589);
nand U8122 (N_8122,N_4408,N_4316);
or U8123 (N_8123,N_2056,N_1565);
nor U8124 (N_8124,N_3295,N_404);
nand U8125 (N_8125,N_2932,N_4551);
or U8126 (N_8126,N_2669,N_2052);
and U8127 (N_8127,N_2839,N_644);
xor U8128 (N_8128,N_1858,N_4294);
and U8129 (N_8129,N_4460,N_236);
nand U8130 (N_8130,N_4135,N_3965);
and U8131 (N_8131,N_2373,N_510);
nor U8132 (N_8132,N_964,N_3601);
and U8133 (N_8133,N_1328,N_2743);
nand U8134 (N_8134,N_122,N_2174);
and U8135 (N_8135,N_4633,N_2416);
nand U8136 (N_8136,N_3703,N_975);
and U8137 (N_8137,N_4495,N_4736);
xnor U8138 (N_8138,N_636,N_3974);
nor U8139 (N_8139,N_2388,N_2641);
nor U8140 (N_8140,N_3988,N_931);
and U8141 (N_8141,N_490,N_115);
and U8142 (N_8142,N_4380,N_2113);
nor U8143 (N_8143,N_4444,N_3912);
xor U8144 (N_8144,N_3894,N_2478);
and U8145 (N_8145,N_4997,N_4545);
nor U8146 (N_8146,N_2482,N_2053);
nand U8147 (N_8147,N_2188,N_2479);
or U8148 (N_8148,N_2808,N_1261);
nand U8149 (N_8149,N_3144,N_2168);
and U8150 (N_8150,N_4608,N_524);
or U8151 (N_8151,N_3831,N_3459);
xnor U8152 (N_8152,N_2321,N_3816);
xnor U8153 (N_8153,N_337,N_4334);
nand U8154 (N_8154,N_335,N_3998);
nor U8155 (N_8155,N_1417,N_267);
or U8156 (N_8156,N_1108,N_4905);
nor U8157 (N_8157,N_285,N_1374);
xor U8158 (N_8158,N_3139,N_3433);
nor U8159 (N_8159,N_3154,N_991);
or U8160 (N_8160,N_2148,N_4393);
nand U8161 (N_8161,N_2511,N_1229);
and U8162 (N_8162,N_4384,N_822);
nand U8163 (N_8163,N_1693,N_1996);
nor U8164 (N_8164,N_3614,N_4083);
or U8165 (N_8165,N_4286,N_2109);
xnor U8166 (N_8166,N_2000,N_4234);
nor U8167 (N_8167,N_1183,N_3085);
or U8168 (N_8168,N_1006,N_3800);
and U8169 (N_8169,N_2378,N_983);
and U8170 (N_8170,N_4798,N_205);
and U8171 (N_8171,N_3878,N_4931);
and U8172 (N_8172,N_4824,N_1029);
xnor U8173 (N_8173,N_585,N_2206);
and U8174 (N_8174,N_120,N_846);
nor U8175 (N_8175,N_3813,N_1766);
nand U8176 (N_8176,N_2702,N_30);
xnor U8177 (N_8177,N_3789,N_2798);
nand U8178 (N_8178,N_3621,N_978);
or U8179 (N_8179,N_3528,N_797);
nand U8180 (N_8180,N_4553,N_2299);
or U8181 (N_8181,N_2830,N_3786);
nor U8182 (N_8182,N_3185,N_2045);
or U8183 (N_8183,N_3052,N_1005);
nor U8184 (N_8184,N_3559,N_2949);
or U8185 (N_8185,N_3791,N_820);
xor U8186 (N_8186,N_1090,N_593);
or U8187 (N_8187,N_2019,N_4245);
nand U8188 (N_8188,N_3447,N_2182);
and U8189 (N_8189,N_611,N_914);
xnor U8190 (N_8190,N_4357,N_2737);
nand U8191 (N_8191,N_3411,N_3554);
nand U8192 (N_8192,N_793,N_1285);
or U8193 (N_8193,N_1536,N_1989);
xnor U8194 (N_8194,N_1468,N_957);
nand U8195 (N_8195,N_136,N_4055);
nand U8196 (N_8196,N_3848,N_2695);
or U8197 (N_8197,N_3908,N_183);
or U8198 (N_8198,N_1139,N_1925);
xnor U8199 (N_8199,N_108,N_701);
nor U8200 (N_8200,N_4572,N_3426);
nand U8201 (N_8201,N_891,N_4171);
nand U8202 (N_8202,N_1521,N_3781);
nor U8203 (N_8203,N_2760,N_2901);
and U8204 (N_8204,N_854,N_791);
or U8205 (N_8205,N_231,N_1454);
nand U8206 (N_8206,N_1233,N_4568);
or U8207 (N_8207,N_2820,N_109);
nor U8208 (N_8208,N_3644,N_3817);
and U8209 (N_8209,N_1742,N_3428);
and U8210 (N_8210,N_2269,N_3802);
or U8211 (N_8211,N_981,N_3927);
or U8212 (N_8212,N_489,N_2146);
and U8213 (N_8213,N_1643,N_1162);
and U8214 (N_8214,N_3425,N_2022);
nand U8215 (N_8215,N_3545,N_2016);
nor U8216 (N_8216,N_4734,N_96);
xor U8217 (N_8217,N_1136,N_80);
and U8218 (N_8218,N_3628,N_1595);
nor U8219 (N_8219,N_1007,N_4461);
xor U8220 (N_8220,N_1500,N_4673);
or U8221 (N_8221,N_3314,N_4255);
and U8222 (N_8222,N_4099,N_2664);
nor U8223 (N_8223,N_3233,N_950);
or U8224 (N_8224,N_2787,N_4983);
nand U8225 (N_8225,N_4029,N_44);
or U8226 (N_8226,N_3605,N_2506);
xor U8227 (N_8227,N_808,N_1601);
xnor U8228 (N_8228,N_3969,N_3158);
nor U8229 (N_8229,N_2879,N_3747);
nor U8230 (N_8230,N_4520,N_1055);
nand U8231 (N_8231,N_1887,N_3062);
or U8232 (N_8232,N_749,N_2049);
xor U8233 (N_8233,N_3993,N_1530);
or U8234 (N_8234,N_2102,N_3933);
nand U8235 (N_8235,N_501,N_2319);
nor U8236 (N_8236,N_1438,N_555);
nor U8237 (N_8237,N_2776,N_2772);
xnor U8238 (N_8238,N_3373,N_3405);
nand U8239 (N_8239,N_4316,N_1934);
nor U8240 (N_8240,N_4346,N_484);
or U8241 (N_8241,N_4129,N_1737);
and U8242 (N_8242,N_585,N_1025);
nand U8243 (N_8243,N_4295,N_1304);
xor U8244 (N_8244,N_2575,N_2);
or U8245 (N_8245,N_2195,N_3837);
xnor U8246 (N_8246,N_3423,N_1546);
nand U8247 (N_8247,N_3448,N_2764);
or U8248 (N_8248,N_3090,N_1354);
and U8249 (N_8249,N_3497,N_3663);
nor U8250 (N_8250,N_98,N_4789);
nand U8251 (N_8251,N_957,N_369);
nor U8252 (N_8252,N_1195,N_1096);
and U8253 (N_8253,N_1145,N_1567);
nor U8254 (N_8254,N_1370,N_2991);
nor U8255 (N_8255,N_3656,N_1884);
nand U8256 (N_8256,N_3244,N_3901);
or U8257 (N_8257,N_2198,N_1887);
and U8258 (N_8258,N_3209,N_3925);
xor U8259 (N_8259,N_3914,N_3992);
or U8260 (N_8260,N_4649,N_4492);
or U8261 (N_8261,N_2818,N_1521);
and U8262 (N_8262,N_1390,N_4108);
xnor U8263 (N_8263,N_1934,N_2738);
and U8264 (N_8264,N_4575,N_2160);
and U8265 (N_8265,N_1042,N_2498);
and U8266 (N_8266,N_4875,N_3908);
or U8267 (N_8267,N_4817,N_1129);
xnor U8268 (N_8268,N_3874,N_1607);
and U8269 (N_8269,N_2899,N_1282);
nand U8270 (N_8270,N_826,N_1178);
xor U8271 (N_8271,N_2471,N_1083);
nor U8272 (N_8272,N_1715,N_1714);
or U8273 (N_8273,N_4105,N_365);
and U8274 (N_8274,N_2398,N_1819);
nor U8275 (N_8275,N_4114,N_1555);
nor U8276 (N_8276,N_4635,N_1758);
and U8277 (N_8277,N_4261,N_1736);
and U8278 (N_8278,N_3580,N_4433);
or U8279 (N_8279,N_3070,N_3861);
xnor U8280 (N_8280,N_976,N_3254);
nor U8281 (N_8281,N_2817,N_397);
xnor U8282 (N_8282,N_3942,N_1794);
xor U8283 (N_8283,N_1060,N_1099);
xnor U8284 (N_8284,N_2823,N_3849);
and U8285 (N_8285,N_2156,N_3604);
nor U8286 (N_8286,N_1812,N_4599);
xor U8287 (N_8287,N_2140,N_4893);
xnor U8288 (N_8288,N_2887,N_4023);
and U8289 (N_8289,N_4807,N_1598);
nand U8290 (N_8290,N_1437,N_3897);
nand U8291 (N_8291,N_4645,N_4803);
xnor U8292 (N_8292,N_4158,N_3429);
nand U8293 (N_8293,N_2155,N_1883);
nor U8294 (N_8294,N_2100,N_4600);
nand U8295 (N_8295,N_2966,N_3111);
xor U8296 (N_8296,N_4202,N_142);
nor U8297 (N_8297,N_2363,N_649);
xor U8298 (N_8298,N_4257,N_807);
xnor U8299 (N_8299,N_2637,N_4900);
and U8300 (N_8300,N_1265,N_1495);
nand U8301 (N_8301,N_1127,N_4597);
nor U8302 (N_8302,N_2004,N_1950);
xnor U8303 (N_8303,N_1645,N_4034);
nor U8304 (N_8304,N_4637,N_3853);
or U8305 (N_8305,N_4716,N_4674);
and U8306 (N_8306,N_381,N_3344);
nand U8307 (N_8307,N_1753,N_1836);
nand U8308 (N_8308,N_2474,N_4778);
nor U8309 (N_8309,N_942,N_2901);
and U8310 (N_8310,N_1919,N_3830);
or U8311 (N_8311,N_3165,N_592);
or U8312 (N_8312,N_4006,N_3573);
nand U8313 (N_8313,N_623,N_2610);
and U8314 (N_8314,N_1128,N_323);
or U8315 (N_8315,N_4794,N_3407);
and U8316 (N_8316,N_4108,N_4244);
or U8317 (N_8317,N_4842,N_4230);
xor U8318 (N_8318,N_1097,N_948);
and U8319 (N_8319,N_3514,N_736);
or U8320 (N_8320,N_1145,N_2434);
and U8321 (N_8321,N_2781,N_3608);
nand U8322 (N_8322,N_84,N_2622);
or U8323 (N_8323,N_4053,N_4557);
xor U8324 (N_8324,N_478,N_3443);
nand U8325 (N_8325,N_1598,N_736);
xnor U8326 (N_8326,N_1000,N_4725);
nor U8327 (N_8327,N_767,N_2005);
or U8328 (N_8328,N_1497,N_4102);
and U8329 (N_8329,N_4192,N_4751);
nor U8330 (N_8330,N_4946,N_2510);
and U8331 (N_8331,N_713,N_3154);
nor U8332 (N_8332,N_1892,N_4213);
or U8333 (N_8333,N_583,N_3627);
and U8334 (N_8334,N_3295,N_2226);
nor U8335 (N_8335,N_2772,N_313);
xor U8336 (N_8336,N_1435,N_4736);
and U8337 (N_8337,N_2701,N_1170);
or U8338 (N_8338,N_1308,N_527);
and U8339 (N_8339,N_2303,N_3533);
nor U8340 (N_8340,N_4870,N_4369);
or U8341 (N_8341,N_2220,N_687);
xor U8342 (N_8342,N_288,N_1862);
or U8343 (N_8343,N_3338,N_679);
nor U8344 (N_8344,N_275,N_4958);
nand U8345 (N_8345,N_987,N_4320);
or U8346 (N_8346,N_3662,N_3207);
nand U8347 (N_8347,N_311,N_555);
and U8348 (N_8348,N_518,N_2111);
nor U8349 (N_8349,N_3629,N_53);
nand U8350 (N_8350,N_568,N_558);
nor U8351 (N_8351,N_4851,N_4914);
or U8352 (N_8352,N_2521,N_3169);
or U8353 (N_8353,N_2932,N_15);
xor U8354 (N_8354,N_2021,N_860);
nor U8355 (N_8355,N_3099,N_126);
or U8356 (N_8356,N_4341,N_4629);
or U8357 (N_8357,N_78,N_3652);
and U8358 (N_8358,N_2782,N_4673);
and U8359 (N_8359,N_4033,N_1356);
and U8360 (N_8360,N_2029,N_4538);
or U8361 (N_8361,N_1331,N_709);
and U8362 (N_8362,N_203,N_4486);
nor U8363 (N_8363,N_2855,N_4095);
or U8364 (N_8364,N_3843,N_2240);
nand U8365 (N_8365,N_4577,N_4068);
and U8366 (N_8366,N_308,N_4102);
or U8367 (N_8367,N_3258,N_1239);
nor U8368 (N_8368,N_4087,N_775);
or U8369 (N_8369,N_630,N_4415);
or U8370 (N_8370,N_2970,N_884);
nand U8371 (N_8371,N_379,N_98);
or U8372 (N_8372,N_1418,N_3432);
nand U8373 (N_8373,N_766,N_874);
nor U8374 (N_8374,N_4504,N_1412);
nor U8375 (N_8375,N_4272,N_4145);
or U8376 (N_8376,N_2323,N_4809);
nand U8377 (N_8377,N_3695,N_549);
xor U8378 (N_8378,N_1106,N_1251);
nor U8379 (N_8379,N_4226,N_681);
xor U8380 (N_8380,N_2304,N_367);
nand U8381 (N_8381,N_4134,N_2616);
nor U8382 (N_8382,N_4649,N_2666);
or U8383 (N_8383,N_3555,N_699);
or U8384 (N_8384,N_2009,N_3797);
nor U8385 (N_8385,N_194,N_1278);
xnor U8386 (N_8386,N_4291,N_86);
nor U8387 (N_8387,N_1841,N_203);
xor U8388 (N_8388,N_3961,N_2951);
and U8389 (N_8389,N_2105,N_1496);
xor U8390 (N_8390,N_944,N_4573);
or U8391 (N_8391,N_403,N_4709);
and U8392 (N_8392,N_1337,N_53);
xor U8393 (N_8393,N_711,N_4121);
nand U8394 (N_8394,N_2920,N_2703);
or U8395 (N_8395,N_1662,N_4218);
or U8396 (N_8396,N_3840,N_549);
nor U8397 (N_8397,N_2443,N_4193);
or U8398 (N_8398,N_2459,N_854);
nand U8399 (N_8399,N_1920,N_4899);
nand U8400 (N_8400,N_1695,N_939);
nand U8401 (N_8401,N_1101,N_1056);
or U8402 (N_8402,N_4830,N_2552);
xnor U8403 (N_8403,N_2985,N_317);
nand U8404 (N_8404,N_4153,N_158);
or U8405 (N_8405,N_4100,N_4314);
nor U8406 (N_8406,N_1672,N_3712);
xnor U8407 (N_8407,N_2139,N_3098);
xor U8408 (N_8408,N_2628,N_3002);
or U8409 (N_8409,N_4035,N_1028);
xor U8410 (N_8410,N_217,N_931);
and U8411 (N_8411,N_1777,N_1799);
xnor U8412 (N_8412,N_3031,N_83);
nand U8413 (N_8413,N_498,N_2619);
or U8414 (N_8414,N_1942,N_3296);
and U8415 (N_8415,N_3869,N_4647);
nand U8416 (N_8416,N_1759,N_2351);
xnor U8417 (N_8417,N_4794,N_4393);
and U8418 (N_8418,N_3443,N_3862);
nand U8419 (N_8419,N_3030,N_4082);
or U8420 (N_8420,N_2779,N_3255);
or U8421 (N_8421,N_1031,N_2986);
and U8422 (N_8422,N_2870,N_2008);
nand U8423 (N_8423,N_4576,N_3959);
nor U8424 (N_8424,N_3894,N_117);
or U8425 (N_8425,N_1609,N_4672);
xnor U8426 (N_8426,N_4813,N_3313);
xor U8427 (N_8427,N_3009,N_4228);
or U8428 (N_8428,N_4136,N_3648);
nor U8429 (N_8429,N_2106,N_590);
and U8430 (N_8430,N_2883,N_4649);
and U8431 (N_8431,N_1121,N_4302);
nand U8432 (N_8432,N_1942,N_4273);
or U8433 (N_8433,N_3546,N_804);
nand U8434 (N_8434,N_2758,N_3250);
or U8435 (N_8435,N_2095,N_4537);
nand U8436 (N_8436,N_1183,N_4708);
nand U8437 (N_8437,N_3948,N_3123);
nor U8438 (N_8438,N_2238,N_200);
xor U8439 (N_8439,N_3322,N_4769);
or U8440 (N_8440,N_2872,N_2481);
nand U8441 (N_8441,N_453,N_3643);
xor U8442 (N_8442,N_4311,N_3519);
nand U8443 (N_8443,N_2654,N_1899);
or U8444 (N_8444,N_4821,N_629);
nand U8445 (N_8445,N_4845,N_3629);
nor U8446 (N_8446,N_71,N_3653);
nand U8447 (N_8447,N_2995,N_114);
or U8448 (N_8448,N_633,N_4179);
or U8449 (N_8449,N_2231,N_2946);
nor U8450 (N_8450,N_1665,N_3328);
nor U8451 (N_8451,N_358,N_3577);
and U8452 (N_8452,N_2330,N_766);
xnor U8453 (N_8453,N_4185,N_4286);
nor U8454 (N_8454,N_4661,N_3875);
xnor U8455 (N_8455,N_2392,N_3391);
nand U8456 (N_8456,N_3482,N_4783);
and U8457 (N_8457,N_1925,N_971);
and U8458 (N_8458,N_1235,N_3731);
nand U8459 (N_8459,N_4171,N_3992);
and U8460 (N_8460,N_4673,N_1863);
nor U8461 (N_8461,N_737,N_686);
nor U8462 (N_8462,N_1677,N_4545);
or U8463 (N_8463,N_211,N_800);
xnor U8464 (N_8464,N_859,N_3746);
nand U8465 (N_8465,N_225,N_832);
nand U8466 (N_8466,N_2210,N_2310);
and U8467 (N_8467,N_663,N_790);
nor U8468 (N_8468,N_3661,N_4488);
xnor U8469 (N_8469,N_2271,N_1946);
nand U8470 (N_8470,N_2581,N_3824);
or U8471 (N_8471,N_777,N_1251);
or U8472 (N_8472,N_1655,N_4189);
or U8473 (N_8473,N_3457,N_613);
xor U8474 (N_8474,N_1977,N_4027);
nor U8475 (N_8475,N_2551,N_3111);
nand U8476 (N_8476,N_4273,N_4572);
nand U8477 (N_8477,N_3859,N_2931);
and U8478 (N_8478,N_576,N_1004);
nand U8479 (N_8479,N_1064,N_3912);
or U8480 (N_8480,N_3491,N_2345);
xor U8481 (N_8481,N_3438,N_1027);
nand U8482 (N_8482,N_935,N_2208);
or U8483 (N_8483,N_3345,N_1175);
xor U8484 (N_8484,N_2278,N_578);
nand U8485 (N_8485,N_3524,N_2714);
or U8486 (N_8486,N_1198,N_2286);
nand U8487 (N_8487,N_2737,N_227);
and U8488 (N_8488,N_4809,N_2873);
nor U8489 (N_8489,N_2648,N_2571);
nor U8490 (N_8490,N_1808,N_4462);
nand U8491 (N_8491,N_3676,N_31);
and U8492 (N_8492,N_3308,N_525);
nor U8493 (N_8493,N_655,N_160);
nor U8494 (N_8494,N_4478,N_1137);
xnor U8495 (N_8495,N_2551,N_2097);
and U8496 (N_8496,N_1322,N_2639);
or U8497 (N_8497,N_1172,N_4504);
and U8498 (N_8498,N_2099,N_4609);
nor U8499 (N_8499,N_2412,N_3466);
nor U8500 (N_8500,N_3970,N_4661);
nor U8501 (N_8501,N_4315,N_1727);
xor U8502 (N_8502,N_4905,N_2297);
xor U8503 (N_8503,N_4339,N_1144);
or U8504 (N_8504,N_4307,N_1897);
xnor U8505 (N_8505,N_4655,N_3241);
xnor U8506 (N_8506,N_2488,N_1280);
and U8507 (N_8507,N_2477,N_4881);
nand U8508 (N_8508,N_1576,N_1710);
or U8509 (N_8509,N_4843,N_1057);
or U8510 (N_8510,N_4271,N_2830);
and U8511 (N_8511,N_1645,N_969);
and U8512 (N_8512,N_24,N_841);
xor U8513 (N_8513,N_2486,N_2098);
or U8514 (N_8514,N_70,N_3251);
xor U8515 (N_8515,N_2122,N_4588);
nand U8516 (N_8516,N_416,N_2037);
or U8517 (N_8517,N_4732,N_3986);
nand U8518 (N_8518,N_2683,N_1812);
nand U8519 (N_8519,N_1236,N_1427);
and U8520 (N_8520,N_3777,N_780);
and U8521 (N_8521,N_3963,N_2298);
nand U8522 (N_8522,N_3946,N_1134);
and U8523 (N_8523,N_4791,N_3780);
and U8524 (N_8524,N_4491,N_1404);
xnor U8525 (N_8525,N_3284,N_1411);
and U8526 (N_8526,N_3667,N_342);
or U8527 (N_8527,N_2179,N_3567);
and U8528 (N_8528,N_1873,N_3940);
nor U8529 (N_8529,N_1188,N_384);
nand U8530 (N_8530,N_4908,N_4444);
nand U8531 (N_8531,N_1775,N_3771);
nand U8532 (N_8532,N_3999,N_1752);
or U8533 (N_8533,N_910,N_2818);
or U8534 (N_8534,N_239,N_1152);
or U8535 (N_8535,N_3775,N_611);
and U8536 (N_8536,N_2568,N_210);
xor U8537 (N_8537,N_3061,N_1548);
xnor U8538 (N_8538,N_1244,N_658);
and U8539 (N_8539,N_1663,N_2962);
nor U8540 (N_8540,N_3850,N_1255);
or U8541 (N_8541,N_3833,N_1270);
nor U8542 (N_8542,N_4682,N_1724);
and U8543 (N_8543,N_482,N_4273);
nand U8544 (N_8544,N_2962,N_4004);
and U8545 (N_8545,N_1669,N_2753);
nand U8546 (N_8546,N_4766,N_3576);
xor U8547 (N_8547,N_3923,N_1136);
nand U8548 (N_8548,N_4299,N_4219);
xor U8549 (N_8549,N_3092,N_1734);
xnor U8550 (N_8550,N_4034,N_2231);
or U8551 (N_8551,N_1334,N_3709);
nor U8552 (N_8552,N_1560,N_4832);
or U8553 (N_8553,N_511,N_1856);
or U8554 (N_8554,N_1360,N_4229);
nor U8555 (N_8555,N_2640,N_3100);
or U8556 (N_8556,N_3086,N_1531);
and U8557 (N_8557,N_4551,N_953);
xnor U8558 (N_8558,N_4992,N_710);
nor U8559 (N_8559,N_938,N_277);
xor U8560 (N_8560,N_4656,N_4507);
and U8561 (N_8561,N_838,N_331);
nor U8562 (N_8562,N_4109,N_2144);
and U8563 (N_8563,N_3175,N_1533);
nand U8564 (N_8564,N_3172,N_2682);
nand U8565 (N_8565,N_1742,N_114);
xor U8566 (N_8566,N_2571,N_4555);
nor U8567 (N_8567,N_2614,N_4448);
or U8568 (N_8568,N_3381,N_2312);
nand U8569 (N_8569,N_571,N_1813);
xnor U8570 (N_8570,N_1449,N_1411);
and U8571 (N_8571,N_903,N_589);
xor U8572 (N_8572,N_3284,N_3328);
xor U8573 (N_8573,N_1765,N_397);
nand U8574 (N_8574,N_158,N_3920);
nand U8575 (N_8575,N_900,N_2434);
or U8576 (N_8576,N_4164,N_3824);
xor U8577 (N_8577,N_1218,N_988);
xnor U8578 (N_8578,N_242,N_3255);
nand U8579 (N_8579,N_315,N_385);
nand U8580 (N_8580,N_3892,N_4987);
or U8581 (N_8581,N_3257,N_1066);
nor U8582 (N_8582,N_650,N_3853);
nand U8583 (N_8583,N_1285,N_1168);
and U8584 (N_8584,N_3522,N_1779);
nor U8585 (N_8585,N_1900,N_939);
nand U8586 (N_8586,N_1521,N_256);
nor U8587 (N_8587,N_4639,N_3914);
xnor U8588 (N_8588,N_4279,N_1289);
or U8589 (N_8589,N_4374,N_4077);
or U8590 (N_8590,N_1646,N_1056);
and U8591 (N_8591,N_318,N_4366);
or U8592 (N_8592,N_1532,N_1557);
nor U8593 (N_8593,N_3285,N_3739);
and U8594 (N_8594,N_3819,N_2603);
xor U8595 (N_8595,N_3056,N_2125);
nand U8596 (N_8596,N_2037,N_1464);
or U8597 (N_8597,N_4671,N_305);
and U8598 (N_8598,N_3104,N_2472);
nor U8599 (N_8599,N_2340,N_59);
nand U8600 (N_8600,N_2784,N_3471);
and U8601 (N_8601,N_1772,N_250);
nor U8602 (N_8602,N_3472,N_2057);
or U8603 (N_8603,N_1516,N_1742);
or U8604 (N_8604,N_4720,N_4304);
and U8605 (N_8605,N_1371,N_1958);
nand U8606 (N_8606,N_1181,N_2467);
xor U8607 (N_8607,N_4822,N_3749);
nand U8608 (N_8608,N_4744,N_298);
or U8609 (N_8609,N_4177,N_3010);
xnor U8610 (N_8610,N_3089,N_2758);
nor U8611 (N_8611,N_4072,N_3489);
nand U8612 (N_8612,N_939,N_420);
nand U8613 (N_8613,N_982,N_2746);
or U8614 (N_8614,N_3036,N_194);
and U8615 (N_8615,N_4034,N_730);
xor U8616 (N_8616,N_3487,N_2100);
and U8617 (N_8617,N_392,N_2478);
nand U8618 (N_8618,N_1412,N_553);
xor U8619 (N_8619,N_169,N_2037);
and U8620 (N_8620,N_1030,N_1719);
and U8621 (N_8621,N_1616,N_3685);
and U8622 (N_8622,N_1248,N_1193);
or U8623 (N_8623,N_772,N_59);
and U8624 (N_8624,N_4300,N_689);
nand U8625 (N_8625,N_297,N_3823);
nor U8626 (N_8626,N_1516,N_754);
nand U8627 (N_8627,N_918,N_748);
or U8628 (N_8628,N_518,N_4608);
nand U8629 (N_8629,N_262,N_3381);
nor U8630 (N_8630,N_579,N_1163);
nand U8631 (N_8631,N_4485,N_4872);
or U8632 (N_8632,N_2132,N_2902);
nor U8633 (N_8633,N_3630,N_2627);
nand U8634 (N_8634,N_303,N_2107);
xor U8635 (N_8635,N_211,N_1427);
or U8636 (N_8636,N_2784,N_4354);
xor U8637 (N_8637,N_4230,N_701);
nor U8638 (N_8638,N_4826,N_2873);
xor U8639 (N_8639,N_3283,N_4937);
or U8640 (N_8640,N_1934,N_2251);
nor U8641 (N_8641,N_715,N_4475);
and U8642 (N_8642,N_4885,N_247);
nor U8643 (N_8643,N_1072,N_4739);
nor U8644 (N_8644,N_1595,N_215);
nor U8645 (N_8645,N_711,N_3740);
and U8646 (N_8646,N_3889,N_273);
or U8647 (N_8647,N_3861,N_3621);
nand U8648 (N_8648,N_2026,N_74);
nand U8649 (N_8649,N_4557,N_669);
or U8650 (N_8650,N_766,N_3523);
nand U8651 (N_8651,N_3402,N_778);
xor U8652 (N_8652,N_3399,N_2366);
nor U8653 (N_8653,N_113,N_4177);
xnor U8654 (N_8654,N_2799,N_2105);
or U8655 (N_8655,N_2662,N_187);
and U8656 (N_8656,N_2763,N_803);
nor U8657 (N_8657,N_1172,N_2099);
or U8658 (N_8658,N_2769,N_2260);
xor U8659 (N_8659,N_2122,N_2658);
nor U8660 (N_8660,N_3912,N_2364);
or U8661 (N_8661,N_668,N_3609);
or U8662 (N_8662,N_4132,N_3997);
xnor U8663 (N_8663,N_3414,N_2672);
xnor U8664 (N_8664,N_3051,N_4488);
nand U8665 (N_8665,N_3601,N_1275);
or U8666 (N_8666,N_295,N_2573);
nand U8667 (N_8667,N_1341,N_3491);
and U8668 (N_8668,N_1129,N_2121);
nor U8669 (N_8669,N_1668,N_1906);
nor U8670 (N_8670,N_4822,N_4915);
xor U8671 (N_8671,N_1232,N_4217);
and U8672 (N_8672,N_151,N_1493);
xnor U8673 (N_8673,N_818,N_1488);
nand U8674 (N_8674,N_2354,N_167);
or U8675 (N_8675,N_2719,N_1336);
nand U8676 (N_8676,N_3832,N_1547);
nand U8677 (N_8677,N_188,N_3421);
or U8678 (N_8678,N_2876,N_2228);
and U8679 (N_8679,N_94,N_241);
xnor U8680 (N_8680,N_3452,N_2694);
or U8681 (N_8681,N_2904,N_1813);
and U8682 (N_8682,N_1891,N_2752);
nand U8683 (N_8683,N_361,N_3382);
or U8684 (N_8684,N_3174,N_3969);
or U8685 (N_8685,N_1873,N_2207);
or U8686 (N_8686,N_1159,N_2698);
xnor U8687 (N_8687,N_1746,N_4359);
and U8688 (N_8688,N_1070,N_3214);
nor U8689 (N_8689,N_2223,N_522);
and U8690 (N_8690,N_1669,N_2110);
xor U8691 (N_8691,N_1399,N_2352);
nand U8692 (N_8692,N_262,N_3715);
nand U8693 (N_8693,N_3927,N_3345);
nor U8694 (N_8694,N_666,N_155);
or U8695 (N_8695,N_4906,N_4089);
nor U8696 (N_8696,N_526,N_948);
or U8697 (N_8697,N_752,N_1281);
or U8698 (N_8698,N_433,N_2667);
nand U8699 (N_8699,N_2833,N_4388);
nand U8700 (N_8700,N_2028,N_4584);
xnor U8701 (N_8701,N_4125,N_704);
and U8702 (N_8702,N_1899,N_3201);
nor U8703 (N_8703,N_3709,N_4552);
nor U8704 (N_8704,N_4273,N_4862);
xor U8705 (N_8705,N_3872,N_1966);
xor U8706 (N_8706,N_2983,N_4862);
or U8707 (N_8707,N_3873,N_1055);
or U8708 (N_8708,N_1311,N_3060);
and U8709 (N_8709,N_2810,N_3597);
xnor U8710 (N_8710,N_2265,N_3766);
or U8711 (N_8711,N_3525,N_4462);
nor U8712 (N_8712,N_3275,N_4602);
or U8713 (N_8713,N_1589,N_1217);
and U8714 (N_8714,N_2652,N_3001);
or U8715 (N_8715,N_4011,N_197);
nand U8716 (N_8716,N_1237,N_4731);
nor U8717 (N_8717,N_389,N_3356);
xor U8718 (N_8718,N_1200,N_1633);
nand U8719 (N_8719,N_1147,N_1680);
xnor U8720 (N_8720,N_856,N_1037);
or U8721 (N_8721,N_2591,N_1009);
or U8722 (N_8722,N_3845,N_3408);
and U8723 (N_8723,N_2897,N_4033);
nand U8724 (N_8724,N_4215,N_4954);
xor U8725 (N_8725,N_2834,N_3162);
xor U8726 (N_8726,N_4307,N_3661);
or U8727 (N_8727,N_639,N_1904);
xor U8728 (N_8728,N_3223,N_3893);
and U8729 (N_8729,N_3918,N_2814);
xnor U8730 (N_8730,N_2311,N_2043);
or U8731 (N_8731,N_3294,N_4774);
nor U8732 (N_8732,N_4818,N_2384);
nor U8733 (N_8733,N_2014,N_2999);
or U8734 (N_8734,N_2128,N_574);
and U8735 (N_8735,N_3475,N_4201);
nand U8736 (N_8736,N_1410,N_1728);
or U8737 (N_8737,N_4544,N_4610);
nand U8738 (N_8738,N_2025,N_3171);
xor U8739 (N_8739,N_874,N_3629);
xnor U8740 (N_8740,N_3498,N_209);
or U8741 (N_8741,N_613,N_4642);
and U8742 (N_8742,N_4169,N_1298);
nand U8743 (N_8743,N_3227,N_3226);
or U8744 (N_8744,N_4854,N_2458);
nor U8745 (N_8745,N_1817,N_229);
or U8746 (N_8746,N_204,N_4038);
and U8747 (N_8747,N_804,N_3575);
or U8748 (N_8748,N_916,N_2528);
nand U8749 (N_8749,N_2193,N_101);
nand U8750 (N_8750,N_1679,N_1526);
or U8751 (N_8751,N_930,N_2589);
nor U8752 (N_8752,N_2799,N_969);
nor U8753 (N_8753,N_3619,N_3370);
nand U8754 (N_8754,N_4605,N_1718);
xnor U8755 (N_8755,N_2916,N_4666);
nand U8756 (N_8756,N_2236,N_31);
xor U8757 (N_8757,N_643,N_3370);
xor U8758 (N_8758,N_4504,N_4463);
nand U8759 (N_8759,N_2142,N_3142);
xnor U8760 (N_8760,N_2895,N_484);
and U8761 (N_8761,N_3323,N_3092);
nor U8762 (N_8762,N_586,N_4998);
xnor U8763 (N_8763,N_3451,N_154);
xor U8764 (N_8764,N_1485,N_936);
nor U8765 (N_8765,N_1253,N_1805);
nand U8766 (N_8766,N_4041,N_1942);
nand U8767 (N_8767,N_1788,N_1576);
nand U8768 (N_8768,N_1279,N_629);
xor U8769 (N_8769,N_4344,N_4096);
or U8770 (N_8770,N_1318,N_1172);
nand U8771 (N_8771,N_534,N_3473);
and U8772 (N_8772,N_4222,N_4433);
or U8773 (N_8773,N_4607,N_2169);
and U8774 (N_8774,N_1700,N_837);
nand U8775 (N_8775,N_3293,N_1697);
nand U8776 (N_8776,N_2862,N_1348);
and U8777 (N_8777,N_3258,N_983);
nand U8778 (N_8778,N_250,N_2490);
nor U8779 (N_8779,N_504,N_4741);
nor U8780 (N_8780,N_4899,N_4292);
nor U8781 (N_8781,N_4610,N_2959);
nand U8782 (N_8782,N_727,N_4914);
or U8783 (N_8783,N_2323,N_2278);
or U8784 (N_8784,N_1472,N_857);
and U8785 (N_8785,N_3202,N_971);
nand U8786 (N_8786,N_3440,N_1124);
or U8787 (N_8787,N_1437,N_1196);
and U8788 (N_8788,N_3064,N_3699);
and U8789 (N_8789,N_812,N_1523);
nand U8790 (N_8790,N_4582,N_3797);
nand U8791 (N_8791,N_1239,N_3663);
or U8792 (N_8792,N_4325,N_3627);
or U8793 (N_8793,N_4167,N_1334);
nand U8794 (N_8794,N_4036,N_2620);
xnor U8795 (N_8795,N_561,N_4694);
nor U8796 (N_8796,N_991,N_4735);
and U8797 (N_8797,N_628,N_1426);
xnor U8798 (N_8798,N_424,N_2501);
nor U8799 (N_8799,N_147,N_2866);
or U8800 (N_8800,N_261,N_4098);
nor U8801 (N_8801,N_1367,N_3273);
nor U8802 (N_8802,N_2474,N_1328);
or U8803 (N_8803,N_3215,N_3692);
nand U8804 (N_8804,N_2553,N_448);
xor U8805 (N_8805,N_938,N_3980);
nand U8806 (N_8806,N_4680,N_2792);
and U8807 (N_8807,N_199,N_953);
xnor U8808 (N_8808,N_1939,N_4598);
or U8809 (N_8809,N_489,N_117);
nor U8810 (N_8810,N_1690,N_382);
xnor U8811 (N_8811,N_4468,N_3660);
or U8812 (N_8812,N_1806,N_2821);
nand U8813 (N_8813,N_1406,N_4922);
and U8814 (N_8814,N_1386,N_3907);
and U8815 (N_8815,N_3288,N_4949);
nand U8816 (N_8816,N_479,N_907);
or U8817 (N_8817,N_1243,N_3274);
nor U8818 (N_8818,N_4327,N_4117);
and U8819 (N_8819,N_859,N_669);
and U8820 (N_8820,N_4282,N_1221);
nand U8821 (N_8821,N_4575,N_1399);
nor U8822 (N_8822,N_1241,N_2161);
nor U8823 (N_8823,N_1278,N_6);
xor U8824 (N_8824,N_4881,N_1117);
and U8825 (N_8825,N_4136,N_4944);
xnor U8826 (N_8826,N_453,N_3500);
nor U8827 (N_8827,N_1179,N_4342);
or U8828 (N_8828,N_3371,N_1946);
nor U8829 (N_8829,N_622,N_3996);
nor U8830 (N_8830,N_21,N_3568);
nand U8831 (N_8831,N_445,N_4493);
nor U8832 (N_8832,N_405,N_3695);
xor U8833 (N_8833,N_548,N_555);
xnor U8834 (N_8834,N_1162,N_992);
xor U8835 (N_8835,N_1786,N_1557);
nand U8836 (N_8836,N_2800,N_2496);
xor U8837 (N_8837,N_4585,N_3299);
nor U8838 (N_8838,N_3912,N_4033);
xnor U8839 (N_8839,N_3173,N_4031);
and U8840 (N_8840,N_4343,N_4162);
xor U8841 (N_8841,N_4776,N_1963);
or U8842 (N_8842,N_943,N_4934);
nor U8843 (N_8843,N_1972,N_973);
nor U8844 (N_8844,N_734,N_3625);
xor U8845 (N_8845,N_1654,N_1154);
nor U8846 (N_8846,N_1248,N_3210);
nor U8847 (N_8847,N_40,N_4687);
or U8848 (N_8848,N_4408,N_4175);
xor U8849 (N_8849,N_4339,N_928);
or U8850 (N_8850,N_3468,N_3819);
nand U8851 (N_8851,N_2592,N_1526);
xnor U8852 (N_8852,N_3238,N_2098);
xor U8853 (N_8853,N_4478,N_1364);
or U8854 (N_8854,N_260,N_1521);
nor U8855 (N_8855,N_3515,N_2483);
xor U8856 (N_8856,N_2158,N_2822);
xnor U8857 (N_8857,N_1159,N_3966);
and U8858 (N_8858,N_4485,N_843);
nand U8859 (N_8859,N_2792,N_3823);
and U8860 (N_8860,N_4924,N_1894);
or U8861 (N_8861,N_551,N_3875);
nor U8862 (N_8862,N_198,N_4163);
xnor U8863 (N_8863,N_3926,N_1616);
nor U8864 (N_8864,N_2251,N_2013);
xnor U8865 (N_8865,N_2877,N_4055);
nand U8866 (N_8866,N_1146,N_4412);
or U8867 (N_8867,N_1365,N_796);
xnor U8868 (N_8868,N_4912,N_4834);
nand U8869 (N_8869,N_2914,N_230);
nor U8870 (N_8870,N_1739,N_63);
or U8871 (N_8871,N_1449,N_2175);
and U8872 (N_8872,N_2928,N_4007);
and U8873 (N_8873,N_4598,N_4679);
nor U8874 (N_8874,N_3785,N_3536);
nand U8875 (N_8875,N_4298,N_3437);
or U8876 (N_8876,N_2669,N_4358);
xor U8877 (N_8877,N_1791,N_4929);
xor U8878 (N_8878,N_4339,N_2915);
or U8879 (N_8879,N_681,N_2764);
nand U8880 (N_8880,N_3480,N_2330);
or U8881 (N_8881,N_1870,N_3777);
nor U8882 (N_8882,N_1344,N_2904);
or U8883 (N_8883,N_163,N_1451);
and U8884 (N_8884,N_3936,N_2230);
nor U8885 (N_8885,N_2031,N_3674);
nand U8886 (N_8886,N_3711,N_2199);
xor U8887 (N_8887,N_842,N_3385);
xor U8888 (N_8888,N_898,N_1544);
or U8889 (N_8889,N_2755,N_1633);
and U8890 (N_8890,N_3377,N_4960);
nand U8891 (N_8891,N_2671,N_2506);
nor U8892 (N_8892,N_2555,N_353);
or U8893 (N_8893,N_3431,N_770);
nor U8894 (N_8894,N_2969,N_1105);
xor U8895 (N_8895,N_4049,N_3072);
or U8896 (N_8896,N_4922,N_2311);
or U8897 (N_8897,N_1220,N_2169);
nor U8898 (N_8898,N_3685,N_2433);
xor U8899 (N_8899,N_4086,N_489);
nand U8900 (N_8900,N_3104,N_4580);
xor U8901 (N_8901,N_4557,N_4791);
or U8902 (N_8902,N_375,N_3298);
nand U8903 (N_8903,N_3177,N_1689);
nor U8904 (N_8904,N_4710,N_1370);
nand U8905 (N_8905,N_1425,N_1662);
or U8906 (N_8906,N_427,N_2608);
nand U8907 (N_8907,N_4736,N_2237);
nor U8908 (N_8908,N_999,N_2317);
and U8909 (N_8909,N_4793,N_3171);
nor U8910 (N_8910,N_2901,N_626);
nor U8911 (N_8911,N_3482,N_1849);
xor U8912 (N_8912,N_2677,N_1220);
xor U8913 (N_8913,N_4110,N_2319);
nor U8914 (N_8914,N_1029,N_229);
nor U8915 (N_8915,N_2133,N_2915);
nor U8916 (N_8916,N_3347,N_4741);
nand U8917 (N_8917,N_1021,N_2533);
or U8918 (N_8918,N_4655,N_456);
xnor U8919 (N_8919,N_2392,N_3119);
nor U8920 (N_8920,N_1063,N_1710);
nor U8921 (N_8921,N_4396,N_2610);
and U8922 (N_8922,N_4273,N_2581);
nand U8923 (N_8923,N_4019,N_8);
and U8924 (N_8924,N_1222,N_1171);
xor U8925 (N_8925,N_1776,N_3625);
or U8926 (N_8926,N_4832,N_1079);
xor U8927 (N_8927,N_1660,N_833);
nand U8928 (N_8928,N_4985,N_4255);
nand U8929 (N_8929,N_1072,N_87);
or U8930 (N_8930,N_2206,N_4053);
or U8931 (N_8931,N_3131,N_3825);
nand U8932 (N_8932,N_3938,N_3761);
or U8933 (N_8933,N_774,N_78);
nand U8934 (N_8934,N_602,N_2875);
nor U8935 (N_8935,N_1805,N_2084);
and U8936 (N_8936,N_948,N_2096);
nor U8937 (N_8937,N_63,N_1591);
or U8938 (N_8938,N_4407,N_3960);
or U8939 (N_8939,N_226,N_3039);
or U8940 (N_8940,N_2393,N_251);
nor U8941 (N_8941,N_881,N_2669);
xnor U8942 (N_8942,N_2563,N_4790);
or U8943 (N_8943,N_1760,N_3413);
or U8944 (N_8944,N_2877,N_4179);
xnor U8945 (N_8945,N_1884,N_4983);
xor U8946 (N_8946,N_2430,N_4205);
nand U8947 (N_8947,N_8,N_1505);
nand U8948 (N_8948,N_1045,N_993);
nand U8949 (N_8949,N_779,N_3693);
xnor U8950 (N_8950,N_3411,N_1831);
xnor U8951 (N_8951,N_3632,N_725);
xnor U8952 (N_8952,N_1869,N_4920);
nand U8953 (N_8953,N_92,N_355);
xnor U8954 (N_8954,N_1357,N_4814);
and U8955 (N_8955,N_2175,N_2753);
xor U8956 (N_8956,N_1712,N_4263);
and U8957 (N_8957,N_164,N_2929);
nor U8958 (N_8958,N_1651,N_195);
xnor U8959 (N_8959,N_2099,N_1597);
and U8960 (N_8960,N_1305,N_3506);
or U8961 (N_8961,N_417,N_4970);
or U8962 (N_8962,N_3055,N_2485);
nor U8963 (N_8963,N_824,N_4325);
and U8964 (N_8964,N_1590,N_445);
or U8965 (N_8965,N_3767,N_4347);
nand U8966 (N_8966,N_1841,N_2966);
nor U8967 (N_8967,N_1747,N_1522);
nand U8968 (N_8968,N_908,N_646);
and U8969 (N_8969,N_4220,N_3668);
and U8970 (N_8970,N_4409,N_3386);
nand U8971 (N_8971,N_4689,N_11);
nand U8972 (N_8972,N_722,N_1358);
nor U8973 (N_8973,N_1509,N_237);
xor U8974 (N_8974,N_2603,N_2779);
nor U8975 (N_8975,N_3636,N_4846);
or U8976 (N_8976,N_1897,N_4369);
or U8977 (N_8977,N_4102,N_1801);
or U8978 (N_8978,N_587,N_738);
xnor U8979 (N_8979,N_1103,N_919);
nand U8980 (N_8980,N_4564,N_2632);
xor U8981 (N_8981,N_4218,N_3225);
and U8982 (N_8982,N_3175,N_4686);
xnor U8983 (N_8983,N_3415,N_4622);
or U8984 (N_8984,N_2267,N_3509);
or U8985 (N_8985,N_2158,N_1769);
nand U8986 (N_8986,N_3727,N_1508);
and U8987 (N_8987,N_3183,N_1331);
and U8988 (N_8988,N_2108,N_4853);
nor U8989 (N_8989,N_3464,N_2106);
or U8990 (N_8990,N_2404,N_3045);
nand U8991 (N_8991,N_1359,N_4573);
and U8992 (N_8992,N_3218,N_4312);
and U8993 (N_8993,N_1881,N_4693);
nand U8994 (N_8994,N_2426,N_2660);
nand U8995 (N_8995,N_4620,N_4942);
nand U8996 (N_8996,N_2595,N_1882);
nor U8997 (N_8997,N_4523,N_2085);
nand U8998 (N_8998,N_2048,N_4615);
or U8999 (N_8999,N_2102,N_2062);
xnor U9000 (N_9000,N_1634,N_1071);
and U9001 (N_9001,N_1886,N_2415);
nor U9002 (N_9002,N_3984,N_52);
xnor U9003 (N_9003,N_539,N_1114);
or U9004 (N_9004,N_1790,N_1352);
xor U9005 (N_9005,N_1861,N_381);
or U9006 (N_9006,N_527,N_3992);
xnor U9007 (N_9007,N_2724,N_2588);
or U9008 (N_9008,N_1701,N_2556);
nand U9009 (N_9009,N_1198,N_68);
nor U9010 (N_9010,N_3297,N_3765);
nand U9011 (N_9011,N_34,N_3544);
nor U9012 (N_9012,N_2531,N_4953);
or U9013 (N_9013,N_1334,N_4046);
xnor U9014 (N_9014,N_1032,N_2815);
nand U9015 (N_9015,N_1378,N_473);
and U9016 (N_9016,N_2940,N_2120);
xnor U9017 (N_9017,N_4838,N_2377);
nand U9018 (N_9018,N_3377,N_1491);
or U9019 (N_9019,N_4479,N_2809);
nor U9020 (N_9020,N_828,N_205);
and U9021 (N_9021,N_2634,N_4268);
and U9022 (N_9022,N_2225,N_2806);
xnor U9023 (N_9023,N_1951,N_1171);
nor U9024 (N_9024,N_3358,N_3201);
nor U9025 (N_9025,N_1282,N_2496);
nor U9026 (N_9026,N_2273,N_2115);
xor U9027 (N_9027,N_4779,N_4917);
or U9028 (N_9028,N_2244,N_3349);
nand U9029 (N_9029,N_2290,N_2990);
or U9030 (N_9030,N_1517,N_2616);
xnor U9031 (N_9031,N_1856,N_897);
nand U9032 (N_9032,N_2921,N_127);
nor U9033 (N_9033,N_788,N_4706);
xor U9034 (N_9034,N_4610,N_3321);
nand U9035 (N_9035,N_760,N_4300);
and U9036 (N_9036,N_1399,N_1257);
or U9037 (N_9037,N_1694,N_1811);
xnor U9038 (N_9038,N_2530,N_3571);
xnor U9039 (N_9039,N_3625,N_2903);
and U9040 (N_9040,N_4554,N_1758);
xnor U9041 (N_9041,N_3338,N_1846);
and U9042 (N_9042,N_4092,N_463);
and U9043 (N_9043,N_2171,N_218);
nor U9044 (N_9044,N_2400,N_2482);
and U9045 (N_9045,N_2523,N_362);
nor U9046 (N_9046,N_2656,N_4194);
or U9047 (N_9047,N_3297,N_564);
nand U9048 (N_9048,N_3033,N_2018);
or U9049 (N_9049,N_3738,N_802);
xor U9050 (N_9050,N_4735,N_3899);
nor U9051 (N_9051,N_1672,N_2901);
nand U9052 (N_9052,N_3317,N_4625);
nor U9053 (N_9053,N_1106,N_4337);
xor U9054 (N_9054,N_2341,N_1912);
and U9055 (N_9055,N_4881,N_1123);
nand U9056 (N_9056,N_2355,N_946);
nor U9057 (N_9057,N_4169,N_2913);
nor U9058 (N_9058,N_4687,N_207);
nand U9059 (N_9059,N_52,N_1854);
nor U9060 (N_9060,N_3684,N_687);
xnor U9061 (N_9061,N_2566,N_481);
nor U9062 (N_9062,N_793,N_991);
xor U9063 (N_9063,N_4792,N_2702);
nor U9064 (N_9064,N_4169,N_4135);
or U9065 (N_9065,N_565,N_447);
xor U9066 (N_9066,N_2465,N_1232);
nor U9067 (N_9067,N_1994,N_3193);
nand U9068 (N_9068,N_1482,N_3375);
nor U9069 (N_9069,N_1743,N_2976);
nand U9070 (N_9070,N_492,N_4763);
and U9071 (N_9071,N_2645,N_4536);
or U9072 (N_9072,N_1412,N_974);
nand U9073 (N_9073,N_4469,N_1818);
nand U9074 (N_9074,N_1311,N_651);
nor U9075 (N_9075,N_3977,N_4187);
nand U9076 (N_9076,N_738,N_3535);
nor U9077 (N_9077,N_1276,N_3911);
xnor U9078 (N_9078,N_689,N_632);
and U9079 (N_9079,N_1482,N_3278);
nor U9080 (N_9080,N_4070,N_2355);
xnor U9081 (N_9081,N_70,N_3110);
nor U9082 (N_9082,N_2971,N_4373);
and U9083 (N_9083,N_1670,N_2689);
or U9084 (N_9084,N_3527,N_1495);
xor U9085 (N_9085,N_408,N_2569);
nand U9086 (N_9086,N_3574,N_2754);
or U9087 (N_9087,N_171,N_4115);
nor U9088 (N_9088,N_1990,N_2749);
or U9089 (N_9089,N_2335,N_1232);
nand U9090 (N_9090,N_3420,N_4947);
xnor U9091 (N_9091,N_476,N_3798);
nand U9092 (N_9092,N_4996,N_2987);
and U9093 (N_9093,N_1005,N_3420);
xnor U9094 (N_9094,N_605,N_1698);
and U9095 (N_9095,N_4115,N_1695);
nor U9096 (N_9096,N_2846,N_3852);
and U9097 (N_9097,N_4552,N_3527);
and U9098 (N_9098,N_3478,N_4245);
or U9099 (N_9099,N_4233,N_3880);
nor U9100 (N_9100,N_2569,N_2516);
and U9101 (N_9101,N_182,N_2330);
and U9102 (N_9102,N_3158,N_1781);
and U9103 (N_9103,N_4939,N_4430);
or U9104 (N_9104,N_1742,N_301);
nor U9105 (N_9105,N_242,N_1422);
nor U9106 (N_9106,N_4745,N_1929);
xor U9107 (N_9107,N_4269,N_1459);
nand U9108 (N_9108,N_3564,N_4694);
and U9109 (N_9109,N_4915,N_110);
nand U9110 (N_9110,N_3740,N_1560);
xnor U9111 (N_9111,N_3061,N_1999);
and U9112 (N_9112,N_2446,N_4753);
nand U9113 (N_9113,N_2595,N_3075);
xor U9114 (N_9114,N_4535,N_2555);
or U9115 (N_9115,N_1337,N_1963);
nor U9116 (N_9116,N_275,N_1534);
xor U9117 (N_9117,N_3258,N_1988);
or U9118 (N_9118,N_466,N_3091);
xnor U9119 (N_9119,N_1176,N_4443);
xor U9120 (N_9120,N_1691,N_4003);
or U9121 (N_9121,N_4220,N_579);
nor U9122 (N_9122,N_2439,N_3506);
or U9123 (N_9123,N_1090,N_1296);
nor U9124 (N_9124,N_2641,N_2033);
nor U9125 (N_9125,N_4053,N_934);
xnor U9126 (N_9126,N_1841,N_4826);
and U9127 (N_9127,N_1496,N_3677);
nand U9128 (N_9128,N_828,N_709);
nor U9129 (N_9129,N_2044,N_462);
nand U9130 (N_9130,N_3111,N_4042);
xnor U9131 (N_9131,N_3906,N_4591);
or U9132 (N_9132,N_1584,N_2221);
xnor U9133 (N_9133,N_1318,N_3209);
nor U9134 (N_9134,N_4106,N_411);
xnor U9135 (N_9135,N_1040,N_564);
nand U9136 (N_9136,N_2170,N_2581);
xor U9137 (N_9137,N_4972,N_3231);
xnor U9138 (N_9138,N_2899,N_3271);
xnor U9139 (N_9139,N_326,N_4772);
or U9140 (N_9140,N_3003,N_2051);
or U9141 (N_9141,N_2709,N_2571);
nand U9142 (N_9142,N_4676,N_4182);
and U9143 (N_9143,N_1814,N_3910);
or U9144 (N_9144,N_3291,N_4871);
nand U9145 (N_9145,N_1775,N_1712);
xnor U9146 (N_9146,N_2922,N_1523);
or U9147 (N_9147,N_927,N_4369);
nor U9148 (N_9148,N_1972,N_4125);
nand U9149 (N_9149,N_2470,N_2163);
nand U9150 (N_9150,N_3935,N_3210);
nand U9151 (N_9151,N_515,N_3465);
nor U9152 (N_9152,N_1056,N_4246);
or U9153 (N_9153,N_463,N_617);
or U9154 (N_9154,N_640,N_940);
nor U9155 (N_9155,N_778,N_696);
and U9156 (N_9156,N_4001,N_3433);
xor U9157 (N_9157,N_3510,N_2392);
or U9158 (N_9158,N_1339,N_2217);
and U9159 (N_9159,N_3082,N_2901);
and U9160 (N_9160,N_3088,N_3205);
nor U9161 (N_9161,N_1928,N_2748);
nand U9162 (N_9162,N_724,N_4664);
nor U9163 (N_9163,N_3138,N_4286);
nand U9164 (N_9164,N_4862,N_4095);
nand U9165 (N_9165,N_430,N_2550);
nand U9166 (N_9166,N_2771,N_3211);
and U9167 (N_9167,N_4409,N_4039);
nor U9168 (N_9168,N_855,N_365);
and U9169 (N_9169,N_1931,N_568);
or U9170 (N_9170,N_1109,N_3554);
or U9171 (N_9171,N_1095,N_51);
xor U9172 (N_9172,N_3135,N_3999);
or U9173 (N_9173,N_4048,N_520);
nand U9174 (N_9174,N_4606,N_3984);
and U9175 (N_9175,N_3150,N_3718);
nand U9176 (N_9176,N_1141,N_3094);
and U9177 (N_9177,N_692,N_2170);
xor U9178 (N_9178,N_2082,N_2296);
or U9179 (N_9179,N_200,N_4690);
or U9180 (N_9180,N_1099,N_1261);
xnor U9181 (N_9181,N_1784,N_2031);
or U9182 (N_9182,N_3984,N_3798);
nor U9183 (N_9183,N_4154,N_1700);
nor U9184 (N_9184,N_4716,N_2321);
nand U9185 (N_9185,N_2977,N_1115);
xor U9186 (N_9186,N_1923,N_4742);
nand U9187 (N_9187,N_4227,N_759);
nor U9188 (N_9188,N_2438,N_3190);
and U9189 (N_9189,N_1869,N_4780);
and U9190 (N_9190,N_2052,N_279);
or U9191 (N_9191,N_3256,N_3924);
nand U9192 (N_9192,N_2623,N_3952);
nand U9193 (N_9193,N_2196,N_4990);
and U9194 (N_9194,N_3732,N_542);
or U9195 (N_9195,N_2042,N_172);
xor U9196 (N_9196,N_3946,N_2516);
xor U9197 (N_9197,N_1912,N_2423);
and U9198 (N_9198,N_1315,N_3720);
and U9199 (N_9199,N_414,N_4145);
or U9200 (N_9200,N_4336,N_2215);
nand U9201 (N_9201,N_1226,N_2611);
nor U9202 (N_9202,N_4397,N_1015);
nand U9203 (N_9203,N_2450,N_379);
xor U9204 (N_9204,N_595,N_2414);
or U9205 (N_9205,N_2385,N_249);
xor U9206 (N_9206,N_751,N_3353);
xor U9207 (N_9207,N_2853,N_0);
nor U9208 (N_9208,N_374,N_2211);
nor U9209 (N_9209,N_761,N_2545);
xnor U9210 (N_9210,N_4940,N_2309);
or U9211 (N_9211,N_1971,N_3430);
nor U9212 (N_9212,N_4272,N_3863);
or U9213 (N_9213,N_4741,N_4273);
xnor U9214 (N_9214,N_4618,N_1119);
nor U9215 (N_9215,N_4042,N_3339);
xnor U9216 (N_9216,N_3731,N_3689);
nor U9217 (N_9217,N_1431,N_4778);
nor U9218 (N_9218,N_2061,N_2632);
or U9219 (N_9219,N_4922,N_2980);
nor U9220 (N_9220,N_4681,N_2211);
xnor U9221 (N_9221,N_3522,N_4175);
nor U9222 (N_9222,N_3903,N_4788);
or U9223 (N_9223,N_3022,N_2328);
and U9224 (N_9224,N_2020,N_1283);
nor U9225 (N_9225,N_1636,N_3420);
nand U9226 (N_9226,N_2249,N_2570);
xor U9227 (N_9227,N_1420,N_4782);
or U9228 (N_9228,N_2889,N_1634);
nor U9229 (N_9229,N_1021,N_3957);
xor U9230 (N_9230,N_2512,N_4114);
nor U9231 (N_9231,N_3680,N_720);
xnor U9232 (N_9232,N_2653,N_1197);
nor U9233 (N_9233,N_2034,N_2269);
xnor U9234 (N_9234,N_3189,N_4819);
or U9235 (N_9235,N_3428,N_3189);
and U9236 (N_9236,N_3401,N_2333);
or U9237 (N_9237,N_896,N_3200);
and U9238 (N_9238,N_1038,N_3783);
and U9239 (N_9239,N_394,N_30);
nand U9240 (N_9240,N_1891,N_3572);
nor U9241 (N_9241,N_4484,N_621);
xor U9242 (N_9242,N_4563,N_30);
nor U9243 (N_9243,N_406,N_978);
nor U9244 (N_9244,N_3806,N_3959);
or U9245 (N_9245,N_3324,N_1602);
and U9246 (N_9246,N_676,N_650);
nand U9247 (N_9247,N_3178,N_1695);
or U9248 (N_9248,N_4276,N_2522);
nor U9249 (N_9249,N_2240,N_1601);
nand U9250 (N_9250,N_4240,N_2540);
and U9251 (N_9251,N_1761,N_3718);
nand U9252 (N_9252,N_3071,N_1102);
or U9253 (N_9253,N_160,N_3138);
nor U9254 (N_9254,N_4355,N_2952);
or U9255 (N_9255,N_4713,N_3869);
xor U9256 (N_9256,N_3341,N_162);
or U9257 (N_9257,N_2744,N_1732);
and U9258 (N_9258,N_3561,N_4454);
xor U9259 (N_9259,N_59,N_1140);
xor U9260 (N_9260,N_2217,N_4816);
and U9261 (N_9261,N_751,N_2858);
nand U9262 (N_9262,N_2870,N_991);
xor U9263 (N_9263,N_2379,N_3788);
or U9264 (N_9264,N_1664,N_218);
xnor U9265 (N_9265,N_4860,N_4224);
nand U9266 (N_9266,N_618,N_4251);
nand U9267 (N_9267,N_369,N_1890);
or U9268 (N_9268,N_863,N_1513);
nand U9269 (N_9269,N_1419,N_3409);
and U9270 (N_9270,N_213,N_2580);
xor U9271 (N_9271,N_259,N_1981);
and U9272 (N_9272,N_1753,N_3796);
xnor U9273 (N_9273,N_3549,N_4592);
nand U9274 (N_9274,N_105,N_701);
nor U9275 (N_9275,N_4349,N_1153);
and U9276 (N_9276,N_3516,N_1186);
or U9277 (N_9277,N_3437,N_3427);
xnor U9278 (N_9278,N_2161,N_39);
nand U9279 (N_9279,N_1413,N_4819);
nor U9280 (N_9280,N_4208,N_3572);
nand U9281 (N_9281,N_3815,N_3190);
or U9282 (N_9282,N_701,N_4876);
or U9283 (N_9283,N_1001,N_595);
nor U9284 (N_9284,N_437,N_4315);
xor U9285 (N_9285,N_4996,N_943);
xor U9286 (N_9286,N_4664,N_2200);
nand U9287 (N_9287,N_4375,N_1096);
or U9288 (N_9288,N_660,N_4709);
nand U9289 (N_9289,N_3899,N_955);
and U9290 (N_9290,N_1378,N_147);
nand U9291 (N_9291,N_409,N_709);
and U9292 (N_9292,N_1865,N_2083);
nor U9293 (N_9293,N_527,N_4124);
nor U9294 (N_9294,N_1843,N_4548);
xnor U9295 (N_9295,N_1042,N_3016);
and U9296 (N_9296,N_3122,N_1752);
and U9297 (N_9297,N_754,N_949);
xor U9298 (N_9298,N_4113,N_3930);
xor U9299 (N_9299,N_3399,N_4671);
nand U9300 (N_9300,N_3235,N_1935);
or U9301 (N_9301,N_2779,N_4749);
and U9302 (N_9302,N_1607,N_144);
nand U9303 (N_9303,N_2728,N_367);
nor U9304 (N_9304,N_718,N_3252);
or U9305 (N_9305,N_3125,N_2327);
nand U9306 (N_9306,N_2426,N_3978);
nor U9307 (N_9307,N_29,N_1912);
xnor U9308 (N_9308,N_3700,N_3573);
and U9309 (N_9309,N_4053,N_447);
nand U9310 (N_9310,N_1428,N_3313);
nand U9311 (N_9311,N_4305,N_4530);
nor U9312 (N_9312,N_2649,N_312);
or U9313 (N_9313,N_10,N_4334);
nand U9314 (N_9314,N_407,N_1036);
xor U9315 (N_9315,N_2714,N_105);
nor U9316 (N_9316,N_1748,N_706);
xnor U9317 (N_9317,N_326,N_3287);
or U9318 (N_9318,N_528,N_2319);
or U9319 (N_9319,N_4991,N_4457);
nand U9320 (N_9320,N_167,N_2052);
or U9321 (N_9321,N_841,N_135);
and U9322 (N_9322,N_3525,N_2685);
and U9323 (N_9323,N_4471,N_328);
nor U9324 (N_9324,N_2287,N_815);
and U9325 (N_9325,N_2823,N_3802);
and U9326 (N_9326,N_2613,N_4497);
or U9327 (N_9327,N_2827,N_4650);
nand U9328 (N_9328,N_3974,N_276);
xor U9329 (N_9329,N_4244,N_2896);
xnor U9330 (N_9330,N_3461,N_3579);
xor U9331 (N_9331,N_1375,N_2099);
and U9332 (N_9332,N_212,N_3177);
nor U9333 (N_9333,N_819,N_3559);
nor U9334 (N_9334,N_3955,N_703);
and U9335 (N_9335,N_4132,N_2507);
nor U9336 (N_9336,N_3320,N_1500);
nand U9337 (N_9337,N_4805,N_4934);
nand U9338 (N_9338,N_415,N_1514);
xnor U9339 (N_9339,N_4582,N_3570);
nor U9340 (N_9340,N_3266,N_491);
and U9341 (N_9341,N_3219,N_405);
or U9342 (N_9342,N_1452,N_1390);
xor U9343 (N_9343,N_2328,N_3127);
xnor U9344 (N_9344,N_4674,N_4402);
nor U9345 (N_9345,N_1824,N_1466);
or U9346 (N_9346,N_300,N_3722);
and U9347 (N_9347,N_2950,N_3570);
xnor U9348 (N_9348,N_1107,N_1898);
nor U9349 (N_9349,N_3789,N_1519);
nor U9350 (N_9350,N_2493,N_1648);
nor U9351 (N_9351,N_1429,N_3874);
nand U9352 (N_9352,N_1286,N_3050);
and U9353 (N_9353,N_278,N_4685);
nand U9354 (N_9354,N_3629,N_2571);
nor U9355 (N_9355,N_4606,N_3024);
and U9356 (N_9356,N_654,N_3099);
nand U9357 (N_9357,N_1501,N_4400);
or U9358 (N_9358,N_3947,N_4096);
and U9359 (N_9359,N_2929,N_3329);
nand U9360 (N_9360,N_1779,N_4139);
xnor U9361 (N_9361,N_2715,N_2655);
xnor U9362 (N_9362,N_1270,N_3655);
nor U9363 (N_9363,N_1329,N_2220);
or U9364 (N_9364,N_369,N_3770);
and U9365 (N_9365,N_314,N_893);
xnor U9366 (N_9366,N_2260,N_3674);
and U9367 (N_9367,N_667,N_2315);
and U9368 (N_9368,N_2331,N_460);
or U9369 (N_9369,N_3065,N_4167);
nor U9370 (N_9370,N_3438,N_1657);
xnor U9371 (N_9371,N_581,N_4874);
nand U9372 (N_9372,N_1483,N_150);
nor U9373 (N_9373,N_2516,N_3999);
nand U9374 (N_9374,N_3530,N_4409);
and U9375 (N_9375,N_2056,N_533);
nor U9376 (N_9376,N_2531,N_3152);
and U9377 (N_9377,N_3003,N_2576);
nor U9378 (N_9378,N_442,N_1533);
or U9379 (N_9379,N_4223,N_4525);
xnor U9380 (N_9380,N_2850,N_4815);
xor U9381 (N_9381,N_4855,N_4294);
and U9382 (N_9382,N_4830,N_4924);
or U9383 (N_9383,N_1817,N_2400);
nand U9384 (N_9384,N_766,N_2226);
and U9385 (N_9385,N_2630,N_3702);
xnor U9386 (N_9386,N_1886,N_4237);
nor U9387 (N_9387,N_3051,N_2177);
xnor U9388 (N_9388,N_321,N_3370);
or U9389 (N_9389,N_2502,N_3046);
nand U9390 (N_9390,N_3274,N_3941);
nand U9391 (N_9391,N_3829,N_2086);
or U9392 (N_9392,N_4725,N_218);
nand U9393 (N_9393,N_2353,N_4403);
nand U9394 (N_9394,N_2569,N_4164);
nor U9395 (N_9395,N_1383,N_168);
nand U9396 (N_9396,N_2344,N_2084);
nor U9397 (N_9397,N_4230,N_2008);
nor U9398 (N_9398,N_1444,N_3162);
xnor U9399 (N_9399,N_189,N_3294);
or U9400 (N_9400,N_3674,N_1286);
xor U9401 (N_9401,N_716,N_1493);
and U9402 (N_9402,N_1881,N_1328);
and U9403 (N_9403,N_3430,N_1164);
nor U9404 (N_9404,N_4729,N_4925);
xnor U9405 (N_9405,N_2729,N_792);
nor U9406 (N_9406,N_3306,N_1588);
and U9407 (N_9407,N_2701,N_1048);
nand U9408 (N_9408,N_350,N_4551);
and U9409 (N_9409,N_4403,N_513);
or U9410 (N_9410,N_3133,N_72);
nor U9411 (N_9411,N_4542,N_3781);
and U9412 (N_9412,N_3379,N_211);
or U9413 (N_9413,N_550,N_472);
xor U9414 (N_9414,N_3355,N_2076);
xor U9415 (N_9415,N_3600,N_4667);
nor U9416 (N_9416,N_3920,N_4146);
nor U9417 (N_9417,N_1957,N_3022);
nand U9418 (N_9418,N_3682,N_4343);
xnor U9419 (N_9419,N_3400,N_1990);
xor U9420 (N_9420,N_1133,N_17);
or U9421 (N_9421,N_899,N_1177);
and U9422 (N_9422,N_3663,N_3847);
or U9423 (N_9423,N_1533,N_3846);
xnor U9424 (N_9424,N_790,N_3291);
and U9425 (N_9425,N_136,N_1514);
and U9426 (N_9426,N_1725,N_1646);
nand U9427 (N_9427,N_4512,N_3490);
nand U9428 (N_9428,N_1216,N_4290);
nand U9429 (N_9429,N_649,N_3284);
nand U9430 (N_9430,N_1251,N_2997);
nor U9431 (N_9431,N_4745,N_1828);
xnor U9432 (N_9432,N_2200,N_4959);
nor U9433 (N_9433,N_1356,N_2881);
xor U9434 (N_9434,N_3267,N_963);
nor U9435 (N_9435,N_1809,N_115);
xor U9436 (N_9436,N_154,N_1004);
nand U9437 (N_9437,N_1151,N_2575);
or U9438 (N_9438,N_4410,N_2436);
or U9439 (N_9439,N_2222,N_141);
xor U9440 (N_9440,N_102,N_1921);
or U9441 (N_9441,N_1759,N_1301);
nand U9442 (N_9442,N_316,N_4052);
xor U9443 (N_9443,N_470,N_3153);
nand U9444 (N_9444,N_2673,N_2005);
or U9445 (N_9445,N_3759,N_1401);
and U9446 (N_9446,N_1266,N_3207);
and U9447 (N_9447,N_2362,N_3382);
xor U9448 (N_9448,N_1833,N_2268);
nand U9449 (N_9449,N_2398,N_760);
xor U9450 (N_9450,N_4234,N_4323);
or U9451 (N_9451,N_854,N_1820);
or U9452 (N_9452,N_2632,N_4685);
or U9453 (N_9453,N_3422,N_4847);
nor U9454 (N_9454,N_4564,N_4565);
and U9455 (N_9455,N_4225,N_4578);
xor U9456 (N_9456,N_4980,N_864);
nor U9457 (N_9457,N_4750,N_1435);
nor U9458 (N_9458,N_3080,N_2249);
xor U9459 (N_9459,N_772,N_1119);
xor U9460 (N_9460,N_4232,N_4082);
nor U9461 (N_9461,N_4415,N_3617);
xor U9462 (N_9462,N_3528,N_3050);
and U9463 (N_9463,N_1910,N_746);
nand U9464 (N_9464,N_4584,N_2014);
nand U9465 (N_9465,N_1031,N_1791);
and U9466 (N_9466,N_4818,N_3115);
nand U9467 (N_9467,N_1570,N_597);
xnor U9468 (N_9468,N_2666,N_736);
and U9469 (N_9469,N_3059,N_1369);
or U9470 (N_9470,N_327,N_2858);
nand U9471 (N_9471,N_228,N_4574);
and U9472 (N_9472,N_1779,N_2524);
nand U9473 (N_9473,N_2830,N_3328);
xor U9474 (N_9474,N_2696,N_2130);
nor U9475 (N_9475,N_324,N_3416);
nor U9476 (N_9476,N_1097,N_2661);
nor U9477 (N_9477,N_3435,N_4506);
or U9478 (N_9478,N_1492,N_2027);
and U9479 (N_9479,N_2867,N_4527);
nor U9480 (N_9480,N_3643,N_3769);
and U9481 (N_9481,N_3820,N_1515);
or U9482 (N_9482,N_938,N_4840);
nand U9483 (N_9483,N_682,N_2939);
nand U9484 (N_9484,N_3212,N_4705);
nor U9485 (N_9485,N_3605,N_3267);
nand U9486 (N_9486,N_2826,N_630);
nor U9487 (N_9487,N_1720,N_4908);
nor U9488 (N_9488,N_2319,N_4419);
nor U9489 (N_9489,N_4886,N_1048);
xnor U9490 (N_9490,N_1468,N_1379);
xor U9491 (N_9491,N_116,N_1870);
and U9492 (N_9492,N_1529,N_2782);
xor U9493 (N_9493,N_15,N_4344);
nor U9494 (N_9494,N_3078,N_1018);
xor U9495 (N_9495,N_2464,N_1774);
xor U9496 (N_9496,N_882,N_4964);
xor U9497 (N_9497,N_1318,N_3322);
and U9498 (N_9498,N_1506,N_461);
nor U9499 (N_9499,N_2443,N_4901);
nand U9500 (N_9500,N_4035,N_643);
or U9501 (N_9501,N_1151,N_2896);
or U9502 (N_9502,N_4277,N_3792);
xor U9503 (N_9503,N_1596,N_2357);
and U9504 (N_9504,N_3167,N_821);
or U9505 (N_9505,N_52,N_4928);
xor U9506 (N_9506,N_2356,N_2451);
and U9507 (N_9507,N_53,N_3189);
or U9508 (N_9508,N_2661,N_1677);
nor U9509 (N_9509,N_3964,N_1789);
nor U9510 (N_9510,N_672,N_2542);
nand U9511 (N_9511,N_4316,N_4972);
xnor U9512 (N_9512,N_4108,N_4818);
and U9513 (N_9513,N_2331,N_942);
or U9514 (N_9514,N_3060,N_2846);
xor U9515 (N_9515,N_1312,N_2727);
xnor U9516 (N_9516,N_213,N_4267);
and U9517 (N_9517,N_3629,N_2518);
xor U9518 (N_9518,N_3313,N_1156);
nand U9519 (N_9519,N_4530,N_4228);
and U9520 (N_9520,N_3860,N_770);
or U9521 (N_9521,N_3894,N_2985);
nand U9522 (N_9522,N_4839,N_2830);
and U9523 (N_9523,N_2959,N_1168);
nand U9524 (N_9524,N_2036,N_3619);
nand U9525 (N_9525,N_3396,N_2345);
nand U9526 (N_9526,N_4922,N_813);
and U9527 (N_9527,N_3595,N_2537);
xor U9528 (N_9528,N_1369,N_1944);
nand U9529 (N_9529,N_2918,N_2148);
nor U9530 (N_9530,N_3433,N_3646);
and U9531 (N_9531,N_4880,N_418);
or U9532 (N_9532,N_2619,N_4653);
xor U9533 (N_9533,N_4768,N_1843);
or U9534 (N_9534,N_1034,N_834);
nand U9535 (N_9535,N_2752,N_3235);
and U9536 (N_9536,N_2221,N_2371);
and U9537 (N_9537,N_470,N_4152);
and U9538 (N_9538,N_4870,N_1233);
xnor U9539 (N_9539,N_4411,N_3552);
or U9540 (N_9540,N_1577,N_1726);
nand U9541 (N_9541,N_1292,N_1683);
nor U9542 (N_9542,N_2607,N_473);
and U9543 (N_9543,N_551,N_1284);
xnor U9544 (N_9544,N_2226,N_4426);
or U9545 (N_9545,N_3672,N_2609);
nand U9546 (N_9546,N_4092,N_2108);
xor U9547 (N_9547,N_1411,N_4114);
xnor U9548 (N_9548,N_3019,N_1232);
xor U9549 (N_9549,N_1015,N_1447);
and U9550 (N_9550,N_1341,N_4253);
nand U9551 (N_9551,N_603,N_2423);
or U9552 (N_9552,N_2750,N_4405);
nor U9553 (N_9553,N_4527,N_600);
nand U9554 (N_9554,N_785,N_2193);
nand U9555 (N_9555,N_2182,N_220);
or U9556 (N_9556,N_721,N_4454);
xor U9557 (N_9557,N_1683,N_4378);
or U9558 (N_9558,N_1514,N_3830);
nor U9559 (N_9559,N_4817,N_1877);
and U9560 (N_9560,N_3748,N_2958);
xor U9561 (N_9561,N_764,N_3363);
xor U9562 (N_9562,N_676,N_4949);
nor U9563 (N_9563,N_3328,N_450);
and U9564 (N_9564,N_2641,N_4303);
nand U9565 (N_9565,N_16,N_4709);
nor U9566 (N_9566,N_3284,N_2603);
xnor U9567 (N_9567,N_4930,N_1461);
or U9568 (N_9568,N_4243,N_3576);
nand U9569 (N_9569,N_3480,N_679);
nor U9570 (N_9570,N_2694,N_2148);
xor U9571 (N_9571,N_1627,N_4749);
nor U9572 (N_9572,N_263,N_1235);
xor U9573 (N_9573,N_2735,N_4535);
or U9574 (N_9574,N_859,N_1626);
or U9575 (N_9575,N_3138,N_2840);
nor U9576 (N_9576,N_3244,N_237);
nor U9577 (N_9577,N_3578,N_984);
xor U9578 (N_9578,N_2930,N_864);
nand U9579 (N_9579,N_3165,N_4199);
and U9580 (N_9580,N_2122,N_4189);
and U9581 (N_9581,N_392,N_2311);
or U9582 (N_9582,N_4565,N_603);
and U9583 (N_9583,N_3054,N_647);
nand U9584 (N_9584,N_3266,N_4823);
and U9585 (N_9585,N_3764,N_806);
xor U9586 (N_9586,N_3806,N_3109);
and U9587 (N_9587,N_2355,N_4432);
and U9588 (N_9588,N_353,N_1857);
or U9589 (N_9589,N_1655,N_319);
and U9590 (N_9590,N_4348,N_1561);
nor U9591 (N_9591,N_1224,N_4366);
xor U9592 (N_9592,N_2161,N_3444);
or U9593 (N_9593,N_1283,N_2618);
or U9594 (N_9594,N_2884,N_1166);
nor U9595 (N_9595,N_1458,N_3167);
or U9596 (N_9596,N_1678,N_3347);
nor U9597 (N_9597,N_2431,N_543);
or U9598 (N_9598,N_4444,N_4784);
and U9599 (N_9599,N_2033,N_2214);
and U9600 (N_9600,N_2739,N_2345);
nor U9601 (N_9601,N_2792,N_2106);
or U9602 (N_9602,N_1766,N_3816);
and U9603 (N_9603,N_4605,N_4404);
and U9604 (N_9604,N_2608,N_67);
and U9605 (N_9605,N_1322,N_559);
nor U9606 (N_9606,N_314,N_4007);
or U9607 (N_9607,N_116,N_1158);
nor U9608 (N_9608,N_282,N_4909);
xor U9609 (N_9609,N_3524,N_2156);
xnor U9610 (N_9610,N_3459,N_3333);
or U9611 (N_9611,N_3943,N_1738);
and U9612 (N_9612,N_4022,N_1313);
nor U9613 (N_9613,N_1398,N_2153);
nor U9614 (N_9614,N_18,N_395);
or U9615 (N_9615,N_494,N_4944);
and U9616 (N_9616,N_3414,N_576);
or U9617 (N_9617,N_491,N_84);
and U9618 (N_9618,N_3830,N_4648);
nor U9619 (N_9619,N_1593,N_2964);
xnor U9620 (N_9620,N_2120,N_4653);
or U9621 (N_9621,N_4677,N_3155);
or U9622 (N_9622,N_1540,N_2409);
and U9623 (N_9623,N_4616,N_3198);
or U9624 (N_9624,N_297,N_1133);
xnor U9625 (N_9625,N_1343,N_4803);
xnor U9626 (N_9626,N_361,N_1075);
and U9627 (N_9627,N_2673,N_2177);
xor U9628 (N_9628,N_4924,N_1269);
or U9629 (N_9629,N_2239,N_1327);
nand U9630 (N_9630,N_981,N_1039);
nand U9631 (N_9631,N_2646,N_2659);
nor U9632 (N_9632,N_4105,N_1830);
nand U9633 (N_9633,N_4799,N_4115);
xnor U9634 (N_9634,N_1344,N_1974);
nor U9635 (N_9635,N_3198,N_1722);
and U9636 (N_9636,N_4139,N_4987);
nor U9637 (N_9637,N_2957,N_1647);
nor U9638 (N_9638,N_1534,N_298);
and U9639 (N_9639,N_1371,N_4590);
or U9640 (N_9640,N_392,N_3341);
or U9641 (N_9641,N_676,N_2382);
nor U9642 (N_9642,N_2545,N_2998);
xor U9643 (N_9643,N_750,N_3609);
nor U9644 (N_9644,N_67,N_3063);
nand U9645 (N_9645,N_791,N_3355);
and U9646 (N_9646,N_1437,N_3530);
nor U9647 (N_9647,N_1364,N_2320);
nand U9648 (N_9648,N_3704,N_3505);
or U9649 (N_9649,N_3197,N_3143);
nor U9650 (N_9650,N_2306,N_2950);
nor U9651 (N_9651,N_2712,N_1156);
nand U9652 (N_9652,N_295,N_6);
nand U9653 (N_9653,N_2207,N_1304);
nand U9654 (N_9654,N_2705,N_1562);
nor U9655 (N_9655,N_720,N_853);
and U9656 (N_9656,N_2650,N_782);
xor U9657 (N_9657,N_415,N_4236);
or U9658 (N_9658,N_2867,N_4102);
nor U9659 (N_9659,N_3366,N_3206);
and U9660 (N_9660,N_1041,N_1773);
xor U9661 (N_9661,N_4766,N_1658);
and U9662 (N_9662,N_3009,N_48);
xor U9663 (N_9663,N_1579,N_2359);
or U9664 (N_9664,N_3091,N_4334);
nor U9665 (N_9665,N_323,N_954);
and U9666 (N_9666,N_1431,N_1899);
xor U9667 (N_9667,N_3338,N_3096);
and U9668 (N_9668,N_593,N_2834);
nand U9669 (N_9669,N_838,N_2310);
xor U9670 (N_9670,N_323,N_2216);
nor U9671 (N_9671,N_233,N_1448);
nand U9672 (N_9672,N_902,N_2397);
and U9673 (N_9673,N_889,N_3188);
xor U9674 (N_9674,N_1984,N_2519);
xnor U9675 (N_9675,N_2936,N_1391);
or U9676 (N_9676,N_2066,N_1403);
or U9677 (N_9677,N_3479,N_1584);
nand U9678 (N_9678,N_4697,N_4744);
nand U9679 (N_9679,N_1598,N_2945);
and U9680 (N_9680,N_1515,N_3422);
nand U9681 (N_9681,N_3644,N_3589);
xnor U9682 (N_9682,N_4565,N_1429);
xor U9683 (N_9683,N_3488,N_543);
nand U9684 (N_9684,N_4541,N_1748);
and U9685 (N_9685,N_3672,N_2103);
nor U9686 (N_9686,N_3225,N_365);
or U9687 (N_9687,N_3644,N_1873);
nor U9688 (N_9688,N_537,N_3840);
and U9689 (N_9689,N_3235,N_4197);
or U9690 (N_9690,N_2695,N_4363);
nor U9691 (N_9691,N_4241,N_4829);
nor U9692 (N_9692,N_2644,N_4931);
nand U9693 (N_9693,N_3739,N_1422);
and U9694 (N_9694,N_4026,N_3088);
or U9695 (N_9695,N_1168,N_3460);
xor U9696 (N_9696,N_65,N_112);
nor U9697 (N_9697,N_615,N_3341);
nand U9698 (N_9698,N_4791,N_946);
and U9699 (N_9699,N_3037,N_3145);
nor U9700 (N_9700,N_4464,N_3681);
and U9701 (N_9701,N_262,N_2822);
nand U9702 (N_9702,N_1503,N_541);
nand U9703 (N_9703,N_2616,N_3944);
and U9704 (N_9704,N_1858,N_4686);
nor U9705 (N_9705,N_1876,N_2168);
xnor U9706 (N_9706,N_4972,N_1862);
or U9707 (N_9707,N_2755,N_605);
nand U9708 (N_9708,N_16,N_1215);
and U9709 (N_9709,N_2902,N_4784);
nand U9710 (N_9710,N_157,N_1713);
xor U9711 (N_9711,N_4851,N_4512);
xor U9712 (N_9712,N_511,N_2415);
or U9713 (N_9713,N_1562,N_2610);
nor U9714 (N_9714,N_2655,N_3439);
or U9715 (N_9715,N_685,N_1509);
or U9716 (N_9716,N_3562,N_3508);
and U9717 (N_9717,N_846,N_4571);
xor U9718 (N_9718,N_2816,N_4847);
nor U9719 (N_9719,N_1508,N_4718);
xor U9720 (N_9720,N_851,N_3986);
nor U9721 (N_9721,N_956,N_4838);
or U9722 (N_9722,N_3474,N_4648);
and U9723 (N_9723,N_4333,N_4526);
nand U9724 (N_9724,N_60,N_232);
xnor U9725 (N_9725,N_957,N_3498);
or U9726 (N_9726,N_2735,N_332);
or U9727 (N_9727,N_890,N_4058);
nand U9728 (N_9728,N_2704,N_3795);
and U9729 (N_9729,N_2730,N_1916);
or U9730 (N_9730,N_4018,N_3424);
xnor U9731 (N_9731,N_1867,N_4219);
nand U9732 (N_9732,N_235,N_3009);
nor U9733 (N_9733,N_3396,N_2710);
or U9734 (N_9734,N_3507,N_297);
xnor U9735 (N_9735,N_847,N_2847);
xnor U9736 (N_9736,N_3851,N_2740);
nand U9737 (N_9737,N_944,N_940);
and U9738 (N_9738,N_530,N_641);
xor U9739 (N_9739,N_2508,N_1470);
nor U9740 (N_9740,N_919,N_4298);
and U9741 (N_9741,N_3129,N_4019);
xnor U9742 (N_9742,N_1290,N_3958);
xor U9743 (N_9743,N_2163,N_1893);
xor U9744 (N_9744,N_3218,N_2637);
and U9745 (N_9745,N_3022,N_4443);
nor U9746 (N_9746,N_843,N_1601);
or U9747 (N_9747,N_460,N_2948);
xnor U9748 (N_9748,N_4739,N_1748);
xor U9749 (N_9749,N_827,N_4959);
and U9750 (N_9750,N_1327,N_1718);
nand U9751 (N_9751,N_3364,N_110);
nor U9752 (N_9752,N_2334,N_3808);
nor U9753 (N_9753,N_3139,N_1218);
or U9754 (N_9754,N_2964,N_531);
or U9755 (N_9755,N_2724,N_4980);
and U9756 (N_9756,N_4535,N_1587);
xnor U9757 (N_9757,N_52,N_4389);
nand U9758 (N_9758,N_4656,N_770);
and U9759 (N_9759,N_3767,N_1323);
nand U9760 (N_9760,N_2599,N_3293);
xnor U9761 (N_9761,N_3226,N_2231);
or U9762 (N_9762,N_2513,N_1709);
xor U9763 (N_9763,N_3001,N_4394);
nand U9764 (N_9764,N_4301,N_143);
nor U9765 (N_9765,N_4135,N_2130);
nor U9766 (N_9766,N_2738,N_3959);
and U9767 (N_9767,N_4897,N_1825);
xnor U9768 (N_9768,N_4948,N_1903);
nand U9769 (N_9769,N_1180,N_1462);
and U9770 (N_9770,N_3975,N_845);
nand U9771 (N_9771,N_2668,N_3146);
and U9772 (N_9772,N_1951,N_2841);
nor U9773 (N_9773,N_2624,N_4056);
and U9774 (N_9774,N_2289,N_2342);
xnor U9775 (N_9775,N_2997,N_1303);
xnor U9776 (N_9776,N_2752,N_4514);
nor U9777 (N_9777,N_894,N_3402);
and U9778 (N_9778,N_3906,N_2210);
nor U9779 (N_9779,N_793,N_797);
and U9780 (N_9780,N_2640,N_1943);
or U9781 (N_9781,N_3806,N_733);
or U9782 (N_9782,N_2601,N_3719);
nor U9783 (N_9783,N_1506,N_4132);
nor U9784 (N_9784,N_3559,N_4045);
and U9785 (N_9785,N_533,N_4742);
nor U9786 (N_9786,N_4880,N_3482);
xor U9787 (N_9787,N_1208,N_4115);
xor U9788 (N_9788,N_797,N_3252);
nor U9789 (N_9789,N_3793,N_3987);
or U9790 (N_9790,N_1492,N_1045);
nor U9791 (N_9791,N_2732,N_3213);
and U9792 (N_9792,N_3205,N_3502);
xnor U9793 (N_9793,N_1759,N_3015);
or U9794 (N_9794,N_4555,N_1364);
or U9795 (N_9795,N_502,N_4683);
nor U9796 (N_9796,N_1413,N_4902);
nor U9797 (N_9797,N_3933,N_993);
xnor U9798 (N_9798,N_1430,N_4036);
xor U9799 (N_9799,N_429,N_2349);
or U9800 (N_9800,N_2603,N_3219);
or U9801 (N_9801,N_4510,N_2564);
nor U9802 (N_9802,N_4015,N_4885);
nand U9803 (N_9803,N_4201,N_2543);
nor U9804 (N_9804,N_2142,N_1130);
and U9805 (N_9805,N_1580,N_4751);
nand U9806 (N_9806,N_4595,N_3947);
nand U9807 (N_9807,N_4822,N_1937);
nand U9808 (N_9808,N_4638,N_2500);
and U9809 (N_9809,N_4381,N_2138);
or U9810 (N_9810,N_3294,N_3524);
and U9811 (N_9811,N_1308,N_973);
nor U9812 (N_9812,N_2692,N_800);
nand U9813 (N_9813,N_1224,N_2587);
xor U9814 (N_9814,N_444,N_2592);
or U9815 (N_9815,N_554,N_1976);
or U9816 (N_9816,N_4413,N_1945);
or U9817 (N_9817,N_3972,N_3937);
or U9818 (N_9818,N_4123,N_3503);
and U9819 (N_9819,N_1122,N_1716);
nand U9820 (N_9820,N_237,N_3279);
xnor U9821 (N_9821,N_3330,N_2917);
nor U9822 (N_9822,N_3843,N_3987);
or U9823 (N_9823,N_4780,N_3790);
nand U9824 (N_9824,N_3243,N_2837);
and U9825 (N_9825,N_4976,N_4694);
xor U9826 (N_9826,N_460,N_4759);
xnor U9827 (N_9827,N_64,N_1791);
nand U9828 (N_9828,N_2785,N_2902);
nand U9829 (N_9829,N_704,N_2188);
nor U9830 (N_9830,N_2852,N_2365);
nor U9831 (N_9831,N_4966,N_2951);
and U9832 (N_9832,N_1897,N_1583);
nand U9833 (N_9833,N_3672,N_1688);
or U9834 (N_9834,N_2119,N_1642);
and U9835 (N_9835,N_1461,N_455);
nor U9836 (N_9836,N_488,N_196);
nand U9837 (N_9837,N_4256,N_528);
or U9838 (N_9838,N_2140,N_15);
and U9839 (N_9839,N_3997,N_1861);
nor U9840 (N_9840,N_2178,N_3073);
nand U9841 (N_9841,N_1697,N_1801);
xnor U9842 (N_9842,N_253,N_4179);
nor U9843 (N_9843,N_2322,N_423);
nor U9844 (N_9844,N_2013,N_2174);
or U9845 (N_9845,N_36,N_4363);
nor U9846 (N_9846,N_886,N_1637);
and U9847 (N_9847,N_578,N_1299);
and U9848 (N_9848,N_1092,N_4371);
xor U9849 (N_9849,N_3944,N_2411);
xor U9850 (N_9850,N_1174,N_2554);
xor U9851 (N_9851,N_1113,N_4462);
nand U9852 (N_9852,N_2882,N_2913);
nand U9853 (N_9853,N_2054,N_2033);
or U9854 (N_9854,N_1461,N_3183);
nand U9855 (N_9855,N_2861,N_3747);
and U9856 (N_9856,N_4052,N_3932);
nor U9857 (N_9857,N_1276,N_2947);
or U9858 (N_9858,N_4825,N_4789);
nor U9859 (N_9859,N_4839,N_3580);
or U9860 (N_9860,N_1579,N_2440);
and U9861 (N_9861,N_1780,N_2324);
and U9862 (N_9862,N_2398,N_1596);
nand U9863 (N_9863,N_611,N_3348);
or U9864 (N_9864,N_2745,N_1072);
and U9865 (N_9865,N_740,N_4859);
xnor U9866 (N_9866,N_1679,N_4080);
and U9867 (N_9867,N_3421,N_2068);
nor U9868 (N_9868,N_3878,N_4337);
or U9869 (N_9869,N_3707,N_1714);
and U9870 (N_9870,N_4070,N_1610);
nand U9871 (N_9871,N_1355,N_1279);
and U9872 (N_9872,N_2413,N_1903);
xor U9873 (N_9873,N_4331,N_2241);
or U9874 (N_9874,N_4433,N_3542);
nand U9875 (N_9875,N_58,N_583);
or U9876 (N_9876,N_3317,N_2070);
nand U9877 (N_9877,N_3031,N_1495);
nand U9878 (N_9878,N_2270,N_4507);
nand U9879 (N_9879,N_3541,N_4572);
nor U9880 (N_9880,N_598,N_1394);
nor U9881 (N_9881,N_4215,N_768);
xor U9882 (N_9882,N_2479,N_2048);
and U9883 (N_9883,N_4188,N_3118);
nor U9884 (N_9884,N_2047,N_1517);
or U9885 (N_9885,N_1474,N_4179);
and U9886 (N_9886,N_1373,N_4147);
nand U9887 (N_9887,N_2716,N_3036);
xor U9888 (N_9888,N_3776,N_554);
and U9889 (N_9889,N_3247,N_3602);
nand U9890 (N_9890,N_2068,N_3029);
and U9891 (N_9891,N_3528,N_902);
and U9892 (N_9892,N_2571,N_1581);
nand U9893 (N_9893,N_3142,N_4162);
and U9894 (N_9894,N_531,N_2783);
and U9895 (N_9895,N_4801,N_4725);
and U9896 (N_9896,N_4563,N_1161);
nand U9897 (N_9897,N_3746,N_486);
or U9898 (N_9898,N_2655,N_600);
nor U9899 (N_9899,N_2383,N_564);
xnor U9900 (N_9900,N_94,N_2991);
or U9901 (N_9901,N_3310,N_2123);
xnor U9902 (N_9902,N_605,N_1520);
nand U9903 (N_9903,N_1718,N_3772);
nand U9904 (N_9904,N_2882,N_505);
nor U9905 (N_9905,N_2910,N_2379);
nor U9906 (N_9906,N_611,N_4979);
xor U9907 (N_9907,N_459,N_240);
and U9908 (N_9908,N_3001,N_1081);
nor U9909 (N_9909,N_3184,N_16);
xnor U9910 (N_9910,N_2831,N_4611);
xnor U9911 (N_9911,N_4204,N_3053);
and U9912 (N_9912,N_2496,N_1911);
and U9913 (N_9913,N_1505,N_787);
and U9914 (N_9914,N_1937,N_2678);
nor U9915 (N_9915,N_1052,N_3523);
nor U9916 (N_9916,N_4584,N_1321);
nor U9917 (N_9917,N_4058,N_523);
and U9918 (N_9918,N_871,N_4860);
xnor U9919 (N_9919,N_1307,N_4459);
and U9920 (N_9920,N_1714,N_4115);
or U9921 (N_9921,N_2880,N_2121);
and U9922 (N_9922,N_3594,N_4219);
nor U9923 (N_9923,N_747,N_2179);
xnor U9924 (N_9924,N_2617,N_1545);
nand U9925 (N_9925,N_3526,N_1565);
nor U9926 (N_9926,N_1714,N_2212);
nand U9927 (N_9927,N_822,N_2425);
nand U9928 (N_9928,N_3008,N_1649);
or U9929 (N_9929,N_55,N_1130);
and U9930 (N_9930,N_3794,N_3387);
nand U9931 (N_9931,N_1968,N_481);
or U9932 (N_9932,N_3994,N_2175);
nand U9933 (N_9933,N_2836,N_4401);
and U9934 (N_9934,N_1881,N_1983);
nor U9935 (N_9935,N_2102,N_102);
and U9936 (N_9936,N_907,N_175);
or U9937 (N_9937,N_1745,N_3091);
nor U9938 (N_9938,N_1627,N_123);
nor U9939 (N_9939,N_3124,N_2266);
nor U9940 (N_9940,N_3259,N_2148);
nand U9941 (N_9941,N_1274,N_4509);
nand U9942 (N_9942,N_715,N_1499);
nand U9943 (N_9943,N_660,N_677);
xor U9944 (N_9944,N_2713,N_3801);
and U9945 (N_9945,N_166,N_3346);
nand U9946 (N_9946,N_3852,N_451);
nand U9947 (N_9947,N_2707,N_1251);
xor U9948 (N_9948,N_3685,N_3552);
nor U9949 (N_9949,N_1299,N_419);
nor U9950 (N_9950,N_3297,N_1809);
nor U9951 (N_9951,N_3027,N_903);
xnor U9952 (N_9952,N_1253,N_3599);
nor U9953 (N_9953,N_1552,N_1536);
xor U9954 (N_9954,N_4773,N_4023);
or U9955 (N_9955,N_4887,N_642);
and U9956 (N_9956,N_1585,N_3652);
nand U9957 (N_9957,N_4181,N_714);
nand U9958 (N_9958,N_1114,N_1662);
xnor U9959 (N_9959,N_4540,N_4537);
nand U9960 (N_9960,N_4670,N_4747);
or U9961 (N_9961,N_4046,N_1985);
or U9962 (N_9962,N_400,N_4104);
and U9963 (N_9963,N_2498,N_685);
nand U9964 (N_9964,N_1136,N_4298);
and U9965 (N_9965,N_3190,N_2594);
nand U9966 (N_9966,N_3922,N_272);
and U9967 (N_9967,N_256,N_4902);
nor U9968 (N_9968,N_2148,N_1752);
nor U9969 (N_9969,N_1194,N_459);
or U9970 (N_9970,N_317,N_723);
or U9971 (N_9971,N_1579,N_623);
xor U9972 (N_9972,N_678,N_3503);
xnor U9973 (N_9973,N_1797,N_3325);
or U9974 (N_9974,N_3194,N_4060);
and U9975 (N_9975,N_3635,N_2043);
nor U9976 (N_9976,N_4607,N_567);
nor U9977 (N_9977,N_558,N_745);
and U9978 (N_9978,N_43,N_3956);
nor U9979 (N_9979,N_3347,N_1956);
xnor U9980 (N_9980,N_2775,N_3683);
nand U9981 (N_9981,N_3114,N_2612);
xnor U9982 (N_9982,N_1821,N_4409);
xor U9983 (N_9983,N_2595,N_3386);
xor U9984 (N_9984,N_4331,N_3638);
nand U9985 (N_9985,N_2280,N_806);
nor U9986 (N_9986,N_1553,N_365);
nor U9987 (N_9987,N_4274,N_4886);
or U9988 (N_9988,N_4618,N_2493);
xnor U9989 (N_9989,N_24,N_2945);
or U9990 (N_9990,N_821,N_587);
nor U9991 (N_9991,N_4189,N_828);
nand U9992 (N_9992,N_3891,N_1485);
and U9993 (N_9993,N_26,N_2384);
or U9994 (N_9994,N_2962,N_740);
and U9995 (N_9995,N_2795,N_3554);
xor U9996 (N_9996,N_1374,N_3931);
nor U9997 (N_9997,N_1437,N_1497);
and U9998 (N_9998,N_3277,N_3122);
and U9999 (N_9999,N_2852,N_1245);
nand UO_0 (O_0,N_9783,N_7777);
nor UO_1 (O_1,N_6848,N_7467);
and UO_2 (O_2,N_9849,N_7095);
xor UO_3 (O_3,N_9173,N_7134);
xnor UO_4 (O_4,N_8443,N_8761);
nand UO_5 (O_5,N_6564,N_6123);
or UO_6 (O_6,N_9210,N_7807);
or UO_7 (O_7,N_9579,N_5260);
or UO_8 (O_8,N_6771,N_9196);
nor UO_9 (O_9,N_7945,N_6670);
nand UO_10 (O_10,N_8398,N_8454);
nor UO_11 (O_11,N_9933,N_9735);
nand UO_12 (O_12,N_7229,N_7489);
nand UO_13 (O_13,N_8850,N_8215);
nor UO_14 (O_14,N_6589,N_8199);
and UO_15 (O_15,N_7495,N_9571);
nor UO_16 (O_16,N_8086,N_6256);
or UO_17 (O_17,N_7233,N_5342);
and UO_18 (O_18,N_9823,N_9494);
xor UO_19 (O_19,N_9772,N_8827);
and UO_20 (O_20,N_8462,N_5554);
nor UO_21 (O_21,N_7916,N_6028);
or UO_22 (O_22,N_8137,N_7282);
or UO_23 (O_23,N_9851,N_6209);
and UO_24 (O_24,N_9737,N_8779);
xnor UO_25 (O_25,N_6737,N_7108);
nor UO_26 (O_26,N_7917,N_8097);
or UO_27 (O_27,N_8396,N_9180);
nand UO_28 (O_28,N_5625,N_7124);
and UO_29 (O_29,N_6794,N_6756);
xnor UO_30 (O_30,N_9288,N_9685);
and UO_31 (O_31,N_7260,N_8860);
nor UO_32 (O_32,N_8116,N_5467);
nand UO_33 (O_33,N_5209,N_8213);
and UO_34 (O_34,N_9816,N_8889);
or UO_35 (O_35,N_7724,N_6269);
or UO_36 (O_36,N_9322,N_6039);
xnor UO_37 (O_37,N_8969,N_6132);
xnor UO_38 (O_38,N_6268,N_8715);
or UO_39 (O_39,N_8266,N_5419);
nand UO_40 (O_40,N_5519,N_8988);
and UO_41 (O_41,N_8432,N_8301);
nand UO_42 (O_42,N_8660,N_8845);
or UO_43 (O_43,N_8773,N_6533);
xnor UO_44 (O_44,N_5032,N_7771);
xnor UO_45 (O_45,N_9666,N_6480);
xnor UO_46 (O_46,N_9682,N_9371);
nand UO_47 (O_47,N_8930,N_6705);
xor UO_48 (O_48,N_8236,N_5992);
or UO_49 (O_49,N_7283,N_8746);
xnor UO_50 (O_50,N_9044,N_7276);
or UO_51 (O_51,N_6647,N_5296);
and UO_52 (O_52,N_9214,N_9502);
nor UO_53 (O_53,N_8562,N_5488);
or UO_54 (O_54,N_5479,N_9527);
nor UO_55 (O_55,N_8849,N_7364);
nand UO_56 (O_56,N_5060,N_6286);
nand UO_57 (O_57,N_7319,N_6747);
or UO_58 (O_58,N_7429,N_6566);
or UO_59 (O_59,N_8110,N_8856);
or UO_60 (O_60,N_8305,N_5168);
nor UO_61 (O_61,N_6287,N_7119);
or UO_62 (O_62,N_8468,N_8232);
and UO_63 (O_63,N_9123,N_9340);
nor UO_64 (O_64,N_8571,N_5264);
nor UO_65 (O_65,N_8934,N_8203);
nor UO_66 (O_66,N_8322,N_5427);
and UO_67 (O_67,N_8308,N_8494);
or UO_68 (O_68,N_5784,N_8261);
or UO_69 (O_69,N_9576,N_7605);
and UO_70 (O_70,N_5319,N_9319);
nand UO_71 (O_71,N_5336,N_5098);
or UO_72 (O_72,N_9108,N_5478);
nand UO_73 (O_73,N_8575,N_8388);
and UO_74 (O_74,N_9402,N_5019);
nand UO_75 (O_75,N_7372,N_7047);
nand UO_76 (O_76,N_6746,N_7991);
or UO_77 (O_77,N_6248,N_5258);
and UO_78 (O_78,N_6847,N_6278);
and UO_79 (O_79,N_5562,N_8258);
or UO_80 (O_80,N_5146,N_7543);
or UO_81 (O_81,N_8582,N_9528);
xor UO_82 (O_82,N_8231,N_6522);
xnor UO_83 (O_83,N_9374,N_6651);
nor UO_84 (O_84,N_8502,N_6327);
nor UO_85 (O_85,N_7726,N_5266);
xnor UO_86 (O_86,N_8688,N_9820);
nor UO_87 (O_87,N_9827,N_8723);
and UO_88 (O_88,N_8159,N_5603);
xnor UO_89 (O_89,N_6546,N_7506);
or UO_90 (O_90,N_9852,N_6553);
or UO_91 (O_91,N_8573,N_5181);
nand UO_92 (O_92,N_6141,N_9657);
and UO_93 (O_93,N_9891,N_9395);
nand UO_94 (O_94,N_9648,N_5800);
nor UO_95 (O_95,N_8354,N_7510);
nor UO_96 (O_96,N_5775,N_6816);
nand UO_97 (O_97,N_5681,N_8346);
nand UO_98 (O_98,N_7426,N_7740);
and UO_99 (O_99,N_8880,N_7598);
nand UO_100 (O_100,N_8712,N_7719);
or UO_101 (O_101,N_5429,N_9093);
nor UO_102 (O_102,N_8531,N_5579);
xor UO_103 (O_103,N_9638,N_7413);
or UO_104 (O_104,N_8523,N_7066);
and UO_105 (O_105,N_7897,N_7511);
nand UO_106 (O_106,N_5069,N_7599);
or UO_107 (O_107,N_6795,N_7321);
or UO_108 (O_108,N_5668,N_5398);
and UO_109 (O_109,N_9581,N_8138);
or UO_110 (O_110,N_8057,N_7383);
nor UO_111 (O_111,N_8903,N_7035);
nor UO_112 (O_112,N_5552,N_5542);
nand UO_113 (O_113,N_8430,N_6215);
and UO_114 (O_114,N_6012,N_5107);
and UO_115 (O_115,N_8557,N_9751);
and UO_116 (O_116,N_6359,N_7353);
nor UO_117 (O_117,N_6375,N_9197);
xnor UO_118 (O_118,N_9013,N_5437);
and UO_119 (O_119,N_8153,N_8998);
nor UO_120 (O_120,N_6017,N_7361);
or UO_121 (O_121,N_7018,N_8777);
nor UO_122 (O_122,N_6512,N_9138);
xnor UO_123 (O_123,N_8947,N_7278);
and UO_124 (O_124,N_6184,N_5269);
nor UO_125 (O_125,N_5178,N_5307);
or UO_126 (O_126,N_5555,N_7985);
nand UO_127 (O_127,N_9854,N_7877);
and UO_128 (O_128,N_9904,N_6629);
nand UO_129 (O_129,N_9635,N_9667);
nor UO_130 (O_130,N_9895,N_6750);
nand UO_131 (O_131,N_7316,N_8371);
xnor UO_132 (O_132,N_8657,N_7631);
and UO_133 (O_133,N_8599,N_8074);
nor UO_134 (O_134,N_7459,N_9928);
nand UO_135 (O_135,N_8942,N_9015);
nor UO_136 (O_136,N_9315,N_5637);
nor UO_137 (O_137,N_5163,N_5829);
and UO_138 (O_138,N_7126,N_8264);
xnor UO_139 (O_139,N_7268,N_7038);
nor UO_140 (O_140,N_9177,N_8940);
xnor UO_141 (O_141,N_6621,N_7349);
and UO_142 (O_142,N_7000,N_9894);
or UO_143 (O_143,N_6718,N_8931);
or UO_144 (O_144,N_5950,N_5027);
or UO_145 (O_145,N_5983,N_7552);
and UO_146 (O_146,N_7781,N_8379);
xnor UO_147 (O_147,N_6446,N_7017);
xor UO_148 (O_148,N_7325,N_6097);
or UO_149 (O_149,N_7892,N_8616);
nand UO_150 (O_150,N_5566,N_5255);
nor UO_151 (O_151,N_8710,N_9716);
or UO_152 (O_152,N_8944,N_9232);
or UO_153 (O_153,N_6971,N_9194);
nand UO_154 (O_154,N_7711,N_5638);
nand UO_155 (O_155,N_6473,N_8742);
or UO_156 (O_156,N_5687,N_8185);
nand UO_157 (O_157,N_7527,N_8709);
xnor UO_158 (O_158,N_9313,N_9719);
or UO_159 (O_159,N_7910,N_8395);
xnor UO_160 (O_160,N_8771,N_9726);
nand UO_161 (O_161,N_6901,N_7259);
nor UO_162 (O_162,N_5219,N_8209);
nor UO_163 (O_163,N_8149,N_9411);
nand UO_164 (O_164,N_9375,N_5618);
xnor UO_165 (O_165,N_8971,N_8658);
or UO_166 (O_166,N_8578,N_7405);
nand UO_167 (O_167,N_9385,N_8267);
and UO_168 (O_168,N_6314,N_5104);
or UO_169 (O_169,N_6585,N_5725);
nand UO_170 (O_170,N_6265,N_6875);
xnor UO_171 (O_171,N_7439,N_7295);
xnor UO_172 (O_172,N_6103,N_8525);
and UO_173 (O_173,N_5564,N_5626);
or UO_174 (O_174,N_8839,N_6685);
or UO_175 (O_175,N_7257,N_5058);
nor UO_176 (O_176,N_9048,N_7672);
and UO_177 (O_177,N_7125,N_5030);
xor UO_178 (O_178,N_8281,N_9830);
and UO_179 (O_179,N_5330,N_6069);
xnor UO_180 (O_180,N_7773,N_5135);
nand UO_181 (O_181,N_7064,N_9506);
and UO_182 (O_182,N_8999,N_6145);
or UO_183 (O_183,N_7694,N_5007);
nand UO_184 (O_184,N_5623,N_7576);
nand UO_185 (O_185,N_6385,N_7216);
xor UO_186 (O_186,N_9591,N_9547);
nand UO_187 (O_187,N_6174,N_5537);
nor UO_188 (O_188,N_9961,N_7201);
or UO_189 (O_189,N_6457,N_7468);
or UO_190 (O_190,N_5823,N_7195);
or UO_191 (O_191,N_8581,N_8418);
or UO_192 (O_192,N_9066,N_5981);
and UO_193 (O_193,N_7953,N_6923);
xnor UO_194 (O_194,N_9717,N_9788);
and UO_195 (O_195,N_9062,N_8592);
nand UO_196 (O_196,N_5409,N_6187);
nand UO_197 (O_197,N_8191,N_5943);
nor UO_198 (O_198,N_5432,N_6855);
nand UO_199 (O_199,N_9223,N_7148);
or UO_200 (O_200,N_6300,N_6603);
or UO_201 (O_201,N_8897,N_8996);
nor UO_202 (O_202,N_7692,N_7374);
xor UO_203 (O_203,N_7399,N_5352);
xor UO_204 (O_204,N_9865,N_9909);
and UO_205 (O_205,N_5177,N_6760);
nor UO_206 (O_206,N_7084,N_8019);
or UO_207 (O_207,N_7474,N_5571);
xor UO_208 (O_208,N_6736,N_6404);
or UO_209 (O_209,N_5796,N_6530);
nor UO_210 (O_210,N_8133,N_8604);
xnor UO_211 (O_211,N_6462,N_9713);
and UO_212 (O_212,N_6351,N_5561);
nand UO_213 (O_213,N_6600,N_8207);
or UO_214 (O_214,N_9723,N_7752);
nor UO_215 (O_215,N_7322,N_8275);
nand UO_216 (O_216,N_6360,N_6606);
and UO_217 (O_217,N_9388,N_9773);
and UO_218 (O_218,N_6073,N_8627);
nand UO_219 (O_219,N_7291,N_9991);
xnor UO_220 (O_220,N_7835,N_9099);
nand UO_221 (O_221,N_9111,N_8725);
nor UO_222 (O_222,N_9507,N_5522);
xnor UO_223 (O_223,N_8680,N_6284);
xor UO_224 (O_224,N_8912,N_9003);
xor UO_225 (O_225,N_9623,N_7859);
and UO_226 (O_226,N_9328,N_5344);
and UO_227 (O_227,N_5746,N_8026);
xor UO_228 (O_228,N_7805,N_5397);
nor UO_229 (O_229,N_5938,N_9668);
nor UO_230 (O_230,N_8227,N_9834);
or UO_231 (O_231,N_8458,N_7833);
nand UO_232 (O_232,N_9777,N_6988);
nor UO_233 (O_233,N_5878,N_5227);
nand UO_234 (O_234,N_8561,N_6658);
nand UO_235 (O_235,N_9530,N_7267);
nand UO_236 (O_236,N_8666,N_9208);
xor UO_237 (O_237,N_9779,N_9963);
xnor UO_238 (O_238,N_7443,N_5204);
or UO_239 (O_239,N_5837,N_8062);
or UO_240 (O_240,N_7002,N_6762);
xnor UO_241 (O_241,N_8645,N_5463);
and UO_242 (O_242,N_8326,N_6406);
nor UO_243 (O_243,N_5399,N_8685);
nor UO_244 (O_244,N_6147,N_5317);
or UO_245 (O_245,N_6733,N_7465);
xor UO_246 (O_246,N_5291,N_5117);
xor UO_247 (O_247,N_6008,N_9833);
nor UO_248 (O_248,N_9286,N_9573);
or UO_249 (O_249,N_7785,N_7435);
nand UO_250 (O_250,N_9290,N_6180);
nor UO_251 (O_251,N_8948,N_7493);
and UO_252 (O_252,N_8800,N_9642);
and UO_253 (O_253,N_8318,N_5541);
nor UO_254 (O_254,N_9239,N_6241);
xnor UO_255 (O_255,N_9094,N_7749);
and UO_256 (O_256,N_5088,N_5734);
and UO_257 (O_257,N_9131,N_7022);
and UO_258 (O_258,N_7544,N_5528);
and UO_259 (O_259,N_5029,N_8123);
nor UO_260 (O_260,N_5639,N_9250);
or UO_261 (O_261,N_6144,N_8529);
and UO_262 (O_262,N_8718,N_9059);
or UO_263 (O_263,N_5842,N_8390);
or UO_264 (O_264,N_9978,N_5076);
nor UO_265 (O_265,N_8960,N_6197);
nor UO_266 (O_266,N_8050,N_9531);
nand UO_267 (O_267,N_8155,N_8358);
xor UO_268 (O_268,N_9790,N_7850);
nand UO_269 (O_269,N_5224,N_7779);
nor UO_270 (O_270,N_8134,N_8569);
nor UO_271 (O_271,N_8887,N_6015);
nand UO_272 (O_272,N_8970,N_5388);
and UO_273 (O_273,N_5436,N_6934);
nor UO_274 (O_274,N_5935,N_7469);
nand UO_275 (O_275,N_6263,N_7354);
and UO_276 (O_276,N_7901,N_6995);
xnor UO_277 (O_277,N_8438,N_6087);
nand UO_278 (O_278,N_6191,N_5780);
nand UO_279 (O_279,N_8896,N_6018);
nand UO_280 (O_280,N_8141,N_6161);
nor UO_281 (O_281,N_9391,N_7554);
xor UO_282 (O_282,N_6814,N_6458);
nand UO_283 (O_283,N_8894,N_7614);
and UO_284 (O_284,N_6790,N_9121);
or UO_285 (O_285,N_7876,N_6518);
nor UO_286 (O_286,N_5661,N_7989);
nand UO_287 (O_287,N_7896,N_7592);
nor UO_288 (O_288,N_6099,N_9162);
or UO_289 (O_289,N_8670,N_5169);
or UO_290 (O_290,N_9349,N_7100);
xor UO_291 (O_291,N_8778,N_8882);
or UO_292 (O_292,N_6997,N_5290);
or UO_293 (O_293,N_6500,N_7816);
nor UO_294 (O_294,N_8169,N_7478);
and UO_295 (O_295,N_8898,N_7856);
and UO_296 (O_296,N_9417,N_9167);
nor UO_297 (O_297,N_7546,N_5894);
or UO_298 (O_298,N_9526,N_7998);
and UO_299 (O_299,N_9333,N_5414);
and UO_300 (O_300,N_5699,N_8362);
xnor UO_301 (O_301,N_9207,N_6235);
nand UO_302 (O_302,N_6569,N_7776);
nor UO_303 (O_303,N_6975,N_9699);
xor UO_304 (O_304,N_5621,N_9932);
and UO_305 (O_305,N_5184,N_5162);
nand UO_306 (O_306,N_8600,N_6973);
xor UO_307 (O_307,N_6739,N_5675);
nand UO_308 (O_308,N_7457,N_7667);
xnor UO_309 (O_309,N_6489,N_7331);
nor UO_310 (O_310,N_5691,N_5462);
and UO_311 (O_311,N_5951,N_7815);
xor UO_312 (O_312,N_5103,N_8437);
or UO_313 (O_313,N_9996,N_7674);
and UO_314 (O_314,N_9873,N_8423);
and UO_315 (O_315,N_8586,N_5836);
nand UO_316 (O_316,N_7738,N_6730);
and UO_317 (O_317,N_6166,N_5695);
nand UO_318 (O_318,N_7230,N_9169);
xnor UO_319 (O_319,N_7098,N_6767);
nor UO_320 (O_320,N_8349,N_9786);
nand UO_321 (O_321,N_6834,N_8551);
xnor UO_322 (O_322,N_8117,N_6939);
or UO_323 (O_323,N_6806,N_7220);
nand UO_324 (O_324,N_5111,N_8309);
xnor UO_325 (O_325,N_8373,N_5359);
nand UO_326 (O_326,N_9944,N_9263);
and UO_327 (O_327,N_9559,N_7450);
or UO_328 (O_328,N_5267,N_9273);
and UO_329 (O_329,N_5171,N_7867);
or UO_330 (O_330,N_6797,N_5712);
nand UO_331 (O_331,N_5387,N_7822);
nand UO_332 (O_332,N_8406,N_5971);
nand UO_333 (O_333,N_5788,N_9413);
nor UO_334 (O_334,N_5892,N_9255);
xor UO_335 (O_335,N_9578,N_5349);
and UO_336 (O_336,N_7551,N_9951);
and UO_337 (O_337,N_7109,N_8279);
or UO_338 (O_338,N_5927,N_6267);
nor UO_339 (O_339,N_8489,N_6067);
nor UO_340 (O_340,N_7303,N_8467);
and UO_341 (O_341,N_5670,N_6216);
and UO_342 (O_342,N_9275,N_8517);
or UO_343 (O_343,N_6148,N_8703);
or UO_344 (O_344,N_7913,N_9874);
nand UO_345 (O_345,N_7863,N_6239);
nand UO_346 (O_346,N_8350,N_6565);
nor UO_347 (O_347,N_6993,N_5074);
nand UO_348 (O_348,N_9082,N_8165);
nor UO_349 (O_349,N_5294,N_6996);
or UO_350 (O_350,N_5790,N_9143);
nand UO_351 (O_351,N_9549,N_5608);
nor UO_352 (O_352,N_7957,N_5254);
xnor UO_353 (O_353,N_5080,N_6125);
nand UO_354 (O_354,N_6143,N_9317);
and UO_355 (O_355,N_8714,N_5934);
and UO_356 (O_356,N_5191,N_9922);
nor UO_357 (O_357,N_7590,N_5116);
xor UO_358 (O_358,N_6292,N_6656);
nand UO_359 (O_359,N_5082,N_8615);
xnor UO_360 (O_360,N_8507,N_6998);
and UO_361 (O_361,N_5186,N_6571);
nor UO_362 (O_362,N_6904,N_7209);
nor UO_363 (O_363,N_5509,N_8828);
or UO_364 (O_364,N_7149,N_9761);
nor UO_365 (O_365,N_6021,N_7128);
nor UO_366 (O_366,N_6649,N_9246);
or UO_367 (O_367,N_8324,N_9989);
nor UO_368 (O_368,N_7828,N_8164);
xnor UO_369 (O_369,N_9681,N_6529);
and UO_370 (O_370,N_9534,N_6042);
xnor UO_371 (O_371,N_5018,N_7794);
nor UO_372 (O_372,N_9660,N_9198);
nor UO_373 (O_373,N_7410,N_6341);
and UO_374 (O_374,N_5979,N_9014);
nand UO_375 (O_375,N_7171,N_9536);
nor UO_376 (O_376,N_5277,N_9728);
xnor UO_377 (O_377,N_7241,N_6786);
xor UO_378 (O_378,N_8935,N_8296);
nand UO_379 (O_379,N_8484,N_5010);
xor UO_380 (O_380,N_7427,N_8422);
and UO_381 (O_381,N_8696,N_6418);
or UO_382 (O_382,N_9278,N_8793);
nor UO_383 (O_383,N_9064,N_8862);
nand UO_384 (O_384,N_6802,N_5716);
xor UO_385 (O_385,N_6772,N_7697);
nand UO_386 (O_386,N_6727,N_9353);
and UO_387 (O_387,N_7366,N_5354);
and UO_388 (O_388,N_6009,N_8152);
nand UO_389 (O_389,N_5331,N_9347);
nor UO_390 (O_390,N_5764,N_9204);
xor UO_391 (O_391,N_5744,N_5001);
and UO_392 (O_392,N_6865,N_6006);
xor UO_393 (O_393,N_8424,N_7763);
nand UO_394 (O_394,N_6678,N_8020);
and UO_395 (O_395,N_7003,N_8994);
or UO_396 (O_396,N_5651,N_8452);
and UO_397 (O_397,N_8810,N_9881);
nand UO_398 (O_398,N_9613,N_9752);
nor UO_399 (O_399,N_8799,N_8351);
nand UO_400 (O_400,N_7327,N_7226);
xor UO_401 (O_401,N_9125,N_9425);
nor UO_402 (O_402,N_5249,N_6837);
xnor UO_403 (O_403,N_8105,N_5108);
or UO_404 (O_404,N_8391,N_7351);
xor UO_405 (O_405,N_5361,N_9035);
nand UO_406 (O_406,N_7416,N_8878);
nand UO_407 (O_407,N_7541,N_5962);
xor UO_408 (O_408,N_5487,N_9176);
xnor UO_409 (O_409,N_8389,N_9351);
nor UO_410 (O_410,N_9965,N_6506);
or UO_411 (O_411,N_8697,N_8824);
nand UO_412 (O_412,N_5396,N_9342);
xnor UO_413 (O_413,N_7415,N_6635);
and UO_414 (O_414,N_8353,N_5762);
and UO_415 (O_415,N_8447,N_5990);
and UO_416 (O_416,N_8536,N_5589);
nor UO_417 (O_417,N_8114,N_5248);
or UO_418 (O_418,N_7836,N_5025);
or UO_419 (O_419,N_5070,N_6773);
or UO_420 (O_420,N_8633,N_5891);
and UO_421 (O_421,N_7296,N_7509);
nand UO_422 (O_422,N_5014,N_9563);
and UO_423 (O_423,N_6376,N_7869);
xor UO_424 (O_424,N_5413,N_6349);
or UO_425 (O_425,N_6504,N_5631);
nor UO_426 (O_426,N_5506,N_6270);
xor UO_427 (O_427,N_8817,N_7471);
nand UO_428 (O_428,N_6403,N_6048);
or UO_429 (O_429,N_8417,N_8776);
or UO_430 (O_430,N_5289,N_5480);
nor UO_431 (O_431,N_9089,N_9508);
nor UO_432 (O_432,N_5718,N_9810);
nor UO_433 (O_433,N_7646,N_5996);
and UO_434 (O_434,N_8890,N_8440);
nand UO_435 (O_435,N_9046,N_8166);
xnor UO_436 (O_436,N_5306,N_5926);
nor UO_437 (O_437,N_8115,N_5126);
or UO_438 (O_438,N_6430,N_6306);
xnor UO_439 (O_439,N_7845,N_9252);
xor UO_440 (O_440,N_6610,N_5558);
and UO_441 (O_441,N_5524,N_9566);
and UO_442 (O_442,N_7213,N_5874);
xor UO_443 (O_443,N_7961,N_6684);
and UO_444 (O_444,N_8108,N_5987);
xor UO_445 (O_445,N_8588,N_5050);
and UO_446 (O_446,N_8366,N_9809);
and UO_447 (O_447,N_5355,N_6254);
or UO_448 (O_448,N_8510,N_9267);
or UO_449 (O_449,N_8472,N_9864);
and UO_450 (O_450,N_9597,N_5031);
xor UO_451 (O_451,N_9758,N_5508);
nor UO_452 (O_452,N_9858,N_7715);
and UO_453 (O_453,N_8087,N_6260);
or UO_454 (O_454,N_9495,N_7787);
xnor UO_455 (O_455,N_8073,N_9714);
and UO_456 (O_456,N_9546,N_5949);
nand UO_457 (O_457,N_9750,N_7995);
and UO_458 (O_458,N_5977,N_9696);
and UO_459 (O_459,N_6877,N_9447);
nor UO_460 (O_460,N_7540,N_7602);
nand UO_461 (O_461,N_9535,N_9725);
nand UO_462 (O_462,N_5363,N_5520);
or UO_463 (O_463,N_9557,N_9945);
nand UO_464 (O_464,N_7580,N_6829);
or UO_465 (O_465,N_9988,N_5362);
and UO_466 (O_466,N_9952,N_9017);
or UO_467 (O_467,N_6022,N_8984);
or UO_468 (O_468,N_8919,N_9670);
nand UO_469 (O_469,N_8297,N_7420);
or UO_470 (O_470,N_8084,N_5000);
or UO_471 (O_471,N_8727,N_7640);
or UO_472 (O_472,N_6780,N_8478);
xnor UO_473 (O_473,N_6242,N_8566);
nor UO_474 (O_474,N_6671,N_5513);
xor UO_475 (O_475,N_9977,N_7363);
or UO_476 (O_476,N_6987,N_7205);
xnor UO_477 (O_477,N_8997,N_7442);
or UO_478 (O_478,N_9747,N_9363);
nor UO_479 (O_479,N_7811,N_8242);
and UO_480 (O_480,N_8330,N_7504);
and UO_481 (O_481,N_6507,N_5348);
or UO_482 (O_482,N_8687,N_7051);
and UO_483 (O_483,N_6538,N_9456);
nor UO_484 (O_484,N_6648,N_5701);
nand UO_485 (O_485,N_5075,N_5905);
or UO_486 (O_486,N_8435,N_9439);
or UO_487 (O_487,N_6843,N_7880);
nand UO_488 (O_488,N_5740,N_8345);
xnor UO_489 (O_489,N_6870,N_9229);
nand UO_490 (O_490,N_6702,N_9856);
or UO_491 (O_491,N_9541,N_7750);
nand UO_492 (O_492,N_5028,N_6915);
nand UO_493 (O_493,N_6893,N_7446);
nor UO_494 (O_494,N_6159,N_7755);
nor UO_495 (O_495,N_9020,N_5866);
or UO_496 (O_496,N_9754,N_5474);
nor UO_497 (O_497,N_5011,N_7742);
nand UO_498 (O_498,N_9480,N_5105);
nor UO_499 (O_499,N_6395,N_5741);
and UO_500 (O_500,N_5335,N_6298);
and UO_501 (O_501,N_7834,N_8005);
nand UO_502 (O_502,N_6700,N_7846);
nor UO_503 (O_503,N_7021,N_9599);
or UO_504 (O_504,N_5672,N_9485);
and UO_505 (O_505,N_6461,N_8642);
and UO_506 (O_506,N_7315,N_5123);
and UO_507 (O_507,N_9513,N_7829);
or UO_508 (O_508,N_7183,N_6983);
and UO_509 (O_509,N_8426,N_5145);
or UO_510 (O_510,N_7492,N_9692);
and UO_511 (O_511,N_8397,N_6070);
or UO_512 (O_512,N_8719,N_8081);
nor UO_513 (O_513,N_9329,N_8542);
or UO_514 (O_514,N_6886,N_6778);
nor UO_515 (O_515,N_8690,N_9918);
nand UO_516 (O_516,N_8598,N_9806);
xor UO_517 (O_517,N_8061,N_5641);
and UO_518 (O_518,N_9216,N_9585);
xnor UO_519 (O_519,N_9938,N_6568);
and UO_520 (O_520,N_7094,N_6689);
nor UO_521 (O_521,N_8950,N_7406);
xor UO_522 (O_522,N_6981,N_6057);
nor UO_523 (O_523,N_6472,N_8549);
and UO_524 (O_524,N_9624,N_9796);
xor UO_525 (O_525,N_9943,N_6692);
xor UO_526 (O_526,N_5925,N_8991);
nand UO_527 (O_527,N_9913,N_8590);
nand UO_528 (O_528,N_6146,N_9980);
nor UO_529 (O_529,N_6397,N_9112);
and UO_530 (O_530,N_8886,N_7110);
xor UO_531 (O_531,N_6475,N_6768);
nand UO_532 (O_532,N_8289,N_7984);
xnor UO_533 (O_533,N_9056,N_8752);
nor UO_534 (O_534,N_8744,N_8623);
nor UO_535 (O_535,N_7538,N_6181);
nand UO_536 (O_536,N_6523,N_5507);
or UO_537 (O_537,N_5565,N_5611);
or UO_538 (O_538,N_9946,N_5898);
nor UO_539 (O_539,N_6019,N_9344);
xor UO_540 (O_540,N_8954,N_5311);
nor UO_541 (O_541,N_7861,N_8338);
xnor UO_542 (O_542,N_5980,N_9600);
xnor UO_543 (O_543,N_6101,N_6672);
nand UO_544 (O_544,N_7431,N_8804);
or UO_545 (O_545,N_8869,N_8023);
xor UO_546 (O_546,N_7765,N_8728);
xnor UO_547 (O_547,N_6043,N_6226);
nand UO_548 (O_548,N_8501,N_7871);
nor UO_549 (O_549,N_9958,N_9191);
nand UO_550 (O_550,N_8796,N_6832);
nand UO_551 (O_551,N_8235,N_9440);
or UO_552 (O_552,N_7797,N_8365);
xor UO_553 (O_553,N_7408,N_5609);
nor UO_554 (O_554,N_8790,N_7612);
nor UO_555 (O_555,N_9798,N_5262);
or UO_556 (O_556,N_6743,N_9669);
nand UO_557 (O_557,N_9900,N_7981);
nand UO_558 (O_558,N_6305,N_9791);
xor UO_559 (O_559,N_7947,N_5583);
nand UO_560 (O_560,N_8433,N_9802);
nor UO_561 (O_561,N_8593,N_6563);
or UO_562 (O_562,N_7369,N_7786);
nor UO_563 (O_563,N_7454,N_6251);
xor UO_564 (O_564,N_8323,N_5867);
or UO_565 (O_565,N_5821,N_8131);
or UO_566 (O_566,N_5465,N_7117);
xnor UO_567 (O_567,N_7934,N_6119);
nand UO_568 (O_568,N_7542,N_8533);
nand UO_569 (O_569,N_9259,N_6954);
nand UO_570 (O_570,N_8080,N_7687);
nor UO_571 (O_571,N_5833,N_7398);
nand UO_572 (O_572,N_9023,N_8981);
and UO_573 (O_573,N_6366,N_8363);
and UO_574 (O_574,N_9588,N_7419);
nor UO_575 (O_575,N_8361,N_5459);
nor UO_576 (O_576,N_5662,N_5131);
or UO_577 (O_577,N_8993,N_8967);
and UO_578 (O_578,N_5752,N_7914);
and UO_579 (O_579,N_5346,N_6902);
xor UO_580 (O_580,N_7448,N_6989);
xor UO_581 (O_581,N_8273,N_6626);
xor UO_582 (O_582,N_8001,N_7272);
and UO_583 (O_583,N_9462,N_8069);
or UO_584 (O_584,N_7091,N_6336);
or UO_585 (O_585,N_9985,N_5855);
xnor UO_586 (O_586,N_9415,N_7270);
or UO_587 (O_587,N_9866,N_8337);
nor UO_588 (O_588,N_5659,N_7801);
or UO_589 (O_589,N_6082,N_5669);
xnor UO_590 (O_590,N_8722,N_6390);
or UO_591 (O_591,N_8949,N_5286);
xor UO_592 (O_592,N_8120,N_6978);
xor UO_593 (O_593,N_8126,N_7654);
or UO_594 (O_594,N_6370,N_7887);
xnor UO_595 (O_595,N_6266,N_8737);
and UO_596 (O_596,N_8254,N_9962);
xnor UO_597 (O_597,N_7502,N_6081);
xnor UO_598 (O_598,N_8527,N_5057);
xnor UO_599 (O_599,N_5605,N_8000);
and UO_600 (O_600,N_8585,N_7340);
or UO_601 (O_601,N_9200,N_9970);
and UO_602 (O_602,N_9763,N_8769);
nand UO_603 (O_603,N_9760,N_8927);
or UO_604 (O_604,N_8492,N_9925);
nand UO_605 (O_605,N_6830,N_6963);
xor UO_606 (O_606,N_6804,N_6346);
and UO_607 (O_607,N_8014,N_8701);
or UO_608 (O_608,N_9244,N_7891);
and UO_609 (O_609,N_6272,N_5195);
xor UO_610 (O_610,N_6435,N_5930);
or UO_611 (O_611,N_8922,N_7154);
nand UO_612 (O_612,N_9929,N_6167);
and UO_613 (O_613,N_5339,N_8072);
nor UO_614 (O_614,N_5854,N_8076);
and UO_615 (O_615,N_9247,N_7147);
nand UO_616 (O_616,N_6849,N_6770);
nor UO_617 (O_617,N_6495,N_9129);
and UO_618 (O_618,N_8698,N_8332);
nand UO_619 (O_619,N_6127,N_9381);
nor UO_620 (O_620,N_6367,N_5481);
or UO_621 (O_621,N_6405,N_9924);
xor UO_622 (O_622,N_5160,N_8135);
nor UO_623 (O_623,N_7087,N_7875);
and UO_624 (O_624,N_6044,N_6204);
nor UO_625 (O_625,N_9935,N_6195);
nand UO_626 (O_626,N_6463,N_5222);
xor UO_627 (O_627,N_5004,N_5646);
and UO_628 (O_628,N_7210,N_7472);
nor UO_629 (O_629,N_7432,N_6655);
nor UO_630 (O_630,N_7900,N_7460);
nand UO_631 (O_631,N_6642,N_9323);
and UO_632 (O_632,N_9033,N_5149);
or UO_633 (O_633,N_8056,N_6699);
or UO_634 (O_634,N_5440,N_9915);
nand UO_635 (O_635,N_7182,N_9853);
nor UO_636 (O_636,N_7935,N_8461);
nor UO_637 (O_637,N_9283,N_7952);
or UO_638 (O_638,N_7744,N_7425);
xnor UO_639 (O_639,N_7207,N_6482);
nor UO_640 (O_640,N_6502,N_9756);
nor UO_641 (O_641,N_8290,N_9299);
nand UO_642 (O_642,N_6907,N_5736);
nand UO_643 (O_643,N_7378,N_7754);
nand UO_644 (O_644,N_8870,N_6961);
and UO_645 (O_645,N_8033,N_6706);
and UO_646 (O_646,N_5984,N_9110);
and UO_647 (O_647,N_8833,N_9912);
and UO_648 (O_648,N_7737,N_6484);
or UO_649 (O_649,N_7421,N_6368);
nor UO_650 (O_650,N_6499,N_6679);
and UO_651 (O_651,N_5830,N_9358);
xor UO_652 (O_652,N_9042,N_9262);
nor UO_653 (O_653,N_8004,N_7564);
nand UO_654 (O_654,N_7299,N_6944);
nand UO_655 (O_655,N_8786,N_7655);
xnor UO_656 (O_656,N_5619,N_8808);
xor UO_657 (O_657,N_7508,N_9540);
or UO_658 (O_658,N_8780,N_9293);
nand UO_659 (O_659,N_6299,N_8847);
or UO_660 (O_660,N_9616,N_5472);
nor UO_661 (O_661,N_7127,N_6691);
nand UO_662 (O_662,N_8622,N_8781);
xor UO_663 (O_663,N_7650,N_8902);
or UO_664 (O_664,N_6659,N_5496);
nor UO_665 (O_665,N_8568,N_7057);
or UO_666 (O_666,N_7758,N_8522);
or UO_667 (O_667,N_6320,N_8920);
and UO_668 (O_668,N_7573,N_8634);
nor UO_669 (O_669,N_9225,N_6527);
and UO_670 (O_670,N_7774,N_5203);
nand UO_671 (O_671,N_8002,N_9457);
nand UO_672 (O_672,N_5077,N_5580);
and UO_673 (O_673,N_5393,N_8317);
or UO_674 (O_674,N_9618,N_5857);
or UO_675 (O_675,N_9813,N_7168);
nor UO_676 (O_676,N_5406,N_7888);
nand UO_677 (O_677,N_7618,N_5747);
and UO_678 (O_678,N_6861,N_7946);
or UO_679 (O_679,N_6005,N_5827);
nor UO_680 (O_680,N_6796,N_5553);
and UO_681 (O_681,N_9704,N_9749);
or UO_682 (O_682,N_9677,N_7885);
and UO_683 (O_683,N_9748,N_7707);
and UO_684 (O_684,N_8720,N_5758);
or UO_685 (O_685,N_5719,N_9300);
and UO_686 (O_686,N_8060,N_9927);
xnor UO_687 (O_687,N_5815,N_9795);
xnor UO_688 (O_688,N_9568,N_9930);
and UO_689 (O_689,N_7456,N_6783);
or UO_690 (O_690,N_7525,N_6152);
xor UO_691 (O_691,N_5805,N_7761);
and UO_692 (O_692,N_6126,N_6941);
nor UO_693 (O_693,N_7924,N_7054);
nand UO_694 (O_694,N_9867,N_7996);
and UO_695 (O_695,N_9399,N_7868);
and UO_696 (O_696,N_9238,N_8321);
or UO_697 (O_697,N_8343,N_6213);
xor UO_698 (O_698,N_6131,N_6665);
nand UO_699 (O_699,N_5710,N_9320);
nand UO_700 (O_700,N_5415,N_6520);
or UO_701 (O_701,N_9258,N_9684);
and UO_702 (O_702,N_7476,N_6850);
nor UO_703 (O_703,N_7937,N_9794);
and UO_704 (O_704,N_7256,N_7008);
and UO_705 (O_705,N_8916,N_9153);
or UO_706 (O_706,N_6844,N_5148);
and UO_707 (O_707,N_5645,N_8884);
nor UO_708 (O_708,N_6609,N_7417);
nand UO_709 (O_709,N_9040,N_5375);
and UO_710 (O_710,N_9672,N_5584);
nor UO_711 (O_711,N_6304,N_9145);
or UO_712 (O_712,N_5383,N_6836);
xor UO_713 (O_713,N_9947,N_8537);
and UO_714 (O_714,N_5771,N_9742);
and UO_715 (O_715,N_5792,N_7607);
or UO_716 (O_716,N_6090,N_7653);
xnor UO_717 (O_717,N_6838,N_8918);
or UO_718 (O_718,N_7122,N_9161);
xor UO_719 (O_719,N_8589,N_7648);
or UO_720 (O_720,N_6443,N_5494);
nor UO_721 (O_721,N_7014,N_7645);
and UO_722 (O_722,N_7516,N_5514);
nor UO_723 (O_723,N_9316,N_6232);
or UO_724 (O_724,N_7379,N_7277);
and UO_725 (O_725,N_9957,N_6862);
xor UO_726 (O_726,N_5256,N_9201);
xnor UO_727 (O_727,N_6535,N_5642);
nor UO_728 (O_728,N_6010,N_5159);
and UO_729 (O_729,N_7572,N_9118);
nor UO_730 (O_730,N_6644,N_9390);
xnor UO_731 (O_731,N_7265,N_5709);
or UO_732 (O_732,N_5380,N_5840);
xnor UO_733 (O_733,N_7809,N_9632);
nor UO_734 (O_734,N_7284,N_6542);
xor UO_735 (O_735,N_5114,N_7804);
nand UO_736 (O_736,N_6697,N_5121);
and UO_737 (O_737,N_5883,N_5353);
or UO_738 (O_738,N_5134,N_9680);
and UO_739 (O_739,N_8130,N_8090);
nand UO_740 (O_740,N_6183,N_7466);
xnor UO_741 (O_741,N_5982,N_5975);
nand UO_742 (O_742,N_6333,N_7865);
and UO_743 (O_743,N_7960,N_9807);
and UO_744 (O_744,N_5220,N_8956);
xnor UO_745 (O_745,N_6434,N_6866);
xnor UO_746 (O_746,N_6449,N_6912);
nor UO_747 (O_747,N_8671,N_9107);
and UO_748 (O_748,N_6608,N_6719);
or UO_749 (O_749,N_8140,N_8584);
nor UO_750 (O_750,N_5677,N_7800);
nor UO_751 (O_751,N_7926,N_7644);
and UO_752 (O_752,N_7958,N_8039);
xnor UO_753 (O_753,N_8606,N_8731);
or UO_754 (O_754,N_9501,N_9377);
nor UO_755 (O_755,N_8837,N_9026);
nand UO_756 (O_756,N_6348,N_5343);
or UO_757 (O_757,N_5865,N_5819);
or UO_758 (O_758,N_9165,N_5377);
nand UO_759 (O_759,N_5721,N_5818);
and UO_760 (O_760,N_5456,N_7445);
or UO_761 (O_761,N_5213,N_9661);
and UO_762 (O_762,N_5902,N_5092);
or UO_763 (O_763,N_5644,N_7453);
or UO_764 (O_764,N_9734,N_8803);
nand UO_765 (O_765,N_9671,N_7718);
xnor UO_766 (O_766,N_7422,N_6076);
and UO_767 (O_767,N_9181,N_9355);
nand UO_768 (O_768,N_5652,N_9832);
and UO_769 (O_769,N_6122,N_5688);
and UO_770 (O_770,N_5132,N_9269);
and UO_771 (O_771,N_7940,N_5500);
nand UO_772 (O_772,N_9679,N_5316);
or UO_773 (O_773,N_8612,N_5686);
nand UO_774 (O_774,N_5968,N_8407);
nand UO_775 (O_775,N_5850,N_6433);
and UO_776 (O_776,N_5613,N_5431);
nor UO_777 (O_777,N_6815,N_8758);
nand UO_778 (O_778,N_5382,N_5443);
or UO_779 (O_779,N_6384,N_5140);
nand UO_780 (O_780,N_8142,N_6052);
nor UO_781 (O_781,N_8875,N_8764);
nor UO_782 (O_782,N_5392,N_7062);
nand UO_783 (O_783,N_6809,N_9718);
nor UO_784 (O_784,N_7521,N_8691);
nand UO_785 (O_785,N_5706,N_8621);
and UO_786 (O_786,N_5274,N_5188);
nand UO_787 (O_787,N_6675,N_7083);
and UO_788 (O_788,N_7882,N_5461);
nand UO_789 (O_789,N_5664,N_7751);
xor UO_790 (O_790,N_8809,N_6663);
or UO_791 (O_791,N_8319,N_7342);
nor UO_792 (O_792,N_6620,N_5281);
and UO_793 (O_793,N_9078,N_6466);
nor UO_794 (O_794,N_9512,N_8286);
nor UO_795 (O_795,N_6558,N_6785);
and UO_796 (O_796,N_7263,N_6918);
or UO_797 (O_797,N_5851,N_5997);
and UO_798 (O_798,N_8907,N_6534);
nand UO_799 (O_799,N_7915,N_7853);
or UO_800 (O_800,N_8190,N_9338);
nor UO_801 (O_801,N_6258,N_7073);
and UO_802 (O_802,N_9289,N_6554);
xor UO_803 (O_803,N_7772,N_8831);
and UO_804 (O_804,N_9553,N_7015);
nand UO_805 (O_805,N_8486,N_7536);
xor UO_806 (O_806,N_6496,N_9675);
and UO_807 (O_807,N_7392,N_6238);
nand UO_808 (O_808,N_6986,N_9006);
nor UO_809 (O_809,N_5152,N_9292);
or UO_810 (O_810,N_8619,N_6420);
nand UO_811 (O_811,N_5732,N_8179);
or UO_812 (O_812,N_6460,N_8876);
nand UO_813 (O_813,N_8180,N_5323);
or UO_814 (O_814,N_9147,N_6483);
or UO_815 (O_815,N_7596,N_7235);
nand UO_816 (O_816,N_9073,N_7889);
or UO_817 (O_817,N_5726,N_9722);
or UO_818 (O_818,N_6325,N_9720);
nor UO_819 (O_819,N_5606,N_8552);
or UO_820 (O_820,N_8933,N_8444);
or UO_821 (O_821,N_8243,N_8618);
nand UO_822 (O_822,N_8654,N_9203);
nor UO_823 (O_823,N_5612,N_9736);
xnor UO_824 (O_824,N_7178,N_7052);
nand UO_825 (O_825,N_7463,N_9464);
xnor UO_826 (O_826,N_7732,N_9926);
nor UO_827 (O_827,N_7630,N_9793);
nor UO_828 (O_828,N_5705,N_6088);
nor UO_829 (O_829,N_8370,N_8754);
xnor UO_830 (O_830,N_9206,N_7044);
or UO_831 (O_831,N_8846,N_7548);
xor UO_832 (O_832,N_5482,N_6567);
nand UO_833 (O_833,N_6481,N_6826);
nand UO_834 (O_834,N_9997,N_5728);
xnor UO_835 (O_835,N_7533,N_9438);
xnor UO_836 (O_836,N_7290,N_7515);
xor UO_837 (O_837,N_5090,N_6025);
nand UO_838 (O_838,N_5887,N_7324);
nor UO_839 (O_839,N_7582,N_7255);
or UO_840 (O_840,N_7994,N_6079);
nand UO_841 (O_841,N_9228,N_6488);
xor UO_842 (O_842,N_7414,N_5557);
nor UO_843 (O_843,N_7623,N_5628);
nor UO_844 (O_844,N_6262,N_8964);
nand UO_845 (O_845,N_9421,N_8481);
nor UO_846 (O_846,N_5787,N_9400);
nor UO_847 (O_847,N_8476,N_9998);
or UO_848 (O_848,N_8962,N_6196);
xnor UO_849 (O_849,N_6026,N_7486);
nand UO_850 (O_850,N_9039,N_7006);
or UO_851 (O_851,N_6003,N_5067);
or UO_852 (O_852,N_5278,N_8538);
xor UO_853 (O_853,N_5089,N_5965);
nand UO_854 (O_854,N_8524,N_6083);
and UO_855 (O_855,N_8506,N_8233);
nand UO_856 (O_856,N_9036,N_5051);
nor UO_857 (O_857,N_7335,N_5693);
nor UO_858 (O_858,N_7371,N_8410);
nor UO_859 (O_859,N_6639,N_5757);
nand UO_860 (O_860,N_8348,N_9448);
nand UO_861 (O_861,N_5877,N_5530);
nand UO_862 (O_862,N_9960,N_5896);
nand UO_863 (O_863,N_7600,N_5073);
and UO_864 (O_864,N_9132,N_5216);
and UO_865 (O_865,N_6176,N_8577);
xnor UO_866 (O_866,N_7424,N_8649);
or UO_867 (O_867,N_5791,N_5947);
xor UO_868 (O_868,N_5326,N_7135);
xor UO_869 (O_869,N_8535,N_8664);
and UO_870 (O_870,N_8157,N_9373);
xnor UO_871 (O_871,N_8352,N_8470);
and UO_872 (O_872,N_5420,N_8450);
nand UO_873 (O_873,N_7196,N_9301);
xor UO_874 (O_874,N_9921,N_9814);
nand UO_875 (O_875,N_6051,N_6095);
nor UO_876 (O_876,N_5422,N_6835);
nand UO_877 (O_877,N_8013,N_7012);
xor UO_878 (O_878,N_8936,N_8943);
or UO_879 (O_879,N_7317,N_9151);
or UO_880 (O_880,N_7187,N_7441);
and UO_881 (O_881,N_9542,N_6399);
and UO_882 (O_882,N_6245,N_9324);
nor UO_883 (O_883,N_7795,N_7962);
nor UO_884 (O_884,N_9172,N_6597);
nor UO_885 (O_885,N_9733,N_7227);
nand UO_886 (O_886,N_9759,N_8576);
and UO_887 (O_887,N_8342,N_6810);
and UO_888 (O_888,N_6974,N_8904);
nand UO_889 (O_889,N_6704,N_6261);
and UO_890 (O_890,N_9170,N_6091);
nand UO_891 (O_891,N_9074,N_9942);
and UO_892 (O_892,N_6874,N_8419);
or UO_893 (O_893,N_9226,N_5239);
or UO_894 (O_894,N_9739,N_7485);
and UO_895 (O_895,N_6050,N_6764);
nand UO_896 (O_896,N_8413,N_7499);
and UO_897 (O_897,N_7034,N_8255);
nand UO_898 (O_898,N_7237,N_9028);
and UO_899 (O_899,N_8198,N_7997);
or UO_900 (O_900,N_6058,N_7238);
nand UO_901 (O_901,N_5253,N_7503);
or UO_902 (O_902,N_6402,N_5733);
nand UO_903 (O_903,N_5110,N_8145);
xnor UO_904 (O_904,N_6948,N_5371);
or UO_905 (O_905,N_7568,N_6930);
nand UO_906 (O_906,N_9484,N_7610);
nor UO_907 (O_907,N_5229,N_5164);
nand UO_908 (O_908,N_7451,N_5430);
xnor UO_909 (O_909,N_7156,N_9590);
xnor UO_910 (O_910,N_7959,N_6839);
or UO_911 (O_911,N_7903,N_6602);
nor UO_912 (O_912,N_5955,N_9309);
and UO_913 (O_913,N_6416,N_7684);
or UO_914 (O_914,N_5279,N_8699);
xor UO_915 (O_915,N_8730,N_7905);
or UO_916 (O_916,N_7860,N_8224);
xor UO_917 (O_917,N_5526,N_6717);
nand UO_918 (O_918,N_8037,N_5994);
xor UO_919 (O_919,N_8204,N_9800);
nand UO_920 (O_920,N_5425,N_5534);
nor UO_921 (O_921,N_8036,N_6919);
xor UO_922 (O_922,N_8819,N_9785);
nor UO_923 (O_923,N_8978,N_5826);
or UO_924 (O_924,N_5270,N_5231);
or UO_925 (O_925,N_6813,N_6661);
xnor UO_926 (O_926,N_9157,N_6616);
nor UO_927 (O_927,N_6316,N_9803);
or UO_928 (O_928,N_7713,N_6863);
nand UO_929 (O_929,N_8556,N_9466);
and UO_930 (O_930,N_6133,N_8059);
nand UO_931 (O_931,N_6757,N_8250);
nor UO_932 (O_932,N_8403,N_5379);
nor UO_933 (O_933,N_5663,N_5401);
nand UO_934 (O_934,N_9314,N_9478);
xor UO_935 (O_935,N_6623,N_7992);
nand UO_936 (O_936,N_7462,N_5903);
and UO_937 (O_937,N_6129,N_9156);
nor UO_938 (O_938,N_5308,N_6641);
or UO_939 (O_939,N_7753,N_7832);
and UO_940 (O_940,N_7532,N_7565);
or UO_941 (O_941,N_7616,N_7025);
nand UO_942 (O_942,N_5370,N_8716);
or UO_943 (O_943,N_9474,N_9767);
xnor UO_944 (O_944,N_6725,N_8613);
xor UO_945 (O_945,N_9029,N_5864);
nand UO_946 (O_946,N_5853,N_9243);
xnor UO_947 (O_947,N_8146,N_9022);
or UO_948 (O_948,N_8214,N_9847);
or UO_949 (O_949,N_9133,N_7314);
nand UO_950 (O_950,N_7673,N_9135);
nand UO_951 (O_951,N_9504,N_6652);
xnor UO_952 (O_952,N_9562,N_6169);
and UO_953 (O_953,N_6959,N_7566);
and UO_954 (O_954,N_6929,N_5586);
nor UO_955 (O_955,N_9248,N_5199);
or UO_956 (O_956,N_8068,N_8184);
nand UO_957 (O_957,N_6885,N_7107);
xnor UO_958 (O_958,N_6636,N_6096);
xor UO_959 (O_959,N_5748,N_6259);
xor UO_960 (O_960,N_5109,N_8183);
xnor UO_961 (O_961,N_7387,N_6887);
nor UO_962 (O_962,N_5529,N_6734);
or UO_963 (O_963,N_8749,N_9879);
and UO_964 (O_964,N_6960,N_8088);
xor UO_965 (O_965,N_9394,N_7103);
and UO_966 (O_966,N_5208,N_7556);
nor UO_967 (O_967,N_5304,N_6253);
nand UO_968 (O_968,N_6102,N_5384);
or UO_969 (O_969,N_7385,N_5005);
nor UO_970 (O_970,N_7247,N_8830);
or UO_971 (O_971,N_9337,N_5717);
xnor UO_972 (O_972,N_7136,N_8821);
or UO_973 (O_973,N_7367,N_5189);
and UO_974 (O_974,N_6198,N_7433);
nand UO_975 (O_975,N_5045,N_6357);
nor UO_976 (O_976,N_8823,N_6992);
xnor UO_977 (O_977,N_6549,N_6598);
or UO_978 (O_978,N_9975,N_5647);
or UO_979 (O_979,N_8464,N_6289);
or UO_980 (O_980,N_8244,N_6172);
xnor UO_981 (O_981,N_5475,N_7939);
nor UO_982 (O_982,N_9631,N_7949);
or UO_983 (O_983,N_9937,N_8661);
xor UO_984 (O_984,N_8293,N_8665);
nand UO_985 (O_985,N_6696,N_5426);
or UO_986 (O_986,N_5447,N_7562);
nand UO_987 (O_987,N_5417,N_9034);
and UO_988 (O_988,N_5094,N_7180);
nand UO_989 (O_989,N_5908,N_5763);
or UO_990 (O_990,N_7292,N_6340);
or UO_991 (O_991,N_5044,N_7971);
and UO_992 (O_992,N_8883,N_5081);
nand UO_993 (O_993,N_8740,N_8228);
xnor UO_994 (O_994,N_6444,N_7248);
and UO_995 (O_995,N_6698,N_5096);
nand UO_996 (O_996,N_5793,N_9298);
and UO_997 (O_997,N_7261,N_9209);
nor UO_998 (O_998,N_9237,N_6163);
or UO_999 (O_999,N_7203,N_5958);
or UO_1000 (O_1000,N_8811,N_9475);
nand UO_1001 (O_1001,N_5678,N_5366);
nor UO_1002 (O_1002,N_7320,N_6324);
nor UO_1003 (O_1003,N_8836,N_9686);
or UO_1004 (O_1004,N_8482,N_8054);
nor UO_1005 (O_1005,N_7192,N_8456);
nor UO_1006 (O_1006,N_8640,N_5989);
and UO_1007 (O_1007,N_6999,N_8528);
xor UO_1008 (O_1008,N_9346,N_9326);
xnor UO_1009 (O_1009,N_9369,N_5237);
nand UO_1010 (O_1010,N_6157,N_5141);
nor UO_1011 (O_1011,N_8448,N_5671);
nand UO_1012 (O_1012,N_9755,N_5424);
xnor UO_1013 (O_1013,N_6142,N_8044);
or UO_1014 (O_1014,N_6151,N_8302);
nand UO_1015 (O_1015,N_7153,N_5329);
xnor UO_1016 (O_1016,N_9412,N_6190);
or UO_1017 (O_1017,N_9215,N_6358);
and UO_1018 (O_1018,N_6720,N_8291);
nor UO_1019 (O_1019,N_9649,N_7225);
nand UO_1020 (O_1020,N_7799,N_5122);
and UO_1021 (O_1021,N_5454,N_8844);
nor UO_1022 (O_1022,N_8067,N_5458);
xor UO_1023 (O_1023,N_5421,N_6840);
or UO_1024 (O_1024,N_5054,N_8911);
nor UO_1025 (O_1025,N_5567,N_5974);
nand UO_1026 (O_1026,N_5912,N_9857);
nor UO_1027 (O_1027,N_8385,N_6828);
nand UO_1028 (O_1028,N_7668,N_8774);
or UO_1029 (O_1029,N_5442,N_6230);
or UO_1030 (O_1030,N_5808,N_5629);
and UO_1031 (O_1031,N_5696,N_7980);
or UO_1032 (O_1032,N_7031,N_9828);
xnor UO_1033 (O_1033,N_7709,N_5812);
or UO_1034 (O_1034,N_8979,N_9359);
and UO_1035 (O_1035,N_7185,N_5347);
xor UO_1036 (O_1036,N_6742,N_8441);
xor UO_1037 (O_1037,N_5410,N_6509);
and UO_1038 (O_1038,N_5265,N_6425);
nand UO_1039 (O_1039,N_6326,N_9117);
xnor UO_1040 (O_1040,N_5450,N_9659);
xor UO_1041 (O_1041,N_9986,N_8545);
and UO_1042 (O_1042,N_9905,N_9936);
nand UO_1043 (O_1043,N_9305,N_6712);
or UO_1044 (O_1044,N_6541,N_8863);
or UO_1045 (O_1045,N_8867,N_7588);
xnor UO_1046 (O_1046,N_7403,N_9981);
xor UO_1047 (O_1047,N_7788,N_5360);
and UO_1048 (O_1048,N_9451,N_9306);
nor UO_1049 (O_1049,N_9075,N_8368);
nand UO_1050 (O_1050,N_6846,N_8614);
nand UO_1051 (O_1051,N_9903,N_9189);
nand UO_1052 (O_1052,N_8514,N_5438);
and UO_1053 (O_1053,N_9159,N_9651);
nor UO_1054 (O_1054,N_9764,N_8865);
or UO_1055 (O_1055,N_8043,N_5139);
nand UO_1056 (O_1056,N_7377,N_9976);
or UO_1057 (O_1057,N_8595,N_6414);
xnor UO_1058 (O_1058,N_6423,N_8439);
or UO_1059 (O_1059,N_8854,N_7685);
xor UO_1060 (O_1060,N_9297,N_9840);
nor UO_1061 (O_1061,N_8055,N_6991);
and UO_1062 (O_1062,N_6153,N_7177);
xnor UO_1063 (O_1063,N_5801,N_5215);
or UO_1064 (O_1064,N_8763,N_6508);
nor UO_1065 (O_1065,N_6503,N_8574);
nor UO_1066 (O_1066,N_6588,N_9397);
nor UO_1067 (O_1067,N_9069,N_8905);
and UO_1068 (O_1068,N_6295,N_5797);
or UO_1069 (O_1069,N_8974,N_7162);
or UO_1070 (O_1070,N_7111,N_8172);
nand UO_1071 (O_1071,N_8269,N_6497);
xnor UO_1072 (O_1072,N_8929,N_6250);
xnor UO_1073 (O_1073,N_9304,N_8900);
xnor UO_1074 (O_1074,N_9769,N_6014);
xnor UO_1075 (O_1075,N_7483,N_7181);
and UO_1076 (O_1076,N_6693,N_5960);
nor UO_1077 (O_1077,N_6976,N_7855);
and UO_1078 (O_1078,N_8491,N_6905);
and UO_1079 (O_1079,N_7526,N_6913);
or UO_1080 (O_1080,N_8700,N_8768);
and UO_1081 (O_1081,N_6781,N_5043);
and UO_1082 (O_1082,N_7919,N_5674);
and UO_1083 (O_1083,N_9876,N_5283);
nand UO_1084 (O_1084,N_9995,N_5634);
and UO_1085 (O_1085,N_9656,N_7964);
xor UO_1086 (O_1086,N_8765,N_8431);
nor UO_1087 (O_1087,N_5310,N_9310);
xnor UO_1088 (O_1088,N_9010,N_6676);
and UO_1089 (O_1089,N_9605,N_9134);
or UO_1090 (O_1090,N_6908,N_8866);
nor UO_1091 (O_1091,N_7090,N_5276);
or UO_1092 (O_1092,N_6206,N_9640);
xnor UO_1093 (O_1093,N_9091,N_5835);
xnor UO_1094 (O_1094,N_6765,N_5911);
xnor UO_1095 (O_1095,N_7904,N_7714);
xnor UO_1096 (O_1096,N_5280,N_5233);
nand UO_1097 (O_1097,N_6412,N_9465);
and UO_1098 (O_1098,N_9594,N_8558);
or UO_1099 (O_1099,N_6900,N_7373);
or UO_1100 (O_1100,N_7308,N_8806);
and UO_1101 (O_1101,N_8705,N_5499);
xnor UO_1102 (O_1102,N_5156,N_9055);
or UO_1103 (O_1103,N_8611,N_6407);
and UO_1104 (O_1104,N_5617,N_6759);
nand UO_1105 (O_1105,N_9572,N_9030);
nor UO_1106 (O_1106,N_7727,N_5999);
and UO_1107 (O_1107,N_7118,N_7329);
or UO_1108 (O_1108,N_7577,N_8583);
and UO_1109 (O_1109,N_9520,N_6798);
or UO_1110 (O_1110,N_9444,N_7444);
nand UO_1111 (O_1111,N_9382,N_9627);
nand UO_1112 (O_1112,N_6592,N_9979);
nor UO_1113 (O_1113,N_9429,N_5785);
or UO_1114 (O_1114,N_5038,N_8334);
or UO_1115 (O_1115,N_6646,N_7817);
and UO_1116 (O_1116,N_6803,N_8331);
nand UO_1117 (O_1117,N_6078,N_9916);
and UO_1118 (O_1118,N_6532,N_6189);
or UO_1119 (O_1119,N_5843,N_8683);
nor UO_1120 (O_1120,N_7473,N_6290);
nand UO_1121 (O_1121,N_8008,N_7622);
xnor UO_1122 (O_1122,N_5015,N_5033);
nor UO_1123 (O_1123,N_8151,N_9220);
or UO_1124 (O_1124,N_6066,N_8853);
xnor UO_1125 (O_1125,N_6873,N_7053);
nand UO_1126 (O_1126,N_7312,N_6972);
or UO_1127 (O_1127,N_7042,N_6222);
nand UO_1128 (O_1128,N_5907,N_9364);
and UO_1129 (O_1129,N_5445,N_5055);
or UO_1130 (O_1130,N_9569,N_7531);
or UO_1131 (O_1131,N_6118,N_5034);
and UO_1132 (O_1132,N_7986,N_9443);
or UO_1133 (O_1133,N_7132,N_7912);
nand UO_1134 (O_1134,N_8483,N_8729);
or UO_1135 (O_1135,N_8003,N_5180);
and UO_1136 (O_1136,N_8329,N_7251);
nand UO_1137 (O_1137,N_9430,N_6510);
xnor UO_1138 (O_1138,N_7242,N_7966);
or UO_1139 (O_1139,N_9969,N_9119);
nand UO_1140 (O_1140,N_9859,N_8792);
nor UO_1141 (O_1141,N_7619,N_7106);
and UO_1142 (O_1142,N_7368,N_9175);
or UO_1143 (O_1143,N_6454,N_5133);
nand UO_1144 (O_1144,N_5574,N_6208);
nor UO_1145 (O_1145,N_7092,N_8162);
or UO_1146 (O_1146,N_6000,N_7401);
nand UO_1147 (O_1147,N_9245,N_5825);
xnor UO_1148 (O_1148,N_9492,N_9518);
or UO_1149 (O_1149,N_5351,N_9948);
and UO_1150 (O_1150,N_5469,N_8629);
and UO_1151 (O_1151,N_6452,N_9277);
or UO_1152 (O_1152,N_6294,N_5400);
nor UO_1153 (O_1153,N_9136,N_5694);
or UO_1154 (O_1154,N_6323,N_9678);
xnor UO_1155 (O_1155,N_8938,N_8226);
and UO_1156 (O_1156,N_5312,N_6138);
nor UO_1157 (O_1157,N_8753,N_7206);
and UO_1158 (O_1158,N_5889,N_5587);
and UO_1159 (O_1159,N_9939,N_7902);
xor UO_1160 (O_1160,N_7933,N_6313);
xor UO_1161 (O_1161,N_5303,N_5200);
and UO_1162 (O_1162,N_9971,N_8208);
and UO_1163 (O_1163,N_8271,N_9431);
and UO_1164 (O_1164,N_7063,N_5803);
or UO_1165 (O_1165,N_7657,N_9780);
xor UO_1166 (O_1166,N_8066,N_8104);
and UO_1167 (O_1167,N_7488,N_5995);
nand UO_1168 (O_1168,N_8834,N_6859);
nor UO_1169 (O_1169,N_8855,N_8251);
and UO_1170 (O_1170,N_6925,N_8386);
xnor UO_1171 (O_1171,N_5372,N_6409);
or UO_1172 (O_1172,N_6137,N_6851);
nand UO_1173 (O_1173,N_8992,N_8229);
nand UO_1174 (O_1174,N_9387,N_8872);
nor UO_1175 (O_1175,N_7438,N_6957);
or UO_1176 (O_1176,N_7734,N_6888);
and UO_1177 (O_1177,N_5337,N_5112);
and UO_1178 (O_1178,N_7193,N_8017);
or UO_1179 (O_1179,N_8260,N_8843);
or UO_1180 (O_1180,N_8565,N_6459);
and UO_1181 (O_1181,N_7624,N_6024);
nor UO_1182 (O_1182,N_8651,N_6494);
nand UO_1183 (O_1183,N_5834,N_9193);
nand UO_1184 (O_1184,N_9630,N_8409);
nand UO_1185 (O_1185,N_8499,N_5125);
xor UO_1186 (O_1186,N_5101,N_7884);
nand UO_1187 (O_1187,N_7701,N_7231);
nor UO_1188 (O_1188,N_9919,N_7641);
nor UO_1189 (O_1189,N_6883,N_8223);
or UO_1190 (O_1190,N_9500,N_9450);
and UO_1191 (O_1191,N_5206,N_9334);
and UO_1192 (O_1192,N_8311,N_8101);
xor UO_1193 (O_1193,N_6513,N_7343);
and UO_1194 (O_1194,N_5923,N_6653);
xor UO_1195 (O_1195,N_9701,N_9449);
and UO_1196 (O_1196,N_6596,N_7879);
xor UO_1197 (O_1197,N_9461,N_7032);
nand UO_1198 (O_1198,N_7589,N_9653);
and UO_1199 (O_1199,N_9514,N_8732);
and UO_1200 (O_1200,N_6465,N_6068);
nand UO_1201 (O_1201,N_7825,N_7628);
and UO_1202 (O_1202,N_5610,N_6493);
nand UO_1203 (O_1203,N_9213,N_7626);
and UO_1204 (O_1204,N_9525,N_5035);
nor UO_1205 (O_1205,N_9423,N_9729);
or UO_1206 (O_1206,N_9144,N_6643);
xor UO_1207 (O_1207,N_6640,N_6867);
nand UO_1208 (O_1208,N_9380,N_5102);
xnor UO_1209 (O_1209,N_6227,N_6601);
or UO_1210 (O_1210,N_9992,N_8316);
nand UO_1211 (O_1211,N_9910,N_9109);
and UO_1212 (O_1212,N_6818,N_6424);
nand UO_1213 (O_1213,N_6124,N_8910);
nand UO_1214 (O_1214,N_7404,N_7050);
and UO_1215 (O_1215,N_7391,N_9544);
and UO_1216 (O_1216,N_6236,N_8280);
or UO_1217 (O_1217,N_6089,N_7769);
and UO_1218 (O_1218,N_6617,N_8733);
or UO_1219 (O_1219,N_9096,N_6139);
or UO_1220 (O_1220,N_8921,N_9265);
nand UO_1221 (O_1221,N_8797,N_5257);
xnor UO_1222 (O_1222,N_9521,N_7394);
nand UO_1223 (O_1223,N_9473,N_5404);
nand UO_1224 (O_1224,N_5768,N_6038);
nor UO_1225 (O_1225,N_8702,N_6769);
xor UO_1226 (O_1226,N_5314,N_6824);
xor UO_1227 (O_1227,N_6966,N_7150);
xnor UO_1228 (O_1228,N_5236,N_6618);
and UO_1229 (O_1229,N_9509,N_6744);
xnor UO_1230 (O_1230,N_5773,N_6940);
xnor UO_1231 (O_1231,N_6634,N_9537);
xor UO_1232 (O_1232,N_9920,N_8471);
nor UO_1233 (O_1233,N_5933,N_6293);
and UO_1234 (O_1234,N_8695,N_7729);
and UO_1235 (O_1235,N_7287,N_8504);
or UO_1236 (O_1236,N_7070,N_7928);
xor UO_1237 (O_1237,N_9990,N_8038);
or UO_1238 (O_1238,N_8957,N_8968);
and UO_1239 (O_1239,N_9116,N_7418);
nand UO_1240 (O_1240,N_9710,N_7505);
xor UO_1241 (O_1241,N_7033,N_9805);
xor UO_1242 (O_1242,N_6808,N_7144);
or UO_1243 (O_1243,N_5581,N_5405);
nor UO_1244 (O_1244,N_7096,N_5847);
and UO_1245 (O_1245,N_9860,N_7059);
and UO_1246 (O_1246,N_9776,N_8344);
nor UO_1247 (O_1247,N_8704,N_6577);
or UO_1248 (O_1248,N_6398,N_8336);
and UO_1249 (O_1249,N_5932,N_9184);
nand UO_1250 (O_1250,N_9602,N_9368);
and UO_1251 (O_1251,N_8519,N_8063);
nor UO_1252 (O_1252,N_9045,N_5635);
and UO_1253 (O_1253,N_6246,N_9254);
nor UO_1254 (O_1254,N_6551,N_8877);
nor UO_1255 (O_1255,N_7381,N_6111);
xnor UO_1256 (O_1256,N_7810,N_8168);
and UO_1257 (O_1257,N_8077,N_7883);
nand UO_1258 (O_1258,N_5751,N_8143);
and UO_1259 (O_1259,N_5988,N_9235);
and UO_1260 (O_1260,N_9829,N_6726);
nor UO_1261 (O_1261,N_8757,N_8473);
nand UO_1262 (O_1262,N_8333,N_9984);
and UO_1263 (O_1263,N_5909,N_6917);
nor UO_1264 (O_1264,N_8457,N_6871);
or UO_1265 (O_1265,N_6607,N_6381);
nand UO_1266 (O_1266,N_6920,N_7494);
nor UO_1267 (O_1267,N_8359,N_6799);
xnor UO_1268 (O_1268,N_5772,N_6531);
xor UO_1269 (O_1269,N_9515,N_7659);
or UO_1270 (O_1270,N_8802,N_6361);
or UO_1271 (O_1271,N_9953,N_8972);
or UO_1272 (O_1272,N_9647,N_5305);
nand UO_1273 (O_1273,N_7142,N_5838);
nor UO_1274 (O_1274,N_7840,N_5369);
nand UO_1275 (O_1275,N_7175,N_7269);
xnor UO_1276 (O_1276,N_5624,N_7274);
nor UO_1277 (O_1277,N_8031,N_6979);
nand UO_1278 (O_1278,N_8040,N_8818);
nand UO_1279 (O_1279,N_7518,N_9356);
or UO_1280 (O_1280,N_8983,N_5916);
and UO_1281 (O_1281,N_5546,N_9279);
xnor UO_1282 (O_1282,N_8990,N_6297);
nand UO_1283 (O_1283,N_5774,N_9987);
and UO_1284 (O_1284,N_5658,N_5046);
nand UO_1285 (O_1285,N_7872,N_5735);
and UO_1286 (O_1286,N_6117,N_8913);
or UO_1287 (O_1287,N_8427,N_6108);
nor UO_1288 (O_1288,N_6935,N_7490);
nand UO_1289 (O_1289,N_8641,N_9202);
nor UO_1290 (O_1290,N_8873,N_9804);
xor UO_1291 (O_1291,N_6001,N_5357);
nor UO_1292 (O_1292,N_6547,N_6953);
nor UO_1293 (O_1293,N_6787,N_7629);
xnor UO_1294 (O_1294,N_9959,N_7412);
xnor UO_1295 (O_1295,N_7561,N_6279);
nor UO_1296 (O_1296,N_9580,N_8567);
and UO_1297 (O_1297,N_6202,N_9318);
nor UO_1298 (O_1298,N_5511,N_7725);
or UO_1299 (O_1299,N_7131,N_5512);
nor UO_1300 (O_1300,N_5196,N_5954);
nor UO_1301 (O_1301,N_7487,N_6074);
xor UO_1302 (O_1302,N_7068,N_9884);
and UO_1303 (O_1303,N_5176,N_5945);
and UO_1304 (O_1304,N_6748,N_9517);
nand UO_1305 (O_1305,N_6487,N_6664);
nor UO_1306 (O_1306,N_7844,N_6694);
nand UO_1307 (O_1307,N_6624,N_7236);
and UO_1308 (O_1308,N_5525,N_6105);
or UO_1309 (O_1309,N_9251,N_6330);
nor UO_1310 (O_1310,N_7790,N_8194);
or UO_1311 (O_1311,N_7522,N_9564);
xnor UO_1312 (O_1312,N_7249,N_5952);
xor UO_1313 (O_1313,N_6895,N_9967);
or UO_1314 (O_1314,N_7080,N_8007);
nand UO_1315 (O_1315,N_6205,N_6779);
and UO_1316 (O_1316,N_7334,N_8544);
nand UO_1317 (O_1317,N_9614,N_5551);
or UO_1318 (O_1318,N_7976,N_6104);
and UO_1319 (O_1319,N_8205,N_7165);
or UO_1320 (O_1320,N_7748,N_8546);
nor UO_1321 (O_1321,N_9950,N_6422);
nand UO_1322 (O_1322,N_8783,N_5452);
and UO_1323 (O_1323,N_8150,N_7783);
and UO_1324 (O_1324,N_5723,N_7764);
nor UO_1325 (O_1325,N_9850,N_7625);
or UO_1326 (O_1326,N_8976,N_5386);
nor UO_1327 (O_1327,N_9280,N_6047);
nor UO_1328 (O_1328,N_7560,N_8505);
nand UO_1329 (O_1329,N_5918,N_6924);
xor UO_1330 (O_1330,N_5970,N_6175);
nand UO_1331 (O_1331,N_7601,N_8564);
xnor UO_1332 (O_1332,N_5556,N_8547);
nor UO_1333 (O_1333,N_6356,N_8453);
or UO_1334 (O_1334,N_6890,N_7146);
nand UO_1335 (O_1335,N_7024,N_8357);
nand UO_1336 (O_1336,N_8684,N_6982);
xnor UO_1337 (O_1337,N_9032,N_8295);
xor UO_1338 (O_1338,N_8405,N_8977);
xor UO_1339 (O_1339,N_8107,N_8859);
xor UO_1340 (O_1340,N_8047,N_5811);
or UO_1341 (O_1341,N_7710,N_6301);
nand UO_1342 (O_1342,N_7326,N_8539);
xor UO_1343 (O_1343,N_9441,N_7716);
or UO_1344 (O_1344,N_9097,N_8689);
and UO_1345 (O_1345,N_6595,N_9270);
xnor UO_1346 (O_1346,N_8526,N_5373);
or UO_1347 (O_1347,N_8374,N_8364);
and UO_1348 (O_1348,N_8734,N_9011);
and UO_1349 (O_1349,N_7613,N_7130);
nor UO_1350 (O_1350,N_8852,N_9875);
nand UO_1351 (O_1351,N_5548,N_5860);
xor UO_1352 (O_1352,N_9454,N_8113);
nand UO_1353 (O_1353,N_6707,N_8864);
nand UO_1354 (O_1354,N_8851,N_9178);
or UO_1355 (O_1355,N_9222,N_5468);
or UO_1356 (O_1356,N_6793,N_8377);
or UO_1357 (O_1357,N_5722,N_9543);
or UO_1358 (O_1358,N_9090,N_7043);
and UO_1359 (O_1359,N_5841,N_7559);
nand UO_1360 (O_1360,N_6853,N_9195);
nand UO_1361 (O_1361,N_6860,N_9266);
nand UO_1362 (O_1362,N_6470,N_8278);
or UO_1363 (O_1363,N_8085,N_5095);
xor UO_1364 (O_1364,N_7010,N_7636);
nor UO_1365 (O_1365,N_9687,N_6128);
nor UO_1366 (O_1366,N_5059,N_7918);
and UO_1367 (O_1367,N_6328,N_9689);
nand UO_1368 (O_1368,N_6436,N_8791);
nand UO_1369 (O_1369,N_7698,N_5846);
nand UO_1370 (O_1370,N_9715,N_5476);
and UO_1371 (O_1371,N_9993,N_7077);
nor UO_1372 (O_1372,N_8893,N_7818);
nor UO_1373 (O_1373,N_6612,N_9071);
xnor UO_1374 (O_1374,N_5590,N_9683);
xnor UO_1375 (O_1375,N_7682,N_5428);
nand UO_1376 (O_1376,N_6556,N_5673);
nand UO_1377 (O_1377,N_8384,N_6419);
nand UO_1378 (O_1378,N_7683,N_6910);
nor UO_1379 (O_1379,N_8294,N_8303);
xor UO_1380 (O_1380,N_6516,N_6632);
nor UO_1381 (O_1381,N_7252,N_9268);
xor UO_1382 (O_1382,N_5516,N_6914);
nand UO_1383 (O_1383,N_7239,N_5190);
and UO_1384 (O_1384,N_9738,N_7055);
nand UO_1385 (O_1385,N_6630,N_8376);
xor UO_1386 (O_1386,N_9160,N_5232);
or UO_1387 (O_1387,N_8075,N_5358);
nand UO_1388 (O_1388,N_5753,N_9914);
nor UO_1389 (O_1389,N_9824,N_8404);
or UO_1390 (O_1390,N_9016,N_5737);
nand UO_1391 (O_1391,N_5884,N_5592);
nor UO_1392 (O_1392,N_9907,N_7217);
nand UO_1393 (O_1393,N_9365,N_7569);
xnor UO_1394 (O_1394,N_7803,N_8249);
xnor UO_1395 (O_1395,N_7159,N_5570);
or UO_1396 (O_1396,N_5240,N_6355);
xor UO_1397 (O_1397,N_7250,N_9414);
and UO_1398 (O_1398,N_7827,N_7030);
xor UO_1399 (O_1399,N_5136,N_7428);
and UO_1400 (O_1400,N_8449,N_8360);
nor UO_1401 (O_1401,N_5704,N_7743);
xor UO_1402 (O_1402,N_5385,N_5175);
nand UO_1403 (O_1403,N_5991,N_9361);
and UO_1404 (O_1404,N_8161,N_6002);
nor UO_1405 (O_1405,N_9080,N_7411);
or UO_1406 (O_1406,N_8247,N_7011);
nor UO_1407 (O_1407,N_9148,N_6037);
nand UO_1408 (O_1408,N_6317,N_9625);
and UO_1409 (O_1409,N_6394,N_7830);
xor UO_1410 (O_1410,N_8313,N_5538);
nor UO_1411 (O_1411,N_7948,N_7155);
or UO_1412 (O_1412,N_7188,N_5147);
or UO_1413 (O_1413,N_5715,N_8591);
nor UO_1414 (O_1414,N_6899,N_6791);
nand UO_1415 (O_1415,N_5099,N_6949);
and UO_1416 (O_1416,N_7086,N_9533);
xnor UO_1417 (O_1417,N_7886,N_5020);
xnor UO_1418 (O_1418,N_5755,N_5368);
and UO_1419 (O_1419,N_7402,N_6408);
nor UO_1420 (O_1420,N_5897,N_5490);
xor UO_1421 (O_1421,N_9479,N_9049);
nand UO_1422 (O_1422,N_5682,N_6249);
and UO_1423 (O_1423,N_7045,N_6911);
or UO_1424 (O_1424,N_8310,N_5144);
nor UO_1425 (O_1425,N_9940,N_7430);
or UO_1426 (O_1426,N_7854,N_9308);
or UO_1427 (O_1427,N_8914,N_9744);
or UO_1428 (O_1428,N_8096,N_7634);
or UO_1429 (O_1429,N_7358,N_8466);
or UO_1430 (O_1430,N_8248,N_7384);
or UO_1431 (O_1431,N_7741,N_7731);
or UO_1432 (O_1432,N_7362,N_6536);
nand UO_1433 (O_1433,N_7376,N_5885);
or UO_1434 (O_1434,N_8952,N_9888);
xnor UO_1435 (O_1435,N_8805,N_6036);
or UO_1436 (O_1436,N_9384,N_7909);
or UO_1437 (O_1437,N_5713,N_6754);
xnor UO_1438 (O_1438,N_7160,N_9187);
and UO_1439 (O_1439,N_6240,N_8848);
xnor UO_1440 (O_1440,N_8751,N_8795);
nand UO_1441 (O_1441,N_9486,N_8200);
xnor UO_1442 (O_1442,N_9724,N_8497);
and UO_1443 (O_1443,N_8211,N_8382);
or UO_1444 (O_1444,N_6100,N_9708);
nor UO_1445 (O_1445,N_9592,N_6194);
and UO_1446 (O_1446,N_5569,N_5198);
nand UO_1447 (O_1447,N_8743,N_6410);
and UO_1448 (O_1448,N_8011,N_5061);
xor UO_1449 (O_1449,N_6514,N_8234);
xor UO_1450 (O_1450,N_8485,N_7987);
nor UO_1451 (O_1451,N_6055,N_8553);
and UO_1452 (O_1452,N_7831,N_6372);
nand UO_1453 (O_1453,N_5536,N_7534);
nand UO_1454 (O_1454,N_5234,N_9705);
nor UO_1455 (O_1455,N_5956,N_8436);
nor UO_1456 (O_1456,N_6660,N_5929);
and UO_1457 (O_1457,N_8838,N_5985);
xnor UO_1458 (O_1458,N_7355,N_6439);
xor UO_1459 (O_1459,N_9285,N_9205);
and UO_1460 (O_1460,N_6032,N_7700);
nor UO_1461 (O_1461,N_8772,N_5313);
nor UO_1462 (O_1462,N_5504,N_6667);
nand UO_1463 (O_1463,N_8868,N_8325);
nor UO_1464 (O_1464,N_7423,N_8189);
nand UO_1465 (O_1465,N_8182,N_5521);
and UO_1466 (O_1466,N_6841,N_8263);
nor UO_1467 (O_1467,N_8206,N_6543);
and UO_1468 (O_1468,N_6080,N_9782);
nand UO_1469 (O_1469,N_8171,N_8635);
nand UO_1470 (O_1470,N_9341,N_7074);
and UO_1471 (O_1471,N_9554,N_6092);
nand UO_1472 (O_1472,N_9092,N_7857);
nand UO_1473 (O_1473,N_7759,N_8738);
or UO_1474 (O_1474,N_8177,N_6594);
xnor UO_1475 (O_1475,N_6968,N_9335);
xnor UO_1476 (O_1476,N_5093,N_5172);
xnor UO_1477 (O_1477,N_5332,N_6150);
nor UO_1478 (O_1478,N_7048,N_5795);
and UO_1479 (O_1479,N_9770,N_9639);
xor UO_1480 (O_1480,N_5615,N_8049);
nor UO_1481 (O_1481,N_6276,N_5859);
xor UO_1482 (O_1482,N_6223,N_9106);
and UO_1483 (O_1483,N_7266,N_6492);
xnor UO_1484 (O_1484,N_8814,N_7058);
and UO_1485 (O_1485,N_8042,N_7514);
and UO_1486 (O_1486,N_6115,N_7847);
nor UO_1487 (O_1487,N_5292,N_7396);
or UO_1488 (O_1488,N_6252,N_9047);
or UO_1489 (O_1489,N_6879,N_7906);
xnor UO_1490 (O_1490,N_6380,N_5202);
xnor UO_1491 (O_1491,N_8794,N_7076);
nand UO_1492 (O_1492,N_6942,N_9072);
nand UO_1493 (O_1493,N_6210,N_8394);
xnor UO_1494 (O_1494,N_6788,N_9233);
nand UO_1495 (O_1495,N_6578,N_5484);
xor UO_1496 (O_1496,N_5197,N_5794);
or UO_1497 (O_1497,N_6927,N_5435);
nand UO_1498 (O_1498,N_8284,N_7470);
xnor UO_1499 (O_1499,N_7647,N_8857);
endmodule