module basic_1000_10000_1500_4_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_218,In_740);
nand U1 (N_1,In_594,In_683);
or U2 (N_2,In_892,In_510);
nand U3 (N_3,In_405,In_123);
nor U4 (N_4,In_917,In_628);
xor U5 (N_5,In_209,In_626);
or U6 (N_6,In_623,In_860);
or U7 (N_7,In_494,In_202);
nand U8 (N_8,In_965,In_841);
and U9 (N_9,In_125,In_290);
xor U10 (N_10,In_978,In_586);
and U11 (N_11,In_29,In_276);
or U12 (N_12,In_447,In_338);
nor U13 (N_13,In_739,In_831);
and U14 (N_14,In_307,In_729);
and U15 (N_15,In_62,In_435);
nand U16 (N_16,In_100,In_787);
nand U17 (N_17,In_908,In_489);
nor U18 (N_18,In_808,In_262);
nor U19 (N_19,In_764,In_737);
xnor U20 (N_20,In_482,In_185);
nor U21 (N_21,In_52,In_884);
or U22 (N_22,In_108,In_678);
xnor U23 (N_23,In_958,In_189);
nand U24 (N_24,In_96,In_725);
nand U25 (N_25,In_190,In_599);
and U26 (N_26,In_502,In_56);
and U27 (N_27,In_520,In_508);
nor U28 (N_28,In_661,In_771);
or U29 (N_29,In_631,In_972);
nand U30 (N_30,In_676,In_156);
nor U31 (N_31,In_864,In_608);
nor U32 (N_32,In_797,In_442);
nor U33 (N_33,In_610,In_298);
nand U34 (N_34,In_387,In_408);
nor U35 (N_35,In_653,In_893);
nor U36 (N_36,In_264,In_689);
or U37 (N_37,In_110,In_412);
and U38 (N_38,In_135,In_322);
nor U39 (N_39,In_15,In_675);
xor U40 (N_40,In_0,In_762);
nand U41 (N_41,In_17,In_138);
xor U42 (N_42,In_803,In_187);
and U43 (N_43,In_553,In_27);
and U44 (N_44,In_369,In_778);
nand U45 (N_45,In_57,In_229);
or U46 (N_46,In_756,In_147);
or U47 (N_47,In_145,In_713);
nand U48 (N_48,In_934,In_310);
or U49 (N_49,In_732,In_559);
nor U50 (N_50,In_14,In_227);
xor U51 (N_51,In_681,In_664);
nand U52 (N_52,In_235,In_160);
nor U53 (N_53,In_411,In_195);
or U54 (N_54,In_593,In_548);
nand U55 (N_55,In_943,In_854);
xor U56 (N_56,In_106,In_550);
or U57 (N_57,In_567,In_380);
and U58 (N_58,In_281,In_614);
nor U59 (N_59,In_461,In_761);
and U60 (N_60,In_730,In_24);
nor U61 (N_61,In_840,In_4);
or U62 (N_62,In_319,In_748);
or U63 (N_63,In_643,In_544);
and U64 (N_64,In_485,In_533);
and U65 (N_65,In_248,In_388);
nor U66 (N_66,In_902,In_541);
nand U67 (N_67,In_691,In_634);
nand U68 (N_68,In_871,In_257);
nor U69 (N_69,In_896,In_796);
nand U70 (N_70,In_220,In_144);
nand U71 (N_71,In_970,In_486);
nor U72 (N_72,In_981,In_383);
or U73 (N_73,In_204,In_804);
or U74 (N_74,In_582,In_392);
and U75 (N_75,In_309,In_980);
nand U76 (N_76,In_844,In_308);
or U77 (N_77,In_942,In_382);
xor U78 (N_78,In_351,In_684);
or U79 (N_79,In_720,In_763);
nor U80 (N_80,In_811,In_241);
nor U81 (N_81,In_90,In_199);
or U82 (N_82,In_196,In_346);
and U83 (N_83,In_930,In_872);
xor U84 (N_84,In_999,In_563);
nand U85 (N_85,In_933,In_478);
nand U86 (N_86,In_759,In_617);
nor U87 (N_87,In_237,In_311);
nor U88 (N_88,In_546,In_105);
xor U89 (N_89,In_894,In_613);
xor U90 (N_90,In_172,In_774);
nand U91 (N_91,In_979,In_534);
xor U92 (N_92,In_260,In_747);
and U93 (N_93,In_252,In_306);
nand U94 (N_94,In_506,In_604);
and U95 (N_95,In_517,In_356);
or U96 (N_96,In_873,In_366);
nor U97 (N_97,In_294,In_54);
or U98 (N_98,In_480,In_651);
xor U99 (N_99,In_107,In_846);
or U100 (N_100,In_746,In_420);
nor U101 (N_101,In_279,In_742);
nor U102 (N_102,In_184,In_149);
nand U103 (N_103,In_124,In_75);
and U104 (N_104,In_950,In_445);
nor U105 (N_105,In_368,In_80);
nor U106 (N_106,In_361,In_710);
xor U107 (N_107,In_398,In_292);
or U108 (N_108,In_39,In_216);
or U109 (N_109,In_556,In_900);
nand U110 (N_110,In_84,In_636);
nand U111 (N_111,In_179,In_698);
or U112 (N_112,In_230,In_436);
nand U113 (N_113,In_829,In_606);
xnor U114 (N_114,In_321,In_772);
nand U115 (N_115,In_513,In_878);
nand U116 (N_116,In_73,In_268);
or U117 (N_117,In_512,In_21);
or U118 (N_118,In_335,In_245);
nor U119 (N_119,In_41,In_326);
nor U120 (N_120,In_460,In_537);
and U121 (N_121,In_527,In_519);
or U122 (N_122,In_33,In_285);
nand U123 (N_123,In_704,In_985);
nand U124 (N_124,In_72,In_440);
and U125 (N_125,In_669,In_745);
and U126 (N_126,In_74,In_165);
xnor U127 (N_127,In_801,In_845);
nor U128 (N_128,In_425,In_858);
nand U129 (N_129,In_575,In_466);
and U130 (N_130,In_629,In_496);
and U131 (N_131,In_953,In_814);
or U132 (N_132,In_35,In_407);
and U133 (N_133,In_856,In_528);
or U134 (N_134,In_153,In_826);
nand U135 (N_135,In_112,In_386);
nand U136 (N_136,In_421,In_265);
nor U137 (N_137,In_837,In_602);
nand U138 (N_138,In_552,In_931);
or U139 (N_139,In_869,In_142);
nor U140 (N_140,In_749,In_818);
or U141 (N_141,In_399,In_379);
nand U142 (N_142,In_810,In_148);
or U143 (N_143,In_79,In_484);
or U144 (N_144,In_194,In_956);
or U145 (N_145,In_848,In_775);
or U146 (N_146,In_518,In_3);
and U147 (N_147,In_34,In_441);
or U148 (N_148,In_549,In_201);
nand U149 (N_149,In_340,In_540);
nand U150 (N_150,In_462,In_794);
nand U151 (N_151,In_899,In_444);
or U152 (N_152,In_259,In_654);
nor U153 (N_153,In_768,In_198);
and U154 (N_154,In_781,In_648);
and U155 (N_155,In_897,In_477);
and U156 (N_156,In_94,In_757);
or U157 (N_157,In_36,In_104);
or U158 (N_158,In_585,In_672);
nand U159 (N_159,In_755,In_996);
xor U160 (N_160,In_936,In_402);
xor U161 (N_161,In_906,In_109);
nand U162 (N_162,In_152,In_139);
nor U163 (N_163,In_385,In_941);
xor U164 (N_164,In_70,In_882);
or U165 (N_165,In_963,In_525);
nor U166 (N_166,In_984,In_850);
nor U167 (N_167,In_497,In_171);
nor U168 (N_168,In_339,In_325);
or U169 (N_169,In_577,In_935);
or U170 (N_170,In_700,In_721);
and U171 (N_171,In_918,In_994);
nor U172 (N_172,In_914,In_371);
and U173 (N_173,In_315,In_622);
nor U174 (N_174,In_291,In_955);
and U175 (N_175,In_9,In_469);
nor U176 (N_176,In_688,In_859);
nand U177 (N_177,In_250,In_587);
nor U178 (N_178,In_674,In_31);
xnor U179 (N_179,In_473,In_451);
and U180 (N_180,In_913,In_287);
nand U181 (N_181,In_652,In_716);
and U182 (N_182,In_313,In_116);
nor U183 (N_183,In_303,In_212);
nand U184 (N_184,In_64,In_790);
and U185 (N_185,In_30,In_946);
and U186 (N_186,In_952,In_452);
or U187 (N_187,In_875,In_671);
nand U188 (N_188,In_802,In_373);
or U189 (N_189,In_66,In_481);
and U190 (N_190,In_524,In_855);
or U191 (N_191,In_87,In_211);
or U192 (N_192,In_971,In_573);
or U193 (N_193,In_706,In_58);
nand U194 (N_194,In_719,In_687);
nand U195 (N_195,In_42,In_224);
and U196 (N_196,In_920,In_718);
xor U197 (N_197,In_734,In_616);
or U198 (N_198,In_673,In_103);
xor U199 (N_199,In_532,In_538);
nor U200 (N_200,In_709,In_680);
nand U201 (N_201,In_127,In_113);
nand U202 (N_202,In_120,In_722);
xor U203 (N_203,In_465,In_28);
or U204 (N_204,In_364,In_800);
xnor U205 (N_205,In_503,In_498);
and U206 (N_206,In_428,In_505);
nand U207 (N_207,In_483,In_375);
and U208 (N_208,In_244,In_522);
and U209 (N_209,In_945,In_487);
nand U210 (N_210,In_565,In_403);
or U211 (N_211,In_492,In_342);
or U212 (N_212,In_446,In_887);
and U213 (N_213,In_434,In_865);
nor U214 (N_214,In_923,In_557);
nor U215 (N_215,In_320,In_773);
or U216 (N_216,In_377,In_547);
nor U217 (N_217,In_419,In_170);
nand U218 (N_218,In_238,In_679);
or U219 (N_219,In_246,In_154);
nand U220 (N_220,In_381,In_961);
nor U221 (N_221,In_666,In_530);
or U222 (N_222,In_588,In_59);
nor U223 (N_223,In_347,In_592);
nand U224 (N_224,In_667,In_659);
nand U225 (N_225,In_545,In_48);
or U226 (N_226,In_430,In_944);
xor U227 (N_227,In_889,In_574);
or U228 (N_228,In_901,In_830);
xnor U229 (N_229,In_690,In_886);
or U230 (N_230,In_630,In_870);
and U231 (N_231,In_429,In_214);
or U232 (N_232,In_866,In_861);
and U233 (N_233,In_959,In_891);
nor U234 (N_234,In_514,In_874);
and U235 (N_235,In_345,In_331);
nor U236 (N_236,In_359,In_785);
or U237 (N_237,In_969,In_828);
xnor U238 (N_238,In_293,In_738);
or U239 (N_239,In_81,In_182);
xor U240 (N_240,In_877,In_798);
or U241 (N_241,In_11,In_554);
nand U242 (N_242,In_267,In_376);
and U243 (N_243,In_584,In_349);
or U244 (N_244,In_976,In_910);
nor U245 (N_245,In_205,In_668);
and U246 (N_246,In_711,In_133);
nor U247 (N_247,In_777,In_314);
and U248 (N_248,In_370,In_779);
nor U249 (N_249,In_805,In_611);
nand U250 (N_250,In_752,In_714);
and U251 (N_251,In_449,In_543);
nor U252 (N_252,In_221,In_601);
and U253 (N_253,In_459,In_677);
nor U254 (N_254,In_975,In_397);
nor U255 (N_255,In_605,In_880);
xnor U256 (N_256,In_507,In_280);
xnor U257 (N_257,In_633,In_694);
nor U258 (N_258,In_438,In_23);
nand U259 (N_259,In_389,In_467);
and U260 (N_260,In_159,In_836);
or U261 (N_261,In_355,In_115);
and U262 (N_262,In_932,In_903);
nor U263 (N_263,In_197,In_400);
nand U264 (N_264,In_362,In_409);
and U265 (N_265,In_60,In_7);
and U266 (N_266,In_266,In_639);
and U267 (N_267,In_839,In_566);
nor U268 (N_268,In_61,In_735);
and U269 (N_269,In_164,In_927);
and U270 (N_270,In_558,In_101);
nor U271 (N_271,In_589,In_219);
nand U272 (N_272,In_301,In_578);
nor U273 (N_273,In_997,In_300);
or U274 (N_274,In_753,In_770);
or U275 (N_275,In_278,In_993);
or U276 (N_276,In_863,In_51);
nand U277 (N_277,In_472,In_323);
and U278 (N_278,In_283,In_333);
or U279 (N_279,In_650,In_744);
nand U280 (N_280,In_8,In_157);
nand U281 (N_281,In_213,In_288);
or U282 (N_282,In_568,In_327);
nor U283 (N_283,In_820,In_715);
nor U284 (N_284,In_600,In_210);
or U285 (N_285,In_535,In_134);
nand U286 (N_286,In_925,In_807);
nor U287 (N_287,In_769,In_596);
and U288 (N_288,In_853,In_119);
nand U289 (N_289,In_168,In_200);
nand U290 (N_290,In_663,In_114);
or U291 (N_291,In_962,In_426);
or U292 (N_292,In_20,In_305);
and U293 (N_293,In_849,In_263);
and U294 (N_294,In_418,In_655);
nor U295 (N_295,In_641,In_986);
or U296 (N_296,In_146,In_390);
or U297 (N_297,In_223,In_624);
nor U298 (N_298,In_766,In_329);
nor U299 (N_299,In_560,In_95);
nor U300 (N_300,In_271,In_470);
nand U301 (N_301,In_647,In_504);
nor U302 (N_302,In_111,In_46);
nor U303 (N_303,In_843,In_295);
and U304 (N_304,In_618,In_312);
and U305 (N_305,In_780,In_431);
nor U306 (N_306,In_922,In_130);
nand U307 (N_307,In_26,In_16);
nor U308 (N_308,In_712,In_63);
nor U309 (N_309,In_819,In_708);
nand U310 (N_310,In_247,In_343);
or U311 (N_311,In_93,In_928);
or U312 (N_312,In_609,In_921);
or U313 (N_313,In_423,In_581);
nand U314 (N_314,In_226,In_177);
nor U315 (N_315,In_118,In_905);
and U316 (N_316,In_948,In_348);
and U317 (N_317,In_37,In_49);
and U318 (N_318,In_367,In_523);
or U319 (N_319,In_394,In_458);
nor U320 (N_320,In_916,In_580);
or U321 (N_321,In_324,In_572);
or U322 (N_322,In_55,In_401);
nand U323 (N_323,In_43,In_253);
and U324 (N_324,In_274,In_137);
or U325 (N_325,In_699,In_261);
nand U326 (N_326,In_5,In_888);
and U327 (N_327,In_992,In_131);
nor U328 (N_328,In_957,In_50);
nand U329 (N_329,In_173,In_562);
and U330 (N_330,In_539,In_776);
or U331 (N_331,In_646,In_432);
or U332 (N_332,In_242,In_12);
nor U333 (N_333,In_121,In_98);
nand U334 (N_334,In_175,In_474);
xor U335 (N_335,In_561,In_236);
or U336 (N_336,In_85,In_254);
nand U337 (N_337,In_316,In_181);
or U338 (N_338,In_702,In_475);
nor U339 (N_339,In_670,In_83);
or U340 (N_340,In_22,In_968);
xor U341 (N_341,In_526,In_951);
and U342 (N_342,In_272,In_966);
nor U343 (N_343,In_89,In_332);
or U344 (N_344,In_750,In_792);
or U345 (N_345,In_296,In_217);
nand U346 (N_346,In_838,In_1);
or U347 (N_347,In_847,In_615);
nand U348 (N_348,In_868,In_2);
nand U349 (N_349,In_102,In_82);
and U350 (N_350,In_232,In_571);
and U351 (N_351,In_842,In_126);
and U352 (N_352,In_363,In_717);
or U353 (N_353,In_693,In_354);
and U354 (N_354,In_977,In_192);
or U355 (N_355,In_169,In_649);
or U356 (N_356,In_396,In_117);
or U357 (N_357,In_256,In_337);
and U358 (N_358,In_812,In_76);
and U359 (N_359,In_161,In_988);
or U360 (N_360,In_555,In_695);
or U361 (N_361,In_140,In_612);
nand U362 (N_362,In_823,In_821);
xor U363 (N_363,In_68,In_53);
and U364 (N_364,In_454,In_607);
and U365 (N_365,In_417,In_964);
nor U366 (N_366,In_912,In_591);
or U367 (N_367,In_372,In_299);
or U368 (N_368,In_193,In_10);
or U369 (N_369,In_907,In_783);
nand U370 (N_370,In_542,In_334);
and U371 (N_371,In_178,In_491);
or U372 (N_372,In_645,In_989);
and U373 (N_373,In_833,In_176);
nor U374 (N_374,In_476,In_825);
and U375 (N_375,In_141,In_915);
and U376 (N_376,In_40,In_471);
nand U377 (N_377,In_44,In_625);
and U378 (N_378,In_728,In_45);
or U379 (N_379,In_515,In_191);
and U380 (N_380,In_464,In_665);
nand U381 (N_381,In_97,In_697);
or U382 (N_382,In_286,In_270);
nor U383 (N_383,In_795,In_974);
xnor U384 (N_384,In_686,In_88);
nor U385 (N_385,In_637,In_413);
and U386 (N_386,In_162,In_576);
nor U387 (N_387,In_132,In_495);
or U388 (N_388,In_806,In_437);
or U389 (N_389,In_282,In_188);
nor U390 (N_390,In_439,In_136);
nor U391 (N_391,In_570,In_318);
and U392 (N_392,In_457,In_816);
xor U393 (N_393,In_603,In_788);
and U394 (N_394,In_949,In_167);
and U395 (N_395,In_357,In_304);
nand U396 (N_396,In_391,In_658);
nor U397 (N_397,In_701,In_341);
nand U398 (N_398,In_410,In_32);
or U399 (N_399,In_404,In_597);
nor U400 (N_400,In_758,In_302);
or U401 (N_401,In_143,In_289);
or U402 (N_402,In_983,In_789);
nor U403 (N_403,In_222,In_277);
and U404 (N_404,In_6,In_330);
xnor U405 (N_405,In_71,In_904);
or U406 (N_406,In_509,In_727);
and U407 (N_407,In_743,In_511);
nor U408 (N_408,In_365,In_939);
and U409 (N_409,In_249,In_215);
or U410 (N_410,In_638,In_867);
xnor U411 (N_411,In_521,In_590);
nand U412 (N_412,In_852,In_973);
and U413 (N_413,In_493,In_987);
xor U414 (N_414,In_583,In_621);
and U415 (N_415,In_851,In_809);
and U416 (N_416,In_551,In_751);
nor U417 (N_417,In_427,In_374);
or U418 (N_418,In_862,In_705);
nor U419 (N_419,In_273,In_817);
nor U420 (N_420,In_344,In_662);
nand U421 (N_421,In_536,In_500);
or U422 (N_422,In_832,In_453);
xor U423 (N_423,In_909,In_642);
and U424 (N_424,In_685,In_151);
and U425 (N_425,In_206,In_378);
and U426 (N_426,In_174,In_929);
nand U427 (N_427,In_239,In_898);
nand U428 (N_428,In_724,In_468);
and U429 (N_429,In_657,In_947);
or U430 (N_430,In_251,In_824);
or U431 (N_431,In_919,In_233);
nor U432 (N_432,In_240,In_47);
nor U433 (N_433,In_490,In_879);
nor U434 (N_434,In_982,In_569);
nand U435 (N_435,In_696,In_65);
or U436 (N_436,In_703,In_960);
and U437 (N_437,In_726,In_450);
nor U438 (N_438,In_627,In_424);
nor U439 (N_439,In_353,In_317);
nand U440 (N_440,In_18,In_765);
xnor U441 (N_441,In_736,In_406);
nand U442 (N_442,In_883,In_516);
nand U443 (N_443,In_86,In_660);
nor U444 (N_444,In_122,In_183);
nor U445 (N_445,In_938,In_336);
nand U446 (N_446,In_479,In_741);
nand U447 (N_447,In_350,In_640);
and U448 (N_448,In_998,In_297);
and U449 (N_449,In_754,In_225);
and U450 (N_450,In_876,In_815);
and U451 (N_451,In_924,In_499);
nor U452 (N_452,In_155,In_19);
and U453 (N_453,In_414,In_707);
and U454 (N_454,In_67,In_448);
and U455 (N_455,In_433,In_895);
or U456 (N_456,In_456,In_635);
xor U457 (N_457,In_38,In_619);
nand U458 (N_458,In_443,In_990);
and U459 (N_459,In_284,In_991);
nand U460 (N_460,In_455,In_163);
and U461 (N_461,In_463,In_834);
and U462 (N_462,In_731,In_269);
nor U463 (N_463,In_91,In_358);
and U464 (N_464,In_231,In_128);
xor U465 (N_465,In_733,In_393);
or U466 (N_466,In_793,In_501);
nand U467 (N_467,In_395,In_208);
or U468 (N_468,In_835,In_786);
nand U469 (N_469,In_78,In_275);
and U470 (N_470,In_822,In_595);
and U471 (N_471,In_881,In_416);
and U472 (N_472,In_827,In_258);
and U473 (N_473,In_228,In_644);
or U474 (N_474,In_967,In_692);
or U475 (N_475,In_656,In_415);
nor U476 (N_476,In_911,In_529);
and U477 (N_477,In_180,In_760);
nand U478 (N_478,In_937,In_234);
and U479 (N_479,In_813,In_723);
nor U480 (N_480,In_564,In_77);
and U481 (N_481,In_531,In_579);
nand U482 (N_482,In_158,In_940);
nor U483 (N_483,In_782,In_620);
nand U484 (N_484,In_954,In_890);
or U485 (N_485,In_799,In_186);
nand U486 (N_486,In_99,In_207);
nor U487 (N_487,In_384,In_360);
or U488 (N_488,In_92,In_632);
nor U489 (N_489,In_488,In_995);
and U490 (N_490,In_13,In_69);
or U491 (N_491,In_255,In_857);
or U492 (N_492,In_682,In_129);
or U493 (N_493,In_598,In_784);
and U494 (N_494,In_422,In_203);
nand U495 (N_495,In_328,In_791);
or U496 (N_496,In_352,In_767);
or U497 (N_497,In_243,In_166);
nor U498 (N_498,In_926,In_885);
or U499 (N_499,In_150,In_25);
nand U500 (N_500,In_671,In_634);
nand U501 (N_501,In_140,In_553);
nor U502 (N_502,In_165,In_225);
nor U503 (N_503,In_201,In_974);
nor U504 (N_504,In_654,In_283);
or U505 (N_505,In_177,In_597);
and U506 (N_506,In_365,In_813);
xor U507 (N_507,In_21,In_118);
nand U508 (N_508,In_803,In_662);
xnor U509 (N_509,In_606,In_373);
nor U510 (N_510,In_894,In_985);
or U511 (N_511,In_395,In_69);
xor U512 (N_512,In_99,In_709);
xnor U513 (N_513,In_299,In_876);
or U514 (N_514,In_274,In_573);
or U515 (N_515,In_85,In_822);
nand U516 (N_516,In_515,In_863);
and U517 (N_517,In_865,In_629);
xor U518 (N_518,In_552,In_722);
nand U519 (N_519,In_856,In_625);
and U520 (N_520,In_584,In_119);
nand U521 (N_521,In_661,In_90);
or U522 (N_522,In_482,In_201);
and U523 (N_523,In_948,In_77);
or U524 (N_524,In_843,In_949);
or U525 (N_525,In_612,In_61);
nand U526 (N_526,In_294,In_358);
nand U527 (N_527,In_776,In_364);
nand U528 (N_528,In_627,In_362);
xnor U529 (N_529,In_372,In_688);
or U530 (N_530,In_228,In_943);
nor U531 (N_531,In_77,In_648);
nand U532 (N_532,In_495,In_632);
nor U533 (N_533,In_372,In_504);
nor U534 (N_534,In_244,In_664);
or U535 (N_535,In_302,In_670);
and U536 (N_536,In_54,In_858);
nand U537 (N_537,In_158,In_57);
or U538 (N_538,In_46,In_342);
and U539 (N_539,In_825,In_398);
xor U540 (N_540,In_52,In_747);
nor U541 (N_541,In_740,In_469);
or U542 (N_542,In_769,In_373);
nand U543 (N_543,In_721,In_997);
nor U544 (N_544,In_274,In_752);
xor U545 (N_545,In_274,In_16);
nand U546 (N_546,In_665,In_773);
and U547 (N_547,In_270,In_855);
or U548 (N_548,In_732,In_38);
or U549 (N_549,In_854,In_324);
or U550 (N_550,In_197,In_49);
nand U551 (N_551,In_11,In_223);
nand U552 (N_552,In_858,In_700);
nand U553 (N_553,In_685,In_366);
and U554 (N_554,In_950,In_468);
nand U555 (N_555,In_190,In_85);
nor U556 (N_556,In_448,In_909);
xnor U557 (N_557,In_92,In_754);
xor U558 (N_558,In_13,In_799);
nand U559 (N_559,In_901,In_491);
or U560 (N_560,In_517,In_593);
or U561 (N_561,In_905,In_480);
and U562 (N_562,In_773,In_844);
nor U563 (N_563,In_497,In_365);
nand U564 (N_564,In_151,In_797);
and U565 (N_565,In_460,In_675);
nor U566 (N_566,In_859,In_134);
and U567 (N_567,In_630,In_80);
and U568 (N_568,In_496,In_349);
xnor U569 (N_569,In_119,In_409);
or U570 (N_570,In_838,In_912);
nor U571 (N_571,In_592,In_633);
xor U572 (N_572,In_229,In_557);
or U573 (N_573,In_894,In_704);
nor U574 (N_574,In_110,In_328);
or U575 (N_575,In_965,In_359);
nand U576 (N_576,In_996,In_583);
nand U577 (N_577,In_350,In_289);
nor U578 (N_578,In_46,In_806);
or U579 (N_579,In_198,In_516);
nor U580 (N_580,In_314,In_416);
nor U581 (N_581,In_844,In_353);
nand U582 (N_582,In_961,In_902);
nand U583 (N_583,In_496,In_291);
xnor U584 (N_584,In_249,In_584);
nor U585 (N_585,In_586,In_377);
and U586 (N_586,In_802,In_269);
nand U587 (N_587,In_953,In_535);
nor U588 (N_588,In_481,In_731);
and U589 (N_589,In_921,In_807);
nor U590 (N_590,In_573,In_946);
and U591 (N_591,In_454,In_155);
nor U592 (N_592,In_701,In_933);
nand U593 (N_593,In_464,In_489);
or U594 (N_594,In_253,In_849);
nand U595 (N_595,In_94,In_217);
nor U596 (N_596,In_362,In_58);
nand U597 (N_597,In_943,In_276);
nand U598 (N_598,In_369,In_370);
nor U599 (N_599,In_329,In_377);
nor U600 (N_600,In_345,In_971);
and U601 (N_601,In_650,In_23);
xor U602 (N_602,In_862,In_455);
and U603 (N_603,In_487,In_747);
nor U604 (N_604,In_955,In_301);
and U605 (N_605,In_422,In_711);
nand U606 (N_606,In_726,In_51);
and U607 (N_607,In_172,In_132);
nor U608 (N_608,In_718,In_601);
xnor U609 (N_609,In_15,In_50);
or U610 (N_610,In_399,In_7);
nor U611 (N_611,In_152,In_232);
nand U612 (N_612,In_86,In_419);
and U613 (N_613,In_508,In_527);
or U614 (N_614,In_554,In_958);
or U615 (N_615,In_742,In_97);
xnor U616 (N_616,In_101,In_586);
nor U617 (N_617,In_503,In_260);
nand U618 (N_618,In_9,In_287);
or U619 (N_619,In_204,In_346);
or U620 (N_620,In_760,In_216);
or U621 (N_621,In_67,In_334);
nand U622 (N_622,In_938,In_974);
and U623 (N_623,In_890,In_919);
nand U624 (N_624,In_460,In_669);
nand U625 (N_625,In_100,In_348);
nand U626 (N_626,In_128,In_506);
nand U627 (N_627,In_679,In_374);
nor U628 (N_628,In_82,In_578);
and U629 (N_629,In_683,In_366);
nand U630 (N_630,In_943,In_500);
or U631 (N_631,In_442,In_932);
nor U632 (N_632,In_107,In_268);
nand U633 (N_633,In_13,In_141);
xor U634 (N_634,In_160,In_72);
xor U635 (N_635,In_405,In_9);
or U636 (N_636,In_604,In_738);
nor U637 (N_637,In_399,In_876);
nand U638 (N_638,In_582,In_96);
nand U639 (N_639,In_482,In_58);
nand U640 (N_640,In_170,In_928);
nor U641 (N_641,In_956,In_930);
nor U642 (N_642,In_756,In_802);
nor U643 (N_643,In_350,In_801);
nor U644 (N_644,In_146,In_532);
or U645 (N_645,In_369,In_331);
or U646 (N_646,In_859,In_433);
or U647 (N_647,In_945,In_289);
xor U648 (N_648,In_934,In_29);
or U649 (N_649,In_729,In_211);
xnor U650 (N_650,In_876,In_818);
nand U651 (N_651,In_225,In_213);
or U652 (N_652,In_926,In_67);
and U653 (N_653,In_620,In_45);
or U654 (N_654,In_102,In_229);
and U655 (N_655,In_306,In_955);
or U656 (N_656,In_789,In_623);
nand U657 (N_657,In_785,In_942);
nand U658 (N_658,In_613,In_430);
or U659 (N_659,In_393,In_94);
nor U660 (N_660,In_680,In_397);
or U661 (N_661,In_699,In_827);
nor U662 (N_662,In_209,In_196);
xnor U663 (N_663,In_285,In_869);
nor U664 (N_664,In_809,In_38);
and U665 (N_665,In_184,In_249);
and U666 (N_666,In_334,In_842);
and U667 (N_667,In_17,In_142);
and U668 (N_668,In_63,In_359);
xnor U669 (N_669,In_753,In_561);
nor U670 (N_670,In_914,In_229);
xnor U671 (N_671,In_781,In_877);
nor U672 (N_672,In_545,In_858);
nor U673 (N_673,In_804,In_88);
nand U674 (N_674,In_113,In_682);
nor U675 (N_675,In_311,In_705);
nor U676 (N_676,In_462,In_679);
and U677 (N_677,In_195,In_453);
and U678 (N_678,In_85,In_759);
or U679 (N_679,In_126,In_669);
nand U680 (N_680,In_333,In_818);
and U681 (N_681,In_440,In_488);
nor U682 (N_682,In_489,In_788);
nor U683 (N_683,In_236,In_192);
nand U684 (N_684,In_502,In_798);
and U685 (N_685,In_660,In_135);
xnor U686 (N_686,In_593,In_786);
or U687 (N_687,In_561,In_411);
xor U688 (N_688,In_648,In_148);
nand U689 (N_689,In_753,In_244);
or U690 (N_690,In_155,In_579);
xnor U691 (N_691,In_615,In_420);
and U692 (N_692,In_588,In_586);
nand U693 (N_693,In_653,In_160);
and U694 (N_694,In_726,In_275);
and U695 (N_695,In_662,In_419);
xnor U696 (N_696,In_97,In_208);
or U697 (N_697,In_674,In_709);
or U698 (N_698,In_989,In_339);
and U699 (N_699,In_442,In_354);
nand U700 (N_700,In_615,In_981);
and U701 (N_701,In_50,In_644);
or U702 (N_702,In_717,In_27);
or U703 (N_703,In_640,In_711);
and U704 (N_704,In_990,In_119);
nor U705 (N_705,In_912,In_958);
or U706 (N_706,In_687,In_325);
nand U707 (N_707,In_141,In_235);
nand U708 (N_708,In_318,In_395);
nor U709 (N_709,In_185,In_971);
and U710 (N_710,In_977,In_40);
and U711 (N_711,In_490,In_498);
or U712 (N_712,In_22,In_652);
and U713 (N_713,In_825,In_582);
nor U714 (N_714,In_128,In_690);
and U715 (N_715,In_220,In_920);
xor U716 (N_716,In_281,In_487);
xnor U717 (N_717,In_279,In_249);
or U718 (N_718,In_365,In_36);
or U719 (N_719,In_501,In_126);
xor U720 (N_720,In_834,In_639);
xor U721 (N_721,In_207,In_387);
xor U722 (N_722,In_548,In_756);
or U723 (N_723,In_743,In_868);
or U724 (N_724,In_212,In_891);
nand U725 (N_725,In_183,In_645);
nand U726 (N_726,In_502,In_982);
nand U727 (N_727,In_700,In_90);
nand U728 (N_728,In_834,In_792);
xnor U729 (N_729,In_118,In_749);
nand U730 (N_730,In_348,In_625);
nor U731 (N_731,In_970,In_854);
nand U732 (N_732,In_124,In_617);
or U733 (N_733,In_654,In_443);
or U734 (N_734,In_387,In_594);
nor U735 (N_735,In_524,In_289);
nand U736 (N_736,In_74,In_694);
or U737 (N_737,In_757,In_97);
and U738 (N_738,In_906,In_638);
and U739 (N_739,In_150,In_647);
nor U740 (N_740,In_904,In_310);
or U741 (N_741,In_260,In_782);
nand U742 (N_742,In_351,In_307);
or U743 (N_743,In_247,In_423);
or U744 (N_744,In_985,In_6);
nor U745 (N_745,In_694,In_722);
nand U746 (N_746,In_926,In_187);
or U747 (N_747,In_629,In_842);
or U748 (N_748,In_836,In_766);
nor U749 (N_749,In_183,In_778);
nand U750 (N_750,In_965,In_832);
nand U751 (N_751,In_418,In_866);
nor U752 (N_752,In_580,In_788);
or U753 (N_753,In_334,In_86);
nor U754 (N_754,In_822,In_706);
or U755 (N_755,In_619,In_915);
nor U756 (N_756,In_295,In_453);
and U757 (N_757,In_583,In_850);
nand U758 (N_758,In_55,In_823);
or U759 (N_759,In_310,In_675);
nand U760 (N_760,In_175,In_274);
nand U761 (N_761,In_729,In_966);
nor U762 (N_762,In_909,In_301);
and U763 (N_763,In_752,In_14);
xnor U764 (N_764,In_171,In_8);
nor U765 (N_765,In_735,In_3);
xnor U766 (N_766,In_129,In_412);
and U767 (N_767,In_868,In_394);
and U768 (N_768,In_874,In_498);
and U769 (N_769,In_391,In_289);
xnor U770 (N_770,In_615,In_307);
or U771 (N_771,In_208,In_740);
nor U772 (N_772,In_216,In_236);
and U773 (N_773,In_892,In_952);
and U774 (N_774,In_214,In_544);
nand U775 (N_775,In_835,In_602);
or U776 (N_776,In_670,In_777);
or U777 (N_777,In_654,In_218);
nor U778 (N_778,In_684,In_935);
or U779 (N_779,In_66,In_889);
nor U780 (N_780,In_942,In_27);
and U781 (N_781,In_876,In_853);
or U782 (N_782,In_255,In_726);
nand U783 (N_783,In_426,In_855);
or U784 (N_784,In_505,In_60);
or U785 (N_785,In_124,In_228);
and U786 (N_786,In_958,In_69);
xnor U787 (N_787,In_43,In_352);
nand U788 (N_788,In_106,In_185);
or U789 (N_789,In_962,In_303);
and U790 (N_790,In_424,In_701);
or U791 (N_791,In_641,In_960);
nor U792 (N_792,In_365,In_896);
xnor U793 (N_793,In_347,In_430);
or U794 (N_794,In_165,In_865);
nand U795 (N_795,In_256,In_983);
or U796 (N_796,In_91,In_969);
nand U797 (N_797,In_65,In_351);
nand U798 (N_798,In_889,In_282);
and U799 (N_799,In_549,In_216);
nand U800 (N_800,In_527,In_316);
nand U801 (N_801,In_438,In_917);
or U802 (N_802,In_756,In_95);
and U803 (N_803,In_687,In_172);
nand U804 (N_804,In_837,In_757);
nor U805 (N_805,In_265,In_806);
and U806 (N_806,In_828,In_374);
or U807 (N_807,In_741,In_565);
nand U808 (N_808,In_197,In_282);
and U809 (N_809,In_273,In_13);
nor U810 (N_810,In_968,In_548);
and U811 (N_811,In_399,In_634);
nand U812 (N_812,In_668,In_296);
nand U813 (N_813,In_533,In_974);
xnor U814 (N_814,In_472,In_743);
xor U815 (N_815,In_194,In_630);
or U816 (N_816,In_580,In_443);
and U817 (N_817,In_473,In_642);
or U818 (N_818,In_574,In_430);
or U819 (N_819,In_990,In_23);
nor U820 (N_820,In_887,In_286);
or U821 (N_821,In_167,In_585);
nor U822 (N_822,In_263,In_658);
nand U823 (N_823,In_681,In_929);
nor U824 (N_824,In_206,In_230);
or U825 (N_825,In_793,In_138);
or U826 (N_826,In_493,In_13);
nor U827 (N_827,In_446,In_387);
nor U828 (N_828,In_738,In_411);
and U829 (N_829,In_15,In_491);
nand U830 (N_830,In_37,In_615);
or U831 (N_831,In_672,In_470);
or U832 (N_832,In_488,In_476);
or U833 (N_833,In_707,In_95);
xor U834 (N_834,In_316,In_834);
or U835 (N_835,In_475,In_150);
or U836 (N_836,In_494,In_991);
nor U837 (N_837,In_49,In_559);
nand U838 (N_838,In_860,In_871);
or U839 (N_839,In_100,In_663);
nand U840 (N_840,In_380,In_118);
and U841 (N_841,In_85,In_567);
nor U842 (N_842,In_679,In_288);
nand U843 (N_843,In_564,In_696);
nor U844 (N_844,In_348,In_223);
or U845 (N_845,In_74,In_697);
nor U846 (N_846,In_875,In_674);
nand U847 (N_847,In_210,In_641);
nor U848 (N_848,In_901,In_59);
nand U849 (N_849,In_171,In_242);
or U850 (N_850,In_114,In_205);
xnor U851 (N_851,In_410,In_444);
nor U852 (N_852,In_568,In_577);
nor U853 (N_853,In_959,In_274);
nand U854 (N_854,In_813,In_711);
nor U855 (N_855,In_822,In_666);
or U856 (N_856,In_990,In_926);
nor U857 (N_857,In_974,In_192);
and U858 (N_858,In_585,In_990);
and U859 (N_859,In_232,In_46);
nand U860 (N_860,In_771,In_281);
nor U861 (N_861,In_284,In_87);
or U862 (N_862,In_435,In_711);
nand U863 (N_863,In_353,In_111);
or U864 (N_864,In_984,In_86);
nand U865 (N_865,In_434,In_192);
nor U866 (N_866,In_429,In_567);
nand U867 (N_867,In_6,In_555);
nor U868 (N_868,In_541,In_822);
nor U869 (N_869,In_864,In_508);
or U870 (N_870,In_229,In_496);
nand U871 (N_871,In_873,In_65);
and U872 (N_872,In_695,In_907);
nand U873 (N_873,In_437,In_933);
nor U874 (N_874,In_938,In_29);
or U875 (N_875,In_224,In_221);
or U876 (N_876,In_962,In_422);
or U877 (N_877,In_516,In_50);
or U878 (N_878,In_164,In_263);
nor U879 (N_879,In_96,In_113);
and U880 (N_880,In_763,In_612);
nand U881 (N_881,In_944,In_571);
nor U882 (N_882,In_794,In_638);
nor U883 (N_883,In_706,In_546);
or U884 (N_884,In_762,In_190);
or U885 (N_885,In_423,In_258);
or U886 (N_886,In_704,In_552);
xnor U887 (N_887,In_824,In_764);
nor U888 (N_888,In_135,In_521);
nand U889 (N_889,In_993,In_652);
or U890 (N_890,In_246,In_354);
or U891 (N_891,In_252,In_664);
or U892 (N_892,In_559,In_763);
nor U893 (N_893,In_773,In_207);
nand U894 (N_894,In_187,In_797);
nand U895 (N_895,In_317,In_726);
and U896 (N_896,In_44,In_1);
and U897 (N_897,In_27,In_973);
nor U898 (N_898,In_214,In_265);
or U899 (N_899,In_565,In_242);
nand U900 (N_900,In_895,In_507);
nor U901 (N_901,In_803,In_524);
nor U902 (N_902,In_994,In_702);
or U903 (N_903,In_731,In_664);
nor U904 (N_904,In_672,In_194);
or U905 (N_905,In_675,In_828);
and U906 (N_906,In_379,In_80);
and U907 (N_907,In_154,In_343);
or U908 (N_908,In_236,In_698);
and U909 (N_909,In_744,In_532);
nand U910 (N_910,In_711,In_980);
and U911 (N_911,In_875,In_990);
and U912 (N_912,In_305,In_972);
nand U913 (N_913,In_60,In_429);
and U914 (N_914,In_553,In_814);
and U915 (N_915,In_52,In_161);
nor U916 (N_916,In_671,In_684);
nor U917 (N_917,In_616,In_440);
or U918 (N_918,In_76,In_967);
or U919 (N_919,In_321,In_643);
and U920 (N_920,In_480,In_596);
nor U921 (N_921,In_88,In_504);
xnor U922 (N_922,In_214,In_202);
and U923 (N_923,In_474,In_670);
nand U924 (N_924,In_206,In_521);
and U925 (N_925,In_500,In_830);
nand U926 (N_926,In_719,In_397);
nor U927 (N_927,In_602,In_641);
xor U928 (N_928,In_338,In_269);
and U929 (N_929,In_886,In_697);
and U930 (N_930,In_120,In_771);
nor U931 (N_931,In_188,In_555);
and U932 (N_932,In_710,In_715);
nor U933 (N_933,In_755,In_476);
and U934 (N_934,In_258,In_153);
and U935 (N_935,In_927,In_795);
or U936 (N_936,In_35,In_367);
nor U937 (N_937,In_6,In_251);
and U938 (N_938,In_732,In_673);
or U939 (N_939,In_706,In_8);
nand U940 (N_940,In_208,In_233);
and U941 (N_941,In_553,In_244);
or U942 (N_942,In_307,In_919);
xor U943 (N_943,In_185,In_386);
nor U944 (N_944,In_693,In_83);
xnor U945 (N_945,In_911,In_242);
nand U946 (N_946,In_3,In_540);
nor U947 (N_947,In_574,In_820);
nand U948 (N_948,In_860,In_740);
nor U949 (N_949,In_103,In_938);
or U950 (N_950,In_282,In_384);
and U951 (N_951,In_442,In_6);
and U952 (N_952,In_954,In_377);
and U953 (N_953,In_732,In_237);
nand U954 (N_954,In_14,In_633);
or U955 (N_955,In_255,In_392);
xnor U956 (N_956,In_198,In_164);
and U957 (N_957,In_590,In_943);
nand U958 (N_958,In_775,In_843);
xor U959 (N_959,In_974,In_591);
nand U960 (N_960,In_422,In_767);
nand U961 (N_961,In_524,In_211);
and U962 (N_962,In_730,In_280);
and U963 (N_963,In_471,In_262);
or U964 (N_964,In_49,In_269);
or U965 (N_965,In_373,In_547);
and U966 (N_966,In_858,In_855);
nor U967 (N_967,In_870,In_611);
or U968 (N_968,In_583,In_339);
and U969 (N_969,In_327,In_875);
xor U970 (N_970,In_769,In_232);
or U971 (N_971,In_609,In_173);
and U972 (N_972,In_455,In_972);
nand U973 (N_973,In_225,In_345);
nand U974 (N_974,In_109,In_44);
nor U975 (N_975,In_169,In_415);
and U976 (N_976,In_376,In_369);
or U977 (N_977,In_654,In_393);
and U978 (N_978,In_201,In_845);
xor U979 (N_979,In_544,In_415);
nor U980 (N_980,In_90,In_223);
nand U981 (N_981,In_734,In_977);
nand U982 (N_982,In_213,In_986);
nand U983 (N_983,In_768,In_218);
nand U984 (N_984,In_738,In_897);
or U985 (N_985,In_285,In_817);
and U986 (N_986,In_648,In_294);
nand U987 (N_987,In_328,In_402);
nand U988 (N_988,In_394,In_860);
nor U989 (N_989,In_688,In_168);
nor U990 (N_990,In_715,In_66);
nand U991 (N_991,In_158,In_425);
or U992 (N_992,In_13,In_647);
nand U993 (N_993,In_467,In_119);
nand U994 (N_994,In_130,In_631);
and U995 (N_995,In_259,In_52);
or U996 (N_996,In_782,In_844);
nor U997 (N_997,In_527,In_878);
nor U998 (N_998,In_67,In_818);
or U999 (N_999,In_552,In_385);
nand U1000 (N_1000,In_321,In_396);
or U1001 (N_1001,In_251,In_358);
nand U1002 (N_1002,In_158,In_120);
nor U1003 (N_1003,In_462,In_579);
and U1004 (N_1004,In_408,In_214);
nor U1005 (N_1005,In_847,In_876);
nor U1006 (N_1006,In_926,In_329);
and U1007 (N_1007,In_535,In_261);
or U1008 (N_1008,In_732,In_943);
nor U1009 (N_1009,In_411,In_183);
and U1010 (N_1010,In_111,In_423);
nor U1011 (N_1011,In_190,In_108);
or U1012 (N_1012,In_677,In_346);
nand U1013 (N_1013,In_707,In_808);
nor U1014 (N_1014,In_798,In_169);
nand U1015 (N_1015,In_777,In_70);
xnor U1016 (N_1016,In_618,In_636);
nand U1017 (N_1017,In_817,In_499);
and U1018 (N_1018,In_77,In_525);
or U1019 (N_1019,In_666,In_834);
or U1020 (N_1020,In_155,In_53);
nand U1021 (N_1021,In_272,In_932);
or U1022 (N_1022,In_430,In_768);
nand U1023 (N_1023,In_927,In_647);
nor U1024 (N_1024,In_792,In_681);
nand U1025 (N_1025,In_447,In_701);
or U1026 (N_1026,In_922,In_983);
or U1027 (N_1027,In_371,In_421);
nor U1028 (N_1028,In_222,In_302);
or U1029 (N_1029,In_497,In_742);
or U1030 (N_1030,In_565,In_971);
or U1031 (N_1031,In_726,In_250);
nand U1032 (N_1032,In_292,In_62);
nand U1033 (N_1033,In_358,In_142);
and U1034 (N_1034,In_391,In_877);
and U1035 (N_1035,In_846,In_303);
and U1036 (N_1036,In_185,In_180);
and U1037 (N_1037,In_403,In_136);
xor U1038 (N_1038,In_902,In_890);
nand U1039 (N_1039,In_679,In_421);
xor U1040 (N_1040,In_439,In_90);
nor U1041 (N_1041,In_403,In_336);
nor U1042 (N_1042,In_155,In_866);
nor U1043 (N_1043,In_364,In_740);
nor U1044 (N_1044,In_675,In_774);
or U1045 (N_1045,In_631,In_63);
nor U1046 (N_1046,In_504,In_153);
nand U1047 (N_1047,In_73,In_174);
and U1048 (N_1048,In_979,In_414);
nand U1049 (N_1049,In_696,In_627);
nand U1050 (N_1050,In_584,In_887);
or U1051 (N_1051,In_607,In_582);
and U1052 (N_1052,In_925,In_548);
nor U1053 (N_1053,In_157,In_902);
or U1054 (N_1054,In_762,In_545);
and U1055 (N_1055,In_552,In_743);
nand U1056 (N_1056,In_749,In_3);
and U1057 (N_1057,In_695,In_964);
or U1058 (N_1058,In_909,In_110);
nand U1059 (N_1059,In_558,In_611);
nor U1060 (N_1060,In_768,In_693);
or U1061 (N_1061,In_475,In_448);
or U1062 (N_1062,In_948,In_786);
xor U1063 (N_1063,In_356,In_728);
or U1064 (N_1064,In_993,In_558);
xor U1065 (N_1065,In_213,In_783);
xor U1066 (N_1066,In_327,In_815);
nor U1067 (N_1067,In_363,In_486);
nor U1068 (N_1068,In_393,In_44);
or U1069 (N_1069,In_480,In_181);
nand U1070 (N_1070,In_989,In_108);
or U1071 (N_1071,In_747,In_607);
nor U1072 (N_1072,In_471,In_599);
nor U1073 (N_1073,In_265,In_316);
or U1074 (N_1074,In_624,In_106);
nand U1075 (N_1075,In_472,In_754);
or U1076 (N_1076,In_463,In_395);
and U1077 (N_1077,In_25,In_268);
nand U1078 (N_1078,In_106,In_693);
nor U1079 (N_1079,In_588,In_503);
and U1080 (N_1080,In_100,In_874);
and U1081 (N_1081,In_393,In_93);
nor U1082 (N_1082,In_439,In_584);
nor U1083 (N_1083,In_728,In_460);
nor U1084 (N_1084,In_474,In_232);
nand U1085 (N_1085,In_539,In_102);
and U1086 (N_1086,In_812,In_740);
nor U1087 (N_1087,In_972,In_196);
or U1088 (N_1088,In_593,In_465);
nor U1089 (N_1089,In_810,In_251);
or U1090 (N_1090,In_363,In_916);
and U1091 (N_1091,In_179,In_865);
nand U1092 (N_1092,In_399,In_241);
nand U1093 (N_1093,In_578,In_850);
and U1094 (N_1094,In_266,In_645);
or U1095 (N_1095,In_761,In_689);
xnor U1096 (N_1096,In_465,In_78);
or U1097 (N_1097,In_61,In_851);
and U1098 (N_1098,In_724,In_373);
or U1099 (N_1099,In_606,In_837);
and U1100 (N_1100,In_830,In_891);
nor U1101 (N_1101,In_531,In_516);
and U1102 (N_1102,In_390,In_863);
or U1103 (N_1103,In_177,In_423);
or U1104 (N_1104,In_860,In_362);
xor U1105 (N_1105,In_42,In_242);
nand U1106 (N_1106,In_154,In_210);
nor U1107 (N_1107,In_266,In_936);
nand U1108 (N_1108,In_826,In_189);
nor U1109 (N_1109,In_161,In_725);
xnor U1110 (N_1110,In_127,In_949);
nor U1111 (N_1111,In_642,In_159);
xnor U1112 (N_1112,In_635,In_522);
and U1113 (N_1113,In_554,In_336);
or U1114 (N_1114,In_955,In_361);
and U1115 (N_1115,In_314,In_208);
nand U1116 (N_1116,In_445,In_69);
nand U1117 (N_1117,In_706,In_376);
nand U1118 (N_1118,In_577,In_576);
and U1119 (N_1119,In_57,In_912);
nor U1120 (N_1120,In_155,In_175);
nor U1121 (N_1121,In_52,In_408);
nand U1122 (N_1122,In_716,In_730);
or U1123 (N_1123,In_995,In_48);
and U1124 (N_1124,In_254,In_265);
nor U1125 (N_1125,In_160,In_680);
nand U1126 (N_1126,In_396,In_602);
nand U1127 (N_1127,In_586,In_173);
or U1128 (N_1128,In_108,In_559);
nand U1129 (N_1129,In_492,In_361);
xor U1130 (N_1130,In_942,In_747);
and U1131 (N_1131,In_189,In_461);
nor U1132 (N_1132,In_0,In_659);
or U1133 (N_1133,In_603,In_80);
xor U1134 (N_1134,In_814,In_558);
and U1135 (N_1135,In_777,In_894);
nand U1136 (N_1136,In_13,In_246);
nand U1137 (N_1137,In_592,In_840);
and U1138 (N_1138,In_958,In_718);
or U1139 (N_1139,In_946,In_228);
or U1140 (N_1140,In_133,In_390);
or U1141 (N_1141,In_307,In_912);
or U1142 (N_1142,In_566,In_510);
or U1143 (N_1143,In_739,In_650);
or U1144 (N_1144,In_594,In_655);
and U1145 (N_1145,In_721,In_481);
nor U1146 (N_1146,In_952,In_118);
and U1147 (N_1147,In_619,In_976);
or U1148 (N_1148,In_670,In_698);
nor U1149 (N_1149,In_625,In_959);
or U1150 (N_1150,In_453,In_603);
nand U1151 (N_1151,In_619,In_513);
or U1152 (N_1152,In_393,In_342);
nand U1153 (N_1153,In_750,In_559);
and U1154 (N_1154,In_394,In_688);
nand U1155 (N_1155,In_933,In_328);
xnor U1156 (N_1156,In_962,In_388);
nand U1157 (N_1157,In_610,In_839);
and U1158 (N_1158,In_381,In_152);
xor U1159 (N_1159,In_638,In_992);
and U1160 (N_1160,In_382,In_879);
nor U1161 (N_1161,In_739,In_468);
or U1162 (N_1162,In_500,In_142);
nor U1163 (N_1163,In_626,In_651);
nand U1164 (N_1164,In_999,In_572);
and U1165 (N_1165,In_253,In_743);
nand U1166 (N_1166,In_609,In_713);
nor U1167 (N_1167,In_717,In_854);
and U1168 (N_1168,In_193,In_664);
nor U1169 (N_1169,In_141,In_602);
nand U1170 (N_1170,In_588,In_435);
nor U1171 (N_1171,In_484,In_195);
or U1172 (N_1172,In_874,In_722);
nand U1173 (N_1173,In_979,In_809);
nand U1174 (N_1174,In_159,In_744);
or U1175 (N_1175,In_542,In_778);
nand U1176 (N_1176,In_452,In_862);
nor U1177 (N_1177,In_454,In_209);
and U1178 (N_1178,In_407,In_478);
and U1179 (N_1179,In_693,In_650);
or U1180 (N_1180,In_168,In_488);
xnor U1181 (N_1181,In_608,In_386);
nand U1182 (N_1182,In_615,In_146);
or U1183 (N_1183,In_129,In_209);
and U1184 (N_1184,In_674,In_195);
or U1185 (N_1185,In_961,In_781);
nand U1186 (N_1186,In_705,In_377);
nand U1187 (N_1187,In_465,In_53);
and U1188 (N_1188,In_930,In_62);
and U1189 (N_1189,In_891,In_25);
xor U1190 (N_1190,In_813,In_925);
or U1191 (N_1191,In_913,In_543);
nand U1192 (N_1192,In_838,In_368);
and U1193 (N_1193,In_832,In_985);
xor U1194 (N_1194,In_778,In_860);
xor U1195 (N_1195,In_173,In_83);
or U1196 (N_1196,In_934,In_159);
and U1197 (N_1197,In_736,In_593);
or U1198 (N_1198,In_626,In_406);
or U1199 (N_1199,In_740,In_61);
nand U1200 (N_1200,In_680,In_919);
and U1201 (N_1201,In_258,In_952);
nand U1202 (N_1202,In_664,In_457);
or U1203 (N_1203,In_670,In_561);
nand U1204 (N_1204,In_735,In_417);
nor U1205 (N_1205,In_458,In_659);
and U1206 (N_1206,In_500,In_600);
xnor U1207 (N_1207,In_958,In_792);
nor U1208 (N_1208,In_677,In_535);
nand U1209 (N_1209,In_152,In_965);
or U1210 (N_1210,In_478,In_799);
nor U1211 (N_1211,In_371,In_182);
nand U1212 (N_1212,In_546,In_78);
nand U1213 (N_1213,In_898,In_205);
or U1214 (N_1214,In_870,In_4);
nand U1215 (N_1215,In_758,In_110);
nor U1216 (N_1216,In_496,In_798);
xor U1217 (N_1217,In_848,In_671);
nand U1218 (N_1218,In_41,In_68);
and U1219 (N_1219,In_774,In_618);
nor U1220 (N_1220,In_653,In_738);
or U1221 (N_1221,In_377,In_730);
nor U1222 (N_1222,In_559,In_337);
or U1223 (N_1223,In_265,In_150);
and U1224 (N_1224,In_88,In_323);
and U1225 (N_1225,In_304,In_514);
nand U1226 (N_1226,In_547,In_223);
and U1227 (N_1227,In_920,In_112);
nand U1228 (N_1228,In_827,In_520);
and U1229 (N_1229,In_395,In_717);
xnor U1230 (N_1230,In_932,In_803);
or U1231 (N_1231,In_687,In_639);
nor U1232 (N_1232,In_733,In_363);
or U1233 (N_1233,In_993,In_145);
nand U1234 (N_1234,In_21,In_17);
nand U1235 (N_1235,In_272,In_233);
nor U1236 (N_1236,In_783,In_836);
and U1237 (N_1237,In_33,In_388);
or U1238 (N_1238,In_498,In_960);
xor U1239 (N_1239,In_649,In_547);
and U1240 (N_1240,In_206,In_83);
nor U1241 (N_1241,In_974,In_682);
nor U1242 (N_1242,In_107,In_49);
nor U1243 (N_1243,In_994,In_347);
and U1244 (N_1244,In_285,In_745);
or U1245 (N_1245,In_922,In_790);
xor U1246 (N_1246,In_767,In_909);
nand U1247 (N_1247,In_13,In_168);
and U1248 (N_1248,In_815,In_959);
or U1249 (N_1249,In_24,In_761);
nand U1250 (N_1250,In_195,In_668);
and U1251 (N_1251,In_575,In_716);
or U1252 (N_1252,In_548,In_28);
or U1253 (N_1253,In_323,In_424);
or U1254 (N_1254,In_243,In_194);
nor U1255 (N_1255,In_159,In_752);
nand U1256 (N_1256,In_136,In_150);
nand U1257 (N_1257,In_532,In_936);
xor U1258 (N_1258,In_906,In_57);
and U1259 (N_1259,In_325,In_978);
and U1260 (N_1260,In_406,In_685);
nand U1261 (N_1261,In_29,In_774);
or U1262 (N_1262,In_324,In_111);
nor U1263 (N_1263,In_732,In_426);
and U1264 (N_1264,In_399,In_695);
or U1265 (N_1265,In_47,In_840);
nand U1266 (N_1266,In_915,In_307);
nand U1267 (N_1267,In_838,In_83);
nand U1268 (N_1268,In_660,In_419);
nor U1269 (N_1269,In_833,In_942);
xnor U1270 (N_1270,In_145,In_849);
or U1271 (N_1271,In_593,In_925);
and U1272 (N_1272,In_796,In_809);
and U1273 (N_1273,In_102,In_848);
nor U1274 (N_1274,In_617,In_892);
and U1275 (N_1275,In_467,In_572);
nor U1276 (N_1276,In_447,In_118);
or U1277 (N_1277,In_877,In_273);
and U1278 (N_1278,In_468,In_88);
nand U1279 (N_1279,In_425,In_207);
or U1280 (N_1280,In_517,In_850);
or U1281 (N_1281,In_580,In_466);
xor U1282 (N_1282,In_504,In_932);
nor U1283 (N_1283,In_571,In_348);
nor U1284 (N_1284,In_376,In_811);
nor U1285 (N_1285,In_750,In_489);
or U1286 (N_1286,In_755,In_386);
nand U1287 (N_1287,In_752,In_185);
and U1288 (N_1288,In_892,In_41);
nand U1289 (N_1289,In_937,In_945);
and U1290 (N_1290,In_83,In_408);
or U1291 (N_1291,In_488,In_53);
and U1292 (N_1292,In_244,In_432);
xnor U1293 (N_1293,In_786,In_880);
nand U1294 (N_1294,In_226,In_436);
nand U1295 (N_1295,In_125,In_46);
and U1296 (N_1296,In_151,In_849);
or U1297 (N_1297,In_294,In_186);
or U1298 (N_1298,In_972,In_582);
nand U1299 (N_1299,In_133,In_449);
and U1300 (N_1300,In_371,In_39);
nand U1301 (N_1301,In_899,In_258);
and U1302 (N_1302,In_741,In_53);
or U1303 (N_1303,In_748,In_678);
or U1304 (N_1304,In_460,In_76);
and U1305 (N_1305,In_63,In_494);
nand U1306 (N_1306,In_309,In_922);
nand U1307 (N_1307,In_92,In_122);
and U1308 (N_1308,In_863,In_567);
nor U1309 (N_1309,In_403,In_36);
nor U1310 (N_1310,In_222,In_269);
nand U1311 (N_1311,In_57,In_740);
or U1312 (N_1312,In_74,In_833);
or U1313 (N_1313,In_274,In_358);
or U1314 (N_1314,In_716,In_371);
and U1315 (N_1315,In_35,In_980);
nor U1316 (N_1316,In_549,In_306);
nand U1317 (N_1317,In_50,In_149);
and U1318 (N_1318,In_416,In_955);
nand U1319 (N_1319,In_832,In_309);
and U1320 (N_1320,In_10,In_938);
and U1321 (N_1321,In_916,In_146);
nand U1322 (N_1322,In_732,In_211);
and U1323 (N_1323,In_494,In_861);
or U1324 (N_1324,In_61,In_461);
nor U1325 (N_1325,In_303,In_464);
and U1326 (N_1326,In_561,In_873);
and U1327 (N_1327,In_334,In_589);
nor U1328 (N_1328,In_995,In_976);
or U1329 (N_1329,In_701,In_541);
and U1330 (N_1330,In_754,In_735);
or U1331 (N_1331,In_597,In_600);
nor U1332 (N_1332,In_241,In_583);
or U1333 (N_1333,In_800,In_515);
xor U1334 (N_1334,In_121,In_437);
and U1335 (N_1335,In_48,In_901);
nand U1336 (N_1336,In_5,In_324);
nor U1337 (N_1337,In_243,In_59);
nor U1338 (N_1338,In_345,In_594);
and U1339 (N_1339,In_954,In_657);
and U1340 (N_1340,In_455,In_116);
nand U1341 (N_1341,In_840,In_769);
xor U1342 (N_1342,In_786,In_633);
nand U1343 (N_1343,In_918,In_38);
or U1344 (N_1344,In_225,In_921);
or U1345 (N_1345,In_353,In_222);
and U1346 (N_1346,In_125,In_586);
nand U1347 (N_1347,In_498,In_44);
or U1348 (N_1348,In_261,In_640);
and U1349 (N_1349,In_148,In_41);
and U1350 (N_1350,In_440,In_847);
or U1351 (N_1351,In_311,In_96);
nand U1352 (N_1352,In_229,In_780);
xor U1353 (N_1353,In_902,In_468);
and U1354 (N_1354,In_165,In_651);
and U1355 (N_1355,In_116,In_325);
or U1356 (N_1356,In_247,In_912);
and U1357 (N_1357,In_637,In_831);
and U1358 (N_1358,In_36,In_258);
or U1359 (N_1359,In_580,In_708);
nand U1360 (N_1360,In_533,In_688);
and U1361 (N_1361,In_785,In_383);
nand U1362 (N_1362,In_767,In_54);
nor U1363 (N_1363,In_474,In_235);
nor U1364 (N_1364,In_604,In_97);
nor U1365 (N_1365,In_279,In_114);
nand U1366 (N_1366,In_498,In_643);
nand U1367 (N_1367,In_298,In_897);
and U1368 (N_1368,In_260,In_501);
or U1369 (N_1369,In_654,In_547);
or U1370 (N_1370,In_573,In_301);
xor U1371 (N_1371,In_139,In_839);
and U1372 (N_1372,In_824,In_269);
nand U1373 (N_1373,In_542,In_394);
and U1374 (N_1374,In_68,In_58);
or U1375 (N_1375,In_261,In_402);
or U1376 (N_1376,In_29,In_84);
nor U1377 (N_1377,In_667,In_699);
and U1378 (N_1378,In_567,In_278);
and U1379 (N_1379,In_415,In_871);
and U1380 (N_1380,In_878,In_154);
xnor U1381 (N_1381,In_963,In_957);
or U1382 (N_1382,In_859,In_464);
or U1383 (N_1383,In_732,In_86);
nand U1384 (N_1384,In_977,In_706);
nor U1385 (N_1385,In_266,In_239);
and U1386 (N_1386,In_984,In_879);
and U1387 (N_1387,In_609,In_281);
nor U1388 (N_1388,In_419,In_28);
and U1389 (N_1389,In_809,In_687);
nand U1390 (N_1390,In_291,In_559);
or U1391 (N_1391,In_350,In_943);
or U1392 (N_1392,In_256,In_541);
nor U1393 (N_1393,In_784,In_250);
and U1394 (N_1394,In_722,In_851);
nand U1395 (N_1395,In_209,In_550);
and U1396 (N_1396,In_111,In_750);
nor U1397 (N_1397,In_214,In_58);
nand U1398 (N_1398,In_121,In_391);
and U1399 (N_1399,In_234,In_693);
nand U1400 (N_1400,In_634,In_814);
or U1401 (N_1401,In_124,In_357);
nor U1402 (N_1402,In_805,In_235);
nand U1403 (N_1403,In_206,In_841);
and U1404 (N_1404,In_177,In_775);
or U1405 (N_1405,In_561,In_420);
nor U1406 (N_1406,In_628,In_391);
or U1407 (N_1407,In_202,In_654);
nand U1408 (N_1408,In_131,In_985);
and U1409 (N_1409,In_217,In_120);
nor U1410 (N_1410,In_468,In_728);
or U1411 (N_1411,In_326,In_160);
or U1412 (N_1412,In_584,In_989);
and U1413 (N_1413,In_395,In_182);
or U1414 (N_1414,In_929,In_764);
or U1415 (N_1415,In_825,In_737);
nor U1416 (N_1416,In_830,In_707);
nand U1417 (N_1417,In_557,In_285);
or U1418 (N_1418,In_497,In_739);
nor U1419 (N_1419,In_370,In_612);
or U1420 (N_1420,In_945,In_542);
nor U1421 (N_1421,In_127,In_856);
nand U1422 (N_1422,In_735,In_475);
nor U1423 (N_1423,In_173,In_554);
and U1424 (N_1424,In_878,In_157);
or U1425 (N_1425,In_990,In_537);
nand U1426 (N_1426,In_743,In_783);
nor U1427 (N_1427,In_722,In_297);
nand U1428 (N_1428,In_239,In_585);
or U1429 (N_1429,In_192,In_584);
nor U1430 (N_1430,In_821,In_621);
nand U1431 (N_1431,In_132,In_679);
or U1432 (N_1432,In_29,In_114);
nor U1433 (N_1433,In_616,In_227);
nand U1434 (N_1434,In_771,In_908);
nor U1435 (N_1435,In_867,In_336);
nand U1436 (N_1436,In_483,In_571);
or U1437 (N_1437,In_593,In_221);
or U1438 (N_1438,In_138,In_701);
and U1439 (N_1439,In_634,In_657);
or U1440 (N_1440,In_574,In_687);
nor U1441 (N_1441,In_55,In_607);
or U1442 (N_1442,In_386,In_397);
and U1443 (N_1443,In_765,In_586);
nor U1444 (N_1444,In_269,In_948);
and U1445 (N_1445,In_513,In_584);
nor U1446 (N_1446,In_714,In_401);
or U1447 (N_1447,In_545,In_139);
and U1448 (N_1448,In_361,In_98);
nand U1449 (N_1449,In_349,In_688);
nor U1450 (N_1450,In_763,In_125);
and U1451 (N_1451,In_587,In_929);
or U1452 (N_1452,In_933,In_487);
and U1453 (N_1453,In_371,In_912);
nand U1454 (N_1454,In_206,In_987);
or U1455 (N_1455,In_570,In_464);
nand U1456 (N_1456,In_916,In_206);
or U1457 (N_1457,In_484,In_945);
nand U1458 (N_1458,In_45,In_329);
and U1459 (N_1459,In_652,In_994);
nor U1460 (N_1460,In_198,In_423);
nor U1461 (N_1461,In_145,In_532);
or U1462 (N_1462,In_92,In_95);
nor U1463 (N_1463,In_952,In_692);
nand U1464 (N_1464,In_750,In_479);
and U1465 (N_1465,In_380,In_903);
and U1466 (N_1466,In_91,In_528);
or U1467 (N_1467,In_305,In_686);
nor U1468 (N_1468,In_412,In_490);
and U1469 (N_1469,In_340,In_997);
nand U1470 (N_1470,In_606,In_105);
or U1471 (N_1471,In_812,In_115);
xor U1472 (N_1472,In_402,In_814);
and U1473 (N_1473,In_923,In_744);
and U1474 (N_1474,In_375,In_463);
nand U1475 (N_1475,In_119,In_477);
or U1476 (N_1476,In_514,In_307);
nor U1477 (N_1477,In_394,In_959);
and U1478 (N_1478,In_970,In_307);
nor U1479 (N_1479,In_130,In_133);
and U1480 (N_1480,In_58,In_522);
xor U1481 (N_1481,In_779,In_139);
xor U1482 (N_1482,In_75,In_482);
nor U1483 (N_1483,In_118,In_682);
nand U1484 (N_1484,In_871,In_717);
or U1485 (N_1485,In_703,In_418);
xor U1486 (N_1486,In_830,In_229);
nor U1487 (N_1487,In_898,In_767);
nor U1488 (N_1488,In_591,In_780);
nand U1489 (N_1489,In_784,In_191);
nand U1490 (N_1490,In_30,In_362);
nor U1491 (N_1491,In_882,In_147);
nor U1492 (N_1492,In_282,In_489);
xor U1493 (N_1493,In_459,In_950);
nor U1494 (N_1494,In_201,In_739);
or U1495 (N_1495,In_993,In_23);
and U1496 (N_1496,In_145,In_527);
nand U1497 (N_1497,In_800,In_605);
xor U1498 (N_1498,In_565,In_137);
nor U1499 (N_1499,In_380,In_659);
and U1500 (N_1500,In_984,In_215);
xnor U1501 (N_1501,In_618,In_339);
nor U1502 (N_1502,In_973,In_353);
nand U1503 (N_1503,In_849,In_767);
nor U1504 (N_1504,In_688,In_670);
or U1505 (N_1505,In_969,In_917);
nor U1506 (N_1506,In_573,In_837);
nor U1507 (N_1507,In_328,In_183);
xnor U1508 (N_1508,In_574,In_892);
and U1509 (N_1509,In_942,In_409);
and U1510 (N_1510,In_381,In_431);
nand U1511 (N_1511,In_554,In_957);
and U1512 (N_1512,In_521,In_425);
nand U1513 (N_1513,In_484,In_138);
and U1514 (N_1514,In_780,In_712);
nand U1515 (N_1515,In_779,In_481);
nor U1516 (N_1516,In_313,In_182);
nand U1517 (N_1517,In_617,In_502);
and U1518 (N_1518,In_638,In_642);
and U1519 (N_1519,In_412,In_810);
nor U1520 (N_1520,In_868,In_609);
nand U1521 (N_1521,In_480,In_512);
xnor U1522 (N_1522,In_578,In_415);
and U1523 (N_1523,In_537,In_703);
or U1524 (N_1524,In_872,In_337);
nand U1525 (N_1525,In_40,In_441);
and U1526 (N_1526,In_516,In_949);
and U1527 (N_1527,In_920,In_877);
or U1528 (N_1528,In_556,In_8);
xor U1529 (N_1529,In_167,In_953);
nand U1530 (N_1530,In_562,In_34);
xor U1531 (N_1531,In_46,In_963);
xnor U1532 (N_1532,In_617,In_12);
xor U1533 (N_1533,In_767,In_448);
and U1534 (N_1534,In_701,In_218);
nor U1535 (N_1535,In_260,In_103);
nor U1536 (N_1536,In_938,In_232);
nand U1537 (N_1537,In_1,In_319);
nor U1538 (N_1538,In_796,In_351);
nand U1539 (N_1539,In_226,In_86);
or U1540 (N_1540,In_565,In_877);
xnor U1541 (N_1541,In_69,In_107);
nand U1542 (N_1542,In_389,In_565);
and U1543 (N_1543,In_569,In_917);
nand U1544 (N_1544,In_361,In_686);
nand U1545 (N_1545,In_320,In_84);
nand U1546 (N_1546,In_878,In_833);
nand U1547 (N_1547,In_191,In_467);
or U1548 (N_1548,In_37,In_566);
nand U1549 (N_1549,In_465,In_556);
xnor U1550 (N_1550,In_274,In_14);
and U1551 (N_1551,In_240,In_620);
nand U1552 (N_1552,In_914,In_31);
and U1553 (N_1553,In_675,In_365);
or U1554 (N_1554,In_794,In_64);
or U1555 (N_1555,In_860,In_301);
and U1556 (N_1556,In_227,In_490);
or U1557 (N_1557,In_165,In_132);
nor U1558 (N_1558,In_556,In_947);
and U1559 (N_1559,In_72,In_983);
or U1560 (N_1560,In_638,In_518);
and U1561 (N_1561,In_523,In_141);
xnor U1562 (N_1562,In_610,In_801);
xnor U1563 (N_1563,In_981,In_448);
or U1564 (N_1564,In_562,In_784);
and U1565 (N_1565,In_470,In_562);
and U1566 (N_1566,In_908,In_129);
nand U1567 (N_1567,In_179,In_615);
nand U1568 (N_1568,In_836,In_442);
xnor U1569 (N_1569,In_406,In_827);
and U1570 (N_1570,In_743,In_904);
and U1571 (N_1571,In_16,In_195);
nand U1572 (N_1572,In_472,In_662);
or U1573 (N_1573,In_851,In_980);
nor U1574 (N_1574,In_880,In_750);
xor U1575 (N_1575,In_62,In_552);
nor U1576 (N_1576,In_640,In_772);
or U1577 (N_1577,In_781,In_630);
nand U1578 (N_1578,In_191,In_702);
and U1579 (N_1579,In_482,In_653);
or U1580 (N_1580,In_934,In_848);
or U1581 (N_1581,In_819,In_631);
nand U1582 (N_1582,In_833,In_387);
nand U1583 (N_1583,In_273,In_415);
and U1584 (N_1584,In_397,In_249);
or U1585 (N_1585,In_13,In_36);
nor U1586 (N_1586,In_355,In_507);
nand U1587 (N_1587,In_673,In_460);
or U1588 (N_1588,In_518,In_993);
nor U1589 (N_1589,In_840,In_467);
and U1590 (N_1590,In_753,In_343);
and U1591 (N_1591,In_20,In_804);
xnor U1592 (N_1592,In_274,In_194);
or U1593 (N_1593,In_96,In_202);
or U1594 (N_1594,In_673,In_749);
nand U1595 (N_1595,In_265,In_911);
and U1596 (N_1596,In_860,In_253);
or U1597 (N_1597,In_371,In_604);
and U1598 (N_1598,In_875,In_308);
or U1599 (N_1599,In_62,In_984);
and U1600 (N_1600,In_75,In_911);
nor U1601 (N_1601,In_829,In_30);
and U1602 (N_1602,In_714,In_559);
nand U1603 (N_1603,In_13,In_193);
nand U1604 (N_1604,In_14,In_501);
nor U1605 (N_1605,In_293,In_392);
nand U1606 (N_1606,In_568,In_997);
nand U1607 (N_1607,In_184,In_744);
or U1608 (N_1608,In_874,In_275);
or U1609 (N_1609,In_734,In_688);
and U1610 (N_1610,In_165,In_458);
nor U1611 (N_1611,In_700,In_937);
and U1612 (N_1612,In_965,In_889);
nand U1613 (N_1613,In_290,In_20);
xnor U1614 (N_1614,In_23,In_559);
and U1615 (N_1615,In_31,In_5);
nor U1616 (N_1616,In_790,In_525);
nor U1617 (N_1617,In_146,In_93);
nor U1618 (N_1618,In_843,In_589);
or U1619 (N_1619,In_782,In_956);
or U1620 (N_1620,In_196,In_911);
nand U1621 (N_1621,In_924,In_576);
or U1622 (N_1622,In_787,In_324);
xnor U1623 (N_1623,In_601,In_517);
nand U1624 (N_1624,In_265,In_571);
nor U1625 (N_1625,In_532,In_921);
or U1626 (N_1626,In_748,In_269);
or U1627 (N_1627,In_787,In_824);
nand U1628 (N_1628,In_696,In_762);
or U1629 (N_1629,In_239,In_615);
or U1630 (N_1630,In_252,In_410);
or U1631 (N_1631,In_896,In_949);
or U1632 (N_1632,In_887,In_531);
nand U1633 (N_1633,In_29,In_143);
nor U1634 (N_1634,In_205,In_864);
xnor U1635 (N_1635,In_249,In_671);
nor U1636 (N_1636,In_386,In_767);
and U1637 (N_1637,In_285,In_74);
and U1638 (N_1638,In_798,In_364);
nor U1639 (N_1639,In_953,In_125);
nor U1640 (N_1640,In_374,In_481);
and U1641 (N_1641,In_888,In_734);
or U1642 (N_1642,In_182,In_895);
and U1643 (N_1643,In_997,In_233);
and U1644 (N_1644,In_816,In_364);
xnor U1645 (N_1645,In_291,In_31);
nor U1646 (N_1646,In_464,In_13);
and U1647 (N_1647,In_32,In_230);
or U1648 (N_1648,In_207,In_196);
and U1649 (N_1649,In_136,In_822);
or U1650 (N_1650,In_642,In_640);
or U1651 (N_1651,In_87,In_385);
or U1652 (N_1652,In_804,In_109);
nor U1653 (N_1653,In_403,In_890);
nor U1654 (N_1654,In_799,In_937);
or U1655 (N_1655,In_888,In_52);
nand U1656 (N_1656,In_292,In_312);
nor U1657 (N_1657,In_665,In_440);
nand U1658 (N_1658,In_597,In_820);
and U1659 (N_1659,In_557,In_361);
and U1660 (N_1660,In_345,In_114);
or U1661 (N_1661,In_911,In_692);
nand U1662 (N_1662,In_342,In_388);
nor U1663 (N_1663,In_463,In_27);
nand U1664 (N_1664,In_550,In_326);
or U1665 (N_1665,In_645,In_125);
nand U1666 (N_1666,In_602,In_184);
nor U1667 (N_1667,In_397,In_264);
nor U1668 (N_1668,In_932,In_586);
and U1669 (N_1669,In_648,In_927);
and U1670 (N_1670,In_513,In_213);
nor U1671 (N_1671,In_74,In_611);
or U1672 (N_1672,In_85,In_620);
or U1673 (N_1673,In_365,In_235);
nor U1674 (N_1674,In_15,In_668);
nor U1675 (N_1675,In_33,In_116);
nor U1676 (N_1676,In_882,In_132);
nand U1677 (N_1677,In_212,In_631);
nand U1678 (N_1678,In_887,In_970);
and U1679 (N_1679,In_820,In_940);
nand U1680 (N_1680,In_235,In_234);
or U1681 (N_1681,In_309,In_385);
nand U1682 (N_1682,In_133,In_554);
and U1683 (N_1683,In_8,In_451);
or U1684 (N_1684,In_273,In_525);
nor U1685 (N_1685,In_263,In_181);
xor U1686 (N_1686,In_879,In_519);
xor U1687 (N_1687,In_932,In_425);
or U1688 (N_1688,In_801,In_925);
and U1689 (N_1689,In_646,In_377);
nand U1690 (N_1690,In_352,In_426);
xor U1691 (N_1691,In_159,In_901);
nor U1692 (N_1692,In_631,In_117);
and U1693 (N_1693,In_967,In_271);
nand U1694 (N_1694,In_697,In_726);
or U1695 (N_1695,In_543,In_420);
or U1696 (N_1696,In_294,In_166);
nand U1697 (N_1697,In_12,In_760);
or U1698 (N_1698,In_912,In_888);
nand U1699 (N_1699,In_671,In_319);
nand U1700 (N_1700,In_328,In_216);
or U1701 (N_1701,In_995,In_205);
or U1702 (N_1702,In_384,In_657);
and U1703 (N_1703,In_838,In_24);
nand U1704 (N_1704,In_914,In_670);
xnor U1705 (N_1705,In_433,In_379);
or U1706 (N_1706,In_24,In_16);
and U1707 (N_1707,In_834,In_254);
or U1708 (N_1708,In_254,In_559);
and U1709 (N_1709,In_22,In_178);
xor U1710 (N_1710,In_798,In_737);
nor U1711 (N_1711,In_936,In_470);
and U1712 (N_1712,In_591,In_701);
nor U1713 (N_1713,In_806,In_584);
nand U1714 (N_1714,In_19,In_310);
xnor U1715 (N_1715,In_631,In_683);
or U1716 (N_1716,In_121,In_170);
and U1717 (N_1717,In_20,In_730);
nor U1718 (N_1718,In_265,In_374);
or U1719 (N_1719,In_61,In_412);
nand U1720 (N_1720,In_889,In_692);
nor U1721 (N_1721,In_160,In_867);
or U1722 (N_1722,In_826,In_666);
nand U1723 (N_1723,In_747,In_390);
or U1724 (N_1724,In_971,In_596);
and U1725 (N_1725,In_684,In_825);
nor U1726 (N_1726,In_486,In_67);
xor U1727 (N_1727,In_857,In_315);
nor U1728 (N_1728,In_278,In_352);
nor U1729 (N_1729,In_616,In_886);
nand U1730 (N_1730,In_106,In_569);
or U1731 (N_1731,In_222,In_988);
and U1732 (N_1732,In_885,In_798);
and U1733 (N_1733,In_766,In_595);
nor U1734 (N_1734,In_569,In_277);
and U1735 (N_1735,In_512,In_577);
nor U1736 (N_1736,In_585,In_984);
nand U1737 (N_1737,In_507,In_154);
and U1738 (N_1738,In_539,In_536);
nor U1739 (N_1739,In_216,In_673);
nor U1740 (N_1740,In_71,In_326);
and U1741 (N_1741,In_634,In_232);
nor U1742 (N_1742,In_952,In_792);
and U1743 (N_1743,In_168,In_170);
nor U1744 (N_1744,In_676,In_495);
or U1745 (N_1745,In_326,In_647);
or U1746 (N_1746,In_609,In_481);
and U1747 (N_1747,In_783,In_427);
nand U1748 (N_1748,In_492,In_398);
nor U1749 (N_1749,In_982,In_619);
and U1750 (N_1750,In_172,In_988);
nor U1751 (N_1751,In_891,In_883);
or U1752 (N_1752,In_540,In_426);
nand U1753 (N_1753,In_465,In_58);
and U1754 (N_1754,In_23,In_15);
nand U1755 (N_1755,In_524,In_958);
nor U1756 (N_1756,In_181,In_277);
or U1757 (N_1757,In_192,In_211);
and U1758 (N_1758,In_46,In_798);
xor U1759 (N_1759,In_674,In_565);
nor U1760 (N_1760,In_193,In_672);
and U1761 (N_1761,In_973,In_821);
nor U1762 (N_1762,In_703,In_39);
nor U1763 (N_1763,In_350,In_923);
nand U1764 (N_1764,In_747,In_355);
xor U1765 (N_1765,In_488,In_389);
or U1766 (N_1766,In_929,In_667);
or U1767 (N_1767,In_668,In_959);
or U1768 (N_1768,In_221,In_376);
nor U1769 (N_1769,In_382,In_585);
and U1770 (N_1770,In_452,In_275);
and U1771 (N_1771,In_682,In_469);
nand U1772 (N_1772,In_813,In_137);
or U1773 (N_1773,In_606,In_814);
or U1774 (N_1774,In_614,In_276);
nor U1775 (N_1775,In_314,In_412);
nand U1776 (N_1776,In_413,In_538);
xnor U1777 (N_1777,In_530,In_644);
nor U1778 (N_1778,In_314,In_331);
xnor U1779 (N_1779,In_999,In_818);
nand U1780 (N_1780,In_983,In_588);
nor U1781 (N_1781,In_536,In_134);
and U1782 (N_1782,In_558,In_664);
and U1783 (N_1783,In_724,In_542);
nand U1784 (N_1784,In_739,In_488);
and U1785 (N_1785,In_408,In_588);
nor U1786 (N_1786,In_447,In_45);
nor U1787 (N_1787,In_746,In_564);
nor U1788 (N_1788,In_972,In_645);
and U1789 (N_1789,In_924,In_48);
or U1790 (N_1790,In_788,In_101);
or U1791 (N_1791,In_321,In_653);
or U1792 (N_1792,In_388,In_177);
or U1793 (N_1793,In_621,In_895);
or U1794 (N_1794,In_739,In_729);
nand U1795 (N_1795,In_187,In_664);
or U1796 (N_1796,In_618,In_366);
nand U1797 (N_1797,In_597,In_966);
and U1798 (N_1798,In_147,In_1);
or U1799 (N_1799,In_515,In_635);
nand U1800 (N_1800,In_84,In_849);
and U1801 (N_1801,In_849,In_975);
xnor U1802 (N_1802,In_498,In_214);
nand U1803 (N_1803,In_159,In_724);
and U1804 (N_1804,In_872,In_870);
and U1805 (N_1805,In_608,In_446);
or U1806 (N_1806,In_564,In_964);
nand U1807 (N_1807,In_704,In_528);
or U1808 (N_1808,In_292,In_129);
and U1809 (N_1809,In_638,In_535);
nor U1810 (N_1810,In_209,In_286);
or U1811 (N_1811,In_745,In_398);
and U1812 (N_1812,In_369,In_643);
and U1813 (N_1813,In_426,In_234);
xnor U1814 (N_1814,In_884,In_262);
nand U1815 (N_1815,In_240,In_993);
xnor U1816 (N_1816,In_71,In_203);
nor U1817 (N_1817,In_17,In_90);
or U1818 (N_1818,In_51,In_252);
nor U1819 (N_1819,In_794,In_725);
nor U1820 (N_1820,In_180,In_863);
nand U1821 (N_1821,In_870,In_766);
and U1822 (N_1822,In_584,In_469);
nor U1823 (N_1823,In_525,In_370);
nor U1824 (N_1824,In_365,In_433);
or U1825 (N_1825,In_451,In_6);
and U1826 (N_1826,In_307,In_464);
or U1827 (N_1827,In_361,In_743);
xor U1828 (N_1828,In_171,In_176);
xnor U1829 (N_1829,In_772,In_916);
nand U1830 (N_1830,In_724,In_329);
nor U1831 (N_1831,In_650,In_258);
nor U1832 (N_1832,In_864,In_9);
xnor U1833 (N_1833,In_42,In_246);
or U1834 (N_1834,In_876,In_115);
nand U1835 (N_1835,In_625,In_279);
nand U1836 (N_1836,In_810,In_925);
nand U1837 (N_1837,In_236,In_239);
nand U1838 (N_1838,In_31,In_929);
nor U1839 (N_1839,In_475,In_21);
nor U1840 (N_1840,In_792,In_357);
and U1841 (N_1841,In_724,In_319);
nor U1842 (N_1842,In_158,In_993);
xnor U1843 (N_1843,In_350,In_210);
nor U1844 (N_1844,In_425,In_38);
or U1845 (N_1845,In_192,In_113);
and U1846 (N_1846,In_796,In_602);
nand U1847 (N_1847,In_117,In_0);
and U1848 (N_1848,In_235,In_381);
nor U1849 (N_1849,In_321,In_610);
and U1850 (N_1850,In_782,In_338);
nand U1851 (N_1851,In_362,In_645);
or U1852 (N_1852,In_357,In_530);
nor U1853 (N_1853,In_159,In_312);
nand U1854 (N_1854,In_299,In_627);
or U1855 (N_1855,In_499,In_554);
nor U1856 (N_1856,In_262,In_676);
xnor U1857 (N_1857,In_174,In_843);
or U1858 (N_1858,In_593,In_557);
and U1859 (N_1859,In_605,In_498);
nor U1860 (N_1860,In_354,In_262);
nand U1861 (N_1861,In_61,In_556);
nor U1862 (N_1862,In_479,In_390);
and U1863 (N_1863,In_616,In_101);
and U1864 (N_1864,In_967,In_982);
and U1865 (N_1865,In_794,In_858);
nand U1866 (N_1866,In_151,In_560);
xnor U1867 (N_1867,In_295,In_610);
nor U1868 (N_1868,In_159,In_71);
nand U1869 (N_1869,In_527,In_699);
nand U1870 (N_1870,In_615,In_902);
and U1871 (N_1871,In_451,In_22);
or U1872 (N_1872,In_553,In_12);
nor U1873 (N_1873,In_526,In_964);
or U1874 (N_1874,In_198,In_496);
and U1875 (N_1875,In_665,In_460);
nor U1876 (N_1876,In_976,In_285);
and U1877 (N_1877,In_224,In_967);
nand U1878 (N_1878,In_918,In_468);
nor U1879 (N_1879,In_140,In_445);
xnor U1880 (N_1880,In_196,In_194);
nor U1881 (N_1881,In_709,In_663);
or U1882 (N_1882,In_653,In_368);
xnor U1883 (N_1883,In_613,In_457);
nor U1884 (N_1884,In_422,In_349);
and U1885 (N_1885,In_791,In_746);
and U1886 (N_1886,In_343,In_164);
nand U1887 (N_1887,In_0,In_742);
nor U1888 (N_1888,In_433,In_844);
nand U1889 (N_1889,In_893,In_809);
or U1890 (N_1890,In_8,In_312);
or U1891 (N_1891,In_863,In_78);
nand U1892 (N_1892,In_996,In_628);
or U1893 (N_1893,In_441,In_454);
or U1894 (N_1894,In_13,In_27);
or U1895 (N_1895,In_93,In_384);
and U1896 (N_1896,In_833,In_20);
or U1897 (N_1897,In_954,In_144);
and U1898 (N_1898,In_641,In_228);
xor U1899 (N_1899,In_399,In_435);
nand U1900 (N_1900,In_119,In_13);
nand U1901 (N_1901,In_325,In_964);
nor U1902 (N_1902,In_573,In_411);
or U1903 (N_1903,In_448,In_999);
or U1904 (N_1904,In_227,In_324);
and U1905 (N_1905,In_389,In_534);
or U1906 (N_1906,In_191,In_873);
xnor U1907 (N_1907,In_111,In_587);
nor U1908 (N_1908,In_444,In_641);
and U1909 (N_1909,In_317,In_787);
and U1910 (N_1910,In_384,In_690);
or U1911 (N_1911,In_839,In_470);
or U1912 (N_1912,In_75,In_861);
and U1913 (N_1913,In_268,In_643);
and U1914 (N_1914,In_214,In_219);
and U1915 (N_1915,In_118,In_637);
and U1916 (N_1916,In_654,In_415);
nand U1917 (N_1917,In_511,In_425);
nand U1918 (N_1918,In_679,In_123);
nor U1919 (N_1919,In_390,In_933);
or U1920 (N_1920,In_705,In_310);
or U1921 (N_1921,In_193,In_217);
nand U1922 (N_1922,In_984,In_517);
and U1923 (N_1923,In_25,In_217);
nor U1924 (N_1924,In_801,In_946);
or U1925 (N_1925,In_507,In_472);
xor U1926 (N_1926,In_516,In_898);
and U1927 (N_1927,In_621,In_488);
nor U1928 (N_1928,In_872,In_51);
or U1929 (N_1929,In_257,In_629);
nand U1930 (N_1930,In_406,In_816);
nand U1931 (N_1931,In_98,In_381);
and U1932 (N_1932,In_751,In_484);
nor U1933 (N_1933,In_143,In_973);
or U1934 (N_1934,In_319,In_39);
and U1935 (N_1935,In_449,In_192);
nor U1936 (N_1936,In_445,In_578);
and U1937 (N_1937,In_958,In_43);
nor U1938 (N_1938,In_938,In_182);
or U1939 (N_1939,In_790,In_194);
or U1940 (N_1940,In_550,In_57);
and U1941 (N_1941,In_894,In_481);
or U1942 (N_1942,In_90,In_759);
nor U1943 (N_1943,In_527,In_24);
or U1944 (N_1944,In_421,In_752);
nor U1945 (N_1945,In_224,In_315);
or U1946 (N_1946,In_825,In_17);
or U1947 (N_1947,In_792,In_400);
and U1948 (N_1948,In_72,In_4);
or U1949 (N_1949,In_30,In_700);
or U1950 (N_1950,In_924,In_530);
nand U1951 (N_1951,In_780,In_156);
nand U1952 (N_1952,In_763,In_382);
nand U1953 (N_1953,In_960,In_147);
nor U1954 (N_1954,In_898,In_487);
and U1955 (N_1955,In_548,In_57);
or U1956 (N_1956,In_424,In_263);
nor U1957 (N_1957,In_601,In_79);
and U1958 (N_1958,In_141,In_356);
and U1959 (N_1959,In_114,In_910);
nand U1960 (N_1960,In_518,In_593);
nor U1961 (N_1961,In_655,In_552);
or U1962 (N_1962,In_860,In_992);
or U1963 (N_1963,In_958,In_450);
nor U1964 (N_1964,In_769,In_228);
nand U1965 (N_1965,In_932,In_712);
or U1966 (N_1966,In_377,In_427);
and U1967 (N_1967,In_351,In_579);
or U1968 (N_1968,In_372,In_167);
and U1969 (N_1969,In_656,In_929);
or U1970 (N_1970,In_525,In_271);
xor U1971 (N_1971,In_185,In_123);
or U1972 (N_1972,In_19,In_148);
and U1973 (N_1973,In_936,In_598);
or U1974 (N_1974,In_503,In_824);
nand U1975 (N_1975,In_264,In_30);
nor U1976 (N_1976,In_668,In_650);
nor U1977 (N_1977,In_813,In_66);
and U1978 (N_1978,In_40,In_954);
nor U1979 (N_1979,In_9,In_227);
or U1980 (N_1980,In_191,In_102);
xnor U1981 (N_1981,In_255,In_802);
or U1982 (N_1982,In_856,In_3);
nor U1983 (N_1983,In_650,In_107);
and U1984 (N_1984,In_971,In_986);
nand U1985 (N_1985,In_953,In_918);
or U1986 (N_1986,In_862,In_560);
or U1987 (N_1987,In_791,In_513);
or U1988 (N_1988,In_801,In_470);
and U1989 (N_1989,In_967,In_59);
nand U1990 (N_1990,In_833,In_738);
nand U1991 (N_1991,In_867,In_611);
nor U1992 (N_1992,In_406,In_41);
xnor U1993 (N_1993,In_119,In_96);
and U1994 (N_1994,In_839,In_942);
nand U1995 (N_1995,In_925,In_425);
nor U1996 (N_1996,In_535,In_825);
or U1997 (N_1997,In_558,In_581);
xor U1998 (N_1998,In_632,In_471);
or U1999 (N_1999,In_984,In_315);
or U2000 (N_2000,In_149,In_517);
xor U2001 (N_2001,In_670,In_175);
xnor U2002 (N_2002,In_398,In_541);
or U2003 (N_2003,In_950,In_87);
nor U2004 (N_2004,In_578,In_93);
nand U2005 (N_2005,In_605,In_330);
nand U2006 (N_2006,In_862,In_23);
nor U2007 (N_2007,In_612,In_299);
and U2008 (N_2008,In_741,In_266);
or U2009 (N_2009,In_471,In_573);
and U2010 (N_2010,In_309,In_619);
or U2011 (N_2011,In_135,In_170);
nand U2012 (N_2012,In_719,In_685);
nor U2013 (N_2013,In_11,In_390);
nor U2014 (N_2014,In_672,In_888);
and U2015 (N_2015,In_25,In_878);
or U2016 (N_2016,In_291,In_882);
and U2017 (N_2017,In_57,In_909);
nand U2018 (N_2018,In_970,In_91);
and U2019 (N_2019,In_75,In_436);
or U2020 (N_2020,In_531,In_232);
nor U2021 (N_2021,In_7,In_391);
nor U2022 (N_2022,In_971,In_76);
nor U2023 (N_2023,In_82,In_921);
or U2024 (N_2024,In_548,In_844);
nor U2025 (N_2025,In_751,In_157);
nor U2026 (N_2026,In_117,In_133);
xor U2027 (N_2027,In_937,In_395);
and U2028 (N_2028,In_751,In_818);
and U2029 (N_2029,In_438,In_763);
nand U2030 (N_2030,In_756,In_951);
nand U2031 (N_2031,In_577,In_926);
or U2032 (N_2032,In_678,In_834);
and U2033 (N_2033,In_722,In_886);
and U2034 (N_2034,In_489,In_101);
and U2035 (N_2035,In_793,In_302);
nor U2036 (N_2036,In_440,In_124);
and U2037 (N_2037,In_881,In_69);
and U2038 (N_2038,In_147,In_204);
or U2039 (N_2039,In_153,In_617);
nor U2040 (N_2040,In_206,In_104);
nand U2041 (N_2041,In_317,In_526);
nor U2042 (N_2042,In_75,In_442);
nor U2043 (N_2043,In_691,In_186);
or U2044 (N_2044,In_910,In_327);
xor U2045 (N_2045,In_2,In_228);
and U2046 (N_2046,In_557,In_601);
and U2047 (N_2047,In_461,In_242);
and U2048 (N_2048,In_63,In_963);
and U2049 (N_2049,In_104,In_616);
and U2050 (N_2050,In_217,In_74);
and U2051 (N_2051,In_134,In_981);
nand U2052 (N_2052,In_461,In_184);
and U2053 (N_2053,In_414,In_486);
and U2054 (N_2054,In_32,In_564);
nand U2055 (N_2055,In_95,In_260);
nor U2056 (N_2056,In_638,In_281);
nand U2057 (N_2057,In_955,In_175);
nor U2058 (N_2058,In_267,In_663);
nor U2059 (N_2059,In_46,In_968);
or U2060 (N_2060,In_487,In_944);
xnor U2061 (N_2061,In_955,In_88);
nand U2062 (N_2062,In_490,In_605);
nand U2063 (N_2063,In_373,In_392);
nand U2064 (N_2064,In_909,In_552);
or U2065 (N_2065,In_425,In_349);
nand U2066 (N_2066,In_969,In_821);
nand U2067 (N_2067,In_438,In_249);
and U2068 (N_2068,In_520,In_205);
xnor U2069 (N_2069,In_781,In_698);
xnor U2070 (N_2070,In_762,In_492);
nand U2071 (N_2071,In_243,In_692);
or U2072 (N_2072,In_404,In_738);
nor U2073 (N_2073,In_187,In_146);
and U2074 (N_2074,In_39,In_243);
or U2075 (N_2075,In_266,In_402);
xnor U2076 (N_2076,In_105,In_853);
and U2077 (N_2077,In_175,In_845);
and U2078 (N_2078,In_137,In_322);
nor U2079 (N_2079,In_164,In_455);
nor U2080 (N_2080,In_576,In_790);
nand U2081 (N_2081,In_286,In_338);
nor U2082 (N_2082,In_996,In_865);
and U2083 (N_2083,In_92,In_475);
and U2084 (N_2084,In_347,In_477);
xor U2085 (N_2085,In_52,In_610);
nor U2086 (N_2086,In_746,In_510);
or U2087 (N_2087,In_441,In_140);
or U2088 (N_2088,In_428,In_940);
or U2089 (N_2089,In_215,In_163);
or U2090 (N_2090,In_344,In_79);
nor U2091 (N_2091,In_132,In_442);
and U2092 (N_2092,In_842,In_340);
xnor U2093 (N_2093,In_376,In_489);
and U2094 (N_2094,In_181,In_954);
nand U2095 (N_2095,In_140,In_311);
and U2096 (N_2096,In_286,In_972);
nand U2097 (N_2097,In_334,In_754);
nand U2098 (N_2098,In_818,In_34);
or U2099 (N_2099,In_613,In_446);
nor U2100 (N_2100,In_347,In_375);
nor U2101 (N_2101,In_484,In_645);
or U2102 (N_2102,In_486,In_114);
or U2103 (N_2103,In_212,In_838);
nand U2104 (N_2104,In_411,In_143);
xnor U2105 (N_2105,In_352,In_607);
nor U2106 (N_2106,In_239,In_499);
xnor U2107 (N_2107,In_790,In_442);
nor U2108 (N_2108,In_401,In_40);
or U2109 (N_2109,In_30,In_592);
or U2110 (N_2110,In_779,In_731);
and U2111 (N_2111,In_275,In_468);
and U2112 (N_2112,In_854,In_638);
xnor U2113 (N_2113,In_315,In_885);
and U2114 (N_2114,In_146,In_246);
nand U2115 (N_2115,In_736,In_541);
nand U2116 (N_2116,In_660,In_250);
or U2117 (N_2117,In_60,In_791);
nor U2118 (N_2118,In_532,In_442);
or U2119 (N_2119,In_949,In_552);
nand U2120 (N_2120,In_903,In_440);
xnor U2121 (N_2121,In_231,In_487);
nand U2122 (N_2122,In_648,In_315);
nand U2123 (N_2123,In_425,In_387);
and U2124 (N_2124,In_529,In_594);
or U2125 (N_2125,In_46,In_881);
nand U2126 (N_2126,In_530,In_514);
or U2127 (N_2127,In_975,In_549);
and U2128 (N_2128,In_533,In_509);
and U2129 (N_2129,In_227,In_292);
nand U2130 (N_2130,In_747,In_490);
or U2131 (N_2131,In_651,In_394);
nand U2132 (N_2132,In_418,In_721);
nor U2133 (N_2133,In_422,In_952);
nand U2134 (N_2134,In_567,In_588);
xor U2135 (N_2135,In_465,In_801);
nand U2136 (N_2136,In_541,In_553);
nand U2137 (N_2137,In_125,In_822);
nor U2138 (N_2138,In_464,In_950);
nand U2139 (N_2139,In_495,In_535);
nand U2140 (N_2140,In_186,In_138);
and U2141 (N_2141,In_496,In_970);
xor U2142 (N_2142,In_556,In_73);
or U2143 (N_2143,In_195,In_35);
or U2144 (N_2144,In_874,In_836);
xnor U2145 (N_2145,In_730,In_711);
nor U2146 (N_2146,In_392,In_104);
nand U2147 (N_2147,In_198,In_196);
nand U2148 (N_2148,In_358,In_236);
nor U2149 (N_2149,In_579,In_850);
nor U2150 (N_2150,In_497,In_941);
or U2151 (N_2151,In_494,In_51);
xnor U2152 (N_2152,In_650,In_604);
nor U2153 (N_2153,In_268,In_396);
nand U2154 (N_2154,In_992,In_87);
or U2155 (N_2155,In_942,In_345);
or U2156 (N_2156,In_732,In_679);
or U2157 (N_2157,In_106,In_896);
or U2158 (N_2158,In_908,In_714);
or U2159 (N_2159,In_330,In_821);
or U2160 (N_2160,In_223,In_460);
nand U2161 (N_2161,In_758,In_553);
nor U2162 (N_2162,In_911,In_420);
or U2163 (N_2163,In_504,In_99);
nand U2164 (N_2164,In_481,In_761);
nor U2165 (N_2165,In_222,In_906);
nor U2166 (N_2166,In_967,In_928);
nor U2167 (N_2167,In_722,In_383);
xnor U2168 (N_2168,In_868,In_446);
nand U2169 (N_2169,In_966,In_492);
nor U2170 (N_2170,In_905,In_866);
or U2171 (N_2171,In_908,In_179);
nor U2172 (N_2172,In_827,In_237);
nand U2173 (N_2173,In_185,In_947);
nor U2174 (N_2174,In_260,In_421);
nor U2175 (N_2175,In_444,In_281);
nor U2176 (N_2176,In_658,In_723);
xor U2177 (N_2177,In_290,In_773);
or U2178 (N_2178,In_931,In_86);
nor U2179 (N_2179,In_835,In_10);
nor U2180 (N_2180,In_323,In_458);
nor U2181 (N_2181,In_771,In_605);
nor U2182 (N_2182,In_317,In_696);
nand U2183 (N_2183,In_637,In_562);
xnor U2184 (N_2184,In_892,In_307);
and U2185 (N_2185,In_510,In_192);
or U2186 (N_2186,In_225,In_698);
or U2187 (N_2187,In_549,In_709);
and U2188 (N_2188,In_293,In_828);
xnor U2189 (N_2189,In_155,In_168);
and U2190 (N_2190,In_738,In_573);
nand U2191 (N_2191,In_706,In_245);
xor U2192 (N_2192,In_84,In_101);
nor U2193 (N_2193,In_859,In_121);
and U2194 (N_2194,In_105,In_525);
nand U2195 (N_2195,In_781,In_470);
and U2196 (N_2196,In_789,In_490);
nand U2197 (N_2197,In_81,In_744);
nor U2198 (N_2198,In_177,In_439);
nand U2199 (N_2199,In_876,In_199);
nor U2200 (N_2200,In_661,In_487);
nor U2201 (N_2201,In_258,In_997);
or U2202 (N_2202,In_821,In_321);
and U2203 (N_2203,In_321,In_485);
nand U2204 (N_2204,In_784,In_316);
or U2205 (N_2205,In_268,In_614);
nor U2206 (N_2206,In_435,In_224);
and U2207 (N_2207,In_234,In_636);
and U2208 (N_2208,In_392,In_708);
or U2209 (N_2209,In_339,In_942);
nor U2210 (N_2210,In_637,In_580);
or U2211 (N_2211,In_431,In_587);
nor U2212 (N_2212,In_94,In_438);
xor U2213 (N_2213,In_110,In_391);
xor U2214 (N_2214,In_983,In_875);
or U2215 (N_2215,In_348,In_89);
nor U2216 (N_2216,In_327,In_665);
or U2217 (N_2217,In_191,In_285);
xor U2218 (N_2218,In_147,In_797);
or U2219 (N_2219,In_625,In_267);
nor U2220 (N_2220,In_260,In_529);
and U2221 (N_2221,In_381,In_271);
nor U2222 (N_2222,In_681,In_261);
and U2223 (N_2223,In_606,In_881);
nand U2224 (N_2224,In_149,In_243);
nor U2225 (N_2225,In_127,In_415);
nand U2226 (N_2226,In_850,In_721);
and U2227 (N_2227,In_831,In_363);
and U2228 (N_2228,In_796,In_963);
and U2229 (N_2229,In_389,In_915);
nor U2230 (N_2230,In_93,In_472);
nor U2231 (N_2231,In_933,In_355);
or U2232 (N_2232,In_720,In_526);
or U2233 (N_2233,In_913,In_847);
and U2234 (N_2234,In_73,In_392);
nor U2235 (N_2235,In_234,In_208);
and U2236 (N_2236,In_884,In_343);
nand U2237 (N_2237,In_756,In_648);
nor U2238 (N_2238,In_972,In_762);
xnor U2239 (N_2239,In_959,In_831);
or U2240 (N_2240,In_529,In_510);
or U2241 (N_2241,In_534,In_361);
nor U2242 (N_2242,In_737,In_13);
or U2243 (N_2243,In_115,In_102);
or U2244 (N_2244,In_479,In_502);
nor U2245 (N_2245,In_84,In_253);
or U2246 (N_2246,In_407,In_669);
or U2247 (N_2247,In_648,In_135);
nand U2248 (N_2248,In_841,In_596);
or U2249 (N_2249,In_69,In_508);
or U2250 (N_2250,In_648,In_414);
nand U2251 (N_2251,In_428,In_801);
or U2252 (N_2252,In_616,In_711);
or U2253 (N_2253,In_707,In_350);
nand U2254 (N_2254,In_359,In_191);
nand U2255 (N_2255,In_686,In_388);
nor U2256 (N_2256,In_637,In_962);
or U2257 (N_2257,In_349,In_874);
and U2258 (N_2258,In_42,In_961);
nor U2259 (N_2259,In_991,In_115);
or U2260 (N_2260,In_79,In_659);
nand U2261 (N_2261,In_715,In_620);
or U2262 (N_2262,In_770,In_800);
and U2263 (N_2263,In_507,In_23);
nand U2264 (N_2264,In_819,In_500);
or U2265 (N_2265,In_329,In_473);
nor U2266 (N_2266,In_984,In_211);
nor U2267 (N_2267,In_489,In_226);
and U2268 (N_2268,In_372,In_445);
nor U2269 (N_2269,In_553,In_11);
or U2270 (N_2270,In_386,In_53);
nor U2271 (N_2271,In_112,In_248);
or U2272 (N_2272,In_732,In_161);
nand U2273 (N_2273,In_200,In_965);
nand U2274 (N_2274,In_69,In_381);
or U2275 (N_2275,In_912,In_756);
nor U2276 (N_2276,In_196,In_727);
and U2277 (N_2277,In_969,In_581);
and U2278 (N_2278,In_19,In_130);
nand U2279 (N_2279,In_42,In_890);
nand U2280 (N_2280,In_965,In_437);
or U2281 (N_2281,In_702,In_114);
or U2282 (N_2282,In_477,In_62);
or U2283 (N_2283,In_100,In_107);
xnor U2284 (N_2284,In_57,In_873);
and U2285 (N_2285,In_862,In_890);
and U2286 (N_2286,In_112,In_49);
or U2287 (N_2287,In_428,In_789);
nand U2288 (N_2288,In_501,In_731);
and U2289 (N_2289,In_602,In_15);
and U2290 (N_2290,In_870,In_719);
and U2291 (N_2291,In_306,In_13);
or U2292 (N_2292,In_105,In_319);
and U2293 (N_2293,In_710,In_455);
and U2294 (N_2294,In_653,In_714);
nor U2295 (N_2295,In_899,In_38);
nor U2296 (N_2296,In_734,In_389);
or U2297 (N_2297,In_986,In_173);
or U2298 (N_2298,In_91,In_108);
and U2299 (N_2299,In_988,In_930);
nand U2300 (N_2300,In_625,In_463);
and U2301 (N_2301,In_929,In_636);
or U2302 (N_2302,In_764,In_248);
nor U2303 (N_2303,In_841,In_730);
or U2304 (N_2304,In_848,In_615);
or U2305 (N_2305,In_806,In_889);
xnor U2306 (N_2306,In_558,In_500);
nand U2307 (N_2307,In_135,In_407);
or U2308 (N_2308,In_400,In_218);
xor U2309 (N_2309,In_973,In_755);
or U2310 (N_2310,In_985,In_810);
or U2311 (N_2311,In_234,In_748);
or U2312 (N_2312,In_719,In_173);
and U2313 (N_2313,In_467,In_492);
nand U2314 (N_2314,In_99,In_191);
or U2315 (N_2315,In_34,In_177);
nand U2316 (N_2316,In_209,In_253);
and U2317 (N_2317,In_894,In_309);
xor U2318 (N_2318,In_286,In_823);
nor U2319 (N_2319,In_62,In_545);
or U2320 (N_2320,In_435,In_9);
nand U2321 (N_2321,In_790,In_662);
or U2322 (N_2322,In_39,In_423);
nor U2323 (N_2323,In_159,In_979);
nand U2324 (N_2324,In_201,In_544);
xnor U2325 (N_2325,In_295,In_356);
nand U2326 (N_2326,In_998,In_732);
and U2327 (N_2327,In_679,In_892);
nand U2328 (N_2328,In_825,In_77);
nand U2329 (N_2329,In_1,In_690);
or U2330 (N_2330,In_234,In_291);
and U2331 (N_2331,In_348,In_706);
nor U2332 (N_2332,In_255,In_742);
or U2333 (N_2333,In_343,In_949);
nand U2334 (N_2334,In_302,In_204);
nand U2335 (N_2335,In_554,In_261);
and U2336 (N_2336,In_972,In_452);
and U2337 (N_2337,In_316,In_303);
and U2338 (N_2338,In_267,In_642);
xnor U2339 (N_2339,In_873,In_999);
nor U2340 (N_2340,In_472,In_936);
xnor U2341 (N_2341,In_190,In_742);
nand U2342 (N_2342,In_305,In_813);
and U2343 (N_2343,In_798,In_773);
nand U2344 (N_2344,In_348,In_422);
or U2345 (N_2345,In_608,In_966);
nor U2346 (N_2346,In_743,In_263);
nor U2347 (N_2347,In_852,In_786);
nor U2348 (N_2348,In_620,In_848);
or U2349 (N_2349,In_476,In_536);
xor U2350 (N_2350,In_106,In_450);
and U2351 (N_2351,In_351,In_564);
and U2352 (N_2352,In_406,In_146);
or U2353 (N_2353,In_429,In_596);
nand U2354 (N_2354,In_34,In_734);
xor U2355 (N_2355,In_150,In_970);
nand U2356 (N_2356,In_277,In_194);
and U2357 (N_2357,In_329,In_558);
xnor U2358 (N_2358,In_141,In_498);
or U2359 (N_2359,In_155,In_550);
or U2360 (N_2360,In_466,In_879);
xnor U2361 (N_2361,In_84,In_207);
or U2362 (N_2362,In_381,In_229);
or U2363 (N_2363,In_277,In_629);
and U2364 (N_2364,In_768,In_502);
and U2365 (N_2365,In_843,In_904);
and U2366 (N_2366,In_102,In_791);
nor U2367 (N_2367,In_586,In_11);
nand U2368 (N_2368,In_700,In_59);
nor U2369 (N_2369,In_132,In_71);
and U2370 (N_2370,In_293,In_905);
or U2371 (N_2371,In_821,In_61);
xnor U2372 (N_2372,In_794,In_789);
nand U2373 (N_2373,In_177,In_853);
and U2374 (N_2374,In_351,In_405);
nand U2375 (N_2375,In_686,In_93);
nor U2376 (N_2376,In_175,In_467);
and U2377 (N_2377,In_722,In_347);
and U2378 (N_2378,In_799,In_678);
and U2379 (N_2379,In_739,In_975);
nand U2380 (N_2380,In_919,In_704);
or U2381 (N_2381,In_33,In_315);
or U2382 (N_2382,In_791,In_352);
or U2383 (N_2383,In_697,In_523);
xnor U2384 (N_2384,In_479,In_998);
and U2385 (N_2385,In_36,In_810);
and U2386 (N_2386,In_202,In_455);
and U2387 (N_2387,In_768,In_296);
or U2388 (N_2388,In_847,In_186);
or U2389 (N_2389,In_8,In_3);
or U2390 (N_2390,In_494,In_754);
and U2391 (N_2391,In_385,In_261);
nand U2392 (N_2392,In_548,In_17);
or U2393 (N_2393,In_687,In_75);
and U2394 (N_2394,In_674,In_200);
or U2395 (N_2395,In_268,In_767);
or U2396 (N_2396,In_230,In_525);
nor U2397 (N_2397,In_109,In_573);
or U2398 (N_2398,In_580,In_971);
or U2399 (N_2399,In_301,In_749);
nor U2400 (N_2400,In_683,In_212);
nor U2401 (N_2401,In_572,In_717);
nand U2402 (N_2402,In_20,In_532);
and U2403 (N_2403,In_48,In_830);
nor U2404 (N_2404,In_153,In_558);
nand U2405 (N_2405,In_148,In_701);
or U2406 (N_2406,In_970,In_506);
or U2407 (N_2407,In_907,In_484);
nand U2408 (N_2408,In_128,In_465);
and U2409 (N_2409,In_199,In_307);
nor U2410 (N_2410,In_200,In_534);
nor U2411 (N_2411,In_225,In_92);
nor U2412 (N_2412,In_39,In_126);
xor U2413 (N_2413,In_575,In_138);
and U2414 (N_2414,In_857,In_461);
or U2415 (N_2415,In_237,In_760);
and U2416 (N_2416,In_518,In_388);
nand U2417 (N_2417,In_7,In_198);
nor U2418 (N_2418,In_109,In_220);
nand U2419 (N_2419,In_288,In_917);
nand U2420 (N_2420,In_91,In_216);
or U2421 (N_2421,In_794,In_715);
xor U2422 (N_2422,In_244,In_645);
and U2423 (N_2423,In_807,In_765);
and U2424 (N_2424,In_466,In_65);
nand U2425 (N_2425,In_264,In_213);
or U2426 (N_2426,In_643,In_34);
and U2427 (N_2427,In_317,In_245);
nand U2428 (N_2428,In_479,In_532);
or U2429 (N_2429,In_263,In_337);
and U2430 (N_2430,In_379,In_75);
xnor U2431 (N_2431,In_505,In_981);
or U2432 (N_2432,In_388,In_256);
and U2433 (N_2433,In_771,In_131);
or U2434 (N_2434,In_334,In_546);
xnor U2435 (N_2435,In_621,In_158);
and U2436 (N_2436,In_419,In_845);
nand U2437 (N_2437,In_801,In_632);
or U2438 (N_2438,In_834,In_365);
or U2439 (N_2439,In_528,In_97);
or U2440 (N_2440,In_620,In_568);
and U2441 (N_2441,In_505,In_349);
nand U2442 (N_2442,In_295,In_403);
and U2443 (N_2443,In_79,In_480);
nand U2444 (N_2444,In_172,In_192);
nand U2445 (N_2445,In_603,In_100);
or U2446 (N_2446,In_699,In_119);
or U2447 (N_2447,In_934,In_929);
nor U2448 (N_2448,In_299,In_455);
nand U2449 (N_2449,In_601,In_789);
xnor U2450 (N_2450,In_258,In_303);
and U2451 (N_2451,In_517,In_805);
nand U2452 (N_2452,In_962,In_429);
xnor U2453 (N_2453,In_561,In_270);
nand U2454 (N_2454,In_606,In_258);
and U2455 (N_2455,In_70,In_589);
or U2456 (N_2456,In_31,In_976);
xor U2457 (N_2457,In_360,In_975);
xnor U2458 (N_2458,In_525,In_48);
or U2459 (N_2459,In_52,In_509);
nand U2460 (N_2460,In_907,In_138);
nand U2461 (N_2461,In_513,In_0);
nand U2462 (N_2462,In_131,In_955);
nor U2463 (N_2463,In_705,In_399);
and U2464 (N_2464,In_847,In_414);
and U2465 (N_2465,In_232,In_256);
nand U2466 (N_2466,In_98,In_226);
nand U2467 (N_2467,In_387,In_719);
nand U2468 (N_2468,In_441,In_863);
or U2469 (N_2469,In_188,In_272);
or U2470 (N_2470,In_344,In_600);
nand U2471 (N_2471,In_955,In_17);
nor U2472 (N_2472,In_455,In_724);
and U2473 (N_2473,In_946,In_616);
or U2474 (N_2474,In_744,In_409);
nor U2475 (N_2475,In_32,In_254);
xnor U2476 (N_2476,In_979,In_636);
nand U2477 (N_2477,In_98,In_779);
nor U2478 (N_2478,In_582,In_616);
and U2479 (N_2479,In_473,In_279);
nor U2480 (N_2480,In_643,In_237);
or U2481 (N_2481,In_639,In_79);
and U2482 (N_2482,In_166,In_681);
or U2483 (N_2483,In_775,In_544);
xor U2484 (N_2484,In_703,In_481);
nor U2485 (N_2485,In_758,In_339);
or U2486 (N_2486,In_23,In_66);
nand U2487 (N_2487,In_959,In_378);
xnor U2488 (N_2488,In_460,In_314);
nor U2489 (N_2489,In_536,In_809);
nand U2490 (N_2490,In_313,In_174);
nand U2491 (N_2491,In_594,In_259);
nor U2492 (N_2492,In_820,In_837);
or U2493 (N_2493,In_337,In_912);
or U2494 (N_2494,In_308,In_636);
and U2495 (N_2495,In_382,In_524);
nand U2496 (N_2496,In_952,In_166);
nor U2497 (N_2497,In_484,In_639);
nor U2498 (N_2498,In_666,In_156);
nor U2499 (N_2499,In_319,In_470);
and U2500 (N_2500,N_1296,N_2373);
or U2501 (N_2501,N_1270,N_1123);
nor U2502 (N_2502,N_2402,N_1);
nand U2503 (N_2503,N_117,N_2262);
nor U2504 (N_2504,N_1726,N_1260);
or U2505 (N_2505,N_837,N_873);
nand U2506 (N_2506,N_2050,N_2094);
or U2507 (N_2507,N_30,N_1680);
and U2508 (N_2508,N_313,N_1010);
or U2509 (N_2509,N_864,N_390);
or U2510 (N_2510,N_2256,N_2269);
and U2511 (N_2511,N_1429,N_27);
nor U2512 (N_2512,N_2039,N_466);
and U2513 (N_2513,N_1508,N_1178);
nand U2514 (N_2514,N_875,N_2212);
xor U2515 (N_2515,N_2489,N_1062);
and U2516 (N_2516,N_685,N_914);
or U2517 (N_2517,N_1399,N_1543);
or U2518 (N_2518,N_1819,N_274);
and U2519 (N_2519,N_1003,N_1836);
nand U2520 (N_2520,N_2183,N_2225);
nor U2521 (N_2521,N_2281,N_881);
xnor U2522 (N_2522,N_583,N_1762);
or U2523 (N_2523,N_2202,N_64);
nor U2524 (N_2524,N_2163,N_2497);
and U2525 (N_2525,N_1293,N_927);
or U2526 (N_2526,N_1306,N_2318);
or U2527 (N_2527,N_2321,N_306);
and U2528 (N_2528,N_2235,N_1714);
nand U2529 (N_2529,N_1636,N_2303);
nand U2530 (N_2530,N_36,N_188);
nor U2531 (N_2531,N_114,N_2081);
or U2532 (N_2532,N_868,N_421);
and U2533 (N_2533,N_15,N_1447);
nor U2534 (N_2534,N_1881,N_672);
nand U2535 (N_2535,N_1052,N_1326);
nor U2536 (N_2536,N_858,N_1491);
nor U2537 (N_2537,N_2315,N_1054);
or U2538 (N_2538,N_1461,N_998);
or U2539 (N_2539,N_1805,N_225);
xor U2540 (N_2540,N_1152,N_1803);
or U2541 (N_2541,N_369,N_2184);
or U2542 (N_2542,N_897,N_324);
nand U2543 (N_2543,N_2106,N_1316);
nand U2544 (N_2544,N_1251,N_2012);
nor U2545 (N_2545,N_609,N_2140);
and U2546 (N_2546,N_1320,N_1710);
and U2547 (N_2547,N_704,N_2372);
and U2548 (N_2548,N_1654,N_2358);
or U2549 (N_2549,N_1124,N_289);
or U2550 (N_2550,N_2125,N_2363);
or U2551 (N_2551,N_1332,N_162);
and U2552 (N_2552,N_1880,N_2241);
nand U2553 (N_2553,N_1741,N_625);
nand U2554 (N_2554,N_1263,N_979);
nand U2555 (N_2555,N_2267,N_980);
or U2556 (N_2556,N_911,N_1387);
or U2557 (N_2557,N_865,N_1892);
and U2558 (N_2558,N_286,N_295);
nor U2559 (N_2559,N_1191,N_1678);
xnor U2560 (N_2560,N_1267,N_544);
nor U2561 (N_2561,N_438,N_1451);
or U2562 (N_2562,N_165,N_1135);
nand U2563 (N_2563,N_794,N_1432);
nor U2564 (N_2564,N_456,N_1825);
or U2565 (N_2565,N_888,N_2131);
nand U2566 (N_2566,N_1896,N_614);
or U2567 (N_2567,N_1939,N_1347);
nor U2568 (N_2568,N_1905,N_167);
nor U2569 (N_2569,N_627,N_743);
nand U2570 (N_2570,N_2266,N_776);
xor U2571 (N_2571,N_1673,N_517);
nor U2572 (N_2572,N_17,N_807);
and U2573 (N_2573,N_359,N_1945);
nor U2574 (N_2574,N_1407,N_1978);
and U2575 (N_2575,N_370,N_1057);
or U2576 (N_2576,N_108,N_2056);
nor U2577 (N_2577,N_751,N_1583);
or U2578 (N_2578,N_2356,N_637);
or U2579 (N_2579,N_769,N_482);
nand U2580 (N_2580,N_1207,N_284);
and U2581 (N_2581,N_530,N_465);
or U2582 (N_2582,N_1318,N_1639);
or U2583 (N_2583,N_877,N_2434);
nor U2584 (N_2584,N_676,N_1291);
xor U2585 (N_2585,N_354,N_664);
xor U2586 (N_2586,N_132,N_1362);
and U2587 (N_2587,N_643,N_2197);
nor U2588 (N_2588,N_2189,N_1566);
nor U2589 (N_2589,N_512,N_1386);
or U2590 (N_2590,N_2139,N_1404);
nand U2591 (N_2591,N_1129,N_561);
nor U2592 (N_2592,N_2275,N_1088);
nor U2593 (N_2593,N_2117,N_1528);
or U2594 (N_2594,N_58,N_2066);
nand U2595 (N_2595,N_679,N_2157);
xor U2596 (N_2596,N_211,N_978);
and U2597 (N_2597,N_538,N_1145);
nand U2598 (N_2598,N_805,N_1984);
nor U2599 (N_2599,N_107,N_355);
or U2600 (N_2600,N_907,N_1609);
or U2601 (N_2601,N_1834,N_79);
nor U2602 (N_2602,N_1684,N_1554);
nand U2603 (N_2603,N_1952,N_101);
and U2604 (N_2604,N_548,N_608);
xnor U2605 (N_2605,N_700,N_812);
nand U2606 (N_2606,N_2098,N_2462);
or U2607 (N_2607,N_2188,N_1641);
nor U2608 (N_2608,N_2219,N_1338);
nor U2609 (N_2609,N_321,N_90);
nand U2610 (N_2610,N_2046,N_1465);
and U2611 (N_2611,N_1149,N_442);
nand U2612 (N_2612,N_1973,N_240);
or U2613 (N_2613,N_1630,N_641);
and U2614 (N_2614,N_1868,N_754);
and U2615 (N_2615,N_1243,N_65);
nor U2616 (N_2616,N_1108,N_2296);
nand U2617 (N_2617,N_1192,N_792);
or U2618 (N_2618,N_1174,N_66);
xnor U2619 (N_2619,N_537,N_1487);
and U2620 (N_2620,N_362,N_1891);
xor U2621 (N_2621,N_567,N_364);
nor U2622 (N_2622,N_305,N_1083);
and U2623 (N_2623,N_2377,N_2392);
or U2624 (N_2624,N_2343,N_596);
nor U2625 (N_2625,N_554,N_2232);
xor U2626 (N_2626,N_513,N_2437);
and U2627 (N_2627,N_533,N_2379);
and U2628 (N_2628,N_2146,N_1206);
and U2629 (N_2629,N_2319,N_32);
or U2630 (N_2630,N_425,N_692);
nor U2631 (N_2631,N_1948,N_981);
or U2632 (N_2632,N_126,N_1706);
nor U2633 (N_2633,N_1503,N_947);
or U2634 (N_2634,N_1220,N_1640);
nor U2635 (N_2635,N_1701,N_457);
or U2636 (N_2636,N_1979,N_531);
nand U2637 (N_2637,N_2082,N_252);
and U2638 (N_2638,N_1434,N_1685);
nand U2639 (N_2639,N_1278,N_149);
nand U2640 (N_2640,N_584,N_806);
nand U2641 (N_2641,N_1691,N_2419);
nand U2642 (N_2642,N_1466,N_228);
or U2643 (N_2643,N_1513,N_1713);
or U2644 (N_2644,N_1763,N_1959);
nand U2645 (N_2645,N_16,N_1764);
nand U2646 (N_2646,N_1065,N_2279);
and U2647 (N_2647,N_1828,N_291);
nor U2648 (N_2648,N_1228,N_952);
and U2649 (N_2649,N_777,N_655);
nor U2650 (N_2650,N_268,N_1662);
nand U2651 (N_2651,N_417,N_1468);
or U2652 (N_2652,N_1907,N_2313);
or U2653 (N_2653,N_322,N_1666);
nor U2654 (N_2654,N_118,N_8);
or U2655 (N_2655,N_2228,N_2078);
xor U2656 (N_2656,N_1275,N_1522);
xor U2657 (N_2657,N_883,N_633);
xor U2658 (N_2658,N_2052,N_2042);
nor U2659 (N_2659,N_1268,N_1344);
nor U2660 (N_2660,N_387,N_1481);
or U2661 (N_2661,N_1109,N_1148);
nor U2662 (N_2662,N_14,N_588);
xnor U2663 (N_2663,N_358,N_2484);
nor U2664 (N_2664,N_497,N_1046);
nor U2665 (N_2665,N_587,N_1817);
and U2666 (N_2666,N_1127,N_304);
nand U2667 (N_2667,N_1385,N_800);
or U2668 (N_2668,N_1951,N_1203);
nand U2669 (N_2669,N_866,N_136);
nor U2670 (N_2670,N_905,N_1122);
nand U2671 (N_2671,N_1163,N_1551);
nand U2672 (N_2672,N_190,N_904);
nor U2673 (N_2673,N_116,N_1738);
and U2674 (N_2674,N_2449,N_2160);
nor U2675 (N_2675,N_1180,N_1259);
and U2676 (N_2676,N_1564,N_2393);
or U2677 (N_2677,N_1971,N_2457);
and U2678 (N_2678,N_2499,N_176);
nand U2679 (N_2679,N_1589,N_2215);
nor U2680 (N_2680,N_1480,N_1657);
nand U2681 (N_2681,N_529,N_35);
or U2682 (N_2682,N_1297,N_2278);
and U2683 (N_2683,N_686,N_1168);
xnor U2684 (N_2684,N_765,N_652);
and U2685 (N_2685,N_1333,N_1169);
or U2686 (N_2686,N_1028,N_613);
or U2687 (N_2687,N_1443,N_995);
nand U2688 (N_2688,N_2209,N_2474);
or U2689 (N_2689,N_1223,N_180);
and U2690 (N_2690,N_948,N_224);
nand U2691 (N_2691,N_271,N_206);
or U2692 (N_2692,N_536,N_214);
nand U2693 (N_2693,N_1424,N_1492);
and U2694 (N_2694,N_479,N_1234);
nor U2695 (N_2695,N_504,N_183);
nor U2696 (N_2696,N_2331,N_78);
or U2697 (N_2697,N_760,N_1582);
or U2698 (N_2698,N_1911,N_372);
or U2699 (N_2699,N_612,N_2185);
nor U2700 (N_2700,N_2341,N_856);
or U2701 (N_2701,N_1674,N_1150);
or U2702 (N_2702,N_431,N_2247);
nor U2703 (N_2703,N_376,N_1839);
nand U2704 (N_2704,N_1693,N_436);
or U2705 (N_2705,N_467,N_2053);
nand U2706 (N_2706,N_576,N_1542);
nand U2707 (N_2707,N_133,N_2205);
nor U2708 (N_2708,N_1237,N_597);
nor U2709 (N_2709,N_1747,N_1970);
and U2710 (N_2710,N_1051,N_412);
and U2711 (N_2711,N_1705,N_1264);
or U2712 (N_2712,N_582,N_1077);
nand U2713 (N_2713,N_869,N_347);
or U2714 (N_2714,N_871,N_2451);
nand U2715 (N_2715,N_2427,N_96);
nor U2716 (N_2716,N_1627,N_2206);
nand U2717 (N_2717,N_1651,N_62);
or U2718 (N_2718,N_660,N_382);
and U2719 (N_2719,N_202,N_1692);
and U2720 (N_2720,N_1798,N_811);
and U2721 (N_2721,N_257,N_1754);
nand U2722 (N_2722,N_131,N_178);
nor U2723 (N_2723,N_1080,N_1374);
nor U2724 (N_2724,N_1687,N_1698);
and U2725 (N_2725,N_977,N_52);
and U2726 (N_2726,N_1906,N_1511);
and U2727 (N_2727,N_1777,N_1273);
nor U2728 (N_2728,N_2161,N_1111);
nand U2729 (N_2729,N_1142,N_303);
xor U2730 (N_2730,N_1408,N_3);
nand U2731 (N_2731,N_1548,N_1060);
xor U2732 (N_2732,N_486,N_262);
nor U2733 (N_2733,N_2348,N_1188);
nor U2734 (N_2734,N_2310,N_1716);
and U2735 (N_2735,N_1557,N_2062);
nand U2736 (N_2736,N_335,N_2481);
nor U2737 (N_2737,N_2011,N_768);
nor U2738 (N_2738,N_171,N_2420);
nor U2739 (N_2739,N_460,N_445);
or U2740 (N_2740,N_2468,N_265);
and U2741 (N_2741,N_1919,N_1201);
and U2742 (N_2742,N_254,N_2444);
and U2743 (N_2743,N_1717,N_192);
or U2744 (N_2744,N_199,N_846);
or U2745 (N_2745,N_661,N_1596);
nor U2746 (N_2746,N_2155,N_1889);
or U2747 (N_2747,N_1631,N_37);
or U2748 (N_2748,N_1027,N_1914);
or U2749 (N_2749,N_1982,N_1055);
or U2750 (N_2750,N_1894,N_323);
and U2751 (N_2751,N_1916,N_1531);
and U2752 (N_2752,N_1202,N_1755);
or U2753 (N_2753,N_1456,N_752);
nor U2754 (N_2754,N_352,N_1866);
and U2755 (N_2755,N_1025,N_1176);
xnor U2756 (N_2756,N_862,N_42);
nor U2757 (N_2757,N_1463,N_218);
xor U2758 (N_2758,N_51,N_1001);
nor U2759 (N_2759,N_1029,N_1814);
nand U2760 (N_2760,N_487,N_1421);
and U2761 (N_2761,N_1537,N_1658);
and U2762 (N_2762,N_933,N_1702);
or U2763 (N_2763,N_831,N_1329);
nor U2764 (N_2764,N_1298,N_922);
and U2765 (N_2765,N_1890,N_2471);
nand U2766 (N_2766,N_219,N_541);
nor U2767 (N_2767,N_522,N_1963);
xor U2768 (N_2768,N_1390,N_645);
nor U2769 (N_2769,N_1185,N_1784);
xor U2770 (N_2770,N_419,N_60);
nor U2771 (N_2771,N_1041,N_2108);
nor U2772 (N_2772,N_973,N_216);
or U2773 (N_2773,N_1858,N_1768);
and U2774 (N_2774,N_550,N_81);
or U2775 (N_2775,N_418,N_407);
or U2776 (N_2776,N_423,N_515);
and U2777 (N_2777,N_683,N_1356);
xnor U2778 (N_2778,N_647,N_982);
nand U2779 (N_2779,N_1138,N_971);
and U2780 (N_2780,N_745,N_1852);
nor U2781 (N_2781,N_1381,N_814);
and U2782 (N_2782,N_1821,N_70);
nor U2783 (N_2783,N_2065,N_1402);
nand U2784 (N_2784,N_1675,N_518);
or U2785 (N_2785,N_1622,N_737);
nand U2786 (N_2786,N_2021,N_1378);
or U2787 (N_2787,N_1024,N_1930);
nor U2788 (N_2788,N_706,N_2283);
or U2789 (N_2789,N_1056,N_1668);
or U2790 (N_2790,N_985,N_74);
or U2791 (N_2791,N_2493,N_2369);
and U2792 (N_2792,N_840,N_525);
nand U2793 (N_2793,N_2055,N_2043);
or U2794 (N_2794,N_1038,N_658);
and U2795 (N_2795,N_1996,N_1253);
and U2796 (N_2796,N_2110,N_112);
nor U2797 (N_2797,N_429,N_549);
nor U2798 (N_2798,N_2092,N_1807);
nand U2799 (N_2799,N_534,N_2249);
and U2800 (N_2800,N_241,N_2335);
nor U2801 (N_2801,N_1193,N_95);
xor U2802 (N_2802,N_1279,N_248);
and U2803 (N_2803,N_2041,N_2038);
or U2804 (N_2804,N_1249,N_950);
nand U2805 (N_2805,N_2273,N_2274);
nand U2806 (N_2806,N_2162,N_1885);
or U2807 (N_2807,N_2386,N_1290);
nor U2808 (N_2808,N_1783,N_1990);
or U2809 (N_2809,N_1183,N_899);
or U2810 (N_2810,N_1884,N_1966);
and U2811 (N_2811,N_33,N_1128);
nor U2812 (N_2812,N_1946,N_77);
or U2813 (N_2813,N_580,N_130);
and U2814 (N_2814,N_2251,N_2133);
nor U2815 (N_2815,N_1427,N_1863);
nand U2816 (N_2816,N_1954,N_1987);
nand U2817 (N_2817,N_1791,N_1216);
nand U2818 (N_2818,N_1092,N_2391);
nor U2819 (N_2819,N_638,N_1049);
xnor U2820 (N_2820,N_1796,N_1588);
nand U2821 (N_2821,N_1061,N_2009);
and U2822 (N_2822,N_441,N_1878);
nand U2823 (N_2823,N_2143,N_1815);
nor U2824 (N_2824,N_2291,N_602);
or U2825 (N_2825,N_2276,N_635);
or U2826 (N_2826,N_850,N_1559);
or U2827 (N_2827,N_2203,N_1442);
nor U2828 (N_2828,N_106,N_2399);
or U2829 (N_2829,N_1002,N_1526);
nor U2830 (N_2830,N_2192,N_1115);
or U2831 (N_2831,N_1400,N_1085);
nand U2832 (N_2832,N_795,N_636);
nor U2833 (N_2833,N_1350,N_1086);
or U2834 (N_2834,N_175,N_1625);
nand U2835 (N_2835,N_296,N_298);
and U2836 (N_2836,N_1078,N_728);
nor U2837 (N_2837,N_1575,N_375);
and U2838 (N_2838,N_1328,N_845);
nor U2839 (N_2839,N_2260,N_1567);
nor U2840 (N_2840,N_2349,N_1143);
or U2841 (N_2841,N_976,N_1585);
or U2842 (N_2842,N_1758,N_1883);
nor U2843 (N_2843,N_2079,N_586);
nand U2844 (N_2844,N_1156,N_1097);
and U2845 (N_2845,N_1039,N_2023);
xnor U2846 (N_2846,N_815,N_1139);
or U2847 (N_2847,N_1026,N_2230);
or U2848 (N_2848,N_1229,N_1428);
or U2849 (N_2849,N_150,N_270);
nand U2850 (N_2850,N_713,N_464);
or U2851 (N_2851,N_1794,N_2257);
or U2852 (N_2852,N_1426,N_349);
nand U2853 (N_2853,N_2271,N_40);
nand U2854 (N_2854,N_200,N_2180);
nand U2855 (N_2855,N_2304,N_1479);
or U2856 (N_2856,N_2159,N_1009);
or U2857 (N_2857,N_890,N_2416);
nand U2858 (N_2858,N_1597,N_1770);
and U2859 (N_2859,N_1226,N_185);
nor U2860 (N_2860,N_903,N_2365);
nor U2861 (N_2861,N_1909,N_337);
and U2862 (N_2862,N_1967,N_292);
nor U2863 (N_2863,N_440,N_689);
and U2864 (N_2864,N_2101,N_1255);
nor U2865 (N_2865,N_11,N_755);
and U2866 (N_2866,N_1147,N_1732);
and U2867 (N_2867,N_2355,N_1782);
or U2868 (N_2868,N_2049,N_793);
and U2869 (N_2869,N_2430,N_99);
or U2870 (N_2870,N_2494,N_1106);
or U2871 (N_2871,N_2436,N_524);
or U2872 (N_2872,N_1743,N_2147);
nand U2873 (N_2873,N_969,N_314);
and U2874 (N_2874,N_1239,N_88);
nand U2875 (N_2875,N_1493,N_1209);
and U2876 (N_2876,N_2177,N_2034);
and U2877 (N_2877,N_2044,N_1521);
or U2878 (N_2878,N_1934,N_2015);
or U2879 (N_2879,N_1496,N_2289);
nand U2880 (N_2880,N_341,N_119);
or U2881 (N_2881,N_264,N_2288);
or U2882 (N_2882,N_1227,N_1859);
and U2883 (N_2883,N_640,N_1118);
nand U2884 (N_2884,N_590,N_2408);
or U2885 (N_2885,N_480,N_509);
nor U2886 (N_2886,N_2145,N_1235);
nor U2887 (N_2887,N_1076,N_2483);
or U2888 (N_2888,N_1101,N_233);
xor U2889 (N_2889,N_2314,N_1765);
xnor U2890 (N_2890,N_671,N_1430);
xnor U2891 (N_2891,N_796,N_122);
or U2892 (N_2892,N_2467,N_2259);
nand U2893 (N_2893,N_1021,N_2020);
or U2894 (N_2894,N_2024,N_13);
nand U2895 (N_2895,N_2378,N_2317);
nor U2896 (N_2896,N_2253,N_898);
nor U2897 (N_2897,N_1471,N_622);
or U2898 (N_2898,N_1187,N_2074);
nor U2899 (N_2899,N_386,N_1126);
or U2900 (N_2900,N_1120,N_191);
xnor U2901 (N_2901,N_532,N_1353);
nand U2902 (N_2902,N_2120,N_2396);
or U2903 (N_2903,N_259,N_2401);
and U2904 (N_2904,N_2382,N_1960);
and U2905 (N_2905,N_61,N_680);
nor U2906 (N_2906,N_2099,N_1014);
nand U2907 (N_2907,N_1931,N_808);
nand U2908 (N_2908,N_2264,N_678);
or U2909 (N_2909,N_1044,N_1953);
nand U2910 (N_2910,N_791,N_1282);
or U2911 (N_2911,N_618,N_163);
or U2912 (N_2912,N_505,N_1565);
and U2913 (N_2913,N_1547,N_520);
or U2914 (N_2914,N_2223,N_246);
or U2915 (N_2915,N_1391,N_2018);
or U2916 (N_2916,N_2244,N_1198);
nand U2917 (N_2917,N_1766,N_575);
and U2918 (N_2918,N_1072,N_160);
and U2919 (N_2919,N_1327,N_1346);
nor U2920 (N_2920,N_506,N_2033);
nand U2921 (N_2921,N_1540,N_86);
and U2922 (N_2922,N_325,N_1269);
and U2923 (N_2923,N_1406,N_73);
xor U2924 (N_2924,N_521,N_987);
or U2925 (N_2925,N_1477,N_247);
and U2926 (N_2926,N_579,N_2433);
nand U2927 (N_2927,N_2102,N_707);
and U2928 (N_2928,N_253,N_889);
xor U2929 (N_2929,N_779,N_2193);
nand U2930 (N_2930,N_1992,N_1637);
nor U2931 (N_2931,N_2072,N_2429);
nor U2932 (N_2932,N_788,N_1215);
xnor U2933 (N_2933,N_139,N_892);
nor U2934 (N_2934,N_2178,N_1665);
nor U2935 (N_2935,N_2035,N_6);
and U2936 (N_2936,N_668,N_1438);
nor U2937 (N_2937,N_1898,N_508);
nand U2938 (N_2938,N_1162,N_401);
nor U2939 (N_2939,N_2004,N_490);
xnor U2940 (N_2940,N_2323,N_2026);
nand U2941 (N_2941,N_2347,N_1450);
and U2942 (N_2942,N_1319,N_1059);
nor U2943 (N_2943,N_953,N_1601);
or U2944 (N_2944,N_1265,N_1416);
nand U2945 (N_2945,N_1475,N_182);
xnor U2946 (N_2946,N_1200,N_475);
xor U2947 (N_2947,N_5,N_822);
nor U2948 (N_2948,N_957,N_1280);
nor U2949 (N_2949,N_2199,N_849);
nor U2950 (N_2950,N_930,N_377);
nand U2951 (N_2951,N_1112,N_740);
nand U2952 (N_2952,N_631,N_2261);
nor U2953 (N_2953,N_1310,N_825);
nand U2954 (N_2954,N_174,N_1167);
or U2955 (N_2955,N_1944,N_269);
nor U2956 (N_2956,N_766,N_1507);
xnor U2957 (N_2957,N_1047,N_1371);
nand U2958 (N_2958,N_2210,N_226);
or U2959 (N_2959,N_1283,N_2428);
and U2960 (N_2960,N_2421,N_1546);
or U2961 (N_2961,N_10,N_2353);
and U2962 (N_2962,N_1822,N_2479);
nor U2963 (N_2963,N_80,N_1494);
nor U2964 (N_2964,N_860,N_1423);
nand U2965 (N_2965,N_975,N_774);
and U2966 (N_2966,N_1617,N_2466);
or U2967 (N_2967,N_1394,N_2186);
or U2968 (N_2968,N_1608,N_2453);
nor U2969 (N_2969,N_2426,N_2057);
or U2970 (N_2970,N_1274,N_1572);
nand U2971 (N_2971,N_1802,N_278);
nand U2972 (N_2972,N_750,N_1130);
and U2973 (N_2973,N_207,N_28);
and U2974 (N_2974,N_1976,N_1355);
xnor U2975 (N_2975,N_2214,N_1418);
nor U2976 (N_2976,N_1855,N_705);
nand U2977 (N_2977,N_1336,N_1517);
xor U2978 (N_2978,N_699,N_109);
or U2979 (N_2979,N_1584,N_742);
or U2980 (N_2980,N_156,N_1231);
or U2981 (N_2981,N_483,N_2475);
and U2982 (N_2982,N_1037,N_523);
and U2983 (N_2983,N_2179,N_701);
nor U2984 (N_2984,N_272,N_997);
nand U2985 (N_2985,N_1082,N_1431);
or U2986 (N_2986,N_258,N_285);
or U2987 (N_2987,N_1562,N_848);
nor U2988 (N_2988,N_993,N_2263);
or U2989 (N_2989,N_917,N_626);
nor U2990 (N_2990,N_2224,N_315);
or U2991 (N_2991,N_1367,N_154);
nor U2992 (N_2992,N_569,N_2445);
nand U2993 (N_2993,N_1853,N_511);
nor U2994 (N_2994,N_1700,N_916);
and U2995 (N_2995,N_2051,N_255);
nand U2996 (N_2996,N_452,N_1727);
and U2997 (N_2997,N_1211,N_1022);
and U2998 (N_2998,N_453,N_1771);
nand U2999 (N_2999,N_499,N_166);
xnor U3000 (N_3000,N_2406,N_1131);
nor U3001 (N_3001,N_565,N_450);
nand U3002 (N_3002,N_1744,N_2351);
nor U3003 (N_3003,N_786,N_1682);
nor U3004 (N_3004,N_2334,N_634);
nor U3005 (N_3005,N_2472,N_1760);
or U3006 (N_3006,N_830,N_1530);
xnor U3007 (N_3007,N_243,N_437);
nand U3008 (N_3008,N_1560,N_2268);
nor U3009 (N_3009,N_1102,N_909);
nand U3010 (N_3010,N_642,N_1573);
nor U3011 (N_3011,N_552,N_836);
nor U3012 (N_3012,N_2150,N_2328);
or U3013 (N_3013,N_574,N_2405);
or U3014 (N_3014,N_2221,N_2447);
or U3015 (N_3015,N_1064,N_1393);
nor U3016 (N_3016,N_604,N_1594);
nand U3017 (N_3017,N_2171,N_2123);
xor U3018 (N_3018,N_1789,N_2299);
nor U3019 (N_3019,N_413,N_443);
nor U3020 (N_3020,N_47,N_1570);
nor U3021 (N_3021,N_2119,N_827);
and U3022 (N_3022,N_1420,N_1995);
nand U3023 (N_3023,N_1523,N_1236);
and U3024 (N_3024,N_1441,N_1529);
nor U3025 (N_3025,N_502,N_1373);
xor U3026 (N_3026,N_650,N_2285);
nor U3027 (N_3027,N_2217,N_623);
nor U3028 (N_3028,N_2272,N_94);
or U3029 (N_3029,N_628,N_1621);
and U3030 (N_3030,N_1190,N_1874);
and U3031 (N_3031,N_432,N_1832);
and U3032 (N_3032,N_801,N_852);
and U3033 (N_3033,N_2022,N_1224);
or U3034 (N_3034,N_2301,N_900);
and U3035 (N_3035,N_2415,N_1998);
nand U3036 (N_3036,N_2088,N_934);
nor U3037 (N_3037,N_1897,N_1904);
or U3038 (N_3038,N_1154,N_653);
or U3039 (N_3039,N_196,N_489);
nor U3040 (N_3040,N_1312,N_557);
nand U3041 (N_3041,N_1464,N_1170);
nand U3042 (N_3042,N_720,N_334);
and U3043 (N_3043,N_870,N_893);
or U3044 (N_3044,N_826,N_297);
nor U3045 (N_3045,N_1458,N_1460);
nand U3046 (N_3046,N_1715,N_2441);
and U3047 (N_3047,N_1107,N_670);
or U3048 (N_3048,N_857,N_1969);
nor U3049 (N_3049,N_113,N_2340);
xor U3050 (N_3050,N_543,N_1730);
and U3051 (N_3051,N_2337,N_2190);
and U3052 (N_3052,N_1900,N_2403);
nor U3053 (N_3053,N_1396,N_2460);
and U3054 (N_3054,N_1823,N_1797);
nor U3055 (N_3055,N_1864,N_592);
or U3056 (N_3056,N_115,N_874);
and U3057 (N_3057,N_984,N_682);
nor U3058 (N_3058,N_2093,N_2438);
nor U3059 (N_3059,N_838,N_1704);
nor U3060 (N_3060,N_1661,N_1724);
or U3061 (N_3061,N_20,N_55);
nor U3062 (N_3062,N_1376,N_802);
nor U3063 (N_3063,N_2002,N_2322);
nand U3064 (N_3064,N_238,N_2329);
nand U3065 (N_3065,N_2195,N_1292);
xnor U3066 (N_3066,N_2144,N_1829);
nand U3067 (N_3067,N_2149,N_2220);
and U3068 (N_3068,N_1739,N_1840);
nand U3069 (N_3069,N_473,N_581);
xnor U3070 (N_3070,N_919,N_389);
nand U3071 (N_3071,N_1071,N_124);
nor U3072 (N_3072,N_861,N_540);
and U3073 (N_3073,N_1923,N_1773);
and U3074 (N_3074,N_381,N_2422);
nor U3075 (N_3075,N_21,N_2118);
nand U3076 (N_3076,N_1590,N_1875);
or U3077 (N_3077,N_1030,N_2397);
or U3078 (N_3078,N_1246,N_2265);
nand U3079 (N_3079,N_2080,N_1469);
or U3080 (N_3080,N_212,N_208);
or U3081 (N_3081,N_1020,N_2114);
nand U3082 (N_3082,N_923,N_2016);
or U3083 (N_3083,N_703,N_610);
nor U3084 (N_3084,N_1079,N_151);
nand U3085 (N_3085,N_371,N_691);
or U3086 (N_3086,N_2384,N_2488);
nand U3087 (N_3087,N_1801,N_403);
and U3088 (N_3088,N_955,N_1865);
or U3089 (N_3089,N_1591,N_2003);
and U3090 (N_3090,N_128,N_46);
or U3091 (N_3091,N_378,N_1696);
or U3092 (N_3092,N_1699,N_1735);
and U3093 (N_3093,N_733,N_1956);
or U3094 (N_3094,N_834,N_427);
or U3095 (N_3095,N_491,N_213);
xor U3096 (N_3096,N_63,N_1315);
nor U3097 (N_3097,N_784,N_1436);
nand U3098 (N_3098,N_1040,N_876);
or U3099 (N_3099,N_994,N_336);
xor U3100 (N_3100,N_267,N_1091);
nor U3101 (N_3101,N_2005,N_2076);
or U3102 (N_3102,N_1616,N_2325);
nand U3103 (N_3103,N_462,N_2182);
nor U3104 (N_3104,N_693,N_1612);
nor U3105 (N_3105,N_1974,N_1354);
and U3106 (N_3106,N_1555,N_308);
nand U3107 (N_3107,N_1942,N_1140);
nand U3108 (N_3108,N_2435,N_1799);
and U3109 (N_3109,N_646,N_1655);
nor U3110 (N_3110,N_2174,N_1189);
xnor U3111 (N_3111,N_1532,N_1015);
or U3112 (N_3112,N_2395,N_730);
nand U3113 (N_3113,N_344,N_1117);
or U3114 (N_3114,N_332,N_798);
or U3115 (N_3115,N_1778,N_972);
or U3116 (N_3116,N_350,N_164);
or U3117 (N_3117,N_724,N_867);
nand U3118 (N_3118,N_463,N_1324);
and U3119 (N_3119,N_1734,N_2496);
nor U3120 (N_3120,N_2246,N_134);
nor U3121 (N_3121,N_621,N_363);
and U3122 (N_3122,N_2073,N_288);
nor U3123 (N_3123,N_908,N_1177);
or U3124 (N_3124,N_501,N_1248);
or U3125 (N_3125,N_2332,N_2109);
and U3126 (N_3126,N_1595,N_785);
nand U3127 (N_3127,N_1314,N_2170);
nor U3128 (N_3128,N_1645,N_406);
or U3129 (N_3129,N_2007,N_1437);
and U3130 (N_3130,N_312,N_726);
nand U3131 (N_3131,N_1756,N_1094);
nor U3132 (N_3132,N_1070,N_1213);
and U3133 (N_3133,N_1459,N_57);
xnor U3134 (N_3134,N_1409,N_2476);
nand U3135 (N_3135,N_1670,N_1949);
or U3136 (N_3136,N_121,N_170);
nor U3137 (N_3137,N_1633,N_1786);
nor U3138 (N_3138,N_1938,N_1034);
nand U3139 (N_3139,N_277,N_2107);
nand U3140 (N_3140,N_669,N_1197);
nor U3141 (N_3141,N_1516,N_2309);
nor U3142 (N_3142,N_434,N_809);
and U3143 (N_3143,N_2019,N_2067);
nor U3144 (N_3144,N_144,N_790);
nor U3145 (N_3145,N_395,N_946);
nand U3146 (N_3146,N_391,N_85);
and U3147 (N_3147,N_1604,N_1417);
or U3148 (N_3148,N_1488,N_527);
and U3149 (N_3149,N_311,N_1068);
nor U3150 (N_3150,N_1016,N_863);
nand U3151 (N_3151,N_2213,N_1067);
and U3152 (N_3152,N_477,N_1256);
xor U3153 (N_3153,N_2130,N_1181);
nor U3154 (N_3154,N_1000,N_539);
or U3155 (N_3155,N_924,N_965);
nand U3156 (N_3156,N_968,N_573);
nor U3157 (N_3157,N_1415,N_1499);
and U3158 (N_3158,N_1302,N_140);
or U3159 (N_3159,N_2366,N_944);
nor U3160 (N_3160,N_1910,N_1276);
and U3161 (N_3161,N_1618,N_235);
and U3162 (N_3162,N_1013,N_854);
or U3163 (N_3163,N_1238,N_819);
and U3164 (N_3164,N_1932,N_1697);
nand U3165 (N_3165,N_2103,N_367);
nor U3166 (N_3166,N_1876,N_1895);
and U3167 (N_3167,N_1780,N_839);
nand U3168 (N_3168,N_1448,N_198);
or U3169 (N_3169,N_87,N_1382);
or U3170 (N_3170,N_2409,N_1317);
nor U3171 (N_3171,N_1225,N_1957);
or U3172 (N_3172,N_2469,N_2032);
xor U3173 (N_3173,N_974,N_411);
and U3174 (N_3174,N_2167,N_1854);
and U3175 (N_3175,N_1955,N_2196);
and U3176 (N_3176,N_936,N_237);
and U3177 (N_3177,N_1790,N_76);
and U3178 (N_3178,N_910,N_2168);
xnor U3179 (N_3179,N_2362,N_962);
nand U3180 (N_3180,N_723,N_1304);
and U3181 (N_3181,N_138,N_2440);
nand U3182 (N_3182,N_2424,N_2135);
and U3183 (N_3183,N_1377,N_1043);
nor U3184 (N_3184,N_1800,N_1502);
nor U3185 (N_3185,N_476,N_1230);
nor U3186 (N_3186,N_1577,N_992);
or U3187 (N_3187,N_75,N_1624);
nor U3188 (N_3188,N_169,N_963);
and U3189 (N_3189,N_93,N_1389);
and U3190 (N_3190,N_415,N_789);
and U3191 (N_3191,N_353,N_1005);
nand U3192 (N_3192,N_912,N_1476);
and U3193 (N_3193,N_735,N_578);
nor U3194 (N_3194,N_1761,N_2132);
and U3195 (N_3195,N_1776,N_729);
xnor U3196 (N_3196,N_2112,N_2200);
and U3197 (N_3197,N_599,N_1849);
nor U3198 (N_3198,N_615,N_2360);
or U3199 (N_3199,N_722,N_835);
nor U3200 (N_3200,N_1988,N_1847);
nor U3201 (N_3201,N_159,N_1208);
and U3202 (N_3202,N_2122,N_1772);
nand U3203 (N_3203,N_1242,N_1096);
nor U3204 (N_3204,N_2326,N_2037);
and U3205 (N_3205,N_1812,N_2454);
nor U3206 (N_3206,N_256,N_989);
and U3207 (N_3207,N_104,N_2316);
nand U3208 (N_3208,N_696,N_891);
xor U3209 (N_3209,N_98,N_813);
and U3210 (N_3210,N_2237,N_681);
and U3211 (N_3211,N_1490,N_988);
nand U3212 (N_3212,N_665,N_2063);
and U3213 (N_3213,N_187,N_1708);
and U3214 (N_3214,N_496,N_1262);
nand U3215 (N_3215,N_551,N_771);
or U3216 (N_3216,N_1598,N_1470);
nand U3217 (N_3217,N_503,N_1341);
or U3218 (N_3218,N_155,N_2354);
nand U3219 (N_3219,N_1848,N_990);
xnor U3220 (N_3220,N_342,N_1844);
and U3221 (N_3221,N_111,N_894);
nand U3222 (N_3222,N_1364,N_222);
nor U3223 (N_3223,N_1553,N_2394);
or U3224 (N_3224,N_1258,N_1087);
nand U3225 (N_3225,N_1520,N_1411);
or U3226 (N_3226,N_1751,N_1244);
xnor U3227 (N_3227,N_632,N_2456);
or U3228 (N_3228,N_1455,N_405);
nor U3229 (N_3229,N_702,N_731);
or U3230 (N_3230,N_1686,N_161);
nand U3231 (N_3231,N_331,N_1599);
nand U3232 (N_3232,N_2128,N_775);
nor U3233 (N_3233,N_2077,N_45);
nor U3234 (N_3234,N_507,N_1550);
nor U3235 (N_3235,N_2418,N_1349);
nand U3236 (N_3236,N_1222,N_422);
and U3237 (N_3237,N_2485,N_158);
nand U3238 (N_3238,N_145,N_439);
or U3239 (N_3239,N_767,N_2001);
nand U3240 (N_3240,N_2387,N_1011);
and U3241 (N_3241,N_662,N_230);
nor U3242 (N_3242,N_1372,N_2061);
nand U3243 (N_3243,N_181,N_1642);
or U3244 (N_3244,N_478,N_474);
nand U3245 (N_3245,N_1989,N_886);
nor U3246 (N_3246,N_374,N_1842);
nand U3247 (N_3247,N_2006,N_2463);
or U3248 (N_3248,N_2111,N_2308);
nand U3249 (N_3249,N_940,N_1157);
and U3250 (N_3250,N_1482,N_1921);
and U3251 (N_3251,N_2226,N_1742);
nor U3252 (N_3252,N_2000,N_186);
or U3253 (N_3253,N_1250,N_841);
or U3254 (N_3254,N_1527,N_2025);
and U3255 (N_3255,N_1843,N_433);
and U3256 (N_3256,N_1991,N_300);
nand U3257 (N_3257,N_1050,N_595);
nand U3258 (N_3258,N_2207,N_2176);
xnor U3259 (N_3259,N_828,N_1136);
nor U3260 (N_3260,N_1781,N_1902);
or U3261 (N_3261,N_2194,N_1748);
or U3262 (N_3262,N_803,N_1592);
and U3263 (N_3263,N_1449,N_996);
nor U3264 (N_3264,N_1740,N_1787);
nor U3265 (N_3265,N_1105,N_203);
nor U3266 (N_3266,N_2352,N_1089);
nor U3267 (N_3267,N_2227,N_220);
nand U3268 (N_3268,N_1444,N_577);
or U3269 (N_3269,N_1379,N_1261);
nand U3270 (N_3270,N_666,N_2383);
and U3271 (N_3271,N_2216,N_2236);
and U3272 (N_3272,N_2013,N_757);
nor U3273 (N_3273,N_282,N_943);
nand U3274 (N_3274,N_1164,N_600);
xor U3275 (N_3275,N_2464,N_1722);
xor U3276 (N_3276,N_817,N_201);
and U3277 (N_3277,N_1484,N_1792);
or U3278 (N_3278,N_1873,N_594);
and U3279 (N_3279,N_2031,N_2311);
nand U3280 (N_3280,N_2346,N_172);
and U3281 (N_3281,N_1845,N_34);
nor U3282 (N_3282,N_2452,N_1830);
and U3283 (N_3283,N_1485,N_1019);
nand U3284 (N_3284,N_2104,N_545);
or U3285 (N_3285,N_2030,N_92);
nand U3286 (N_3286,N_772,N_67);
nor U3287 (N_3287,N_1915,N_1141);
xor U3288 (N_3288,N_684,N_1846);
and U3289 (N_3289,N_2370,N_1690);
xnor U3290 (N_3290,N_991,N_1694);
or U3291 (N_3291,N_1383,N_1968);
xor U3292 (N_3292,N_1144,N_2473);
or U3293 (N_3293,N_1746,N_2380);
and U3294 (N_3294,N_547,N_2191);
and U3295 (N_3295,N_1729,N_2134);
nor U3296 (N_3296,N_824,N_1361);
nand U3297 (N_3297,N_195,N_2431);
or U3298 (N_3298,N_1534,N_2231);
and U3299 (N_3299,N_2357,N_2439);
nor U3300 (N_3300,N_2115,N_428);
or U3301 (N_3301,N_2069,N_1023);
nor U3302 (N_3302,N_1928,N_142);
and U3303 (N_3303,N_1918,N_1860);
or U3304 (N_3304,N_1950,N_1737);
or U3305 (N_3305,N_326,N_1425);
or U3306 (N_3306,N_2068,N_1788);
and U3307 (N_3307,N_1605,N_1877);
nand U3308 (N_3308,N_1403,N_1663);
xor U3309 (N_3309,N_231,N_2070);
nand U3310 (N_3310,N_695,N_1232);
and U3311 (N_3311,N_2338,N_1495);
xnor U3312 (N_3312,N_1943,N_2327);
nor U3313 (N_3313,N_1677,N_2166);
nand U3314 (N_3314,N_1515,N_571);
nand U3315 (N_3315,N_1719,N_360);
xnor U3316 (N_3316,N_1733,N_1033);
and U3317 (N_3317,N_2064,N_328);
and U3318 (N_3318,N_717,N_2083);
or U3319 (N_3319,N_620,N_424);
nor U3320 (N_3320,N_451,N_2240);
nor U3321 (N_3321,N_931,N_1922);
and U3322 (N_3322,N_1453,N_1712);
and U3323 (N_3323,N_1414,N_317);
or U3324 (N_3324,N_39,N_2432);
and U3325 (N_3325,N_1133,N_1358);
or U3326 (N_3326,N_44,N_2054);
nor U3327 (N_3327,N_1348,N_2127);
or U3328 (N_3328,N_2097,N_1857);
and U3329 (N_3329,N_1750,N_141);
nor U3330 (N_3330,N_1936,N_2284);
or U3331 (N_3331,N_1257,N_558);
nand U3332 (N_3332,N_1506,N_942);
nor U3333 (N_3333,N_797,N_2495);
nor U3334 (N_3334,N_2367,N_951);
nor U3335 (N_3335,N_2404,N_1912);
or U3336 (N_3336,N_1870,N_379);
or U3337 (N_3337,N_1961,N_307);
nand U3338 (N_3338,N_674,N_1983);
nor U3339 (N_3339,N_1384,N_1288);
or U3340 (N_3340,N_1498,N_1769);
xnor U3341 (N_3341,N_1779,N_302);
or U3342 (N_3342,N_585,N_1311);
or U3343 (N_3343,N_2425,N_2295);
nor U3344 (N_3344,N_1218,N_773);
nor U3345 (N_3345,N_2470,N_1929);
nor U3346 (N_3346,N_928,N_1538);
or U3347 (N_3347,N_1165,N_329);
and U3348 (N_3348,N_1247,N_1084);
nand U3349 (N_3349,N_1940,N_2248);
or U3350 (N_3350,N_1035,N_275);
and U3351 (N_3351,N_1300,N_205);
nor U3352 (N_3352,N_2381,N_1667);
and U3353 (N_3353,N_718,N_83);
or U3354 (N_3354,N_215,N_1580);
nand U3355 (N_3355,N_1103,N_49);
or U3356 (N_3356,N_1804,N_639);
and U3357 (N_3357,N_2239,N_2412);
nand U3358 (N_3358,N_1820,N_878);
nor U3359 (N_3359,N_339,N_2400);
and U3360 (N_3360,N_1603,N_2448);
xor U3361 (N_3361,N_2255,N_1439);
and U3362 (N_3362,N_293,N_1339);
and U3363 (N_3363,N_97,N_1933);
nor U3364 (N_3364,N_54,N_1446);
or U3365 (N_3365,N_677,N_1721);
nor U3366 (N_3366,N_560,N_435);
and U3367 (N_3367,N_1472,N_29);
or U3368 (N_3368,N_492,N_2490);
or U3369 (N_3369,N_416,N_239);
or U3370 (N_3370,N_1074,N_2359);
and U3371 (N_3371,N_1676,N_519);
nor U3372 (N_3372,N_2477,N_383);
xnor U3373 (N_3373,N_667,N_844);
nand U3374 (N_3374,N_1160,N_2300);
or U3375 (N_3375,N_143,N_69);
nor U3376 (N_3376,N_2350,N_708);
or U3377 (N_3377,N_1638,N_959);
or U3378 (N_3378,N_711,N_2375);
nand U3379 (N_3379,N_366,N_1808);
nor U3380 (N_3380,N_1179,N_2153);
xnor U3381 (N_3381,N_2320,N_1767);
nor U3382 (N_3382,N_1578,N_1707);
nor U3383 (N_3383,N_1669,N_2487);
nor U3384 (N_3384,N_746,N_1917);
and U3385 (N_3385,N_1619,N_721);
nor U3386 (N_3386,N_2158,N_2086);
nor U3387 (N_3387,N_563,N_399);
and U3388 (N_3388,N_1184,N_310);
nand U3389 (N_3389,N_385,N_2204);
and U3390 (N_3390,N_709,N_896);
and U3391 (N_3391,N_309,N_430);
and U3392 (N_3392,N_1473,N_872);
xnor U3393 (N_3393,N_902,N_1545);
and U3394 (N_3394,N_2333,N_510);
and U3395 (N_3395,N_105,N_1110);
nor U3396 (N_3396,N_832,N_404);
or U3397 (N_3397,N_31,N_630);
nand U3398 (N_3398,N_1709,N_146);
xor U3399 (N_3399,N_261,N_1576);
nand U3400 (N_3400,N_18,N_2342);
xnor U3401 (N_3401,N_227,N_1558);
or U3402 (N_3402,N_528,N_1644);
nand U3403 (N_3403,N_2417,N_901);
and U3404 (N_3404,N_2040,N_110);
nand U3405 (N_3405,N_1941,N_1613);
and U3406 (N_3406,N_1587,N_1660);
or U3407 (N_3407,N_753,N_2172);
and U3408 (N_3408,N_2465,N_967);
nor U3409 (N_3409,N_408,N_127);
nor U3410 (N_3410,N_1901,N_1623);
or U3411 (N_3411,N_1295,N_1462);
nor U3412 (N_3412,N_273,N_1569);
and U3413 (N_3413,N_194,N_1972);
xor U3414 (N_3414,N_1795,N_1204);
nor U3415 (N_3415,N_2164,N_1611);
nor U3416 (N_3416,N_770,N_1869);
nand U3417 (N_3417,N_471,N_1602);
or U3418 (N_3418,N_2486,N_2121);
nor U3419 (N_3419,N_2361,N_1871);
and U3420 (N_3420,N_1175,N_756);
xnor U3421 (N_3421,N_656,N_1058);
or U3422 (N_3422,N_1116,N_1656);
and U3423 (N_3423,N_712,N_2211);
nand U3424 (N_3424,N_1549,N_1410);
nor U3425 (N_3425,N_1098,N_2234);
and U3426 (N_3426,N_1032,N_1161);
nor U3427 (N_3427,N_1571,N_1155);
and U3428 (N_3428,N_1370,N_2461);
nor U3429 (N_3429,N_1606,N_1081);
nor U3430 (N_3430,N_420,N_454);
or U3431 (N_3431,N_276,N_1301);
and U3432 (N_3432,N_1581,N_1245);
nor U3433 (N_3433,N_970,N_1533);
nor U3434 (N_3434,N_2312,N_958);
and U3435 (N_3435,N_1649,N_2085);
or U3436 (N_3436,N_23,N_999);
and U3437 (N_3437,N_1999,N_294);
xnor U3438 (N_3438,N_397,N_1628);
and U3439 (N_3439,N_414,N_675);
nand U3440 (N_3440,N_1063,N_778);
or U3441 (N_3441,N_591,N_694);
or U3442 (N_3442,N_727,N_500);
xor U3443 (N_3443,N_484,N_210);
nor U3444 (N_3444,N_2048,N_1614);
nand U3445 (N_3445,N_847,N_1856);
and U3446 (N_3446,N_1134,N_2169);
nand U3447 (N_3447,N_125,N_448);
xor U3448 (N_3448,N_2407,N_603);
xor U3449 (N_3449,N_2414,N_2492);
nand U3450 (N_3450,N_173,N_741);
nor U3451 (N_3451,N_251,N_2218);
xor U3452 (N_3452,N_2385,N_2293);
nor U3453 (N_3453,N_2258,N_920);
or U3454 (N_3454,N_823,N_2116);
nand U3455 (N_3455,N_1926,N_458);
and U3456 (N_3456,N_734,N_842);
and U3457 (N_3457,N_1993,N_1525);
nor U3458 (N_3458,N_816,N_2222);
or U3459 (N_3459,N_725,N_2058);
xnor U3460 (N_3460,N_148,N_1544);
xor U3461 (N_3461,N_818,N_1752);
nand U3462 (N_3462,N_2100,N_562);
nor U3463 (N_3463,N_56,N_1977);
and U3464 (N_3464,N_2233,N_1212);
and U3465 (N_3465,N_1357,N_949);
nor U3466 (N_3466,N_1749,N_2156);
nand U3467 (N_3467,N_68,N_345);
nor U3468 (N_3468,N_137,N_559);
nand U3469 (N_3469,N_925,N_1478);
nor U3470 (N_3470,N_189,N_59);
or U3471 (N_3471,N_25,N_859);
xor U3472 (N_3472,N_2090,N_1284);
and U3473 (N_3473,N_485,N_495);
xnor U3474 (N_3474,N_526,N_555);
and U3475 (N_3475,N_26,N_747);
xor U3476 (N_3476,N_1745,N_209);
or U3477 (N_3477,N_2047,N_1331);
nor U3478 (N_3478,N_1321,N_217);
and U3479 (N_3479,N_1075,N_2374);
and U3480 (N_3480,N_887,N_1908);
nand U3481 (N_3481,N_710,N_1369);
nand U3482 (N_3482,N_400,N_498);
nand U3483 (N_3483,N_1340,N_236);
or U3484 (N_3484,N_1309,N_91);
xor U3485 (N_3485,N_1277,N_426);
xor U3486 (N_3486,N_1720,N_2450);
nor U3487 (N_3487,N_956,N_983);
and U3488 (N_3488,N_1158,N_103);
nor U3489 (N_3489,N_1899,N_135);
xor U3490 (N_3490,N_1927,N_1287);
or U3491 (N_3491,N_1454,N_732);
xor U3492 (N_3492,N_1233,N_184);
or U3493 (N_3493,N_619,N_1352);
nand U3494 (N_3494,N_229,N_245);
nand U3495 (N_3495,N_394,N_1099);
nor U3496 (N_3496,N_1299,N_1422);
and U3497 (N_3497,N_960,N_1457);
xnor U3498 (N_3498,N_649,N_1536);
nand U3499 (N_3499,N_781,N_1672);
xnor U3500 (N_3500,N_1397,N_1664);
nand U3501 (N_3501,N_1294,N_2089);
or U3502 (N_3502,N_2087,N_2198);
nor U3503 (N_3503,N_1474,N_1806);
and U3504 (N_3504,N_1600,N_1574);
nand U3505 (N_3505,N_409,N_2154);
nor U3506 (N_3506,N_688,N_152);
and U3507 (N_3507,N_986,N_1634);
xor U3508 (N_3508,N_1947,N_384);
nor U3509 (N_3509,N_468,N_1008);
nor U3510 (N_3510,N_1964,N_1345);
and U3511 (N_3511,N_651,N_1629);
or U3512 (N_3512,N_204,N_1997);
nor U3513 (N_3513,N_1535,N_606);
or U3514 (N_3514,N_1395,N_223);
and U3515 (N_3515,N_780,N_2491);
nor U3516 (N_3516,N_1335,N_2364);
or U3517 (N_3517,N_1683,N_2270);
nor U3518 (N_3518,N_2368,N_393);
nor U3519 (N_3519,N_410,N_1100);
and U3520 (N_3520,N_2413,N_553);
or U3521 (N_3521,N_938,N_1615);
xnor U3522 (N_3522,N_1166,N_1252);
and U3523 (N_3523,N_605,N_455);
nand U3524 (N_3524,N_1586,N_1042);
or U3525 (N_3525,N_514,N_1816);
and U3526 (N_3526,N_2388,N_1467);
and U3527 (N_3527,N_853,N_715);
or U3528 (N_3528,N_147,N_1375);
or U3529 (N_3529,N_1392,N_1632);
nor U3530 (N_3530,N_921,N_1872);
and U3531 (N_3531,N_1303,N_1981);
nand U3532 (N_3532,N_697,N_564);
nor U3533 (N_3533,N_2277,N_2410);
nand U3534 (N_3534,N_48,N_657);
nor U3535 (N_3535,N_570,N_72);
and U3536 (N_3536,N_41,N_1886);
or U3537 (N_3537,N_357,N_396);
nor U3538 (N_3538,N_2142,N_494);
xnor U3539 (N_3539,N_459,N_446);
or U3540 (N_3540,N_855,N_279);
and U3541 (N_3541,N_221,N_1723);
nor U3542 (N_3542,N_1119,N_1882);
or U3543 (N_3543,N_913,N_1679);
or U3544 (N_3544,N_1893,N_234);
nand U3545 (N_3545,N_348,N_748);
nand U3546 (N_3546,N_1509,N_1095);
or U3547 (N_3547,N_1240,N_546);
nand U3548 (N_3548,N_2398,N_392);
nor U3549 (N_3549,N_1552,N_1199);
or U3550 (N_3550,N_1323,N_2294);
nand U3551 (N_3551,N_1541,N_1793);
nor U3552 (N_3552,N_1132,N_1271);
xnor U3553 (N_3553,N_1343,N_617);
and U3554 (N_3554,N_1659,N_2376);
and U3555 (N_3555,N_1433,N_749);
and U3556 (N_3556,N_351,N_380);
nand U3557 (N_3557,N_1031,N_954);
and U3558 (N_3558,N_1380,N_1401);
nor U3559 (N_3559,N_2148,N_915);
nand U3560 (N_3560,N_804,N_1635);
and U3561 (N_3561,N_2286,N_1217);
or U3562 (N_3562,N_783,N_1643);
and U3563 (N_3563,N_1325,N_2208);
or U3564 (N_3564,N_556,N_2344);
nor U3565 (N_3565,N_2137,N_2290);
nand U3566 (N_3566,N_2175,N_799);
and U3567 (N_3567,N_1689,N_1958);
nand U3568 (N_3568,N_1307,N_2390);
or U3569 (N_3569,N_2250,N_2498);
nand U3570 (N_3570,N_535,N_1980);
nor U3571 (N_3571,N_2027,N_1671);
nand U3572 (N_3572,N_461,N_2017);
and U3573 (N_3573,N_1137,N_939);
nand U3574 (N_3574,N_1153,N_43);
and U3575 (N_3575,N_719,N_7);
nand U3576 (N_3576,N_1489,N_1850);
nor U3577 (N_3577,N_763,N_648);
xnor U3578 (N_3578,N_1196,N_1861);
nand U3579 (N_3579,N_2336,N_1824);
or U3580 (N_3580,N_53,N_1505);
and U3581 (N_3581,N_2201,N_937);
or U3582 (N_3582,N_1007,N_644);
and U3583 (N_3583,N_1121,N_2187);
nand U3584 (N_3584,N_1975,N_1986);
or U3585 (N_3585,N_1241,N_1113);
xnor U3586 (N_3586,N_2136,N_1486);
or U3587 (N_3587,N_1759,N_1837);
xnor U3588 (N_3588,N_698,N_961);
nor U3589 (N_3589,N_1219,N_343);
and U3590 (N_3590,N_1648,N_820);
or U3591 (N_3591,N_193,N_2252);
and U3592 (N_3592,N_2280,N_1514);
or U3593 (N_3593,N_941,N_1826);
nor U3594 (N_3594,N_2446,N_2173);
and U3595 (N_3595,N_2036,N_966);
nor U3596 (N_3596,N_1405,N_488);
nor U3597 (N_3597,N_177,N_1913);
nand U3598 (N_3598,N_102,N_1388);
nand U3599 (N_3599,N_249,N_759);
and U3600 (N_3600,N_2138,N_1924);
or U3601 (N_3601,N_879,N_2298);
and U3602 (N_3602,N_1500,N_1313);
or U3603 (N_3603,N_895,N_1286);
nor U3604 (N_3604,N_330,N_2480);
nor U3605 (N_3605,N_71,N_1626);
nand U3606 (N_3606,N_1831,N_1090);
nand U3607 (N_3607,N_1398,N_1435);
or U3608 (N_3608,N_762,N_84);
xor U3609 (N_3609,N_624,N_1363);
nand U3610 (N_3610,N_616,N_346);
and U3611 (N_3611,N_572,N_1017);
nor U3612 (N_3612,N_1862,N_1888);
xnor U3613 (N_3613,N_2165,N_1186);
nand U3614 (N_3614,N_1412,N_1841);
or U3615 (N_3615,N_2324,N_0);
nand U3616 (N_3616,N_1593,N_1413);
nor U3617 (N_3617,N_1510,N_472);
nand U3618 (N_3618,N_1066,N_2010);
nor U3619 (N_3619,N_2181,N_929);
nand U3620 (N_3620,N_1653,N_833);
nand U3621 (N_3621,N_1818,N_1607);
nand U3622 (N_3622,N_250,N_1368);
and U3623 (N_3623,N_882,N_1563);
or U3624 (N_3624,N_469,N_821);
nand U3625 (N_3625,N_242,N_1114);
and U3626 (N_3626,N_1785,N_2243);
or U3627 (N_3627,N_593,N_601);
or U3628 (N_3628,N_2113,N_301);
or U3629 (N_3629,N_1561,N_906);
xnor U3630 (N_3630,N_2029,N_1337);
or U3631 (N_3631,N_179,N_1518);
and U3632 (N_3632,N_738,N_1359);
or U3633 (N_3633,N_782,N_2282);
and U3634 (N_3634,N_1334,N_884);
and U3635 (N_3635,N_1937,N_1835);
nor U3636 (N_3636,N_318,N_744);
nand U3637 (N_3637,N_338,N_687);
or U3638 (N_3638,N_1045,N_260);
and U3639 (N_3639,N_1221,N_1330);
or U3640 (N_3640,N_316,N_1053);
and U3641 (N_3641,N_153,N_589);
xnor U3642 (N_3642,N_611,N_2238);
xnor U3643 (N_3643,N_761,N_1004);
nand U3644 (N_3644,N_4,N_964);
nor U3645 (N_3645,N_2482,N_470);
nand U3646 (N_3646,N_1647,N_1366);
and U3647 (N_3647,N_1281,N_654);
or U3648 (N_3648,N_1305,N_89);
nor U3649 (N_3649,N_2242,N_1610);
or U3650 (N_3650,N_2014,N_19);
nand U3651 (N_3651,N_1452,N_2126);
and U3652 (N_3652,N_1753,N_516);
and U3653 (N_3653,N_598,N_1012);
nand U3654 (N_3654,N_2292,N_123);
nand U3655 (N_3655,N_1006,N_232);
and U3656 (N_3656,N_1879,N_2254);
nand U3657 (N_3657,N_1579,N_281);
nand U3658 (N_3658,N_736,N_283);
nor U3659 (N_3659,N_1736,N_481);
xnor U3660 (N_3660,N_629,N_1483);
xor U3661 (N_3661,N_24,N_1272);
or U3662 (N_3662,N_764,N_1254);
nor U3663 (N_3663,N_2245,N_299);
and U3664 (N_3664,N_716,N_2306);
or U3665 (N_3665,N_2455,N_1171);
nor U3666 (N_3666,N_2091,N_1867);
nor U3667 (N_3667,N_100,N_880);
nor U3668 (N_3668,N_398,N_673);
nor U3669 (N_3669,N_2060,N_120);
and U3670 (N_3670,N_2345,N_810);
or U3671 (N_3671,N_1965,N_2443);
nand U3672 (N_3672,N_659,N_280);
nor U3673 (N_3673,N_1652,N_2141);
or U3674 (N_3674,N_542,N_368);
nand U3675 (N_3675,N_739,N_1811);
and U3676 (N_3676,N_945,N_2084);
or U3677 (N_3677,N_1073,N_1159);
or U3678 (N_3678,N_935,N_168);
or U3679 (N_3679,N_2371,N_1360);
or U3680 (N_3680,N_1365,N_365);
nor U3681 (N_3681,N_320,N_1445);
or U3682 (N_3682,N_2478,N_1725);
or U3683 (N_3683,N_1851,N_22);
and U3684 (N_3684,N_758,N_287);
and U3685 (N_3685,N_1289,N_1810);
and U3686 (N_3686,N_1985,N_1695);
nand U3687 (N_3687,N_444,N_1504);
nor U3688 (N_3688,N_2459,N_1646);
and U3689 (N_3689,N_1827,N_82);
and U3690 (N_3690,N_2045,N_829);
or U3691 (N_3691,N_1195,N_340);
or U3692 (N_3692,N_2330,N_1342);
nand U3693 (N_3693,N_1173,N_388);
nor U3694 (N_3694,N_2,N_1775);
or U3695 (N_3695,N_1182,N_1205);
nor U3696 (N_3696,N_1650,N_2008);
or U3697 (N_3697,N_1018,N_244);
or U3698 (N_3698,N_2411,N_1711);
nor U3699 (N_3699,N_2442,N_2129);
or U3700 (N_3700,N_2124,N_1556);
nor U3701 (N_3701,N_333,N_2423);
nor U3702 (N_3702,N_1210,N_1757);
nor U3703 (N_3703,N_787,N_12);
or U3704 (N_3704,N_2297,N_402);
nor U3705 (N_3705,N_493,N_690);
nor U3706 (N_3706,N_843,N_1036);
nor U3707 (N_3707,N_9,N_1501);
nand U3708 (N_3708,N_1903,N_568);
nor U3709 (N_3709,N_1838,N_1512);
nor U3710 (N_3710,N_2305,N_2229);
and U3711 (N_3711,N_1568,N_356);
or U3712 (N_3712,N_1069,N_129);
or U3713 (N_3713,N_2095,N_361);
or U3714 (N_3714,N_447,N_1285);
nand U3715 (N_3715,N_2105,N_38);
nand U3716 (N_3716,N_1104,N_319);
or U3717 (N_3717,N_2096,N_2152);
and U3718 (N_3718,N_2151,N_918);
nor U3719 (N_3719,N_1351,N_263);
nand U3720 (N_3720,N_1994,N_1194);
xnor U3721 (N_3721,N_1419,N_1440);
or U3722 (N_3722,N_1214,N_2059);
or U3723 (N_3723,N_1920,N_1731);
nand U3724 (N_3724,N_1519,N_1146);
or U3725 (N_3725,N_607,N_2458);
nand U3726 (N_3726,N_1308,N_1833);
nor U3727 (N_3727,N_2339,N_2302);
nand U3728 (N_3728,N_1539,N_1887);
and U3729 (N_3729,N_1093,N_1718);
nand U3730 (N_3730,N_2287,N_266);
or U3731 (N_3731,N_851,N_566);
and U3732 (N_3732,N_327,N_1681);
or U3733 (N_3733,N_1172,N_1497);
xnor U3734 (N_3734,N_2075,N_1322);
and U3735 (N_3735,N_1935,N_714);
or U3736 (N_3736,N_50,N_2071);
or U3737 (N_3737,N_1728,N_197);
and U3738 (N_3738,N_2389,N_290);
or U3739 (N_3739,N_449,N_1620);
nand U3740 (N_3740,N_373,N_885);
nand U3741 (N_3741,N_1813,N_1125);
nor U3742 (N_3742,N_2028,N_663);
nand U3743 (N_3743,N_2307,N_1151);
nor U3744 (N_3744,N_1688,N_1266);
xnor U3745 (N_3745,N_157,N_1925);
or U3746 (N_3746,N_1962,N_1048);
and U3747 (N_3747,N_1774,N_926);
nor U3748 (N_3748,N_1524,N_1703);
nor U3749 (N_3749,N_1809,N_932);
or U3750 (N_3750,N_751,N_1087);
and U3751 (N_3751,N_64,N_1134);
nor U3752 (N_3752,N_2241,N_700);
xor U3753 (N_3753,N_1347,N_341);
or U3754 (N_3754,N_328,N_967);
and U3755 (N_3755,N_2260,N_1018);
and U3756 (N_3756,N_280,N_1404);
nand U3757 (N_3757,N_1852,N_903);
nor U3758 (N_3758,N_2241,N_1214);
and U3759 (N_3759,N_202,N_2404);
nand U3760 (N_3760,N_2449,N_1130);
and U3761 (N_3761,N_828,N_1819);
and U3762 (N_3762,N_603,N_1829);
or U3763 (N_3763,N_938,N_1957);
nor U3764 (N_3764,N_187,N_1122);
and U3765 (N_3765,N_381,N_242);
nor U3766 (N_3766,N_2078,N_1567);
nand U3767 (N_3767,N_654,N_886);
and U3768 (N_3768,N_2487,N_2305);
and U3769 (N_3769,N_807,N_1909);
nand U3770 (N_3770,N_1490,N_1001);
nor U3771 (N_3771,N_532,N_1785);
or U3772 (N_3772,N_2005,N_1910);
and U3773 (N_3773,N_94,N_2419);
nor U3774 (N_3774,N_30,N_2224);
and U3775 (N_3775,N_1124,N_2311);
and U3776 (N_3776,N_862,N_2421);
nor U3777 (N_3777,N_2217,N_183);
nand U3778 (N_3778,N_1730,N_1341);
nor U3779 (N_3779,N_328,N_2404);
nand U3780 (N_3780,N_1225,N_617);
or U3781 (N_3781,N_2439,N_2210);
nand U3782 (N_3782,N_663,N_1954);
or U3783 (N_3783,N_2037,N_431);
nand U3784 (N_3784,N_2045,N_1146);
nor U3785 (N_3785,N_1354,N_701);
nand U3786 (N_3786,N_2066,N_1425);
or U3787 (N_3787,N_2007,N_2006);
nand U3788 (N_3788,N_1303,N_587);
nand U3789 (N_3789,N_863,N_896);
nand U3790 (N_3790,N_1985,N_769);
or U3791 (N_3791,N_1343,N_2374);
xnor U3792 (N_3792,N_318,N_1732);
xnor U3793 (N_3793,N_1204,N_797);
or U3794 (N_3794,N_996,N_1115);
nand U3795 (N_3795,N_1514,N_194);
nor U3796 (N_3796,N_775,N_132);
nand U3797 (N_3797,N_1233,N_877);
nor U3798 (N_3798,N_2200,N_2016);
and U3799 (N_3799,N_1741,N_375);
and U3800 (N_3800,N_1159,N_725);
and U3801 (N_3801,N_2383,N_2094);
and U3802 (N_3802,N_645,N_61);
or U3803 (N_3803,N_455,N_1417);
nand U3804 (N_3804,N_477,N_497);
and U3805 (N_3805,N_2097,N_1473);
or U3806 (N_3806,N_2177,N_1808);
nand U3807 (N_3807,N_984,N_649);
or U3808 (N_3808,N_331,N_39);
and U3809 (N_3809,N_146,N_412);
or U3810 (N_3810,N_551,N_2157);
and U3811 (N_3811,N_747,N_1678);
nor U3812 (N_3812,N_834,N_1684);
and U3813 (N_3813,N_1866,N_1534);
or U3814 (N_3814,N_2166,N_557);
nor U3815 (N_3815,N_284,N_205);
and U3816 (N_3816,N_1945,N_272);
and U3817 (N_3817,N_1473,N_1433);
and U3818 (N_3818,N_2122,N_1508);
nand U3819 (N_3819,N_657,N_1273);
or U3820 (N_3820,N_1663,N_2377);
or U3821 (N_3821,N_732,N_121);
or U3822 (N_3822,N_1039,N_47);
nor U3823 (N_3823,N_663,N_280);
and U3824 (N_3824,N_1410,N_2186);
and U3825 (N_3825,N_454,N_61);
xnor U3826 (N_3826,N_221,N_585);
xnor U3827 (N_3827,N_874,N_1785);
and U3828 (N_3828,N_427,N_749);
nand U3829 (N_3829,N_329,N_1327);
nor U3830 (N_3830,N_182,N_30);
or U3831 (N_3831,N_623,N_2114);
nand U3832 (N_3832,N_532,N_122);
or U3833 (N_3833,N_769,N_1923);
or U3834 (N_3834,N_2405,N_554);
and U3835 (N_3835,N_1809,N_267);
and U3836 (N_3836,N_69,N_2377);
and U3837 (N_3837,N_858,N_944);
and U3838 (N_3838,N_2424,N_902);
nand U3839 (N_3839,N_2179,N_2412);
nand U3840 (N_3840,N_23,N_848);
nand U3841 (N_3841,N_333,N_1748);
xnor U3842 (N_3842,N_1493,N_2058);
nor U3843 (N_3843,N_1596,N_1327);
and U3844 (N_3844,N_1879,N_1655);
or U3845 (N_3845,N_298,N_1110);
or U3846 (N_3846,N_2007,N_1209);
nand U3847 (N_3847,N_942,N_197);
and U3848 (N_3848,N_2093,N_2467);
nand U3849 (N_3849,N_2352,N_1974);
or U3850 (N_3850,N_1162,N_1543);
and U3851 (N_3851,N_804,N_1702);
nand U3852 (N_3852,N_1081,N_1592);
or U3853 (N_3853,N_1767,N_1425);
or U3854 (N_3854,N_1801,N_104);
and U3855 (N_3855,N_880,N_2492);
and U3856 (N_3856,N_582,N_115);
nand U3857 (N_3857,N_29,N_375);
nor U3858 (N_3858,N_155,N_948);
and U3859 (N_3859,N_875,N_806);
and U3860 (N_3860,N_209,N_2248);
nand U3861 (N_3861,N_1292,N_1661);
nor U3862 (N_3862,N_1692,N_1176);
xor U3863 (N_3863,N_1021,N_357);
nand U3864 (N_3864,N_1501,N_787);
or U3865 (N_3865,N_516,N_831);
and U3866 (N_3866,N_840,N_838);
and U3867 (N_3867,N_141,N_852);
nor U3868 (N_3868,N_646,N_1498);
xnor U3869 (N_3869,N_60,N_2390);
nor U3870 (N_3870,N_1483,N_2481);
or U3871 (N_3871,N_153,N_2482);
or U3872 (N_3872,N_1311,N_958);
or U3873 (N_3873,N_1771,N_761);
or U3874 (N_3874,N_660,N_225);
or U3875 (N_3875,N_2466,N_1157);
nand U3876 (N_3876,N_179,N_2486);
and U3877 (N_3877,N_1011,N_1833);
and U3878 (N_3878,N_2094,N_807);
and U3879 (N_3879,N_14,N_417);
and U3880 (N_3880,N_741,N_1626);
or U3881 (N_3881,N_1888,N_1326);
nor U3882 (N_3882,N_1803,N_193);
nor U3883 (N_3883,N_1568,N_794);
nor U3884 (N_3884,N_798,N_1879);
and U3885 (N_3885,N_1671,N_1507);
nor U3886 (N_3886,N_837,N_1539);
or U3887 (N_3887,N_1871,N_1021);
nor U3888 (N_3888,N_918,N_1773);
nor U3889 (N_3889,N_2117,N_590);
and U3890 (N_3890,N_300,N_977);
or U3891 (N_3891,N_1123,N_936);
or U3892 (N_3892,N_1843,N_1460);
nor U3893 (N_3893,N_1522,N_1671);
and U3894 (N_3894,N_416,N_1879);
or U3895 (N_3895,N_10,N_694);
and U3896 (N_3896,N_2304,N_2475);
nor U3897 (N_3897,N_512,N_1441);
nor U3898 (N_3898,N_1073,N_2418);
nor U3899 (N_3899,N_2080,N_1302);
and U3900 (N_3900,N_1225,N_2413);
and U3901 (N_3901,N_478,N_1383);
and U3902 (N_3902,N_509,N_227);
or U3903 (N_3903,N_1220,N_1189);
nand U3904 (N_3904,N_1746,N_666);
nand U3905 (N_3905,N_1595,N_1019);
nor U3906 (N_3906,N_270,N_367);
and U3907 (N_3907,N_1625,N_2042);
nand U3908 (N_3908,N_654,N_1801);
or U3909 (N_3909,N_190,N_1925);
xnor U3910 (N_3910,N_248,N_1124);
xnor U3911 (N_3911,N_43,N_907);
nand U3912 (N_3912,N_389,N_2493);
or U3913 (N_3913,N_341,N_193);
and U3914 (N_3914,N_246,N_2409);
or U3915 (N_3915,N_1774,N_2403);
nand U3916 (N_3916,N_2435,N_1065);
or U3917 (N_3917,N_1065,N_1727);
nand U3918 (N_3918,N_1574,N_2293);
nand U3919 (N_3919,N_1297,N_790);
and U3920 (N_3920,N_17,N_1862);
and U3921 (N_3921,N_853,N_1360);
or U3922 (N_3922,N_2080,N_1285);
nor U3923 (N_3923,N_422,N_1571);
or U3924 (N_3924,N_109,N_2426);
nand U3925 (N_3925,N_697,N_1316);
xnor U3926 (N_3926,N_1685,N_251);
xnor U3927 (N_3927,N_1654,N_1774);
nor U3928 (N_3928,N_1664,N_330);
nor U3929 (N_3929,N_773,N_1872);
and U3930 (N_3930,N_2466,N_2005);
or U3931 (N_3931,N_17,N_2217);
and U3932 (N_3932,N_339,N_203);
xor U3933 (N_3933,N_2318,N_2187);
nand U3934 (N_3934,N_2132,N_2331);
nand U3935 (N_3935,N_1807,N_993);
or U3936 (N_3936,N_1892,N_1115);
nand U3937 (N_3937,N_128,N_668);
and U3938 (N_3938,N_803,N_1310);
and U3939 (N_3939,N_812,N_886);
xor U3940 (N_3940,N_107,N_763);
and U3941 (N_3941,N_2396,N_383);
and U3942 (N_3942,N_935,N_1067);
nand U3943 (N_3943,N_1675,N_2095);
and U3944 (N_3944,N_744,N_144);
xor U3945 (N_3945,N_683,N_348);
or U3946 (N_3946,N_1782,N_2138);
nor U3947 (N_3947,N_160,N_861);
or U3948 (N_3948,N_693,N_1241);
nor U3949 (N_3949,N_5,N_204);
and U3950 (N_3950,N_1777,N_756);
and U3951 (N_3951,N_1660,N_2193);
or U3952 (N_3952,N_832,N_1671);
nor U3953 (N_3953,N_1366,N_333);
and U3954 (N_3954,N_2425,N_534);
and U3955 (N_3955,N_29,N_1623);
and U3956 (N_3956,N_1846,N_1954);
nand U3957 (N_3957,N_2140,N_2386);
nand U3958 (N_3958,N_713,N_784);
or U3959 (N_3959,N_1641,N_2201);
nand U3960 (N_3960,N_516,N_4);
nor U3961 (N_3961,N_987,N_1849);
xnor U3962 (N_3962,N_440,N_2109);
and U3963 (N_3963,N_1340,N_1831);
and U3964 (N_3964,N_1780,N_1452);
xor U3965 (N_3965,N_808,N_696);
nor U3966 (N_3966,N_1898,N_1973);
nor U3967 (N_3967,N_2299,N_1538);
or U3968 (N_3968,N_271,N_1858);
and U3969 (N_3969,N_1976,N_1668);
nor U3970 (N_3970,N_2211,N_2206);
nand U3971 (N_3971,N_1987,N_579);
or U3972 (N_3972,N_1521,N_1539);
or U3973 (N_3973,N_819,N_551);
and U3974 (N_3974,N_1665,N_2336);
or U3975 (N_3975,N_857,N_2313);
and U3976 (N_3976,N_842,N_1616);
and U3977 (N_3977,N_2462,N_925);
or U3978 (N_3978,N_672,N_286);
nor U3979 (N_3979,N_1957,N_2466);
nor U3980 (N_3980,N_893,N_2216);
nand U3981 (N_3981,N_1422,N_1515);
and U3982 (N_3982,N_1776,N_577);
nand U3983 (N_3983,N_217,N_1451);
nand U3984 (N_3984,N_2190,N_1475);
nor U3985 (N_3985,N_1524,N_1482);
nor U3986 (N_3986,N_1679,N_1209);
nand U3987 (N_3987,N_2487,N_718);
or U3988 (N_3988,N_2397,N_425);
nor U3989 (N_3989,N_2314,N_1025);
nand U3990 (N_3990,N_1421,N_2432);
nand U3991 (N_3991,N_2499,N_2454);
nand U3992 (N_3992,N_1652,N_1668);
and U3993 (N_3993,N_1365,N_1427);
xnor U3994 (N_3994,N_1672,N_816);
or U3995 (N_3995,N_1163,N_2012);
or U3996 (N_3996,N_2377,N_1065);
nand U3997 (N_3997,N_2278,N_1444);
xnor U3998 (N_3998,N_1133,N_2232);
nand U3999 (N_3999,N_786,N_1510);
or U4000 (N_4000,N_2070,N_2453);
nor U4001 (N_4001,N_882,N_2173);
nand U4002 (N_4002,N_794,N_415);
xor U4003 (N_4003,N_1382,N_1562);
or U4004 (N_4004,N_2451,N_409);
xnor U4005 (N_4005,N_597,N_1302);
and U4006 (N_4006,N_218,N_69);
nor U4007 (N_4007,N_1966,N_967);
xor U4008 (N_4008,N_938,N_1585);
nand U4009 (N_4009,N_732,N_1633);
and U4010 (N_4010,N_211,N_586);
nand U4011 (N_4011,N_1130,N_23);
xnor U4012 (N_4012,N_644,N_1243);
xor U4013 (N_4013,N_1076,N_456);
nand U4014 (N_4014,N_526,N_2080);
or U4015 (N_4015,N_484,N_595);
and U4016 (N_4016,N_853,N_2101);
nor U4017 (N_4017,N_1095,N_1597);
nor U4018 (N_4018,N_213,N_12);
and U4019 (N_4019,N_926,N_1507);
and U4020 (N_4020,N_1921,N_295);
and U4021 (N_4021,N_630,N_774);
nor U4022 (N_4022,N_889,N_693);
or U4023 (N_4023,N_740,N_858);
nor U4024 (N_4024,N_1148,N_503);
nand U4025 (N_4025,N_451,N_2472);
nand U4026 (N_4026,N_46,N_677);
xor U4027 (N_4027,N_642,N_1610);
and U4028 (N_4028,N_625,N_413);
nor U4029 (N_4029,N_1744,N_520);
nand U4030 (N_4030,N_1664,N_1265);
or U4031 (N_4031,N_307,N_999);
and U4032 (N_4032,N_407,N_13);
nand U4033 (N_4033,N_511,N_2252);
or U4034 (N_4034,N_1696,N_2286);
nor U4035 (N_4035,N_2057,N_2422);
or U4036 (N_4036,N_1837,N_855);
and U4037 (N_4037,N_2007,N_135);
and U4038 (N_4038,N_1825,N_81);
xor U4039 (N_4039,N_1866,N_1187);
or U4040 (N_4040,N_1037,N_1350);
or U4041 (N_4041,N_679,N_1907);
and U4042 (N_4042,N_1373,N_832);
nor U4043 (N_4043,N_2062,N_2304);
xnor U4044 (N_4044,N_361,N_2323);
nand U4045 (N_4045,N_1595,N_2450);
nor U4046 (N_4046,N_358,N_730);
nand U4047 (N_4047,N_2417,N_1190);
and U4048 (N_4048,N_2289,N_1986);
nand U4049 (N_4049,N_200,N_1931);
or U4050 (N_4050,N_2493,N_367);
and U4051 (N_4051,N_1842,N_258);
nor U4052 (N_4052,N_132,N_2051);
nand U4053 (N_4053,N_1261,N_927);
nand U4054 (N_4054,N_2243,N_1520);
nand U4055 (N_4055,N_71,N_518);
or U4056 (N_4056,N_2248,N_772);
nand U4057 (N_4057,N_1693,N_983);
nand U4058 (N_4058,N_2337,N_1931);
nor U4059 (N_4059,N_2141,N_205);
nand U4060 (N_4060,N_1490,N_107);
nand U4061 (N_4061,N_2121,N_1140);
nor U4062 (N_4062,N_865,N_2048);
or U4063 (N_4063,N_1869,N_2241);
and U4064 (N_4064,N_2374,N_1901);
nor U4065 (N_4065,N_124,N_2);
nor U4066 (N_4066,N_251,N_1734);
or U4067 (N_4067,N_74,N_1652);
nor U4068 (N_4068,N_632,N_2321);
nand U4069 (N_4069,N_954,N_843);
or U4070 (N_4070,N_436,N_1336);
nor U4071 (N_4071,N_38,N_266);
or U4072 (N_4072,N_8,N_248);
xnor U4073 (N_4073,N_2461,N_1957);
nand U4074 (N_4074,N_720,N_1015);
and U4075 (N_4075,N_487,N_786);
xnor U4076 (N_4076,N_292,N_1691);
or U4077 (N_4077,N_315,N_1449);
and U4078 (N_4078,N_2123,N_2097);
nor U4079 (N_4079,N_1026,N_2427);
or U4080 (N_4080,N_1855,N_1987);
xnor U4081 (N_4081,N_278,N_2357);
nand U4082 (N_4082,N_470,N_1557);
nor U4083 (N_4083,N_2454,N_463);
nor U4084 (N_4084,N_1803,N_2239);
nor U4085 (N_4085,N_1609,N_2371);
or U4086 (N_4086,N_447,N_1038);
xor U4087 (N_4087,N_1417,N_1863);
and U4088 (N_4088,N_1593,N_239);
nor U4089 (N_4089,N_523,N_198);
and U4090 (N_4090,N_770,N_1888);
and U4091 (N_4091,N_419,N_1770);
nor U4092 (N_4092,N_1523,N_1026);
nor U4093 (N_4093,N_1280,N_758);
or U4094 (N_4094,N_7,N_953);
or U4095 (N_4095,N_989,N_298);
xnor U4096 (N_4096,N_15,N_2481);
and U4097 (N_4097,N_2241,N_967);
xnor U4098 (N_4098,N_512,N_2390);
nor U4099 (N_4099,N_1782,N_1834);
or U4100 (N_4100,N_2405,N_278);
nand U4101 (N_4101,N_2137,N_1453);
and U4102 (N_4102,N_1378,N_1919);
nor U4103 (N_4103,N_1741,N_2396);
nand U4104 (N_4104,N_1203,N_2039);
and U4105 (N_4105,N_2455,N_2468);
nor U4106 (N_4106,N_932,N_2278);
nand U4107 (N_4107,N_298,N_2116);
nor U4108 (N_4108,N_2469,N_764);
nor U4109 (N_4109,N_1839,N_7);
and U4110 (N_4110,N_937,N_2000);
nand U4111 (N_4111,N_1841,N_706);
and U4112 (N_4112,N_1739,N_988);
and U4113 (N_4113,N_1039,N_826);
xor U4114 (N_4114,N_944,N_121);
or U4115 (N_4115,N_1889,N_743);
nand U4116 (N_4116,N_51,N_2446);
or U4117 (N_4117,N_1544,N_296);
xor U4118 (N_4118,N_1284,N_2100);
nor U4119 (N_4119,N_1543,N_1034);
nor U4120 (N_4120,N_535,N_153);
nor U4121 (N_4121,N_1967,N_2046);
or U4122 (N_4122,N_2496,N_1122);
nor U4123 (N_4123,N_37,N_130);
and U4124 (N_4124,N_1132,N_1596);
xor U4125 (N_4125,N_704,N_1236);
nand U4126 (N_4126,N_178,N_560);
or U4127 (N_4127,N_259,N_956);
or U4128 (N_4128,N_1318,N_2228);
and U4129 (N_4129,N_196,N_1564);
or U4130 (N_4130,N_7,N_1984);
or U4131 (N_4131,N_2110,N_2007);
and U4132 (N_4132,N_2385,N_90);
nand U4133 (N_4133,N_444,N_2144);
and U4134 (N_4134,N_806,N_989);
or U4135 (N_4135,N_1159,N_234);
nand U4136 (N_4136,N_730,N_407);
or U4137 (N_4137,N_2007,N_1046);
nand U4138 (N_4138,N_700,N_312);
nor U4139 (N_4139,N_841,N_453);
nand U4140 (N_4140,N_2196,N_983);
nor U4141 (N_4141,N_30,N_2094);
or U4142 (N_4142,N_80,N_262);
nand U4143 (N_4143,N_1070,N_1420);
nor U4144 (N_4144,N_2113,N_1881);
nand U4145 (N_4145,N_2496,N_428);
and U4146 (N_4146,N_2186,N_196);
nor U4147 (N_4147,N_1127,N_2018);
xor U4148 (N_4148,N_1613,N_1034);
or U4149 (N_4149,N_1995,N_1553);
nand U4150 (N_4150,N_1825,N_347);
or U4151 (N_4151,N_1701,N_1122);
nor U4152 (N_4152,N_2021,N_1601);
nand U4153 (N_4153,N_2173,N_2012);
and U4154 (N_4154,N_858,N_1790);
nand U4155 (N_4155,N_1694,N_2228);
or U4156 (N_4156,N_885,N_2050);
or U4157 (N_4157,N_643,N_943);
nand U4158 (N_4158,N_441,N_1358);
and U4159 (N_4159,N_1254,N_1829);
or U4160 (N_4160,N_1158,N_1641);
nand U4161 (N_4161,N_234,N_1244);
and U4162 (N_4162,N_2029,N_838);
and U4163 (N_4163,N_2010,N_2264);
nor U4164 (N_4164,N_1017,N_1459);
nand U4165 (N_4165,N_480,N_1193);
xnor U4166 (N_4166,N_1179,N_998);
nand U4167 (N_4167,N_1114,N_1895);
nor U4168 (N_4168,N_201,N_1165);
nor U4169 (N_4169,N_2042,N_2435);
nand U4170 (N_4170,N_934,N_607);
and U4171 (N_4171,N_559,N_1361);
nand U4172 (N_4172,N_167,N_1790);
and U4173 (N_4173,N_2195,N_2424);
or U4174 (N_4174,N_417,N_1806);
and U4175 (N_4175,N_904,N_2091);
nand U4176 (N_4176,N_2050,N_1038);
nand U4177 (N_4177,N_504,N_842);
nor U4178 (N_4178,N_1371,N_2127);
nand U4179 (N_4179,N_1438,N_50);
nor U4180 (N_4180,N_1545,N_1353);
nand U4181 (N_4181,N_2384,N_2307);
nand U4182 (N_4182,N_1168,N_786);
nor U4183 (N_4183,N_58,N_545);
or U4184 (N_4184,N_1715,N_2366);
nand U4185 (N_4185,N_2271,N_1510);
xnor U4186 (N_4186,N_1739,N_1266);
nor U4187 (N_4187,N_491,N_1392);
nand U4188 (N_4188,N_2316,N_2244);
or U4189 (N_4189,N_1301,N_2018);
or U4190 (N_4190,N_1077,N_1391);
nand U4191 (N_4191,N_1690,N_842);
nor U4192 (N_4192,N_2101,N_1001);
nand U4193 (N_4193,N_270,N_136);
nand U4194 (N_4194,N_1033,N_2429);
or U4195 (N_4195,N_1680,N_2114);
and U4196 (N_4196,N_1660,N_309);
or U4197 (N_4197,N_2296,N_2035);
nand U4198 (N_4198,N_2142,N_1208);
nand U4199 (N_4199,N_2183,N_483);
or U4200 (N_4200,N_1066,N_1839);
and U4201 (N_4201,N_2287,N_1638);
xor U4202 (N_4202,N_27,N_761);
and U4203 (N_4203,N_648,N_1341);
nor U4204 (N_4204,N_1433,N_417);
and U4205 (N_4205,N_1982,N_1613);
or U4206 (N_4206,N_1889,N_640);
and U4207 (N_4207,N_647,N_844);
and U4208 (N_4208,N_2323,N_1709);
nor U4209 (N_4209,N_2122,N_222);
nor U4210 (N_4210,N_842,N_1098);
and U4211 (N_4211,N_702,N_1860);
and U4212 (N_4212,N_2312,N_1399);
xnor U4213 (N_4213,N_2041,N_591);
nor U4214 (N_4214,N_1079,N_2429);
and U4215 (N_4215,N_2243,N_412);
nor U4216 (N_4216,N_758,N_2177);
nand U4217 (N_4217,N_2335,N_1365);
nor U4218 (N_4218,N_1699,N_1413);
nor U4219 (N_4219,N_1951,N_372);
and U4220 (N_4220,N_2317,N_1279);
nand U4221 (N_4221,N_2158,N_15);
or U4222 (N_4222,N_21,N_1039);
and U4223 (N_4223,N_156,N_678);
nand U4224 (N_4224,N_1750,N_899);
nor U4225 (N_4225,N_1460,N_1457);
and U4226 (N_4226,N_1030,N_1254);
xor U4227 (N_4227,N_749,N_1030);
nor U4228 (N_4228,N_326,N_2379);
or U4229 (N_4229,N_245,N_1013);
nor U4230 (N_4230,N_1311,N_1494);
xnor U4231 (N_4231,N_1521,N_1184);
and U4232 (N_4232,N_2076,N_2346);
nor U4233 (N_4233,N_1497,N_2119);
nor U4234 (N_4234,N_2210,N_61);
nand U4235 (N_4235,N_1549,N_1419);
and U4236 (N_4236,N_1909,N_1091);
and U4237 (N_4237,N_1150,N_724);
nor U4238 (N_4238,N_1577,N_2467);
or U4239 (N_4239,N_1318,N_566);
nor U4240 (N_4240,N_902,N_217);
or U4241 (N_4241,N_1689,N_416);
nand U4242 (N_4242,N_1900,N_1915);
and U4243 (N_4243,N_2321,N_1709);
or U4244 (N_4244,N_1105,N_450);
xor U4245 (N_4245,N_1985,N_1812);
or U4246 (N_4246,N_1001,N_2233);
or U4247 (N_4247,N_302,N_392);
xor U4248 (N_4248,N_2058,N_55);
or U4249 (N_4249,N_2132,N_2446);
and U4250 (N_4250,N_70,N_792);
and U4251 (N_4251,N_1352,N_496);
and U4252 (N_4252,N_1384,N_248);
nor U4253 (N_4253,N_1054,N_745);
nor U4254 (N_4254,N_1615,N_1168);
nand U4255 (N_4255,N_160,N_1723);
nor U4256 (N_4256,N_389,N_2458);
nand U4257 (N_4257,N_1904,N_2275);
or U4258 (N_4258,N_286,N_2492);
nor U4259 (N_4259,N_583,N_1754);
and U4260 (N_4260,N_1164,N_1107);
nand U4261 (N_4261,N_813,N_553);
and U4262 (N_4262,N_1095,N_1027);
nand U4263 (N_4263,N_1698,N_1534);
and U4264 (N_4264,N_1271,N_609);
nor U4265 (N_4265,N_826,N_1590);
nand U4266 (N_4266,N_148,N_2379);
nand U4267 (N_4267,N_587,N_1397);
or U4268 (N_4268,N_2487,N_1289);
or U4269 (N_4269,N_1052,N_2497);
or U4270 (N_4270,N_842,N_1770);
and U4271 (N_4271,N_522,N_1515);
nand U4272 (N_4272,N_1950,N_1184);
nand U4273 (N_4273,N_1432,N_238);
or U4274 (N_4274,N_1718,N_2242);
or U4275 (N_4275,N_1084,N_81);
and U4276 (N_4276,N_1603,N_2014);
nand U4277 (N_4277,N_2276,N_411);
nand U4278 (N_4278,N_1583,N_506);
and U4279 (N_4279,N_1062,N_2088);
and U4280 (N_4280,N_355,N_872);
nand U4281 (N_4281,N_1924,N_696);
nand U4282 (N_4282,N_1315,N_2048);
and U4283 (N_4283,N_590,N_2016);
nand U4284 (N_4284,N_464,N_1932);
nand U4285 (N_4285,N_46,N_1378);
xor U4286 (N_4286,N_81,N_994);
nand U4287 (N_4287,N_7,N_33);
nor U4288 (N_4288,N_619,N_2451);
nor U4289 (N_4289,N_1639,N_2483);
nand U4290 (N_4290,N_1361,N_1743);
nand U4291 (N_4291,N_1905,N_1603);
nand U4292 (N_4292,N_1904,N_1567);
nor U4293 (N_4293,N_395,N_1005);
nor U4294 (N_4294,N_48,N_1158);
and U4295 (N_4295,N_1297,N_859);
nor U4296 (N_4296,N_64,N_2090);
nor U4297 (N_4297,N_1910,N_196);
nor U4298 (N_4298,N_1589,N_522);
or U4299 (N_4299,N_31,N_999);
nand U4300 (N_4300,N_2441,N_867);
nand U4301 (N_4301,N_2252,N_2137);
and U4302 (N_4302,N_1830,N_1985);
nand U4303 (N_4303,N_2158,N_650);
nand U4304 (N_4304,N_1173,N_1189);
nand U4305 (N_4305,N_1307,N_537);
nor U4306 (N_4306,N_317,N_1886);
nor U4307 (N_4307,N_1767,N_301);
nor U4308 (N_4308,N_406,N_1784);
or U4309 (N_4309,N_766,N_760);
xor U4310 (N_4310,N_1476,N_63);
and U4311 (N_4311,N_2139,N_2342);
or U4312 (N_4312,N_142,N_767);
nand U4313 (N_4313,N_1363,N_96);
and U4314 (N_4314,N_2230,N_612);
nor U4315 (N_4315,N_668,N_1392);
and U4316 (N_4316,N_1352,N_680);
and U4317 (N_4317,N_157,N_2224);
nor U4318 (N_4318,N_990,N_1442);
and U4319 (N_4319,N_1655,N_1415);
nor U4320 (N_4320,N_81,N_1689);
nor U4321 (N_4321,N_1486,N_1316);
nor U4322 (N_4322,N_2259,N_1392);
and U4323 (N_4323,N_190,N_324);
and U4324 (N_4324,N_2083,N_373);
nand U4325 (N_4325,N_125,N_1491);
and U4326 (N_4326,N_1983,N_1381);
xnor U4327 (N_4327,N_940,N_1681);
and U4328 (N_4328,N_1855,N_1933);
or U4329 (N_4329,N_22,N_1941);
nand U4330 (N_4330,N_1151,N_425);
and U4331 (N_4331,N_1365,N_624);
or U4332 (N_4332,N_709,N_493);
nor U4333 (N_4333,N_1469,N_1505);
and U4334 (N_4334,N_2367,N_329);
and U4335 (N_4335,N_165,N_1557);
nand U4336 (N_4336,N_1785,N_590);
nand U4337 (N_4337,N_2031,N_484);
nand U4338 (N_4338,N_631,N_2042);
nand U4339 (N_4339,N_2271,N_229);
nor U4340 (N_4340,N_568,N_2052);
and U4341 (N_4341,N_630,N_27);
nor U4342 (N_4342,N_884,N_1599);
xnor U4343 (N_4343,N_128,N_179);
nand U4344 (N_4344,N_236,N_23);
nor U4345 (N_4345,N_2439,N_967);
nor U4346 (N_4346,N_2429,N_1777);
nor U4347 (N_4347,N_1309,N_1513);
and U4348 (N_4348,N_1531,N_2054);
nand U4349 (N_4349,N_1759,N_2154);
or U4350 (N_4350,N_1787,N_1335);
and U4351 (N_4351,N_120,N_824);
xnor U4352 (N_4352,N_2441,N_154);
or U4353 (N_4353,N_849,N_774);
and U4354 (N_4354,N_1676,N_358);
and U4355 (N_4355,N_1845,N_1238);
nor U4356 (N_4356,N_1653,N_2078);
and U4357 (N_4357,N_2260,N_2477);
and U4358 (N_4358,N_1919,N_2288);
and U4359 (N_4359,N_2317,N_809);
nand U4360 (N_4360,N_760,N_904);
nor U4361 (N_4361,N_1851,N_1017);
nor U4362 (N_4362,N_2259,N_2112);
and U4363 (N_4363,N_2260,N_670);
nor U4364 (N_4364,N_965,N_1195);
nor U4365 (N_4365,N_415,N_1882);
nand U4366 (N_4366,N_1200,N_984);
or U4367 (N_4367,N_87,N_965);
or U4368 (N_4368,N_1984,N_626);
nand U4369 (N_4369,N_160,N_1533);
or U4370 (N_4370,N_415,N_204);
nand U4371 (N_4371,N_1026,N_184);
nand U4372 (N_4372,N_640,N_357);
nor U4373 (N_4373,N_207,N_1599);
or U4374 (N_4374,N_354,N_2114);
and U4375 (N_4375,N_152,N_2264);
nor U4376 (N_4376,N_139,N_1309);
xnor U4377 (N_4377,N_1570,N_257);
or U4378 (N_4378,N_2432,N_1110);
nor U4379 (N_4379,N_1414,N_1038);
nand U4380 (N_4380,N_290,N_1265);
nand U4381 (N_4381,N_1789,N_773);
or U4382 (N_4382,N_996,N_953);
xnor U4383 (N_4383,N_182,N_1021);
xor U4384 (N_4384,N_759,N_890);
nand U4385 (N_4385,N_1640,N_2062);
and U4386 (N_4386,N_2353,N_368);
and U4387 (N_4387,N_2419,N_276);
xnor U4388 (N_4388,N_1285,N_1742);
xor U4389 (N_4389,N_1511,N_1772);
or U4390 (N_4390,N_2474,N_1111);
or U4391 (N_4391,N_2285,N_2295);
or U4392 (N_4392,N_835,N_165);
and U4393 (N_4393,N_288,N_109);
and U4394 (N_4394,N_1536,N_230);
nand U4395 (N_4395,N_1141,N_543);
or U4396 (N_4396,N_1927,N_1504);
xor U4397 (N_4397,N_1087,N_1429);
or U4398 (N_4398,N_277,N_2195);
nand U4399 (N_4399,N_832,N_1094);
and U4400 (N_4400,N_1693,N_1276);
nand U4401 (N_4401,N_378,N_1409);
and U4402 (N_4402,N_793,N_2297);
nand U4403 (N_4403,N_415,N_1437);
and U4404 (N_4404,N_1924,N_730);
xor U4405 (N_4405,N_433,N_2321);
nand U4406 (N_4406,N_1127,N_2307);
and U4407 (N_4407,N_484,N_465);
and U4408 (N_4408,N_1466,N_270);
or U4409 (N_4409,N_992,N_1477);
nand U4410 (N_4410,N_764,N_1245);
nand U4411 (N_4411,N_1871,N_1097);
and U4412 (N_4412,N_972,N_1862);
nand U4413 (N_4413,N_579,N_2061);
and U4414 (N_4414,N_1811,N_677);
and U4415 (N_4415,N_293,N_1503);
and U4416 (N_4416,N_1148,N_2097);
and U4417 (N_4417,N_2064,N_795);
nand U4418 (N_4418,N_328,N_1622);
and U4419 (N_4419,N_200,N_2041);
or U4420 (N_4420,N_779,N_2379);
nand U4421 (N_4421,N_2496,N_782);
nand U4422 (N_4422,N_304,N_303);
nor U4423 (N_4423,N_2458,N_1641);
xnor U4424 (N_4424,N_798,N_1196);
xnor U4425 (N_4425,N_1450,N_654);
xor U4426 (N_4426,N_659,N_2080);
nor U4427 (N_4427,N_584,N_1127);
and U4428 (N_4428,N_2375,N_1083);
and U4429 (N_4429,N_2185,N_1147);
xnor U4430 (N_4430,N_806,N_1282);
xnor U4431 (N_4431,N_639,N_1241);
nand U4432 (N_4432,N_2413,N_2304);
or U4433 (N_4433,N_438,N_561);
nor U4434 (N_4434,N_1306,N_1138);
and U4435 (N_4435,N_262,N_1399);
nand U4436 (N_4436,N_1661,N_1887);
nor U4437 (N_4437,N_727,N_2223);
and U4438 (N_4438,N_2424,N_454);
nor U4439 (N_4439,N_735,N_1366);
or U4440 (N_4440,N_439,N_1973);
or U4441 (N_4441,N_2093,N_2318);
nand U4442 (N_4442,N_1649,N_60);
xnor U4443 (N_4443,N_47,N_1853);
and U4444 (N_4444,N_152,N_740);
nand U4445 (N_4445,N_599,N_1618);
nor U4446 (N_4446,N_1627,N_1111);
nand U4447 (N_4447,N_1082,N_1188);
nand U4448 (N_4448,N_868,N_1753);
nand U4449 (N_4449,N_2256,N_1909);
xor U4450 (N_4450,N_2024,N_1143);
nand U4451 (N_4451,N_1789,N_1637);
or U4452 (N_4452,N_224,N_1443);
nor U4453 (N_4453,N_52,N_947);
or U4454 (N_4454,N_140,N_651);
xnor U4455 (N_4455,N_1896,N_936);
nand U4456 (N_4456,N_699,N_1555);
nor U4457 (N_4457,N_1774,N_542);
and U4458 (N_4458,N_819,N_446);
nor U4459 (N_4459,N_777,N_1683);
nand U4460 (N_4460,N_72,N_2066);
and U4461 (N_4461,N_423,N_560);
nor U4462 (N_4462,N_246,N_1447);
xor U4463 (N_4463,N_1077,N_933);
xor U4464 (N_4464,N_992,N_284);
nor U4465 (N_4465,N_1881,N_1697);
nand U4466 (N_4466,N_2429,N_1383);
xnor U4467 (N_4467,N_23,N_2275);
nand U4468 (N_4468,N_2378,N_892);
nand U4469 (N_4469,N_667,N_1734);
or U4470 (N_4470,N_2395,N_2331);
nand U4471 (N_4471,N_1190,N_942);
and U4472 (N_4472,N_1751,N_2111);
xnor U4473 (N_4473,N_19,N_1172);
nor U4474 (N_4474,N_2184,N_25);
or U4475 (N_4475,N_2271,N_1206);
or U4476 (N_4476,N_229,N_1874);
and U4477 (N_4477,N_1731,N_614);
and U4478 (N_4478,N_1540,N_751);
xor U4479 (N_4479,N_2228,N_1092);
nand U4480 (N_4480,N_1661,N_1956);
or U4481 (N_4481,N_237,N_2210);
nand U4482 (N_4482,N_1875,N_2452);
or U4483 (N_4483,N_2498,N_1955);
nand U4484 (N_4484,N_2235,N_1315);
nand U4485 (N_4485,N_613,N_1222);
or U4486 (N_4486,N_1126,N_1739);
xnor U4487 (N_4487,N_1230,N_2043);
or U4488 (N_4488,N_23,N_2235);
nand U4489 (N_4489,N_2338,N_829);
or U4490 (N_4490,N_2093,N_143);
nor U4491 (N_4491,N_429,N_1194);
nor U4492 (N_4492,N_2253,N_1446);
nor U4493 (N_4493,N_2398,N_1330);
nand U4494 (N_4494,N_2275,N_219);
nor U4495 (N_4495,N_2106,N_1150);
and U4496 (N_4496,N_578,N_7);
and U4497 (N_4497,N_92,N_1175);
nand U4498 (N_4498,N_1713,N_2302);
xor U4499 (N_4499,N_799,N_1742);
or U4500 (N_4500,N_701,N_1750);
nand U4501 (N_4501,N_1177,N_2163);
and U4502 (N_4502,N_98,N_1341);
nor U4503 (N_4503,N_1153,N_740);
nand U4504 (N_4504,N_1453,N_1622);
or U4505 (N_4505,N_105,N_1926);
or U4506 (N_4506,N_1289,N_2213);
or U4507 (N_4507,N_212,N_1780);
or U4508 (N_4508,N_2084,N_1649);
and U4509 (N_4509,N_389,N_250);
and U4510 (N_4510,N_1037,N_2300);
xnor U4511 (N_4511,N_2315,N_866);
xor U4512 (N_4512,N_34,N_279);
and U4513 (N_4513,N_986,N_397);
and U4514 (N_4514,N_123,N_2497);
nand U4515 (N_4515,N_1886,N_1051);
and U4516 (N_4516,N_646,N_244);
or U4517 (N_4517,N_306,N_1555);
or U4518 (N_4518,N_734,N_2292);
nand U4519 (N_4519,N_2332,N_402);
and U4520 (N_4520,N_630,N_107);
and U4521 (N_4521,N_1187,N_546);
nor U4522 (N_4522,N_257,N_745);
xnor U4523 (N_4523,N_1446,N_1338);
and U4524 (N_4524,N_655,N_638);
nor U4525 (N_4525,N_964,N_1266);
and U4526 (N_4526,N_1965,N_465);
nor U4527 (N_4527,N_265,N_1471);
or U4528 (N_4528,N_669,N_2014);
or U4529 (N_4529,N_18,N_2382);
and U4530 (N_4530,N_2150,N_1752);
nor U4531 (N_4531,N_2250,N_1389);
nor U4532 (N_4532,N_597,N_2274);
or U4533 (N_4533,N_997,N_596);
and U4534 (N_4534,N_1292,N_2465);
nor U4535 (N_4535,N_1588,N_2492);
nor U4536 (N_4536,N_1151,N_543);
xor U4537 (N_4537,N_1451,N_1885);
or U4538 (N_4538,N_308,N_914);
or U4539 (N_4539,N_2043,N_377);
or U4540 (N_4540,N_1923,N_1727);
nand U4541 (N_4541,N_1554,N_867);
or U4542 (N_4542,N_323,N_591);
nand U4543 (N_4543,N_279,N_806);
and U4544 (N_4544,N_1818,N_133);
and U4545 (N_4545,N_163,N_1565);
and U4546 (N_4546,N_662,N_2279);
and U4547 (N_4547,N_2061,N_483);
xor U4548 (N_4548,N_436,N_2417);
nor U4549 (N_4549,N_31,N_1317);
nor U4550 (N_4550,N_150,N_353);
nand U4551 (N_4551,N_566,N_236);
and U4552 (N_4552,N_1631,N_700);
or U4553 (N_4553,N_2052,N_243);
nand U4554 (N_4554,N_168,N_912);
and U4555 (N_4555,N_816,N_1658);
nor U4556 (N_4556,N_946,N_910);
or U4557 (N_4557,N_139,N_19);
xnor U4558 (N_4558,N_1339,N_1277);
or U4559 (N_4559,N_1010,N_1410);
or U4560 (N_4560,N_543,N_1753);
nor U4561 (N_4561,N_2036,N_778);
xor U4562 (N_4562,N_1903,N_1099);
nor U4563 (N_4563,N_802,N_54);
and U4564 (N_4564,N_2028,N_499);
nand U4565 (N_4565,N_1403,N_374);
nor U4566 (N_4566,N_1267,N_2465);
or U4567 (N_4567,N_869,N_2216);
nand U4568 (N_4568,N_2343,N_2281);
nor U4569 (N_4569,N_1090,N_2404);
nor U4570 (N_4570,N_2147,N_1271);
nor U4571 (N_4571,N_218,N_2474);
and U4572 (N_4572,N_1736,N_1528);
nand U4573 (N_4573,N_1639,N_474);
xor U4574 (N_4574,N_797,N_1438);
or U4575 (N_4575,N_2359,N_2163);
nand U4576 (N_4576,N_1690,N_783);
nor U4577 (N_4577,N_1868,N_2424);
and U4578 (N_4578,N_436,N_344);
nor U4579 (N_4579,N_1032,N_125);
or U4580 (N_4580,N_1774,N_83);
xor U4581 (N_4581,N_294,N_957);
and U4582 (N_4582,N_334,N_1535);
nand U4583 (N_4583,N_538,N_5);
nor U4584 (N_4584,N_896,N_2417);
or U4585 (N_4585,N_689,N_1898);
or U4586 (N_4586,N_1050,N_584);
nor U4587 (N_4587,N_1442,N_717);
nor U4588 (N_4588,N_2136,N_1432);
and U4589 (N_4589,N_1328,N_904);
nor U4590 (N_4590,N_2040,N_1701);
nand U4591 (N_4591,N_476,N_2157);
xnor U4592 (N_4592,N_1908,N_2212);
or U4593 (N_4593,N_957,N_2014);
xnor U4594 (N_4594,N_1987,N_87);
nand U4595 (N_4595,N_2375,N_1833);
xor U4596 (N_4596,N_1,N_182);
nor U4597 (N_4597,N_42,N_552);
or U4598 (N_4598,N_2267,N_1181);
xnor U4599 (N_4599,N_905,N_1149);
nor U4600 (N_4600,N_512,N_1838);
nor U4601 (N_4601,N_42,N_1729);
and U4602 (N_4602,N_560,N_185);
and U4603 (N_4603,N_1999,N_678);
and U4604 (N_4604,N_990,N_1416);
and U4605 (N_4605,N_1384,N_1919);
nor U4606 (N_4606,N_1650,N_2085);
nand U4607 (N_4607,N_1261,N_1925);
nand U4608 (N_4608,N_912,N_2305);
nor U4609 (N_4609,N_1414,N_761);
nand U4610 (N_4610,N_1423,N_1852);
nand U4611 (N_4611,N_1646,N_6);
nand U4612 (N_4612,N_1398,N_257);
nor U4613 (N_4613,N_439,N_1290);
nor U4614 (N_4614,N_473,N_1959);
nor U4615 (N_4615,N_2387,N_1368);
nand U4616 (N_4616,N_2239,N_2249);
nor U4617 (N_4617,N_1628,N_1415);
and U4618 (N_4618,N_1775,N_2198);
and U4619 (N_4619,N_1324,N_1512);
nand U4620 (N_4620,N_1092,N_1061);
nand U4621 (N_4621,N_1279,N_1927);
nand U4622 (N_4622,N_2230,N_1824);
nor U4623 (N_4623,N_2409,N_1531);
xor U4624 (N_4624,N_1691,N_469);
or U4625 (N_4625,N_1809,N_2420);
nand U4626 (N_4626,N_1554,N_901);
and U4627 (N_4627,N_623,N_162);
xor U4628 (N_4628,N_1775,N_996);
nand U4629 (N_4629,N_1707,N_2312);
nor U4630 (N_4630,N_1807,N_1735);
and U4631 (N_4631,N_2215,N_2092);
or U4632 (N_4632,N_815,N_1969);
xor U4633 (N_4633,N_581,N_188);
nor U4634 (N_4634,N_2227,N_2085);
and U4635 (N_4635,N_1263,N_2048);
or U4636 (N_4636,N_2480,N_2447);
or U4637 (N_4637,N_1730,N_92);
and U4638 (N_4638,N_1996,N_174);
nand U4639 (N_4639,N_116,N_1182);
and U4640 (N_4640,N_2079,N_1776);
or U4641 (N_4641,N_1685,N_2108);
nor U4642 (N_4642,N_320,N_2095);
nand U4643 (N_4643,N_1031,N_1707);
and U4644 (N_4644,N_1126,N_1084);
and U4645 (N_4645,N_178,N_1270);
or U4646 (N_4646,N_1617,N_1004);
nor U4647 (N_4647,N_1322,N_531);
and U4648 (N_4648,N_1404,N_779);
nand U4649 (N_4649,N_1288,N_1710);
and U4650 (N_4650,N_222,N_409);
nor U4651 (N_4651,N_1509,N_159);
and U4652 (N_4652,N_215,N_2059);
nor U4653 (N_4653,N_982,N_0);
or U4654 (N_4654,N_26,N_2174);
nor U4655 (N_4655,N_2258,N_1125);
or U4656 (N_4656,N_2021,N_1364);
nand U4657 (N_4657,N_693,N_2441);
and U4658 (N_4658,N_1641,N_1046);
nand U4659 (N_4659,N_2248,N_1001);
xnor U4660 (N_4660,N_733,N_2115);
or U4661 (N_4661,N_389,N_1978);
nor U4662 (N_4662,N_917,N_573);
nand U4663 (N_4663,N_1962,N_637);
and U4664 (N_4664,N_279,N_715);
and U4665 (N_4665,N_279,N_340);
xor U4666 (N_4666,N_836,N_490);
and U4667 (N_4667,N_1448,N_962);
nand U4668 (N_4668,N_2465,N_2449);
and U4669 (N_4669,N_2345,N_1348);
nand U4670 (N_4670,N_464,N_728);
and U4671 (N_4671,N_28,N_1132);
nor U4672 (N_4672,N_952,N_894);
nor U4673 (N_4673,N_2456,N_1696);
nand U4674 (N_4674,N_1368,N_1787);
or U4675 (N_4675,N_736,N_1185);
or U4676 (N_4676,N_1929,N_1165);
and U4677 (N_4677,N_409,N_2407);
or U4678 (N_4678,N_680,N_248);
xnor U4679 (N_4679,N_388,N_678);
nand U4680 (N_4680,N_1094,N_580);
nand U4681 (N_4681,N_1108,N_1647);
or U4682 (N_4682,N_162,N_1489);
nand U4683 (N_4683,N_2079,N_1067);
or U4684 (N_4684,N_400,N_846);
nand U4685 (N_4685,N_319,N_471);
and U4686 (N_4686,N_2010,N_1617);
and U4687 (N_4687,N_750,N_1750);
or U4688 (N_4688,N_1197,N_442);
nand U4689 (N_4689,N_148,N_1175);
nor U4690 (N_4690,N_25,N_717);
or U4691 (N_4691,N_2486,N_728);
nor U4692 (N_4692,N_1489,N_2363);
or U4693 (N_4693,N_1895,N_1373);
and U4694 (N_4694,N_2127,N_25);
or U4695 (N_4695,N_282,N_2314);
or U4696 (N_4696,N_793,N_92);
nand U4697 (N_4697,N_2200,N_1995);
xor U4698 (N_4698,N_1805,N_2464);
and U4699 (N_4699,N_1465,N_292);
and U4700 (N_4700,N_770,N_516);
and U4701 (N_4701,N_666,N_1408);
or U4702 (N_4702,N_590,N_325);
nor U4703 (N_4703,N_249,N_224);
xor U4704 (N_4704,N_2338,N_688);
and U4705 (N_4705,N_1749,N_2072);
and U4706 (N_4706,N_2390,N_464);
and U4707 (N_4707,N_851,N_121);
xor U4708 (N_4708,N_1517,N_182);
xor U4709 (N_4709,N_1331,N_25);
and U4710 (N_4710,N_481,N_747);
xor U4711 (N_4711,N_746,N_154);
xor U4712 (N_4712,N_2195,N_1630);
nor U4713 (N_4713,N_1868,N_894);
nor U4714 (N_4714,N_369,N_343);
nand U4715 (N_4715,N_2239,N_691);
and U4716 (N_4716,N_459,N_580);
or U4717 (N_4717,N_48,N_2410);
or U4718 (N_4718,N_2167,N_1464);
nor U4719 (N_4719,N_1744,N_1824);
nand U4720 (N_4720,N_954,N_935);
nand U4721 (N_4721,N_181,N_1989);
nand U4722 (N_4722,N_1640,N_2131);
and U4723 (N_4723,N_1054,N_2451);
xor U4724 (N_4724,N_460,N_610);
nor U4725 (N_4725,N_1327,N_2002);
xnor U4726 (N_4726,N_317,N_1072);
nand U4727 (N_4727,N_929,N_2261);
nand U4728 (N_4728,N_271,N_1368);
or U4729 (N_4729,N_842,N_753);
and U4730 (N_4730,N_215,N_497);
xnor U4731 (N_4731,N_1617,N_746);
nand U4732 (N_4732,N_32,N_1852);
or U4733 (N_4733,N_1719,N_6);
nand U4734 (N_4734,N_918,N_1133);
nand U4735 (N_4735,N_602,N_536);
or U4736 (N_4736,N_2413,N_2194);
and U4737 (N_4737,N_1167,N_683);
and U4738 (N_4738,N_297,N_1280);
and U4739 (N_4739,N_2497,N_1780);
nand U4740 (N_4740,N_2499,N_1912);
or U4741 (N_4741,N_401,N_837);
nor U4742 (N_4742,N_236,N_832);
or U4743 (N_4743,N_464,N_1628);
nor U4744 (N_4744,N_2066,N_840);
and U4745 (N_4745,N_2377,N_1772);
or U4746 (N_4746,N_2121,N_1005);
nand U4747 (N_4747,N_670,N_1643);
nand U4748 (N_4748,N_1424,N_2079);
xor U4749 (N_4749,N_1473,N_750);
and U4750 (N_4750,N_1757,N_1501);
nand U4751 (N_4751,N_1651,N_2281);
nor U4752 (N_4752,N_33,N_844);
and U4753 (N_4753,N_408,N_1743);
nor U4754 (N_4754,N_1054,N_160);
nand U4755 (N_4755,N_1126,N_1237);
nor U4756 (N_4756,N_873,N_1188);
and U4757 (N_4757,N_678,N_1989);
and U4758 (N_4758,N_136,N_1179);
or U4759 (N_4759,N_987,N_1420);
nor U4760 (N_4760,N_2094,N_1424);
or U4761 (N_4761,N_2105,N_176);
nor U4762 (N_4762,N_1369,N_1703);
or U4763 (N_4763,N_1156,N_1885);
nor U4764 (N_4764,N_1939,N_1075);
nor U4765 (N_4765,N_1998,N_635);
nand U4766 (N_4766,N_1217,N_1606);
nor U4767 (N_4767,N_1252,N_2263);
or U4768 (N_4768,N_1459,N_955);
nor U4769 (N_4769,N_2210,N_1828);
and U4770 (N_4770,N_2423,N_2269);
nand U4771 (N_4771,N_707,N_1315);
or U4772 (N_4772,N_378,N_478);
or U4773 (N_4773,N_2162,N_1216);
or U4774 (N_4774,N_2405,N_538);
and U4775 (N_4775,N_37,N_461);
and U4776 (N_4776,N_2424,N_2228);
or U4777 (N_4777,N_536,N_775);
or U4778 (N_4778,N_1621,N_1821);
and U4779 (N_4779,N_842,N_1407);
nor U4780 (N_4780,N_1646,N_732);
and U4781 (N_4781,N_1741,N_844);
nor U4782 (N_4782,N_1620,N_2152);
nand U4783 (N_4783,N_992,N_1897);
and U4784 (N_4784,N_635,N_452);
xnor U4785 (N_4785,N_490,N_586);
or U4786 (N_4786,N_936,N_1344);
nand U4787 (N_4787,N_210,N_956);
or U4788 (N_4788,N_1432,N_1991);
or U4789 (N_4789,N_768,N_2108);
nand U4790 (N_4790,N_1030,N_2071);
or U4791 (N_4791,N_2335,N_1866);
nor U4792 (N_4792,N_1341,N_1129);
nand U4793 (N_4793,N_237,N_431);
nor U4794 (N_4794,N_43,N_137);
or U4795 (N_4795,N_1859,N_294);
nand U4796 (N_4796,N_1468,N_460);
or U4797 (N_4797,N_1406,N_1586);
nor U4798 (N_4798,N_2031,N_2207);
nand U4799 (N_4799,N_70,N_2180);
nand U4800 (N_4800,N_1978,N_629);
and U4801 (N_4801,N_307,N_1505);
nor U4802 (N_4802,N_1151,N_257);
xnor U4803 (N_4803,N_1054,N_542);
or U4804 (N_4804,N_2050,N_132);
nor U4805 (N_4805,N_832,N_2448);
and U4806 (N_4806,N_616,N_146);
nand U4807 (N_4807,N_153,N_14);
nor U4808 (N_4808,N_287,N_1956);
nor U4809 (N_4809,N_1652,N_55);
or U4810 (N_4810,N_1918,N_1098);
nand U4811 (N_4811,N_1999,N_1399);
and U4812 (N_4812,N_286,N_2409);
or U4813 (N_4813,N_1961,N_182);
nor U4814 (N_4814,N_2084,N_567);
xnor U4815 (N_4815,N_839,N_1368);
nand U4816 (N_4816,N_1847,N_1893);
nand U4817 (N_4817,N_274,N_528);
nand U4818 (N_4818,N_646,N_2255);
nand U4819 (N_4819,N_1410,N_2103);
nor U4820 (N_4820,N_2307,N_2204);
nand U4821 (N_4821,N_912,N_2207);
xor U4822 (N_4822,N_1277,N_574);
or U4823 (N_4823,N_1693,N_234);
and U4824 (N_4824,N_1910,N_2053);
nor U4825 (N_4825,N_1823,N_873);
nand U4826 (N_4826,N_1816,N_753);
nor U4827 (N_4827,N_828,N_491);
nor U4828 (N_4828,N_564,N_370);
and U4829 (N_4829,N_2067,N_242);
or U4830 (N_4830,N_2465,N_2422);
nor U4831 (N_4831,N_308,N_1939);
nor U4832 (N_4832,N_2,N_1185);
nor U4833 (N_4833,N_1700,N_2372);
nand U4834 (N_4834,N_2198,N_262);
nand U4835 (N_4835,N_488,N_1478);
nor U4836 (N_4836,N_2493,N_516);
nand U4837 (N_4837,N_2125,N_2207);
nand U4838 (N_4838,N_451,N_669);
nor U4839 (N_4839,N_744,N_1855);
nor U4840 (N_4840,N_1632,N_1086);
or U4841 (N_4841,N_1523,N_2116);
and U4842 (N_4842,N_2240,N_66);
nand U4843 (N_4843,N_726,N_470);
nor U4844 (N_4844,N_1596,N_1968);
nor U4845 (N_4845,N_1835,N_494);
nor U4846 (N_4846,N_1782,N_993);
and U4847 (N_4847,N_1339,N_2229);
or U4848 (N_4848,N_610,N_1508);
nor U4849 (N_4849,N_1769,N_2382);
nand U4850 (N_4850,N_1156,N_1962);
or U4851 (N_4851,N_1051,N_2348);
nand U4852 (N_4852,N_1093,N_466);
xor U4853 (N_4853,N_910,N_653);
and U4854 (N_4854,N_2002,N_252);
nand U4855 (N_4855,N_1553,N_1105);
nand U4856 (N_4856,N_2431,N_1343);
and U4857 (N_4857,N_2300,N_776);
nand U4858 (N_4858,N_96,N_2438);
or U4859 (N_4859,N_2039,N_1374);
nand U4860 (N_4860,N_235,N_1823);
or U4861 (N_4861,N_2005,N_1377);
nor U4862 (N_4862,N_2194,N_450);
and U4863 (N_4863,N_36,N_2301);
and U4864 (N_4864,N_699,N_415);
nor U4865 (N_4865,N_362,N_1110);
nor U4866 (N_4866,N_1648,N_676);
and U4867 (N_4867,N_2489,N_1447);
and U4868 (N_4868,N_840,N_58);
nor U4869 (N_4869,N_1692,N_180);
or U4870 (N_4870,N_1663,N_1356);
and U4871 (N_4871,N_1386,N_670);
nor U4872 (N_4872,N_409,N_1364);
and U4873 (N_4873,N_2000,N_2289);
xor U4874 (N_4874,N_982,N_113);
or U4875 (N_4875,N_731,N_859);
or U4876 (N_4876,N_717,N_1406);
xnor U4877 (N_4877,N_301,N_1561);
nor U4878 (N_4878,N_1463,N_544);
xor U4879 (N_4879,N_2191,N_2074);
nand U4880 (N_4880,N_1718,N_537);
and U4881 (N_4881,N_552,N_1472);
or U4882 (N_4882,N_327,N_991);
or U4883 (N_4883,N_2118,N_701);
or U4884 (N_4884,N_137,N_1610);
nor U4885 (N_4885,N_2415,N_2428);
nand U4886 (N_4886,N_1325,N_2438);
and U4887 (N_4887,N_1720,N_1156);
or U4888 (N_4888,N_798,N_915);
nor U4889 (N_4889,N_659,N_2310);
nand U4890 (N_4890,N_1462,N_997);
nor U4891 (N_4891,N_1425,N_907);
or U4892 (N_4892,N_1395,N_1105);
nand U4893 (N_4893,N_1309,N_83);
and U4894 (N_4894,N_602,N_487);
or U4895 (N_4895,N_1968,N_2490);
or U4896 (N_4896,N_1550,N_1038);
or U4897 (N_4897,N_708,N_1059);
nor U4898 (N_4898,N_464,N_328);
or U4899 (N_4899,N_1967,N_658);
or U4900 (N_4900,N_426,N_1666);
nand U4901 (N_4901,N_951,N_1904);
or U4902 (N_4902,N_1820,N_549);
nor U4903 (N_4903,N_2084,N_1258);
and U4904 (N_4904,N_1305,N_344);
nand U4905 (N_4905,N_1956,N_975);
nand U4906 (N_4906,N_2323,N_1014);
or U4907 (N_4907,N_1151,N_518);
nand U4908 (N_4908,N_562,N_2122);
and U4909 (N_4909,N_123,N_716);
nor U4910 (N_4910,N_410,N_2370);
nand U4911 (N_4911,N_1711,N_2020);
or U4912 (N_4912,N_166,N_1647);
and U4913 (N_4913,N_1712,N_2202);
and U4914 (N_4914,N_2226,N_1455);
and U4915 (N_4915,N_743,N_2207);
and U4916 (N_4916,N_1927,N_566);
nand U4917 (N_4917,N_1567,N_2288);
or U4918 (N_4918,N_2196,N_109);
nor U4919 (N_4919,N_880,N_2455);
or U4920 (N_4920,N_112,N_981);
or U4921 (N_4921,N_455,N_209);
nor U4922 (N_4922,N_1590,N_1451);
nand U4923 (N_4923,N_1936,N_1194);
and U4924 (N_4924,N_2081,N_242);
or U4925 (N_4925,N_2183,N_792);
nor U4926 (N_4926,N_2135,N_1964);
or U4927 (N_4927,N_1538,N_70);
nor U4928 (N_4928,N_227,N_1611);
or U4929 (N_4929,N_2119,N_2488);
and U4930 (N_4930,N_773,N_1586);
or U4931 (N_4931,N_2483,N_1233);
nor U4932 (N_4932,N_2379,N_1034);
nor U4933 (N_4933,N_806,N_1490);
nor U4934 (N_4934,N_998,N_1345);
nand U4935 (N_4935,N_1502,N_1712);
nor U4936 (N_4936,N_112,N_777);
nand U4937 (N_4937,N_155,N_1465);
nand U4938 (N_4938,N_655,N_2296);
nor U4939 (N_4939,N_2317,N_1810);
and U4940 (N_4940,N_1171,N_236);
nor U4941 (N_4941,N_6,N_1959);
xnor U4942 (N_4942,N_980,N_1926);
nor U4943 (N_4943,N_1862,N_964);
xor U4944 (N_4944,N_1990,N_2254);
nor U4945 (N_4945,N_1007,N_1685);
nor U4946 (N_4946,N_2321,N_919);
and U4947 (N_4947,N_1031,N_1255);
and U4948 (N_4948,N_2170,N_1182);
or U4949 (N_4949,N_905,N_1522);
and U4950 (N_4950,N_1374,N_2450);
nand U4951 (N_4951,N_206,N_926);
nand U4952 (N_4952,N_212,N_1371);
nand U4953 (N_4953,N_1799,N_501);
xnor U4954 (N_4954,N_404,N_1739);
and U4955 (N_4955,N_2165,N_1282);
or U4956 (N_4956,N_303,N_1662);
nand U4957 (N_4957,N_1879,N_1833);
xor U4958 (N_4958,N_1414,N_1799);
or U4959 (N_4959,N_2362,N_116);
or U4960 (N_4960,N_1388,N_971);
or U4961 (N_4961,N_2378,N_926);
and U4962 (N_4962,N_2124,N_987);
nor U4963 (N_4963,N_835,N_323);
nand U4964 (N_4964,N_1910,N_1073);
or U4965 (N_4965,N_1122,N_1295);
xnor U4966 (N_4966,N_497,N_2216);
or U4967 (N_4967,N_1554,N_1975);
nand U4968 (N_4968,N_2373,N_149);
and U4969 (N_4969,N_13,N_1095);
nor U4970 (N_4970,N_1560,N_178);
and U4971 (N_4971,N_1144,N_339);
or U4972 (N_4972,N_896,N_2007);
and U4973 (N_4973,N_1707,N_1962);
nor U4974 (N_4974,N_2364,N_921);
nor U4975 (N_4975,N_340,N_2257);
nor U4976 (N_4976,N_358,N_2188);
and U4977 (N_4977,N_1072,N_1243);
and U4978 (N_4978,N_1999,N_305);
nand U4979 (N_4979,N_1144,N_1064);
nand U4980 (N_4980,N_321,N_1026);
xor U4981 (N_4981,N_145,N_99);
xnor U4982 (N_4982,N_915,N_664);
nand U4983 (N_4983,N_714,N_1244);
nor U4984 (N_4984,N_1006,N_1175);
and U4985 (N_4985,N_1704,N_1451);
xnor U4986 (N_4986,N_353,N_453);
or U4987 (N_4987,N_149,N_1691);
and U4988 (N_4988,N_2133,N_2318);
nor U4989 (N_4989,N_2203,N_265);
nor U4990 (N_4990,N_2032,N_1344);
nor U4991 (N_4991,N_2291,N_1539);
nor U4992 (N_4992,N_2276,N_538);
or U4993 (N_4993,N_513,N_1030);
nor U4994 (N_4994,N_837,N_2135);
nand U4995 (N_4995,N_1227,N_544);
nor U4996 (N_4996,N_1421,N_1136);
nor U4997 (N_4997,N_1443,N_929);
nor U4998 (N_4998,N_960,N_618);
nand U4999 (N_4999,N_2251,N_633);
nand U5000 (N_5000,N_4923,N_4584);
or U5001 (N_5001,N_4176,N_4055);
nor U5002 (N_5002,N_2903,N_2672);
xor U5003 (N_5003,N_4899,N_2612);
xor U5004 (N_5004,N_4685,N_3634);
and U5005 (N_5005,N_4776,N_2704);
nand U5006 (N_5006,N_4203,N_3237);
xnor U5007 (N_5007,N_3766,N_3945);
nor U5008 (N_5008,N_3244,N_4528);
nor U5009 (N_5009,N_4819,N_4332);
or U5010 (N_5010,N_4397,N_3386);
or U5011 (N_5011,N_4377,N_2926);
and U5012 (N_5012,N_3043,N_4078);
or U5013 (N_5013,N_2854,N_3291);
xnor U5014 (N_5014,N_4117,N_3466);
nor U5015 (N_5015,N_2951,N_4757);
nor U5016 (N_5016,N_4472,N_4961);
nor U5017 (N_5017,N_3120,N_4667);
xor U5018 (N_5018,N_4887,N_4309);
nand U5019 (N_5019,N_3926,N_2671);
or U5020 (N_5020,N_4022,N_2654);
and U5021 (N_5021,N_4791,N_2602);
nor U5022 (N_5022,N_3863,N_3310);
nand U5023 (N_5023,N_2681,N_4005);
or U5024 (N_5024,N_3369,N_2557);
and U5025 (N_5025,N_3658,N_4914);
or U5026 (N_5026,N_3697,N_2603);
nor U5027 (N_5027,N_3105,N_4829);
nor U5028 (N_5028,N_3363,N_4408);
xnor U5029 (N_5029,N_2942,N_3305);
nor U5030 (N_5030,N_3055,N_3839);
and U5031 (N_5031,N_2614,N_4904);
or U5032 (N_5032,N_2668,N_3206);
nand U5033 (N_5033,N_3478,N_4885);
or U5034 (N_5034,N_4211,N_4698);
nor U5035 (N_5035,N_3711,N_4768);
nor U5036 (N_5036,N_2694,N_2988);
nand U5037 (N_5037,N_4576,N_2724);
nor U5038 (N_5038,N_3250,N_3398);
nand U5039 (N_5039,N_3103,N_3391);
or U5040 (N_5040,N_3734,N_3112);
or U5041 (N_5041,N_4315,N_2791);
or U5042 (N_5042,N_4387,N_2962);
nor U5043 (N_5043,N_2792,N_2841);
nand U5044 (N_5044,N_2892,N_4288);
and U5045 (N_5045,N_4663,N_2787);
nand U5046 (N_5046,N_3018,N_2629);
xor U5047 (N_5047,N_4740,N_4901);
and U5048 (N_5048,N_4912,N_4617);
nand U5049 (N_5049,N_3725,N_3061);
or U5050 (N_5050,N_4338,N_3701);
nor U5051 (N_5051,N_2679,N_3608);
nor U5052 (N_5052,N_4809,N_3272);
and U5053 (N_5053,N_3065,N_2559);
xnor U5054 (N_5054,N_3251,N_3078);
nand U5055 (N_5055,N_4385,N_3284);
or U5056 (N_5056,N_4349,N_4144);
nand U5057 (N_5057,N_2598,N_3439);
or U5058 (N_5058,N_4084,N_3671);
or U5059 (N_5059,N_4872,N_2740);
or U5060 (N_5060,N_4652,N_4200);
or U5061 (N_5061,N_2961,N_3771);
nand U5062 (N_5062,N_3050,N_3510);
and U5063 (N_5063,N_4659,N_3920);
and U5064 (N_5064,N_4687,N_3320);
nor U5065 (N_5065,N_3017,N_4563);
nor U5066 (N_5066,N_4010,N_3451);
nor U5067 (N_5067,N_2851,N_4865);
xor U5068 (N_5068,N_2533,N_3474);
and U5069 (N_5069,N_3803,N_4034);
xor U5070 (N_5070,N_2505,N_2575);
or U5071 (N_5071,N_2738,N_3225);
or U5072 (N_5072,N_3855,N_3768);
nand U5073 (N_5073,N_3410,N_2610);
nand U5074 (N_5074,N_3279,N_4876);
nor U5075 (N_5075,N_3298,N_4559);
nand U5076 (N_5076,N_3495,N_3774);
nor U5077 (N_5077,N_3685,N_4074);
and U5078 (N_5078,N_2566,N_4087);
or U5079 (N_5079,N_3416,N_2577);
nand U5080 (N_5080,N_4875,N_4684);
and U5081 (N_5081,N_4372,N_2673);
or U5082 (N_5082,N_4143,N_4931);
nand U5083 (N_5083,N_3328,N_3249);
or U5084 (N_5084,N_4322,N_3853);
and U5085 (N_5085,N_3502,N_3807);
nand U5086 (N_5086,N_3976,N_3432);
or U5087 (N_5087,N_4379,N_4936);
or U5088 (N_5088,N_3149,N_4655);
and U5089 (N_5089,N_3889,N_3269);
and U5090 (N_5090,N_4162,N_2864);
or U5091 (N_5091,N_3083,N_4123);
nand U5092 (N_5092,N_3998,N_3544);
or U5093 (N_5093,N_2826,N_2924);
nor U5094 (N_5094,N_2959,N_3706);
xnor U5095 (N_5095,N_2811,N_2975);
nor U5096 (N_5096,N_3790,N_3592);
xor U5097 (N_5097,N_4880,N_3951);
nor U5098 (N_5098,N_4314,N_4145);
nor U5099 (N_5099,N_3151,N_3411);
or U5100 (N_5100,N_2808,N_2789);
and U5101 (N_5101,N_4506,N_4966);
and U5102 (N_5102,N_3224,N_2822);
and U5103 (N_5103,N_3735,N_4831);
xor U5104 (N_5104,N_3116,N_4075);
nand U5105 (N_5105,N_4641,N_3750);
nand U5106 (N_5106,N_3869,N_3554);
and U5107 (N_5107,N_3838,N_3381);
or U5108 (N_5108,N_4153,N_4769);
and U5109 (N_5109,N_4194,N_3773);
nand U5110 (N_5110,N_3045,N_4292);
or U5111 (N_5111,N_4008,N_3076);
xor U5112 (N_5112,N_4242,N_3261);
nor U5113 (N_5113,N_4304,N_2928);
nor U5114 (N_5114,N_2894,N_3593);
or U5115 (N_5115,N_3282,N_4575);
and U5116 (N_5116,N_3851,N_4424);
nand U5117 (N_5117,N_4588,N_3236);
nor U5118 (N_5118,N_4308,N_4004);
or U5119 (N_5119,N_3621,N_4488);
nor U5120 (N_5120,N_2540,N_2628);
nor U5121 (N_5121,N_2721,N_2729);
or U5122 (N_5122,N_2813,N_4491);
and U5123 (N_5123,N_4848,N_2706);
nor U5124 (N_5124,N_3082,N_3638);
nor U5125 (N_5125,N_4851,N_2678);
nand U5126 (N_5126,N_4639,N_4275);
nand U5127 (N_5127,N_3005,N_3543);
nor U5128 (N_5128,N_2630,N_3646);
and U5129 (N_5129,N_2597,N_2897);
and U5130 (N_5130,N_3182,N_4997);
nand U5131 (N_5131,N_3559,N_3896);
or U5132 (N_5132,N_3630,N_4501);
nand U5133 (N_5133,N_4594,N_2741);
or U5134 (N_5134,N_2595,N_4411);
or U5135 (N_5135,N_2590,N_3997);
xnor U5136 (N_5136,N_4085,N_3371);
xnor U5137 (N_5137,N_3340,N_3349);
and U5138 (N_5138,N_4765,N_2860);
nor U5139 (N_5139,N_3727,N_4170);
nor U5140 (N_5140,N_3744,N_4628);
or U5141 (N_5141,N_2796,N_4380);
and U5142 (N_5142,N_3358,N_3848);
or U5143 (N_5143,N_4573,N_4622);
and U5144 (N_5144,N_3641,N_3931);
and U5145 (N_5145,N_3792,N_4417);
and U5146 (N_5146,N_3166,N_4969);
nand U5147 (N_5147,N_4933,N_2762);
nor U5148 (N_5148,N_4522,N_3577);
or U5149 (N_5149,N_4076,N_2723);
xor U5150 (N_5150,N_3780,N_4700);
or U5151 (N_5151,N_3343,N_4215);
or U5152 (N_5152,N_2565,N_4538);
nand U5153 (N_5153,N_4447,N_2984);
and U5154 (N_5154,N_4774,N_4129);
or U5155 (N_5155,N_2967,N_4731);
nand U5156 (N_5156,N_4699,N_4516);
nand U5157 (N_5157,N_2698,N_3561);
and U5158 (N_5158,N_3874,N_3021);
nand U5159 (N_5159,N_3689,N_3739);
nand U5160 (N_5160,N_2948,N_3167);
or U5161 (N_5161,N_4883,N_3455);
nor U5162 (N_5162,N_4499,N_4994);
nand U5163 (N_5163,N_3527,N_4250);
xnor U5164 (N_5164,N_2755,N_4982);
xor U5165 (N_5165,N_4859,N_3642);
nor U5166 (N_5166,N_4764,N_3072);
nor U5167 (N_5167,N_4578,N_3453);
nand U5168 (N_5168,N_3223,N_3295);
or U5169 (N_5169,N_2583,N_4492);
and U5170 (N_5170,N_2814,N_4476);
xor U5171 (N_5171,N_2674,N_3423);
and U5172 (N_5172,N_3028,N_4228);
and U5173 (N_5173,N_4011,N_2564);
or U5174 (N_5174,N_4560,N_4240);
xnor U5175 (N_5175,N_2527,N_4734);
nor U5176 (N_5176,N_3899,N_4978);
or U5177 (N_5177,N_2558,N_3024);
and U5178 (N_5178,N_3587,N_2637);
and U5179 (N_5179,N_4513,N_2563);
and U5180 (N_5180,N_4817,N_3507);
nand U5181 (N_5181,N_3387,N_4452);
nor U5182 (N_5182,N_3908,N_3840);
nand U5183 (N_5183,N_4675,N_2799);
nor U5184 (N_5184,N_2749,N_4789);
or U5185 (N_5185,N_3098,N_4786);
xor U5186 (N_5186,N_4404,N_3214);
nand U5187 (N_5187,N_3456,N_3202);
or U5188 (N_5188,N_4673,N_4745);
nor U5189 (N_5189,N_2562,N_4175);
nand U5190 (N_5190,N_3562,N_3486);
or U5191 (N_5191,N_2874,N_4744);
nor U5192 (N_5192,N_3473,N_3514);
and U5193 (N_5193,N_4712,N_3347);
or U5194 (N_5194,N_2617,N_3201);
nand U5195 (N_5195,N_3881,N_3296);
and U5196 (N_5196,N_3664,N_4006);
or U5197 (N_5197,N_3183,N_4450);
nor U5198 (N_5198,N_3163,N_4291);
nor U5199 (N_5199,N_4135,N_4317);
nor U5200 (N_5200,N_3969,N_4775);
nor U5201 (N_5201,N_3170,N_4079);
nand U5202 (N_5202,N_3550,N_4448);
nand U5203 (N_5203,N_2682,N_3267);
nor U5204 (N_5204,N_3604,N_2775);
and U5205 (N_5205,N_2662,N_2898);
nor U5206 (N_5206,N_4344,N_4224);
and U5207 (N_5207,N_2646,N_4024);
nand U5208 (N_5208,N_4846,N_3511);
nor U5209 (N_5209,N_2594,N_4347);
or U5210 (N_5210,N_4165,N_4329);
xnor U5211 (N_5211,N_2700,N_3822);
and U5212 (N_5212,N_4193,N_3304);
nand U5213 (N_5213,N_4965,N_4196);
or U5214 (N_5214,N_2605,N_3912);
nor U5215 (N_5215,N_3069,N_4556);
or U5216 (N_5216,N_3796,N_2691);
nor U5217 (N_5217,N_3487,N_3463);
nor U5218 (N_5218,N_3030,N_3372);
nand U5219 (N_5219,N_4101,N_3203);
xor U5220 (N_5220,N_3230,N_4643);
or U5221 (N_5221,N_3538,N_4742);
and U5222 (N_5222,N_4626,N_3993);
and U5223 (N_5223,N_2536,N_2554);
nor U5224 (N_5224,N_2815,N_4727);
and U5225 (N_5225,N_2686,N_2716);
and U5226 (N_5226,N_2795,N_4231);
or U5227 (N_5227,N_3143,N_4572);
and U5228 (N_5228,N_2838,N_2767);
and U5229 (N_5229,N_2781,N_3057);
nand U5230 (N_5230,N_4577,N_3235);
nand U5231 (N_5231,N_2683,N_4278);
nand U5232 (N_5232,N_3709,N_4947);
and U5233 (N_5233,N_3533,N_2746);
or U5234 (N_5234,N_4987,N_3716);
nand U5235 (N_5235,N_4281,N_4157);
nand U5236 (N_5236,N_3353,N_4726);
or U5237 (N_5237,N_2555,N_2619);
or U5238 (N_5238,N_4721,N_4407);
and U5239 (N_5239,N_3779,N_3273);
or U5240 (N_5240,N_3003,N_4271);
and U5241 (N_5241,N_3414,N_3129);
or U5242 (N_5242,N_4654,N_4457);
and U5243 (N_5243,N_3088,N_2957);
and U5244 (N_5244,N_3321,N_4959);
nand U5245 (N_5245,N_4952,N_4739);
and U5246 (N_5246,N_3266,N_3265);
nor U5247 (N_5247,N_3217,N_2632);
nand U5248 (N_5248,N_3977,N_4390);
nand U5249 (N_5249,N_3285,N_4541);
and U5250 (N_5250,N_4330,N_4386);
nand U5251 (N_5251,N_4456,N_3753);
nor U5252 (N_5252,N_2886,N_4616);
nand U5253 (N_5253,N_4236,N_3929);
nor U5254 (N_5254,N_4102,N_2979);
or U5255 (N_5255,N_2997,N_4625);
or U5256 (N_5256,N_4077,N_4557);
xor U5257 (N_5257,N_4795,N_3812);
xnor U5258 (N_5258,N_3002,N_4061);
nor U5259 (N_5259,N_3615,N_3600);
and U5260 (N_5260,N_3910,N_4767);
and U5261 (N_5261,N_3344,N_3373);
xnor U5262 (N_5262,N_4855,N_3660);
nor U5263 (N_5263,N_2701,N_2506);
nor U5264 (N_5264,N_4527,N_2636);
xnor U5265 (N_5265,N_3429,N_4903);
nor U5266 (N_5266,N_3946,N_4830);
or U5267 (N_5267,N_4723,N_3520);
and U5268 (N_5268,N_3728,N_3232);
xor U5269 (N_5269,N_2908,N_3240);
nor U5270 (N_5270,N_3806,N_4126);
nor U5271 (N_5271,N_3588,N_2965);
nor U5272 (N_5272,N_4574,N_2976);
nor U5273 (N_5273,N_4777,N_3902);
nand U5274 (N_5274,N_3553,N_4551);
or U5275 (N_5275,N_4105,N_3177);
nand U5276 (N_5276,N_4879,N_2776);
xor U5277 (N_5277,N_4790,N_4426);
nor U5278 (N_5278,N_2524,N_3488);
or U5279 (N_5279,N_4239,N_3677);
or U5280 (N_5280,N_4627,N_3556);
nand U5281 (N_5281,N_3521,N_3365);
nand U5282 (N_5282,N_4651,N_4001);
or U5283 (N_5283,N_4542,N_3718);
and U5284 (N_5284,N_2664,N_3092);
nand U5285 (N_5285,N_4653,N_2635);
nor U5286 (N_5286,N_3074,N_4930);
and U5287 (N_5287,N_4052,N_3607);
and U5288 (N_5288,N_2880,N_4218);
xnor U5289 (N_5289,N_4805,N_2818);
or U5290 (N_5290,N_3610,N_2801);
nor U5291 (N_5291,N_4993,N_2896);
nand U5292 (N_5292,N_3574,N_3791);
or U5293 (N_5293,N_2757,N_4898);
nand U5294 (N_5294,N_4313,N_3653);
nand U5295 (N_5295,N_3179,N_4631);
xor U5296 (N_5296,N_3300,N_3268);
nor U5297 (N_5297,N_4439,N_4784);
and U5298 (N_5298,N_4319,N_3764);
or U5299 (N_5299,N_3877,N_4477);
or U5300 (N_5300,N_4695,N_2991);
or U5301 (N_5301,N_2649,N_4917);
or U5302 (N_5302,N_3211,N_3695);
nor U5303 (N_5303,N_4125,N_4216);
or U5304 (N_5304,N_4119,N_4350);
nor U5305 (N_5305,N_3162,N_3324);
nand U5306 (N_5306,N_3811,N_2613);
and U5307 (N_5307,N_2744,N_3060);
nand U5308 (N_5308,N_3142,N_3860);
nor U5309 (N_5309,N_3786,N_2687);
xor U5310 (N_5310,N_4249,N_4039);
or U5311 (N_5311,N_3091,N_3854);
or U5312 (N_5312,N_2836,N_4414);
nand U5313 (N_5313,N_3539,N_4722);
nor U5314 (N_5314,N_3271,N_3081);
nand U5315 (N_5315,N_2621,N_3430);
nor U5316 (N_5316,N_4284,N_3159);
or U5317 (N_5317,N_2653,N_4049);
and U5318 (N_5318,N_3672,N_4031);
nor U5319 (N_5319,N_4610,N_4428);
or U5320 (N_5320,N_3490,N_4591);
and U5321 (N_5321,N_4642,N_4285);
xnor U5322 (N_5322,N_3454,N_3040);
and U5323 (N_5323,N_4012,N_3576);
or U5324 (N_5324,N_4261,N_3821);
or U5325 (N_5325,N_2925,N_2888);
nand U5326 (N_5326,N_4054,N_4946);
or U5327 (N_5327,N_2805,N_2656);
nand U5328 (N_5328,N_4847,N_4369);
xor U5329 (N_5329,N_2504,N_4694);
nand U5330 (N_5330,N_4030,N_2515);
nand U5331 (N_5331,N_3808,N_3276);
nor U5332 (N_5332,N_4394,N_3342);
and U5333 (N_5333,N_3663,N_3622);
and U5334 (N_5334,N_3552,N_3086);
nand U5335 (N_5335,N_4098,N_4918);
or U5336 (N_5336,N_3684,N_4844);
nand U5337 (N_5337,N_4204,N_4048);
nor U5338 (N_5338,N_4913,N_4155);
and U5339 (N_5339,N_3668,N_4188);
nand U5340 (N_5340,N_4137,N_4780);
nand U5341 (N_5341,N_4097,N_3900);
nand U5342 (N_5342,N_3799,N_3311);
and U5343 (N_5343,N_2537,N_4420);
and U5344 (N_5344,N_3783,N_3836);
and U5345 (N_5345,N_3048,N_2503);
and U5346 (N_5346,N_2964,N_4517);
or U5347 (N_5347,N_3168,N_2665);
nand U5348 (N_5348,N_3096,N_3243);
or U5349 (N_5349,N_4127,N_2710);
nand U5350 (N_5350,N_3299,N_4352);
and U5351 (N_5351,N_3443,N_2955);
nor U5352 (N_5352,N_4614,N_2618);
or U5353 (N_5353,N_4986,N_3654);
nor U5354 (N_5354,N_4132,N_3425);
xor U5355 (N_5355,N_4172,N_4571);
nand U5356 (N_5356,N_4185,N_4658);
nand U5357 (N_5357,N_3568,N_2660);
or U5358 (N_5358,N_2571,N_2622);
and U5359 (N_5359,N_3318,N_4804);
and U5360 (N_5360,N_2802,N_3011);
nor U5361 (N_5361,N_4497,N_3397);
or U5362 (N_5362,N_3713,N_4362);
nand U5363 (N_5363,N_2733,N_4106);
and U5364 (N_5364,N_2817,N_3468);
nor U5365 (N_5365,N_4134,N_3359);
and U5366 (N_5366,N_4709,N_2507);
nor U5367 (N_5367,N_4733,N_3756);
nand U5368 (N_5368,N_4148,N_2850);
and U5369 (N_5369,N_4378,N_4587);
xnor U5370 (N_5370,N_4779,N_3705);
nor U5371 (N_5371,N_3944,N_4827);
nand U5372 (N_5372,N_3555,N_3708);
xnor U5373 (N_5373,N_3348,N_4264);
nor U5374 (N_5374,N_3312,N_4714);
nor U5375 (N_5375,N_4824,N_3107);
xnor U5376 (N_5376,N_3191,N_3814);
nor U5377 (N_5377,N_2675,N_2844);
nand U5378 (N_5378,N_3625,N_3837);
or U5379 (N_5379,N_2780,N_4896);
nand U5380 (N_5380,N_2692,N_2752);
and U5381 (N_5381,N_2845,N_3274);
or U5382 (N_5382,N_4432,N_3584);
nor U5383 (N_5383,N_2901,N_4507);
nand U5384 (N_5384,N_2727,N_4579);
xor U5385 (N_5385,N_4995,N_3326);
and U5386 (N_5386,N_4593,N_4253);
xor U5387 (N_5387,N_4130,N_3341);
and U5388 (N_5388,N_3479,N_4437);
or U5389 (N_5389,N_2713,N_3401);
and U5390 (N_5390,N_2914,N_3139);
nor U5391 (N_5391,N_4608,N_3742);
and U5392 (N_5392,N_3313,N_2807);
xnor U5393 (N_5393,N_2819,N_3136);
and U5394 (N_5394,N_3064,N_3886);
and U5395 (N_5395,N_4050,N_3333);
nand U5396 (N_5396,N_4632,N_4038);
nand U5397 (N_5397,N_3563,N_4611);
and U5398 (N_5398,N_4058,N_3797);
or U5399 (N_5399,N_3160,N_3213);
or U5400 (N_5400,N_2772,N_4853);
xnor U5401 (N_5401,N_2648,N_3482);
xor U5402 (N_5402,N_4979,N_3933);
nor U5403 (N_5403,N_2846,N_3334);
nand U5404 (N_5404,N_4635,N_4171);
nor U5405 (N_5405,N_2545,N_3582);
or U5406 (N_5406,N_3194,N_3135);
xnor U5407 (N_5407,N_4567,N_2876);
nand U5408 (N_5408,N_3415,N_4713);
xor U5409 (N_5409,N_3392,N_2812);
nor U5410 (N_5410,N_3963,N_3483);
or U5411 (N_5411,N_4729,N_4139);
nand U5412 (N_5412,N_2939,N_3594);
or U5413 (N_5413,N_3717,N_4435);
or U5414 (N_5414,N_2581,N_3212);
or U5415 (N_5415,N_3459,N_3111);
nor U5416 (N_5416,N_3763,N_4463);
xor U5417 (N_5417,N_2861,N_4656);
nor U5418 (N_5418,N_3572,N_3651);
nand U5419 (N_5419,N_2765,N_2834);
and U5420 (N_5420,N_4920,N_3970);
or U5421 (N_5421,N_3820,N_3809);
and U5422 (N_5422,N_4998,N_3073);
nor U5423 (N_5423,N_4686,N_4014);
and U5424 (N_5424,N_4163,N_4154);
nor U5425 (N_5425,N_3955,N_3173);
and U5426 (N_5426,N_2661,N_2714);
nand U5427 (N_5427,N_4895,N_4690);
and U5428 (N_5428,N_3053,N_3119);
xor U5429 (N_5429,N_3571,N_4521);
nor U5430 (N_5430,N_4479,N_2719);
nand U5431 (N_5431,N_4187,N_4564);
xnor U5432 (N_5432,N_3719,N_4482);
nand U5433 (N_5433,N_4182,N_4149);
xor U5434 (N_5434,N_2731,N_3505);
and U5435 (N_5435,N_4464,N_2549);
and U5436 (N_5436,N_3252,N_3759);
and U5437 (N_5437,N_2690,N_3408);
nand U5438 (N_5438,N_3937,N_2702);
or U5439 (N_5439,N_2945,N_2883);
nand U5440 (N_5440,N_2875,N_4648);
nand U5441 (N_5441,N_3657,N_3681);
and U5442 (N_5442,N_4983,N_3503);
nor U5443 (N_5443,N_2856,N_4927);
nor U5444 (N_5444,N_3376,N_2981);
and U5445 (N_5445,N_3636,N_3523);
nand U5446 (N_5446,N_3823,N_3567);
nor U5447 (N_5447,N_2972,N_4837);
nand U5448 (N_5448,N_4724,N_4179);
nand U5449 (N_5449,N_4916,N_3974);
and U5450 (N_5450,N_4807,N_3962);
nand U5451 (N_5451,N_2745,N_3442);
nor U5452 (N_5452,N_3176,N_4743);
and U5453 (N_5453,N_3856,N_2935);
nor U5454 (N_5454,N_2950,N_3674);
or U5455 (N_5455,N_2969,N_3366);
nand U5456 (N_5456,N_3772,N_3800);
xor U5457 (N_5457,N_4433,N_2532);
or U5458 (N_5458,N_3145,N_2909);
or U5459 (N_5459,N_2919,N_4856);
xor U5460 (N_5460,N_4558,N_4178);
and U5461 (N_5461,N_4295,N_2978);
xnor U5462 (N_5462,N_3012,N_3936);
xnor U5463 (N_5463,N_3165,N_4060);
nor U5464 (N_5464,N_4888,N_2918);
nand U5465 (N_5465,N_4028,N_4410);
xor U5466 (N_5466,N_4832,N_4247);
xnor U5467 (N_5467,N_4099,N_3435);
nand U5468 (N_5468,N_4057,N_4544);
nor U5469 (N_5469,N_3934,N_4376);
nand U5470 (N_5470,N_3242,N_4519);
nor U5471 (N_5471,N_3732,N_2634);
or U5472 (N_5472,N_2624,N_4301);
nand U5473 (N_5473,N_4666,N_4045);
nor U5474 (N_5474,N_4209,N_4198);
nor U5475 (N_5475,N_4533,N_4802);
or U5476 (N_5476,N_3745,N_2580);
nor U5477 (N_5477,N_2947,N_2728);
nand U5478 (N_5478,N_4881,N_4481);
or U5479 (N_5479,N_3010,N_2879);
and U5480 (N_5480,N_2989,N_4581);
and U5481 (N_5481,N_3013,N_4598);
or U5482 (N_5482,N_3286,N_4681);
and U5483 (N_5483,N_2786,N_2720);
nor U5484 (N_5484,N_2971,N_4677);
and U5485 (N_5485,N_4877,N_3850);
nor U5486 (N_5486,N_4468,N_2857);
xnor U5487 (N_5487,N_2677,N_4202);
nor U5488 (N_5488,N_4088,N_3616);
nor U5489 (N_5489,N_2858,N_4884);
nor U5490 (N_5490,N_3292,N_2530);
and U5491 (N_5491,N_4766,N_2759);
nor U5492 (N_5492,N_4756,N_3586);
nand U5493 (N_5493,N_4116,N_2758);
nand U5494 (N_5494,N_4429,N_4190);
xor U5495 (N_5495,N_2705,N_4040);
or U5496 (N_5496,N_4942,N_4850);
or U5497 (N_5497,N_4366,N_3322);
nand U5498 (N_5498,N_3501,N_3364);
and U5499 (N_5499,N_4430,N_3761);
nor U5500 (N_5500,N_4976,N_3661);
xor U5501 (N_5501,N_4266,N_4273);
or U5502 (N_5502,N_3885,N_3597);
nand U5503 (N_5503,N_3475,N_4719);
or U5504 (N_5504,N_4928,N_4825);
and U5505 (N_5505,N_3404,N_3508);
xnor U5506 (N_5506,N_4661,N_4421);
nor U5507 (N_5507,N_4523,N_2693);
nand U5508 (N_5508,N_4630,N_3470);
nand U5509 (N_5509,N_3990,N_4715);
xor U5510 (N_5510,N_3733,N_3513);
xor U5511 (N_5511,N_4967,N_4431);
and U5512 (N_5512,N_3181,N_3583);
nor U5513 (N_5513,N_4181,N_4728);
and U5514 (N_5514,N_3618,N_4445);
nor U5515 (N_5515,N_4502,N_4364);
nor U5516 (N_5516,N_4570,N_4036);
or U5517 (N_5517,N_3500,N_2611);
xor U5518 (N_5518,N_3027,N_3380);
nand U5519 (N_5519,N_4787,N_3694);
or U5520 (N_5520,N_3825,N_2788);
and U5521 (N_5521,N_3743,N_4670);
or U5522 (N_5522,N_4554,N_3585);
nand U5523 (N_5523,N_4037,N_4401);
or U5524 (N_5524,N_3765,N_3884);
and U5525 (N_5525,N_4939,N_4867);
and U5526 (N_5526,N_4945,N_3897);
and U5527 (N_5527,N_3703,N_3180);
nor U5528 (N_5528,N_3611,N_4835);
nor U5529 (N_5529,N_4371,N_3019);
nand U5530 (N_5530,N_3288,N_2585);
and U5531 (N_5531,N_3873,N_3147);
nor U5532 (N_5532,N_4358,N_2553);
nand U5533 (N_5533,N_4298,N_3542);
xor U5534 (N_5534,N_3154,N_3015);
or U5535 (N_5535,N_3384,N_3991);
and U5536 (N_5536,N_2800,N_3026);
nand U5537 (N_5537,N_3782,N_3323);
nand U5538 (N_5538,N_4660,N_4629);
and U5539 (N_5539,N_3314,N_3988);
xnor U5540 (N_5540,N_4638,N_2751);
or U5541 (N_5541,N_2525,N_2821);
xor U5542 (N_5542,N_3484,N_3126);
nor U5543 (N_5543,N_2993,N_3516);
or U5544 (N_5544,N_3370,N_3606);
or U5545 (N_5545,N_3834,N_4033);
xor U5546 (N_5546,N_4064,N_4138);
or U5547 (N_5547,N_4669,N_4268);
and U5548 (N_5548,N_3109,N_3751);
nor U5549 (N_5549,N_4612,N_2785);
nor U5550 (N_5550,N_4836,N_2626);
nor U5551 (N_5551,N_3345,N_3099);
and U5552 (N_5552,N_4356,N_4640);
and U5553 (N_5553,N_4514,N_3731);
nor U5554 (N_5554,N_3198,N_3054);
nor U5555 (N_5555,N_3009,N_4886);
nor U5556 (N_5556,N_2514,N_3256);
xor U5557 (N_5557,N_2608,N_3631);
nor U5558 (N_5558,N_3972,N_4255);
nand U5559 (N_5559,N_4158,N_4299);
nor U5560 (N_5560,N_4806,N_4046);
or U5561 (N_5561,N_2638,N_4173);
or U5562 (N_5562,N_2520,N_4500);
or U5563 (N_5563,N_3648,N_4672);
nand U5564 (N_5564,N_3623,N_4282);
xnor U5565 (N_5565,N_3210,N_3127);
nand U5566 (N_5566,N_2828,N_2916);
nor U5567 (N_5567,N_4526,N_4906);
nor U5568 (N_5568,N_2519,N_3595);
and U5569 (N_5569,N_2803,N_4941);
and U5570 (N_5570,N_3499,N_4725);
nor U5571 (N_5571,N_4136,N_4749);
nand U5572 (N_5572,N_3234,N_3827);
nand U5573 (N_5573,N_3164,N_3958);
or U5574 (N_5574,N_2512,N_2528);
nor U5575 (N_5575,N_3535,N_4343);
and U5576 (N_5576,N_4618,N_3652);
and U5577 (N_5577,N_3208,N_3248);
nand U5578 (N_5578,N_4915,N_4549);
nand U5579 (N_5579,N_4702,N_2849);
and U5580 (N_5580,N_3833,N_4258);
nand U5581 (N_5581,N_3316,N_4217);
xnor U5582 (N_5582,N_4161,N_2542);
xor U5583 (N_5583,N_3257,N_3767);
nor U5584 (N_5584,N_4552,N_4662);
and U5585 (N_5585,N_3609,N_2770);
or U5586 (N_5586,N_4160,N_2666);
nand U5587 (N_5587,N_4484,N_3506);
or U5588 (N_5588,N_4341,N_3828);
nor U5589 (N_5589,N_3222,N_3729);
nand U5590 (N_5590,N_4246,N_4826);
and U5591 (N_5591,N_4537,N_3575);
xor U5592 (N_5592,N_4813,N_3412);
xor U5593 (N_5593,N_4934,N_3428);
or U5594 (N_5594,N_4736,N_3868);
nand U5595 (N_5595,N_4580,N_4370);
nor U5596 (N_5596,N_4512,N_4985);
nand U5597 (N_5597,N_3356,N_4168);
nor U5598 (N_5598,N_3117,N_3346);
nand U5599 (N_5599,N_4707,N_4373);
or U5600 (N_5600,N_4260,N_3847);
and U5601 (N_5601,N_4693,N_4355);
nor U5602 (N_5602,N_4243,N_3400);
and U5603 (N_5603,N_3522,N_4335);
nor U5604 (N_5604,N_3068,N_2631);
and U5605 (N_5605,N_2680,N_3038);
and U5606 (N_5606,N_2640,N_4297);
nand U5607 (N_5607,N_4383,N_3130);
or U5608 (N_5608,N_3667,N_3132);
or U5609 (N_5609,N_3605,N_3862);
nand U5610 (N_5610,N_3351,N_2607);
xnor U5611 (N_5611,N_2806,N_3650);
or U5612 (N_5612,N_3540,N_4839);
xor U5613 (N_5613,N_2726,N_4925);
nand U5614 (N_5614,N_3699,N_3205);
nor U5615 (N_5615,N_3368,N_4027);
or U5616 (N_5616,N_3984,N_3941);
xnor U5617 (N_5617,N_2778,N_4657);
or U5618 (N_5618,N_4409,N_4703);
and U5619 (N_5619,N_3262,N_4307);
nor U5620 (N_5620,N_3953,N_3079);
and U5621 (N_5621,N_3961,N_2754);
or U5622 (N_5622,N_3949,N_2823);
or U5623 (N_5623,N_4316,N_3156);
nor U5624 (N_5624,N_4763,N_3871);
or U5625 (N_5625,N_4490,N_2932);
or U5626 (N_5626,N_4938,N_4873);
xnor U5627 (N_5627,N_2970,N_4760);
nand U5628 (N_5628,N_3619,N_4440);
nand U5629 (N_5629,N_3283,N_3327);
nand U5630 (N_5630,N_3805,N_3148);
and U5631 (N_5631,N_2768,N_3188);
nor U5632 (N_5632,N_2543,N_3966);
and U5633 (N_5633,N_2810,N_3128);
or U5634 (N_5634,N_4086,N_4320);
nand U5635 (N_5635,N_3329,N_4682);
or U5636 (N_5636,N_4056,N_4991);
xor U5637 (N_5637,N_4140,N_2589);
nor U5638 (N_5638,N_2987,N_4107);
nand U5639 (N_5639,N_3254,N_2995);
or U5640 (N_5640,N_3158,N_3125);
nand U5641 (N_5641,N_3246,N_3987);
or U5642 (N_5642,N_2912,N_2866);
and U5643 (N_5643,N_3730,N_3378);
nor U5644 (N_5644,N_3921,N_2921);
or U5645 (N_5645,N_3355,N_4592);
nor U5646 (N_5646,N_3231,N_3867);
or U5647 (N_5647,N_4494,N_3085);
nand U5648 (N_5648,N_3193,N_3883);
and U5649 (N_5649,N_3865,N_2839);
nand U5650 (N_5650,N_2958,N_3888);
and U5651 (N_5651,N_2560,N_3157);
and U5652 (N_5652,N_2940,N_2885);
xor U5653 (N_5653,N_2592,N_4794);
and U5654 (N_5654,N_3419,N_4676);
xor U5655 (N_5655,N_4645,N_4167);
nand U5656 (N_5656,N_3121,N_4555);
or U5657 (N_5657,N_4483,N_2552);
and U5658 (N_5658,N_4759,N_4065);
or U5659 (N_5659,N_4585,N_3440);
xnor U5660 (N_5660,N_4305,N_3992);
and U5661 (N_5661,N_2963,N_4334);
and U5662 (N_5662,N_4094,N_4436);
or U5663 (N_5663,N_2996,N_4461);
and U5664 (N_5664,N_3448,N_3629);
nor U5665 (N_5665,N_3080,N_3995);
nand U5666 (N_5666,N_4232,N_2994);
and U5667 (N_5667,N_4346,N_2907);
nor U5668 (N_5668,N_4720,N_4838);
nand U5669 (N_5669,N_3335,N_3260);
or U5670 (N_5670,N_2761,N_3377);
nor U5671 (N_5671,N_4423,N_2582);
and U5672 (N_5672,N_4459,N_4073);
nor U5673 (N_5673,N_3633,N_3656);
or U5674 (N_5674,N_3557,N_2625);
and U5675 (N_5675,N_2663,N_3978);
nand U5676 (N_5676,N_4324,N_3841);
nand U5677 (N_5677,N_3438,N_4705);
and U5678 (N_5678,N_3049,N_3207);
or U5679 (N_5679,N_2734,N_3673);
or U5680 (N_5680,N_3996,N_2865);
nand U5681 (N_5681,N_3187,N_4546);
and U5682 (N_5682,N_3239,N_3748);
or U5683 (N_5683,N_3287,N_4751);
and U5684 (N_5684,N_3784,N_2534);
or U5685 (N_5685,N_3545,N_4841);
nand U5686 (N_5686,N_3645,N_3426);
and U5687 (N_5687,N_2824,N_3515);
and U5688 (N_5688,N_3547,N_4843);
nand U5689 (N_5689,N_3123,N_2938);
or U5690 (N_5690,N_4926,N_2627);
or U5691 (N_5691,N_4023,N_3626);
or U5692 (N_5692,N_4957,N_4988);
nand U5693 (N_5693,N_4539,N_2531);
nor U5694 (N_5694,N_4002,N_2910);
xor U5695 (N_5695,N_4783,N_3035);
or U5696 (N_5696,N_2853,N_4532);
nand U5697 (N_5697,N_2526,N_3564);
and U5698 (N_5698,N_3935,N_3357);
nor U5699 (N_5699,N_4327,N_4475);
xnor U5700 (N_5700,N_4808,N_3361);
nand U5701 (N_5701,N_4637,N_4274);
nor U5702 (N_5702,N_3022,N_3033);
nand U5703 (N_5703,N_3031,N_3532);
xor U5704 (N_5704,N_3472,N_4692);
nand U5705 (N_5705,N_3476,N_3385);
nand U5706 (N_5706,N_3036,N_3110);
or U5707 (N_5707,N_3491,N_3209);
or U5708 (N_5708,N_4368,N_3518);
nor U5709 (N_5709,N_3039,N_3566);
nand U5710 (N_5710,N_4321,N_3815);
or U5711 (N_5711,N_4213,N_2871);
nand U5712 (N_5712,N_2756,N_3044);
nor U5713 (N_5713,N_4954,N_3952);
nand U5714 (N_5714,N_2837,N_4265);
xor U5715 (N_5715,N_4943,N_2842);
nor U5716 (N_5716,N_3957,N_4089);
or U5717 (N_5717,N_2609,N_4974);
xnor U5718 (N_5718,N_3452,N_3598);
nand U5719 (N_5719,N_3670,N_4907);
nand U5720 (N_5720,N_2923,N_4191);
xor U5721 (N_5721,N_3882,N_2578);
and U5722 (N_5722,N_4469,N_4345);
or U5723 (N_5723,N_2830,N_3736);
nor U5724 (N_5724,N_2547,N_2588);
and U5725 (N_5725,N_4940,N_4186);
and U5726 (N_5726,N_4035,N_4755);
nand U5727 (N_5727,N_4972,N_4133);
or U5728 (N_5728,N_3894,N_3712);
nor U5729 (N_5729,N_4683,N_2927);
and U5730 (N_5730,N_4531,N_2877);
xnor U5731 (N_5731,N_2510,N_3270);
and U5732 (N_5732,N_4897,N_2829);
or U5733 (N_5733,N_2695,N_4220);
nand U5734 (N_5734,N_2774,N_3427);
and U5735 (N_5735,N_3436,N_3691);
nor U5736 (N_5736,N_3915,N_3570);
nor U5737 (N_5737,N_3534,N_3084);
and U5738 (N_5738,N_3190,N_3388);
nand U5739 (N_5739,N_4908,N_4530);
and U5740 (N_5740,N_4003,N_4900);
nor U5741 (N_5741,N_2872,N_3985);
and U5742 (N_5742,N_3383,N_4256);
and U5743 (N_5743,N_3923,N_4624);
nor U5744 (N_5744,N_3560,N_3457);
nor U5745 (N_5745,N_4398,N_3245);
nor U5746 (N_5746,N_3445,N_2884);
nand U5747 (N_5747,N_4294,N_3858);
xnor U5748 (N_5748,N_3857,N_3647);
nand U5749 (N_5749,N_4233,N_4164);
and U5750 (N_5750,N_3549,N_4263);
xor U5751 (N_5751,N_3032,N_3447);
and U5752 (N_5752,N_2769,N_2937);
or U5753 (N_5753,N_4878,N_3757);
and U5754 (N_5754,N_3496,N_4509);
and U5755 (N_5755,N_2707,N_3950);
or U5756 (N_5756,N_4834,N_4212);
nand U5757 (N_5757,N_4984,N_4525);
xor U5758 (N_5758,N_3973,N_4454);
nand U5759 (N_5759,N_4801,N_3956);
or U5760 (N_5760,N_4621,N_3810);
nor U5761 (N_5761,N_3537,N_4465);
nor U5762 (N_5762,N_3911,N_2977);
nor U5763 (N_5763,N_4964,N_4367);
and U5764 (N_5764,N_3059,N_2882);
nor U5765 (N_5765,N_3186,N_2717);
or U5766 (N_5766,N_4623,N_4403);
or U5767 (N_5767,N_4785,N_4405);
nand U5768 (N_5768,N_4388,N_3339);
or U5769 (N_5769,N_4221,N_3512);
and U5770 (N_5770,N_3666,N_3590);
or U5771 (N_5771,N_4455,N_4029);
or U5772 (N_5772,N_4811,N_3090);
and U5773 (N_5773,N_4467,N_4510);
nor U5774 (N_5774,N_4602,N_4326);
and U5775 (N_5775,N_4151,N_3338);
and U5776 (N_5776,N_2538,N_4778);
and U5777 (N_5777,N_4547,N_3200);
nand U5778 (N_5778,N_2804,N_4237);
and U5779 (N_5779,N_2954,N_3693);
and U5780 (N_5780,N_3723,N_2868);
xnor U5781 (N_5781,N_3063,N_2591);
or U5782 (N_5782,N_3948,N_3067);
and U5783 (N_5783,N_3189,N_3999);
nand U5784 (N_5784,N_4810,N_4091);
nor U5785 (N_5785,N_2922,N_4112);
xnor U5786 (N_5786,N_4152,N_4664);
or U5787 (N_5787,N_2952,N_3140);
nor U5788 (N_5788,N_2670,N_4741);
and U5789 (N_5789,N_4582,N_4845);
nand U5790 (N_5790,N_4636,N_3620);
and U5791 (N_5791,N_4691,N_3494);
or U5792 (N_5792,N_2990,N_4762);
nor U5793 (N_5793,N_4968,N_4478);
xnor U5794 (N_5794,N_3379,N_4069);
or U5795 (N_5795,N_3460,N_4267);
nor U5796 (N_5796,N_3940,N_3787);
xor U5797 (N_5797,N_3016,N_4100);
and U5798 (N_5798,N_4192,N_3354);
xnor U5799 (N_5799,N_3924,N_4496);
nand U5800 (N_5800,N_2760,N_4821);
nor U5801 (N_5801,N_2936,N_4999);
xnor U5802 (N_5802,N_3124,N_4399);
or U5803 (N_5803,N_4644,N_2567);
and U5804 (N_5804,N_4814,N_3104);
or U5805 (N_5805,N_4815,N_4451);
and U5806 (N_5806,N_3898,N_3906);
and U5807 (N_5807,N_3892,N_4406);
nand U5808 (N_5808,N_4828,N_3307);
nor U5809 (N_5809,N_3662,N_3880);
xor U5810 (N_5810,N_3465,N_2579);
nand U5811 (N_5811,N_3409,N_3614);
or U5812 (N_5812,N_3578,N_3101);
xnor U5813 (N_5813,N_2798,N_4799);
nor U5814 (N_5814,N_3102,N_4619);
xor U5815 (N_5815,N_2832,N_4063);
nor U5816 (N_5816,N_3034,N_3859);
and U5817 (N_5817,N_2831,N_2985);
nand U5818 (N_5818,N_3433,N_2794);
and U5819 (N_5819,N_4493,N_3724);
nand U5820 (N_5820,N_4222,N_2658);
nand U5821 (N_5821,N_3336,N_4796);
and U5822 (N_5822,N_3895,N_3175);
nor U5823 (N_5823,N_3793,N_2905);
nand U5824 (N_5824,N_3192,N_4601);
or U5825 (N_5825,N_3216,N_4360);
nand U5826 (N_5826,N_4565,N_2501);
nor U5827 (N_5827,N_4981,N_2642);
nand U5828 (N_5828,N_3441,N_3758);
and U5829 (N_5829,N_3389,N_3399);
and U5830 (N_5830,N_3804,N_3644);
and U5831 (N_5831,N_2873,N_3277);
and U5832 (N_5832,N_3220,N_2688);
nor U5833 (N_5833,N_4990,N_4545);
or U5834 (N_5834,N_4374,N_4400);
nor U5835 (N_5835,N_3070,N_4059);
nor U5836 (N_5836,N_4146,N_3367);
and U5837 (N_5837,N_4816,N_3832);
xor U5838 (N_5838,N_4095,N_4485);
nor U5839 (N_5839,N_3303,N_3077);
xnor U5840 (N_5840,N_3437,N_4753);
nor U5841 (N_5841,N_3041,N_3150);
and U5842 (N_5842,N_3983,N_4166);
or U5843 (N_5843,N_4124,N_3922);
nand U5844 (N_5844,N_4861,N_4070);
and U5845 (N_5845,N_2576,N_3485);
or U5846 (N_5846,N_2569,N_3337);
nor U5847 (N_5847,N_3602,N_3655);
nor U5848 (N_5848,N_4025,N_4583);
nand U5849 (N_5849,N_4348,N_4286);
or U5850 (N_5850,N_4393,N_3617);
nor U5851 (N_5851,N_3259,N_3481);
xor U5852 (N_5852,N_3916,N_4323);
nor U5853 (N_5853,N_2522,N_4852);
or U5854 (N_5854,N_3954,N_4891);
or U5855 (N_5855,N_3826,N_3197);
nor U5856 (N_5856,N_4115,N_2715);
or U5857 (N_5857,N_4021,N_3687);
nand U5858 (N_5858,N_3319,N_4989);
nor U5859 (N_5859,N_3612,N_3781);
nor U5860 (N_5860,N_2667,N_2550);
nor U5861 (N_5861,N_4833,N_2867);
xnor U5862 (N_5862,N_3184,N_4384);
or U5863 (N_5863,N_2712,N_3627);
nor U5864 (N_5864,N_4858,N_4473);
nand U5865 (N_5865,N_3403,N_4812);
and U5866 (N_5866,N_2513,N_2753);
nor U5867 (N_5867,N_3795,N_4929);
and U5868 (N_5868,N_3794,N_3178);
or U5869 (N_5869,N_4996,N_2584);
or U5870 (N_5870,N_3565,N_2750);
nor U5871 (N_5871,N_4781,N_3959);
nand U5872 (N_5872,N_4665,N_3238);
nand U5873 (N_5873,N_4910,N_2586);
or U5874 (N_5874,N_3122,N_2944);
and U5875 (N_5875,N_4026,N_4863);
and U5876 (N_5876,N_2887,N_2902);
nor U5877 (N_5877,N_4402,N_4548);
nor U5878 (N_5878,N_3579,N_3603);
nand U5879 (N_5879,N_2718,N_2790);
or U5880 (N_5880,N_3887,N_3402);
nor U5881 (N_5881,N_4293,N_3219);
and U5882 (N_5882,N_4633,N_2644);
or U5883 (N_5883,N_3971,N_3306);
xor U5884 (N_5884,N_2779,N_4518);
xor U5885 (N_5885,N_2777,N_4062);
nand U5886 (N_5886,N_3227,N_4032);
nor U5887 (N_5887,N_3255,N_4053);
or U5888 (N_5888,N_4890,N_2915);
nor U5889 (N_5889,N_4892,N_3393);
or U5890 (N_5890,N_3087,N_2895);
and U5891 (N_5891,N_3264,N_3153);
or U5892 (N_5892,N_4909,N_3449);
nor U5893 (N_5893,N_3960,N_3875);
and U5894 (N_5894,N_3981,N_4540);
xor U5895 (N_5895,N_3395,N_2913);
xor U5896 (N_5896,N_3907,N_4474);
xor U5897 (N_5897,N_2784,N_3682);
nand U5898 (N_5898,N_3052,N_4708);
or U5899 (N_5899,N_4363,N_2986);
nand U5900 (N_5900,N_4797,N_2771);
nand U5901 (N_5901,N_4710,N_4415);
nand U5902 (N_5902,N_4634,N_2544);
nor U5903 (N_5903,N_4357,N_3928);
nor U5904 (N_5904,N_2900,N_4980);
and U5905 (N_5905,N_4018,N_4051);
or U5906 (N_5906,N_3406,N_4870);
or U5907 (N_5907,N_4092,N_2904);
nor U5908 (N_5908,N_4044,N_2652);
nand U5909 (N_5909,N_3903,N_4771);
nand U5910 (N_5910,N_4646,N_4121);
and U5911 (N_5911,N_4871,N_3639);
and U5912 (N_5912,N_4303,N_3581);
nor U5913 (N_5913,N_3525,N_3692);
and U5914 (N_5914,N_2973,N_3526);
and U5915 (N_5915,N_4090,N_4416);
or U5916 (N_5916,N_4550,N_4043);
and U5917 (N_5917,N_2843,N_4515);
and U5918 (N_5918,N_4949,N_4331);
and U5919 (N_5919,N_3185,N_4842);
nand U5920 (N_5920,N_2643,N_4180);
or U5921 (N_5921,N_2615,N_4568);
xor U5922 (N_5922,N_3390,N_2891);
or U5923 (N_5923,N_2669,N_3754);
and U5924 (N_5924,N_3573,N_4822);
nor U5925 (N_5925,N_3925,N_4520);
nor U5926 (N_5926,N_3738,N_4613);
and U5927 (N_5927,N_2593,N_3891);
xor U5928 (N_5928,N_3008,N_2743);
nand U5929 (N_5929,N_3446,N_3613);
nand U5930 (N_5930,N_4306,N_2639);
or U5931 (N_5931,N_2766,N_4607);
nand U5932 (N_5932,N_3094,N_3640);
nor U5933 (N_5933,N_4508,N_2732);
or U5934 (N_5934,N_4015,N_2933);
nor U5935 (N_5935,N_4754,N_3051);
nor U5936 (N_5936,N_3161,N_3062);
and U5937 (N_5937,N_3517,N_2604);
or U5938 (N_5938,N_4849,N_2941);
nand U5939 (N_5939,N_3293,N_4604);
nor U5940 (N_5940,N_4460,N_4489);
or U5941 (N_5941,N_3659,N_2847);
nor U5942 (N_5942,N_3675,N_4948);
nand U5943 (N_5943,N_4184,N_4016);
nor U5944 (N_5944,N_4109,N_4458);
and U5945 (N_5945,N_2982,N_3601);
and U5946 (N_5946,N_4000,N_4820);
and U5947 (N_5947,N_3986,N_4312);
nor U5948 (N_5948,N_3317,N_3762);
xor U5949 (N_5949,N_3769,N_3146);
nor U5950 (N_5950,N_2934,N_4586);
nand U5951 (N_5951,N_2570,N_4718);
nand U5952 (N_5952,N_3325,N_3352);
nand U5953 (N_5953,N_4128,N_3422);
and U5954 (N_5954,N_2889,N_4595);
or U5955 (N_5955,N_3632,N_3174);
and U5956 (N_5956,N_3943,N_3737);
and U5957 (N_5957,N_4911,N_3967);
and U5958 (N_5958,N_4534,N_2623);
or U5959 (N_5959,N_4296,N_2783);
and U5960 (N_5960,N_4889,N_3014);
and U5961 (N_5961,N_3760,N_4206);
or U5962 (N_5962,N_3524,N_4620);
nand U5963 (N_5963,N_3536,N_3362);
xor U5964 (N_5964,N_4953,N_3290);
nor U5965 (N_5965,N_3846,N_4750);
nand U5966 (N_5966,N_4277,N_2816);
nand U5967 (N_5967,N_3749,N_3531);
xor U5968 (N_5968,N_3919,N_3669);
and U5969 (N_5969,N_4442,N_4391);
nor U5970 (N_5970,N_2676,N_4860);
nor U5971 (N_5971,N_4992,N_4716);
nand U5972 (N_5972,N_3417,N_4142);
nor U5973 (N_5973,N_3721,N_3551);
or U5974 (N_5974,N_4189,N_3913);
nor U5975 (N_5975,N_4262,N_3819);
or U5976 (N_5976,N_4717,N_3144);
and U5977 (N_5977,N_3047,N_2827);
and U5978 (N_5978,N_3866,N_3628);
nand U5979 (N_5979,N_3872,N_2606);
nand U5980 (N_5980,N_2949,N_3680);
xnor U5981 (N_5981,N_3665,N_4932);
and U5982 (N_5982,N_3114,N_3247);
nor U5983 (N_5983,N_3001,N_3994);
nand U5984 (N_5984,N_2699,N_4302);
or U5985 (N_5985,N_2881,N_4392);
or U5986 (N_5986,N_3498,N_3492);
or U5987 (N_5987,N_3006,N_4080);
nand U5988 (N_5988,N_2647,N_4605);
or U5989 (N_5989,N_3813,N_4287);
nor U5990 (N_5990,N_3226,N_4970);
and U5991 (N_5991,N_2655,N_2998);
or U5992 (N_5992,N_3108,N_4019);
nand U5993 (N_5993,N_2946,N_4083);
and U5994 (N_5994,N_4590,N_4449);
and U5995 (N_5995,N_3979,N_3678);
or U5996 (N_5996,N_3480,N_4792);
nand U5997 (N_5997,N_4207,N_3818);
nand U5998 (N_5998,N_4259,N_3093);
nand U5999 (N_5999,N_2573,N_2722);
or U6000 (N_6000,N_2685,N_4205);
and U6001 (N_6001,N_3471,N_4328);
nand U6002 (N_6002,N_4396,N_3233);
or U6003 (N_6003,N_4219,N_4788);
nor U6004 (N_6004,N_3519,N_4113);
nor U6005 (N_6005,N_2983,N_3007);
nand U6006 (N_6006,N_3914,N_2502);
or U6007 (N_6007,N_2899,N_2529);
nand U6008 (N_6008,N_4066,N_3700);
or U6009 (N_6009,N_3830,N_2508);
nor U6010 (N_6010,N_2855,N_4921);
or U6011 (N_6011,N_3528,N_3870);
nor U6012 (N_6012,N_3530,N_3350);
and U6013 (N_6013,N_4902,N_3141);
xnor U6014 (N_6014,N_2725,N_3253);
nor U6015 (N_6015,N_2742,N_4480);
xnor U6016 (N_6016,N_4351,N_4427);
xor U6017 (N_6017,N_3702,N_4419);
xor U6018 (N_6018,N_3058,N_4919);
nor U6019 (N_6019,N_4504,N_2600);
nor U6020 (N_6020,N_4337,N_4730);
or U6021 (N_6021,N_4020,N_4111);
nand U6022 (N_6022,N_4680,N_4679);
nand U6023 (N_6023,N_4752,N_4963);
nor U6024 (N_6024,N_3942,N_3643);
or U6025 (N_6025,N_3688,N_2509);
and U6026 (N_6026,N_4120,N_3968);
and U6027 (N_6027,N_2730,N_4067);
nor U6028 (N_6028,N_2763,N_3747);
or U6029 (N_6029,N_2862,N_4894);
nand U6030 (N_6030,N_3228,N_2709);
or U6031 (N_6031,N_3683,N_4823);
and U6032 (N_6032,N_3097,N_3776);
and U6033 (N_6033,N_3301,N_4425);
nand U6034 (N_6034,N_3294,N_4462);
or U6035 (N_6035,N_3421,N_3195);
nand U6036 (N_6036,N_2999,N_4696);
nor U6037 (N_6037,N_4245,N_2736);
nand U6038 (N_6038,N_3489,N_4893);
nand U6039 (N_6039,N_3785,N_3927);
nor U6040 (N_6040,N_2601,N_2992);
and U6041 (N_6041,N_4874,N_4543);
nand U6042 (N_6042,N_4864,N_2793);
nand U6043 (N_6043,N_4441,N_3497);
and U6044 (N_6044,N_3788,N_3509);
nand U6045 (N_6045,N_4503,N_2539);
nor U6046 (N_6046,N_4649,N_3420);
and U6047 (N_6047,N_2561,N_4269);
and U6048 (N_6048,N_3965,N_3467);
and U6049 (N_6049,N_3493,N_3308);
or U6050 (N_6050,N_4104,N_4017);
nor U6051 (N_6051,N_3280,N_4773);
and U6052 (N_6052,N_4336,N_4395);
and U6053 (N_6053,N_3686,N_4668);
xor U6054 (N_6054,N_4177,N_4096);
or U6055 (N_6055,N_4747,N_4770);
and U6056 (N_6056,N_3890,N_4251);
nand U6057 (N_6057,N_3546,N_4093);
or U6058 (N_6058,N_4487,N_4955);
and U6059 (N_6059,N_3878,N_4937);
nand U6060 (N_6060,N_4569,N_4840);
xnor U6061 (N_6061,N_4214,N_4183);
nand U6062 (N_6062,N_4041,N_4013);
nor U6063 (N_6063,N_4195,N_4466);
or U6064 (N_6064,N_2878,N_2840);
nand U6065 (N_6065,N_4782,N_2930);
and U6066 (N_6066,N_3029,N_2863);
nor U6067 (N_6067,N_3844,N_4359);
and U6068 (N_6068,N_2848,N_4229);
nor U6069 (N_6069,N_4800,N_3746);
xor U6070 (N_6070,N_4922,N_4241);
nand U6071 (N_6071,N_2546,N_4958);
nand U6072 (N_6072,N_4798,N_4536);
or U6073 (N_6073,N_4761,N_4862);
nor U6074 (N_6074,N_4470,N_2929);
nor U6075 (N_6075,N_3461,N_4868);
and U6076 (N_6076,N_3777,N_3042);
xnor U6077 (N_6077,N_2764,N_4226);
nand U6078 (N_6078,N_4169,N_3964);
nand U6079 (N_6079,N_2616,N_3982);
nor U6080 (N_6080,N_3726,N_4956);
or U6081 (N_6081,N_4325,N_4647);
or U6082 (N_6082,N_3020,N_4342);
nor U6083 (N_6083,N_3315,N_3134);
or U6084 (N_6084,N_3396,N_4944);
xnor U6085 (N_6085,N_3113,N_4047);
nor U6086 (N_6086,N_4068,N_4866);
nand U6087 (N_6087,N_4678,N_3131);
nor U6088 (N_6088,N_4118,N_4042);
nor U6089 (N_6089,N_2911,N_2968);
nand U6090 (N_6090,N_3462,N_4434);
or U6091 (N_6091,N_3374,N_2697);
nor U6092 (N_6092,N_4793,N_4772);
or U6093 (N_6093,N_4147,N_3281);
nand U6094 (N_6094,N_2535,N_3829);
and U6095 (N_6095,N_3529,N_2541);
and U6096 (N_6096,N_2516,N_3331);
nand U6097 (N_6097,N_2572,N_3275);
or U6098 (N_6098,N_4596,N_3548);
nand U6099 (N_6099,N_3025,N_3909);
and U6100 (N_6100,N_2906,N_3196);
nand U6101 (N_6101,N_4244,N_3106);
nand U6102 (N_6102,N_3802,N_4615);
nor U6103 (N_6103,N_2703,N_3221);
or U6104 (N_6104,N_4310,N_4365);
or U6105 (N_6105,N_3431,N_4758);
and U6106 (N_6106,N_2747,N_4748);
or U6107 (N_6107,N_4706,N_3278);
nand U6108 (N_6108,N_4072,N_4254);
or U6109 (N_6109,N_3707,N_4272);
nand U6110 (N_6110,N_4141,N_4960);
nand U6111 (N_6111,N_3649,N_3596);
nor U6112 (N_6112,N_2689,N_3450);
nor U6113 (N_6113,N_4290,N_3741);
xor U6114 (N_6114,N_4276,N_4711);
or U6115 (N_6115,N_2651,N_4857);
or U6116 (N_6116,N_4671,N_2859);
and U6117 (N_6117,N_2974,N_2711);
xor U6118 (N_6118,N_4422,N_4361);
nand U6119 (N_6119,N_3589,N_4561);
nand U6120 (N_6120,N_4505,N_4524);
or U6121 (N_6121,N_4495,N_4975);
nor U6122 (N_6122,N_3133,N_3477);
or U6123 (N_6123,N_3199,N_3115);
and U6124 (N_6124,N_3842,N_4869);
nor U6125 (N_6125,N_3075,N_4650);
and U6126 (N_6126,N_3375,N_4283);
and U6127 (N_6127,N_2748,N_3824);
or U6128 (N_6128,N_3722,N_3394);
and U6129 (N_6129,N_2960,N_3752);
xor U6130 (N_6130,N_3690,N_3424);
nand U6131 (N_6131,N_4704,N_3789);
and U6132 (N_6132,N_3095,N_4689);
and U6133 (N_6133,N_4882,N_3755);
or U6134 (N_6134,N_4950,N_4535);
nand U6135 (N_6135,N_3469,N_2782);
or U6136 (N_6136,N_3258,N_3843);
and U6137 (N_6137,N_3580,N_3172);
or U6138 (N_6138,N_4609,N_3801);
nand U6139 (N_6139,N_2659,N_2551);
or U6140 (N_6140,N_3330,N_4951);
or U6141 (N_6141,N_2835,N_2809);
or U6142 (N_6142,N_4234,N_3023);
nor U6143 (N_6143,N_4498,N_4697);
nor U6144 (N_6144,N_3698,N_2511);
and U6145 (N_6145,N_2966,N_3635);
nor U6146 (N_6146,N_3171,N_3714);
nor U6147 (N_6147,N_2518,N_2587);
or U6148 (N_6148,N_3599,N_2920);
or U6149 (N_6149,N_4150,N_4103);
and U6150 (N_6150,N_3817,N_3413);
nand U6151 (N_6151,N_3939,N_4333);
nand U6152 (N_6152,N_3778,N_4381);
nand U6153 (N_6153,N_3893,N_4131);
and U6154 (N_6154,N_4412,N_3715);
nor U6155 (N_6155,N_4553,N_3138);
or U6156 (N_6156,N_2641,N_3835);
or U6157 (N_6157,N_2869,N_3676);
nand U6158 (N_6158,N_4340,N_4446);
nand U6159 (N_6159,N_4444,N_4973);
nor U6160 (N_6160,N_2657,N_4156);
or U6161 (N_6161,N_3775,N_4223);
nor U6162 (N_6162,N_2825,N_4935);
and U6163 (N_6163,N_4197,N_4589);
nand U6164 (N_6164,N_2696,N_2500);
and U6165 (N_6165,N_3938,N_3215);
nor U6166 (N_6166,N_2517,N_3137);
or U6167 (N_6167,N_3504,N_2620);
and U6168 (N_6168,N_4413,N_4235);
and U6169 (N_6169,N_2521,N_3405);
nand U6170 (N_6170,N_4300,N_3770);
nor U6171 (N_6171,N_3637,N_2852);
nor U6172 (N_6172,N_3849,N_4443);
nor U6173 (N_6173,N_2556,N_3852);
xor U6174 (N_6174,N_3798,N_4311);
nand U6175 (N_6175,N_3241,N_3947);
or U6176 (N_6176,N_3155,N_3332);
nor U6177 (N_6177,N_4600,N_3696);
or U6178 (N_6178,N_4210,N_3901);
and U6179 (N_6179,N_2650,N_4471);
nand U6180 (N_6180,N_4353,N_4009);
or U6181 (N_6181,N_4738,N_3458);
nand U6182 (N_6182,N_2893,N_3218);
or U6183 (N_6183,N_3464,N_4732);
and U6184 (N_6184,N_4248,N_2548);
and U6185 (N_6185,N_3845,N_3297);
nand U6186 (N_6186,N_4279,N_4511);
xnor U6187 (N_6187,N_3118,N_3740);
or U6188 (N_6188,N_3263,N_3046);
nor U6189 (N_6189,N_2739,N_3989);
xor U6190 (N_6190,N_4701,N_4257);
xor U6191 (N_6191,N_3037,N_3541);
nand U6192 (N_6192,N_3679,N_4201);
or U6193 (N_6193,N_4159,N_3710);
or U6194 (N_6194,N_4081,N_3864);
nor U6195 (N_6195,N_3071,N_4599);
and U6196 (N_6196,N_4199,N_2797);
or U6197 (N_6197,N_4007,N_4225);
nor U6198 (N_6198,N_2820,N_4280);
nand U6199 (N_6199,N_2633,N_4071);
and U6200 (N_6200,N_3980,N_4962);
or U6201 (N_6201,N_2599,N_4270);
nor U6202 (N_6202,N_3444,N_3169);
and U6203 (N_6203,N_4529,N_3876);
nand U6204 (N_6204,N_3975,N_3930);
and U6205 (N_6205,N_4122,N_4603);
and U6206 (N_6206,N_4289,N_2568);
xor U6207 (N_6207,N_2773,N_2917);
nand U6208 (N_6208,N_2980,N_4230);
xor U6209 (N_6209,N_4971,N_2645);
xnor U6210 (N_6210,N_3904,N_2890);
nor U6211 (N_6211,N_3816,N_4905);
xnor U6212 (N_6212,N_4418,N_3879);
nor U6213 (N_6213,N_4375,N_3152);
xnor U6214 (N_6214,N_2708,N_3407);
nand U6215 (N_6215,N_4688,N_2596);
nand U6216 (N_6216,N_3000,N_4566);
nor U6217 (N_6217,N_3302,N_4208);
and U6218 (N_6218,N_3229,N_3569);
and U6219 (N_6219,N_4854,N_3720);
nand U6220 (N_6220,N_3382,N_4108);
or U6221 (N_6221,N_3861,N_4803);
or U6222 (N_6222,N_3004,N_3289);
nor U6223 (N_6223,N_2523,N_2737);
nor U6224 (N_6224,N_2931,N_3624);
and U6225 (N_6225,N_4746,N_4597);
and U6226 (N_6226,N_4114,N_4318);
nand U6227 (N_6227,N_4606,N_4389);
xnor U6228 (N_6228,N_4354,N_4674);
nor U6229 (N_6229,N_3932,N_4562);
nand U6230 (N_6230,N_4438,N_3917);
or U6231 (N_6231,N_4737,N_3591);
nand U6232 (N_6232,N_2956,N_3204);
and U6233 (N_6233,N_2684,N_4252);
or U6234 (N_6234,N_4227,N_4382);
or U6235 (N_6235,N_2870,N_3918);
xnor U6236 (N_6236,N_2735,N_3360);
and U6237 (N_6237,N_3309,N_2953);
or U6238 (N_6238,N_4110,N_4453);
nor U6239 (N_6239,N_3056,N_4339);
and U6240 (N_6240,N_3831,N_2574);
and U6241 (N_6241,N_4486,N_4238);
nand U6242 (N_6242,N_4977,N_4082);
or U6243 (N_6243,N_2943,N_3704);
and U6244 (N_6244,N_4924,N_3905);
and U6245 (N_6245,N_2833,N_3100);
xor U6246 (N_6246,N_3418,N_4174);
nand U6247 (N_6247,N_3066,N_3434);
nand U6248 (N_6248,N_3089,N_3558);
and U6249 (N_6249,N_4818,N_4735);
nand U6250 (N_6250,N_2942,N_3177);
or U6251 (N_6251,N_3503,N_3984);
nor U6252 (N_6252,N_3665,N_3215);
and U6253 (N_6253,N_4891,N_4303);
nand U6254 (N_6254,N_4250,N_4197);
xnor U6255 (N_6255,N_4255,N_3312);
or U6256 (N_6256,N_2851,N_4017);
or U6257 (N_6257,N_3935,N_3234);
and U6258 (N_6258,N_3346,N_2988);
or U6259 (N_6259,N_3344,N_3424);
nor U6260 (N_6260,N_3896,N_4084);
nor U6261 (N_6261,N_4018,N_4646);
or U6262 (N_6262,N_4026,N_4800);
nor U6263 (N_6263,N_2926,N_3409);
nand U6264 (N_6264,N_3376,N_2881);
xor U6265 (N_6265,N_3897,N_2798);
xnor U6266 (N_6266,N_3630,N_4474);
nand U6267 (N_6267,N_2559,N_4031);
nor U6268 (N_6268,N_2990,N_2613);
nor U6269 (N_6269,N_4326,N_2945);
and U6270 (N_6270,N_3030,N_3446);
xor U6271 (N_6271,N_3669,N_3534);
nor U6272 (N_6272,N_4856,N_4155);
nor U6273 (N_6273,N_4297,N_3267);
nand U6274 (N_6274,N_2573,N_3812);
or U6275 (N_6275,N_4078,N_4789);
nor U6276 (N_6276,N_2772,N_4815);
xor U6277 (N_6277,N_4824,N_3547);
or U6278 (N_6278,N_4685,N_3795);
and U6279 (N_6279,N_2638,N_4461);
nor U6280 (N_6280,N_2972,N_2569);
or U6281 (N_6281,N_3593,N_4888);
and U6282 (N_6282,N_2614,N_4624);
or U6283 (N_6283,N_3643,N_4871);
nor U6284 (N_6284,N_4196,N_4812);
and U6285 (N_6285,N_4841,N_4574);
xor U6286 (N_6286,N_3641,N_4508);
and U6287 (N_6287,N_3700,N_2644);
and U6288 (N_6288,N_3242,N_2834);
nand U6289 (N_6289,N_2652,N_3981);
and U6290 (N_6290,N_4256,N_4262);
or U6291 (N_6291,N_3028,N_2602);
and U6292 (N_6292,N_3094,N_4627);
xnor U6293 (N_6293,N_3565,N_3491);
nand U6294 (N_6294,N_4620,N_3185);
and U6295 (N_6295,N_3007,N_2715);
nor U6296 (N_6296,N_4712,N_3331);
nor U6297 (N_6297,N_3614,N_4810);
nor U6298 (N_6298,N_3123,N_4837);
nor U6299 (N_6299,N_4458,N_4654);
nor U6300 (N_6300,N_3627,N_3394);
nand U6301 (N_6301,N_3868,N_2727);
and U6302 (N_6302,N_3572,N_4746);
nor U6303 (N_6303,N_4104,N_2763);
or U6304 (N_6304,N_4756,N_4524);
nor U6305 (N_6305,N_4881,N_3144);
and U6306 (N_6306,N_3152,N_3084);
nor U6307 (N_6307,N_3009,N_4141);
xor U6308 (N_6308,N_3624,N_3682);
nand U6309 (N_6309,N_3394,N_4311);
or U6310 (N_6310,N_2670,N_2554);
and U6311 (N_6311,N_4568,N_3732);
nor U6312 (N_6312,N_3087,N_3654);
and U6313 (N_6313,N_3002,N_4849);
nor U6314 (N_6314,N_3894,N_2881);
xor U6315 (N_6315,N_4740,N_3535);
nand U6316 (N_6316,N_2970,N_3200);
nand U6317 (N_6317,N_2800,N_3542);
nor U6318 (N_6318,N_2852,N_4350);
nand U6319 (N_6319,N_3372,N_4131);
nor U6320 (N_6320,N_3079,N_3026);
nor U6321 (N_6321,N_2998,N_4003);
nand U6322 (N_6322,N_3091,N_2600);
and U6323 (N_6323,N_2662,N_4023);
nand U6324 (N_6324,N_4477,N_2581);
nand U6325 (N_6325,N_2719,N_4357);
xnor U6326 (N_6326,N_3820,N_3728);
nand U6327 (N_6327,N_4502,N_3812);
and U6328 (N_6328,N_2861,N_4681);
or U6329 (N_6329,N_4357,N_3986);
xnor U6330 (N_6330,N_4289,N_3382);
or U6331 (N_6331,N_3545,N_3677);
nand U6332 (N_6332,N_3906,N_4716);
and U6333 (N_6333,N_4468,N_4572);
or U6334 (N_6334,N_4463,N_2912);
nand U6335 (N_6335,N_2851,N_4802);
and U6336 (N_6336,N_4278,N_3667);
and U6337 (N_6337,N_2639,N_3447);
nand U6338 (N_6338,N_3839,N_2651);
nand U6339 (N_6339,N_2703,N_4367);
xor U6340 (N_6340,N_3241,N_3451);
or U6341 (N_6341,N_2858,N_4530);
nor U6342 (N_6342,N_3707,N_4515);
nor U6343 (N_6343,N_4665,N_4340);
xnor U6344 (N_6344,N_4392,N_4312);
nor U6345 (N_6345,N_2563,N_4587);
xnor U6346 (N_6346,N_3246,N_3423);
and U6347 (N_6347,N_2571,N_3638);
xnor U6348 (N_6348,N_2632,N_3156);
nand U6349 (N_6349,N_4530,N_3283);
and U6350 (N_6350,N_4658,N_3531);
nor U6351 (N_6351,N_3389,N_2923);
or U6352 (N_6352,N_3241,N_4510);
nand U6353 (N_6353,N_2586,N_4676);
and U6354 (N_6354,N_4876,N_3312);
or U6355 (N_6355,N_4493,N_4369);
nand U6356 (N_6356,N_4018,N_3132);
nor U6357 (N_6357,N_3718,N_4287);
nor U6358 (N_6358,N_4291,N_3027);
nor U6359 (N_6359,N_3164,N_4395);
and U6360 (N_6360,N_3367,N_4423);
or U6361 (N_6361,N_4126,N_3902);
nor U6362 (N_6362,N_4027,N_3938);
nor U6363 (N_6363,N_4476,N_2868);
and U6364 (N_6364,N_4408,N_3773);
or U6365 (N_6365,N_2920,N_4432);
nor U6366 (N_6366,N_3609,N_4440);
and U6367 (N_6367,N_4331,N_4525);
or U6368 (N_6368,N_4766,N_3473);
nor U6369 (N_6369,N_2549,N_4771);
nand U6370 (N_6370,N_3756,N_4675);
or U6371 (N_6371,N_4358,N_3655);
nand U6372 (N_6372,N_3013,N_3995);
nor U6373 (N_6373,N_2668,N_2506);
and U6374 (N_6374,N_2605,N_4915);
or U6375 (N_6375,N_3431,N_2860);
nand U6376 (N_6376,N_4006,N_4083);
and U6377 (N_6377,N_4490,N_3387);
or U6378 (N_6378,N_2904,N_4596);
or U6379 (N_6379,N_3554,N_4807);
xnor U6380 (N_6380,N_2787,N_3674);
and U6381 (N_6381,N_4741,N_4614);
and U6382 (N_6382,N_3676,N_2775);
or U6383 (N_6383,N_4405,N_3209);
xnor U6384 (N_6384,N_3407,N_2575);
and U6385 (N_6385,N_3331,N_3234);
or U6386 (N_6386,N_3317,N_4663);
nor U6387 (N_6387,N_4535,N_3546);
nor U6388 (N_6388,N_2936,N_3675);
nand U6389 (N_6389,N_4880,N_4950);
nand U6390 (N_6390,N_2703,N_4430);
or U6391 (N_6391,N_3039,N_4095);
and U6392 (N_6392,N_4002,N_4304);
nor U6393 (N_6393,N_4164,N_4081);
and U6394 (N_6394,N_3363,N_4975);
and U6395 (N_6395,N_4392,N_4088);
nor U6396 (N_6396,N_3275,N_4420);
and U6397 (N_6397,N_3868,N_2849);
nor U6398 (N_6398,N_3810,N_3862);
or U6399 (N_6399,N_4083,N_3350);
or U6400 (N_6400,N_2950,N_2648);
and U6401 (N_6401,N_4745,N_3891);
xor U6402 (N_6402,N_4818,N_3942);
and U6403 (N_6403,N_4348,N_4791);
and U6404 (N_6404,N_4839,N_4853);
nand U6405 (N_6405,N_2902,N_4076);
nand U6406 (N_6406,N_4401,N_2566);
nand U6407 (N_6407,N_3654,N_3981);
or U6408 (N_6408,N_3779,N_3854);
nand U6409 (N_6409,N_2971,N_4359);
xnor U6410 (N_6410,N_3732,N_3258);
nor U6411 (N_6411,N_3704,N_4135);
or U6412 (N_6412,N_3755,N_3318);
nand U6413 (N_6413,N_4190,N_3278);
nand U6414 (N_6414,N_3968,N_4027);
and U6415 (N_6415,N_4280,N_3489);
nor U6416 (N_6416,N_3528,N_3426);
nor U6417 (N_6417,N_4560,N_2718);
nor U6418 (N_6418,N_4725,N_4700);
nand U6419 (N_6419,N_3308,N_3774);
or U6420 (N_6420,N_4281,N_2667);
xor U6421 (N_6421,N_4938,N_2864);
or U6422 (N_6422,N_3627,N_3102);
or U6423 (N_6423,N_4739,N_4010);
nand U6424 (N_6424,N_3915,N_3874);
nor U6425 (N_6425,N_4626,N_4625);
nand U6426 (N_6426,N_3378,N_4356);
nor U6427 (N_6427,N_4221,N_4480);
nor U6428 (N_6428,N_4495,N_4032);
or U6429 (N_6429,N_4490,N_3143);
nor U6430 (N_6430,N_3366,N_4419);
or U6431 (N_6431,N_3416,N_2938);
nand U6432 (N_6432,N_2631,N_3926);
nor U6433 (N_6433,N_2930,N_2900);
nand U6434 (N_6434,N_4054,N_3920);
nor U6435 (N_6435,N_2726,N_3854);
nand U6436 (N_6436,N_3220,N_4889);
nor U6437 (N_6437,N_4063,N_2820);
nor U6438 (N_6438,N_3914,N_3215);
xnor U6439 (N_6439,N_3210,N_3567);
and U6440 (N_6440,N_3441,N_3764);
and U6441 (N_6441,N_2558,N_4638);
and U6442 (N_6442,N_3629,N_4473);
or U6443 (N_6443,N_3183,N_2519);
nand U6444 (N_6444,N_3525,N_3738);
and U6445 (N_6445,N_3067,N_3520);
xnor U6446 (N_6446,N_4675,N_4851);
nor U6447 (N_6447,N_3815,N_3216);
and U6448 (N_6448,N_4542,N_4500);
and U6449 (N_6449,N_4290,N_3995);
or U6450 (N_6450,N_2790,N_3500);
nor U6451 (N_6451,N_4495,N_3912);
and U6452 (N_6452,N_4327,N_4925);
nand U6453 (N_6453,N_3527,N_4485);
xor U6454 (N_6454,N_4769,N_3376);
or U6455 (N_6455,N_2802,N_3472);
or U6456 (N_6456,N_3426,N_3749);
or U6457 (N_6457,N_3857,N_3990);
or U6458 (N_6458,N_2621,N_2728);
xor U6459 (N_6459,N_3672,N_2880);
and U6460 (N_6460,N_3653,N_4244);
xor U6461 (N_6461,N_2665,N_3715);
nor U6462 (N_6462,N_4052,N_4108);
nor U6463 (N_6463,N_4895,N_3451);
nor U6464 (N_6464,N_3593,N_4695);
xnor U6465 (N_6465,N_3916,N_3912);
and U6466 (N_6466,N_3223,N_4146);
nor U6467 (N_6467,N_2663,N_3189);
nand U6468 (N_6468,N_3763,N_3335);
xor U6469 (N_6469,N_3891,N_4856);
nand U6470 (N_6470,N_3203,N_2913);
nand U6471 (N_6471,N_3622,N_2715);
nand U6472 (N_6472,N_3611,N_4294);
or U6473 (N_6473,N_4469,N_2545);
or U6474 (N_6474,N_2625,N_2919);
or U6475 (N_6475,N_3042,N_3890);
or U6476 (N_6476,N_3792,N_3544);
and U6477 (N_6477,N_4402,N_3663);
and U6478 (N_6478,N_4315,N_4944);
and U6479 (N_6479,N_2531,N_3653);
nor U6480 (N_6480,N_2666,N_4567);
or U6481 (N_6481,N_4832,N_3113);
xnor U6482 (N_6482,N_3774,N_2545);
nand U6483 (N_6483,N_3150,N_3005);
and U6484 (N_6484,N_4398,N_4273);
or U6485 (N_6485,N_2845,N_3387);
nor U6486 (N_6486,N_2585,N_2988);
nand U6487 (N_6487,N_4751,N_4675);
xor U6488 (N_6488,N_3782,N_2678);
and U6489 (N_6489,N_3043,N_3941);
nand U6490 (N_6490,N_4348,N_3369);
nor U6491 (N_6491,N_2808,N_4338);
or U6492 (N_6492,N_2613,N_2988);
nor U6493 (N_6493,N_3094,N_3007);
xnor U6494 (N_6494,N_3491,N_4240);
nand U6495 (N_6495,N_4286,N_3799);
or U6496 (N_6496,N_4427,N_4949);
nand U6497 (N_6497,N_3769,N_3375);
nand U6498 (N_6498,N_4256,N_4066);
nor U6499 (N_6499,N_2637,N_3778);
nor U6500 (N_6500,N_2786,N_3485);
nor U6501 (N_6501,N_2632,N_4005);
nor U6502 (N_6502,N_4474,N_2567);
and U6503 (N_6503,N_3922,N_3822);
nand U6504 (N_6504,N_3064,N_3366);
or U6505 (N_6505,N_2500,N_4289);
nand U6506 (N_6506,N_3595,N_2528);
xnor U6507 (N_6507,N_3268,N_2808);
xor U6508 (N_6508,N_2639,N_4313);
xor U6509 (N_6509,N_3853,N_2930);
nand U6510 (N_6510,N_3048,N_3507);
nand U6511 (N_6511,N_3228,N_3121);
and U6512 (N_6512,N_3814,N_4569);
or U6513 (N_6513,N_4571,N_3778);
nand U6514 (N_6514,N_2987,N_4503);
and U6515 (N_6515,N_3761,N_2816);
and U6516 (N_6516,N_4497,N_3275);
nor U6517 (N_6517,N_3769,N_3871);
or U6518 (N_6518,N_4473,N_3666);
or U6519 (N_6519,N_2853,N_3101);
nor U6520 (N_6520,N_3466,N_3316);
nor U6521 (N_6521,N_4550,N_2740);
and U6522 (N_6522,N_4465,N_2544);
nor U6523 (N_6523,N_3085,N_3934);
nor U6524 (N_6524,N_4471,N_3142);
nor U6525 (N_6525,N_4226,N_4638);
and U6526 (N_6526,N_3331,N_3250);
or U6527 (N_6527,N_3959,N_4515);
nand U6528 (N_6528,N_2786,N_2544);
nand U6529 (N_6529,N_3942,N_2802);
nand U6530 (N_6530,N_3233,N_4625);
xor U6531 (N_6531,N_4770,N_2538);
nor U6532 (N_6532,N_4971,N_4502);
xnor U6533 (N_6533,N_3702,N_2580);
xor U6534 (N_6534,N_4876,N_4543);
nand U6535 (N_6535,N_2985,N_2862);
or U6536 (N_6536,N_3070,N_3722);
nor U6537 (N_6537,N_4690,N_3796);
and U6538 (N_6538,N_3214,N_3709);
nor U6539 (N_6539,N_3729,N_4275);
or U6540 (N_6540,N_2532,N_3009);
or U6541 (N_6541,N_3120,N_3332);
xnor U6542 (N_6542,N_2828,N_3214);
nor U6543 (N_6543,N_2888,N_3918);
xor U6544 (N_6544,N_3032,N_3974);
or U6545 (N_6545,N_4742,N_3280);
nand U6546 (N_6546,N_4126,N_2883);
and U6547 (N_6547,N_3847,N_3320);
nand U6548 (N_6548,N_3827,N_4009);
and U6549 (N_6549,N_2902,N_4481);
xnor U6550 (N_6550,N_4933,N_3706);
nand U6551 (N_6551,N_2805,N_4973);
nand U6552 (N_6552,N_4489,N_3745);
nor U6553 (N_6553,N_3950,N_4086);
nor U6554 (N_6554,N_4987,N_4605);
nor U6555 (N_6555,N_3530,N_3012);
or U6556 (N_6556,N_3520,N_2680);
or U6557 (N_6557,N_4281,N_4460);
or U6558 (N_6558,N_4299,N_4504);
or U6559 (N_6559,N_4062,N_4433);
and U6560 (N_6560,N_3078,N_3224);
and U6561 (N_6561,N_4939,N_2644);
nor U6562 (N_6562,N_4636,N_3290);
nor U6563 (N_6563,N_3144,N_4429);
or U6564 (N_6564,N_3501,N_3907);
xnor U6565 (N_6565,N_2790,N_3627);
and U6566 (N_6566,N_4949,N_4013);
nand U6567 (N_6567,N_4672,N_4324);
nand U6568 (N_6568,N_3223,N_4008);
nor U6569 (N_6569,N_4354,N_4859);
xor U6570 (N_6570,N_3006,N_3316);
nor U6571 (N_6571,N_3187,N_2603);
xor U6572 (N_6572,N_3097,N_4695);
and U6573 (N_6573,N_4364,N_4991);
and U6574 (N_6574,N_3522,N_3865);
or U6575 (N_6575,N_3349,N_3645);
xor U6576 (N_6576,N_2853,N_2876);
and U6577 (N_6577,N_2987,N_3825);
nor U6578 (N_6578,N_3116,N_4523);
nor U6579 (N_6579,N_4988,N_4806);
and U6580 (N_6580,N_3795,N_4460);
nand U6581 (N_6581,N_4986,N_3867);
or U6582 (N_6582,N_2895,N_2565);
nand U6583 (N_6583,N_2919,N_3257);
nand U6584 (N_6584,N_3623,N_4050);
and U6585 (N_6585,N_3498,N_2575);
nand U6586 (N_6586,N_4265,N_4458);
and U6587 (N_6587,N_2911,N_3457);
or U6588 (N_6588,N_4581,N_3460);
nor U6589 (N_6589,N_4489,N_4839);
and U6590 (N_6590,N_4053,N_2896);
nand U6591 (N_6591,N_2955,N_3594);
or U6592 (N_6592,N_2506,N_2871);
nor U6593 (N_6593,N_4778,N_4393);
nor U6594 (N_6594,N_3065,N_4252);
nand U6595 (N_6595,N_4586,N_4360);
nand U6596 (N_6596,N_2721,N_2627);
nand U6597 (N_6597,N_3016,N_2571);
nor U6598 (N_6598,N_3579,N_3336);
and U6599 (N_6599,N_4530,N_4362);
and U6600 (N_6600,N_3643,N_4524);
nor U6601 (N_6601,N_3419,N_4147);
nand U6602 (N_6602,N_4216,N_3206);
and U6603 (N_6603,N_4669,N_2954);
nor U6604 (N_6604,N_3108,N_3789);
and U6605 (N_6605,N_3921,N_4709);
nor U6606 (N_6606,N_4993,N_4127);
nor U6607 (N_6607,N_4657,N_4679);
nor U6608 (N_6608,N_3119,N_4822);
and U6609 (N_6609,N_2926,N_3048);
and U6610 (N_6610,N_2771,N_4248);
or U6611 (N_6611,N_3170,N_2643);
nor U6612 (N_6612,N_3083,N_3723);
or U6613 (N_6613,N_4128,N_2800);
nor U6614 (N_6614,N_3758,N_4877);
xor U6615 (N_6615,N_4721,N_3147);
nor U6616 (N_6616,N_3641,N_3066);
nor U6617 (N_6617,N_4623,N_3001);
nor U6618 (N_6618,N_3161,N_3043);
or U6619 (N_6619,N_2554,N_3958);
or U6620 (N_6620,N_3773,N_2657);
nand U6621 (N_6621,N_2875,N_3931);
or U6622 (N_6622,N_2614,N_3931);
nor U6623 (N_6623,N_3376,N_3783);
and U6624 (N_6624,N_2659,N_3660);
nand U6625 (N_6625,N_3805,N_4528);
and U6626 (N_6626,N_3096,N_2787);
nor U6627 (N_6627,N_3794,N_2964);
nor U6628 (N_6628,N_4556,N_3585);
and U6629 (N_6629,N_4701,N_3835);
or U6630 (N_6630,N_2944,N_4122);
and U6631 (N_6631,N_3870,N_2757);
nor U6632 (N_6632,N_3888,N_2623);
and U6633 (N_6633,N_3855,N_3669);
or U6634 (N_6634,N_4690,N_4765);
nor U6635 (N_6635,N_4684,N_2798);
nor U6636 (N_6636,N_2717,N_3773);
nand U6637 (N_6637,N_2983,N_2844);
nor U6638 (N_6638,N_2798,N_2783);
and U6639 (N_6639,N_4594,N_3382);
or U6640 (N_6640,N_2784,N_2845);
nand U6641 (N_6641,N_4608,N_3250);
and U6642 (N_6642,N_4683,N_2891);
and U6643 (N_6643,N_4065,N_2515);
or U6644 (N_6644,N_2578,N_3713);
and U6645 (N_6645,N_2740,N_3941);
nand U6646 (N_6646,N_2533,N_2808);
or U6647 (N_6647,N_4834,N_3729);
nor U6648 (N_6648,N_2935,N_2670);
nand U6649 (N_6649,N_4551,N_3211);
or U6650 (N_6650,N_4660,N_4090);
and U6651 (N_6651,N_4975,N_4188);
and U6652 (N_6652,N_4139,N_3772);
or U6653 (N_6653,N_2746,N_3635);
or U6654 (N_6654,N_2712,N_2683);
nand U6655 (N_6655,N_2844,N_4598);
xor U6656 (N_6656,N_4477,N_2663);
nand U6657 (N_6657,N_4284,N_4599);
nor U6658 (N_6658,N_4258,N_3688);
or U6659 (N_6659,N_3767,N_4324);
or U6660 (N_6660,N_3749,N_3514);
nor U6661 (N_6661,N_2718,N_2935);
and U6662 (N_6662,N_4441,N_4929);
or U6663 (N_6663,N_2962,N_3720);
and U6664 (N_6664,N_2875,N_3952);
nand U6665 (N_6665,N_3600,N_4794);
and U6666 (N_6666,N_3415,N_3823);
nand U6667 (N_6667,N_2683,N_2576);
or U6668 (N_6668,N_3917,N_2975);
nor U6669 (N_6669,N_4453,N_4995);
nor U6670 (N_6670,N_2767,N_2977);
xnor U6671 (N_6671,N_3710,N_4473);
nor U6672 (N_6672,N_3076,N_3328);
nand U6673 (N_6673,N_3983,N_3914);
and U6674 (N_6674,N_3779,N_4616);
or U6675 (N_6675,N_3586,N_2816);
nand U6676 (N_6676,N_4253,N_3466);
nor U6677 (N_6677,N_4853,N_4496);
nor U6678 (N_6678,N_2794,N_3772);
nor U6679 (N_6679,N_4484,N_2874);
nand U6680 (N_6680,N_4155,N_4461);
nand U6681 (N_6681,N_3872,N_2564);
or U6682 (N_6682,N_2825,N_4132);
nor U6683 (N_6683,N_2972,N_4589);
nor U6684 (N_6684,N_3991,N_3409);
and U6685 (N_6685,N_4603,N_4785);
or U6686 (N_6686,N_3734,N_4510);
and U6687 (N_6687,N_3636,N_2583);
nor U6688 (N_6688,N_2668,N_4698);
nand U6689 (N_6689,N_4989,N_3199);
xnor U6690 (N_6690,N_3727,N_3123);
xnor U6691 (N_6691,N_4780,N_4329);
nand U6692 (N_6692,N_3204,N_4247);
nand U6693 (N_6693,N_3381,N_4081);
and U6694 (N_6694,N_3735,N_4157);
and U6695 (N_6695,N_3224,N_4318);
nand U6696 (N_6696,N_4084,N_3320);
nor U6697 (N_6697,N_4331,N_3608);
nor U6698 (N_6698,N_2592,N_2522);
or U6699 (N_6699,N_3821,N_4550);
xor U6700 (N_6700,N_3904,N_3864);
and U6701 (N_6701,N_3999,N_4418);
nor U6702 (N_6702,N_3682,N_3072);
nor U6703 (N_6703,N_3972,N_3539);
and U6704 (N_6704,N_4321,N_4384);
and U6705 (N_6705,N_4228,N_2550);
nor U6706 (N_6706,N_2741,N_3005);
nand U6707 (N_6707,N_3346,N_4466);
and U6708 (N_6708,N_3635,N_2650);
and U6709 (N_6709,N_3119,N_4824);
nor U6710 (N_6710,N_4325,N_3493);
and U6711 (N_6711,N_4724,N_4126);
nand U6712 (N_6712,N_4386,N_4840);
or U6713 (N_6713,N_4911,N_4110);
nand U6714 (N_6714,N_2587,N_4141);
or U6715 (N_6715,N_2599,N_4256);
nand U6716 (N_6716,N_2615,N_3462);
nor U6717 (N_6717,N_4160,N_4227);
nand U6718 (N_6718,N_3631,N_3695);
xor U6719 (N_6719,N_2648,N_3934);
nor U6720 (N_6720,N_2994,N_3279);
nor U6721 (N_6721,N_3897,N_4124);
nor U6722 (N_6722,N_4311,N_3016);
nand U6723 (N_6723,N_4222,N_4917);
nor U6724 (N_6724,N_4693,N_2687);
or U6725 (N_6725,N_4184,N_4165);
or U6726 (N_6726,N_3423,N_3726);
xor U6727 (N_6727,N_3695,N_4683);
nor U6728 (N_6728,N_4740,N_3691);
nor U6729 (N_6729,N_4659,N_3345);
and U6730 (N_6730,N_3049,N_4667);
nand U6731 (N_6731,N_3968,N_2905);
and U6732 (N_6732,N_4675,N_4486);
and U6733 (N_6733,N_4292,N_4924);
and U6734 (N_6734,N_4066,N_3767);
nand U6735 (N_6735,N_4438,N_4513);
xnor U6736 (N_6736,N_4363,N_3970);
and U6737 (N_6737,N_2706,N_4085);
nor U6738 (N_6738,N_4398,N_4749);
or U6739 (N_6739,N_2520,N_3719);
or U6740 (N_6740,N_3528,N_3210);
nand U6741 (N_6741,N_3333,N_4557);
nand U6742 (N_6742,N_4283,N_3977);
nor U6743 (N_6743,N_2729,N_2952);
xnor U6744 (N_6744,N_3479,N_2802);
nand U6745 (N_6745,N_3577,N_4174);
nor U6746 (N_6746,N_2801,N_4775);
or U6747 (N_6747,N_4925,N_3772);
nor U6748 (N_6748,N_4845,N_4714);
nor U6749 (N_6749,N_4357,N_3284);
or U6750 (N_6750,N_3254,N_4260);
and U6751 (N_6751,N_4495,N_4655);
or U6752 (N_6752,N_3178,N_4438);
and U6753 (N_6753,N_3806,N_2516);
nand U6754 (N_6754,N_4060,N_2960);
xnor U6755 (N_6755,N_2985,N_2774);
nand U6756 (N_6756,N_2870,N_3640);
xnor U6757 (N_6757,N_3390,N_3562);
or U6758 (N_6758,N_3366,N_4502);
nand U6759 (N_6759,N_3929,N_3943);
xnor U6760 (N_6760,N_3501,N_2615);
or U6761 (N_6761,N_4414,N_4426);
nand U6762 (N_6762,N_4885,N_3307);
xor U6763 (N_6763,N_3380,N_3459);
or U6764 (N_6764,N_3544,N_2695);
xor U6765 (N_6765,N_3315,N_4212);
nor U6766 (N_6766,N_3582,N_2878);
nor U6767 (N_6767,N_4009,N_2930);
nand U6768 (N_6768,N_4006,N_4628);
xnor U6769 (N_6769,N_4841,N_2823);
xor U6770 (N_6770,N_3866,N_4086);
or U6771 (N_6771,N_3448,N_2748);
nand U6772 (N_6772,N_2730,N_4374);
and U6773 (N_6773,N_3686,N_3483);
nor U6774 (N_6774,N_3033,N_3566);
nor U6775 (N_6775,N_4676,N_4702);
nand U6776 (N_6776,N_2594,N_3419);
nand U6777 (N_6777,N_4019,N_4160);
xor U6778 (N_6778,N_4462,N_4658);
xor U6779 (N_6779,N_2601,N_2999);
nand U6780 (N_6780,N_2556,N_4287);
nor U6781 (N_6781,N_3464,N_4018);
and U6782 (N_6782,N_3971,N_3482);
or U6783 (N_6783,N_4321,N_4520);
or U6784 (N_6784,N_4455,N_2817);
nor U6785 (N_6785,N_4331,N_3569);
and U6786 (N_6786,N_2563,N_3993);
or U6787 (N_6787,N_2849,N_4915);
or U6788 (N_6788,N_4188,N_4769);
and U6789 (N_6789,N_3298,N_3142);
nand U6790 (N_6790,N_3368,N_4819);
or U6791 (N_6791,N_3209,N_2695);
nor U6792 (N_6792,N_3341,N_4623);
or U6793 (N_6793,N_4357,N_3492);
or U6794 (N_6794,N_2919,N_3329);
nor U6795 (N_6795,N_3289,N_2681);
nand U6796 (N_6796,N_4956,N_2534);
or U6797 (N_6797,N_2867,N_3359);
nor U6798 (N_6798,N_3033,N_3223);
xor U6799 (N_6799,N_4972,N_2791);
xor U6800 (N_6800,N_3038,N_4063);
nand U6801 (N_6801,N_2552,N_3240);
nor U6802 (N_6802,N_2561,N_2703);
or U6803 (N_6803,N_2821,N_3717);
and U6804 (N_6804,N_3996,N_4199);
and U6805 (N_6805,N_3235,N_3692);
nor U6806 (N_6806,N_3939,N_3278);
nor U6807 (N_6807,N_4539,N_4118);
nor U6808 (N_6808,N_3021,N_4365);
and U6809 (N_6809,N_4162,N_4302);
nand U6810 (N_6810,N_2710,N_4871);
or U6811 (N_6811,N_3544,N_3650);
nor U6812 (N_6812,N_3142,N_3004);
or U6813 (N_6813,N_3506,N_3189);
or U6814 (N_6814,N_4140,N_3236);
nor U6815 (N_6815,N_2708,N_3238);
and U6816 (N_6816,N_2765,N_3673);
nor U6817 (N_6817,N_4042,N_3352);
nand U6818 (N_6818,N_4431,N_3788);
and U6819 (N_6819,N_3018,N_3109);
and U6820 (N_6820,N_4785,N_4262);
and U6821 (N_6821,N_4048,N_2721);
nand U6822 (N_6822,N_3775,N_3655);
and U6823 (N_6823,N_3391,N_2624);
nand U6824 (N_6824,N_4241,N_3232);
and U6825 (N_6825,N_3466,N_4464);
xor U6826 (N_6826,N_4289,N_4390);
nor U6827 (N_6827,N_4567,N_3520);
nand U6828 (N_6828,N_4667,N_3637);
nand U6829 (N_6829,N_3449,N_3719);
nor U6830 (N_6830,N_4675,N_4767);
nor U6831 (N_6831,N_3510,N_2799);
and U6832 (N_6832,N_3727,N_3439);
or U6833 (N_6833,N_4340,N_4756);
and U6834 (N_6834,N_2711,N_4797);
and U6835 (N_6835,N_2951,N_2569);
or U6836 (N_6836,N_4405,N_4734);
nand U6837 (N_6837,N_2738,N_4696);
and U6838 (N_6838,N_4846,N_3216);
nor U6839 (N_6839,N_4440,N_4884);
xnor U6840 (N_6840,N_3040,N_4942);
or U6841 (N_6841,N_4333,N_2585);
or U6842 (N_6842,N_2778,N_3234);
or U6843 (N_6843,N_4848,N_4405);
or U6844 (N_6844,N_4123,N_4051);
nor U6845 (N_6845,N_4168,N_4554);
or U6846 (N_6846,N_4664,N_4178);
nand U6847 (N_6847,N_3830,N_4097);
nand U6848 (N_6848,N_3521,N_4693);
nand U6849 (N_6849,N_4914,N_4302);
and U6850 (N_6850,N_4757,N_3270);
nand U6851 (N_6851,N_4933,N_3301);
xnor U6852 (N_6852,N_3837,N_2921);
and U6853 (N_6853,N_4284,N_3595);
and U6854 (N_6854,N_4213,N_2600);
or U6855 (N_6855,N_3240,N_3469);
or U6856 (N_6856,N_3342,N_2962);
and U6857 (N_6857,N_3373,N_3260);
nor U6858 (N_6858,N_4003,N_4546);
or U6859 (N_6859,N_4491,N_3486);
nand U6860 (N_6860,N_4317,N_4912);
nand U6861 (N_6861,N_3887,N_4893);
nand U6862 (N_6862,N_4408,N_3268);
and U6863 (N_6863,N_3148,N_4848);
nand U6864 (N_6864,N_3237,N_3189);
nor U6865 (N_6865,N_3332,N_4050);
nand U6866 (N_6866,N_2965,N_2564);
and U6867 (N_6867,N_3950,N_3108);
nor U6868 (N_6868,N_3549,N_3339);
nand U6869 (N_6869,N_4112,N_4614);
nand U6870 (N_6870,N_4700,N_2540);
or U6871 (N_6871,N_4419,N_2916);
or U6872 (N_6872,N_4900,N_3606);
or U6873 (N_6873,N_2997,N_3888);
nand U6874 (N_6874,N_4790,N_4302);
nor U6875 (N_6875,N_4649,N_4393);
xnor U6876 (N_6876,N_4061,N_2741);
or U6877 (N_6877,N_2801,N_4812);
xor U6878 (N_6878,N_2565,N_3779);
nor U6879 (N_6879,N_3966,N_4150);
or U6880 (N_6880,N_3947,N_4783);
nand U6881 (N_6881,N_4151,N_3156);
nor U6882 (N_6882,N_4812,N_4978);
or U6883 (N_6883,N_4291,N_2542);
and U6884 (N_6884,N_3170,N_2665);
nor U6885 (N_6885,N_3388,N_3928);
nand U6886 (N_6886,N_4970,N_4022);
nand U6887 (N_6887,N_4829,N_3334);
and U6888 (N_6888,N_3936,N_4871);
xor U6889 (N_6889,N_4043,N_3544);
or U6890 (N_6890,N_3450,N_3625);
nor U6891 (N_6891,N_4376,N_4763);
nand U6892 (N_6892,N_3505,N_2648);
and U6893 (N_6893,N_3862,N_2697);
nand U6894 (N_6894,N_3911,N_4235);
nor U6895 (N_6895,N_4349,N_4361);
and U6896 (N_6896,N_2919,N_4765);
nor U6897 (N_6897,N_4117,N_4191);
or U6898 (N_6898,N_4054,N_3629);
nand U6899 (N_6899,N_3406,N_2847);
nand U6900 (N_6900,N_3554,N_2503);
and U6901 (N_6901,N_3539,N_3857);
nand U6902 (N_6902,N_3670,N_3470);
nand U6903 (N_6903,N_2514,N_3927);
nand U6904 (N_6904,N_3372,N_3333);
or U6905 (N_6905,N_3905,N_4762);
nand U6906 (N_6906,N_4813,N_4279);
xor U6907 (N_6907,N_3883,N_2588);
or U6908 (N_6908,N_2912,N_4758);
nand U6909 (N_6909,N_3856,N_4408);
or U6910 (N_6910,N_4910,N_3183);
nor U6911 (N_6911,N_2558,N_4244);
or U6912 (N_6912,N_4835,N_2927);
xnor U6913 (N_6913,N_4119,N_3315);
and U6914 (N_6914,N_3656,N_3735);
nand U6915 (N_6915,N_4350,N_4579);
nor U6916 (N_6916,N_4951,N_3993);
and U6917 (N_6917,N_4671,N_4882);
or U6918 (N_6918,N_4358,N_4233);
and U6919 (N_6919,N_3158,N_3665);
xor U6920 (N_6920,N_4633,N_3839);
xnor U6921 (N_6921,N_4565,N_4038);
nor U6922 (N_6922,N_4136,N_2693);
nor U6923 (N_6923,N_2580,N_4484);
nand U6924 (N_6924,N_4512,N_2582);
or U6925 (N_6925,N_3122,N_3313);
xor U6926 (N_6926,N_4286,N_3143);
or U6927 (N_6927,N_3019,N_4664);
xor U6928 (N_6928,N_3968,N_2682);
nor U6929 (N_6929,N_3318,N_3329);
nor U6930 (N_6930,N_4867,N_4989);
or U6931 (N_6931,N_2510,N_4123);
nor U6932 (N_6932,N_3433,N_2856);
or U6933 (N_6933,N_4853,N_3359);
or U6934 (N_6934,N_3844,N_4656);
and U6935 (N_6935,N_3530,N_3656);
or U6936 (N_6936,N_2597,N_2759);
nor U6937 (N_6937,N_4323,N_3672);
nand U6938 (N_6938,N_4027,N_3455);
and U6939 (N_6939,N_4563,N_3841);
nor U6940 (N_6940,N_3854,N_3832);
nor U6941 (N_6941,N_2759,N_3673);
nor U6942 (N_6942,N_4629,N_4812);
and U6943 (N_6943,N_2657,N_4509);
and U6944 (N_6944,N_4213,N_4012);
nor U6945 (N_6945,N_4424,N_2590);
nand U6946 (N_6946,N_2679,N_3364);
nand U6947 (N_6947,N_3740,N_3497);
or U6948 (N_6948,N_4262,N_4360);
nor U6949 (N_6949,N_4916,N_2594);
nor U6950 (N_6950,N_2502,N_3463);
nor U6951 (N_6951,N_4730,N_3164);
or U6952 (N_6952,N_3527,N_4326);
or U6953 (N_6953,N_3534,N_3936);
nor U6954 (N_6954,N_3094,N_3284);
and U6955 (N_6955,N_4760,N_4578);
or U6956 (N_6956,N_3953,N_3587);
nand U6957 (N_6957,N_3341,N_4479);
or U6958 (N_6958,N_4689,N_4861);
and U6959 (N_6959,N_4114,N_3701);
nor U6960 (N_6960,N_4290,N_2705);
or U6961 (N_6961,N_4425,N_2930);
nor U6962 (N_6962,N_2689,N_3078);
or U6963 (N_6963,N_4376,N_3870);
and U6964 (N_6964,N_2950,N_4035);
xor U6965 (N_6965,N_4267,N_2915);
or U6966 (N_6966,N_4267,N_3178);
nand U6967 (N_6967,N_3550,N_4207);
nor U6968 (N_6968,N_4799,N_3619);
or U6969 (N_6969,N_2917,N_4187);
xor U6970 (N_6970,N_3567,N_2864);
nand U6971 (N_6971,N_2861,N_4026);
nor U6972 (N_6972,N_3324,N_2503);
nor U6973 (N_6973,N_2626,N_2932);
nor U6974 (N_6974,N_4447,N_4378);
nand U6975 (N_6975,N_3396,N_3859);
and U6976 (N_6976,N_3574,N_4911);
nand U6977 (N_6977,N_2592,N_4022);
or U6978 (N_6978,N_3372,N_3195);
nand U6979 (N_6979,N_2934,N_3414);
or U6980 (N_6980,N_3208,N_4541);
and U6981 (N_6981,N_4306,N_4589);
or U6982 (N_6982,N_4139,N_4043);
nand U6983 (N_6983,N_2975,N_3659);
nand U6984 (N_6984,N_4714,N_3420);
nor U6985 (N_6985,N_4037,N_4337);
nand U6986 (N_6986,N_4932,N_4586);
nor U6987 (N_6987,N_4861,N_2543);
nor U6988 (N_6988,N_4566,N_3548);
or U6989 (N_6989,N_3876,N_3993);
or U6990 (N_6990,N_3269,N_3543);
nor U6991 (N_6991,N_3584,N_4187);
nor U6992 (N_6992,N_4469,N_4154);
or U6993 (N_6993,N_4833,N_3906);
nor U6994 (N_6994,N_4106,N_2637);
xnor U6995 (N_6995,N_2972,N_3256);
nor U6996 (N_6996,N_4070,N_2684);
nor U6997 (N_6997,N_4202,N_3687);
or U6998 (N_6998,N_3773,N_4502);
xnor U6999 (N_6999,N_3353,N_3482);
and U7000 (N_7000,N_3345,N_4057);
nand U7001 (N_7001,N_3065,N_4632);
nand U7002 (N_7002,N_3771,N_3843);
xnor U7003 (N_7003,N_4539,N_4318);
nor U7004 (N_7004,N_4221,N_4467);
or U7005 (N_7005,N_2869,N_4587);
or U7006 (N_7006,N_3598,N_4790);
or U7007 (N_7007,N_3304,N_2986);
nor U7008 (N_7008,N_4247,N_4425);
or U7009 (N_7009,N_4807,N_3765);
nor U7010 (N_7010,N_3033,N_2715);
and U7011 (N_7011,N_3902,N_2691);
nand U7012 (N_7012,N_2652,N_3287);
and U7013 (N_7013,N_2508,N_4605);
nand U7014 (N_7014,N_2866,N_3106);
xnor U7015 (N_7015,N_2997,N_2500);
and U7016 (N_7016,N_4697,N_3575);
nor U7017 (N_7017,N_4310,N_4576);
xnor U7018 (N_7018,N_3098,N_3496);
or U7019 (N_7019,N_4447,N_3190);
and U7020 (N_7020,N_4261,N_2866);
and U7021 (N_7021,N_2992,N_2790);
nor U7022 (N_7022,N_4079,N_2547);
and U7023 (N_7023,N_3656,N_3577);
or U7024 (N_7024,N_2525,N_2786);
or U7025 (N_7025,N_4416,N_4859);
nor U7026 (N_7026,N_3115,N_4505);
or U7027 (N_7027,N_3382,N_2687);
or U7028 (N_7028,N_4715,N_3645);
or U7029 (N_7029,N_4230,N_2794);
and U7030 (N_7030,N_4855,N_3989);
and U7031 (N_7031,N_3178,N_3375);
nand U7032 (N_7032,N_4011,N_4130);
nand U7033 (N_7033,N_2572,N_4290);
or U7034 (N_7034,N_3806,N_4046);
and U7035 (N_7035,N_3652,N_4499);
and U7036 (N_7036,N_4008,N_3023);
and U7037 (N_7037,N_3127,N_4777);
or U7038 (N_7038,N_2866,N_4455);
nor U7039 (N_7039,N_3588,N_3884);
xor U7040 (N_7040,N_3426,N_3790);
nand U7041 (N_7041,N_2572,N_4562);
nor U7042 (N_7042,N_4182,N_3600);
or U7043 (N_7043,N_2883,N_4318);
nor U7044 (N_7044,N_2504,N_4950);
or U7045 (N_7045,N_4710,N_3664);
nor U7046 (N_7046,N_3862,N_4128);
and U7047 (N_7047,N_4160,N_2516);
or U7048 (N_7048,N_3659,N_3933);
and U7049 (N_7049,N_2734,N_2943);
nand U7050 (N_7050,N_3927,N_3110);
nand U7051 (N_7051,N_2555,N_2711);
and U7052 (N_7052,N_3810,N_4990);
or U7053 (N_7053,N_3883,N_4237);
or U7054 (N_7054,N_3940,N_4275);
and U7055 (N_7055,N_3930,N_3092);
and U7056 (N_7056,N_3042,N_3887);
or U7057 (N_7057,N_3777,N_3279);
nand U7058 (N_7058,N_3586,N_4217);
or U7059 (N_7059,N_3882,N_3556);
nand U7060 (N_7060,N_3847,N_3201);
nand U7061 (N_7061,N_2717,N_4190);
and U7062 (N_7062,N_2741,N_3817);
nand U7063 (N_7063,N_4586,N_3420);
nor U7064 (N_7064,N_3012,N_4257);
xnor U7065 (N_7065,N_2756,N_4165);
and U7066 (N_7066,N_3128,N_4986);
nand U7067 (N_7067,N_3923,N_4212);
or U7068 (N_7068,N_3110,N_3087);
nand U7069 (N_7069,N_4422,N_2597);
or U7070 (N_7070,N_2880,N_4894);
and U7071 (N_7071,N_3612,N_2641);
and U7072 (N_7072,N_4990,N_4471);
nor U7073 (N_7073,N_4518,N_2581);
xor U7074 (N_7074,N_3863,N_3343);
nand U7075 (N_7075,N_4034,N_4690);
and U7076 (N_7076,N_2913,N_2926);
and U7077 (N_7077,N_4919,N_4230);
or U7078 (N_7078,N_3542,N_3880);
or U7079 (N_7079,N_4374,N_2623);
and U7080 (N_7080,N_4480,N_4308);
and U7081 (N_7081,N_3263,N_3980);
and U7082 (N_7082,N_3826,N_2799);
and U7083 (N_7083,N_2965,N_3998);
nor U7084 (N_7084,N_4251,N_3617);
xor U7085 (N_7085,N_2851,N_4843);
and U7086 (N_7086,N_3990,N_3594);
or U7087 (N_7087,N_4834,N_4871);
and U7088 (N_7088,N_4089,N_4651);
and U7089 (N_7089,N_3284,N_4979);
nor U7090 (N_7090,N_2716,N_4443);
nand U7091 (N_7091,N_2644,N_3648);
and U7092 (N_7092,N_3108,N_3593);
and U7093 (N_7093,N_4715,N_3131);
or U7094 (N_7094,N_4969,N_2779);
and U7095 (N_7095,N_4011,N_4586);
xnor U7096 (N_7096,N_4182,N_2889);
xnor U7097 (N_7097,N_2929,N_4794);
and U7098 (N_7098,N_3779,N_4999);
and U7099 (N_7099,N_2544,N_4594);
or U7100 (N_7100,N_3176,N_2605);
nor U7101 (N_7101,N_2768,N_2652);
or U7102 (N_7102,N_2778,N_4895);
or U7103 (N_7103,N_3040,N_4241);
or U7104 (N_7104,N_4655,N_3010);
nand U7105 (N_7105,N_2962,N_3944);
or U7106 (N_7106,N_3690,N_4434);
or U7107 (N_7107,N_3468,N_4559);
or U7108 (N_7108,N_4259,N_2534);
nand U7109 (N_7109,N_3534,N_2727);
nand U7110 (N_7110,N_2589,N_4089);
nand U7111 (N_7111,N_4454,N_2616);
nand U7112 (N_7112,N_3802,N_3011);
nor U7113 (N_7113,N_4600,N_4508);
nor U7114 (N_7114,N_3361,N_2581);
nor U7115 (N_7115,N_2927,N_4858);
or U7116 (N_7116,N_2896,N_3060);
nand U7117 (N_7117,N_4750,N_2851);
and U7118 (N_7118,N_3797,N_2542);
and U7119 (N_7119,N_3357,N_4870);
and U7120 (N_7120,N_4274,N_3657);
nor U7121 (N_7121,N_3879,N_2766);
nor U7122 (N_7122,N_3476,N_3668);
or U7123 (N_7123,N_3746,N_3840);
xor U7124 (N_7124,N_4308,N_3329);
nand U7125 (N_7125,N_4651,N_4047);
and U7126 (N_7126,N_4914,N_2952);
and U7127 (N_7127,N_3081,N_4854);
nor U7128 (N_7128,N_4697,N_2930);
xnor U7129 (N_7129,N_3274,N_2617);
or U7130 (N_7130,N_2816,N_3242);
and U7131 (N_7131,N_3066,N_2524);
or U7132 (N_7132,N_4439,N_3112);
xor U7133 (N_7133,N_2949,N_3230);
nor U7134 (N_7134,N_3820,N_2716);
and U7135 (N_7135,N_3497,N_2554);
nor U7136 (N_7136,N_2633,N_3473);
nor U7137 (N_7137,N_3834,N_3842);
nor U7138 (N_7138,N_4204,N_3356);
or U7139 (N_7139,N_2598,N_3997);
or U7140 (N_7140,N_4124,N_3949);
nand U7141 (N_7141,N_4167,N_3848);
nor U7142 (N_7142,N_4394,N_3524);
and U7143 (N_7143,N_4326,N_4319);
or U7144 (N_7144,N_2894,N_3263);
nor U7145 (N_7145,N_3707,N_4416);
xor U7146 (N_7146,N_3306,N_3355);
or U7147 (N_7147,N_4929,N_3912);
or U7148 (N_7148,N_4621,N_4336);
and U7149 (N_7149,N_3359,N_2950);
nor U7150 (N_7150,N_4838,N_3010);
and U7151 (N_7151,N_3663,N_3262);
nor U7152 (N_7152,N_2805,N_2847);
xor U7153 (N_7153,N_3656,N_3376);
nor U7154 (N_7154,N_2697,N_4748);
or U7155 (N_7155,N_2911,N_4572);
nand U7156 (N_7156,N_4058,N_3849);
and U7157 (N_7157,N_3662,N_4408);
or U7158 (N_7158,N_2964,N_2734);
nand U7159 (N_7159,N_3137,N_2736);
nor U7160 (N_7160,N_3017,N_4820);
xor U7161 (N_7161,N_3180,N_4662);
nor U7162 (N_7162,N_2863,N_4432);
nand U7163 (N_7163,N_3206,N_2600);
and U7164 (N_7164,N_4629,N_3071);
xnor U7165 (N_7165,N_3008,N_4323);
and U7166 (N_7166,N_3670,N_2974);
or U7167 (N_7167,N_3167,N_4326);
or U7168 (N_7168,N_3866,N_4599);
and U7169 (N_7169,N_4240,N_4796);
nor U7170 (N_7170,N_4431,N_3938);
nand U7171 (N_7171,N_2562,N_3991);
xnor U7172 (N_7172,N_4437,N_3880);
or U7173 (N_7173,N_3791,N_3795);
nand U7174 (N_7174,N_4492,N_2896);
nor U7175 (N_7175,N_4880,N_4184);
nand U7176 (N_7176,N_4060,N_4606);
or U7177 (N_7177,N_4578,N_4157);
nand U7178 (N_7178,N_3504,N_2813);
nand U7179 (N_7179,N_3826,N_3125);
or U7180 (N_7180,N_3297,N_2506);
nand U7181 (N_7181,N_4273,N_3923);
nand U7182 (N_7182,N_4348,N_4985);
nor U7183 (N_7183,N_3413,N_4435);
xnor U7184 (N_7184,N_3578,N_4698);
and U7185 (N_7185,N_4056,N_2857);
or U7186 (N_7186,N_3789,N_4018);
nor U7187 (N_7187,N_4989,N_4695);
or U7188 (N_7188,N_3820,N_4794);
xor U7189 (N_7189,N_4783,N_3892);
nor U7190 (N_7190,N_4478,N_4474);
nand U7191 (N_7191,N_2617,N_2621);
nand U7192 (N_7192,N_3778,N_4599);
and U7193 (N_7193,N_4224,N_3900);
nand U7194 (N_7194,N_4820,N_3324);
nor U7195 (N_7195,N_3750,N_3743);
and U7196 (N_7196,N_4515,N_4909);
and U7197 (N_7197,N_4442,N_4071);
and U7198 (N_7198,N_4496,N_4724);
nand U7199 (N_7199,N_2715,N_3734);
nor U7200 (N_7200,N_4822,N_3104);
or U7201 (N_7201,N_3006,N_4681);
nand U7202 (N_7202,N_3438,N_4182);
and U7203 (N_7203,N_4981,N_4365);
nor U7204 (N_7204,N_4619,N_4008);
or U7205 (N_7205,N_4083,N_4857);
or U7206 (N_7206,N_2887,N_3988);
or U7207 (N_7207,N_3598,N_2618);
nand U7208 (N_7208,N_3426,N_2663);
or U7209 (N_7209,N_4238,N_3632);
and U7210 (N_7210,N_4002,N_2578);
xnor U7211 (N_7211,N_3270,N_4135);
or U7212 (N_7212,N_4647,N_4833);
xor U7213 (N_7213,N_4836,N_3262);
nand U7214 (N_7214,N_4049,N_4573);
nand U7215 (N_7215,N_4636,N_2543);
and U7216 (N_7216,N_2748,N_3073);
or U7217 (N_7217,N_4971,N_4302);
and U7218 (N_7218,N_4750,N_3681);
and U7219 (N_7219,N_2692,N_3692);
or U7220 (N_7220,N_2699,N_3859);
and U7221 (N_7221,N_3688,N_3385);
or U7222 (N_7222,N_4280,N_3138);
or U7223 (N_7223,N_4878,N_4451);
or U7224 (N_7224,N_4726,N_3049);
and U7225 (N_7225,N_2984,N_3151);
or U7226 (N_7226,N_3302,N_3587);
and U7227 (N_7227,N_4521,N_4227);
and U7228 (N_7228,N_3918,N_4978);
or U7229 (N_7229,N_3847,N_3401);
nand U7230 (N_7230,N_4868,N_4207);
or U7231 (N_7231,N_3133,N_3151);
xnor U7232 (N_7232,N_4306,N_4449);
or U7233 (N_7233,N_4293,N_3600);
and U7234 (N_7234,N_4555,N_2579);
or U7235 (N_7235,N_2892,N_2595);
and U7236 (N_7236,N_3906,N_4855);
nand U7237 (N_7237,N_3932,N_4287);
and U7238 (N_7238,N_3838,N_3462);
and U7239 (N_7239,N_3142,N_4955);
nor U7240 (N_7240,N_3146,N_4275);
and U7241 (N_7241,N_2924,N_4584);
nand U7242 (N_7242,N_3886,N_2815);
nand U7243 (N_7243,N_4170,N_3578);
and U7244 (N_7244,N_2791,N_3902);
nor U7245 (N_7245,N_2975,N_2614);
nor U7246 (N_7246,N_3652,N_4451);
nor U7247 (N_7247,N_4679,N_3803);
or U7248 (N_7248,N_3673,N_3684);
and U7249 (N_7249,N_3945,N_3140);
and U7250 (N_7250,N_3732,N_3751);
and U7251 (N_7251,N_3377,N_3852);
nand U7252 (N_7252,N_3362,N_4495);
or U7253 (N_7253,N_2896,N_2718);
and U7254 (N_7254,N_3484,N_4723);
and U7255 (N_7255,N_3984,N_3609);
nor U7256 (N_7256,N_3818,N_3283);
nand U7257 (N_7257,N_2591,N_3821);
nor U7258 (N_7258,N_4306,N_4335);
and U7259 (N_7259,N_2886,N_2550);
nor U7260 (N_7260,N_4246,N_4988);
and U7261 (N_7261,N_4110,N_2602);
nand U7262 (N_7262,N_2655,N_4833);
or U7263 (N_7263,N_2551,N_4788);
or U7264 (N_7264,N_3883,N_3799);
and U7265 (N_7265,N_3957,N_3398);
nor U7266 (N_7266,N_3367,N_3018);
or U7267 (N_7267,N_4330,N_3686);
xor U7268 (N_7268,N_2800,N_2876);
and U7269 (N_7269,N_2920,N_4600);
nor U7270 (N_7270,N_2711,N_4545);
nor U7271 (N_7271,N_4590,N_3786);
nand U7272 (N_7272,N_4809,N_3498);
nand U7273 (N_7273,N_4863,N_3082);
nand U7274 (N_7274,N_4225,N_3665);
and U7275 (N_7275,N_3302,N_2513);
nor U7276 (N_7276,N_4811,N_3800);
nand U7277 (N_7277,N_4636,N_3657);
nor U7278 (N_7278,N_3235,N_4817);
and U7279 (N_7279,N_3616,N_4831);
nor U7280 (N_7280,N_4446,N_4126);
nor U7281 (N_7281,N_3352,N_3462);
nor U7282 (N_7282,N_4984,N_4560);
and U7283 (N_7283,N_3789,N_4528);
nor U7284 (N_7284,N_3440,N_4411);
xor U7285 (N_7285,N_4404,N_4318);
or U7286 (N_7286,N_2583,N_3783);
or U7287 (N_7287,N_4447,N_3437);
nor U7288 (N_7288,N_3033,N_3785);
nor U7289 (N_7289,N_3864,N_4577);
xor U7290 (N_7290,N_4396,N_4980);
or U7291 (N_7291,N_3106,N_3126);
or U7292 (N_7292,N_2862,N_4337);
or U7293 (N_7293,N_3694,N_2890);
xor U7294 (N_7294,N_4762,N_3745);
and U7295 (N_7295,N_2998,N_3609);
and U7296 (N_7296,N_3940,N_3363);
nand U7297 (N_7297,N_4443,N_3024);
nand U7298 (N_7298,N_4704,N_4519);
nand U7299 (N_7299,N_4088,N_4878);
nand U7300 (N_7300,N_4587,N_4768);
or U7301 (N_7301,N_2629,N_4884);
or U7302 (N_7302,N_3613,N_4426);
or U7303 (N_7303,N_3781,N_2769);
nand U7304 (N_7304,N_2628,N_4358);
nor U7305 (N_7305,N_3455,N_4313);
nor U7306 (N_7306,N_3180,N_4963);
nor U7307 (N_7307,N_4625,N_4679);
nor U7308 (N_7308,N_2701,N_4595);
or U7309 (N_7309,N_3253,N_3488);
or U7310 (N_7310,N_2683,N_2621);
and U7311 (N_7311,N_3527,N_4643);
xor U7312 (N_7312,N_2941,N_3579);
or U7313 (N_7313,N_4055,N_4738);
nand U7314 (N_7314,N_4530,N_4171);
and U7315 (N_7315,N_3538,N_2871);
nand U7316 (N_7316,N_2746,N_3459);
nand U7317 (N_7317,N_3896,N_3773);
and U7318 (N_7318,N_4921,N_4402);
or U7319 (N_7319,N_2936,N_4474);
and U7320 (N_7320,N_2744,N_3700);
or U7321 (N_7321,N_4505,N_4980);
and U7322 (N_7322,N_3751,N_4456);
or U7323 (N_7323,N_4258,N_4407);
nor U7324 (N_7324,N_3578,N_3744);
nor U7325 (N_7325,N_4836,N_4258);
and U7326 (N_7326,N_2622,N_4073);
or U7327 (N_7327,N_4429,N_2742);
and U7328 (N_7328,N_4059,N_3138);
xor U7329 (N_7329,N_4353,N_3685);
xnor U7330 (N_7330,N_3571,N_3692);
nor U7331 (N_7331,N_3222,N_3554);
and U7332 (N_7332,N_4829,N_4381);
or U7333 (N_7333,N_4024,N_3160);
nor U7334 (N_7334,N_4116,N_3754);
and U7335 (N_7335,N_3778,N_4780);
nor U7336 (N_7336,N_3892,N_4004);
nor U7337 (N_7337,N_4761,N_3394);
nand U7338 (N_7338,N_4636,N_3105);
and U7339 (N_7339,N_3618,N_4303);
and U7340 (N_7340,N_3663,N_4290);
nand U7341 (N_7341,N_4944,N_3423);
xor U7342 (N_7342,N_4902,N_3667);
nor U7343 (N_7343,N_2646,N_3899);
and U7344 (N_7344,N_3657,N_3226);
nand U7345 (N_7345,N_3621,N_4932);
nand U7346 (N_7346,N_3937,N_2725);
and U7347 (N_7347,N_4785,N_3281);
nor U7348 (N_7348,N_4513,N_4854);
nand U7349 (N_7349,N_4923,N_2541);
nand U7350 (N_7350,N_3246,N_4836);
nor U7351 (N_7351,N_4244,N_4423);
and U7352 (N_7352,N_3514,N_3218);
and U7353 (N_7353,N_4191,N_3588);
xor U7354 (N_7354,N_3036,N_4369);
or U7355 (N_7355,N_4684,N_3576);
or U7356 (N_7356,N_3717,N_4030);
nor U7357 (N_7357,N_3691,N_3687);
nor U7358 (N_7358,N_4901,N_3122);
and U7359 (N_7359,N_3046,N_3708);
xnor U7360 (N_7360,N_4228,N_4317);
and U7361 (N_7361,N_4517,N_3640);
and U7362 (N_7362,N_4981,N_4499);
nand U7363 (N_7363,N_3752,N_4616);
or U7364 (N_7364,N_2965,N_2663);
and U7365 (N_7365,N_4360,N_2914);
and U7366 (N_7366,N_4448,N_2546);
and U7367 (N_7367,N_3610,N_4946);
nand U7368 (N_7368,N_4981,N_4412);
or U7369 (N_7369,N_2764,N_3938);
and U7370 (N_7370,N_2546,N_4347);
nand U7371 (N_7371,N_3845,N_4422);
xnor U7372 (N_7372,N_4219,N_2617);
nor U7373 (N_7373,N_4133,N_4942);
xor U7374 (N_7374,N_2690,N_4628);
or U7375 (N_7375,N_3422,N_4701);
nor U7376 (N_7376,N_2512,N_3139);
nor U7377 (N_7377,N_2613,N_3695);
nand U7378 (N_7378,N_4311,N_4511);
nand U7379 (N_7379,N_3849,N_3093);
nand U7380 (N_7380,N_4503,N_2543);
nor U7381 (N_7381,N_4260,N_4934);
nand U7382 (N_7382,N_4709,N_3951);
or U7383 (N_7383,N_4739,N_3069);
nor U7384 (N_7384,N_3589,N_2932);
nor U7385 (N_7385,N_4954,N_2858);
nor U7386 (N_7386,N_4047,N_3527);
xnor U7387 (N_7387,N_2563,N_4698);
and U7388 (N_7388,N_3518,N_4589);
nand U7389 (N_7389,N_4047,N_2635);
nand U7390 (N_7390,N_3350,N_3031);
nor U7391 (N_7391,N_3183,N_3394);
xnor U7392 (N_7392,N_3518,N_4498);
and U7393 (N_7393,N_2617,N_4133);
nor U7394 (N_7394,N_3324,N_4617);
nor U7395 (N_7395,N_3716,N_3970);
and U7396 (N_7396,N_3849,N_3347);
or U7397 (N_7397,N_4931,N_4611);
nor U7398 (N_7398,N_4719,N_3094);
or U7399 (N_7399,N_4817,N_3352);
nand U7400 (N_7400,N_4706,N_4218);
nor U7401 (N_7401,N_4495,N_4314);
or U7402 (N_7402,N_2897,N_3150);
xnor U7403 (N_7403,N_4334,N_4541);
nand U7404 (N_7404,N_2865,N_3223);
nand U7405 (N_7405,N_3097,N_3229);
and U7406 (N_7406,N_4897,N_3072);
nand U7407 (N_7407,N_3720,N_3242);
nor U7408 (N_7408,N_3124,N_4136);
nor U7409 (N_7409,N_2727,N_3827);
nor U7410 (N_7410,N_3300,N_4052);
or U7411 (N_7411,N_4929,N_3249);
or U7412 (N_7412,N_3469,N_3269);
and U7413 (N_7413,N_2965,N_2751);
or U7414 (N_7414,N_3626,N_2780);
and U7415 (N_7415,N_2753,N_3602);
nand U7416 (N_7416,N_3556,N_4738);
and U7417 (N_7417,N_4170,N_4321);
or U7418 (N_7418,N_3430,N_4416);
nor U7419 (N_7419,N_2515,N_3447);
xor U7420 (N_7420,N_4124,N_2906);
nand U7421 (N_7421,N_4686,N_4885);
and U7422 (N_7422,N_4184,N_3811);
and U7423 (N_7423,N_4460,N_3502);
and U7424 (N_7424,N_4555,N_4482);
and U7425 (N_7425,N_2868,N_4379);
or U7426 (N_7426,N_3216,N_3413);
or U7427 (N_7427,N_3267,N_3462);
or U7428 (N_7428,N_3432,N_4410);
or U7429 (N_7429,N_4444,N_4407);
or U7430 (N_7430,N_4837,N_4581);
nor U7431 (N_7431,N_3340,N_2503);
nor U7432 (N_7432,N_3281,N_3395);
nor U7433 (N_7433,N_2963,N_4430);
or U7434 (N_7434,N_4675,N_3475);
or U7435 (N_7435,N_4851,N_3667);
xnor U7436 (N_7436,N_4892,N_4236);
nor U7437 (N_7437,N_2861,N_3385);
or U7438 (N_7438,N_3249,N_3799);
nand U7439 (N_7439,N_4080,N_3492);
xnor U7440 (N_7440,N_2865,N_3274);
and U7441 (N_7441,N_3538,N_2661);
nand U7442 (N_7442,N_3857,N_3344);
nand U7443 (N_7443,N_3369,N_4267);
or U7444 (N_7444,N_3956,N_3884);
or U7445 (N_7445,N_2979,N_3901);
nand U7446 (N_7446,N_3935,N_3481);
xor U7447 (N_7447,N_3987,N_4651);
nor U7448 (N_7448,N_2569,N_3195);
nand U7449 (N_7449,N_3591,N_4113);
xor U7450 (N_7450,N_4953,N_4800);
xnor U7451 (N_7451,N_4746,N_3837);
or U7452 (N_7452,N_4369,N_2791);
nor U7453 (N_7453,N_2753,N_2854);
or U7454 (N_7454,N_3341,N_3964);
or U7455 (N_7455,N_3658,N_4183);
nand U7456 (N_7456,N_4230,N_4286);
nand U7457 (N_7457,N_2654,N_3745);
xor U7458 (N_7458,N_3594,N_3005);
or U7459 (N_7459,N_4280,N_3145);
nand U7460 (N_7460,N_4585,N_4746);
or U7461 (N_7461,N_4173,N_4436);
or U7462 (N_7462,N_4041,N_4723);
nor U7463 (N_7463,N_2823,N_2763);
or U7464 (N_7464,N_4711,N_4197);
or U7465 (N_7465,N_4269,N_4743);
nand U7466 (N_7466,N_3521,N_3057);
nor U7467 (N_7467,N_3120,N_3511);
nand U7468 (N_7468,N_3623,N_3186);
nand U7469 (N_7469,N_4445,N_4398);
nand U7470 (N_7470,N_4905,N_4132);
or U7471 (N_7471,N_3021,N_4932);
or U7472 (N_7472,N_4710,N_3217);
nor U7473 (N_7473,N_3720,N_3227);
xnor U7474 (N_7474,N_3245,N_4934);
nor U7475 (N_7475,N_4635,N_4832);
nand U7476 (N_7476,N_3493,N_3657);
nand U7477 (N_7477,N_3920,N_3353);
xnor U7478 (N_7478,N_3575,N_2576);
and U7479 (N_7479,N_3974,N_2909);
nand U7480 (N_7480,N_3950,N_2765);
nand U7481 (N_7481,N_2847,N_4854);
nor U7482 (N_7482,N_2613,N_3676);
nand U7483 (N_7483,N_3317,N_2900);
nor U7484 (N_7484,N_4799,N_3743);
xor U7485 (N_7485,N_3863,N_3446);
nand U7486 (N_7486,N_4662,N_3797);
nand U7487 (N_7487,N_4112,N_3506);
or U7488 (N_7488,N_3867,N_4165);
nor U7489 (N_7489,N_3918,N_3561);
nor U7490 (N_7490,N_4694,N_3427);
nand U7491 (N_7491,N_2623,N_2922);
nand U7492 (N_7492,N_3551,N_2974);
nand U7493 (N_7493,N_3335,N_4997);
or U7494 (N_7494,N_3811,N_3192);
and U7495 (N_7495,N_4253,N_4872);
nand U7496 (N_7496,N_3609,N_3783);
and U7497 (N_7497,N_3162,N_4736);
nand U7498 (N_7498,N_4927,N_4469);
nand U7499 (N_7499,N_3145,N_4948);
and U7500 (N_7500,N_7365,N_5933);
nand U7501 (N_7501,N_6552,N_7007);
nor U7502 (N_7502,N_6204,N_6818);
and U7503 (N_7503,N_6613,N_7164);
nand U7504 (N_7504,N_6437,N_7122);
and U7505 (N_7505,N_5244,N_7278);
and U7506 (N_7506,N_5109,N_5205);
nand U7507 (N_7507,N_7429,N_5118);
or U7508 (N_7508,N_5092,N_5782);
and U7509 (N_7509,N_5268,N_6207);
nand U7510 (N_7510,N_7125,N_5369);
and U7511 (N_7511,N_6206,N_5880);
or U7512 (N_7512,N_6029,N_7126);
and U7513 (N_7513,N_7499,N_7115);
nand U7514 (N_7514,N_6002,N_6975);
nor U7515 (N_7515,N_6122,N_5073);
nor U7516 (N_7516,N_6268,N_6234);
and U7517 (N_7517,N_5129,N_6737);
and U7518 (N_7518,N_6454,N_7079);
nor U7519 (N_7519,N_7140,N_5425);
nand U7520 (N_7520,N_6535,N_5280);
nand U7521 (N_7521,N_5327,N_7009);
nor U7522 (N_7522,N_6840,N_5962);
or U7523 (N_7523,N_6428,N_5547);
xor U7524 (N_7524,N_5945,N_6313);
and U7525 (N_7525,N_6369,N_6302);
nand U7526 (N_7526,N_5502,N_5778);
nand U7527 (N_7527,N_5054,N_7432);
xor U7528 (N_7528,N_6800,N_7151);
nand U7529 (N_7529,N_5628,N_7333);
nand U7530 (N_7530,N_5605,N_7399);
nor U7531 (N_7531,N_6291,N_5768);
xnor U7532 (N_7532,N_5656,N_6203);
nand U7533 (N_7533,N_5952,N_5906);
or U7534 (N_7534,N_6598,N_6601);
nand U7535 (N_7535,N_5214,N_7442);
and U7536 (N_7536,N_5598,N_6399);
nor U7537 (N_7537,N_7202,N_5913);
or U7538 (N_7538,N_7014,N_5686);
nor U7539 (N_7539,N_5183,N_5811);
nor U7540 (N_7540,N_5653,N_7242);
and U7541 (N_7541,N_5055,N_5433);
nor U7542 (N_7542,N_6509,N_5397);
nor U7543 (N_7543,N_6823,N_5245);
nor U7544 (N_7544,N_5527,N_5114);
and U7545 (N_7545,N_6325,N_6726);
nor U7546 (N_7546,N_6030,N_6735);
and U7547 (N_7547,N_6844,N_6046);
or U7548 (N_7548,N_6086,N_5878);
xnor U7549 (N_7549,N_5080,N_6950);
nor U7550 (N_7550,N_7401,N_7434);
and U7551 (N_7551,N_6470,N_7404);
or U7552 (N_7552,N_6690,N_5204);
and U7553 (N_7553,N_5248,N_7400);
nand U7554 (N_7554,N_5925,N_6721);
or U7555 (N_7555,N_7344,N_6825);
nand U7556 (N_7556,N_6792,N_5446);
nor U7557 (N_7557,N_7327,N_6553);
or U7558 (N_7558,N_6315,N_5478);
or U7559 (N_7559,N_5134,N_6247);
or U7560 (N_7560,N_5780,N_5312);
and U7561 (N_7561,N_7004,N_6281);
and U7562 (N_7562,N_6216,N_7392);
nor U7563 (N_7563,N_6843,N_6926);
and U7564 (N_7564,N_6557,N_6431);
and U7565 (N_7565,N_6150,N_6117);
xnor U7566 (N_7566,N_7003,N_6514);
or U7567 (N_7567,N_6661,N_6245);
nand U7568 (N_7568,N_7339,N_6044);
nor U7569 (N_7569,N_5013,N_6688);
and U7570 (N_7570,N_5383,N_6426);
nor U7571 (N_7571,N_6838,N_5039);
or U7572 (N_7572,N_7065,N_6039);
nor U7573 (N_7573,N_6169,N_5572);
and U7574 (N_7574,N_5717,N_6516);
or U7575 (N_7575,N_5824,N_5172);
and U7576 (N_7576,N_7116,N_5938);
or U7577 (N_7577,N_7270,N_7256);
nor U7578 (N_7578,N_6615,N_6013);
nor U7579 (N_7579,N_7388,N_7258);
nor U7580 (N_7580,N_6263,N_5899);
xor U7581 (N_7581,N_5164,N_5875);
or U7582 (N_7582,N_6213,N_5870);
nand U7583 (N_7583,N_6802,N_5489);
nor U7584 (N_7584,N_6362,N_5479);
and U7585 (N_7585,N_7483,N_7194);
and U7586 (N_7586,N_6765,N_6682);
and U7587 (N_7587,N_5901,N_6376);
nand U7588 (N_7588,N_6318,N_6253);
xnor U7589 (N_7589,N_6812,N_6907);
or U7590 (N_7590,N_6215,N_6532);
nor U7591 (N_7591,N_6005,N_5390);
nand U7592 (N_7592,N_5001,N_5398);
nor U7593 (N_7593,N_5530,N_6074);
nand U7594 (N_7594,N_6968,N_5708);
and U7595 (N_7595,N_5148,N_6816);
or U7596 (N_7596,N_7480,N_6444);
nand U7597 (N_7597,N_6242,N_6421);
and U7598 (N_7598,N_5087,N_7058);
or U7599 (N_7599,N_6286,N_5872);
or U7600 (N_7600,N_7317,N_5517);
xor U7601 (N_7601,N_6036,N_5744);
and U7602 (N_7602,N_5061,N_7135);
nand U7603 (N_7603,N_6712,N_7496);
xnor U7604 (N_7604,N_5677,N_6109);
xor U7605 (N_7605,N_6507,N_7201);
and U7606 (N_7606,N_5184,N_6893);
or U7607 (N_7607,N_7376,N_6579);
nor U7608 (N_7608,N_7269,N_5252);
and U7609 (N_7609,N_6224,N_5888);
xor U7610 (N_7610,N_7448,N_7186);
nand U7611 (N_7611,N_5596,N_7109);
or U7612 (N_7612,N_7280,N_6389);
and U7613 (N_7613,N_6231,N_6547);
and U7614 (N_7614,N_6282,N_6577);
nor U7615 (N_7615,N_5178,N_6487);
and U7616 (N_7616,N_5570,N_6011);
and U7617 (N_7617,N_5706,N_7359);
or U7618 (N_7618,N_5269,N_5541);
or U7619 (N_7619,N_7019,N_5625);
nand U7620 (N_7620,N_7106,N_5958);
nand U7621 (N_7621,N_5841,N_6715);
or U7622 (N_7622,N_5429,N_5325);
nand U7623 (N_7623,N_5917,N_5518);
nor U7624 (N_7624,N_7132,N_5132);
nor U7625 (N_7625,N_6931,N_5549);
nand U7626 (N_7626,N_6987,N_5281);
nor U7627 (N_7627,N_5259,N_7431);
and U7628 (N_7628,N_5593,N_5033);
nor U7629 (N_7629,N_5051,N_7463);
nand U7630 (N_7630,N_6772,N_5275);
nand U7631 (N_7631,N_6149,N_5698);
or U7632 (N_7632,N_5186,N_5045);
nor U7633 (N_7633,N_5975,N_5759);
or U7634 (N_7634,N_5763,N_6955);
or U7635 (N_7635,N_6602,N_5781);
nor U7636 (N_7636,N_6774,N_5128);
nor U7637 (N_7637,N_6728,N_5139);
nor U7638 (N_7638,N_6064,N_6394);
nand U7639 (N_7639,N_5602,N_5492);
and U7640 (N_7640,N_7488,N_6422);
and U7641 (N_7641,N_7096,N_6141);
and U7642 (N_7642,N_7435,N_5908);
and U7643 (N_7643,N_7152,N_5816);
xor U7644 (N_7644,N_5828,N_5236);
or U7645 (N_7645,N_6903,N_5652);
xnor U7646 (N_7646,N_6945,N_5179);
nor U7647 (N_7647,N_5820,N_5400);
or U7648 (N_7648,N_5626,N_5904);
nor U7649 (N_7649,N_5600,N_6279);
nor U7650 (N_7650,N_5848,N_5505);
or U7651 (N_7651,N_6189,N_7041);
or U7652 (N_7652,N_5861,N_7255);
or U7653 (N_7653,N_5126,N_5189);
nor U7654 (N_7654,N_6618,N_5322);
nand U7655 (N_7655,N_6533,N_7322);
or U7656 (N_7656,N_7320,N_6947);
and U7657 (N_7657,N_5030,N_5165);
nor U7658 (N_7658,N_5578,N_6808);
nand U7659 (N_7659,N_5443,N_5403);
and U7660 (N_7660,N_7485,N_6841);
nand U7661 (N_7661,N_5480,N_6961);
and U7662 (N_7662,N_6548,N_5002);
nand U7663 (N_7663,N_6071,N_6218);
and U7664 (N_7664,N_7154,N_5557);
or U7665 (N_7665,N_6730,N_5910);
or U7666 (N_7666,N_5347,N_7038);
nand U7667 (N_7667,N_5162,N_6745);
or U7668 (N_7668,N_7010,N_6382);
nor U7669 (N_7669,N_5751,N_5903);
and U7670 (N_7670,N_5599,N_7261);
xnor U7671 (N_7671,N_7063,N_5069);
or U7672 (N_7672,N_5950,N_5218);
or U7673 (N_7673,N_5451,N_7074);
nand U7674 (N_7674,N_5897,N_5997);
and U7675 (N_7675,N_6519,N_5378);
and U7676 (N_7676,N_5113,N_7073);
nor U7677 (N_7677,N_6580,N_5332);
or U7678 (N_7678,N_5972,N_7110);
nor U7679 (N_7679,N_7185,N_7313);
and U7680 (N_7680,N_5770,N_7301);
nor U7681 (N_7681,N_6156,N_5146);
nand U7682 (N_7682,N_6966,N_5743);
nand U7683 (N_7683,N_7217,N_5724);
nand U7684 (N_7684,N_7482,N_6722);
xnor U7685 (N_7685,N_5388,N_5583);
or U7686 (N_7686,N_5298,N_6790);
or U7687 (N_7687,N_5696,N_5589);
or U7688 (N_7688,N_6473,N_5188);
and U7689 (N_7689,N_7390,N_5417);
nor U7690 (N_7690,N_7120,N_6828);
and U7691 (N_7691,N_5854,N_7484);
xor U7692 (N_7692,N_5334,N_5331);
nor U7693 (N_7693,N_6752,N_7205);
nor U7694 (N_7694,N_6095,N_6290);
nand U7695 (N_7695,N_6022,N_5983);
or U7696 (N_7696,N_6283,N_5320);
xor U7697 (N_7697,N_6767,N_7118);
nor U7698 (N_7698,N_6536,N_5984);
nand U7699 (N_7699,N_6352,N_5927);
and U7700 (N_7700,N_6391,N_7229);
and U7701 (N_7701,N_5260,N_6671);
and U7702 (N_7702,N_7143,N_6185);
or U7703 (N_7703,N_7139,N_6214);
or U7704 (N_7704,N_6942,N_6177);
or U7705 (N_7705,N_6517,N_6972);
nand U7706 (N_7706,N_7117,N_6757);
xnor U7707 (N_7707,N_6933,N_5765);
and U7708 (N_7708,N_6639,N_6296);
nand U7709 (N_7709,N_6070,N_6622);
nor U7710 (N_7710,N_5261,N_6104);
nand U7711 (N_7711,N_6641,N_5454);
and U7712 (N_7712,N_5858,N_7450);
and U7713 (N_7713,N_6293,N_6904);
xor U7714 (N_7714,N_5890,N_7002);
xor U7715 (N_7715,N_6403,N_5684);
nand U7716 (N_7716,N_6559,N_5258);
nand U7717 (N_7717,N_5427,N_6385);
and U7718 (N_7718,N_7291,N_6465);
nand U7719 (N_7719,N_7391,N_5660);
or U7720 (N_7720,N_6289,N_5832);
and U7721 (N_7721,N_5104,N_6845);
xnor U7722 (N_7722,N_5771,N_6694);
or U7723 (N_7723,N_5584,N_6978);
and U7724 (N_7724,N_6549,N_5201);
nor U7725 (N_7725,N_6928,N_5376);
nor U7726 (N_7726,N_5728,N_6298);
and U7727 (N_7727,N_5253,N_5629);
or U7728 (N_7728,N_5267,N_6355);
nand U7729 (N_7729,N_6175,N_5086);
nor U7730 (N_7730,N_5068,N_7461);
or U7731 (N_7731,N_7408,N_6921);
xnor U7732 (N_7732,N_6162,N_5675);
and U7733 (N_7733,N_7092,N_7479);
and U7734 (N_7734,N_5532,N_5877);
nand U7735 (N_7735,N_7209,N_7295);
nor U7736 (N_7736,N_6451,N_6753);
nor U7737 (N_7737,N_5971,N_5441);
and U7738 (N_7738,N_5710,N_5075);
nand U7739 (N_7739,N_6392,N_7316);
nand U7740 (N_7740,N_6967,N_6919);
nor U7741 (N_7741,N_5673,N_5024);
nand U7742 (N_7742,N_5745,N_7015);
or U7743 (N_7743,N_5430,N_6578);
and U7744 (N_7744,N_6692,N_5381);
nor U7745 (N_7745,N_6448,N_6301);
nor U7746 (N_7746,N_6604,N_6855);
nand U7747 (N_7747,N_5539,N_5469);
and U7748 (N_7748,N_5767,N_6525);
or U7749 (N_7749,N_5922,N_6733);
and U7750 (N_7750,N_6822,N_7153);
or U7751 (N_7751,N_5709,N_5367);
nand U7752 (N_7752,N_5773,N_7474);
xor U7753 (N_7753,N_5894,N_5548);
nand U7754 (N_7754,N_5955,N_5392);
nor U7755 (N_7755,N_6550,N_6665);
and U7756 (N_7756,N_6925,N_7175);
nand U7757 (N_7757,N_6527,N_6440);
nor U7758 (N_7758,N_7080,N_6648);
and U7759 (N_7759,N_7283,N_5876);
xor U7760 (N_7760,N_5703,N_6161);
and U7761 (N_7761,N_6568,N_6138);
and U7762 (N_7762,N_6986,N_6300);
and U7763 (N_7763,N_6126,N_6344);
nand U7764 (N_7764,N_6927,N_6436);
nor U7765 (N_7765,N_5834,N_6048);
and U7766 (N_7766,N_7159,N_5431);
and U7767 (N_7767,N_6883,N_5546);
nor U7768 (N_7768,N_5554,N_6824);
nand U7769 (N_7769,N_7337,N_6646);
xor U7770 (N_7770,N_5019,N_6427);
and U7771 (N_7771,N_5130,N_7006);
and U7772 (N_7772,N_7310,N_6856);
or U7773 (N_7773,N_5350,N_6131);
or U7774 (N_7774,N_7213,N_6564);
or U7775 (N_7775,N_7146,N_6495);
and U7776 (N_7776,N_5807,N_6676);
or U7777 (N_7777,N_6699,N_6211);
xor U7778 (N_7778,N_6847,N_6670);
nor U7779 (N_7779,N_6793,N_7389);
or U7780 (N_7780,N_5500,N_6130);
xnor U7781 (N_7781,N_6941,N_6991);
nor U7782 (N_7782,N_5704,N_6877);
nand U7783 (N_7783,N_7037,N_6572);
nor U7784 (N_7784,N_6652,N_7182);
nor U7785 (N_7785,N_7356,N_5364);
nor U7786 (N_7786,N_7150,N_6693);
and U7787 (N_7787,N_7200,N_6546);
or U7788 (N_7788,N_6880,N_7158);
nor U7789 (N_7789,N_6007,N_5101);
and U7790 (N_7790,N_7239,N_6743);
and U7791 (N_7791,N_5912,N_5806);
or U7792 (N_7792,N_6689,N_5302);
or U7793 (N_7793,N_5868,N_6179);
xnor U7794 (N_7794,N_5345,N_5304);
nand U7795 (N_7795,N_5453,N_5223);
and U7796 (N_7796,N_6981,N_5813);
and U7797 (N_7797,N_6713,N_7222);
nor U7798 (N_7798,N_5682,N_5141);
and U7799 (N_7799,N_7147,N_6455);
or U7800 (N_7800,N_5005,N_5991);
and U7801 (N_7801,N_6152,N_5800);
or U7802 (N_7802,N_5730,N_7456);
nor U7803 (N_7803,N_5817,N_7308);
or U7804 (N_7804,N_7381,N_7180);
nor U7805 (N_7805,N_5452,N_5022);
and U7806 (N_7806,N_6186,N_5107);
xor U7807 (N_7807,N_6090,N_6062);
and U7808 (N_7808,N_5420,N_7378);
nor U7809 (N_7809,N_5789,N_6839);
or U7810 (N_7810,N_7325,N_5127);
or U7811 (N_7811,N_7028,N_5566);
nor U7812 (N_7812,N_5419,N_6043);
xor U7813 (N_7813,N_6383,N_7067);
nor U7814 (N_7814,N_5697,N_6583);
nor U7815 (N_7815,N_6178,N_5216);
nor U7816 (N_7816,N_5929,N_5103);
and U7817 (N_7817,N_5029,N_7324);
or U7818 (N_7818,N_6626,N_7166);
or U7819 (N_7819,N_6112,N_5402);
nand U7820 (N_7820,N_6796,N_5520);
or U7821 (N_7821,N_6401,N_5230);
nand U7822 (N_7822,N_6960,N_6969);
nand U7823 (N_7823,N_5519,N_5764);
or U7824 (N_7824,N_5616,N_7419);
and U7825 (N_7825,N_6098,N_7297);
and U7826 (N_7826,N_5718,N_6780);
xnor U7827 (N_7827,N_7494,N_6660);
nor U7828 (N_7828,N_5956,N_5822);
nor U7829 (N_7829,N_6309,N_6478);
or U7830 (N_7830,N_6000,N_5353);
nor U7831 (N_7831,N_6053,N_6288);
nor U7832 (N_7832,N_6351,N_6170);
nor U7833 (N_7833,N_6603,N_6848);
or U7834 (N_7834,N_6526,N_7328);
or U7835 (N_7835,N_6678,N_5330);
nor U7836 (N_7836,N_5873,N_6241);
and U7837 (N_7837,N_6277,N_6266);
and U7838 (N_7838,N_7095,N_5284);
or U7839 (N_7839,N_5377,N_5758);
or U7840 (N_7840,N_5565,N_5173);
xor U7841 (N_7841,N_6782,N_6939);
or U7842 (N_7842,N_5799,N_5457);
or U7843 (N_7843,N_5814,N_7338);
nor U7844 (N_7844,N_5556,N_6248);
nor U7845 (N_7845,N_6240,N_5380);
nor U7846 (N_7846,N_7260,N_6540);
and U7847 (N_7847,N_5159,N_5082);
or U7848 (N_7848,N_7197,N_5891);
nand U7849 (N_7849,N_5902,N_5911);
or U7850 (N_7850,N_5643,N_6915);
or U7851 (N_7851,N_6619,N_5874);
nand U7852 (N_7852,N_5472,N_6166);
nor U7853 (N_7853,N_7347,N_5319);
and U7854 (N_7854,N_6027,N_5211);
and U7855 (N_7855,N_5825,N_6677);
nand U7856 (N_7856,N_5646,N_7394);
or U7857 (N_7857,N_6799,N_5083);
nor U7858 (N_7858,N_5671,N_7412);
nor U7859 (N_7859,N_5761,N_5299);
or U7860 (N_7860,N_7462,N_6498);
and U7861 (N_7861,N_7179,N_5169);
or U7862 (N_7862,N_5976,N_6786);
nor U7863 (N_7863,N_6510,N_6065);
nand U7864 (N_7864,N_6347,N_5639);
nand U7865 (N_7865,N_6106,N_5752);
and U7866 (N_7866,N_5559,N_5138);
nand U7867 (N_7867,N_5294,N_6054);
or U7868 (N_7868,N_6851,N_5613);
nand U7869 (N_7869,N_6373,N_5034);
and U7870 (N_7870,N_7299,N_5746);
nor U7871 (N_7871,N_5049,N_6265);
nor U7872 (N_7872,N_7066,N_6205);
and U7873 (N_7873,N_5734,N_6124);
or U7874 (N_7874,N_7421,N_5667);
nor U7875 (N_7875,N_6669,N_6238);
nand U7876 (N_7876,N_7346,N_5043);
xnor U7877 (N_7877,N_7195,N_6445);
or U7878 (N_7878,N_5097,N_5805);
nor U7879 (N_7879,N_5349,N_6212);
nor U7880 (N_7880,N_6810,N_6135);
nor U7881 (N_7881,N_6711,N_5644);
nor U7882 (N_7882,N_6999,N_6791);
nand U7883 (N_7883,N_7001,N_5050);
nor U7884 (N_7884,N_6685,N_6929);
and U7885 (N_7885,N_6001,N_5270);
nor U7886 (N_7886,N_5409,N_5098);
and U7887 (N_7887,N_5048,N_5462);
or U7888 (N_7888,N_7398,N_5898);
and U7889 (N_7889,N_7133,N_6795);
nor U7890 (N_7890,N_6709,N_6537);
xnor U7891 (N_7891,N_5823,N_7384);
nor U7892 (N_7892,N_6346,N_5100);
nor U7893 (N_7893,N_6555,N_5028);
xnor U7894 (N_7894,N_6311,N_7387);
nand U7895 (N_7895,N_6585,N_6217);
nand U7896 (N_7896,N_5683,N_7061);
or U7897 (N_7897,N_7443,N_6989);
and U7898 (N_7898,N_5670,N_6593);
nor U7899 (N_7899,N_6600,N_5206);
or U7900 (N_7900,N_7332,N_6763);
nand U7901 (N_7901,N_5849,N_5919);
and U7902 (N_7902,N_6785,N_7465);
nor U7903 (N_7903,N_5166,N_5707);
and U7904 (N_7904,N_5287,N_6879);
and U7905 (N_7905,N_6332,N_5610);
nand U7906 (N_7906,N_7174,N_6457);
and U7907 (N_7907,N_6631,N_5046);
nand U7908 (N_7908,N_5798,N_6751);
or U7909 (N_7909,N_6861,N_7413);
nor U7910 (N_7910,N_5635,N_5209);
or U7911 (N_7911,N_6460,N_5833);
nand U7912 (N_7912,N_6082,N_5732);
nand U7913 (N_7913,N_6228,N_7241);
nor U7914 (N_7914,N_5265,N_6481);
or U7915 (N_7915,N_6591,N_5081);
and U7916 (N_7916,N_6147,N_7259);
nor U7917 (N_7917,N_6020,N_6333);
nand U7918 (N_7918,N_6038,N_6042);
or U7919 (N_7919,N_7246,N_6337);
and U7920 (N_7920,N_6538,N_5213);
and U7921 (N_7921,N_6008,N_6673);
nor U7922 (N_7922,N_6881,N_5257);
or U7923 (N_7923,N_5323,N_5998);
or U7924 (N_7924,N_5526,N_6384);
nor U7925 (N_7925,N_5543,N_6625);
nand U7926 (N_7926,N_5064,N_6884);
and U7927 (N_7927,N_5089,N_5150);
nand U7928 (N_7928,N_5731,N_5301);
or U7929 (N_7929,N_6348,N_6486);
and U7930 (N_7930,N_7097,N_6472);
nand U7931 (N_7931,N_7234,N_6438);
xnor U7932 (N_7932,N_6303,N_6061);
or U7933 (N_7933,N_6443,N_6696);
and U7934 (N_7934,N_5315,N_6869);
nand U7935 (N_7935,N_5266,N_6127);
nor U7936 (N_7936,N_6654,N_5797);
xor U7937 (N_7937,N_6803,N_5227);
nor U7938 (N_7938,N_5246,N_5882);
nand U7939 (N_7939,N_5993,N_7459);
or U7940 (N_7940,N_5968,N_7319);
xnor U7941 (N_7941,N_7071,N_5008);
or U7942 (N_7942,N_5685,N_7128);
or U7943 (N_7943,N_5283,N_7350);
or U7944 (N_7944,N_5791,N_6917);
nand U7945 (N_7945,N_6187,N_5511);
nor U7946 (N_7946,N_5180,N_6252);
or U7947 (N_7947,N_6396,N_6698);
or U7948 (N_7948,N_6873,N_5442);
nor U7949 (N_7949,N_5966,N_6645);
or U7950 (N_7950,N_5658,N_7207);
nor U7951 (N_7951,N_7363,N_5663);
and U7952 (N_7952,N_6829,N_6256);
nand U7953 (N_7953,N_5934,N_5513);
nor U7954 (N_7954,N_6662,N_7176);
and U7955 (N_7955,N_6747,N_5640);
nand U7956 (N_7956,N_7077,N_6870);
and U7957 (N_7957,N_6273,N_7351);
nor U7958 (N_7958,N_5642,N_5581);
nor U7959 (N_7959,N_5242,N_7123);
and U7960 (N_7960,N_6599,N_6260);
or U7961 (N_7961,N_5953,N_6125);
nor U7962 (N_7962,N_6110,N_7455);
or U7963 (N_7963,N_7342,N_5406);
nand U7964 (N_7964,N_5052,N_7248);
nand U7965 (N_7965,N_5175,N_6462);
or U7966 (N_7966,N_6980,N_5914);
nor U7967 (N_7967,N_6172,N_6154);
and U7968 (N_7968,N_5449,N_6041);
nor U7969 (N_7969,N_5949,N_5025);
nor U7970 (N_7970,N_6140,N_7440);
or U7971 (N_7971,N_6723,N_5607);
xor U7972 (N_7972,N_5931,N_5305);
xnor U7973 (N_7973,N_6541,N_5755);
nor U7974 (N_7974,N_6305,N_7298);
or U7975 (N_7975,N_5085,N_6350);
nor U7976 (N_7976,N_5404,N_7414);
nand U7977 (N_7977,N_5156,N_5631);
and U7978 (N_7978,N_6637,N_5515);
or U7979 (N_7979,N_7268,N_6805);
nand U7980 (N_7980,N_5516,N_7288);
and U7981 (N_7981,N_5338,N_6387);
nand U7982 (N_7982,N_5009,N_5212);
nor U7983 (N_7983,N_6534,N_6359);
nand U7984 (N_7984,N_7476,N_7075);
nand U7985 (N_7985,N_7049,N_7296);
and U7986 (N_7986,N_5006,N_7021);
and U7987 (N_7987,N_6418,N_6983);
or U7988 (N_7988,N_6226,N_6529);
nand U7989 (N_7989,N_5926,N_5438);
or U7990 (N_7990,N_5318,N_5487);
nand U7991 (N_7991,N_6237,N_7045);
and U7992 (N_7992,N_6562,N_5292);
nand U7993 (N_7993,N_5310,N_7102);
or U7994 (N_7994,N_6916,N_5142);
nand U7995 (N_7995,N_5387,N_6115);
nor U7996 (N_7996,N_5120,N_6764);
and U7997 (N_7997,N_5535,N_5149);
and U7998 (N_7998,N_7084,N_5405);
nor U7999 (N_7999,N_5247,N_5440);
and U8000 (N_8000,N_5688,N_6372);
and U8001 (N_8001,N_7486,N_6321);
and U8002 (N_8002,N_7190,N_6412);
and U8003 (N_8003,N_6632,N_5503);
xor U8004 (N_8004,N_7254,N_6116);
and U8005 (N_8005,N_6787,N_6932);
or U8006 (N_8006,N_6679,N_5428);
or U8007 (N_8007,N_6964,N_7372);
nand U8008 (N_8008,N_5285,N_6775);
or U8009 (N_8009,N_6833,N_6993);
nor U8010 (N_8010,N_6378,N_6836);
xor U8011 (N_8011,N_5273,N_5741);
or U8012 (N_8012,N_5328,N_7373);
nor U8013 (N_8013,N_5468,N_7302);
and U8014 (N_8014,N_5587,N_7043);
or U8015 (N_8015,N_6539,N_6118);
nand U8016 (N_8016,N_5721,N_6731);
nand U8017 (N_8017,N_7478,N_5344);
and U8018 (N_8018,N_7034,N_7068);
and U8019 (N_8019,N_6614,N_7072);
and U8020 (N_8020,N_5679,N_6108);
or U8021 (N_8021,N_5573,N_7424);
nand U8022 (N_8022,N_5634,N_5220);
xnor U8023 (N_8023,N_5176,N_7444);
or U8024 (N_8024,N_6623,N_5356);
or U8025 (N_8025,N_6734,N_5057);
and U8026 (N_8026,N_6595,N_6949);
or U8027 (N_8027,N_6413,N_6336);
and U8028 (N_8028,N_5932,N_6868);
and U8029 (N_8029,N_7409,N_6640);
nor U8030 (N_8030,N_7385,N_5011);
or U8031 (N_8031,N_5809,N_6377);
or U8032 (N_8032,N_5125,N_6948);
nor U8033 (N_8033,N_5358,N_6209);
and U8034 (N_8034,N_7334,N_5542);
and U8035 (N_8035,N_6184,N_6894);
nor U8036 (N_8036,N_5694,N_6105);
or U8037 (N_8037,N_5296,N_7156);
nand U8038 (N_8038,N_5579,N_6119);
and U8039 (N_8039,N_5990,N_5382);
or U8040 (N_8040,N_7335,N_7364);
and U8041 (N_8041,N_5666,N_6566);
nor U8042 (N_8042,N_5608,N_6905);
nand U8043 (N_8043,N_6484,N_5368);
nor U8044 (N_8044,N_5262,N_6867);
nand U8045 (N_8045,N_6900,N_5742);
xor U8046 (N_8046,N_5137,N_5256);
nor U8047 (N_8047,N_6294,N_6997);
or U8048 (N_8048,N_6627,N_6159);
and U8049 (N_8049,N_7108,N_5649);
or U8050 (N_8050,N_5720,N_5847);
xnor U8051 (N_8051,N_5612,N_5617);
nor U8052 (N_8052,N_5477,N_7247);
and U8053 (N_8053,N_6067,N_5357);
xor U8054 (N_8054,N_6560,N_7368);
nor U8055 (N_8055,N_6176,N_5152);
and U8056 (N_8056,N_5592,N_5041);
xnor U8057 (N_8057,N_7212,N_6653);
or U8058 (N_8058,N_6310,N_5193);
xor U8059 (N_8059,N_6956,N_7145);
nor U8060 (N_8060,N_5222,N_7477);
or U8061 (N_8061,N_5947,N_5979);
and U8062 (N_8062,N_6363,N_6466);
xnor U8063 (N_8063,N_6656,N_6133);
xor U8064 (N_8064,N_6695,N_7464);
xor U8065 (N_8065,N_7249,N_5432);
nand U8066 (N_8066,N_5994,N_5558);
nor U8067 (N_8067,N_6299,N_7018);
nor U8068 (N_8068,N_6866,N_7131);
nor U8069 (N_8069,N_5249,N_6827);
nor U8070 (N_8070,N_5831,N_5636);
nand U8071 (N_8071,N_6196,N_5412);
and U8072 (N_8072,N_6442,N_7447);
nor U8073 (N_8073,N_5853,N_6137);
nand U8074 (N_8074,N_7050,N_5396);
xnor U8075 (N_8075,N_7138,N_5341);
xor U8076 (N_8076,N_5753,N_7008);
or U8077 (N_8077,N_6930,N_6643);
nand U8078 (N_8078,N_7460,N_5713);
or U8079 (N_8079,N_5016,N_7357);
and U8080 (N_8080,N_7360,N_7467);
nand U8081 (N_8081,N_5916,N_7183);
and U8082 (N_8082,N_5907,N_5736);
and U8083 (N_8083,N_5389,N_6582);
and U8084 (N_8084,N_6094,N_7196);
nor U8085 (N_8085,N_5633,N_7204);
nand U8086 (N_8086,N_5112,N_7091);
nand U8087 (N_8087,N_7040,N_6411);
and U8088 (N_8088,N_5460,N_6702);
nor U8089 (N_8089,N_7157,N_5884);
or U8090 (N_8090,N_7489,N_5066);
nand U8091 (N_8091,N_5363,N_5313);
or U8092 (N_8092,N_6024,N_5115);
nand U8093 (N_8093,N_5650,N_5648);
nand U8094 (N_8094,N_5210,N_5444);
and U8095 (N_8095,N_6895,N_6229);
nor U8096 (N_8096,N_7290,N_6806);
nor U8097 (N_8097,N_5977,N_7148);
nand U8098 (N_8098,N_5072,N_7418);
nor U8099 (N_8099,N_7046,N_5749);
or U8100 (N_8100,N_6756,N_6181);
and U8101 (N_8101,N_6406,N_6794);
nand U8102 (N_8102,N_6778,N_5422);
nor U8103 (N_8103,N_6590,N_6477);
nor U8104 (N_8104,N_7417,N_5739);
or U8105 (N_8105,N_5110,N_7407);
or U8106 (N_8106,N_6239,N_7305);
nand U8107 (N_8107,N_6164,N_7470);
xor U8108 (N_8108,N_6033,N_5842);
xnor U8109 (N_8109,N_5174,N_5754);
nand U8110 (N_8110,N_5915,N_7468);
or U8111 (N_8111,N_7027,N_5748);
xnor U8112 (N_8112,N_6766,N_6554);
or U8113 (N_8113,N_6663,N_6842);
and U8114 (N_8114,N_5194,N_5905);
and U8115 (N_8115,N_7142,N_7416);
nand U8116 (N_8116,N_5091,N_5232);
and U8117 (N_8117,N_5601,N_7345);
nor U8118 (N_8118,N_6714,N_5133);
nand U8119 (N_8119,N_6979,N_6724);
and U8120 (N_8120,N_5669,N_6821);
xnor U8121 (N_8121,N_6817,N_7438);
and U8122 (N_8122,N_6704,N_5326);
nand U8123 (N_8123,N_6173,N_6633);
nor U8124 (N_8124,N_6261,N_6143);
and U8125 (N_8125,N_5215,N_6958);
xor U8126 (N_8126,N_5415,N_6901);
nor U8127 (N_8127,N_5031,N_6023);
and U8128 (N_8128,N_5514,N_5394);
or U8129 (N_8129,N_6129,N_7383);
nor U8130 (N_8130,N_5808,N_6334);
and U8131 (N_8131,N_5537,N_5254);
and U8132 (N_8132,N_5655,N_6849);
or U8133 (N_8133,N_7315,N_6317);
nor U8134 (N_8134,N_5552,N_5935);
nor U8135 (N_8135,N_7025,N_5131);
and U8136 (N_8136,N_5944,N_7451);
nor U8137 (N_8137,N_5886,N_6744);
and U8138 (N_8138,N_6647,N_7111);
nor U8139 (N_8139,N_7481,N_6269);
and U8140 (N_8140,N_5940,N_6819);
nor U8141 (N_8141,N_7005,N_5837);
nand U8142 (N_8142,N_6468,N_5439);
and U8143 (N_8143,N_6761,N_6439);
nor U8144 (N_8144,N_5482,N_6542);
nand U8145 (N_8145,N_5574,N_5591);
nor U8146 (N_8146,N_6314,N_5538);
nor U8147 (N_8147,N_6227,N_5255);
or U8148 (N_8148,N_7292,N_5196);
nand U8149 (N_8149,N_7210,N_6081);
and U8150 (N_8150,N_6551,N_5866);
or U8151 (N_8151,N_6419,N_5918);
and U8152 (N_8152,N_7032,N_5803);
xnor U8153 (N_8153,N_6057,N_6762);
nand U8154 (N_8154,N_6093,N_7426);
nand U8155 (N_8155,N_6198,N_6732);
nor U8156 (N_8156,N_7059,N_5423);
and U8157 (N_8157,N_5603,N_5491);
and U8158 (N_8158,N_7044,N_7087);
nor U8159 (N_8159,N_6474,N_5399);
nor U8160 (N_8160,N_5893,N_5145);
and U8161 (N_8161,N_6191,N_7172);
xor U8162 (N_8162,N_5859,N_6911);
nor U8163 (N_8163,N_6319,N_7031);
and U8164 (N_8164,N_6236,N_5498);
and U8165 (N_8165,N_6078,N_6666);
nor U8166 (N_8166,N_6429,N_7362);
nor U8167 (N_8167,N_7012,N_6746);
and U8168 (N_8168,N_5819,N_7446);
xor U8169 (N_8169,N_5827,N_6779);
and U8170 (N_8170,N_6434,N_5668);
and U8171 (N_8171,N_5941,N_6890);
nor U8172 (N_8172,N_5860,N_6099);
nor U8173 (N_8173,N_5198,N_7013);
nand U8174 (N_8174,N_7165,N_6188);
or U8175 (N_8175,N_6609,N_6028);
and U8176 (N_8176,N_6397,N_5116);
nand U8177 (N_8177,N_6897,N_6258);
nand U8178 (N_8178,N_6010,N_5776);
nand U8179 (N_8179,N_7208,N_7441);
nand U8180 (N_8180,N_5279,N_7427);
nand U8181 (N_8181,N_6621,N_6749);
and U8182 (N_8182,N_5681,N_5020);
and U8183 (N_8183,N_5769,N_6493);
nand U8184 (N_8184,N_6607,N_6617);
nor U8185 (N_8185,N_5727,N_6075);
or U8186 (N_8186,N_6530,N_5495);
nor U8187 (N_8187,N_5867,N_6584);
nor U8188 (N_8188,N_5306,N_6973);
and U8189 (N_8189,N_6331,N_7240);
and U8190 (N_8190,N_6040,N_5965);
nor U8191 (N_8191,N_7062,N_5464);
and U8192 (N_8192,N_6853,N_5657);
xnor U8193 (N_8193,N_7300,N_5093);
nor U8194 (N_8194,N_5986,N_6658);
xnor U8195 (N_8195,N_5471,N_6606);
or U8196 (N_8196,N_5014,N_5786);
nand U8197 (N_8197,N_5693,N_6644);
xor U8198 (N_8198,N_7490,N_5411);
xor U8199 (N_8199,N_6329,N_7094);
and U8200 (N_8200,N_5119,N_6463);
and U8201 (N_8201,N_6461,N_7033);
and U8202 (N_8202,N_6515,N_6707);
nor U8203 (N_8203,N_6080,N_5522);
and U8204 (N_8204,N_5843,N_6136);
xnor U8205 (N_8205,N_5641,N_5700);
or U8206 (N_8206,N_6091,N_6852);
nor U8207 (N_8207,N_5692,N_7199);
xor U8208 (N_8208,N_5497,N_6479);
xor U8209 (N_8209,N_7191,N_6769);
and U8210 (N_8210,N_5414,N_5037);
nand U8211 (N_8211,N_6938,N_5735);
nor U8212 (N_8212,N_7469,N_7056);
xor U8213 (N_8213,N_6449,N_7103);
and U8214 (N_8214,N_5621,N_5942);
or U8215 (N_8215,N_6183,N_7343);
nor U8216 (N_8216,N_6045,N_6748);
and U8217 (N_8217,N_7130,N_5200);
or U8218 (N_8218,N_7303,N_6287);
and U8219 (N_8219,N_5370,N_6922);
or U8220 (N_8220,N_5544,N_7035);
nand U8221 (N_8221,N_6850,N_5835);
or U8222 (N_8222,N_5960,N_6854);
and U8223 (N_8223,N_5158,N_6642);
nand U8224 (N_8224,N_7177,N_5090);
xnor U8225 (N_8225,N_5863,N_6423);
nor U8226 (N_8226,N_5384,N_6503);
xor U8227 (N_8227,N_6285,N_6543);
nand U8228 (N_8228,N_5623,N_5711);
nand U8229 (N_8229,N_6518,N_5475);
nand U8230 (N_8230,N_5488,N_6157);
and U8231 (N_8231,N_6937,N_5340);
xnor U8232 (N_8232,N_7306,N_5740);
nand U8233 (N_8233,N_6345,N_6755);
nand U8234 (N_8234,N_6655,N_5190);
nand U8235 (N_8235,N_7244,N_5408);
nor U8236 (N_8236,N_6996,N_5102);
and U8237 (N_8237,N_7104,N_6912);
or U8238 (N_8238,N_5716,N_6073);
nand U8239 (N_8239,N_7082,N_5638);
xor U8240 (N_8240,N_7060,N_7187);
and U8241 (N_8241,N_5564,N_5026);
nand U8242 (N_8242,N_5937,N_6367);
or U8243 (N_8243,N_7184,N_7493);
and U8244 (N_8244,N_5059,N_6142);
xor U8245 (N_8245,N_6798,N_7265);
or U8246 (N_8246,N_5372,N_6977);
nand U8247 (N_8247,N_5714,N_6417);
and U8248 (N_8248,N_6343,N_5857);
or U8249 (N_8249,N_6107,N_5963);
xor U8250 (N_8250,N_6657,N_5851);
and U8251 (N_8251,N_5274,N_6971);
xnor U8252 (N_8252,N_5307,N_5199);
nor U8253 (N_8253,N_6740,N_5225);
or U8254 (N_8254,N_6934,N_6923);
or U8255 (N_8255,N_5999,N_6596);
and U8256 (N_8256,N_6742,N_5241);
and U8257 (N_8257,N_6416,N_7445);
or U8258 (N_8258,N_7171,N_7193);
nor U8259 (N_8259,N_7000,N_6597);
or U8260 (N_8260,N_5555,N_6837);
or U8261 (N_8261,N_7277,N_7433);
or U8262 (N_8262,N_6402,N_6797);
nand U8263 (N_8263,N_6943,N_5490);
and U8264 (N_8264,N_6674,N_7223);
and U8265 (N_8265,N_5531,N_5772);
xor U8266 (N_8266,N_7101,N_6499);
or U8267 (N_8267,N_5379,N_5750);
and U8268 (N_8268,N_5794,N_6528);
or U8269 (N_8269,N_7422,N_6862);
and U8270 (N_8270,N_5995,N_6182);
or U8271 (N_8271,N_6019,N_5787);
nor U8272 (N_8272,N_6210,N_6066);
and U8273 (N_8273,N_5982,N_5191);
nor U8274 (N_8274,N_6274,N_5909);
nand U8275 (N_8275,N_6146,N_7341);
nand U8276 (N_8276,N_6490,N_6876);
or U8277 (N_8277,N_6990,N_5303);
nand U8278 (N_8278,N_6031,N_7330);
xor U8279 (N_8279,N_7160,N_5035);
xor U8280 (N_8280,N_6611,N_6508);
or U8281 (N_8281,N_5810,N_6494);
and U8282 (N_8282,N_5140,N_6857);
nor U8283 (N_8283,N_5348,N_7367);
nand U8284 (N_8284,N_5551,N_7088);
or U8285 (N_8285,N_7030,N_5637);
nor U8286 (N_8286,N_5992,N_7051);
and U8287 (N_8287,N_5435,N_6860);
and U8288 (N_8288,N_7458,N_5970);
or U8289 (N_8289,N_5346,N_6558);
or U8290 (N_8290,N_6563,N_6379);
nand U8291 (N_8291,N_6328,N_6612);
nor U8292 (N_8292,N_6326,N_5774);
or U8293 (N_8293,N_5852,N_7425);
or U8294 (N_8294,N_5844,N_6052);
or U8295 (N_8295,N_6395,N_7406);
or U8296 (N_8296,N_7136,N_7105);
nor U8297 (N_8297,N_5366,N_5954);
nand U8298 (N_8298,N_6447,N_6267);
nor U8299 (N_8299,N_6316,N_7457);
or U8300 (N_8300,N_6195,N_7267);
and U8301 (N_8301,N_5691,N_5424);
nor U8302 (N_8302,N_6976,N_6664);
nand U8303 (N_8303,N_6565,N_6680);
and U8304 (N_8304,N_6088,N_7178);
nand U8305 (N_8305,N_5153,N_6390);
nand U8306 (N_8306,N_5760,N_7386);
xnor U8307 (N_8307,N_7215,N_5939);
nand U8308 (N_8308,N_5445,N_5337);
and U8309 (N_8309,N_5117,N_6335);
xnor U8310 (N_8310,N_7411,N_6284);
nand U8311 (N_8311,N_5410,N_6914);
xnor U8312 (N_8312,N_6686,N_5078);
and U8313 (N_8313,N_6092,N_6908);
nor U8314 (N_8314,N_5336,N_5987);
nor U8315 (N_8315,N_6349,N_5135);
nor U8316 (N_8316,N_6232,N_6491);
and U8317 (N_8317,N_6243,N_5494);
nor U8318 (N_8318,N_5881,N_5609);
or U8319 (N_8319,N_5855,N_6924);
nand U8320 (N_8320,N_6414,N_6936);
nor U8321 (N_8321,N_7272,N_5756);
or U8322 (N_8322,N_5595,N_7081);
nor U8323 (N_8323,N_5985,N_6452);
nor U8324 (N_8324,N_6888,N_7119);
xor U8325 (N_8325,N_5463,N_6570);
nand U8326 (N_8326,N_5796,N_6158);
and U8327 (N_8327,N_6920,N_6768);
nand U8328 (N_8328,N_7189,N_5582);
nand U8329 (N_8329,N_6251,N_7036);
and U8330 (N_8330,N_7168,N_6651);
or U8331 (N_8331,N_6244,N_6255);
and U8332 (N_8332,N_7206,N_5804);
and U8333 (N_8333,N_6407,N_5436);
nand U8334 (N_8334,N_7011,N_7017);
nor U8335 (N_8335,N_5959,N_5862);
nor U8336 (N_8336,N_5506,N_6725);
nand U8337 (N_8337,N_6035,N_6047);
nor U8338 (N_8338,N_7395,N_5036);
and U8339 (N_8339,N_7113,N_6174);
or U8340 (N_8340,N_6327,N_7273);
and U8341 (N_8341,N_6180,N_7352);
or U8342 (N_8342,N_6758,N_6221);
xor U8343 (N_8343,N_5615,N_6544);
nor U8344 (N_8344,N_5989,N_7243);
or U8345 (N_8345,N_5715,N_6858);
and U8346 (N_8346,N_6364,N_6573);
xor U8347 (N_8347,N_7403,N_7366);
or U8348 (N_8348,N_7393,N_5004);
nor U8349 (N_8349,N_5373,N_5680);
or U8350 (N_8350,N_5447,N_5067);
or U8351 (N_8351,N_5996,N_6716);
or U8352 (N_8352,N_7331,N_5007);
nand U8353 (N_8353,N_5385,N_7214);
and U8354 (N_8354,N_5314,N_7078);
nand U8355 (N_8355,N_6691,N_5355);
nor U8356 (N_8356,N_5620,N_6155);
nor U8357 (N_8357,N_6323,N_6885);
or U8358 (N_8358,N_6505,N_6741);
nor U8359 (N_8359,N_7279,N_6831);
nor U8360 (N_8360,N_6965,N_6500);
xor U8361 (N_8361,N_7377,N_6087);
nor U8362 (N_8362,N_5943,N_7064);
nand U8363 (N_8363,N_6259,N_6718);
nand U8364 (N_8364,N_6032,N_5459);
xor U8365 (N_8365,N_5264,N_6381);
and U8366 (N_8366,N_5096,N_7452);
nor U8367 (N_8367,N_5978,N_5630);
and U8368 (N_8368,N_6814,N_5512);
nor U8369 (N_8369,N_5614,N_6497);
nand U8370 (N_8370,N_7253,N_7252);
nand U8371 (N_8371,N_6103,N_6489);
nand U8372 (N_8372,N_7144,N_6341);
nand U8373 (N_8373,N_5567,N_6820);
nor U8374 (N_8374,N_5836,N_6194);
xnor U8375 (N_8375,N_5757,N_6523);
nand U8376 (N_8376,N_7251,N_5571);
xor U8377 (N_8377,N_7107,N_6736);
and U8378 (N_8378,N_5553,N_7323);
nand U8379 (N_8379,N_6026,N_5775);
xor U8380 (N_8380,N_7326,N_5229);
and U8381 (N_8381,N_6910,N_5865);
and U8382 (N_8382,N_6220,N_7149);
nand U8383 (N_8383,N_6132,N_6012);
or U8384 (N_8384,N_7161,N_5042);
nor U8385 (N_8385,N_7238,N_7304);
nor U8386 (N_8386,N_6635,N_5015);
and U8387 (N_8387,N_6368,N_6700);
or U8388 (N_8388,N_7225,N_7220);
nand U8389 (N_8389,N_5108,N_6441);
and U8390 (N_8390,N_6006,N_6404);
and U8391 (N_8391,N_5665,N_6340);
or U8392 (N_8392,N_7262,N_7230);
xnor U8393 (N_8393,N_6594,N_5365);
nand U8394 (N_8394,N_6223,N_7275);
nand U8395 (N_8395,N_6272,N_6683);
nand U8396 (N_8396,N_5003,N_6909);
xnor U8397 (N_8397,N_6018,N_6063);
nand U8398 (N_8398,N_7358,N_6219);
nand U8399 (N_8399,N_6168,N_6144);
xor U8400 (N_8400,N_5961,N_5359);
nand U8401 (N_8401,N_6102,N_7020);
nor U8402 (N_8402,N_6592,N_7263);
nand U8403 (N_8403,N_6512,N_6304);
nand U8404 (N_8404,N_7487,N_6225);
and U8405 (N_8405,N_5964,N_5058);
nor U8406 (N_8406,N_7475,N_5622);
and U8407 (N_8407,N_5830,N_6072);
nand U8408 (N_8408,N_5659,N_5568);
nand U8409 (N_8409,N_7042,N_7236);
and U8410 (N_8410,N_6634,N_5618);
and U8411 (N_8411,N_6249,N_5951);
or U8412 (N_8412,N_6306,N_6610);
or U8413 (N_8413,N_6015,N_5762);
xor U8414 (N_8414,N_6420,N_6400);
or U8415 (N_8415,N_5590,N_5333);
nand U8416 (N_8416,N_7047,N_6097);
nand U8417 (N_8417,N_5509,N_5674);
and U8418 (N_8418,N_6875,N_6037);
or U8419 (N_8419,N_7282,N_7321);
or U8420 (N_8420,N_6830,N_5339);
nand U8421 (N_8421,N_6230,N_5228);
or U8422 (N_8422,N_5234,N_6954);
or U8423 (N_8423,N_7397,N_6060);
nor U8424 (N_8424,N_6636,N_7472);
or U8425 (N_8425,N_7219,N_5545);
and U8426 (N_8426,N_6771,N_5540);
or U8427 (N_8427,N_5053,N_6754);
and U8428 (N_8428,N_5077,N_6167);
nor U8429 (N_8429,N_5123,N_5160);
xnor U8430 (N_8430,N_5224,N_6502);
nor U8431 (N_8431,N_6650,N_6101);
nor U8432 (N_8432,N_6366,N_5719);
xor U8433 (N_8433,N_6339,N_5969);
nand U8434 (N_8434,N_7070,N_6356);
nor U8435 (N_8435,N_6160,N_6025);
and U8436 (N_8436,N_5645,N_5157);
nor U8437 (N_8437,N_5790,N_5272);
nand U8438 (N_8438,N_5278,N_5374);
nor U8439 (N_8439,N_6069,N_6681);
nand U8440 (N_8440,N_6902,N_7155);
or U8441 (N_8441,N_5664,N_5343);
and U8442 (N_8442,N_6574,N_5240);
nor U8443 (N_8443,N_6777,N_5662);
nor U8444 (N_8444,N_5864,N_5395);
or U8445 (N_8445,N_5672,N_6330);
nand U8446 (N_8446,N_6781,N_6720);
nand U8447 (N_8447,N_7437,N_5154);
nor U8448 (N_8448,N_5722,N_5235);
or U8449 (N_8449,N_5560,N_5168);
nor U8450 (N_8450,N_5099,N_6371);
nand U8451 (N_8451,N_6151,N_6506);
and U8452 (N_8452,N_6459,N_5879);
nor U8453 (N_8453,N_6496,N_7307);
xor U8454 (N_8454,N_6467,N_7453);
nor U8455 (N_8455,N_6889,N_5455);
xor U8456 (N_8456,N_6393,N_6899);
nor U8457 (N_8457,N_5690,N_5793);
nand U8458 (N_8458,N_7284,N_7348);
nand U8459 (N_8459,N_6322,N_5896);
nand U8460 (N_8460,N_7312,N_5481);
and U8461 (N_8461,N_5695,N_6815);
nor U8462 (N_8462,N_5450,N_7449);
and U8463 (N_8463,N_7137,N_7039);
xnor U8464 (N_8464,N_6863,N_6450);
and U8465 (N_8465,N_5924,N_6134);
nor U8466 (N_8466,N_7124,N_5351);
and U8467 (N_8467,N_6953,N_5562);
or U8468 (N_8468,N_6089,N_7054);
nand U8469 (N_8469,N_5702,N_5948);
or U8470 (N_8470,N_6295,N_5678);
and U8471 (N_8471,N_7294,N_6898);
and U8472 (N_8472,N_6957,N_6208);
nand U8473 (N_8473,N_7023,N_5044);
nand U8474 (N_8474,N_5106,N_5580);
and U8475 (N_8475,N_5895,N_6608);
or U8476 (N_8476,N_5448,N_5084);
nand U8477 (N_8477,N_6083,N_6717);
or U8478 (N_8478,N_6409,N_6051);
and U8479 (N_8479,N_7380,N_5594);
and U8480 (N_8480,N_6992,N_5354);
nor U8481 (N_8481,N_5829,N_6264);
nor U8482 (N_8482,N_6308,N_5465);
nand U8483 (N_8483,N_6446,N_6605);
nor U8484 (N_8484,N_6935,N_5687);
nor U8485 (N_8485,N_5219,N_7016);
and U8486 (N_8486,N_6545,N_6469);
nor U8487 (N_8487,N_7374,N_6320);
xor U8488 (N_8488,N_6050,N_7311);
or U8489 (N_8489,N_6003,N_7371);
nand U8490 (N_8490,N_7127,N_7233);
or U8491 (N_8491,N_7423,N_5856);
xnor U8492 (N_8492,N_6139,N_7293);
nand U8493 (N_8493,N_6859,N_6668);
nor U8494 (N_8494,N_5063,N_5458);
nor U8495 (N_8495,N_5391,N_6719);
xor U8496 (N_8496,N_5550,N_5845);
nor U8497 (N_8497,N_5606,N_7221);
and U8498 (N_8498,N_6324,N_5821);
nand U8499 (N_8499,N_6886,N_6913);
nand U8500 (N_8500,N_7112,N_5818);
nand U8501 (N_8501,N_5071,N_6952);
or U8502 (N_8502,N_7361,N_6408);
nand U8503 (N_8503,N_7309,N_6887);
and U8504 (N_8504,N_5632,N_5712);
nand U8505 (N_8505,N_6988,N_5467);
xor U8506 (N_8506,N_6475,N_5892);
and U8507 (N_8507,N_7100,N_7086);
nor U8508 (N_8508,N_5226,N_5060);
nor U8509 (N_8509,N_6430,N_6882);
nor U8510 (N_8510,N_6079,N_6703);
or U8511 (N_8511,N_5407,N_5074);
xor U8512 (N_8512,N_7402,N_6739);
nor U8513 (N_8513,N_6630,N_7379);
or U8514 (N_8514,N_6826,N_5416);
nand U8515 (N_8515,N_5163,N_6616);
nor U8516 (N_8516,N_5483,N_6388);
nand U8517 (N_8517,N_7271,N_7218);
or U8518 (N_8518,N_6788,N_7492);
xor U8519 (N_8519,N_5699,N_6100);
or U8520 (N_8520,N_5124,N_5508);
and U8521 (N_8521,N_7415,N_7349);
and U8522 (N_8522,N_5575,N_5869);
nand U8523 (N_8523,N_6995,N_5525);
nor U8524 (N_8524,N_7198,N_5263);
or U8525 (N_8525,N_6365,N_6235);
xor U8526 (N_8526,N_5121,N_5167);
or U8527 (N_8527,N_6864,N_7405);
and U8528 (N_8528,N_5012,N_6874);
or U8529 (N_8529,N_6004,N_6750);
or U8530 (N_8530,N_5777,N_7228);
and U8531 (N_8531,N_5563,N_5561);
xor U8532 (N_8532,N_7227,N_5221);
nor U8533 (N_8533,N_7266,N_5456);
nor U8534 (N_8534,N_5957,N_6811);
or U8535 (N_8535,N_5501,N_6375);
and U8536 (N_8536,N_6801,N_7188);
nand U8537 (N_8537,N_7231,N_5282);
or U8538 (N_8538,N_5023,N_6561);
or U8539 (N_8539,N_6201,N_6567);
xnor U8540 (N_8540,N_5887,N_5801);
and U8541 (N_8541,N_5838,N_6896);
nor U8542 (N_8542,N_6405,N_5476);
or U8543 (N_8543,N_6575,N_7052);
nor U8544 (N_8544,N_7287,N_5062);
and U8545 (N_8545,N_6222,N_5737);
nand U8546 (N_8546,N_5421,N_6705);
xor U8547 (N_8547,N_6813,N_6193);
or U8548 (N_8548,N_5361,N_5974);
and U8549 (N_8549,N_5967,N_6974);
nand U8550 (N_8550,N_7085,N_7129);
and U8551 (N_8551,N_6944,N_7026);
and U8552 (N_8552,N_7181,N_5231);
nor U8553 (N_8553,N_6153,N_7454);
or U8554 (N_8554,N_6587,N_6807);
nand U8555 (N_8555,N_6522,N_7375);
xor U8556 (N_8556,N_6684,N_5300);
and U8557 (N_8557,N_5324,N_7121);
nand U8558 (N_8558,N_6846,N_5000);
nand U8559 (N_8559,N_6710,N_6415);
nand U8560 (N_8560,N_6962,N_6556);
or U8561 (N_8561,N_6021,N_7471);
nand U8562 (N_8562,N_5290,N_6738);
xnor U8563 (N_8563,N_7169,N_6342);
or U8564 (N_8564,N_7336,N_7203);
or U8565 (N_8565,N_7076,N_6192);
or U8566 (N_8566,N_6055,N_5426);
and U8567 (N_8567,N_6809,N_5597);
or U8568 (N_8568,N_5237,N_6077);
or U8569 (N_8569,N_6520,N_6398);
nor U8570 (N_8570,N_5725,N_6076);
nand U8571 (N_8571,N_6789,N_6998);
and U8572 (N_8572,N_5651,N_6832);
or U8573 (N_8573,N_5920,N_7495);
and U8574 (N_8574,N_5840,N_6017);
or U8575 (N_8575,N_7163,N_5504);
nor U8576 (N_8576,N_5182,N_5510);
or U8577 (N_8577,N_5523,N_6760);
or U8578 (N_8578,N_6624,N_5783);
and U8579 (N_8579,N_6380,N_5250);
and U8580 (N_8580,N_5624,N_5171);
nand U8581 (N_8581,N_5529,N_7053);
nand U8582 (N_8582,N_5360,N_7353);
nand U8583 (N_8583,N_5207,N_6872);
nor U8584 (N_8584,N_5288,N_6878);
nor U8585 (N_8585,N_6985,N_6649);
and U8586 (N_8586,N_6706,N_5461);
and U8587 (N_8587,N_6511,N_5815);
and U8588 (N_8588,N_5192,N_6009);
and U8589 (N_8589,N_5047,N_5586);
nor U8590 (N_8590,N_5619,N_6165);
nand U8591 (N_8591,N_6951,N_6471);
nor U8592 (N_8592,N_6620,N_7173);
nand U8593 (N_8593,N_6982,N_6357);
nor U8594 (N_8594,N_7029,N_5785);
nor U8595 (N_8595,N_7069,N_7022);
or U8596 (N_8596,N_5238,N_6374);
nor U8597 (N_8597,N_7430,N_6257);
nor U8598 (N_8598,N_5293,N_6581);
or U8599 (N_8599,N_5647,N_7090);
or U8600 (N_8600,N_5276,N_5010);
nand U8601 (N_8601,N_5611,N_7167);
or U8602 (N_8602,N_5889,N_7289);
nor U8603 (N_8603,N_6589,N_7192);
and U8604 (N_8604,N_5493,N_5654);
nor U8605 (N_8605,N_6675,N_5308);
or U8606 (N_8606,N_6485,N_7055);
xor U8607 (N_8607,N_5040,N_7211);
and U8608 (N_8608,N_7498,N_6386);
or U8609 (N_8609,N_5208,N_6360);
nor U8610 (N_8610,N_5705,N_6784);
nand U8611 (N_8611,N_5151,N_6891);
and U8612 (N_8612,N_6697,N_7089);
and U8613 (N_8613,N_6085,N_5329);
nor U8614 (N_8614,N_7274,N_6483);
nand U8615 (N_8615,N_5362,N_6435);
xnor U8616 (N_8616,N_5352,N_7099);
or U8617 (N_8617,N_5070,N_6569);
nor U8618 (N_8618,N_5195,N_7370);
and U8619 (N_8619,N_5585,N_6120);
nor U8620 (N_8620,N_6672,N_7436);
or U8621 (N_8621,N_7264,N_6959);
and U8622 (N_8622,N_7057,N_5177);
and U8623 (N_8623,N_6667,N_6275);
nor U8624 (N_8624,N_5802,N_5018);
nor U8625 (N_8625,N_5170,N_5017);
and U8626 (N_8626,N_7141,N_5335);
nand U8627 (N_8627,N_6128,N_5251);
or U8628 (N_8628,N_7114,N_5788);
nand U8629 (N_8629,N_5485,N_6034);
and U8630 (N_8630,N_6940,N_5846);
nor U8631 (N_8631,N_5507,N_5528);
and U8632 (N_8632,N_6918,N_5277);
and U8633 (N_8633,N_5850,N_5187);
and U8634 (N_8634,N_5466,N_6148);
nand U8635 (N_8635,N_7134,N_5747);
xor U8636 (N_8636,N_5122,N_7224);
nor U8637 (N_8637,N_5795,N_5095);
or U8638 (N_8638,N_5291,N_5766);
and U8639 (N_8639,N_5883,N_5437);
nor U8640 (N_8640,N_6056,N_6727);
nor U8641 (N_8641,N_5988,N_5885);
nand U8642 (N_8642,N_6458,N_7250);
and U8643 (N_8643,N_6361,N_5342);
and U8644 (N_8644,N_6970,N_5661);
and U8645 (N_8645,N_5534,N_6197);
or U8646 (N_8646,N_5604,N_7497);
nand U8647 (N_8647,N_5980,N_6424);
or U8648 (N_8648,N_5701,N_6254);
nand U8649 (N_8649,N_7355,N_5473);
nand U8650 (N_8650,N_6586,N_5689);
and U8651 (N_8651,N_5812,N_5027);
nand U8652 (N_8652,N_7420,N_6480);
nand U8653 (N_8653,N_5726,N_5723);
and U8654 (N_8654,N_5203,N_6531);
nor U8655 (N_8655,N_5470,N_5038);
or U8656 (N_8656,N_6571,N_5738);
nand U8657 (N_8657,N_6835,N_6629);
nand U8658 (N_8658,N_6121,N_7340);
or U8659 (N_8659,N_5588,N_6163);
and U8660 (N_8660,N_5136,N_5094);
or U8661 (N_8661,N_7216,N_6464);
nand U8662 (N_8662,N_5286,N_5056);
or U8663 (N_8663,N_5936,N_5233);
and U8664 (N_8664,N_7226,N_6576);
nor U8665 (N_8665,N_6270,N_7314);
nor U8666 (N_8666,N_7162,N_5923);
and U8667 (N_8667,N_6453,N_5295);
nor U8668 (N_8668,N_6524,N_6262);
nor U8669 (N_8669,N_5144,N_5946);
nor U8670 (N_8670,N_6906,N_7245);
xnor U8671 (N_8671,N_6059,N_5289);
nand U8672 (N_8672,N_7276,N_6338);
and U8673 (N_8673,N_7369,N_7281);
and U8674 (N_8674,N_5733,N_6946);
or U8675 (N_8675,N_6804,N_6708);
nor U8676 (N_8676,N_5413,N_6456);
and U8677 (N_8677,N_5496,N_6307);
nor U8678 (N_8678,N_7048,N_5928);
nand U8679 (N_8679,N_5729,N_6297);
nor U8680 (N_8680,N_6246,N_5499);
nor U8681 (N_8681,N_5316,N_5243);
xor U8682 (N_8682,N_5311,N_5418);
or U8683 (N_8683,N_5111,N_6994);
or U8684 (N_8684,N_5297,N_6588);
nor U8685 (N_8685,N_5239,N_6353);
nor U8686 (N_8686,N_5536,N_5779);
or U8687 (N_8687,N_5533,N_7235);
and U8688 (N_8688,N_5065,N_5371);
nor U8689 (N_8689,N_6068,N_7170);
nor U8690 (N_8690,N_6123,N_6501);
or U8691 (N_8691,N_6114,N_5627);
and U8692 (N_8692,N_5524,N_5147);
and U8693 (N_8693,N_5839,N_6433);
or U8694 (N_8694,N_6701,N_7257);
or U8695 (N_8695,N_6280,N_6776);
and U8696 (N_8696,N_6292,N_6659);
or U8697 (N_8697,N_7285,N_7410);
xor U8698 (N_8698,N_6278,N_5576);
and U8699 (N_8699,N_6984,N_6504);
and U8700 (N_8700,N_7098,N_6963);
or U8701 (N_8701,N_6521,N_5079);
xnor U8702 (N_8702,N_6759,N_5155);
nor U8703 (N_8703,N_6014,N_6312);
and U8704 (N_8704,N_6354,N_6190);
nand U8705 (N_8705,N_5309,N_6202);
nor U8706 (N_8706,N_7466,N_7439);
nand U8707 (N_8707,N_6425,N_7329);
and U8708 (N_8708,N_6871,N_6049);
nand U8709 (N_8709,N_5577,N_6145);
and U8710 (N_8710,N_6783,N_5826);
and U8711 (N_8711,N_7428,N_6016);
and U8712 (N_8712,N_5181,N_5317);
xor U8713 (N_8713,N_6476,N_6276);
and U8714 (N_8714,N_5161,N_6113);
and U8715 (N_8715,N_5401,N_7318);
nand U8716 (N_8716,N_6773,N_6729);
nor U8717 (N_8717,N_5217,N_5185);
nor U8718 (N_8718,N_6892,N_6358);
or U8719 (N_8719,N_5569,N_6271);
xnor U8720 (N_8720,N_5386,N_6687);
and U8721 (N_8721,N_5434,N_5973);
or U8722 (N_8722,N_6058,N_7382);
and U8723 (N_8723,N_7237,N_6111);
nor U8724 (N_8724,N_6250,N_5032);
nand U8725 (N_8725,N_5321,N_5676);
nor U8726 (N_8726,N_5521,N_6770);
or U8727 (N_8727,N_6199,N_5792);
nand U8728 (N_8728,N_5921,N_5105);
nor U8729 (N_8729,N_6482,N_6628);
nand U8730 (N_8730,N_6834,N_6513);
and U8731 (N_8731,N_7093,N_6096);
nor U8732 (N_8732,N_5375,N_5197);
nand U8733 (N_8733,N_5871,N_6084);
nand U8734 (N_8734,N_7491,N_5484);
xor U8735 (N_8735,N_6488,N_5202);
and U8736 (N_8736,N_7232,N_6410);
nand U8737 (N_8737,N_7083,N_6233);
nand U8738 (N_8738,N_5021,N_7396);
or U8739 (N_8739,N_6171,N_6200);
and U8740 (N_8740,N_6865,N_5784);
and U8741 (N_8741,N_5474,N_7024);
or U8742 (N_8742,N_7473,N_5271);
or U8743 (N_8743,N_6492,N_5900);
nand U8744 (N_8744,N_6432,N_5393);
and U8745 (N_8745,N_5143,N_5088);
nor U8746 (N_8746,N_7286,N_7354);
and U8747 (N_8747,N_5930,N_5076);
or U8748 (N_8748,N_6638,N_5981);
xnor U8749 (N_8749,N_5486,N_6370);
and U8750 (N_8750,N_5308,N_6462);
nand U8751 (N_8751,N_5915,N_5909);
nor U8752 (N_8752,N_5668,N_6016);
and U8753 (N_8753,N_5591,N_5713);
nor U8754 (N_8754,N_7434,N_7002);
or U8755 (N_8755,N_5454,N_6632);
nand U8756 (N_8756,N_5630,N_6017);
nand U8757 (N_8757,N_5757,N_5961);
nand U8758 (N_8758,N_5883,N_6571);
and U8759 (N_8759,N_5176,N_5412);
or U8760 (N_8760,N_5030,N_5560);
or U8761 (N_8761,N_6075,N_7067);
nor U8762 (N_8762,N_6430,N_6885);
xnor U8763 (N_8763,N_7353,N_5726);
and U8764 (N_8764,N_6403,N_5904);
nor U8765 (N_8765,N_6934,N_5130);
or U8766 (N_8766,N_5925,N_5230);
nand U8767 (N_8767,N_7171,N_5759);
xnor U8768 (N_8768,N_7013,N_6486);
xor U8769 (N_8769,N_6238,N_6142);
nor U8770 (N_8770,N_6774,N_5742);
and U8771 (N_8771,N_6465,N_6911);
and U8772 (N_8772,N_7294,N_5023);
nor U8773 (N_8773,N_5479,N_6792);
and U8774 (N_8774,N_7238,N_5725);
or U8775 (N_8775,N_5867,N_7104);
nor U8776 (N_8776,N_6536,N_6417);
nand U8777 (N_8777,N_7096,N_5505);
nor U8778 (N_8778,N_7027,N_7426);
or U8779 (N_8779,N_6925,N_6811);
nand U8780 (N_8780,N_5771,N_6194);
and U8781 (N_8781,N_6676,N_6745);
or U8782 (N_8782,N_6539,N_6542);
or U8783 (N_8783,N_7147,N_5447);
nor U8784 (N_8784,N_5724,N_7414);
and U8785 (N_8785,N_5362,N_7386);
nor U8786 (N_8786,N_6946,N_7120);
nor U8787 (N_8787,N_6150,N_7042);
xnor U8788 (N_8788,N_6566,N_5252);
or U8789 (N_8789,N_5400,N_5570);
nor U8790 (N_8790,N_5687,N_6191);
nand U8791 (N_8791,N_6795,N_6489);
nand U8792 (N_8792,N_5865,N_5240);
and U8793 (N_8793,N_6598,N_5427);
xor U8794 (N_8794,N_6685,N_5902);
nor U8795 (N_8795,N_5349,N_6147);
or U8796 (N_8796,N_5596,N_6614);
nand U8797 (N_8797,N_6338,N_6219);
nor U8798 (N_8798,N_5092,N_5008);
nor U8799 (N_8799,N_5357,N_6796);
or U8800 (N_8800,N_7295,N_7349);
or U8801 (N_8801,N_5417,N_7318);
or U8802 (N_8802,N_5193,N_6179);
and U8803 (N_8803,N_5042,N_6925);
nand U8804 (N_8804,N_5005,N_5480);
nor U8805 (N_8805,N_5163,N_5733);
nand U8806 (N_8806,N_6038,N_5448);
and U8807 (N_8807,N_5599,N_5258);
or U8808 (N_8808,N_5331,N_7234);
and U8809 (N_8809,N_5434,N_6848);
nand U8810 (N_8810,N_6703,N_7376);
nand U8811 (N_8811,N_7108,N_5860);
or U8812 (N_8812,N_6871,N_5840);
xor U8813 (N_8813,N_5473,N_5475);
nor U8814 (N_8814,N_5436,N_6952);
nand U8815 (N_8815,N_6328,N_7370);
xnor U8816 (N_8816,N_5548,N_5390);
or U8817 (N_8817,N_6671,N_6827);
nand U8818 (N_8818,N_7118,N_6556);
nor U8819 (N_8819,N_5505,N_6836);
nand U8820 (N_8820,N_7304,N_6155);
or U8821 (N_8821,N_6940,N_6813);
nand U8822 (N_8822,N_6856,N_7257);
nor U8823 (N_8823,N_7301,N_5571);
nand U8824 (N_8824,N_6837,N_6835);
nor U8825 (N_8825,N_6145,N_5779);
nor U8826 (N_8826,N_6431,N_5086);
nand U8827 (N_8827,N_5696,N_6896);
xor U8828 (N_8828,N_7020,N_7392);
and U8829 (N_8829,N_6612,N_6346);
xnor U8830 (N_8830,N_5421,N_6485);
nor U8831 (N_8831,N_6213,N_5880);
and U8832 (N_8832,N_6352,N_5059);
nand U8833 (N_8833,N_6368,N_7062);
nand U8834 (N_8834,N_6751,N_6738);
nor U8835 (N_8835,N_5240,N_5803);
xor U8836 (N_8836,N_6659,N_7201);
or U8837 (N_8837,N_6952,N_6294);
nand U8838 (N_8838,N_6842,N_5360);
or U8839 (N_8839,N_6018,N_7217);
nor U8840 (N_8840,N_5552,N_7444);
and U8841 (N_8841,N_6048,N_7361);
or U8842 (N_8842,N_5610,N_5948);
nor U8843 (N_8843,N_5210,N_6659);
nor U8844 (N_8844,N_5776,N_7039);
xnor U8845 (N_8845,N_5794,N_7353);
nor U8846 (N_8846,N_6990,N_5566);
nand U8847 (N_8847,N_5210,N_5493);
and U8848 (N_8848,N_5826,N_6680);
and U8849 (N_8849,N_5480,N_6126);
nor U8850 (N_8850,N_5643,N_5847);
and U8851 (N_8851,N_6580,N_5753);
and U8852 (N_8852,N_5344,N_6914);
xor U8853 (N_8853,N_6841,N_7385);
nor U8854 (N_8854,N_5523,N_5135);
nand U8855 (N_8855,N_6412,N_5965);
nor U8856 (N_8856,N_5301,N_5773);
and U8857 (N_8857,N_5401,N_6832);
xor U8858 (N_8858,N_6136,N_6352);
nand U8859 (N_8859,N_7210,N_6969);
and U8860 (N_8860,N_6390,N_5801);
nand U8861 (N_8861,N_6926,N_5047);
and U8862 (N_8862,N_5433,N_5323);
nand U8863 (N_8863,N_7421,N_5993);
nand U8864 (N_8864,N_5155,N_6733);
nor U8865 (N_8865,N_5315,N_6151);
nand U8866 (N_8866,N_5658,N_5280);
and U8867 (N_8867,N_6742,N_5904);
or U8868 (N_8868,N_7183,N_5824);
or U8869 (N_8869,N_5919,N_6742);
xor U8870 (N_8870,N_5883,N_5740);
nand U8871 (N_8871,N_7253,N_5982);
nand U8872 (N_8872,N_5986,N_5749);
nor U8873 (N_8873,N_6724,N_7081);
nor U8874 (N_8874,N_5839,N_5831);
and U8875 (N_8875,N_6865,N_5647);
nand U8876 (N_8876,N_7131,N_6169);
and U8877 (N_8877,N_6835,N_5217);
nor U8878 (N_8878,N_6901,N_6942);
nor U8879 (N_8879,N_5766,N_5898);
and U8880 (N_8880,N_5937,N_6387);
nor U8881 (N_8881,N_6067,N_5049);
nor U8882 (N_8882,N_6358,N_5237);
nor U8883 (N_8883,N_7279,N_5221);
nand U8884 (N_8884,N_5137,N_7114);
and U8885 (N_8885,N_5600,N_7049);
and U8886 (N_8886,N_5614,N_5968);
and U8887 (N_8887,N_5585,N_5107);
and U8888 (N_8888,N_5829,N_7293);
nand U8889 (N_8889,N_6915,N_7221);
or U8890 (N_8890,N_7090,N_6835);
nand U8891 (N_8891,N_6328,N_5636);
nand U8892 (N_8892,N_5970,N_6125);
nand U8893 (N_8893,N_6258,N_6503);
and U8894 (N_8894,N_5106,N_5358);
and U8895 (N_8895,N_5848,N_5449);
nand U8896 (N_8896,N_6343,N_5112);
nand U8897 (N_8897,N_7055,N_7085);
and U8898 (N_8898,N_6083,N_6131);
and U8899 (N_8899,N_5068,N_6849);
or U8900 (N_8900,N_5204,N_6640);
and U8901 (N_8901,N_6951,N_6961);
xor U8902 (N_8902,N_5986,N_7024);
nor U8903 (N_8903,N_6417,N_5055);
or U8904 (N_8904,N_5299,N_5249);
xor U8905 (N_8905,N_5200,N_5204);
nand U8906 (N_8906,N_7412,N_5466);
nand U8907 (N_8907,N_6209,N_6831);
and U8908 (N_8908,N_6851,N_5807);
or U8909 (N_8909,N_5616,N_7246);
nand U8910 (N_8910,N_7388,N_7430);
nor U8911 (N_8911,N_5371,N_6115);
nand U8912 (N_8912,N_6630,N_6145);
nor U8913 (N_8913,N_5893,N_5368);
or U8914 (N_8914,N_5615,N_6854);
and U8915 (N_8915,N_5350,N_5262);
nand U8916 (N_8916,N_5083,N_5118);
nor U8917 (N_8917,N_7187,N_5894);
nor U8918 (N_8918,N_5793,N_6983);
or U8919 (N_8919,N_6882,N_6047);
and U8920 (N_8920,N_7147,N_6995);
and U8921 (N_8921,N_5057,N_7417);
and U8922 (N_8922,N_6783,N_5052);
nand U8923 (N_8923,N_5133,N_5503);
or U8924 (N_8924,N_5891,N_7465);
nand U8925 (N_8925,N_6444,N_7420);
xnor U8926 (N_8926,N_6011,N_6603);
and U8927 (N_8927,N_7385,N_5882);
nand U8928 (N_8928,N_5192,N_7202);
nor U8929 (N_8929,N_5287,N_6332);
and U8930 (N_8930,N_5484,N_6368);
or U8931 (N_8931,N_5030,N_5581);
or U8932 (N_8932,N_6375,N_5599);
and U8933 (N_8933,N_6988,N_5267);
xnor U8934 (N_8934,N_5408,N_5346);
or U8935 (N_8935,N_5907,N_5660);
xnor U8936 (N_8936,N_5984,N_5452);
or U8937 (N_8937,N_6749,N_6495);
nand U8938 (N_8938,N_6961,N_5072);
nor U8939 (N_8939,N_5534,N_6509);
xnor U8940 (N_8940,N_6052,N_6273);
nand U8941 (N_8941,N_5773,N_6759);
xnor U8942 (N_8942,N_7144,N_5483);
nand U8943 (N_8943,N_5456,N_5970);
nor U8944 (N_8944,N_5496,N_7040);
nand U8945 (N_8945,N_6675,N_5719);
nor U8946 (N_8946,N_5129,N_5045);
nand U8947 (N_8947,N_6992,N_7026);
nand U8948 (N_8948,N_5990,N_5713);
or U8949 (N_8949,N_5068,N_5102);
nor U8950 (N_8950,N_6162,N_5758);
or U8951 (N_8951,N_6771,N_6745);
xor U8952 (N_8952,N_6165,N_5909);
and U8953 (N_8953,N_6046,N_5800);
or U8954 (N_8954,N_5256,N_6354);
or U8955 (N_8955,N_7217,N_6438);
or U8956 (N_8956,N_5369,N_7185);
nand U8957 (N_8957,N_6064,N_5367);
or U8958 (N_8958,N_5293,N_5640);
nand U8959 (N_8959,N_5148,N_7498);
and U8960 (N_8960,N_6157,N_5472);
nor U8961 (N_8961,N_7073,N_6783);
and U8962 (N_8962,N_6289,N_6614);
nor U8963 (N_8963,N_6887,N_6550);
nor U8964 (N_8964,N_7209,N_7011);
or U8965 (N_8965,N_6730,N_5116);
and U8966 (N_8966,N_5190,N_6239);
nand U8967 (N_8967,N_5197,N_5862);
nand U8968 (N_8968,N_6181,N_5994);
and U8969 (N_8969,N_6922,N_6410);
nand U8970 (N_8970,N_7093,N_6466);
nor U8971 (N_8971,N_6327,N_6912);
and U8972 (N_8972,N_6158,N_6627);
and U8973 (N_8973,N_5718,N_5066);
nand U8974 (N_8974,N_6429,N_6419);
or U8975 (N_8975,N_6188,N_5002);
nand U8976 (N_8976,N_5684,N_6542);
nor U8977 (N_8977,N_6835,N_7233);
and U8978 (N_8978,N_6035,N_5735);
or U8979 (N_8979,N_6609,N_7291);
nand U8980 (N_8980,N_7414,N_5443);
and U8981 (N_8981,N_6387,N_5420);
nor U8982 (N_8982,N_7298,N_6741);
or U8983 (N_8983,N_6344,N_6358);
nor U8984 (N_8984,N_7056,N_7245);
or U8985 (N_8985,N_7265,N_5379);
xor U8986 (N_8986,N_7236,N_7392);
nor U8987 (N_8987,N_6367,N_6680);
nand U8988 (N_8988,N_6687,N_6535);
xnor U8989 (N_8989,N_5305,N_5114);
and U8990 (N_8990,N_7068,N_5109);
or U8991 (N_8991,N_6396,N_5804);
xnor U8992 (N_8992,N_5993,N_6987);
or U8993 (N_8993,N_6379,N_6678);
nand U8994 (N_8994,N_5634,N_5135);
nand U8995 (N_8995,N_6403,N_6431);
and U8996 (N_8996,N_5146,N_5694);
xor U8997 (N_8997,N_7091,N_7363);
nand U8998 (N_8998,N_5719,N_6160);
nor U8999 (N_8999,N_5067,N_7415);
or U9000 (N_9000,N_7394,N_6116);
nor U9001 (N_9001,N_7078,N_7378);
or U9002 (N_9002,N_6230,N_5452);
nand U9003 (N_9003,N_7311,N_5998);
nor U9004 (N_9004,N_5066,N_5609);
and U9005 (N_9005,N_5344,N_5771);
nand U9006 (N_9006,N_5767,N_5187);
or U9007 (N_9007,N_5197,N_7061);
nand U9008 (N_9008,N_5625,N_5856);
nor U9009 (N_9009,N_6746,N_6432);
and U9010 (N_9010,N_7127,N_7409);
or U9011 (N_9011,N_7088,N_7240);
nor U9012 (N_9012,N_6811,N_7138);
nand U9013 (N_9013,N_6770,N_7349);
nor U9014 (N_9014,N_6288,N_5085);
or U9015 (N_9015,N_7143,N_5840);
nand U9016 (N_9016,N_6613,N_7302);
nor U9017 (N_9017,N_7231,N_6763);
nand U9018 (N_9018,N_7308,N_6608);
nand U9019 (N_9019,N_6578,N_5149);
xnor U9020 (N_9020,N_6708,N_6098);
nand U9021 (N_9021,N_6554,N_6220);
or U9022 (N_9022,N_5398,N_5796);
nor U9023 (N_9023,N_7383,N_6589);
or U9024 (N_9024,N_5209,N_7152);
and U9025 (N_9025,N_6136,N_6341);
and U9026 (N_9026,N_5180,N_5691);
nand U9027 (N_9027,N_7000,N_5445);
nand U9028 (N_9028,N_5568,N_6518);
and U9029 (N_9029,N_5294,N_5533);
nor U9030 (N_9030,N_6044,N_6557);
and U9031 (N_9031,N_7017,N_5858);
xor U9032 (N_9032,N_5546,N_6978);
nand U9033 (N_9033,N_6175,N_5807);
and U9034 (N_9034,N_5343,N_6611);
xnor U9035 (N_9035,N_5105,N_5693);
or U9036 (N_9036,N_5302,N_6936);
xor U9037 (N_9037,N_5408,N_5026);
and U9038 (N_9038,N_7092,N_6366);
nor U9039 (N_9039,N_5127,N_6674);
or U9040 (N_9040,N_6487,N_5560);
xnor U9041 (N_9041,N_5758,N_5311);
xor U9042 (N_9042,N_5538,N_5118);
nor U9043 (N_9043,N_5107,N_5552);
and U9044 (N_9044,N_5339,N_6590);
and U9045 (N_9045,N_7453,N_7097);
or U9046 (N_9046,N_5614,N_7269);
nand U9047 (N_9047,N_6350,N_6248);
or U9048 (N_9048,N_5533,N_5207);
xnor U9049 (N_9049,N_5081,N_5996);
xor U9050 (N_9050,N_5899,N_7170);
and U9051 (N_9051,N_6224,N_6972);
or U9052 (N_9052,N_7202,N_5806);
and U9053 (N_9053,N_6705,N_6231);
nand U9054 (N_9054,N_6724,N_5107);
or U9055 (N_9055,N_5879,N_5841);
nor U9056 (N_9056,N_7116,N_6348);
nand U9057 (N_9057,N_6374,N_6505);
and U9058 (N_9058,N_6362,N_7079);
xor U9059 (N_9059,N_7440,N_7254);
and U9060 (N_9060,N_7420,N_5502);
and U9061 (N_9061,N_6609,N_6430);
and U9062 (N_9062,N_6018,N_6796);
xnor U9063 (N_9063,N_5051,N_6042);
and U9064 (N_9064,N_6401,N_7459);
xor U9065 (N_9065,N_5958,N_5464);
nor U9066 (N_9066,N_5737,N_6724);
nand U9067 (N_9067,N_5611,N_5049);
or U9068 (N_9068,N_7344,N_6427);
xnor U9069 (N_9069,N_5729,N_6780);
nand U9070 (N_9070,N_5082,N_6390);
and U9071 (N_9071,N_7466,N_6374);
nand U9072 (N_9072,N_5423,N_5311);
nor U9073 (N_9073,N_6383,N_5568);
and U9074 (N_9074,N_5698,N_7472);
xor U9075 (N_9075,N_5277,N_6589);
xnor U9076 (N_9076,N_5037,N_7496);
nand U9077 (N_9077,N_6347,N_5938);
nor U9078 (N_9078,N_7145,N_6371);
xor U9079 (N_9079,N_5386,N_6888);
and U9080 (N_9080,N_6262,N_6506);
nor U9081 (N_9081,N_7326,N_7361);
nor U9082 (N_9082,N_5844,N_6226);
nand U9083 (N_9083,N_5449,N_6316);
and U9084 (N_9084,N_5734,N_5278);
nand U9085 (N_9085,N_5713,N_6426);
nand U9086 (N_9086,N_5760,N_6530);
and U9087 (N_9087,N_5937,N_6219);
nand U9088 (N_9088,N_6208,N_5903);
nand U9089 (N_9089,N_6368,N_6659);
and U9090 (N_9090,N_7187,N_7202);
or U9091 (N_9091,N_6213,N_5520);
nor U9092 (N_9092,N_7266,N_7415);
nor U9093 (N_9093,N_7064,N_6432);
xnor U9094 (N_9094,N_6906,N_5419);
nand U9095 (N_9095,N_5467,N_7472);
nor U9096 (N_9096,N_6627,N_5618);
nor U9097 (N_9097,N_6938,N_6355);
xnor U9098 (N_9098,N_6450,N_5576);
nor U9099 (N_9099,N_6511,N_5193);
nor U9100 (N_9100,N_6034,N_5817);
or U9101 (N_9101,N_6606,N_5026);
or U9102 (N_9102,N_6761,N_7009);
or U9103 (N_9103,N_5033,N_7134);
nor U9104 (N_9104,N_7059,N_6523);
or U9105 (N_9105,N_7479,N_7104);
nand U9106 (N_9106,N_6650,N_5801);
or U9107 (N_9107,N_6618,N_7283);
or U9108 (N_9108,N_6690,N_6364);
nor U9109 (N_9109,N_5422,N_5391);
nor U9110 (N_9110,N_5615,N_7208);
nor U9111 (N_9111,N_5438,N_5254);
or U9112 (N_9112,N_7087,N_6836);
nand U9113 (N_9113,N_6402,N_7412);
or U9114 (N_9114,N_5899,N_6080);
or U9115 (N_9115,N_7360,N_7135);
or U9116 (N_9116,N_6976,N_6817);
and U9117 (N_9117,N_6694,N_6220);
and U9118 (N_9118,N_6253,N_5927);
nor U9119 (N_9119,N_5259,N_5619);
nor U9120 (N_9120,N_6284,N_5000);
nand U9121 (N_9121,N_5709,N_7390);
nand U9122 (N_9122,N_6471,N_5895);
nand U9123 (N_9123,N_7208,N_6996);
xnor U9124 (N_9124,N_7208,N_7154);
nand U9125 (N_9125,N_5293,N_5191);
or U9126 (N_9126,N_5374,N_6198);
nand U9127 (N_9127,N_5785,N_7398);
nor U9128 (N_9128,N_5577,N_6942);
xnor U9129 (N_9129,N_5124,N_5913);
and U9130 (N_9130,N_7305,N_7128);
nand U9131 (N_9131,N_5580,N_5534);
and U9132 (N_9132,N_5780,N_7494);
and U9133 (N_9133,N_5053,N_5656);
nor U9134 (N_9134,N_7415,N_5577);
or U9135 (N_9135,N_7278,N_6747);
and U9136 (N_9136,N_6843,N_6573);
nor U9137 (N_9137,N_6417,N_5274);
nor U9138 (N_9138,N_7067,N_5950);
nand U9139 (N_9139,N_5918,N_7170);
nor U9140 (N_9140,N_5059,N_7153);
nor U9141 (N_9141,N_5360,N_6182);
nand U9142 (N_9142,N_6789,N_7480);
nor U9143 (N_9143,N_5554,N_7331);
xor U9144 (N_9144,N_6638,N_6287);
nand U9145 (N_9145,N_7132,N_6362);
and U9146 (N_9146,N_6932,N_5489);
xor U9147 (N_9147,N_5408,N_6045);
xor U9148 (N_9148,N_6823,N_6069);
nor U9149 (N_9149,N_7433,N_5119);
nor U9150 (N_9150,N_7032,N_6275);
nand U9151 (N_9151,N_5329,N_5379);
or U9152 (N_9152,N_6903,N_7407);
xor U9153 (N_9153,N_7350,N_5020);
or U9154 (N_9154,N_6503,N_6155);
xnor U9155 (N_9155,N_6298,N_5326);
and U9156 (N_9156,N_7410,N_6950);
and U9157 (N_9157,N_5753,N_6831);
or U9158 (N_9158,N_6647,N_5194);
nand U9159 (N_9159,N_6915,N_5512);
nand U9160 (N_9160,N_5399,N_5470);
xor U9161 (N_9161,N_6149,N_5502);
nand U9162 (N_9162,N_6883,N_5468);
and U9163 (N_9163,N_6879,N_5066);
or U9164 (N_9164,N_6738,N_5570);
or U9165 (N_9165,N_6069,N_5813);
or U9166 (N_9166,N_6243,N_5101);
or U9167 (N_9167,N_6247,N_5450);
xnor U9168 (N_9168,N_5685,N_6878);
or U9169 (N_9169,N_5914,N_5653);
nand U9170 (N_9170,N_6085,N_7018);
nand U9171 (N_9171,N_6255,N_5292);
nand U9172 (N_9172,N_7067,N_6186);
nor U9173 (N_9173,N_5373,N_5791);
nor U9174 (N_9174,N_6378,N_5324);
xnor U9175 (N_9175,N_6715,N_7318);
and U9176 (N_9176,N_6283,N_5570);
nor U9177 (N_9177,N_6833,N_6273);
nor U9178 (N_9178,N_6771,N_7194);
nand U9179 (N_9179,N_5421,N_6622);
nand U9180 (N_9180,N_5179,N_5660);
or U9181 (N_9181,N_7086,N_6475);
nor U9182 (N_9182,N_5574,N_5345);
and U9183 (N_9183,N_5704,N_7355);
and U9184 (N_9184,N_6206,N_6359);
or U9185 (N_9185,N_6968,N_5446);
nand U9186 (N_9186,N_7356,N_6668);
nor U9187 (N_9187,N_7017,N_6123);
nor U9188 (N_9188,N_7229,N_7196);
xor U9189 (N_9189,N_5544,N_5517);
and U9190 (N_9190,N_6813,N_7061);
and U9191 (N_9191,N_5893,N_5728);
nand U9192 (N_9192,N_7188,N_5601);
and U9193 (N_9193,N_7218,N_5538);
or U9194 (N_9194,N_5281,N_7327);
nand U9195 (N_9195,N_5439,N_7439);
and U9196 (N_9196,N_7269,N_5839);
or U9197 (N_9197,N_6158,N_7494);
and U9198 (N_9198,N_5222,N_7068);
nor U9199 (N_9199,N_6369,N_5701);
or U9200 (N_9200,N_5358,N_5885);
nor U9201 (N_9201,N_6528,N_6214);
or U9202 (N_9202,N_5498,N_6960);
and U9203 (N_9203,N_6671,N_5199);
nand U9204 (N_9204,N_6590,N_6052);
xor U9205 (N_9205,N_7377,N_7354);
nor U9206 (N_9206,N_6543,N_7488);
and U9207 (N_9207,N_7000,N_6545);
xor U9208 (N_9208,N_5628,N_7091);
nor U9209 (N_9209,N_5124,N_5230);
xnor U9210 (N_9210,N_7450,N_5190);
nor U9211 (N_9211,N_6201,N_5605);
and U9212 (N_9212,N_6450,N_6499);
nor U9213 (N_9213,N_6735,N_6014);
nand U9214 (N_9214,N_5973,N_6511);
or U9215 (N_9215,N_5032,N_5724);
or U9216 (N_9216,N_7436,N_6911);
xor U9217 (N_9217,N_7084,N_6452);
nor U9218 (N_9218,N_5248,N_6820);
or U9219 (N_9219,N_5412,N_5869);
xor U9220 (N_9220,N_7326,N_5685);
nand U9221 (N_9221,N_7490,N_5499);
and U9222 (N_9222,N_6978,N_7153);
nor U9223 (N_9223,N_5967,N_6570);
nor U9224 (N_9224,N_5064,N_5009);
nand U9225 (N_9225,N_7092,N_5845);
nor U9226 (N_9226,N_5884,N_5534);
and U9227 (N_9227,N_5877,N_6845);
xnor U9228 (N_9228,N_6769,N_6415);
nor U9229 (N_9229,N_5605,N_6181);
nand U9230 (N_9230,N_6905,N_7291);
nand U9231 (N_9231,N_5355,N_5119);
or U9232 (N_9232,N_6365,N_6617);
and U9233 (N_9233,N_5251,N_5838);
nor U9234 (N_9234,N_5740,N_7115);
or U9235 (N_9235,N_6029,N_7000);
nor U9236 (N_9236,N_6415,N_7312);
and U9237 (N_9237,N_6152,N_6046);
nand U9238 (N_9238,N_6268,N_5799);
xor U9239 (N_9239,N_7425,N_6325);
nor U9240 (N_9240,N_6215,N_6273);
or U9241 (N_9241,N_6117,N_6782);
nand U9242 (N_9242,N_5035,N_7433);
and U9243 (N_9243,N_5917,N_5489);
or U9244 (N_9244,N_7486,N_5971);
and U9245 (N_9245,N_6558,N_7079);
nor U9246 (N_9246,N_7022,N_5392);
xor U9247 (N_9247,N_6428,N_5945);
nor U9248 (N_9248,N_6389,N_6507);
nand U9249 (N_9249,N_6460,N_6981);
nand U9250 (N_9250,N_5811,N_6989);
and U9251 (N_9251,N_6161,N_7100);
and U9252 (N_9252,N_7261,N_7309);
xnor U9253 (N_9253,N_5032,N_5947);
or U9254 (N_9254,N_6651,N_5557);
nand U9255 (N_9255,N_6180,N_5270);
or U9256 (N_9256,N_7455,N_7048);
or U9257 (N_9257,N_7319,N_5421);
nor U9258 (N_9258,N_6816,N_7332);
nor U9259 (N_9259,N_5601,N_6447);
and U9260 (N_9260,N_6996,N_6220);
nand U9261 (N_9261,N_5869,N_6860);
nand U9262 (N_9262,N_7318,N_5277);
or U9263 (N_9263,N_5103,N_5401);
nand U9264 (N_9264,N_5911,N_6376);
xor U9265 (N_9265,N_7369,N_6819);
nor U9266 (N_9266,N_6563,N_5221);
nand U9267 (N_9267,N_5736,N_5868);
nor U9268 (N_9268,N_5872,N_5204);
or U9269 (N_9269,N_7089,N_5219);
xnor U9270 (N_9270,N_6850,N_5431);
nand U9271 (N_9271,N_6517,N_5773);
and U9272 (N_9272,N_6703,N_5742);
and U9273 (N_9273,N_6957,N_7421);
nor U9274 (N_9274,N_6894,N_5018);
and U9275 (N_9275,N_5814,N_6497);
nand U9276 (N_9276,N_5448,N_5613);
xor U9277 (N_9277,N_5043,N_5784);
nor U9278 (N_9278,N_6421,N_6468);
and U9279 (N_9279,N_6241,N_5993);
or U9280 (N_9280,N_5526,N_7284);
or U9281 (N_9281,N_5116,N_6115);
xnor U9282 (N_9282,N_6121,N_7328);
and U9283 (N_9283,N_6538,N_7087);
nor U9284 (N_9284,N_6848,N_6607);
or U9285 (N_9285,N_6018,N_6256);
nand U9286 (N_9286,N_5282,N_5150);
and U9287 (N_9287,N_7099,N_6977);
nor U9288 (N_9288,N_7247,N_5279);
nand U9289 (N_9289,N_5761,N_6521);
and U9290 (N_9290,N_7410,N_6122);
and U9291 (N_9291,N_5458,N_5631);
nor U9292 (N_9292,N_6981,N_7071);
nor U9293 (N_9293,N_6717,N_6830);
and U9294 (N_9294,N_6895,N_5775);
and U9295 (N_9295,N_5631,N_5448);
or U9296 (N_9296,N_7344,N_5166);
and U9297 (N_9297,N_5591,N_6623);
or U9298 (N_9298,N_5703,N_6408);
and U9299 (N_9299,N_5443,N_5290);
and U9300 (N_9300,N_6514,N_6226);
xor U9301 (N_9301,N_6359,N_5903);
and U9302 (N_9302,N_5424,N_7451);
or U9303 (N_9303,N_5970,N_6547);
nor U9304 (N_9304,N_7165,N_5912);
nor U9305 (N_9305,N_5397,N_6087);
nand U9306 (N_9306,N_5061,N_5568);
nand U9307 (N_9307,N_5093,N_5843);
nand U9308 (N_9308,N_7145,N_6990);
xnor U9309 (N_9309,N_5216,N_6468);
nor U9310 (N_9310,N_7241,N_7065);
and U9311 (N_9311,N_6162,N_6706);
and U9312 (N_9312,N_7091,N_5331);
or U9313 (N_9313,N_6013,N_5647);
xnor U9314 (N_9314,N_5172,N_7420);
or U9315 (N_9315,N_7234,N_6998);
or U9316 (N_9316,N_6629,N_5440);
nand U9317 (N_9317,N_5186,N_7434);
nor U9318 (N_9318,N_6368,N_5340);
and U9319 (N_9319,N_7000,N_5171);
or U9320 (N_9320,N_6396,N_5729);
or U9321 (N_9321,N_6949,N_6707);
and U9322 (N_9322,N_5551,N_5897);
nor U9323 (N_9323,N_5373,N_7434);
nand U9324 (N_9324,N_5047,N_6198);
nor U9325 (N_9325,N_5955,N_6283);
or U9326 (N_9326,N_7132,N_7119);
nand U9327 (N_9327,N_5540,N_7144);
or U9328 (N_9328,N_6154,N_6476);
and U9329 (N_9329,N_5746,N_7297);
or U9330 (N_9330,N_7004,N_5172);
or U9331 (N_9331,N_5489,N_7330);
nand U9332 (N_9332,N_7367,N_6060);
and U9333 (N_9333,N_6407,N_6342);
nand U9334 (N_9334,N_6008,N_6422);
nand U9335 (N_9335,N_5416,N_7318);
nand U9336 (N_9336,N_6622,N_5634);
and U9337 (N_9337,N_5252,N_7185);
and U9338 (N_9338,N_6227,N_6891);
nand U9339 (N_9339,N_5632,N_5675);
nor U9340 (N_9340,N_6125,N_5055);
nand U9341 (N_9341,N_6180,N_5578);
nor U9342 (N_9342,N_6735,N_5469);
nand U9343 (N_9343,N_7227,N_6688);
and U9344 (N_9344,N_6446,N_6689);
nor U9345 (N_9345,N_7450,N_6610);
xor U9346 (N_9346,N_6925,N_5964);
nand U9347 (N_9347,N_7049,N_5427);
nand U9348 (N_9348,N_5095,N_5802);
nand U9349 (N_9349,N_6364,N_5759);
and U9350 (N_9350,N_7093,N_6026);
xor U9351 (N_9351,N_6049,N_7225);
nor U9352 (N_9352,N_5627,N_6507);
or U9353 (N_9353,N_7214,N_5498);
or U9354 (N_9354,N_6243,N_5187);
xnor U9355 (N_9355,N_5228,N_6450);
xnor U9356 (N_9356,N_5984,N_6817);
or U9357 (N_9357,N_5217,N_7214);
nor U9358 (N_9358,N_5972,N_6591);
and U9359 (N_9359,N_7484,N_7041);
nand U9360 (N_9360,N_7339,N_6636);
or U9361 (N_9361,N_6096,N_5852);
and U9362 (N_9362,N_6603,N_5329);
or U9363 (N_9363,N_6064,N_7406);
nor U9364 (N_9364,N_6165,N_6646);
xor U9365 (N_9365,N_6997,N_6208);
or U9366 (N_9366,N_7068,N_7279);
or U9367 (N_9367,N_7213,N_6041);
nand U9368 (N_9368,N_7292,N_5155);
and U9369 (N_9369,N_6424,N_5321);
nand U9370 (N_9370,N_6647,N_7498);
nor U9371 (N_9371,N_6733,N_6211);
or U9372 (N_9372,N_5999,N_6195);
nand U9373 (N_9373,N_5688,N_5035);
nor U9374 (N_9374,N_6666,N_6211);
and U9375 (N_9375,N_6903,N_6313);
or U9376 (N_9376,N_5031,N_6991);
and U9377 (N_9377,N_6401,N_6768);
nand U9378 (N_9378,N_6179,N_6073);
and U9379 (N_9379,N_7295,N_5390);
xnor U9380 (N_9380,N_5288,N_6823);
and U9381 (N_9381,N_6499,N_6520);
nand U9382 (N_9382,N_5071,N_5168);
nand U9383 (N_9383,N_5460,N_6925);
and U9384 (N_9384,N_5063,N_5245);
and U9385 (N_9385,N_5324,N_6310);
xor U9386 (N_9386,N_6290,N_5989);
nand U9387 (N_9387,N_7328,N_6690);
xnor U9388 (N_9388,N_6063,N_6967);
and U9389 (N_9389,N_5847,N_5877);
nor U9390 (N_9390,N_5712,N_6191);
and U9391 (N_9391,N_5251,N_6895);
nand U9392 (N_9392,N_5248,N_6813);
and U9393 (N_9393,N_6606,N_6138);
and U9394 (N_9394,N_5909,N_6997);
or U9395 (N_9395,N_5907,N_5683);
xnor U9396 (N_9396,N_7021,N_5437);
nand U9397 (N_9397,N_6481,N_6640);
xnor U9398 (N_9398,N_6455,N_7062);
xnor U9399 (N_9399,N_6994,N_6665);
nand U9400 (N_9400,N_5344,N_7410);
nor U9401 (N_9401,N_7412,N_6238);
xnor U9402 (N_9402,N_7001,N_7361);
nand U9403 (N_9403,N_7164,N_6134);
nor U9404 (N_9404,N_5993,N_7135);
nand U9405 (N_9405,N_6817,N_5879);
nand U9406 (N_9406,N_7367,N_6706);
and U9407 (N_9407,N_6318,N_7109);
and U9408 (N_9408,N_5121,N_5868);
or U9409 (N_9409,N_6227,N_6617);
and U9410 (N_9410,N_5560,N_5701);
or U9411 (N_9411,N_5480,N_5501);
or U9412 (N_9412,N_5051,N_5629);
nor U9413 (N_9413,N_7031,N_7374);
nand U9414 (N_9414,N_5830,N_6100);
xnor U9415 (N_9415,N_6225,N_5282);
and U9416 (N_9416,N_6463,N_5061);
and U9417 (N_9417,N_5938,N_5441);
nor U9418 (N_9418,N_6644,N_5326);
nor U9419 (N_9419,N_6848,N_5138);
nor U9420 (N_9420,N_7001,N_6953);
nand U9421 (N_9421,N_5039,N_5779);
nor U9422 (N_9422,N_7264,N_6046);
or U9423 (N_9423,N_6983,N_6912);
xor U9424 (N_9424,N_6772,N_6931);
xor U9425 (N_9425,N_5203,N_5101);
nand U9426 (N_9426,N_6152,N_7304);
nand U9427 (N_9427,N_6709,N_6238);
or U9428 (N_9428,N_6972,N_5673);
or U9429 (N_9429,N_6908,N_5197);
nand U9430 (N_9430,N_7393,N_6878);
nand U9431 (N_9431,N_5039,N_6070);
nor U9432 (N_9432,N_7284,N_6285);
nand U9433 (N_9433,N_7311,N_5263);
nor U9434 (N_9434,N_7431,N_6422);
or U9435 (N_9435,N_6130,N_5584);
nor U9436 (N_9436,N_6026,N_5495);
or U9437 (N_9437,N_7263,N_6987);
and U9438 (N_9438,N_7431,N_5958);
nand U9439 (N_9439,N_5426,N_6935);
and U9440 (N_9440,N_5237,N_7361);
and U9441 (N_9441,N_6402,N_5449);
or U9442 (N_9442,N_6061,N_5961);
nand U9443 (N_9443,N_7294,N_6248);
nor U9444 (N_9444,N_7458,N_7179);
nand U9445 (N_9445,N_6066,N_7403);
nor U9446 (N_9446,N_7060,N_6104);
nor U9447 (N_9447,N_6142,N_7320);
and U9448 (N_9448,N_5481,N_5624);
nand U9449 (N_9449,N_5583,N_5171);
and U9450 (N_9450,N_7174,N_7359);
or U9451 (N_9451,N_6950,N_5426);
nor U9452 (N_9452,N_5055,N_5883);
nor U9453 (N_9453,N_5938,N_6206);
and U9454 (N_9454,N_5552,N_6575);
and U9455 (N_9455,N_5624,N_6194);
or U9456 (N_9456,N_7167,N_6439);
and U9457 (N_9457,N_7279,N_5521);
nand U9458 (N_9458,N_5386,N_6828);
nand U9459 (N_9459,N_6340,N_5682);
or U9460 (N_9460,N_6620,N_5486);
nor U9461 (N_9461,N_5176,N_5434);
xnor U9462 (N_9462,N_5921,N_6174);
and U9463 (N_9463,N_5194,N_7026);
nand U9464 (N_9464,N_6550,N_5665);
and U9465 (N_9465,N_6587,N_7283);
nand U9466 (N_9466,N_6327,N_6035);
nor U9467 (N_9467,N_5170,N_6222);
and U9468 (N_9468,N_5569,N_7482);
and U9469 (N_9469,N_6013,N_5750);
or U9470 (N_9470,N_6507,N_7045);
xnor U9471 (N_9471,N_6774,N_6606);
xor U9472 (N_9472,N_7092,N_6728);
nor U9473 (N_9473,N_5646,N_5409);
nand U9474 (N_9474,N_6024,N_6034);
or U9475 (N_9475,N_5543,N_5289);
nand U9476 (N_9476,N_5079,N_6365);
and U9477 (N_9477,N_6256,N_5822);
nor U9478 (N_9478,N_5283,N_5101);
or U9479 (N_9479,N_5041,N_5764);
nor U9480 (N_9480,N_6818,N_6473);
xor U9481 (N_9481,N_5998,N_5599);
or U9482 (N_9482,N_6356,N_5825);
nand U9483 (N_9483,N_7035,N_6817);
and U9484 (N_9484,N_6362,N_7090);
nor U9485 (N_9485,N_6121,N_7415);
nor U9486 (N_9486,N_6895,N_6409);
or U9487 (N_9487,N_6003,N_5564);
nor U9488 (N_9488,N_6903,N_7490);
nor U9489 (N_9489,N_5813,N_6756);
xnor U9490 (N_9490,N_5579,N_6123);
or U9491 (N_9491,N_5002,N_5397);
nand U9492 (N_9492,N_5077,N_7339);
nand U9493 (N_9493,N_6252,N_6140);
or U9494 (N_9494,N_7432,N_7334);
nand U9495 (N_9495,N_6030,N_5849);
nor U9496 (N_9496,N_6260,N_7393);
or U9497 (N_9497,N_5702,N_6248);
xor U9498 (N_9498,N_6859,N_5462);
xnor U9499 (N_9499,N_5246,N_7062);
nand U9500 (N_9500,N_6954,N_6359);
nor U9501 (N_9501,N_5395,N_6753);
and U9502 (N_9502,N_5384,N_5646);
nor U9503 (N_9503,N_6058,N_5411);
xor U9504 (N_9504,N_7426,N_5357);
and U9505 (N_9505,N_6174,N_7363);
nor U9506 (N_9506,N_5184,N_6931);
or U9507 (N_9507,N_6369,N_5582);
nor U9508 (N_9508,N_5944,N_5233);
nor U9509 (N_9509,N_7151,N_6343);
or U9510 (N_9510,N_5241,N_6830);
and U9511 (N_9511,N_6726,N_6326);
or U9512 (N_9512,N_6809,N_5613);
and U9513 (N_9513,N_5507,N_5602);
nand U9514 (N_9514,N_6587,N_5214);
xor U9515 (N_9515,N_7368,N_5689);
xnor U9516 (N_9516,N_6056,N_6408);
nand U9517 (N_9517,N_6082,N_5825);
xnor U9518 (N_9518,N_5600,N_5120);
xor U9519 (N_9519,N_6741,N_5361);
nand U9520 (N_9520,N_6120,N_5777);
and U9521 (N_9521,N_6534,N_6529);
nor U9522 (N_9522,N_5190,N_6415);
and U9523 (N_9523,N_6217,N_6877);
xor U9524 (N_9524,N_6332,N_6942);
nand U9525 (N_9525,N_6774,N_7458);
or U9526 (N_9526,N_5519,N_6367);
or U9527 (N_9527,N_7257,N_6839);
nor U9528 (N_9528,N_5989,N_7448);
or U9529 (N_9529,N_6917,N_5440);
nand U9530 (N_9530,N_5294,N_6616);
or U9531 (N_9531,N_6751,N_5036);
nor U9532 (N_9532,N_7478,N_5808);
and U9533 (N_9533,N_7393,N_5078);
or U9534 (N_9534,N_5102,N_6418);
nor U9535 (N_9535,N_5611,N_7127);
and U9536 (N_9536,N_6247,N_6451);
and U9537 (N_9537,N_5252,N_6646);
and U9538 (N_9538,N_6593,N_7335);
nand U9539 (N_9539,N_7151,N_5876);
or U9540 (N_9540,N_6354,N_6829);
nor U9541 (N_9541,N_5840,N_5740);
nor U9542 (N_9542,N_7235,N_5028);
nor U9543 (N_9543,N_7274,N_5109);
xor U9544 (N_9544,N_5931,N_5147);
nand U9545 (N_9545,N_5188,N_7083);
or U9546 (N_9546,N_6002,N_6365);
nor U9547 (N_9547,N_6698,N_5602);
nor U9548 (N_9548,N_5666,N_7240);
nand U9549 (N_9549,N_5498,N_7290);
and U9550 (N_9550,N_7229,N_5918);
and U9551 (N_9551,N_5367,N_5542);
or U9552 (N_9552,N_6899,N_6199);
and U9553 (N_9553,N_5704,N_5770);
nor U9554 (N_9554,N_6934,N_5486);
nor U9555 (N_9555,N_5792,N_5428);
nor U9556 (N_9556,N_5916,N_6127);
nor U9557 (N_9557,N_7474,N_5838);
nor U9558 (N_9558,N_5455,N_7304);
and U9559 (N_9559,N_6288,N_7263);
or U9560 (N_9560,N_7443,N_6744);
or U9561 (N_9561,N_5013,N_5915);
or U9562 (N_9562,N_5396,N_6039);
or U9563 (N_9563,N_6037,N_5260);
nand U9564 (N_9564,N_6555,N_6203);
nor U9565 (N_9565,N_7197,N_6522);
nor U9566 (N_9566,N_5134,N_5085);
or U9567 (N_9567,N_5137,N_5954);
nand U9568 (N_9568,N_6004,N_5004);
nand U9569 (N_9569,N_5685,N_5694);
or U9570 (N_9570,N_6547,N_5927);
or U9571 (N_9571,N_6107,N_6806);
and U9572 (N_9572,N_5435,N_5547);
nand U9573 (N_9573,N_6610,N_7300);
or U9574 (N_9574,N_5991,N_6378);
nand U9575 (N_9575,N_6678,N_5234);
and U9576 (N_9576,N_5973,N_5442);
or U9577 (N_9577,N_6701,N_6553);
xor U9578 (N_9578,N_5961,N_5776);
nor U9579 (N_9579,N_5706,N_7293);
nor U9580 (N_9580,N_6595,N_6769);
and U9581 (N_9581,N_7297,N_7146);
nand U9582 (N_9582,N_6632,N_5184);
nand U9583 (N_9583,N_6781,N_6533);
nor U9584 (N_9584,N_5153,N_6474);
nor U9585 (N_9585,N_7057,N_5108);
or U9586 (N_9586,N_6094,N_7109);
xnor U9587 (N_9587,N_7048,N_6049);
and U9588 (N_9588,N_5798,N_5405);
or U9589 (N_9589,N_6749,N_7415);
nor U9590 (N_9590,N_6931,N_5722);
nor U9591 (N_9591,N_6726,N_6198);
xnor U9592 (N_9592,N_7263,N_6148);
and U9593 (N_9593,N_7131,N_7045);
and U9594 (N_9594,N_7482,N_7326);
nand U9595 (N_9595,N_5458,N_5746);
and U9596 (N_9596,N_5817,N_5154);
or U9597 (N_9597,N_7439,N_6276);
or U9598 (N_9598,N_6873,N_6155);
nor U9599 (N_9599,N_5576,N_6262);
nor U9600 (N_9600,N_5712,N_6093);
or U9601 (N_9601,N_5614,N_5280);
nor U9602 (N_9602,N_6735,N_7201);
nand U9603 (N_9603,N_6882,N_6749);
nand U9604 (N_9604,N_5806,N_6740);
nand U9605 (N_9605,N_6159,N_5769);
or U9606 (N_9606,N_5955,N_5564);
xnor U9607 (N_9607,N_6204,N_6300);
nand U9608 (N_9608,N_6448,N_6182);
nand U9609 (N_9609,N_6473,N_7059);
or U9610 (N_9610,N_5986,N_6806);
and U9611 (N_9611,N_6334,N_6246);
nor U9612 (N_9612,N_6890,N_6524);
or U9613 (N_9613,N_6925,N_6899);
xnor U9614 (N_9614,N_5499,N_5033);
nor U9615 (N_9615,N_6671,N_5216);
nand U9616 (N_9616,N_6987,N_5602);
nor U9617 (N_9617,N_6945,N_6582);
nor U9618 (N_9618,N_5749,N_6481);
nand U9619 (N_9619,N_5686,N_6309);
nand U9620 (N_9620,N_5929,N_7440);
and U9621 (N_9621,N_6285,N_7393);
or U9622 (N_9622,N_6592,N_7038);
nand U9623 (N_9623,N_5347,N_6149);
and U9624 (N_9624,N_7112,N_5971);
and U9625 (N_9625,N_5264,N_6974);
and U9626 (N_9626,N_6569,N_6801);
and U9627 (N_9627,N_6715,N_6455);
nand U9628 (N_9628,N_6949,N_5273);
xnor U9629 (N_9629,N_5199,N_5294);
nor U9630 (N_9630,N_7332,N_6720);
nand U9631 (N_9631,N_5413,N_5542);
or U9632 (N_9632,N_6920,N_6037);
nand U9633 (N_9633,N_5895,N_5703);
or U9634 (N_9634,N_6380,N_7050);
xor U9635 (N_9635,N_5637,N_7034);
nand U9636 (N_9636,N_6250,N_5795);
or U9637 (N_9637,N_6966,N_6023);
nor U9638 (N_9638,N_5892,N_6933);
or U9639 (N_9639,N_5716,N_5520);
or U9640 (N_9640,N_5403,N_6368);
nor U9641 (N_9641,N_7137,N_5657);
nor U9642 (N_9642,N_5505,N_5100);
nand U9643 (N_9643,N_5988,N_5063);
nand U9644 (N_9644,N_6757,N_6772);
nor U9645 (N_9645,N_7368,N_7062);
xnor U9646 (N_9646,N_5620,N_7258);
and U9647 (N_9647,N_5983,N_7113);
nor U9648 (N_9648,N_5073,N_6580);
xnor U9649 (N_9649,N_6402,N_5087);
xor U9650 (N_9650,N_5745,N_7371);
nor U9651 (N_9651,N_6306,N_7324);
and U9652 (N_9652,N_6389,N_5602);
nand U9653 (N_9653,N_7206,N_7338);
or U9654 (N_9654,N_5557,N_6813);
and U9655 (N_9655,N_7089,N_5279);
nand U9656 (N_9656,N_5592,N_5050);
nor U9657 (N_9657,N_7081,N_7290);
nand U9658 (N_9658,N_7025,N_7011);
xnor U9659 (N_9659,N_6498,N_5003);
nand U9660 (N_9660,N_7103,N_6765);
nand U9661 (N_9661,N_5945,N_5664);
nor U9662 (N_9662,N_7378,N_6684);
or U9663 (N_9663,N_6200,N_6320);
and U9664 (N_9664,N_6434,N_6148);
nor U9665 (N_9665,N_7222,N_6313);
or U9666 (N_9666,N_7214,N_5376);
nor U9667 (N_9667,N_6442,N_6859);
and U9668 (N_9668,N_5998,N_6515);
nand U9669 (N_9669,N_5802,N_7345);
nand U9670 (N_9670,N_5932,N_5158);
and U9671 (N_9671,N_7139,N_5946);
nor U9672 (N_9672,N_5632,N_6965);
and U9673 (N_9673,N_7414,N_6993);
nor U9674 (N_9674,N_6348,N_7458);
and U9675 (N_9675,N_5410,N_7049);
and U9676 (N_9676,N_5367,N_6684);
nand U9677 (N_9677,N_5648,N_6514);
nand U9678 (N_9678,N_6946,N_6028);
nand U9679 (N_9679,N_6443,N_7036);
or U9680 (N_9680,N_5914,N_5388);
xnor U9681 (N_9681,N_6688,N_5138);
nor U9682 (N_9682,N_5878,N_6627);
or U9683 (N_9683,N_5260,N_7243);
nor U9684 (N_9684,N_7365,N_7129);
or U9685 (N_9685,N_5539,N_5500);
xnor U9686 (N_9686,N_6687,N_5500);
nand U9687 (N_9687,N_6072,N_6318);
or U9688 (N_9688,N_7257,N_5148);
xnor U9689 (N_9689,N_7292,N_5097);
and U9690 (N_9690,N_5610,N_5903);
and U9691 (N_9691,N_5355,N_6986);
xnor U9692 (N_9692,N_7479,N_6969);
or U9693 (N_9693,N_6251,N_6976);
nor U9694 (N_9694,N_7297,N_5264);
or U9695 (N_9695,N_7421,N_5234);
nor U9696 (N_9696,N_7117,N_5939);
nor U9697 (N_9697,N_7394,N_5304);
nand U9698 (N_9698,N_6121,N_5251);
and U9699 (N_9699,N_6396,N_6699);
nand U9700 (N_9700,N_6475,N_5316);
or U9701 (N_9701,N_5649,N_5916);
and U9702 (N_9702,N_5817,N_7147);
or U9703 (N_9703,N_5456,N_5398);
nor U9704 (N_9704,N_7362,N_7180);
and U9705 (N_9705,N_7409,N_6776);
xor U9706 (N_9706,N_5546,N_5771);
nor U9707 (N_9707,N_6832,N_7005);
nand U9708 (N_9708,N_6209,N_5287);
nand U9709 (N_9709,N_5929,N_5770);
and U9710 (N_9710,N_7206,N_6312);
nand U9711 (N_9711,N_6912,N_7450);
or U9712 (N_9712,N_6387,N_5231);
or U9713 (N_9713,N_5156,N_5504);
or U9714 (N_9714,N_6551,N_6838);
or U9715 (N_9715,N_5389,N_7382);
xor U9716 (N_9716,N_5625,N_6745);
nor U9717 (N_9717,N_6299,N_6963);
nand U9718 (N_9718,N_5063,N_7200);
nand U9719 (N_9719,N_5016,N_7348);
nor U9720 (N_9720,N_5344,N_5855);
nand U9721 (N_9721,N_5637,N_5392);
nor U9722 (N_9722,N_7329,N_6807);
nand U9723 (N_9723,N_5745,N_5013);
xor U9724 (N_9724,N_6864,N_5248);
nor U9725 (N_9725,N_5079,N_6742);
and U9726 (N_9726,N_7120,N_5682);
or U9727 (N_9727,N_5043,N_6298);
or U9728 (N_9728,N_7082,N_6911);
and U9729 (N_9729,N_6134,N_5282);
and U9730 (N_9730,N_7269,N_6818);
nor U9731 (N_9731,N_6544,N_6799);
nor U9732 (N_9732,N_6673,N_6974);
and U9733 (N_9733,N_7067,N_6178);
or U9734 (N_9734,N_5557,N_6279);
xnor U9735 (N_9735,N_5412,N_5575);
nand U9736 (N_9736,N_7497,N_5093);
nor U9737 (N_9737,N_5475,N_7355);
nor U9738 (N_9738,N_6921,N_5591);
and U9739 (N_9739,N_6567,N_5698);
xor U9740 (N_9740,N_7416,N_5445);
or U9741 (N_9741,N_5149,N_6676);
and U9742 (N_9742,N_6712,N_6282);
or U9743 (N_9743,N_6752,N_6627);
or U9744 (N_9744,N_5439,N_6624);
and U9745 (N_9745,N_6024,N_5083);
nand U9746 (N_9746,N_5039,N_6991);
xnor U9747 (N_9747,N_6355,N_5403);
nor U9748 (N_9748,N_6088,N_7238);
or U9749 (N_9749,N_6948,N_6207);
nand U9750 (N_9750,N_5086,N_7241);
or U9751 (N_9751,N_6120,N_5679);
or U9752 (N_9752,N_6441,N_5224);
or U9753 (N_9753,N_5873,N_6035);
nand U9754 (N_9754,N_5325,N_5583);
nor U9755 (N_9755,N_5576,N_6569);
or U9756 (N_9756,N_5613,N_5858);
nand U9757 (N_9757,N_7060,N_5259);
or U9758 (N_9758,N_5528,N_5342);
and U9759 (N_9759,N_6300,N_6567);
and U9760 (N_9760,N_6413,N_7210);
nand U9761 (N_9761,N_6744,N_7381);
nand U9762 (N_9762,N_7101,N_5256);
or U9763 (N_9763,N_5570,N_6693);
xor U9764 (N_9764,N_5473,N_5391);
nand U9765 (N_9765,N_6953,N_7217);
and U9766 (N_9766,N_5046,N_5528);
xnor U9767 (N_9767,N_7417,N_6930);
or U9768 (N_9768,N_5169,N_7189);
nor U9769 (N_9769,N_5551,N_6735);
and U9770 (N_9770,N_7370,N_7067);
or U9771 (N_9771,N_5052,N_5839);
xnor U9772 (N_9772,N_6794,N_7221);
nand U9773 (N_9773,N_5838,N_5211);
xor U9774 (N_9774,N_6723,N_6098);
nor U9775 (N_9775,N_6974,N_7372);
nand U9776 (N_9776,N_6793,N_5285);
nor U9777 (N_9777,N_7298,N_5359);
and U9778 (N_9778,N_6309,N_7227);
xor U9779 (N_9779,N_5045,N_6975);
or U9780 (N_9780,N_6883,N_6000);
nor U9781 (N_9781,N_5370,N_5640);
or U9782 (N_9782,N_5636,N_7303);
nor U9783 (N_9783,N_7183,N_5147);
or U9784 (N_9784,N_5055,N_6895);
nand U9785 (N_9785,N_5194,N_5078);
or U9786 (N_9786,N_5751,N_5486);
nor U9787 (N_9787,N_5690,N_7199);
nand U9788 (N_9788,N_7194,N_6518);
and U9789 (N_9789,N_7145,N_5751);
or U9790 (N_9790,N_6834,N_5321);
or U9791 (N_9791,N_5474,N_7443);
and U9792 (N_9792,N_7092,N_5950);
nor U9793 (N_9793,N_6965,N_7421);
xnor U9794 (N_9794,N_6030,N_6139);
or U9795 (N_9795,N_6497,N_6035);
nand U9796 (N_9796,N_5169,N_7383);
xnor U9797 (N_9797,N_5184,N_7090);
or U9798 (N_9798,N_6102,N_6813);
nand U9799 (N_9799,N_5933,N_6463);
xor U9800 (N_9800,N_5655,N_5882);
and U9801 (N_9801,N_5692,N_5364);
nor U9802 (N_9802,N_5898,N_5202);
nand U9803 (N_9803,N_6574,N_7124);
or U9804 (N_9804,N_5451,N_6199);
and U9805 (N_9805,N_6903,N_7168);
nor U9806 (N_9806,N_5841,N_6221);
or U9807 (N_9807,N_6704,N_5045);
and U9808 (N_9808,N_6983,N_7404);
nor U9809 (N_9809,N_7000,N_6582);
nor U9810 (N_9810,N_7349,N_6523);
and U9811 (N_9811,N_7368,N_7078);
xor U9812 (N_9812,N_6437,N_5609);
nand U9813 (N_9813,N_6861,N_6101);
or U9814 (N_9814,N_5406,N_6354);
and U9815 (N_9815,N_7357,N_7047);
or U9816 (N_9816,N_5522,N_7158);
or U9817 (N_9817,N_6254,N_7228);
and U9818 (N_9818,N_5313,N_5609);
nor U9819 (N_9819,N_5850,N_7072);
nor U9820 (N_9820,N_5867,N_6782);
or U9821 (N_9821,N_7185,N_6708);
and U9822 (N_9822,N_6574,N_6556);
or U9823 (N_9823,N_6900,N_7240);
nand U9824 (N_9824,N_5875,N_7467);
xnor U9825 (N_9825,N_6259,N_5946);
and U9826 (N_9826,N_5361,N_5991);
nor U9827 (N_9827,N_5269,N_5926);
and U9828 (N_9828,N_5923,N_7302);
and U9829 (N_9829,N_6024,N_5016);
nor U9830 (N_9830,N_5918,N_6962);
nor U9831 (N_9831,N_7361,N_6651);
and U9832 (N_9832,N_6552,N_5712);
nor U9833 (N_9833,N_6207,N_6705);
nand U9834 (N_9834,N_7120,N_5461);
and U9835 (N_9835,N_7482,N_5767);
nor U9836 (N_9836,N_5726,N_6916);
or U9837 (N_9837,N_6166,N_6535);
or U9838 (N_9838,N_6575,N_6725);
nor U9839 (N_9839,N_7456,N_5176);
nand U9840 (N_9840,N_5257,N_6302);
xor U9841 (N_9841,N_5124,N_7288);
nor U9842 (N_9842,N_6088,N_6115);
and U9843 (N_9843,N_6776,N_6810);
and U9844 (N_9844,N_7091,N_5553);
nor U9845 (N_9845,N_6475,N_7237);
nor U9846 (N_9846,N_6894,N_6117);
or U9847 (N_9847,N_6338,N_7337);
nand U9848 (N_9848,N_6383,N_5301);
nand U9849 (N_9849,N_5316,N_7384);
nor U9850 (N_9850,N_7180,N_5081);
nor U9851 (N_9851,N_6006,N_6980);
and U9852 (N_9852,N_5721,N_5201);
nand U9853 (N_9853,N_7352,N_6982);
nor U9854 (N_9854,N_5341,N_7182);
nand U9855 (N_9855,N_7408,N_5880);
nand U9856 (N_9856,N_5606,N_7253);
and U9857 (N_9857,N_7319,N_6051);
nand U9858 (N_9858,N_6377,N_6270);
nand U9859 (N_9859,N_6007,N_6277);
or U9860 (N_9860,N_7309,N_6995);
and U9861 (N_9861,N_5888,N_5105);
nand U9862 (N_9862,N_5238,N_5146);
nor U9863 (N_9863,N_5067,N_6893);
nor U9864 (N_9864,N_7115,N_6532);
and U9865 (N_9865,N_6615,N_6592);
and U9866 (N_9866,N_6340,N_7359);
or U9867 (N_9867,N_5827,N_6796);
nor U9868 (N_9868,N_6902,N_5168);
or U9869 (N_9869,N_6075,N_5145);
nor U9870 (N_9870,N_5301,N_5739);
nor U9871 (N_9871,N_6548,N_6850);
or U9872 (N_9872,N_5386,N_6694);
nor U9873 (N_9873,N_7254,N_5642);
nor U9874 (N_9874,N_7042,N_5269);
or U9875 (N_9875,N_6588,N_7080);
nand U9876 (N_9876,N_7439,N_5289);
nor U9877 (N_9877,N_6070,N_6549);
or U9878 (N_9878,N_6804,N_6747);
and U9879 (N_9879,N_6248,N_6590);
nor U9880 (N_9880,N_7126,N_5333);
nand U9881 (N_9881,N_6475,N_6358);
and U9882 (N_9882,N_6164,N_6406);
nor U9883 (N_9883,N_6311,N_6095);
nand U9884 (N_9884,N_5472,N_5467);
xor U9885 (N_9885,N_5433,N_5692);
and U9886 (N_9886,N_5387,N_6176);
xor U9887 (N_9887,N_6056,N_7184);
or U9888 (N_9888,N_5086,N_6710);
nand U9889 (N_9889,N_5106,N_5616);
or U9890 (N_9890,N_5404,N_5402);
and U9891 (N_9891,N_5415,N_6463);
nand U9892 (N_9892,N_5006,N_7376);
nand U9893 (N_9893,N_7400,N_7025);
nor U9894 (N_9894,N_6956,N_6601);
and U9895 (N_9895,N_5656,N_6932);
and U9896 (N_9896,N_6422,N_5096);
and U9897 (N_9897,N_7165,N_6896);
nor U9898 (N_9898,N_5173,N_5691);
nand U9899 (N_9899,N_6064,N_5092);
or U9900 (N_9900,N_6021,N_7437);
nor U9901 (N_9901,N_6203,N_5972);
nand U9902 (N_9902,N_5567,N_7256);
nand U9903 (N_9903,N_6902,N_7427);
xor U9904 (N_9904,N_6159,N_5013);
nor U9905 (N_9905,N_5272,N_5592);
nor U9906 (N_9906,N_5906,N_6041);
nand U9907 (N_9907,N_5726,N_6350);
nand U9908 (N_9908,N_6126,N_6943);
or U9909 (N_9909,N_7254,N_6468);
nor U9910 (N_9910,N_7178,N_6963);
nand U9911 (N_9911,N_6358,N_7252);
or U9912 (N_9912,N_5023,N_6357);
nand U9913 (N_9913,N_6254,N_6377);
nand U9914 (N_9914,N_6682,N_5112);
or U9915 (N_9915,N_7092,N_5683);
xnor U9916 (N_9916,N_7080,N_7132);
nor U9917 (N_9917,N_6336,N_7396);
and U9918 (N_9918,N_5544,N_6333);
nand U9919 (N_9919,N_7395,N_7057);
nor U9920 (N_9920,N_5498,N_5541);
nor U9921 (N_9921,N_5418,N_5185);
or U9922 (N_9922,N_6372,N_6592);
nand U9923 (N_9923,N_5668,N_5359);
nand U9924 (N_9924,N_6739,N_5560);
nand U9925 (N_9925,N_6085,N_5359);
or U9926 (N_9926,N_5570,N_6310);
or U9927 (N_9927,N_5975,N_6710);
nand U9928 (N_9928,N_6350,N_6184);
nor U9929 (N_9929,N_5606,N_6198);
and U9930 (N_9930,N_5029,N_6939);
nand U9931 (N_9931,N_7106,N_6489);
or U9932 (N_9932,N_6629,N_5159);
and U9933 (N_9933,N_6602,N_5344);
nor U9934 (N_9934,N_5124,N_5980);
or U9935 (N_9935,N_6217,N_6826);
nand U9936 (N_9936,N_5753,N_5269);
nand U9937 (N_9937,N_6301,N_6321);
xor U9938 (N_9938,N_6772,N_6462);
nand U9939 (N_9939,N_5683,N_6194);
and U9940 (N_9940,N_7025,N_6536);
or U9941 (N_9941,N_6636,N_6951);
nand U9942 (N_9942,N_7285,N_6500);
nor U9943 (N_9943,N_6604,N_7275);
nand U9944 (N_9944,N_5281,N_5913);
and U9945 (N_9945,N_5189,N_7216);
nand U9946 (N_9946,N_6263,N_6319);
nand U9947 (N_9947,N_6257,N_7088);
or U9948 (N_9948,N_6239,N_6994);
xnor U9949 (N_9949,N_6550,N_7431);
nor U9950 (N_9950,N_6549,N_6517);
nand U9951 (N_9951,N_5503,N_6947);
and U9952 (N_9952,N_5351,N_5812);
or U9953 (N_9953,N_6668,N_7145);
and U9954 (N_9954,N_6324,N_6861);
nand U9955 (N_9955,N_6108,N_6126);
nor U9956 (N_9956,N_5973,N_6344);
and U9957 (N_9957,N_7499,N_6757);
or U9958 (N_9958,N_7498,N_6881);
or U9959 (N_9959,N_7492,N_6038);
xnor U9960 (N_9960,N_5757,N_5534);
nand U9961 (N_9961,N_5379,N_6217);
and U9962 (N_9962,N_5013,N_6558);
xor U9963 (N_9963,N_6858,N_6813);
and U9964 (N_9964,N_6020,N_7004);
and U9965 (N_9965,N_7120,N_5670);
nor U9966 (N_9966,N_6608,N_6524);
or U9967 (N_9967,N_6168,N_6962);
and U9968 (N_9968,N_6689,N_6327);
nor U9969 (N_9969,N_6814,N_5274);
or U9970 (N_9970,N_5061,N_5462);
nand U9971 (N_9971,N_5738,N_5595);
and U9972 (N_9972,N_5795,N_5394);
or U9973 (N_9973,N_5570,N_7174);
and U9974 (N_9974,N_5478,N_5570);
nor U9975 (N_9975,N_6041,N_5724);
and U9976 (N_9976,N_6989,N_5074);
xnor U9977 (N_9977,N_6216,N_6817);
nor U9978 (N_9978,N_7153,N_6849);
or U9979 (N_9979,N_5295,N_5819);
nor U9980 (N_9980,N_5879,N_5057);
and U9981 (N_9981,N_5037,N_5640);
nor U9982 (N_9982,N_5750,N_7219);
or U9983 (N_9983,N_6829,N_6167);
and U9984 (N_9984,N_5562,N_7115);
and U9985 (N_9985,N_5506,N_5219);
nand U9986 (N_9986,N_6144,N_6047);
or U9987 (N_9987,N_7221,N_5903);
nand U9988 (N_9988,N_6142,N_5680);
and U9989 (N_9989,N_5333,N_7032);
xor U9990 (N_9990,N_7496,N_6795);
or U9991 (N_9991,N_7473,N_6842);
and U9992 (N_9992,N_6060,N_6907);
and U9993 (N_9993,N_5160,N_5950);
and U9994 (N_9994,N_6316,N_5964);
and U9995 (N_9995,N_5476,N_5213);
or U9996 (N_9996,N_7044,N_6248);
or U9997 (N_9997,N_6392,N_6104);
nand U9998 (N_9998,N_5797,N_6349);
and U9999 (N_9999,N_6922,N_5152);
and UO_0 (O_0,N_9728,N_8948);
or UO_1 (O_1,N_7916,N_9681);
nand UO_2 (O_2,N_8981,N_8430);
nor UO_3 (O_3,N_8201,N_9969);
and UO_4 (O_4,N_8960,N_8015);
nor UO_5 (O_5,N_9921,N_8266);
xnor UO_6 (O_6,N_7563,N_8265);
nor UO_7 (O_7,N_8256,N_8327);
nor UO_8 (O_8,N_7997,N_9642);
xnor UO_9 (O_9,N_9632,N_9889);
nand UO_10 (O_10,N_7522,N_9264);
and UO_11 (O_11,N_9283,N_9291);
nor UO_12 (O_12,N_8363,N_9601);
nand UO_13 (O_13,N_9797,N_9347);
nor UO_14 (O_14,N_7506,N_9688);
nand UO_15 (O_15,N_8945,N_8768);
and UO_16 (O_16,N_8096,N_9447);
nor UO_17 (O_17,N_8445,N_8598);
nor UO_18 (O_18,N_7878,N_9277);
nand UO_19 (O_19,N_9184,N_8062);
nand UO_20 (O_20,N_9121,N_8518);
and UO_21 (O_21,N_7852,N_8980);
nand UO_22 (O_22,N_9458,N_9329);
nand UO_23 (O_23,N_8339,N_8423);
nor UO_24 (O_24,N_8920,N_9285);
or UO_25 (O_25,N_7704,N_8408);
and UO_26 (O_26,N_9685,N_8725);
nand UO_27 (O_27,N_7682,N_9359);
nor UO_28 (O_28,N_8975,N_8837);
nand UO_29 (O_29,N_9843,N_8668);
nor UO_30 (O_30,N_8319,N_9788);
or UO_31 (O_31,N_8578,N_9868);
or UO_32 (O_32,N_9030,N_9813);
or UO_33 (O_33,N_7595,N_8144);
and UO_34 (O_34,N_9314,N_8692);
or UO_35 (O_35,N_8754,N_7600);
nor UO_36 (O_36,N_9172,N_7592);
or UO_37 (O_37,N_7926,N_9647);
and UO_38 (O_38,N_9483,N_9327);
nor UO_39 (O_39,N_8588,N_9017);
or UO_40 (O_40,N_8324,N_9488);
nand UO_41 (O_41,N_9444,N_8184);
or UO_42 (O_42,N_8821,N_8099);
and UO_43 (O_43,N_9584,N_7728);
and UO_44 (O_44,N_7778,N_8384);
and UO_45 (O_45,N_9323,N_8331);
nor UO_46 (O_46,N_9667,N_8538);
or UO_47 (O_47,N_8603,N_9846);
nand UO_48 (O_48,N_9226,N_8621);
and UO_49 (O_49,N_7591,N_8858);
or UO_50 (O_50,N_8278,N_9271);
nand UO_51 (O_51,N_8115,N_7849);
or UO_52 (O_52,N_9893,N_8541);
nand UO_53 (O_53,N_9666,N_8910);
and UO_54 (O_54,N_9441,N_9579);
xor UO_55 (O_55,N_8977,N_7884);
xnor UO_56 (O_56,N_7869,N_7877);
and UO_57 (O_57,N_9103,N_9554);
nor UO_58 (O_58,N_8646,N_8932);
and UO_59 (O_59,N_7891,N_9151);
nor UO_60 (O_60,N_8964,N_7706);
nor UO_61 (O_61,N_9982,N_8552);
or UO_62 (O_62,N_7765,N_9125);
nand UO_63 (O_63,N_7768,N_8593);
xor UO_64 (O_64,N_7590,N_8494);
nand UO_65 (O_65,N_9598,N_9400);
nor UO_66 (O_66,N_7774,N_8466);
or UO_67 (O_67,N_8416,N_8811);
and UO_68 (O_68,N_9092,N_9951);
nor UO_69 (O_69,N_9454,N_9787);
nor UO_70 (O_70,N_9036,N_8205);
nand UO_71 (O_71,N_7629,N_8010);
nand UO_72 (O_72,N_8017,N_9001);
and UO_73 (O_73,N_9418,N_9957);
xnor UO_74 (O_74,N_9145,N_9491);
and UO_75 (O_75,N_9257,N_9494);
and UO_76 (O_76,N_9716,N_7638);
and UO_77 (O_77,N_8845,N_8746);
nor UO_78 (O_78,N_8338,N_8097);
nor UO_79 (O_79,N_9741,N_8889);
xnor UO_80 (O_80,N_9452,N_8671);
and UO_81 (O_81,N_7988,N_8897);
nand UO_82 (O_82,N_8159,N_8002);
and UO_83 (O_83,N_8310,N_8657);
and UO_84 (O_84,N_7707,N_9095);
nor UO_85 (O_85,N_8642,N_9777);
or UO_86 (O_86,N_9504,N_7539);
nand UO_87 (O_87,N_7750,N_8230);
nor UO_88 (O_88,N_9159,N_8069);
nor UO_89 (O_89,N_8297,N_9194);
xnor UO_90 (O_90,N_8501,N_9398);
nor UO_91 (O_91,N_9428,N_9828);
nand UO_92 (O_92,N_9841,N_8576);
xor UO_93 (O_93,N_9793,N_9721);
xnor UO_94 (O_94,N_8506,N_9344);
nand UO_95 (O_95,N_9305,N_8027);
nor UO_96 (O_96,N_8417,N_9438);
and UO_97 (O_97,N_8713,N_9358);
nand UO_98 (O_98,N_8622,N_9161);
and UO_99 (O_99,N_8880,N_9365);
nor UO_100 (O_100,N_8838,N_9354);
xnor UO_101 (O_101,N_8227,N_9590);
or UO_102 (O_102,N_9414,N_8790);
xnor UO_103 (O_103,N_8903,N_9191);
nand UO_104 (O_104,N_9244,N_8074);
nor UO_105 (O_105,N_9656,N_7520);
or UO_106 (O_106,N_7669,N_8413);
nand UO_107 (O_107,N_9732,N_9152);
and UO_108 (O_108,N_9867,N_8833);
or UO_109 (O_109,N_9403,N_8586);
or UO_110 (O_110,N_8401,N_7611);
nand UO_111 (O_111,N_8309,N_8647);
and UO_112 (O_112,N_7566,N_9566);
nand UO_113 (O_113,N_8641,N_7910);
nor UO_114 (O_114,N_9018,N_8885);
nand UO_115 (O_115,N_8128,N_8674);
and UO_116 (O_116,N_9411,N_7685);
nand UO_117 (O_117,N_9267,N_8599);
nand UO_118 (O_118,N_8864,N_7741);
or UO_119 (O_119,N_7537,N_8127);
xnor UO_120 (O_120,N_8420,N_8274);
xor UO_121 (O_121,N_8037,N_8720);
or UO_122 (O_122,N_8276,N_8103);
nor UO_123 (O_123,N_8721,N_9545);
or UO_124 (O_124,N_8066,N_8286);
or UO_125 (O_125,N_9730,N_8165);
nor UO_126 (O_126,N_8996,N_9724);
and UO_127 (O_127,N_8448,N_9210);
nor UO_128 (O_128,N_8602,N_9409);
xor UO_129 (O_129,N_9890,N_9228);
xor UO_130 (O_130,N_9224,N_7676);
xor UO_131 (O_131,N_8369,N_8503);
nand UO_132 (O_132,N_8895,N_7727);
xor UO_133 (O_133,N_7536,N_9179);
and UO_134 (O_134,N_8712,N_8151);
nand UO_135 (O_135,N_8508,N_8601);
and UO_136 (O_136,N_9102,N_8481);
nand UO_137 (O_137,N_8308,N_8397);
nand UO_138 (O_138,N_8925,N_9532);
and UO_139 (O_139,N_8616,N_8209);
and UO_140 (O_140,N_8477,N_8400);
or UO_141 (O_141,N_8831,N_8370);
nor UO_142 (O_142,N_9214,N_8167);
or UO_143 (O_143,N_8939,N_9669);
nand UO_144 (O_144,N_8968,N_8618);
and UO_145 (O_145,N_9789,N_9809);
or UO_146 (O_146,N_9419,N_9778);
and UO_147 (O_147,N_9343,N_7799);
nor UO_148 (O_148,N_9235,N_9000);
or UO_149 (O_149,N_8741,N_8564);
nor UO_150 (O_150,N_9881,N_8187);
nand UO_151 (O_151,N_9934,N_9692);
or UO_152 (O_152,N_9586,N_9613);
and UO_153 (O_153,N_9231,N_8287);
and UO_154 (O_154,N_8590,N_7931);
xnor UO_155 (O_155,N_9296,N_9963);
or UO_156 (O_156,N_9106,N_9582);
or UO_157 (O_157,N_8143,N_8489);
nor UO_158 (O_158,N_9312,N_9311);
and UO_159 (O_159,N_9187,N_8665);
and UO_160 (O_160,N_8553,N_7675);
xor UO_161 (O_161,N_9094,N_9148);
and UO_162 (O_162,N_9623,N_8325);
or UO_163 (O_163,N_8181,N_9236);
and UO_164 (O_164,N_9211,N_9333);
or UO_165 (O_165,N_9270,N_8299);
nand UO_166 (O_166,N_8842,N_9596);
or UO_167 (O_167,N_9895,N_9936);
and UO_168 (O_168,N_7881,N_7882);
nor UO_169 (O_169,N_7726,N_9239);
nor UO_170 (O_170,N_8407,N_8463);
nor UO_171 (O_171,N_9370,N_7983);
or UO_172 (O_172,N_9022,N_8807);
nand UO_173 (O_173,N_7565,N_7989);
or UO_174 (O_174,N_8163,N_8966);
and UO_175 (O_175,N_9091,N_9213);
and UO_176 (O_176,N_8557,N_9521);
xor UO_177 (O_177,N_8937,N_8342);
or UO_178 (O_178,N_7656,N_9743);
nand UO_179 (O_179,N_7894,N_9644);
nor UO_180 (O_180,N_8488,N_9759);
xnor UO_181 (O_181,N_9142,N_8844);
xnor UO_182 (O_182,N_8282,N_7867);
nand UO_183 (O_183,N_7578,N_8350);
nor UO_184 (O_184,N_8328,N_9051);
xor UO_185 (O_185,N_9926,N_8472);
or UO_186 (O_186,N_7545,N_8186);
and UO_187 (O_187,N_8058,N_8882);
or UO_188 (O_188,N_9407,N_8753);
and UO_189 (O_189,N_8149,N_8125);
or UO_190 (O_190,N_7821,N_8063);
or UO_191 (O_191,N_7942,N_7526);
nand UO_192 (O_192,N_9648,N_7610);
nor UO_193 (O_193,N_7571,N_8877);
or UO_194 (O_194,N_8653,N_9563);
and UO_195 (O_195,N_9129,N_8418);
xnor UO_196 (O_196,N_8734,N_7670);
nand UO_197 (O_197,N_8778,N_9351);
or UO_198 (O_198,N_9715,N_7813);
or UO_199 (O_199,N_8531,N_9907);
xor UO_200 (O_200,N_7836,N_8574);
or UO_201 (O_201,N_7885,N_9363);
xor UO_202 (O_202,N_7992,N_9627);
and UO_203 (O_203,N_9386,N_8215);
and UO_204 (O_204,N_8344,N_9469);
nor UO_205 (O_205,N_8801,N_9948);
or UO_206 (O_206,N_8800,N_8750);
nand UO_207 (O_207,N_9261,N_9978);
nand UO_208 (O_208,N_8168,N_7966);
and UO_209 (O_209,N_8556,N_8343);
or UO_210 (O_210,N_9511,N_9466);
nand UO_211 (O_211,N_8815,N_8701);
nand UO_212 (O_212,N_9153,N_9342);
or UO_213 (O_213,N_9147,N_9420);
and UO_214 (O_214,N_8498,N_7691);
nor UO_215 (O_215,N_9256,N_8268);
or UO_216 (O_216,N_7513,N_8060);
nand UO_217 (O_217,N_8927,N_9076);
and UO_218 (O_218,N_8303,N_8345);
nor UO_219 (O_219,N_9714,N_7722);
xor UO_220 (O_220,N_9026,N_9780);
nor UO_221 (O_221,N_7961,N_9585);
or UO_222 (O_222,N_7857,N_9149);
or UO_223 (O_223,N_9263,N_9625);
and UO_224 (O_224,N_7607,N_8860);
nand UO_225 (O_225,N_7860,N_8982);
xor UO_226 (O_226,N_9388,N_9043);
nand UO_227 (O_227,N_7844,N_8210);
and UO_228 (O_228,N_9423,N_8043);
nor UO_229 (O_229,N_9044,N_7964);
or UO_230 (O_230,N_9081,N_9249);
nor UO_231 (O_231,N_7651,N_8051);
nand UO_232 (O_232,N_7808,N_7646);
nor UO_233 (O_233,N_8949,N_9064);
xor UO_234 (O_234,N_8804,N_9706);
xnor UO_235 (O_235,N_7658,N_8719);
or UO_236 (O_236,N_8441,N_9530);
xor UO_237 (O_237,N_8198,N_8562);
nor UO_238 (O_238,N_7889,N_9665);
nor UO_239 (O_239,N_9718,N_8172);
and UO_240 (O_240,N_9956,N_9056);
nor UO_241 (O_241,N_8504,N_7608);
and UO_242 (O_242,N_7922,N_9009);
nand UO_243 (O_243,N_9492,N_9562);
nor UO_244 (O_244,N_8623,N_8783);
and UO_245 (O_245,N_9729,N_8519);
or UO_246 (O_246,N_9550,N_9535);
nand UO_247 (O_247,N_9130,N_9254);
nand UO_248 (O_248,N_9804,N_8579);
or UO_249 (O_249,N_8496,N_9624);
xnor UO_250 (O_250,N_8722,N_7906);
and UO_251 (O_251,N_8180,N_8164);
and UO_252 (O_252,N_8404,N_7825);
xnor UO_253 (O_253,N_9415,N_8883);
nor UO_254 (O_254,N_9731,N_8253);
nor UO_255 (O_255,N_8469,N_8204);
nand UO_256 (O_256,N_8994,N_9294);
and UO_257 (O_257,N_8524,N_8946);
or UO_258 (O_258,N_8707,N_7796);
xor UO_259 (O_259,N_7625,N_8262);
and UO_260 (O_260,N_9357,N_9918);
xnor UO_261 (O_261,N_8374,N_8849);
and UO_262 (O_262,N_9164,N_9872);
and UO_263 (O_263,N_9192,N_8615);
nor UO_264 (O_264,N_7939,N_9929);
and UO_265 (O_265,N_9424,N_7725);
and UO_266 (O_266,N_8312,N_8570);
xor UO_267 (O_267,N_8486,N_8726);
and UO_268 (O_268,N_8183,N_9942);
nand UO_269 (O_269,N_7822,N_9541);
or UO_270 (O_270,N_8305,N_8161);
or UO_271 (O_271,N_8360,N_7540);
nand UO_272 (O_272,N_8951,N_8824);
and UO_273 (O_273,N_8777,N_8738);
nor UO_274 (O_274,N_8387,N_9068);
nor UO_275 (O_275,N_7841,N_9542);
nor UO_276 (O_276,N_9313,N_7810);
or UO_277 (O_277,N_9353,N_9992);
nand UO_278 (O_278,N_8089,N_7950);
or UO_279 (O_279,N_8026,N_9241);
xnor UO_280 (O_280,N_7978,N_8639);
and UO_281 (O_281,N_8853,N_8396);
xor UO_282 (O_282,N_9324,N_8427);
or UO_283 (O_283,N_8866,N_9046);
xor UO_284 (O_284,N_8359,N_9654);
or UO_285 (O_285,N_8390,N_8351);
or UO_286 (O_286,N_9433,N_8704);
nor UO_287 (O_287,N_8697,N_7954);
and UO_288 (O_288,N_7688,N_8747);
or UO_289 (O_289,N_8600,N_9421);
or UO_290 (O_290,N_8545,N_8675);
and UO_291 (O_291,N_8064,N_9537);
or UO_292 (O_292,N_7554,N_9474);
and UO_293 (O_293,N_7692,N_8499);
and UO_294 (O_294,N_9199,N_9886);
or UO_295 (O_295,N_7759,N_9917);
nor UO_296 (O_296,N_9186,N_8284);
and UO_297 (O_297,N_9004,N_9355);
nor UO_298 (O_298,N_9856,N_7957);
nor UO_299 (O_299,N_7987,N_8611);
nand UO_300 (O_300,N_8965,N_8513);
nand UO_301 (O_301,N_8904,N_8008);
nor UO_302 (O_302,N_7873,N_7555);
xnor UO_303 (O_303,N_8688,N_7662);
nor UO_304 (O_304,N_8323,N_8162);
and UO_305 (O_305,N_9811,N_8689);
nor UO_306 (O_306,N_8533,N_7757);
nor UO_307 (O_307,N_8567,N_9146);
or UO_308 (O_308,N_8317,N_9885);
xor UO_309 (O_309,N_9749,N_9442);
and UO_310 (O_310,N_7960,N_8859);
or UO_311 (O_311,N_8648,N_8993);
or UO_312 (O_312,N_7758,N_8592);
and UO_313 (O_313,N_8059,N_9097);
nor UO_314 (O_314,N_8534,N_8666);
nand UO_315 (O_315,N_8435,N_8986);
or UO_316 (O_316,N_7556,N_7667);
nand UO_317 (O_317,N_9059,N_9085);
or UO_318 (O_318,N_9561,N_7781);
or UO_319 (O_319,N_9968,N_8727);
nor UO_320 (O_320,N_8029,N_7708);
and UO_321 (O_321,N_9538,N_8225);
or UO_322 (O_322,N_7888,N_7524);
xor UO_323 (O_323,N_8915,N_8810);
xnor UO_324 (O_324,N_9912,N_8200);
and UO_325 (O_325,N_7854,N_7562);
xnor UO_326 (O_326,N_8879,N_8818);
nand UO_327 (O_327,N_8480,N_9527);
nor UO_328 (O_328,N_8129,N_9865);
and UO_329 (O_329,N_7684,N_8065);
or UO_330 (O_330,N_7868,N_9633);
nand UO_331 (O_331,N_7823,N_9988);
and UO_332 (O_332,N_9998,N_7752);
and UO_333 (O_333,N_8379,N_9941);
and UO_334 (O_334,N_9659,N_9924);
nor UO_335 (O_335,N_9482,N_9110);
xor UO_336 (O_336,N_9171,N_9237);
and UO_337 (O_337,N_8054,N_7927);
nand UO_338 (O_338,N_8763,N_8020);
xor UO_339 (O_339,N_9836,N_8460);
or UO_340 (O_340,N_8145,N_9696);
and UO_341 (O_341,N_8502,N_7529);
or UO_342 (O_342,N_8281,N_9600);
nand UO_343 (O_343,N_9587,N_9638);
nor UO_344 (O_344,N_8854,N_8042);
or UO_345 (O_345,N_9168,N_9795);
and UO_346 (O_346,N_9835,N_9539);
xnor UO_347 (O_347,N_9077,N_7642);
or UO_348 (O_348,N_8431,N_9015);
nand UO_349 (O_349,N_8606,N_7890);
and UO_350 (O_350,N_8523,N_7696);
nand UO_351 (O_351,N_7621,N_7679);
or UO_352 (O_352,N_8153,N_8914);
and UO_353 (O_353,N_9364,N_8375);
nor UO_354 (O_354,N_8073,N_9838);
xor UO_355 (O_355,N_7784,N_9297);
nor UO_356 (O_356,N_8724,N_9269);
nor UO_357 (O_357,N_9485,N_9593);
or UO_358 (O_358,N_9185,N_9552);
and UO_359 (O_359,N_8941,N_8241);
nor UO_360 (O_360,N_8244,N_9122);
nor UO_361 (O_361,N_8372,N_9162);
nor UO_362 (O_362,N_8921,N_9708);
nand UO_363 (O_363,N_7937,N_8613);
nand UO_364 (O_364,N_7870,N_9575);
and UO_365 (O_365,N_9476,N_9352);
nand UO_366 (O_366,N_7904,N_8425);
or UO_367 (O_367,N_8437,N_8710);
xnor UO_368 (O_368,N_7716,N_7598);
nand UO_369 (O_369,N_9246,N_9093);
nor UO_370 (O_370,N_9193,N_9878);
nand UO_371 (O_371,N_8540,N_9750);
xnor UO_372 (O_372,N_8549,N_7570);
or UO_373 (O_373,N_9014,N_9338);
nand UO_374 (O_374,N_9857,N_9111);
and UO_375 (O_375,N_7970,N_8467);
nor UO_376 (O_376,N_9024,N_7635);
nor UO_377 (O_377,N_9131,N_8148);
and UO_378 (O_378,N_9242,N_7971);
nor UO_379 (O_379,N_8944,N_9183);
nand UO_380 (O_380,N_7816,N_8371);
and UO_381 (O_381,N_8507,N_9489);
nor UO_382 (O_382,N_8095,N_9981);
or UO_383 (O_383,N_7948,N_8661);
nand UO_384 (O_384,N_7875,N_8236);
nor UO_385 (O_385,N_8597,N_8764);
nor UO_386 (O_386,N_7895,N_8971);
nand UO_387 (O_387,N_7990,N_8112);
or UO_388 (O_388,N_9742,N_9635);
nand UO_389 (O_389,N_9175,N_7933);
and UO_390 (O_390,N_8812,N_9058);
and UO_391 (O_391,N_7541,N_8684);
nor UO_392 (O_392,N_8544,N_7547);
nor UO_393 (O_393,N_9913,N_8220);
or UO_394 (O_394,N_7649,N_8334);
or UO_395 (O_395,N_9548,N_8723);
xnor UO_396 (O_396,N_8584,N_7531);
and UO_397 (O_397,N_8890,N_8202);
nor UO_398 (O_398,N_8239,N_8156);
and UO_399 (O_399,N_9767,N_7501);
xnor UO_400 (O_400,N_9457,N_7782);
nand UO_401 (O_401,N_8814,N_9345);
and UO_402 (O_402,N_8667,N_8291);
nor UO_403 (O_403,N_9176,N_8378);
or UO_404 (O_404,N_8805,N_9565);
or UO_405 (O_405,N_8650,N_9021);
nand UO_406 (O_406,N_9348,N_9816);
xnor UO_407 (O_407,N_8774,N_9155);
nand UO_408 (O_408,N_9544,N_7930);
and UO_409 (O_409,N_8012,N_9126);
and UO_410 (O_410,N_8388,N_9873);
and UO_411 (O_411,N_8031,N_8123);
and UO_412 (O_412,N_8514,N_7747);
nand UO_413 (O_413,N_9188,N_8940);
nor UO_414 (O_414,N_9072,N_7703);
and UO_415 (O_415,N_9919,N_9053);
or UO_416 (O_416,N_9687,N_8424);
xor UO_417 (O_417,N_9528,N_8683);
or UO_418 (O_418,N_8876,N_7798);
or UO_419 (O_419,N_9299,N_7559);
and UO_420 (O_420,N_9916,N_8687);
nor UO_421 (O_421,N_9914,N_7773);
and UO_422 (O_422,N_8536,N_9276);
nand UO_423 (O_423,N_8314,N_9067);
or UO_424 (O_424,N_7697,N_7709);
xor UO_425 (O_425,N_9570,N_8240);
nor UO_426 (O_426,N_8873,N_7949);
xnor UO_427 (O_427,N_9707,N_9499);
nor UO_428 (O_428,N_7612,N_9055);
nor UO_429 (O_429,N_8742,N_9506);
or UO_430 (O_430,N_7811,N_8452);
or UO_431 (O_431,N_9380,N_7858);
and UO_432 (O_432,N_7627,N_7780);
and UO_433 (O_433,N_9909,N_9603);
nand UO_434 (O_434,N_9098,N_8884);
and UO_435 (O_435,N_7523,N_7623);
xnor UO_436 (O_436,N_8547,N_8373);
or UO_437 (O_437,N_9088,N_8476);
or UO_438 (O_438,N_9831,N_7929);
nand UO_439 (O_439,N_9472,N_9115);
nor UO_440 (O_440,N_7947,N_9005);
and UO_441 (O_441,N_8663,N_8141);
or UO_442 (O_442,N_9473,N_9496);
and UO_443 (O_443,N_8875,N_9855);
nor UO_444 (O_444,N_8119,N_9949);
and UO_445 (O_445,N_8694,N_8298);
and UO_446 (O_446,N_9066,N_9705);
nor UO_447 (O_447,N_9134,N_7505);
and UO_448 (O_448,N_9215,N_8526);
and UO_449 (O_449,N_8108,N_8656);
nor UO_450 (O_450,N_8436,N_9822);
nor UO_451 (O_451,N_9576,N_9771);
nor UO_452 (O_452,N_7665,N_9533);
nor UO_453 (O_453,N_8454,N_9950);
or UO_454 (O_454,N_7982,N_8208);
or UO_455 (O_455,N_7624,N_8958);
or UO_456 (O_456,N_8772,N_8254);
or UO_457 (O_457,N_7995,N_7981);
nand UO_458 (O_458,N_9646,N_9752);
nand UO_459 (O_459,N_9341,N_9863);
nand UO_460 (O_460,N_8751,N_8142);
nand UO_461 (O_461,N_7580,N_9923);
nand UO_462 (O_462,N_9074,N_7575);
or UO_463 (O_463,N_7618,N_8137);
xor UO_464 (O_464,N_7828,N_9736);
nor UO_465 (O_465,N_9905,N_9869);
xnor UO_466 (O_466,N_8522,N_9702);
nor UO_467 (O_467,N_9803,N_8443);
nand UO_468 (O_468,N_9583,N_7577);
nor UO_469 (O_469,N_7746,N_7622);
or UO_470 (O_470,N_9680,N_8685);
or UO_471 (O_471,N_9607,N_9114);
nor UO_472 (O_472,N_9425,N_8223);
or UO_473 (O_473,N_9470,N_8084);
nand UO_474 (O_474,N_9955,N_8983);
and UO_475 (O_475,N_8461,N_9170);
or UO_476 (O_476,N_8221,N_9812);
or UO_477 (O_477,N_9662,N_8038);
or UO_478 (O_478,N_9655,N_8654);
and UO_479 (O_479,N_7533,N_8152);
or UO_480 (O_480,N_9048,N_9478);
nor UO_481 (O_481,N_9925,N_8836);
xnor UO_482 (O_482,N_8662,N_8321);
nor UO_483 (O_483,N_9167,N_7938);
nor UO_484 (O_484,N_9258,N_8124);
nor UO_485 (O_485,N_8698,N_8793);
nand UO_486 (O_486,N_8005,N_7593);
nand UO_487 (O_487,N_9221,N_9765);
nor UO_488 (O_488,N_7788,N_8410);
nand UO_489 (O_489,N_8825,N_8077);
nand UO_490 (O_490,N_9286,N_8147);
or UO_491 (O_491,N_9178,N_9052);
nand UO_492 (O_492,N_9008,N_8700);
nand UO_493 (O_493,N_7699,N_9784);
and UO_494 (O_494,N_9119,N_8318);
nand UO_495 (O_495,N_8251,N_7945);
and UO_496 (O_496,N_9290,N_9894);
xnor UO_497 (O_497,N_9233,N_8006);
and UO_498 (O_498,N_9807,N_9453);
nor UO_499 (O_499,N_9888,N_8224);
or UO_500 (O_500,N_9837,N_7839);
and UO_501 (O_501,N_7614,N_8780);
nand UO_502 (O_502,N_9964,N_7880);
nor UO_503 (O_503,N_8076,N_9935);
nor UO_504 (O_504,N_8677,N_7515);
xor UO_505 (O_505,N_9362,N_8658);
or UO_506 (O_506,N_9675,N_9676);
xnor UO_507 (O_507,N_7806,N_7579);
and UO_508 (O_508,N_9169,N_8714);
and UO_509 (O_509,N_9559,N_9144);
nand UO_510 (O_510,N_8353,N_7574);
nand UO_511 (O_511,N_9079,N_9107);
or UO_512 (O_512,N_8296,N_8930);
nand UO_513 (O_513,N_9628,N_7606);
or UO_514 (O_514,N_8795,N_8446);
and UO_515 (O_515,N_7872,N_8770);
and UO_516 (O_516,N_7560,N_7585);
and UO_517 (O_517,N_9108,N_9281);
nand UO_518 (O_518,N_9574,N_8438);
nor UO_519 (O_519,N_7654,N_9551);
or UO_520 (O_520,N_7792,N_7996);
nor UO_521 (O_521,N_9034,N_8909);
nand UO_522 (O_522,N_9620,N_7829);
nand UO_523 (O_523,N_8779,N_8539);
xor UO_524 (O_524,N_9326,N_9220);
nand UO_525 (O_525,N_8255,N_7833);
or UO_526 (O_526,N_9109,N_9117);
or UO_527 (O_527,N_8030,N_7680);
or UO_528 (O_528,N_9307,N_9084);
xnor UO_529 (O_529,N_9629,N_7609);
or UO_530 (O_530,N_9755,N_8744);
nand UO_531 (O_531,N_8450,N_9123);
or UO_532 (O_532,N_7753,N_7687);
nor UO_533 (O_533,N_8264,N_9356);
nor UO_534 (O_534,N_8235,N_7818);
or UO_535 (O_535,N_9556,N_8900);
nor UO_536 (O_536,N_9695,N_8706);
nor UO_537 (O_537,N_9754,N_8072);
or UO_538 (O_538,N_7994,N_8952);
and UO_539 (O_539,N_8367,N_8640);
or UO_540 (O_540,N_7602,N_7871);
nor UO_541 (O_541,N_9879,N_9062);
nand UO_542 (O_542,N_8933,N_8708);
nor UO_543 (O_543,N_7897,N_9495);
nand UO_544 (O_544,N_7507,N_9884);
nand UO_545 (O_545,N_9581,N_9128);
and UO_546 (O_546,N_8596,N_8068);
nand UO_547 (O_547,N_8293,N_7527);
and UO_548 (O_548,N_7917,N_9880);
xor UO_549 (O_549,N_9922,N_9591);
or UO_550 (O_550,N_7652,N_9761);
nand UO_551 (O_551,N_8792,N_9225);
nand UO_552 (O_552,N_9834,N_9508);
or UO_553 (O_553,N_9137,N_8786);
xnor UO_554 (O_554,N_8179,N_9288);
nand UO_555 (O_555,N_9430,N_8242);
nand UO_556 (O_556,N_8559,N_9135);
and UO_557 (O_557,N_7879,N_8185);
xnor UO_558 (O_558,N_9671,N_8121);
nor UO_559 (O_559,N_9124,N_8326);
nor UO_560 (O_560,N_9783,N_9567);
nand UO_561 (O_561,N_8280,N_8672);
or UO_562 (O_562,N_9522,N_9391);
and UO_563 (O_563,N_9773,N_7892);
xor UO_564 (O_564,N_9772,N_8827);
nor UO_565 (O_565,N_8449,N_9686);
or UO_566 (O_566,N_7775,N_9274);
nand UO_567 (O_567,N_8352,N_8624);
and UO_568 (O_568,N_9477,N_9697);
and UO_569 (O_569,N_7738,N_9513);
nor UO_570 (O_570,N_7830,N_9747);
nor UO_571 (O_571,N_8543,N_8716);
nor UO_572 (O_572,N_8847,N_7918);
nor UO_573 (O_573,N_8113,N_9805);
and UO_574 (O_574,N_9320,N_8620);
nand UO_575 (O_575,N_8341,N_8285);
and UO_576 (O_576,N_9031,N_9975);
and UO_577 (O_577,N_8525,N_9316);
or UO_578 (O_578,N_9976,N_9710);
xor UO_579 (O_579,N_9006,N_8609);
or UO_580 (O_580,N_9367,N_8094);
nor UO_581 (O_581,N_8213,N_8997);
nand UO_582 (O_582,N_9592,N_8034);
xor UO_583 (O_583,N_9459,N_8868);
or UO_584 (O_584,N_7657,N_8558);
or UO_585 (O_585,N_9908,N_9431);
xor UO_586 (O_586,N_7940,N_8969);
nand UO_587 (O_587,N_7793,N_8316);
or UO_588 (O_588,N_9887,N_8175);
nor UO_589 (O_589,N_8560,N_9057);
or UO_590 (O_590,N_8000,N_7965);
xor UO_591 (O_591,N_9664,N_8595);
and UO_592 (O_592,N_9061,N_8483);
or UO_593 (O_593,N_7789,N_7862);
nor UO_594 (O_594,N_8356,N_9825);
nand UO_595 (O_595,N_8403,N_9604);
or UO_596 (O_596,N_7510,N_7751);
or UO_597 (O_597,N_8819,N_8835);
nor UO_598 (O_598,N_9279,N_9674);
nand UO_599 (O_599,N_9163,N_9738);
and UO_600 (O_600,N_8366,N_8748);
or UO_601 (O_601,N_8277,N_8347);
nand UO_602 (O_602,N_8573,N_9766);
and UO_603 (O_603,N_7514,N_7903);
or UO_604 (O_604,N_9768,N_8563);
or UO_605 (O_605,N_7729,N_7500);
xnor UO_606 (O_606,N_9790,N_7672);
and UO_607 (O_607,N_7644,N_8365);
xnor UO_608 (O_608,N_7564,N_7745);
xnor UO_609 (O_609,N_8131,N_9230);
or UO_610 (O_610,N_7743,N_8872);
nor UO_611 (O_611,N_9947,N_7686);
nand UO_612 (O_612,N_9143,N_9204);
nand UO_613 (O_613,N_7534,N_8212);
nand UO_614 (O_614,N_8756,N_9650);
nand UO_615 (O_615,N_8098,N_7700);
or UO_616 (O_616,N_9205,N_7516);
nor UO_617 (O_617,N_8019,N_7613);
and UO_618 (O_618,N_9166,N_9720);
nor UO_619 (O_619,N_7824,N_7866);
nor UO_620 (O_620,N_9756,N_9451);
and UO_621 (O_621,N_9900,N_8368);
or UO_622 (O_622,N_9394,N_8138);
nor UO_623 (O_623,N_8928,N_8848);
nor UO_624 (O_624,N_9801,N_9810);
and UO_625 (O_625,N_8736,N_8957);
nand UO_626 (O_626,N_9791,N_8090);
and UO_627 (O_627,N_9898,N_9927);
nand UO_628 (O_628,N_8867,N_9558);
xnor UO_629 (O_629,N_9943,N_8267);
nand UO_630 (O_630,N_9512,N_8752);
nor UO_631 (O_631,N_7896,N_8765);
or UO_632 (O_632,N_8232,N_8987);
or UO_633 (O_633,N_8512,N_8924);
nor UO_634 (O_634,N_9939,N_9019);
nand UO_635 (O_635,N_8645,N_8510);
xnor UO_636 (O_636,N_8169,N_8625);
nand UO_637 (O_637,N_9526,N_7705);
and UO_638 (O_638,N_8947,N_8492);
xnor UO_639 (O_639,N_8572,N_9547);
nand UO_640 (O_640,N_9012,N_9465);
and UO_641 (O_641,N_8678,N_7710);
or UO_642 (O_642,N_9165,N_9302);
xnor UO_643 (O_643,N_9637,N_8263);
nand UO_644 (O_644,N_8717,N_8479);
or UO_645 (O_645,N_9413,N_9578);
nor UO_646 (O_646,N_8130,N_7999);
and UO_647 (O_647,N_9255,N_8196);
nand UO_648 (O_648,N_9201,N_8962);
nand UO_649 (O_649,N_8619,N_8259);
nand UO_650 (O_650,N_8226,N_9518);
nor UO_651 (O_651,N_7794,N_8739);
nand UO_652 (O_652,N_8101,N_9875);
nand UO_653 (O_653,N_9120,N_9989);
nor UO_654 (O_654,N_9437,N_8745);
xnor UO_655 (O_655,N_7583,N_9769);
nand UO_656 (O_656,N_9849,N_9308);
nand UO_657 (O_657,N_9717,N_9502);
or UO_658 (O_658,N_9450,N_9910);
nand UO_659 (O_659,N_7769,N_9840);
or UO_660 (O_660,N_9839,N_8891);
or UO_661 (O_661,N_7584,N_8532);
nand UO_662 (O_662,N_9284,N_7840);
or UO_663 (O_663,N_7661,N_8389);
nor UO_664 (O_664,N_9977,N_9758);
and UO_665 (O_665,N_8690,N_9086);
or UO_666 (O_666,N_7712,N_8440);
or UO_667 (O_667,N_8203,N_8120);
nand UO_668 (O_668,N_9824,N_8758);
or UO_669 (O_669,N_9737,N_7760);
nor UO_670 (O_670,N_8078,N_9222);
nand UO_671 (O_671,N_9965,N_8785);
or UO_672 (O_672,N_9815,N_8471);
or UO_673 (O_673,N_9979,N_7733);
or UO_674 (O_674,N_8191,N_7739);
nand UO_675 (O_675,N_9614,N_9523);
xnor UO_676 (O_676,N_8465,N_8802);
nand UO_677 (O_677,N_8140,N_9378);
or UO_678 (O_678,N_8245,N_9427);
and UO_679 (O_679,N_7632,N_9972);
xnor UO_680 (O_680,N_8733,N_7831);
and UO_681 (O_681,N_9197,N_8561);
xnor UO_682 (O_682,N_7732,N_8773);
or UO_683 (O_683,N_9608,N_9377);
nor UO_684 (O_684,N_8381,N_9683);
or UO_685 (O_685,N_8491,N_9035);
or UO_686 (O_686,N_8329,N_8660);
or UO_687 (O_687,N_8582,N_9468);
or UO_688 (O_688,N_9640,N_8839);
nor UO_689 (O_689,N_7962,N_8990);
xnor UO_690 (O_690,N_8383,N_9693);
nor UO_691 (O_691,N_8248,N_9027);
xor UO_692 (O_692,N_9287,N_7767);
nor UO_693 (O_693,N_8789,N_9016);
xor UO_694 (O_694,N_9854,N_9540);
or UO_695 (O_695,N_8218,N_8333);
or UO_696 (O_696,N_9723,N_9216);
nand UO_697 (O_697,N_8970,N_9434);
nand UO_698 (O_698,N_8004,N_8136);
or UO_699 (O_699,N_8555,N_7807);
or UO_700 (O_700,N_7558,N_8197);
nand UO_701 (O_701,N_9933,N_8456);
nand UO_702 (O_702,N_8991,N_7655);
nor UO_703 (O_703,N_7573,N_9698);
nor UO_704 (O_704,N_8740,N_8843);
nor UO_705 (O_705,N_9534,N_8070);
or UO_706 (O_706,N_9317,N_9991);
or UO_707 (O_707,N_9218,N_7636);
nand UO_708 (O_708,N_9426,N_9990);
nor UO_709 (O_709,N_9785,N_8357);
and UO_710 (O_710,N_9739,N_7749);
or UO_711 (O_711,N_7951,N_9096);
nor UO_712 (O_712,N_8988,N_9250);
or UO_713 (O_713,N_9641,N_7521);
nor UO_714 (O_714,N_8992,N_9657);
nand UO_715 (O_715,N_9339,N_9634);
and UO_716 (O_716,N_9340,N_9273);
and UO_717 (O_717,N_7856,N_9033);
nor UO_718 (O_718,N_9090,N_7650);
or UO_719 (O_719,N_9332,N_7736);
nor UO_720 (O_720,N_8432,N_7660);
or UO_721 (O_721,N_7604,N_7698);
or UO_722 (O_722,N_7695,N_8632);
nand UO_723 (O_723,N_8178,N_8199);
and UO_724 (O_724,N_9157,N_9003);
nor UO_725 (O_725,N_9065,N_9253);
nor UO_726 (O_726,N_8542,N_8863);
and UO_727 (O_727,N_9786,N_8846);
and UO_728 (O_728,N_9677,N_8973);
and UO_729 (O_729,N_9455,N_8330);
nand UO_730 (O_730,N_9986,N_9691);
nand UO_731 (O_731,N_8637,N_7639);
nor UO_732 (O_732,N_8100,N_9573);
nand UO_733 (O_733,N_9996,N_9206);
and UO_734 (O_734,N_7653,N_8269);
nor UO_735 (O_735,N_9156,N_8049);
nor UO_736 (O_736,N_7640,N_9310);
nand UO_737 (O_737,N_8386,N_8139);
or UO_738 (O_738,N_9814,N_8798);
nand UO_739 (O_739,N_9746,N_7973);
xor UO_740 (O_740,N_9069,N_9970);
xnor UO_741 (O_741,N_8182,N_9658);
nor UO_742 (O_742,N_9384,N_9303);
xor UO_743 (O_743,N_9223,N_7975);
nand UO_744 (O_744,N_7984,N_8036);
and UO_745 (O_745,N_9182,N_7615);
and UO_746 (O_746,N_7968,N_9902);
nor UO_747 (O_747,N_7630,N_7628);
or UO_748 (O_748,N_9381,N_8610);
and UO_749 (O_749,N_8699,N_7557);
or UO_750 (O_750,N_8260,N_9328);
nand UO_751 (O_751,N_8813,N_9678);
nand UO_752 (O_752,N_9181,N_8302);
or UO_753 (O_753,N_8091,N_9445);
and UO_754 (O_754,N_8682,N_8111);
nand UO_755 (O_755,N_8936,N_9652);
nor UO_756 (O_756,N_7837,N_7924);
nand UO_757 (O_757,N_8893,N_7519);
nand UO_758 (O_758,N_9387,N_7838);
or UO_759 (O_759,N_8495,N_9684);
nand UO_760 (O_760,N_8634,N_8822);
nand UO_761 (O_761,N_8775,N_9280);
nand UO_762 (O_762,N_9385,N_8349);
nor UO_763 (O_763,N_8033,N_9138);
nand UO_764 (O_764,N_8464,N_7718);
nor UO_765 (O_765,N_8935,N_8061);
nor UO_766 (O_766,N_9531,N_9379);
and UO_767 (O_767,N_8247,N_8614);
nor UO_768 (O_768,N_8336,N_8289);
and UO_769 (O_769,N_8679,N_7764);
nor UO_770 (O_770,N_8942,N_9023);
nor UO_771 (O_771,N_9699,N_8439);
nor UO_772 (O_772,N_8905,N_9127);
xnor UO_773 (O_773,N_8385,N_9763);
and UO_774 (O_774,N_8021,N_9112);
nand UO_775 (O_775,N_9158,N_8497);
xnor UO_776 (O_776,N_8214,N_8799);
and UO_777 (O_777,N_8731,N_9038);
nand UO_778 (O_778,N_7912,N_9870);
or UO_779 (O_779,N_9487,N_7724);
nor UO_780 (O_780,N_8470,N_8016);
nand UO_781 (O_781,N_8500,N_9238);
and UO_782 (O_782,N_8426,N_8906);
and UO_783 (O_783,N_9486,N_8626);
and UO_784 (O_784,N_8788,N_8453);
and UO_785 (O_785,N_7586,N_8160);
or UO_786 (O_786,N_7955,N_8402);
nand UO_787 (O_787,N_7617,N_7683);
nand UO_788 (O_788,N_8193,N_8411);
or UO_789 (O_789,N_7795,N_9525);
nand UO_790 (O_790,N_9346,N_9748);
or UO_791 (O_791,N_9321,N_7702);
and UO_792 (O_792,N_7923,N_7855);
nand UO_793 (O_793,N_9577,N_8974);
nor UO_794 (O_794,N_9334,N_8870);
and UO_795 (O_795,N_7671,N_9995);
and UO_796 (O_796,N_8332,N_7977);
nor UO_797 (O_797,N_9519,N_7561);
nand UO_798 (O_798,N_9713,N_9572);
or UO_799 (O_799,N_8080,N_9132);
or UO_800 (O_800,N_9876,N_9966);
or UO_801 (O_801,N_8485,N_8393);
and UO_802 (O_802,N_8243,N_9443);
and UO_803 (O_803,N_8482,N_7694);
nand UO_804 (O_804,N_7581,N_9937);
nand UO_805 (O_805,N_8760,N_8629);
nand UO_806 (O_806,N_8850,N_8669);
nand UO_807 (O_807,N_9262,N_9649);
or UO_808 (O_808,N_8631,N_9173);
and UO_809 (O_809,N_8834,N_9259);
or UO_810 (O_810,N_7674,N_8086);
and UO_811 (O_811,N_8311,N_9272);
nand UO_812 (O_812,N_7648,N_9993);
nand UO_813 (O_813,N_8511,N_8771);
xnor UO_814 (O_814,N_8444,N_9891);
or UO_815 (O_815,N_7974,N_8907);
or UO_816 (O_816,N_7805,N_7512);
nand UO_817 (O_817,N_8409,N_9802);
and UO_818 (O_818,N_8219,N_8896);
nor UO_819 (O_819,N_8173,N_8583);
nand UO_820 (O_820,N_9760,N_7980);
and UO_821 (O_821,N_9826,N_8728);
or UO_822 (O_822,N_8358,N_9672);
nor UO_823 (O_823,N_7932,N_7827);
or UO_824 (O_824,N_8871,N_7935);
and UO_825 (O_825,N_9974,N_9503);
nor UO_826 (O_826,N_7779,N_7502);
xnor UO_827 (O_827,N_9774,N_7761);
nand UO_828 (O_828,N_8715,N_7785);
nand UO_829 (O_829,N_9906,N_8954);
nand UO_830 (O_830,N_9198,N_7783);
nand UO_831 (O_831,N_9727,N_8493);
or UO_832 (O_832,N_8442,N_8273);
nor UO_833 (O_833,N_7663,N_8231);
nor UO_834 (O_834,N_8307,N_9037);
nand UO_835 (O_835,N_9406,N_9217);
nand UO_836 (O_836,N_9013,N_7920);
or UO_837 (O_837,N_8109,N_9799);
and UO_838 (O_838,N_7689,N_7525);
nand UO_839 (O_839,N_9212,N_9306);
nand UO_840 (O_840,N_9852,N_7551);
and UO_841 (O_841,N_9954,N_9463);
or UO_842 (O_842,N_8730,N_9243);
nor UO_843 (O_843,N_9557,N_8515);
or UO_844 (O_844,N_7517,N_9827);
nand UO_845 (O_845,N_9725,N_8394);
or UO_846 (O_846,N_8406,N_9440);
and UO_847 (O_847,N_7587,N_9896);
nor UO_848 (O_848,N_8053,N_7900);
and UO_849 (O_849,N_9336,N_7503);
and UO_850 (O_850,N_9432,N_9818);
or UO_851 (O_851,N_7790,N_7991);
nor UO_852 (O_852,N_8451,N_7528);
and UO_853 (O_853,N_9412,N_7643);
and UO_854 (O_854,N_9694,N_8718);
and UO_855 (O_855,N_9753,N_9049);
xor UO_856 (O_856,N_8105,N_9404);
nor UO_857 (O_857,N_8899,N_8150);
nor UO_858 (O_858,N_9589,N_8041);
or UO_859 (O_859,N_8787,N_7846);
and UO_860 (O_860,N_9762,N_9002);
nand UO_861 (O_861,N_9781,N_8749);
nor UO_862 (O_862,N_8794,N_8228);
nor UO_863 (O_863,N_8009,N_8998);
nand UO_864 (O_864,N_7967,N_9800);
nor UO_865 (O_865,N_8826,N_9368);
and UO_866 (O_866,N_7762,N_8761);
or UO_867 (O_867,N_9500,N_8919);
and UO_868 (O_868,N_8023,N_9195);
and UO_869 (O_869,N_8462,N_9248);
and UO_870 (O_870,N_7637,N_9663);
nand UO_871 (O_871,N_8107,N_7943);
nor UO_872 (O_872,N_8571,N_8709);
nor UO_873 (O_873,N_7605,N_8170);
or UO_874 (O_874,N_8122,N_9325);
or UO_875 (O_875,N_9903,N_7572);
nand UO_876 (O_876,N_9040,N_7548);
and UO_877 (O_877,N_7886,N_9569);
or UO_878 (O_878,N_8206,N_9207);
and UO_879 (O_879,N_8422,N_9174);
and UO_880 (O_880,N_9944,N_7754);
and UO_881 (O_881,N_9501,N_7777);
or UO_882 (O_882,N_8364,N_9821);
or UO_883 (O_883,N_8886,N_7504);
nand UO_884 (O_884,N_9507,N_9395);
and UO_885 (O_885,N_8676,N_8898);
and UO_886 (O_886,N_8782,N_7734);
or UO_887 (O_887,N_8929,N_9973);
nor UO_888 (O_888,N_8537,N_9429);
or UO_889 (O_889,N_8320,N_9439);
or UO_890 (O_890,N_7641,N_9645);
nand UO_891 (O_891,N_9374,N_7659);
nand UO_892 (O_892,N_9360,N_7740);
xnor UO_893 (O_893,N_8189,N_9251);
nand UO_894 (O_894,N_8433,N_8548);
nor UO_895 (O_895,N_7956,N_9232);
or UO_896 (O_896,N_8135,N_8527);
or UO_897 (O_897,N_8517,N_8784);
and UO_898 (O_898,N_9393,N_9618);
nor UO_899 (O_899,N_8803,N_8250);
nand UO_900 (O_900,N_9560,N_8565);
and UO_901 (O_901,N_8664,N_8862);
or UO_902 (O_902,N_8052,N_9300);
and UO_903 (O_903,N_7693,N_8934);
or UO_904 (O_904,N_8762,N_7835);
nor UO_905 (O_905,N_8972,N_8888);
nand UO_906 (O_906,N_9704,N_9751);
nor UO_907 (O_907,N_7925,N_7952);
xor UO_908 (O_908,N_9229,N_7913);
nand UO_909 (O_909,N_9757,N_9874);
and UO_910 (O_910,N_7645,N_9490);
nand UO_911 (O_911,N_8190,N_7713);
nor UO_912 (O_912,N_7848,N_8566);
or UO_913 (O_913,N_9605,N_8192);
nor UO_914 (O_914,N_9844,N_7861);
or UO_915 (O_915,N_8638,N_8275);
and UO_916 (O_916,N_7594,N_9260);
nand UO_917 (O_917,N_7902,N_8040);
or UO_918 (O_918,N_9467,N_8313);
or UO_919 (O_919,N_9932,N_9820);
nor UO_920 (O_920,N_9505,N_8087);
and UO_921 (O_921,N_8693,N_9330);
or UO_922 (O_922,N_8056,N_9524);
or UO_923 (O_923,N_7771,N_9883);
nand UO_924 (O_924,N_9612,N_9350);
or UO_925 (O_925,N_8892,N_7801);
or UO_926 (O_926,N_8025,N_9703);
and UO_927 (O_927,N_8816,N_9938);
and UO_928 (O_928,N_7568,N_7666);
and UO_929 (O_929,N_8395,N_8382);
xor UO_930 (O_930,N_8769,N_9497);
and UO_931 (O_931,N_8967,N_8490);
nand UO_932 (O_932,N_9041,N_9549);
or UO_933 (O_933,N_9520,N_9808);
or UO_934 (O_934,N_9029,N_9679);
and UO_935 (O_935,N_7812,N_9331);
xnor UO_936 (O_936,N_7647,N_8840);
nand UO_937 (O_937,N_9177,N_9712);
or UO_938 (O_938,N_7969,N_7543);
or UO_939 (O_939,N_8270,N_7958);
or UO_940 (O_940,N_7899,N_8796);
or UO_941 (O_941,N_8956,N_9643);
nor UO_942 (O_942,N_9113,N_7711);
nand UO_943 (O_943,N_8475,N_9602);
and UO_944 (O_944,N_7941,N_8808);
or UO_945 (O_945,N_9546,N_7719);
nand UO_946 (O_946,N_7596,N_9595);
and UO_947 (O_947,N_7508,N_8415);
nand UO_948 (O_948,N_8233,N_8976);
and UO_949 (O_949,N_7998,N_8014);
and UO_950 (O_950,N_9266,N_9514);
nand UO_951 (O_951,N_7921,N_7979);
nand UO_952 (O_952,N_9099,N_8177);
nor UO_953 (O_953,N_7865,N_9945);
nand UO_954 (O_954,N_7576,N_8766);
nor UO_955 (O_955,N_9136,N_9971);
nand UO_956 (O_956,N_8703,N_8651);
nor UO_957 (O_957,N_7616,N_8743);
and UO_958 (O_958,N_9892,N_8104);
and UO_959 (O_959,N_8155,N_7756);
and UO_960 (O_960,N_9882,N_8055);
nor UO_961 (O_961,N_8234,N_8989);
nor UO_962 (O_962,N_9071,N_9745);
nand UO_963 (O_963,N_9371,N_7876);
nor UO_964 (O_964,N_7864,N_9517);
nand UO_965 (O_965,N_7907,N_8781);
and UO_966 (O_966,N_8229,N_8528);
and UO_967 (O_967,N_9962,N_8686);
nor UO_968 (O_968,N_7815,N_9078);
nand UO_969 (O_969,N_7763,N_9245);
or UO_970 (O_970,N_8911,N_8757);
and UO_971 (O_971,N_7538,N_8458);
nand UO_972 (O_972,N_8628,N_7678);
xor UO_973 (O_973,N_9087,N_7847);
xnor UO_974 (O_974,N_9660,N_7883);
and UO_975 (O_975,N_8680,N_8681);
or UO_976 (O_976,N_8612,N_9899);
nor UO_977 (O_977,N_9200,N_7748);
and UO_978 (O_978,N_8290,N_9408);
and UO_979 (O_979,N_7546,N_7850);
or UO_980 (O_980,N_9920,N_7626);
or UO_981 (O_981,N_9571,N_8841);
nor UO_982 (O_982,N_8405,N_9460);
xor UO_983 (O_983,N_9626,N_9396);
nand UO_984 (O_984,N_8079,N_9651);
nor UO_985 (O_985,N_7550,N_9372);
nor UO_986 (O_986,N_9397,N_8806);
nand UO_987 (O_987,N_8832,N_9776);
xor UO_988 (O_988,N_8114,N_8874);
and UO_989 (O_989,N_9100,N_8473);
nor UO_990 (O_990,N_9133,N_9689);
and UO_991 (O_991,N_8633,N_9025);
nor UO_992 (O_992,N_8082,N_9794);
nand UO_993 (O_993,N_8376,N_8468);
nand UO_994 (O_994,N_9915,N_8102);
nand UO_995 (O_995,N_7766,N_7804);
and UO_996 (O_996,N_8447,N_7936);
or UO_997 (O_997,N_8216,N_9630);
nand UO_998 (O_998,N_9369,N_9740);
or UO_999 (O_999,N_9045,N_8195);
xnor UO_1000 (O_1000,N_8207,N_9337);
nand UO_1001 (O_1001,N_8869,N_8032);
nand UO_1002 (O_1002,N_9080,N_9154);
nand UO_1003 (O_1003,N_9985,N_8950);
nor UO_1004 (O_1004,N_7690,N_7914);
xor UO_1005 (O_1005,N_7723,N_7915);
or UO_1006 (O_1006,N_9862,N_8546);
or UO_1007 (O_1007,N_8047,N_8044);
nor UO_1008 (O_1008,N_9448,N_9318);
nand UO_1009 (O_1009,N_8246,N_8414);
xor UO_1010 (O_1010,N_8046,N_9382);
or UO_1011 (O_1011,N_9622,N_9289);
nand UO_1012 (O_1012,N_8067,N_8354);
and UO_1013 (O_1013,N_9189,N_8995);
nor UO_1014 (O_1014,N_8237,N_8110);
xor UO_1015 (O_1015,N_8050,N_9553);
nor UO_1016 (O_1016,N_9493,N_9366);
nor UO_1017 (O_1017,N_9462,N_8695);
and UO_1018 (O_1018,N_8691,N_8881);
nor UO_1019 (O_1019,N_7509,N_7631);
nand UO_1020 (O_1020,N_8575,N_8391);
or UO_1021 (O_1021,N_9007,N_8516);
and UO_1022 (O_1022,N_7826,N_9543);
xnor UO_1023 (O_1023,N_9484,N_9792);
nor UO_1024 (O_1024,N_7802,N_8171);
nand UO_1025 (O_1025,N_9265,N_8581);
nand UO_1026 (O_1026,N_8071,N_7797);
or UO_1027 (O_1027,N_8908,N_8222);
or UO_1028 (O_1028,N_8003,N_8355);
nand UO_1029 (O_1029,N_9636,N_8217);
and UO_1030 (O_1030,N_9536,N_9295);
and UO_1031 (O_1031,N_9670,N_7681);
or UO_1032 (O_1032,N_8938,N_9621);
nand UO_1033 (O_1033,N_9847,N_7993);
nor UO_1034 (O_1034,N_9475,N_8627);
xnor UO_1035 (O_1035,N_8670,N_7901);
nor UO_1036 (O_1036,N_8580,N_9611);
and UO_1037 (O_1037,N_9278,N_8092);
or UO_1038 (O_1038,N_9735,N_8630);
xor UO_1039 (O_1039,N_8048,N_9515);
xor UO_1040 (O_1040,N_8589,N_8551);
xnor UO_1041 (O_1041,N_9011,N_8673);
or UO_1042 (O_1042,N_8529,N_8399);
and UO_1043 (O_1043,N_8851,N_9104);
nor UO_1044 (O_1044,N_8652,N_9042);
or UO_1045 (O_1045,N_9389,N_8085);
and UO_1046 (O_1046,N_9850,N_8605);
xor UO_1047 (O_1047,N_9292,N_9779);
nand UO_1048 (O_1048,N_8279,N_8705);
and UO_1049 (O_1049,N_8272,N_9842);
or UO_1050 (O_1050,N_7620,N_9160);
nor UO_1051 (O_1051,N_9298,N_9282);
xnor UO_1052 (O_1052,N_9498,N_8817);
and UO_1053 (O_1053,N_9967,N_8861);
and UO_1054 (O_1054,N_9050,N_7673);
or UO_1055 (O_1055,N_7820,N_8755);
or UO_1056 (O_1056,N_8607,N_8735);
and UO_1057 (O_1057,N_9435,N_7963);
or UO_1058 (O_1058,N_9405,N_7853);
and UO_1059 (O_1059,N_9829,N_7946);
nor UO_1060 (O_1060,N_9456,N_9744);
and UO_1061 (O_1061,N_8923,N_7588);
nand UO_1062 (O_1062,N_8081,N_9479);
nor UO_1063 (O_1063,N_9180,N_9959);
nor UO_1064 (O_1064,N_8505,N_7735);
nor UO_1065 (O_1065,N_9032,N_8655);
nand UO_1066 (O_1066,N_8146,N_9823);
nand UO_1067 (O_1067,N_8797,N_8604);
and UO_1068 (O_1068,N_7934,N_9417);
nor UO_1069 (O_1069,N_7809,N_7744);
nor UO_1070 (O_1070,N_8258,N_8083);
nor UO_1071 (O_1071,N_7553,N_7786);
or UO_1072 (O_1072,N_7633,N_8791);
and UO_1073 (O_1073,N_9931,N_7582);
nor UO_1074 (O_1074,N_8922,N_7599);
or UO_1075 (O_1075,N_9866,N_9848);
xnor UO_1076 (O_1076,N_8943,N_8306);
and UO_1077 (O_1077,N_8978,N_9871);
and UO_1078 (O_1078,N_8554,N_7770);
nand UO_1079 (O_1079,N_9410,N_9987);
nor UO_1080 (O_1080,N_9510,N_7972);
nor UO_1081 (O_1081,N_9958,N_7544);
xnor UO_1082 (O_1082,N_8294,N_9980);
or UO_1083 (O_1083,N_8116,N_8644);
xnor UO_1084 (O_1084,N_7634,N_8045);
and UO_1085 (O_1085,N_8348,N_7928);
and UO_1086 (O_1086,N_9606,N_9952);
and UO_1087 (O_1087,N_7549,N_8568);
nor UO_1088 (O_1088,N_9376,N_9617);
nand UO_1089 (O_1089,N_9480,N_9594);
or UO_1090 (O_1090,N_8154,N_9141);
or UO_1091 (O_1091,N_9940,N_7787);
nor UO_1092 (O_1092,N_8166,N_9315);
nor UO_1093 (O_1093,N_8916,N_7664);
or UO_1094 (O_1094,N_7668,N_8194);
nand UO_1095 (O_1095,N_7851,N_8132);
or UO_1096 (O_1096,N_8011,N_7721);
nand UO_1097 (O_1097,N_9564,N_9764);
or UO_1098 (O_1098,N_8018,N_8117);
nor UO_1099 (O_1099,N_8271,N_8088);
or UO_1100 (O_1100,N_9901,N_7908);
nand UO_1101 (O_1101,N_8894,N_8577);
or UO_1102 (O_1102,N_9580,N_8913);
nand UO_1103 (O_1103,N_8315,N_9349);
nand UO_1104 (O_1104,N_8257,N_9700);
nor UO_1105 (O_1105,N_8484,N_8057);
nor UO_1106 (O_1106,N_9568,N_8984);
and UO_1107 (O_1107,N_8340,N_7677);
xor UO_1108 (O_1108,N_9997,N_7535);
xor UO_1109 (O_1109,N_9190,N_9461);
nor UO_1110 (O_1110,N_8429,N_7874);
nand UO_1111 (O_1111,N_9999,N_8926);
and UO_1112 (O_1112,N_8377,N_7953);
xor UO_1113 (O_1113,N_8617,N_8737);
or UO_1114 (O_1114,N_9830,N_8767);
nand UO_1115 (O_1115,N_9116,N_9118);
nor UO_1116 (O_1116,N_9599,N_9070);
xor UO_1117 (O_1117,N_9661,N_9819);
xor UO_1118 (O_1118,N_8412,N_9673);
and UO_1119 (O_1119,N_8252,N_7832);
or UO_1120 (O_1120,N_8594,N_8176);
nand UO_1121 (O_1121,N_7567,N_8075);
nand UO_1122 (O_1122,N_8759,N_9668);
nand UO_1123 (O_1123,N_9140,N_9859);
nand UO_1124 (O_1124,N_8337,N_8901);
nor UO_1125 (O_1125,N_9383,N_7589);
or UO_1126 (O_1126,N_9446,N_8261);
and UO_1127 (O_1127,N_8300,N_9555);
or UO_1128 (O_1128,N_9653,N_8346);
or UO_1129 (O_1129,N_9610,N_9897);
and UO_1130 (O_1130,N_9105,N_8521);
or UO_1131 (O_1131,N_9319,N_9208);
nor UO_1132 (O_1132,N_9726,N_8999);
or UO_1133 (O_1133,N_9639,N_8106);
and UO_1134 (O_1134,N_7976,N_9984);
and UO_1135 (O_1135,N_9911,N_9234);
and UO_1136 (O_1136,N_8398,N_9293);
xor UO_1137 (O_1137,N_9953,N_8028);
xnor UO_1138 (O_1138,N_8301,N_9047);
or UO_1139 (O_1139,N_9010,N_8535);
or UO_1140 (O_1140,N_9516,N_9682);
and UO_1141 (O_1141,N_7985,N_9375);
nor UO_1142 (O_1142,N_8283,N_9202);
nor UO_1143 (O_1143,N_9481,N_7772);
nor UO_1144 (O_1144,N_7737,N_8809);
and UO_1145 (O_1145,N_9219,N_9449);
nor UO_1146 (O_1146,N_9402,N_8474);
or UO_1147 (O_1147,N_9775,N_8520);
and UO_1148 (O_1148,N_8024,N_8392);
or UO_1149 (O_1149,N_7887,N_9101);
and UO_1150 (O_1150,N_9227,N_8380);
and UO_1151 (O_1151,N_7905,N_8188);
nor UO_1152 (O_1152,N_9304,N_8322);
nor UO_1153 (O_1153,N_8295,N_9722);
nor UO_1154 (O_1154,N_8608,N_9833);
nor UO_1155 (O_1155,N_7909,N_9082);
nand UO_1156 (O_1156,N_9877,N_9390);
xnor UO_1157 (O_1157,N_9609,N_9588);
nor UO_1158 (O_1158,N_9083,N_9960);
and UO_1159 (O_1159,N_9930,N_9615);
nand UO_1160 (O_1160,N_8776,N_8126);
and UO_1161 (O_1161,N_8830,N_8238);
and UO_1162 (O_1162,N_8917,N_9309);
nand UO_1163 (O_1163,N_9054,N_7959);
and UO_1164 (O_1164,N_8361,N_8478);
nor UO_1165 (O_1165,N_8569,N_9770);
nor UO_1166 (O_1166,N_8174,N_9690);
nand UO_1167 (O_1167,N_9509,N_7817);
nor UO_1168 (O_1168,N_9782,N_8961);
or UO_1169 (O_1169,N_9734,N_7552);
nand UO_1170 (O_1170,N_8959,N_8878);
nand UO_1171 (O_1171,N_9860,N_7518);
nor UO_1172 (O_1172,N_9139,N_9701);
nand UO_1173 (O_1173,N_7720,N_7715);
or UO_1174 (O_1174,N_8335,N_8732);
nor UO_1175 (O_1175,N_8591,N_7776);
and UO_1176 (O_1176,N_7834,N_8509);
or UO_1177 (O_1177,N_8421,N_8419);
and UO_1178 (O_1178,N_8118,N_7601);
or UO_1179 (O_1179,N_8887,N_9464);
xnor UO_1180 (O_1180,N_9631,N_8157);
nor UO_1181 (O_1181,N_9845,N_9028);
and UO_1182 (O_1182,N_9073,N_9994);
nor UO_1183 (O_1183,N_9401,N_8643);
or UO_1184 (O_1184,N_9075,N_8211);
and UO_1185 (O_1185,N_9089,N_9240);
or UO_1186 (O_1186,N_8428,N_8702);
nor UO_1187 (O_1187,N_7730,N_9711);
or UO_1188 (O_1188,N_7714,N_8902);
or UO_1189 (O_1189,N_7800,N_7863);
nand UO_1190 (O_1190,N_9858,N_9301);
xnor UO_1191 (O_1191,N_9322,N_9983);
nand UO_1192 (O_1192,N_7742,N_7814);
xor UO_1193 (O_1193,N_9796,N_9798);
nand UO_1194 (O_1194,N_8865,N_8530);
nand UO_1195 (O_1195,N_7898,N_7843);
or UO_1196 (O_1196,N_9203,N_9020);
xor UO_1197 (O_1197,N_9399,N_9832);
nand UO_1198 (O_1198,N_8550,N_7597);
nor UO_1199 (O_1199,N_7944,N_9719);
or UO_1200 (O_1200,N_9616,N_8649);
and UO_1201 (O_1201,N_9063,N_8828);
or UO_1202 (O_1202,N_8039,N_7859);
nor UO_1203 (O_1203,N_9851,N_8931);
and UO_1204 (O_1204,N_8249,N_8007);
nand UO_1205 (O_1205,N_9150,N_7701);
nor UO_1206 (O_1206,N_9619,N_8457);
or UO_1207 (O_1207,N_8979,N_8134);
or UO_1208 (O_1208,N_8953,N_7569);
nor UO_1209 (O_1209,N_8855,N_8852);
or UO_1210 (O_1210,N_8856,N_7842);
nand UO_1211 (O_1211,N_7511,N_8434);
xnor UO_1212 (O_1212,N_9196,N_8857);
nor UO_1213 (O_1213,N_7731,N_8985);
and UO_1214 (O_1214,N_7791,N_9392);
or UO_1215 (O_1215,N_8013,N_9436);
or UO_1216 (O_1216,N_8636,N_9817);
xor UO_1217 (O_1217,N_9928,N_8711);
xnor UO_1218 (O_1218,N_8918,N_7603);
and UO_1219 (O_1219,N_8659,N_8304);
or UO_1220 (O_1220,N_9422,N_8288);
and UO_1221 (O_1221,N_9864,N_8362);
or UO_1222 (O_1222,N_8292,N_9961);
and UO_1223 (O_1223,N_7619,N_9247);
nor UO_1224 (O_1224,N_8158,N_8820);
nand UO_1225 (O_1225,N_8635,N_9597);
or UO_1226 (O_1226,N_9209,N_8093);
xor UO_1227 (O_1227,N_9709,N_8587);
xnor UO_1228 (O_1228,N_9733,N_9853);
nor UO_1229 (O_1229,N_9275,N_8955);
nand UO_1230 (O_1230,N_7893,N_9060);
or UO_1231 (O_1231,N_7530,N_7755);
and UO_1232 (O_1232,N_7717,N_9806);
nand UO_1233 (O_1233,N_7911,N_9416);
xor UO_1234 (O_1234,N_8459,N_8729);
and UO_1235 (O_1235,N_8035,N_8585);
nor UO_1236 (O_1236,N_8963,N_9252);
nand UO_1237 (O_1237,N_9529,N_8455);
nor UO_1238 (O_1238,N_7532,N_8022);
nor UO_1239 (O_1239,N_9946,N_9335);
or UO_1240 (O_1240,N_9268,N_7986);
nand UO_1241 (O_1241,N_7845,N_9373);
and UO_1242 (O_1242,N_8823,N_8133);
xnor UO_1243 (O_1243,N_7819,N_8001);
nor UO_1244 (O_1244,N_8829,N_7803);
and UO_1245 (O_1245,N_8696,N_7919);
and UO_1246 (O_1246,N_9861,N_7542);
xnor UO_1247 (O_1247,N_9361,N_8487);
nand UO_1248 (O_1248,N_9039,N_9904);
xnor UO_1249 (O_1249,N_8912,N_9471);
nor UO_1250 (O_1250,N_9134,N_9680);
nand UO_1251 (O_1251,N_7929,N_8233);
nor UO_1252 (O_1252,N_8149,N_8082);
and UO_1253 (O_1253,N_9537,N_8320);
and UO_1254 (O_1254,N_8585,N_8840);
and UO_1255 (O_1255,N_8833,N_9808);
nand UO_1256 (O_1256,N_7596,N_9034);
and UO_1257 (O_1257,N_8505,N_8856);
or UO_1258 (O_1258,N_9904,N_9701);
xor UO_1259 (O_1259,N_9196,N_8563);
xnor UO_1260 (O_1260,N_9963,N_8337);
and UO_1261 (O_1261,N_9406,N_8628);
nor UO_1262 (O_1262,N_9797,N_7631);
nand UO_1263 (O_1263,N_7843,N_9297);
xor UO_1264 (O_1264,N_8226,N_9415);
or UO_1265 (O_1265,N_7624,N_9614);
and UO_1266 (O_1266,N_8634,N_7862);
nand UO_1267 (O_1267,N_7594,N_9262);
xnor UO_1268 (O_1268,N_8672,N_9442);
and UO_1269 (O_1269,N_8367,N_9153);
nand UO_1270 (O_1270,N_9602,N_8700);
nor UO_1271 (O_1271,N_8511,N_8783);
and UO_1272 (O_1272,N_8627,N_9351);
or UO_1273 (O_1273,N_9034,N_8908);
nand UO_1274 (O_1274,N_7965,N_8141);
nor UO_1275 (O_1275,N_8232,N_8989);
or UO_1276 (O_1276,N_8131,N_9220);
and UO_1277 (O_1277,N_8702,N_9700);
nand UO_1278 (O_1278,N_8229,N_9939);
xnor UO_1279 (O_1279,N_8077,N_9575);
nor UO_1280 (O_1280,N_9758,N_9675);
nand UO_1281 (O_1281,N_8193,N_8364);
nand UO_1282 (O_1282,N_7846,N_8492);
nand UO_1283 (O_1283,N_8189,N_9808);
or UO_1284 (O_1284,N_9196,N_9994);
nor UO_1285 (O_1285,N_9243,N_8410);
and UO_1286 (O_1286,N_7678,N_9624);
xnor UO_1287 (O_1287,N_8512,N_8279);
or UO_1288 (O_1288,N_7721,N_7800);
nor UO_1289 (O_1289,N_8501,N_8820);
and UO_1290 (O_1290,N_8589,N_8494);
nand UO_1291 (O_1291,N_9555,N_7736);
nor UO_1292 (O_1292,N_7552,N_8676);
nand UO_1293 (O_1293,N_7968,N_9233);
xnor UO_1294 (O_1294,N_9203,N_9028);
or UO_1295 (O_1295,N_8196,N_7730);
nand UO_1296 (O_1296,N_9461,N_9812);
nor UO_1297 (O_1297,N_7731,N_8007);
nand UO_1298 (O_1298,N_9108,N_9546);
and UO_1299 (O_1299,N_9013,N_9329);
nor UO_1300 (O_1300,N_8309,N_7749);
nand UO_1301 (O_1301,N_9101,N_9039);
xor UO_1302 (O_1302,N_8904,N_9239);
nor UO_1303 (O_1303,N_7774,N_8567);
or UO_1304 (O_1304,N_8529,N_9668);
or UO_1305 (O_1305,N_8762,N_7731);
nand UO_1306 (O_1306,N_8058,N_7691);
and UO_1307 (O_1307,N_9576,N_7910);
nand UO_1308 (O_1308,N_9113,N_7863);
or UO_1309 (O_1309,N_7817,N_8506);
or UO_1310 (O_1310,N_9358,N_9228);
nand UO_1311 (O_1311,N_8095,N_9848);
or UO_1312 (O_1312,N_7744,N_8634);
nor UO_1313 (O_1313,N_9584,N_9332);
nor UO_1314 (O_1314,N_9482,N_8004);
nor UO_1315 (O_1315,N_8337,N_8659);
or UO_1316 (O_1316,N_8280,N_8681);
nand UO_1317 (O_1317,N_9736,N_8952);
xor UO_1318 (O_1318,N_9115,N_7625);
nand UO_1319 (O_1319,N_9080,N_8558);
or UO_1320 (O_1320,N_8952,N_7914);
xor UO_1321 (O_1321,N_7746,N_7541);
nand UO_1322 (O_1322,N_8358,N_9828);
and UO_1323 (O_1323,N_7991,N_8457);
nor UO_1324 (O_1324,N_7557,N_7579);
nand UO_1325 (O_1325,N_7510,N_8633);
nand UO_1326 (O_1326,N_7892,N_8603);
nor UO_1327 (O_1327,N_7747,N_9723);
nor UO_1328 (O_1328,N_8240,N_8476);
nand UO_1329 (O_1329,N_9574,N_7800);
or UO_1330 (O_1330,N_8932,N_8570);
xor UO_1331 (O_1331,N_9326,N_9068);
or UO_1332 (O_1332,N_7966,N_9956);
nand UO_1333 (O_1333,N_9606,N_8528);
nor UO_1334 (O_1334,N_7712,N_9714);
xnor UO_1335 (O_1335,N_8696,N_7521);
or UO_1336 (O_1336,N_8913,N_7715);
or UO_1337 (O_1337,N_8680,N_8353);
or UO_1338 (O_1338,N_8951,N_8346);
nand UO_1339 (O_1339,N_9747,N_8354);
and UO_1340 (O_1340,N_9653,N_8282);
nand UO_1341 (O_1341,N_8695,N_7999);
nor UO_1342 (O_1342,N_7782,N_9595);
and UO_1343 (O_1343,N_9539,N_9622);
nand UO_1344 (O_1344,N_9668,N_8522);
and UO_1345 (O_1345,N_8208,N_7728);
or UO_1346 (O_1346,N_8538,N_8755);
or UO_1347 (O_1347,N_9563,N_8808);
and UO_1348 (O_1348,N_9735,N_9451);
or UO_1349 (O_1349,N_8325,N_9930);
and UO_1350 (O_1350,N_8452,N_7826);
and UO_1351 (O_1351,N_7517,N_8309);
nor UO_1352 (O_1352,N_9116,N_9526);
nor UO_1353 (O_1353,N_7564,N_8348);
nor UO_1354 (O_1354,N_8398,N_8970);
and UO_1355 (O_1355,N_7742,N_9439);
xnor UO_1356 (O_1356,N_8698,N_9644);
and UO_1357 (O_1357,N_8961,N_9711);
or UO_1358 (O_1358,N_8827,N_7819);
nand UO_1359 (O_1359,N_8506,N_9547);
nor UO_1360 (O_1360,N_9201,N_7662);
or UO_1361 (O_1361,N_9730,N_7964);
or UO_1362 (O_1362,N_8914,N_8650);
nand UO_1363 (O_1363,N_8914,N_7707);
or UO_1364 (O_1364,N_8961,N_7706);
nand UO_1365 (O_1365,N_7506,N_8308);
and UO_1366 (O_1366,N_9613,N_8032);
and UO_1367 (O_1367,N_7740,N_9947);
or UO_1368 (O_1368,N_9963,N_8140);
nor UO_1369 (O_1369,N_8957,N_9148);
or UO_1370 (O_1370,N_9341,N_8103);
or UO_1371 (O_1371,N_8476,N_9327);
nor UO_1372 (O_1372,N_9529,N_8257);
and UO_1373 (O_1373,N_9026,N_8092);
nor UO_1374 (O_1374,N_7617,N_8615);
nor UO_1375 (O_1375,N_7727,N_8975);
nor UO_1376 (O_1376,N_9975,N_7583);
nor UO_1377 (O_1377,N_8342,N_8992);
xor UO_1378 (O_1378,N_8066,N_9323);
or UO_1379 (O_1379,N_8300,N_8200);
or UO_1380 (O_1380,N_7809,N_9362);
xnor UO_1381 (O_1381,N_7680,N_7809);
nand UO_1382 (O_1382,N_7756,N_7511);
nor UO_1383 (O_1383,N_9500,N_8055);
or UO_1384 (O_1384,N_9571,N_7880);
nand UO_1385 (O_1385,N_9343,N_8049);
or UO_1386 (O_1386,N_9095,N_8183);
or UO_1387 (O_1387,N_7841,N_9376);
nor UO_1388 (O_1388,N_7797,N_9822);
nor UO_1389 (O_1389,N_8229,N_9007);
nor UO_1390 (O_1390,N_9021,N_9182);
xor UO_1391 (O_1391,N_9743,N_9355);
and UO_1392 (O_1392,N_8768,N_8658);
and UO_1393 (O_1393,N_8155,N_8829);
nor UO_1394 (O_1394,N_8086,N_8696);
nor UO_1395 (O_1395,N_8230,N_8508);
or UO_1396 (O_1396,N_8297,N_9907);
and UO_1397 (O_1397,N_8105,N_8869);
or UO_1398 (O_1398,N_9735,N_9120);
or UO_1399 (O_1399,N_8154,N_9135);
nor UO_1400 (O_1400,N_7742,N_8037);
nor UO_1401 (O_1401,N_9353,N_9399);
nor UO_1402 (O_1402,N_7702,N_9971);
and UO_1403 (O_1403,N_8704,N_7672);
and UO_1404 (O_1404,N_8596,N_8696);
and UO_1405 (O_1405,N_9083,N_8938);
nor UO_1406 (O_1406,N_7595,N_7536);
or UO_1407 (O_1407,N_8198,N_7960);
and UO_1408 (O_1408,N_9083,N_7689);
nand UO_1409 (O_1409,N_8357,N_9728);
or UO_1410 (O_1410,N_7828,N_9711);
nor UO_1411 (O_1411,N_7954,N_8188);
or UO_1412 (O_1412,N_8253,N_8016);
and UO_1413 (O_1413,N_8028,N_8588);
nand UO_1414 (O_1414,N_7635,N_9561);
nor UO_1415 (O_1415,N_9713,N_8508);
xor UO_1416 (O_1416,N_7634,N_7617);
nand UO_1417 (O_1417,N_9796,N_8956);
nor UO_1418 (O_1418,N_8774,N_8786);
or UO_1419 (O_1419,N_9852,N_8900);
or UO_1420 (O_1420,N_8439,N_9714);
xnor UO_1421 (O_1421,N_8273,N_8551);
and UO_1422 (O_1422,N_8838,N_8532);
nor UO_1423 (O_1423,N_8761,N_9423);
nand UO_1424 (O_1424,N_7979,N_9625);
or UO_1425 (O_1425,N_9331,N_9603);
nor UO_1426 (O_1426,N_8890,N_8006);
and UO_1427 (O_1427,N_9635,N_8863);
xor UO_1428 (O_1428,N_7538,N_7747);
nand UO_1429 (O_1429,N_8209,N_9069);
nor UO_1430 (O_1430,N_7905,N_7717);
or UO_1431 (O_1431,N_7867,N_9555);
nand UO_1432 (O_1432,N_8534,N_8168);
nand UO_1433 (O_1433,N_8116,N_8513);
nand UO_1434 (O_1434,N_9338,N_7707);
nand UO_1435 (O_1435,N_8638,N_9623);
nand UO_1436 (O_1436,N_9943,N_9922);
and UO_1437 (O_1437,N_9930,N_8919);
xnor UO_1438 (O_1438,N_9682,N_7904);
nor UO_1439 (O_1439,N_7535,N_7978);
and UO_1440 (O_1440,N_8660,N_7792);
or UO_1441 (O_1441,N_8686,N_9014);
or UO_1442 (O_1442,N_7900,N_7958);
or UO_1443 (O_1443,N_7663,N_8715);
nand UO_1444 (O_1444,N_7878,N_9619);
xnor UO_1445 (O_1445,N_8237,N_9034);
or UO_1446 (O_1446,N_9475,N_9646);
xnor UO_1447 (O_1447,N_7844,N_8535);
nor UO_1448 (O_1448,N_9192,N_8588);
or UO_1449 (O_1449,N_8131,N_9408);
and UO_1450 (O_1450,N_7830,N_9612);
nand UO_1451 (O_1451,N_8906,N_8265);
or UO_1452 (O_1452,N_9560,N_7552);
or UO_1453 (O_1453,N_9571,N_8778);
or UO_1454 (O_1454,N_9815,N_8699);
and UO_1455 (O_1455,N_8307,N_8315);
xnor UO_1456 (O_1456,N_7897,N_7864);
and UO_1457 (O_1457,N_8377,N_7940);
and UO_1458 (O_1458,N_9484,N_8314);
and UO_1459 (O_1459,N_9519,N_9591);
or UO_1460 (O_1460,N_7600,N_8685);
and UO_1461 (O_1461,N_7999,N_9477);
or UO_1462 (O_1462,N_9743,N_7556);
nor UO_1463 (O_1463,N_8845,N_9134);
nand UO_1464 (O_1464,N_8044,N_8568);
nor UO_1465 (O_1465,N_8794,N_8710);
nand UO_1466 (O_1466,N_8611,N_7626);
xnor UO_1467 (O_1467,N_9736,N_9168);
nand UO_1468 (O_1468,N_7654,N_9498);
or UO_1469 (O_1469,N_8682,N_9050);
nand UO_1470 (O_1470,N_8312,N_8617);
xnor UO_1471 (O_1471,N_7879,N_8517);
nand UO_1472 (O_1472,N_7888,N_8275);
and UO_1473 (O_1473,N_9177,N_9192);
nor UO_1474 (O_1474,N_9530,N_8324);
or UO_1475 (O_1475,N_8550,N_8900);
or UO_1476 (O_1476,N_8641,N_8854);
and UO_1477 (O_1477,N_9646,N_8842);
nand UO_1478 (O_1478,N_8411,N_9620);
or UO_1479 (O_1479,N_9390,N_8049);
nor UO_1480 (O_1480,N_9304,N_9908);
nor UO_1481 (O_1481,N_9998,N_9915);
and UO_1482 (O_1482,N_9641,N_9589);
and UO_1483 (O_1483,N_8405,N_8600);
or UO_1484 (O_1484,N_9922,N_9800);
nand UO_1485 (O_1485,N_8156,N_8358);
or UO_1486 (O_1486,N_8319,N_9759);
and UO_1487 (O_1487,N_9247,N_7922);
and UO_1488 (O_1488,N_9420,N_7606);
xnor UO_1489 (O_1489,N_9853,N_9277);
nand UO_1490 (O_1490,N_9409,N_7500);
or UO_1491 (O_1491,N_9157,N_9487);
nor UO_1492 (O_1492,N_9432,N_9005);
nor UO_1493 (O_1493,N_9416,N_9381);
nand UO_1494 (O_1494,N_9122,N_9862);
nor UO_1495 (O_1495,N_8948,N_8501);
xnor UO_1496 (O_1496,N_8169,N_9599);
and UO_1497 (O_1497,N_8326,N_9244);
nor UO_1498 (O_1498,N_9909,N_9776);
or UO_1499 (O_1499,N_9258,N_7761);
endmodule