module basic_3000_30000_3500_30_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2289,In_490);
nand U1 (N_1,In_2024,In_2507);
or U2 (N_2,In_2245,In_2145);
xnor U3 (N_3,In_2862,In_1118);
or U4 (N_4,In_1885,In_204);
nor U5 (N_5,In_2674,In_1276);
nor U6 (N_6,In_179,In_2470);
or U7 (N_7,In_2391,In_2200);
xnor U8 (N_8,In_1107,In_938);
xnor U9 (N_9,In_928,In_1673);
or U10 (N_10,In_1985,In_361);
xor U11 (N_11,In_2805,In_797);
xnor U12 (N_12,In_2929,In_321);
nand U13 (N_13,In_811,In_651);
nand U14 (N_14,In_2705,In_1551);
or U15 (N_15,In_2201,In_1873);
xor U16 (N_16,In_2804,In_1761);
or U17 (N_17,In_160,In_1709);
and U18 (N_18,In_2396,In_1462);
and U19 (N_19,In_1793,In_488);
and U20 (N_20,In_1725,In_727);
or U21 (N_21,In_925,In_301);
xnor U22 (N_22,In_427,In_932);
nand U23 (N_23,In_2652,In_2189);
nor U24 (N_24,In_763,In_1598);
and U25 (N_25,In_2136,In_1362);
or U26 (N_26,In_1190,In_871);
and U27 (N_27,In_470,In_2659);
xor U28 (N_28,In_1596,In_2184);
xnor U29 (N_29,In_323,In_237);
xnor U30 (N_30,In_971,In_1760);
and U31 (N_31,In_662,In_135);
and U32 (N_32,In_1788,In_1677);
and U33 (N_33,In_2643,In_2056);
nand U34 (N_34,In_1218,In_977);
xnor U35 (N_35,In_2259,In_789);
nor U36 (N_36,In_2103,In_182);
or U37 (N_37,In_650,In_1973);
and U38 (N_38,In_1925,In_497);
and U39 (N_39,In_1879,In_2119);
or U40 (N_40,In_2653,In_436);
nor U41 (N_41,In_2198,In_2355);
nor U42 (N_42,In_259,In_67);
nand U43 (N_43,In_2222,In_1783);
and U44 (N_44,In_1251,In_2413);
or U45 (N_45,In_2008,In_1972);
and U46 (N_46,In_1641,In_2320);
or U47 (N_47,In_2953,In_1238);
nor U48 (N_48,In_1071,In_1003);
or U49 (N_49,In_996,In_2793);
or U50 (N_50,In_1244,In_760);
nor U51 (N_51,In_743,In_2131);
xnor U52 (N_52,In_1241,In_424);
nand U53 (N_53,In_1356,In_2279);
xor U54 (N_54,In_2416,In_2577);
or U55 (N_55,In_523,In_1085);
or U56 (N_56,In_737,In_2051);
xnor U57 (N_57,In_2149,In_799);
and U58 (N_58,In_2133,In_107);
and U59 (N_59,In_324,In_1390);
xnor U60 (N_60,In_2752,In_2387);
or U61 (N_61,In_1737,In_954);
nor U62 (N_62,In_1047,In_715);
xnor U63 (N_63,In_2760,In_2171);
and U64 (N_64,In_2802,In_61);
and U65 (N_65,In_350,In_1888);
nor U66 (N_66,In_1833,In_1215);
xnor U67 (N_67,In_1548,In_446);
and U68 (N_68,In_1515,In_2064);
and U69 (N_69,In_585,In_1541);
xnor U70 (N_70,In_998,In_2376);
or U71 (N_71,In_1736,In_1120);
and U72 (N_72,In_1379,In_2300);
or U73 (N_73,In_1899,In_58);
xnor U74 (N_74,In_381,In_1773);
and U75 (N_75,In_352,In_2233);
nand U76 (N_76,In_1337,In_2878);
and U77 (N_77,In_1167,In_2780);
nand U78 (N_78,In_1662,In_586);
nor U79 (N_79,In_487,In_567);
and U80 (N_80,In_2987,In_1850);
and U81 (N_81,In_1139,In_731);
or U82 (N_82,In_607,In_1346);
nor U83 (N_83,In_1625,In_2126);
or U84 (N_84,In_2580,In_2276);
or U85 (N_85,In_2829,In_876);
nand U86 (N_86,In_1691,In_2003);
and U87 (N_87,In_1511,In_2697);
xor U88 (N_88,In_1978,In_1381);
nor U89 (N_89,In_686,In_1028);
and U90 (N_90,In_706,In_1470);
or U91 (N_91,In_1395,In_883);
nor U92 (N_92,In_2498,In_2431);
nor U93 (N_93,In_874,In_262);
xnor U94 (N_94,In_1839,In_1552);
and U95 (N_95,In_2016,In_1780);
and U96 (N_96,In_1956,In_1112);
and U97 (N_97,In_441,In_1207);
or U98 (N_98,In_113,In_120);
or U99 (N_99,In_2671,In_1684);
nand U100 (N_100,In_1225,In_2027);
xnor U101 (N_101,In_2499,In_27);
nand U102 (N_102,In_1353,In_1295);
and U103 (N_103,In_2723,In_209);
or U104 (N_104,In_20,In_2563);
and U105 (N_105,In_543,In_440);
or U106 (N_106,In_1815,In_2465);
and U107 (N_107,In_1794,In_1382);
and U108 (N_108,In_222,In_455);
nand U109 (N_109,In_1606,In_765);
nand U110 (N_110,In_2576,In_2587);
or U111 (N_111,In_2812,In_2273);
and U112 (N_112,In_2540,In_1611);
or U113 (N_113,In_2579,In_792);
or U114 (N_114,In_943,In_249);
or U115 (N_115,In_2806,In_322);
or U116 (N_116,In_518,In_2374);
or U117 (N_117,In_1876,In_754);
nor U118 (N_118,In_1664,In_126);
nand U119 (N_119,In_2473,In_1796);
xor U120 (N_120,In_2515,In_357);
nand U121 (N_121,In_1584,In_1954);
and U122 (N_122,In_2477,In_1465);
or U123 (N_123,In_1124,In_41);
and U124 (N_124,In_1443,In_1667);
xnor U125 (N_125,In_1425,In_2039);
and U126 (N_126,In_1051,In_2196);
xnor U127 (N_127,In_2637,In_2090);
and U128 (N_128,In_38,In_377);
or U129 (N_129,In_1307,In_302);
or U130 (N_130,In_327,In_1571);
or U131 (N_131,In_389,In_1715);
or U132 (N_132,In_2322,In_87);
nand U133 (N_133,In_1593,In_1367);
and U134 (N_134,In_2859,In_335);
nor U135 (N_135,In_1083,In_1280);
and U136 (N_136,In_1575,In_1073);
and U137 (N_137,In_830,In_1233);
and U138 (N_138,In_690,In_1319);
xnor U139 (N_139,In_341,In_1690);
or U140 (N_140,In_1679,In_2831);
xor U141 (N_141,In_1312,In_2611);
nor U142 (N_142,In_458,In_2510);
or U143 (N_143,In_1623,In_356);
xor U144 (N_144,In_177,In_1519);
or U145 (N_145,In_2927,In_2231);
and U146 (N_146,In_1363,In_1048);
or U147 (N_147,In_2796,In_495);
nor U148 (N_148,In_2010,In_1479);
or U149 (N_149,In_100,In_1779);
xnor U150 (N_150,In_850,In_620);
nand U151 (N_151,In_2963,In_1430);
nand U152 (N_152,In_911,In_700);
nor U153 (N_153,In_2025,In_157);
xnor U154 (N_154,In_2779,In_2028);
and U155 (N_155,In_1079,In_906);
nor U156 (N_156,In_1705,In_2047);
nor U157 (N_157,In_527,In_2932);
xor U158 (N_158,In_2712,In_935);
xnor U159 (N_159,In_1916,In_2714);
nand U160 (N_160,In_206,In_2380);
nor U161 (N_161,In_344,In_499);
nand U162 (N_162,In_288,In_2216);
nor U163 (N_163,In_376,In_1461);
nand U164 (N_164,In_997,In_717);
nand U165 (N_165,In_1608,In_2741);
nand U166 (N_166,In_1277,In_2573);
or U167 (N_167,In_1650,In_2106);
or U168 (N_168,In_2340,In_2140);
and U169 (N_169,In_858,In_2241);
nand U170 (N_170,In_2899,In_143);
or U171 (N_171,In_273,In_86);
nor U172 (N_172,In_309,In_1924);
xor U173 (N_173,In_1492,In_299);
nand U174 (N_174,In_2651,In_2130);
xnor U175 (N_175,In_168,In_2698);
or U176 (N_176,In_2182,In_286);
or U177 (N_177,In_1640,In_1365);
nand U178 (N_178,In_116,In_1132);
xnor U179 (N_179,In_2942,In_910);
and U180 (N_180,In_2732,In_485);
nor U181 (N_181,In_2619,In_2132);
and U182 (N_182,In_2301,In_2173);
or U183 (N_183,In_2744,In_439);
nand U184 (N_184,In_852,In_1106);
nor U185 (N_185,In_203,In_1377);
nand U186 (N_186,In_1039,In_2811);
and U187 (N_187,In_0,In_656);
xor U188 (N_188,In_132,In_807);
or U189 (N_189,In_189,In_820);
nor U190 (N_190,In_1834,In_1142);
nand U191 (N_191,In_106,In_2377);
nor U192 (N_192,In_1370,In_1439);
and U193 (N_193,In_474,In_90);
or U194 (N_194,In_919,In_857);
nor U195 (N_195,In_263,In_46);
xor U196 (N_196,In_1901,In_550);
nand U197 (N_197,In_2020,In_1865);
xnor U198 (N_198,In_88,In_1351);
nor U199 (N_199,In_1302,In_278);
or U200 (N_200,In_2801,In_1749);
xnor U201 (N_201,In_677,In_2411);
nand U202 (N_202,In_18,In_1521);
nor U203 (N_203,In_2737,In_1448);
and U204 (N_204,In_172,In_2917);
nand U205 (N_205,In_1620,In_1836);
nor U206 (N_206,In_2467,In_2740);
and U207 (N_207,In_465,In_1052);
or U208 (N_208,In_962,In_959);
xnor U209 (N_209,In_2581,In_877);
nand U210 (N_210,In_1605,In_1510);
or U211 (N_211,In_1756,In_1245);
nand U212 (N_212,In_1560,In_145);
xor U213 (N_213,In_663,In_313);
xor U214 (N_214,In_42,In_564);
and U215 (N_215,In_1955,In_2695);
and U216 (N_216,In_853,In_2738);
nand U217 (N_217,In_2041,In_755);
nor U218 (N_218,In_2819,In_461);
and U219 (N_219,In_1971,In_1153);
and U220 (N_220,In_1660,In_636);
nand U221 (N_221,In_1629,In_2493);
xor U222 (N_222,In_2835,In_886);
nor U223 (N_223,In_450,In_2965);
xor U224 (N_224,In_2000,In_2975);
nand U225 (N_225,In_1601,In_942);
nand U226 (N_226,In_60,In_2494);
nand U227 (N_227,In_1556,In_473);
or U228 (N_228,In_824,In_1713);
xnor U229 (N_229,In_2441,In_534);
or U230 (N_230,In_2366,In_510);
and U231 (N_231,In_2154,In_171);
or U232 (N_232,In_1587,In_1219);
nor U233 (N_233,In_909,In_1402);
or U234 (N_234,In_1919,In_1930);
nand U235 (N_235,In_334,In_720);
and U236 (N_236,In_29,In_821);
nand U237 (N_237,In_1842,In_1098);
or U238 (N_238,In_1852,In_788);
xor U239 (N_239,In_2326,In_808);
and U240 (N_240,In_2995,In_2262);
xnor U241 (N_241,In_1292,In_1333);
nand U242 (N_242,In_1758,In_2203);
or U243 (N_243,In_2762,In_268);
nand U244 (N_244,In_1661,In_21);
xor U245 (N_245,In_1375,In_383);
xor U246 (N_246,In_2770,In_2209);
nand U247 (N_247,In_804,In_181);
or U248 (N_248,In_2933,In_2827);
or U249 (N_249,In_1845,In_867);
xnor U250 (N_250,In_2316,In_664);
nand U251 (N_251,In_1180,In_669);
nor U252 (N_252,In_1838,In_1922);
xor U253 (N_253,In_380,In_2795);
or U254 (N_254,In_317,In_544);
or U255 (N_255,In_672,In_2797);
or U256 (N_256,In_868,In_1844);
nand U257 (N_257,In_696,In_2688);
nor U258 (N_258,In_1745,In_463);
and U259 (N_259,In_657,In_2113);
and U260 (N_260,In_2252,In_566);
nand U261 (N_261,In_2313,In_2172);
or U262 (N_262,In_598,In_981);
or U263 (N_263,In_134,In_1045);
and U264 (N_264,In_956,In_912);
nand U265 (N_265,In_716,In_2962);
and U266 (N_266,In_1393,In_622);
xnor U267 (N_267,In_1624,In_330);
xor U268 (N_268,In_1591,In_1210);
or U269 (N_269,In_414,In_2769);
and U270 (N_270,In_1422,In_1198);
nor U271 (N_271,In_169,In_1820);
nand U272 (N_272,In_2570,In_751);
nand U273 (N_273,In_1798,In_1261);
xor U274 (N_274,In_1772,In_870);
and U275 (N_275,In_2404,In_2562);
nor U276 (N_276,In_2602,In_884);
xor U277 (N_277,In_2828,In_2244);
and U278 (N_278,In_1696,In_326);
xor U279 (N_279,In_1615,In_2684);
or U280 (N_280,In_1848,In_2403);
nor U281 (N_281,In_538,In_831);
or U282 (N_282,In_2733,In_2751);
nand U283 (N_283,In_2254,In_809);
nor U284 (N_284,In_1847,In_1424);
nor U285 (N_285,In_922,In_2143);
nor U286 (N_286,In_192,In_668);
nor U287 (N_287,In_2521,In_632);
xnor U288 (N_288,In_1406,In_1494);
xnor U289 (N_289,In_1723,In_2379);
nand U290 (N_290,In_363,In_1887);
nor U291 (N_291,In_1604,In_1750);
or U292 (N_292,In_773,In_2075);
nor U293 (N_293,In_1600,In_1114);
and U294 (N_294,In_14,In_255);
or U295 (N_295,In_2144,In_43);
and U296 (N_296,In_2531,In_2050);
nand U297 (N_297,In_583,In_2836);
and U298 (N_298,In_2676,In_7);
and U299 (N_299,In_422,In_1417);
and U300 (N_300,In_1271,In_2870);
or U301 (N_301,In_2682,In_1903);
xor U302 (N_302,In_1332,In_1025);
or U303 (N_303,In_1298,In_2863);
nand U304 (N_304,In_1603,In_2922);
nor U305 (N_305,In_1171,In_2551);
nand U306 (N_306,In_1057,In_834);
or U307 (N_307,In_1474,In_644);
xnor U308 (N_308,In_2857,In_1666);
nand U309 (N_309,In_584,In_1259);
nand U310 (N_310,In_1914,In_2825);
nand U311 (N_311,In_2636,In_1050);
and U312 (N_312,In_1979,In_2307);
and U313 (N_313,In_1341,In_835);
and U314 (N_314,In_841,In_2469);
and U315 (N_315,In_2937,In_127);
and U316 (N_316,In_983,In_641);
or U317 (N_317,In_674,In_2755);
and U318 (N_318,In_1636,In_1969);
or U319 (N_319,In_532,In_698);
nand U320 (N_320,In_119,In_2009);
nand U321 (N_321,In_1654,In_1096);
xor U322 (N_322,In_2640,In_572);
xnor U323 (N_323,In_679,In_1187);
nand U324 (N_324,In_80,In_32);
and U325 (N_325,In_2461,In_325);
nor U326 (N_326,In_2260,In_1310);
nor U327 (N_327,In_71,In_2156);
and U328 (N_328,In_823,In_1965);
nand U329 (N_329,In_2014,In_2622);
and U330 (N_330,In_1119,In_980);
nand U331 (N_331,In_1463,In_1009);
or U332 (N_332,In_2206,In_1316);
or U333 (N_333,In_2523,In_749);
nor U334 (N_334,In_1966,In_957);
nand U335 (N_335,In_2188,In_2291);
nor U336 (N_336,In_149,In_2485);
nor U337 (N_337,In_1987,In_568);
and U338 (N_338,In_1669,In_2794);
or U339 (N_339,In_660,In_571);
and U340 (N_340,In_2620,In_129);
xnor U341 (N_341,In_864,In_2315);
or U342 (N_342,In_2815,In_1350);
nor U343 (N_343,In_1069,In_8);
xnor U344 (N_344,In_1910,In_1934);
xor U345 (N_345,In_1621,In_2710);
nand U346 (N_346,In_2706,In_399);
nand U347 (N_347,In_1748,In_635);
and U348 (N_348,In_2284,In_2389);
xnor U349 (N_349,In_2765,In_2429);
xor U350 (N_350,In_2181,In_1391);
or U351 (N_351,In_1131,In_1704);
or U352 (N_352,In_724,In_999);
xor U353 (N_353,In_89,In_873);
nor U354 (N_354,In_2505,In_2897);
and U355 (N_355,In_1893,In_2046);
nand U356 (N_356,In_480,In_2639);
nand U357 (N_357,In_1249,In_2193);
xnor U358 (N_358,In_846,In_2972);
nor U359 (N_359,In_2263,In_2838);
nand U360 (N_360,In_2536,In_2912);
nand U361 (N_361,In_1097,In_1599);
or U362 (N_362,In_1436,In_2135);
or U363 (N_363,In_319,In_2719);
nand U364 (N_364,In_12,In_2518);
xor U365 (N_365,In_945,In_1209);
nand U366 (N_366,In_2585,In_1173);
nand U367 (N_367,In_1030,In_51);
xnor U368 (N_368,In_1813,In_613);
xnor U369 (N_369,In_756,In_2333);
nor U370 (N_370,In_2165,In_2109);
nor U371 (N_371,In_343,In_551);
xnor U372 (N_372,In_2680,In_2596);
nand U373 (N_373,In_947,In_2270);
or U374 (N_374,In_1567,In_2419);
nand U375 (N_375,In_1670,In_721);
nor U376 (N_376,In_2353,In_1076);
and U377 (N_377,In_2210,In_515);
or U378 (N_378,In_2550,In_711);
xnor U379 (N_379,In_2123,In_454);
or U380 (N_380,In_1435,In_1138);
xor U381 (N_381,In_777,In_2754);
nand U382 (N_382,In_2675,In_2809);
and U383 (N_383,In_2974,In_1746);
or U384 (N_384,In_307,In_1081);
xor U385 (N_385,In_1962,In_1905);
or U386 (N_386,In_2527,In_1299);
xnor U387 (N_387,In_1970,In_2178);
xor U388 (N_388,In_1383,In_508);
nor U389 (N_389,In_443,In_581);
or U390 (N_390,In_898,In_1147);
nand U391 (N_391,In_1027,In_2455);
nand U392 (N_392,In_1067,In_1143);
and U393 (N_393,In_2820,In_1314);
or U394 (N_394,In_2186,In_1508);
or U395 (N_395,In_2655,In_289);
nor U396 (N_396,In_1545,In_1357);
and U397 (N_397,In_2250,In_2327);
xor U398 (N_398,In_2854,In_62);
nand U399 (N_399,In_1540,In_1411);
and U400 (N_400,In_2978,In_1222);
xor U401 (N_401,In_516,In_2115);
nor U402 (N_402,In_1897,In_879);
nand U403 (N_403,In_899,In_2157);
or U404 (N_404,In_1331,In_2454);
nand U405 (N_405,In_779,In_124);
xnor U406 (N_406,In_570,In_882);
or U407 (N_407,In_196,In_1082);
and U408 (N_408,In_2246,In_1270);
or U409 (N_409,In_1646,In_382);
and U410 (N_410,In_2873,In_1123);
xnor U411 (N_411,In_2775,In_2761);
and U412 (N_412,In_863,In_22);
and U413 (N_413,In_2945,In_1931);
and U414 (N_414,In_1227,In_2928);
or U415 (N_415,In_2557,In_1185);
xnor U416 (N_416,In_2408,In_953);
or U417 (N_417,In_2446,In_546);
and U418 (N_418,In_2893,In_565);
or U419 (N_419,In_2763,In_2021);
xor U420 (N_420,In_2624,In_822);
or U421 (N_421,In_1695,In_2920);
nor U422 (N_422,In_153,In_2384);
nand U423 (N_423,In_2954,In_2669);
xnor U424 (N_424,In_2532,In_1294);
nand U425 (N_425,In_2544,In_1005);
or U426 (N_426,In_2708,In_1090);
nor U427 (N_427,In_705,In_2220);
and U428 (N_428,In_599,In_59);
nand U429 (N_429,In_643,In_270);
nor U430 (N_430,In_791,In_44);
or U431 (N_431,In_216,In_1616);
or U432 (N_432,In_994,In_1140);
and U433 (N_433,In_245,In_869);
nor U434 (N_434,In_2537,In_2789);
and U435 (N_435,In_57,In_2558);
nand U436 (N_436,In_429,In_103);
nand U437 (N_437,In_854,In_2439);
xor U438 (N_438,In_1401,In_2073);
nand U439 (N_439,In_2683,In_1655);
xor U440 (N_440,In_464,In_2524);
and U441 (N_441,In_2459,In_2402);
nor U442 (N_442,In_2331,In_2997);
xor U443 (N_443,In_2992,In_1824);
xnor U444 (N_444,In_2299,In_560);
nor U445 (N_445,In_2490,In_597);
xnor U446 (N_446,In_1301,In_1843);
and U447 (N_447,In_2079,In_1255);
nor U448 (N_448,In_97,In_55);
and U449 (N_449,In_915,In_2038);
and U450 (N_450,In_1054,In_1246);
xnor U451 (N_451,In_320,In_2716);
and U452 (N_452,In_2287,In_378);
nand U453 (N_453,In_2807,In_1317);
nor U454 (N_454,In_1759,In_2590);
nand U455 (N_455,In_1493,In_2930);
nor U456 (N_456,In_1200,In_1323);
and U457 (N_457,In_923,In_372);
or U458 (N_458,In_1205,In_240);
nand U459 (N_459,In_1376,In_2709);
or U460 (N_460,In_391,In_374);
nand U461 (N_461,In_1447,In_2269);
nor U462 (N_462,In_2642,In_2613);
xnor U463 (N_463,In_2035,In_741);
nor U464 (N_464,In_23,In_1522);
nor U465 (N_465,In_631,In_1906);
or U466 (N_466,In_2895,In_2187);
nand U467 (N_467,In_1480,In_496);
xnor U468 (N_468,In_2907,In_848);
or U469 (N_469,In_667,In_1340);
and U470 (N_470,In_1547,In_1714);
nand U471 (N_471,In_1170,In_2348);
or U472 (N_472,In_2884,In_1473);
or U473 (N_473,In_2512,In_2955);
and U474 (N_474,In_2139,In_772);
nor U475 (N_475,In_2378,In_842);
nand U476 (N_476,In_1823,In_233);
or U477 (N_477,In_1019,In_2633);
xnor U478 (N_478,In_2480,In_628);
and U479 (N_479,In_2692,In_689);
nand U480 (N_480,In_1647,In_2179);
nor U481 (N_481,In_1789,In_2615);
or U482 (N_482,In_437,In_881);
xnor U483 (N_483,In_1991,In_10);
nor U484 (N_484,In_253,In_1495);
nor U485 (N_485,In_2964,In_1819);
or U486 (N_486,In_2100,In_342);
nand U487 (N_487,In_2813,In_2853);
nor U488 (N_488,In_780,In_633);
nand U489 (N_489,In_503,In_1950);
nor U490 (N_490,In_1303,In_2871);
and U491 (N_491,In_1216,In_1908);
xnor U492 (N_492,In_1127,In_1944);
xnor U493 (N_493,In_193,In_1656);
and U494 (N_494,In_2204,In_2935);
and U495 (N_495,In_2832,In_2420);
xor U496 (N_496,In_2368,In_2229);
nand U497 (N_497,In_2033,In_2840);
or U498 (N_498,In_1457,In_274);
xnor U499 (N_499,In_456,In_759);
nand U500 (N_500,In_1989,In_995);
or U501 (N_501,In_1104,In_2717);
or U502 (N_502,In_475,In_961);
nor U503 (N_503,In_2561,In_590);
nor U504 (N_504,In_1487,In_1380);
nor U505 (N_505,In_525,In_444);
or U506 (N_506,In_1016,In_2294);
nor U507 (N_507,In_861,In_1863);
nand U508 (N_508,In_800,In_2324);
xor U509 (N_509,In_2541,In_2511);
and U510 (N_510,In_2919,In_384);
and U511 (N_511,In_2625,In_2606);
and U512 (N_512,In_1053,In_2077);
and U513 (N_513,In_1658,In_531);
and U514 (N_514,In_50,In_1403);
and U515 (N_515,In_333,In_1634);
nor U516 (N_516,In_2383,In_2730);
nor U517 (N_517,In_1012,In_2004);
nand U518 (N_518,In_1570,In_2437);
nor U519 (N_519,In_2589,In_162);
nand U520 (N_520,In_747,In_927);
nor U521 (N_521,In_1297,In_1676);
or U522 (N_522,In_2554,In_2711);
and U523 (N_523,In_1755,In_1364);
or U524 (N_524,In_984,In_476);
xnor U525 (N_525,In_1037,In_1652);
nand U526 (N_526,In_2808,In_2721);
xnor U527 (N_527,In_2860,In_1775);
or U528 (N_528,In_2739,In_1583);
nor U529 (N_529,In_1717,In_1400);
xnor U530 (N_530,In_1892,In_2913);
nor U531 (N_531,In_315,In_2423);
or U532 (N_532,In_1049,In_648);
nand U533 (N_533,In_2756,In_2373);
nor U534 (N_534,In_845,In_1498);
nor U535 (N_535,In_2479,In_2901);
nand U536 (N_536,In_2704,In_2357);
nor U537 (N_537,In_1553,In_1702);
nand U538 (N_538,In_371,In_851);
or U539 (N_539,In_2567,In_1203);
xor U540 (N_540,In_542,In_260);
nand U541 (N_541,In_576,In_2170);
and U542 (N_542,In_2247,In_1361);
nor U543 (N_543,In_1534,In_896);
nand U544 (N_544,In_1388,In_477);
and U545 (N_545,In_802,In_2350);
nand U546 (N_546,In_2332,In_517);
and U547 (N_547,In_174,In_671);
nand U548 (N_548,In_1055,In_331);
and U549 (N_549,In_2595,In_359);
nor U550 (N_550,In_2724,In_2658);
xor U551 (N_551,In_2234,In_2161);
and U552 (N_552,In_596,In_2169);
and U553 (N_553,In_2725,In_2983);
and U554 (N_554,In_1559,In_2497);
nor U555 (N_555,In_2013,In_2317);
nand U556 (N_556,In_2146,In_1774);
or U557 (N_557,In_768,In_616);
nand U558 (N_558,In_2834,In_1806);
nand U559 (N_559,In_1420,In_1369);
nand U560 (N_560,In_2506,In_2235);
and U561 (N_561,In_2956,In_5);
or U562 (N_562,In_1633,In_2528);
or U563 (N_563,In_2823,In_128);
or U564 (N_564,In_819,In_1042);
xnor U565 (N_565,In_1324,In_1609);
nand U566 (N_566,In_1161,In_292);
nand U567 (N_567,In_466,In_2628);
nor U568 (N_568,In_252,In_2285);
nor U569 (N_569,In_2991,In_1164);
nor U570 (N_570,In_1100,In_2646);
nor U571 (N_571,In_1146,In_1113);
and U572 (N_572,In_1995,In_277);
xor U573 (N_573,In_99,In_1898);
nand U574 (N_574,In_362,In_1024);
nor U575 (N_575,In_2369,In_2876);
nand U576 (N_576,In_549,In_236);
nand U577 (N_577,In_2335,In_2892);
xnor U578 (N_578,In_2395,In_1546);
and U579 (N_579,In_1993,In_612);
or U580 (N_580,In_778,In_2830);
and U581 (N_581,In_2722,In_2852);
or U582 (N_582,In_349,In_1983);
xor U583 (N_583,In_1329,In_165);
or U584 (N_584,In_920,In_2142);
or U585 (N_585,In_77,In_1087);
xor U586 (N_586,In_593,In_2654);
xnor U587 (N_587,In_1169,In_2598);
nand U588 (N_588,In_2608,In_2272);
or U589 (N_589,In_606,In_2783);
and U590 (N_590,In_2001,In_2005);
nor U591 (N_591,In_1926,In_306);
nand U592 (N_592,In_1144,In_2283);
xor U593 (N_593,In_2996,In_83);
nand U594 (N_594,In_1674,In_2215);
nand U595 (N_595,In_167,In_275);
nor U596 (N_596,In_1536,In_872);
xnor U597 (N_597,In_1555,In_1912);
or U598 (N_598,In_1861,In_2514);
nor U599 (N_599,In_2701,In_2686);
or U600 (N_600,In_2614,In_1288);
and U601 (N_601,In_1345,In_1786);
or U602 (N_602,In_2082,In_484);
xnor U603 (N_603,In_729,In_1174);
xor U604 (N_604,In_2508,In_692);
nor U605 (N_605,In_2338,In_2026);
nand U606 (N_606,In_2087,In_2151);
nand U607 (N_607,In_199,In_680);
and U608 (N_608,In_579,In_710);
nand U609 (N_609,In_2844,In_180);
nor U610 (N_610,In_2427,In_790);
nor U611 (N_611,In_946,In_552);
and U612 (N_612,In_2902,In_707);
nand U613 (N_613,In_2998,In_1882);
nor U614 (N_614,In_2310,In_188);
xor U615 (N_615,In_2183,In_730);
nand U616 (N_616,In_2500,In_2104);
and U617 (N_617,In_370,In_105);
nand U618 (N_618,In_1243,In_1102);
and U619 (N_619,In_1657,In_1730);
or U620 (N_620,In_2817,In_665);
nand U621 (N_621,In_2464,In_2883);
and U622 (N_622,In_666,In_1869);
nor U623 (N_623,In_1451,In_210);
xnor U624 (N_624,In_862,In_1507);
nor U625 (N_625,In_2948,In_2286);
nand U626 (N_626,In_1721,In_2406);
or U627 (N_627,In_2773,In_1751);
xnor U628 (N_628,In_300,In_2476);
or U629 (N_629,In_951,In_1352);
nor U630 (N_630,In_2810,In_1242);
nand U631 (N_631,In_1974,In_2522);
or U632 (N_632,In_960,In_1980);
nand U633 (N_633,In_248,In_1384);
nor U634 (N_634,In_1909,In_2742);
or U635 (N_635,In_1221,In_833);
and U636 (N_636,In_685,In_761);
and U637 (N_637,In_1267,In_1692);
and U638 (N_638,In_2826,In_426);
nor U639 (N_639,In_2358,In_557);
xnor U640 (N_640,In_1825,In_2586);
and U641 (N_641,In_186,In_2941);
xnor U642 (N_642,In_2398,In_1450);
nor U643 (N_643,In_1366,In_269);
nand U644 (N_644,In_1781,In_2600);
or U645 (N_645,In_1273,In_434);
or U646 (N_646,In_1535,In_2303);
nand U647 (N_647,In_2980,In_354);
nand U648 (N_648,In_1046,In_1405);
nand U649 (N_649,In_1300,In_340);
nand U650 (N_650,In_2034,In_2985);
nand U651 (N_651,In_2472,In_615);
or U652 (N_652,In_2474,In_2070);
nand U653 (N_653,In_695,In_1687);
nor U654 (N_654,In_2939,In_148);
xor U655 (N_655,In_2594,In_1484);
nor U656 (N_656,In_279,In_1472);
xor U657 (N_657,In_629,In_1582);
nand U658 (N_658,In_2471,In_1008);
nor U659 (N_659,In_173,In_2176);
nand U660 (N_660,In_1023,In_1444);
or U661 (N_661,In_782,In_1921);
nand U662 (N_662,In_1533,In_2288);
nor U663 (N_663,In_175,In_108);
or U664 (N_664,In_1642,In_1328);
nor U665 (N_665,In_661,In_1946);
nor U666 (N_666,In_1020,In_958);
xor U667 (N_667,In_888,In_649);
xnor U668 (N_668,In_524,In_2124);
nand U669 (N_669,In_433,In_812);
or U670 (N_670,In_2153,In_2572);
nand U671 (N_671,In_1196,In_1126);
and U672 (N_672,In_766,In_709);
nand U673 (N_673,In_1856,In_17);
xnor U674 (N_674,In_930,In_195);
nor U675 (N_675,In_2022,In_2120);
xnor U676 (N_676,In_197,In_1618);
xnor U677 (N_677,In_1563,In_985);
and U678 (N_678,In_1110,In_703);
nor U679 (N_679,In_2257,In_924);
nor U680 (N_680,In_224,In_13);
or U681 (N_681,In_223,In_417);
nand U682 (N_682,In_2069,In_1031);
xor U683 (N_683,In_592,In_2148);
and U684 (N_684,In_2059,In_1999);
and U685 (N_685,In_2816,In_2597);
xnor U686 (N_686,In_2890,In_25);
xor U687 (N_687,In_505,In_1967);
nor U688 (N_688,In_1006,In_2509);
or U689 (N_689,In_2372,In_2105);
nor U690 (N_690,In_250,In_678);
or U691 (N_691,In_226,In_856);
xnor U692 (N_692,In_1631,In_1454);
xnor U693 (N_693,In_1475,In_1639);
xor U694 (N_694,In_1220,In_2006);
nor U695 (N_695,In_2782,In_2715);
and U696 (N_696,In_2647,In_258);
or U697 (N_697,In_104,In_806);
and U698 (N_698,In_2743,In_2914);
and U699 (N_699,In_2970,In_653);
nor U700 (N_700,In_630,In_507);
nand U701 (N_701,In_2221,In_621);
nor U702 (N_702,In_784,In_1549);
nor U703 (N_703,In_547,In_1182);
nor U704 (N_704,In_1805,In_1681);
xor U705 (N_705,In_2097,In_2781);
nor U706 (N_706,In_318,In_2539);
or U707 (N_707,In_1858,In_2155);
and U708 (N_708,In_2915,In_2650);
xnor U709 (N_709,In_825,In_1528);
or U710 (N_710,In_1075,In_2066);
and U711 (N_711,In_1742,In_112);
nor U712 (N_712,In_1335,In_1231);
xor U713 (N_713,In_2689,In_604);
and U714 (N_714,In_1026,In_639);
nand U715 (N_715,In_1342,In_522);
and U716 (N_716,In_9,In_73);
nor U717 (N_717,In_283,In_266);
or U718 (N_718,In_589,In_54);
or U719 (N_719,In_1141,In_2091);
or U720 (N_720,In_500,In_2356);
xnor U721 (N_721,In_2410,In_1886);
nand U722 (N_722,In_2354,In_1506);
nand U723 (N_723,In_569,In_1043);
nor U724 (N_724,In_1826,In_601);
xor U725 (N_725,In_1372,In_1557);
and U726 (N_726,In_2425,In_2575);
or U727 (N_727,In_2891,In_1374);
nand U728 (N_728,In_457,In_1428);
or U729 (N_729,In_1949,In_2949);
and U730 (N_730,In_2645,In_1483);
nand U731 (N_731,In_1263,In_2971);
xor U732 (N_732,In_1645,In_2243);
xnor U733 (N_733,In_1389,In_2565);
and U734 (N_734,In_2342,In_2931);
nor U735 (N_735,In_2344,In_1753);
nor U736 (N_736,In_425,In_2213);
xnor U737 (N_737,In_191,In_79);
nand U738 (N_738,In_2319,In_2502);
nor U739 (N_739,In_2750,In_2442);
xnor U740 (N_740,In_2874,In_238);
nor U741 (N_741,In_244,In_704);
xor U742 (N_742,In_2681,In_1602);
xor U743 (N_743,In_358,In_2483);
nor U744 (N_744,In_448,In_1531);
nor U745 (N_745,In_1460,In_2202);
xor U746 (N_746,In_2588,In_623);
nand U747 (N_747,In_794,In_1686);
and U748 (N_748,In_251,In_2424);
xnor U749 (N_749,In_1550,In_304);
and U750 (N_750,In_2031,In_2609);
and U751 (N_751,In_40,In_1449);
nand U752 (N_752,In_1524,In_1410);
nor U753 (N_753,In_1735,In_1638);
and U754 (N_754,In_141,In_1194);
and U755 (N_755,In_1822,In_987);
nor U756 (N_756,In_1157,In_744);
nor U757 (N_757,In_1033,In_1343);
xor U758 (N_758,In_2764,In_646);
or U759 (N_759,In_933,In_98);
nand U760 (N_760,In_1577,In_285);
or U761 (N_761,In_1088,In_2076);
and U762 (N_762,In_1168,In_1763);
nand U763 (N_763,In_2460,In_990);
nand U764 (N_764,In_468,In_719);
nor U765 (N_765,In_2278,In_1940);
nand U766 (N_766,In_2693,In_1320);
xnor U767 (N_767,In_117,In_1849);
or U768 (N_768,In_2534,In_1708);
or U769 (N_769,In_2434,In_1918);
xnor U770 (N_770,In_256,In_1757);
or U771 (N_771,In_494,In_2592);
nor U772 (N_772,In_220,In_2295);
nor U773 (N_773,In_2685,In_1150);
xnor U774 (N_774,In_1201,In_902);
xnor U775 (N_775,In_1041,In_795);
xnor U776 (N_776,In_2555,In_1290);
or U777 (N_777,In_161,In_645);
and U778 (N_778,In_1941,In_78);
nor U779 (N_779,In_2661,In_2496);
nor U780 (N_780,In_2923,In_1179);
and U781 (N_781,In_1223,In_2851);
and U782 (N_782,In_228,In_39);
nand U783 (N_783,In_2036,In_561);
xor U784 (N_784,In_591,In_832);
and U785 (N_785,In_890,In_365);
nor U786 (N_786,In_2994,In_1226);
nor U787 (N_787,In_1626,In_816);
xnor U788 (N_788,In_889,In_1426);
nor U789 (N_789,In_2433,In_2277);
and U790 (N_790,In_2060,In_682);
xnor U791 (N_791,In_843,In_625);
and U792 (N_792,In_895,In_2936);
and U793 (N_793,In_303,In_2280);
and U794 (N_794,In_2239,In_2699);
nor U795 (N_795,In_676,In_74);
and U796 (N_796,In_280,In_2947);
or U797 (N_797,In_2968,In_2386);
and U798 (N_798,In_1080,In_2879);
or U799 (N_799,In_836,In_2160);
nand U800 (N_800,In_1257,In_2162);
or U801 (N_801,In_2167,In_904);
and U802 (N_802,In_2607,In_1874);
and U803 (N_803,In_2989,In_555);
nand U804 (N_804,In_1942,In_144);
nand U805 (N_805,In_56,In_211);
nand U806 (N_806,In_619,In_1778);
or U807 (N_807,In_1035,In_271);
or U808 (N_808,In_1151,In_452);
xor U809 (N_809,In_1589,In_762);
nand U810 (N_810,In_2771,In_880);
or U811 (N_811,In_699,In_1013);
nand U812 (N_812,In_1262,In_2397);
xor U813 (N_813,In_2375,In_347);
nor U814 (N_814,In_1935,In_1722);
nor U815 (N_815,In_467,In_941);
or U816 (N_816,In_2435,In_1588);
and U817 (N_817,In_486,In_2045);
and U818 (N_818,In_305,In_2885);
nand U819 (N_819,In_2800,In_1189);
and U820 (N_820,In_600,In_2309);
nor U821 (N_821,In_2086,In_2281);
nand U822 (N_822,In_1373,In_1707);
and U823 (N_823,In_916,In_1321);
nand U824 (N_824,In_2211,In_2456);
nand U825 (N_825,In_1576,In_2248);
xor U826 (N_826,In_1418,In_1700);
nand U827 (N_827,In_445,In_1197);
nor U828 (N_828,In_2067,In_397);
and U829 (N_829,In_1538,In_805);
nor U830 (N_830,In_849,In_1175);
and U831 (N_831,In_652,In_420);
nor U832 (N_832,In_541,In_2792);
nor U833 (N_833,In_1948,In_1719);
or U834 (N_834,In_548,In_1386);
or U835 (N_835,In_1099,In_102);
and U836 (N_836,In_1911,In_2703);
xnor U837 (N_837,In_2547,In_2138);
xnor U838 (N_838,In_1236,In_2488);
nor U839 (N_839,In_1315,In_976);
or U840 (N_840,In_929,In_1121);
or U841 (N_841,In_1868,In_1091);
and U842 (N_842,In_2776,In_1204);
nand U843 (N_843,In_1269,In_2337);
or U844 (N_844,In_2924,In_2667);
nor U845 (N_845,In_1371,In_2869);
xor U846 (N_846,In_2966,In_1776);
or U847 (N_847,In_2381,In_459);
or U848 (N_848,In_1787,In_2638);
and U849 (N_849,In_2478,In_2224);
nand U850 (N_850,In_1133,In_2687);
xor U851 (N_851,In_1501,In_2520);
and U852 (N_852,In_2631,In_2894);
nand U853 (N_853,In_1811,In_410);
xor U854 (N_854,In_2768,In_2925);
and U855 (N_855,In_2767,In_2088);
nor U856 (N_856,In_2205,In_580);
nand U857 (N_857,In_125,In_1562);
nand U858 (N_858,In_37,In_713);
and U859 (N_859,In_2040,In_801);
and U860 (N_860,In_2057,In_2858);
and U861 (N_861,In_2981,In_1523);
nor U862 (N_862,In_2484,In_728);
nor U863 (N_863,In_1412,In_1505);
or U864 (N_864,In_2037,In_339);
and U865 (N_865,In_133,In_595);
nand U866 (N_866,In_2296,In_1070);
nand U867 (N_867,In_1928,In_337);
nor U868 (N_868,In_2940,In_2938);
and U869 (N_869,In_894,In_926);
or U870 (N_870,In_1149,In_1963);
or U871 (N_871,In_2855,In_658);
xor U872 (N_872,In_693,In_66);
xnor U873 (N_873,In_282,In_1056);
nor U874 (N_874,In_1491,In_1471);
or U875 (N_875,In_1952,In_2848);
xnor U876 (N_876,In_2977,In_2195);
nand U877 (N_877,In_2414,In_781);
or U878 (N_878,In_1877,In_739);
nor U879 (N_879,In_491,In_140);
nor U880 (N_880,In_154,In_247);
or U881 (N_881,In_1902,In_1040);
or U882 (N_882,In_2905,In_2909);
xnor U883 (N_883,In_1431,In_1101);
xnor U884 (N_884,In_2486,In_702);
xor U885 (N_885,In_1036,In_2530);
and U886 (N_886,In_2626,In_65);
nand U887 (N_887,In_1857,In_582);
xnor U888 (N_888,In_2265,In_1632);
xor U889 (N_889,In_2462,In_609);
nand U890 (N_890,In_2242,In_1866);
and U891 (N_891,In_19,In_787);
nand U892 (N_892,In_431,In_1558);
and U893 (N_893,In_2116,In_1871);
and U894 (N_894,In_2833,In_1671);
nand U895 (N_895,In_1414,In_1566);
and U896 (N_896,In_2649,In_733);
or U897 (N_897,In_1982,In_1803);
xnor U898 (N_898,In_936,In_1232);
nor U899 (N_899,In_1957,In_205);
nor U900 (N_900,In_1693,In_35);
nor U901 (N_901,In_2617,In_2621);
nand U902 (N_902,In_2491,In_1694);
xnor U903 (N_903,In_2641,In_2696);
nor U904 (N_904,In_2030,In_1900);
and U905 (N_905,In_1467,In_2657);
nor U906 (N_906,In_2886,In_758);
nor U907 (N_907,In_1234,In_395);
nand U908 (N_908,In_2290,In_1701);
xnor U909 (N_909,In_2542,In_2566);
xnor U910 (N_910,In_1754,In_2101);
nor U911 (N_911,In_146,In_2785);
xor U912 (N_912,In_1339,In_2092);
nor U913 (N_913,In_2943,In_2784);
nand U914 (N_914,In_1581,In_2430);
and U915 (N_915,In_368,In_785);
or U916 (N_916,In_1360,In_1015);
xnor U917 (N_917,In_2112,In_514);
and U918 (N_918,In_2728,In_114);
and U919 (N_919,In_2668,In_691);
and U920 (N_920,In_992,In_2111);
nor U921 (N_921,In_900,In_764);
xnor U922 (N_922,In_2282,In_2432);
nand U923 (N_923,In_2535,In_1413);
xor U924 (N_924,In_2412,In_683);
nor U925 (N_925,In_963,In_1607);
xor U926 (N_926,In_1228,In_221);
nand U927 (N_927,In_1145,In_1500);
xnor U928 (N_928,In_164,In_2864);
xor U929 (N_929,In_829,In_2990);
xnor U930 (N_930,In_2982,In_1630);
nor U931 (N_931,In_796,In_26);
xnor U932 (N_932,In_2129,In_2392);
xnor U933 (N_933,In_2952,In_241);
nand U934 (N_934,In_1407,In_1230);
nor U935 (N_935,In_2236,In_2102);
and U936 (N_936,In_1038,In_752);
and U937 (N_937,In_934,In_1306);
or U938 (N_938,In_1784,In_2325);
xor U939 (N_939,In_1817,In_526);
nand U940 (N_940,In_1808,In_1398);
xnor U941 (N_941,In_575,In_2556);
nand U942 (N_942,In_2746,In_346);
xnor U943 (N_943,In_2048,In_366);
and U944 (N_944,In_2495,In_328);
nor U945 (N_945,In_2264,In_979);
nor U946 (N_946,In_2753,In_2988);
or U947 (N_947,In_2426,In_2672);
and U948 (N_948,In_1663,In_840);
or U949 (N_949,In_1738,In_2818);
xor U950 (N_950,In_970,In_68);
nand U951 (N_951,In_398,In_614);
nand U952 (N_952,In_545,In_2559);
nor U953 (N_953,In_1094,In_155);
or U954 (N_954,In_574,In_2158);
nor U955 (N_955,In_227,In_212);
and U956 (N_956,In_624,In_2266);
nor U957 (N_957,In_2359,In_573);
nand U958 (N_958,In_369,In_1018);
or U959 (N_959,In_2147,In_2271);
nand U960 (N_960,In_2175,In_2249);
and U961 (N_961,In_1044,In_1733);
xor U962 (N_962,In_2644,In_2839);
or U963 (N_963,In_748,In_1421);
xnor U964 (N_964,In_2385,In_1077);
and U965 (N_965,In_1569,In_1812);
and U966 (N_966,In_2916,In_2192);
nor U967 (N_967,In_783,In_215);
or U968 (N_968,In_298,In_2582);
or U969 (N_969,In_24,In_944);
or U970 (N_970,In_2062,In_2993);
and U971 (N_971,In_1409,In_242);
or U972 (N_972,In_423,In_2043);
nand U973 (N_973,In_1539,In_28);
nor U974 (N_974,In_2261,In_1111);
xor U975 (N_975,In_2846,In_234);
or U976 (N_976,In_1427,In_2117);
nor U977 (N_977,In_131,In_1959);
and U978 (N_978,In_447,In_798);
nand U979 (N_979,In_2311,In_1565);
or U980 (N_980,In_2065,In_2632);
nand U981 (N_981,In_1441,In_659);
nor U982 (N_982,In_1532,In_1516);
and U983 (N_983,In_940,In_2399);
nor U984 (N_984,In_1984,In_1181);
and U985 (N_985,In_2516,In_1841);
nor U986 (N_986,In_640,In_738);
and U987 (N_987,In_1831,In_69);
xnor U988 (N_988,In_421,In_471);
nand U989 (N_989,In_1387,In_687);
or U990 (N_990,In_2438,In_1489);
or U991 (N_991,In_2517,In_2543);
nand U992 (N_992,In_770,In_875);
nand U993 (N_993,In_76,In_2847);
nand U994 (N_994,In_1453,In_435);
and U995 (N_995,In_1572,In_1172);
nand U996 (N_996,In_403,In_1913);
nand U997 (N_997,In_2786,In_1394);
or U998 (N_998,In_379,In_974);
nor U999 (N_999,In_1517,In_950);
xor U1000 (N_1000,N_413,In_2177);
and U1001 (N_1001,In_405,N_243);
xnor U1002 (N_1002,N_734,N_180);
nand U1003 (N_1003,In_63,In_2174);
nor U1004 (N_1004,N_195,N_602);
nand U1005 (N_1005,In_767,In_1011);
and U1006 (N_1006,In_1915,In_2166);
nor U1007 (N_1007,N_597,In_1867);
xnor U1008 (N_1008,In_2553,N_307);
nand U1009 (N_1009,N_783,N_309);
nor U1010 (N_1010,In_1272,N_666);
and U1011 (N_1011,In_509,N_650);
nand U1012 (N_1012,N_760,In_2098);
nand U1013 (N_1013,N_313,In_201);
nand U1014 (N_1014,In_1291,In_967);
nand U1015 (N_1015,In_1064,In_1192);
nor U1016 (N_1016,N_792,N_172);
or U1017 (N_1017,In_348,N_619);
nand U1018 (N_1018,In_290,N_160);
nor U1019 (N_1019,N_516,In_1136);
nand U1020 (N_1020,In_479,In_2445);
nand U1021 (N_1021,In_1177,In_2950);
and U1022 (N_1022,N_963,In_2900);
nor U1023 (N_1023,N_794,In_1002);
and U1024 (N_1024,N_782,In_529);
xnor U1025 (N_1025,N_627,In_937);
xnor U1026 (N_1026,N_838,In_535);
or U1027 (N_1027,N_441,N_349);
and U1028 (N_1028,N_612,N_337);
nor U1029 (N_1029,N_940,In_416);
nor U1030 (N_1030,N_480,In_1637);
nand U1031 (N_1031,N_559,N_374);
nor U1032 (N_1032,N_442,In_803);
nor U1033 (N_1033,In_734,N_984);
xor U1034 (N_1034,In_1809,In_2824);
xnor U1035 (N_1035,N_862,N_887);
and U1036 (N_1036,N_410,N_434);
nor U1037 (N_1037,N_819,In_1990);
or U1038 (N_1038,N_118,In_2841);
nand U1039 (N_1039,N_467,N_250);
and U1040 (N_1040,N_644,N_146);
nand U1041 (N_1041,In_2872,N_830);
xnor U1042 (N_1042,N_424,N_561);
or U1043 (N_1043,In_988,N_923);
nand U1044 (N_1044,In_2552,N_563);
xnor U1045 (N_1045,In_1542,In_2388);
xor U1046 (N_1046,N_755,N_385);
xor U1047 (N_1047,In_2778,In_701);
nor U1048 (N_1048,In_708,In_1322);
nand U1049 (N_1049,In_1933,N_883);
and U1050 (N_1050,N_124,N_71);
or U1051 (N_1051,In_498,In_1953);
nand U1052 (N_1052,N_197,In_1862);
nor U1053 (N_1053,N_431,N_128);
nor U1054 (N_1054,In_121,In_1782);
nor U1055 (N_1055,In_712,In_2468);
nand U1056 (N_1056,In_2875,In_297);
xor U1057 (N_1057,In_2255,In_2141);
xor U1058 (N_1058,N_852,N_658);
and U1059 (N_1059,In_402,N_873);
nor U1060 (N_1060,N_73,N_111);
xor U1061 (N_1061,In_1459,N_556);
or U1062 (N_1062,N_969,N_170);
and U1063 (N_1063,In_1355,N_452);
and U1064 (N_1064,N_248,N_227);
xor U1065 (N_1065,N_70,N_870);
or U1066 (N_1066,In_603,N_475);
xnor U1067 (N_1067,N_922,In_1739);
nand U1068 (N_1068,In_694,N_564);
or U1069 (N_1069,In_1610,N_19);
or U1070 (N_1070,In_1937,In_1309);
nand U1071 (N_1071,In_2083,In_411);
nand U1072 (N_1072,In_818,In_2346);
nand U1073 (N_1073,N_395,In_1152);
and U1074 (N_1074,In_1699,N_295);
nand U1075 (N_1075,In_726,In_2934);
nor U1076 (N_1076,In_2921,In_482);
nor U1077 (N_1077,In_1183,In_1768);
and U1078 (N_1078,N_353,In_2777);
xnor U1079 (N_1079,In_418,In_1253);
nand U1080 (N_1080,N_24,In_740);
nor U1081 (N_1081,In_1832,In_1084);
or U1082 (N_1082,In_2908,N_525);
nor U1083 (N_1083,N_29,In_225);
or U1084 (N_1084,In_2673,In_921);
and U1085 (N_1085,In_2440,N_554);
xor U1086 (N_1086,N_292,In_847);
xnor U1087 (N_1087,N_266,N_7);
nor U1088 (N_1088,In_775,In_745);
or U1089 (N_1089,N_207,In_2308);
nor U1090 (N_1090,N_801,In_1875);
nand U1091 (N_1091,N_457,In_2803);
xnor U1092 (N_1092,In_1496,N_506);
or U1093 (N_1093,In_1125,N_526);
nor U1094 (N_1094,N_717,N_171);
nor U1095 (N_1095,In_2318,In_2545);
nand U1096 (N_1096,In_1502,In_1668);
nand U1097 (N_1097,In_1554,In_294);
and U1098 (N_1098,In_142,N_583);
nand U1099 (N_1099,N_25,In_2702);
nor U1100 (N_1100,In_839,N_610);
and U1101 (N_1101,In_1643,N_636);
xnor U1102 (N_1102,N_592,In_2095);
and U1103 (N_1103,In_2969,N_121);
nand U1104 (N_1104,In_2911,In_2623);
xor U1105 (N_1105,N_150,N_509);
nor U1106 (N_1106,In_897,In_1325);
or U1107 (N_1107,In_11,In_2616);
nor U1108 (N_1108,In_1520,N_296);
xnor U1109 (N_1109,In_404,In_725);
or U1110 (N_1110,N_481,In_1208);
or U1111 (N_1111,In_1790,N_803);
or U1112 (N_1112,N_914,In_2304);
nand U1113 (N_1113,N_703,N_331);
nor U1114 (N_1114,N_420,In_170);
and U1115 (N_1115,N_897,In_1499);
nor U1116 (N_1116,In_1093,N_938);
nor U1117 (N_1117,N_977,In_973);
nor U1118 (N_1118,N_934,N_761);
nand U1119 (N_1119,In_1017,N_302);
or U1120 (N_1120,N_912,N_59);
and U1121 (N_1121,N_367,In_1810);
nor U1122 (N_1122,N_728,In_2343);
xor U1123 (N_1123,In_147,N_909);
xnor U1124 (N_1124,In_1509,In_2012);
nor U1125 (N_1125,N_138,In_675);
nor U1126 (N_1126,In_2305,In_2360);
nor U1127 (N_1127,N_461,In_1711);
nor U1128 (N_1128,N_492,In_2513);
or U1129 (N_1129,N_901,In_1264);
nand U1130 (N_1130,N_341,N_642);
nor U1131 (N_1131,N_244,N_523);
or U1132 (N_1132,N_423,N_436);
or U1133 (N_1133,In_1992,In_412);
xor U1134 (N_1134,In_1837,N_918);
nor U1135 (N_1135,In_1108,N_289);
and U1136 (N_1136,N_291,In_815);
nor U1137 (N_1137,N_212,N_188);
or U1138 (N_1138,In_1481,In_407);
nor U1139 (N_1139,N_275,In_1021);
and U1140 (N_1140,N_571,N_677);
or U1141 (N_1141,In_2849,N_74);
or U1142 (N_1142,In_742,N_57);
or U1143 (N_1143,N_399,In_2529);
xnor U1144 (N_1144,In_1486,In_786);
nor U1145 (N_1145,In_281,N_850);
xnor U1146 (N_1146,In_1260,In_1296);
and U1147 (N_1147,In_2487,N_818);
nand U1148 (N_1148,In_2345,In_396);
xor U1149 (N_1149,In_2664,N_384);
nand U1150 (N_1150,N_412,In_1468);
or U1151 (N_1151,In_1308,N_355);
xor U1152 (N_1152,N_380,N_368);
xnor U1153 (N_1153,In_1814,N_470);
nor U1154 (N_1154,In_1497,N_867);
nand U1155 (N_1155,N_672,In_563);
nor U1156 (N_1156,In_118,N_694);
nand U1157 (N_1157,In_2274,In_31);
xor U1158 (N_1158,In_194,N_647);
xnor U1159 (N_1159,In_2078,N_864);
or U1160 (N_1160,In_2,N_750);
or U1161 (N_1161,N_298,N_109);
nor U1162 (N_1162,In_2503,In_1853);
nor U1163 (N_1163,N_992,In_49);
xor U1164 (N_1164,In_91,N_406);
nor U1165 (N_1165,N_795,In_828);
or U1166 (N_1166,N_369,In_2134);
and U1167 (N_1167,N_305,N_884);
nor U1168 (N_1168,In_1846,In_360);
and U1169 (N_1169,N_344,N_787);
nor U1170 (N_1170,N_811,N_371);
xor U1171 (N_1171,N_686,In_913);
nand U1172 (N_1172,In_627,In_413);
nor U1173 (N_1173,In_2227,N_796);
and U1174 (N_1174,N_542,In_966);
and U1175 (N_1175,In_1977,In_1433);
or U1176 (N_1176,In_1022,N_455);
nand U1177 (N_1177,N_774,N_55);
xor U1178 (N_1178,N_215,N_387);
nand U1179 (N_1179,In_2180,In_1062);
nand U1180 (N_1180,N_237,N_351);
xnor U1181 (N_1181,N_967,N_615);
and U1182 (N_1182,N_165,N_235);
nand U1183 (N_1183,In_519,In_901);
nor U1184 (N_1184,N_518,In_1743);
nor U1185 (N_1185,N_28,In_2605);
nand U1186 (N_1186,In_1830,N_613);
nor U1187 (N_1187,N_360,N_324);
xor U1188 (N_1188,In_2569,In_520);
and U1189 (N_1189,N_20,N_725);
nand U1190 (N_1190,N_638,N_426);
or U1191 (N_1191,N_913,In_2418);
or U1192 (N_1192,N_190,N_907);
nand U1193 (N_1193,N_568,In_478);
nand U1194 (N_1194,In_481,In_2749);
or U1195 (N_1195,N_837,In_151);
or U1196 (N_1196,N_102,In_2110);
and U1197 (N_1197,In_1224,N_553);
and U1198 (N_1198,In_198,In_1951);
and U1199 (N_1199,In_1095,In_2063);
and U1200 (N_1200,N_193,N_714);
and U1201 (N_1201,N_508,N_567);
or U1202 (N_1202,N_256,In_2293);
nand U1203 (N_1203,In_430,N_692);
xnor U1204 (N_1204,In_1344,N_974);
or U1205 (N_1205,N_252,In_265);
nor U1206 (N_1206,In_2328,N_231);
nand U1207 (N_1207,N_505,N_290);
or U1208 (N_1208,In_1156,N_723);
xnor U1209 (N_1209,In_2713,N_893);
or U1210 (N_1210,In_2666,In_2463);
or U1211 (N_1211,N_328,N_683);
xor U1212 (N_1212,In_1574,N_94);
or U1213 (N_1213,In_163,In_688);
or U1214 (N_1214,N_268,In_1612);
xor U1215 (N_1215,In_166,In_964);
and U1216 (N_1216,N_765,N_283);
xor U1217 (N_1217,In_1154,In_2837);
xor U1218 (N_1218,In_351,In_254);
or U1219 (N_1219,N_575,In_2772);
and U1220 (N_1220,N_817,In_2019);
nand U1221 (N_1221,N_404,In_1440);
nand U1222 (N_1222,N_320,N_317);
nand U1223 (N_1223,In_2089,N_531);
and U1224 (N_1224,N_821,In_1368);
nor U1225 (N_1225,N_958,N_414);
and U1226 (N_1226,In_1304,N_507);
and U1227 (N_1227,N_641,N_225);
or U1228 (N_1228,In_375,N_18);
nor U1229 (N_1229,N_679,In_2367);
and U1230 (N_1230,N_286,N_46);
and U1231 (N_1231,In_53,N_285);
nor U1232 (N_1232,N_859,N_186);
and U1233 (N_1233,N_136,In_2225);
nand U1234 (N_1234,In_2058,In_2788);
nor U1235 (N_1235,N_595,In_1191);
and U1236 (N_1236,In_952,In_1438);
or U1237 (N_1237,In_2362,N_620);
or U1238 (N_1238,N_594,In_2492);
nor U1239 (N_1239,In_2856,N_955);
and U1240 (N_1240,In_2268,In_2329);
and U1241 (N_1241,N_366,N_125);
nand U1242 (N_1242,In_2583,In_1827);
xnor U1243 (N_1243,In_885,N_996);
nor U1244 (N_1244,N_216,N_739);
and U1245 (N_1245,N_562,N_100);
or U1246 (N_1246,N_75,In_2096);
or U1247 (N_1247,In_2747,In_1229);
nor U1248 (N_1248,N_336,N_468);
or U1249 (N_1249,N_975,In_2866);
or U1250 (N_1250,N_157,In_2085);
xnor U1251 (N_1251,N_411,In_261);
nor U1252 (N_1252,N_823,In_2748);
xnor U1253 (N_1253,In_2237,In_2648);
xor U1254 (N_1254,In_2054,In_1728);
and U1255 (N_1255,In_1176,N_314);
nor U1256 (N_1256,N_22,In_2049);
xor U1257 (N_1257,N_578,N_780);
nand U1258 (N_1258,In_1799,In_2164);
nor U1259 (N_1259,N_898,In_1579);
nand U1260 (N_1260,In_2334,In_200);
xor U1261 (N_1261,N_885,N_98);
or U1262 (N_1262,N_529,In_2791);
nor U1263 (N_1263,In_243,N_822);
or U1264 (N_1264,In_1103,N_653);
and U1265 (N_1265,In_1680,N_515);
and U1266 (N_1266,N_980,In_611);
nor U1267 (N_1267,In_3,N_142);
or U1268 (N_1268,In_2436,N_629);
xnor U1269 (N_1269,N_645,N_702);
nor U1270 (N_1270,N_236,In_2482);
nor U1271 (N_1271,In_219,In_2766);
or U1272 (N_1272,In_1060,N_425);
nor U1273 (N_1273,In_587,N_373);
xnor U1274 (N_1274,In_159,In_750);
xor U1275 (N_1275,In_355,In_1678);
nand U1276 (N_1276,N_152,In_1729);
or U1277 (N_1277,In_2292,N_855);
xor U1278 (N_1278,In_1258,In_2843);
nor U1279 (N_1279,In_94,N_886);
xnor U1280 (N_1280,N_931,In_2861);
and U1281 (N_1281,N_663,In_989);
and U1282 (N_1282,In_81,In_1766);
xor U1283 (N_1283,In_1936,N_941);
or U1284 (N_1284,N_416,N_97);
xor U1285 (N_1285,N_483,N_700);
nand U1286 (N_1286,N_630,N_26);
xor U1287 (N_1287,N_635,N_119);
xnor U1288 (N_1288,In_1543,In_955);
nor U1289 (N_1289,N_533,In_386);
nand U1290 (N_1290,In_34,N_306);
nand U1291 (N_1291,N_789,In_122);
nand U1292 (N_1292,N_430,N_989);
and U1293 (N_1293,In_1184,N_319);
nor U1294 (N_1294,N_107,N_271);
and U1295 (N_1295,In_887,N_246);
nand U1296 (N_1296,N_668,N_742);
and U1297 (N_1297,In_1195,N_372);
xnor U1298 (N_1298,N_450,N_64);
and U1299 (N_1299,In_2591,N_920);
or U1300 (N_1300,In_1432,N_741);
nor U1301 (N_1301,In_528,N_463);
nor U1302 (N_1302,N_697,N_340);
or U1303 (N_1303,N_935,In_2450);
or U1304 (N_1304,In_394,In_2691);
nor U1305 (N_1305,In_2223,In_47);
and U1306 (N_1306,N_987,N_878);
nand U1307 (N_1307,In_2199,N_948);
nand U1308 (N_1308,In_387,N_764);
nor U1309 (N_1309,In_1122,N_359);
and U1310 (N_1310,In_432,N_498);
and U1311 (N_1311,N_528,In_390);
and U1312 (N_1312,In_1456,N_421);
and U1313 (N_1313,In_1330,N_998);
or U1314 (N_1314,In_2850,In_1282);
nor U1315 (N_1315,N_217,In_602);
nand U1316 (N_1316,In_1477,In_1718);
and U1317 (N_1317,In_771,In_512);
nor U1318 (N_1318,In_2007,N_952);
and U1319 (N_1319,N_191,In_1014);
nand U1320 (N_1320,N_134,N_776);
xor U1321 (N_1321,In_554,N_813);
xor U1322 (N_1322,N_655,N_464);
xor U1323 (N_1323,N_144,N_173);
xnor U1324 (N_1324,N_962,N_79);
or U1325 (N_1325,In_2564,N_633);
nor U1326 (N_1326,In_1960,N_705);
nor U1327 (N_1327,N_433,In_2421);
xor U1328 (N_1328,N_99,In_1105);
or U1329 (N_1329,N_875,N_863);
or U1330 (N_1330,In_415,In_1927);
xnor U1331 (N_1331,N_902,N_218);
nand U1332 (N_1332,In_2394,In_2452);
nand U1333 (N_1333,In_1648,N_383);
and U1334 (N_1334,In_1595,In_556);
nor U1335 (N_1335,In_1162,N_249);
nor U1336 (N_1336,N_435,N_12);
nor U1337 (N_1337,In_1651,In_408);
nand U1338 (N_1338,N_345,N_131);
and U1339 (N_1339,N_799,N_66);
nand U1340 (N_1340,N_767,N_730);
nand U1341 (N_1341,N_36,N_365);
nand U1342 (N_1342,In_2417,In_1313);
nand U1343 (N_1343,In_1004,In_1415);
xor U1344 (N_1344,N_68,In_1932);
nor U1345 (N_1345,N_701,N_978);
and U1346 (N_1346,N_4,N_281);
nor U1347 (N_1347,N_652,N_745);
and U1348 (N_1348,N_634,N_133);
or U1349 (N_1349,In_1327,In_2790);
xnor U1350 (N_1350,In_2601,In_1923);
nand U1351 (N_1351,N_851,In_723);
nor U1352 (N_1352,In_64,In_2526);
or U1353 (N_1353,In_1943,In_1274);
xor U1354 (N_1354,In_2986,In_2238);
or U1355 (N_1355,N_370,In_264);
or U1356 (N_1356,In_1061,N_866);
and U1357 (N_1357,In_2612,In_483);
and U1358 (N_1358,In_813,N_514);
and U1359 (N_1359,N_649,N_824);
nor U1360 (N_1360,N_582,N_82);
and U1361 (N_1361,N_791,N_151);
xor U1362 (N_1362,In_905,In_1199);
xnor U1363 (N_1363,N_392,N_440);
nand U1364 (N_1364,In_150,N_105);
xor U1365 (N_1365,N_600,In_1423);
and U1366 (N_1366,N_788,N_673);
or U1367 (N_1367,N_260,In_2256);
and U1368 (N_1368,N_226,N_569);
or U1369 (N_1369,N_202,N_985);
nor U1370 (N_1370,N_660,In_2729);
and U1371 (N_1371,N_535,N_80);
nand U1372 (N_1372,N_756,N_954);
nor U1373 (N_1373,N_143,N_189);
nand U1374 (N_1374,In_272,N_311);
nand U1375 (N_1375,In_462,In_1284);
xor U1376 (N_1376,In_1880,N_735);
nor U1377 (N_1377,In_2798,In_1976);
nor U1378 (N_1378,In_392,In_2444);
nand U1379 (N_1379,N_607,In_2593);
and U1380 (N_1380,N_727,N_882);
and U1381 (N_1381,In_1458,N_713);
or U1382 (N_1382,In_1442,N_240);
nor U1383 (N_1383,N_681,In_1392);
nand U1384 (N_1384,N_536,N_388);
nand U1385 (N_1385,N_971,In_267);
nand U1386 (N_1386,In_178,N_40);
nor U1387 (N_1387,In_2745,N_112);
nand U1388 (N_1388,In_1279,In_859);
and U1389 (N_1389,In_610,N_228);
nand U1390 (N_1390,In_1904,In_972);
xnor U1391 (N_1391,N_409,N_988);
xnor U1392 (N_1392,In_2447,In_2546);
nor U1393 (N_1393,N_844,N_565);
or U1394 (N_1394,In_1254,In_2364);
nand U1395 (N_1395,In_1938,In_533);
nand U1396 (N_1396,N_106,In_1464);
nand U1397 (N_1397,In_1594,In_2208);
nand U1398 (N_1398,In_1452,N_917);
nand U1399 (N_1399,N_579,N_141);
nand U1400 (N_1400,N_691,In_501);
xor U1401 (N_1401,N_77,In_2336);
xor U1402 (N_1402,N_263,In_2799);
nand U1403 (N_1403,In_2108,In_284);
nand U1404 (N_1404,In_1,In_2443);
or U1405 (N_1405,In_314,N_720);
nand U1406 (N_1406,In_2670,N_826);
or U1407 (N_1407,In_1268,N_347);
xnor U1408 (N_1408,In_2999,In_2029);
xor U1409 (N_1409,N_454,N_890);
and U1410 (N_1410,In_1851,In_1685);
nand U1411 (N_1411,N_871,N_364);
or U1412 (N_1412,N_443,In_2787);
and U1413 (N_1413,In_1476,N_995);
and U1414 (N_1414,N_698,N_773);
nand U1415 (N_1415,In_817,N_339);
or U1416 (N_1416,In_239,In_2489);
or U1417 (N_1417,In_2212,N_417);
nor U1418 (N_1418,N_675,In_1840);
and U1419 (N_1419,In_774,N_447);
or U1420 (N_1420,In_2604,N_103);
and U1421 (N_1421,N_881,N_192);
xor U1422 (N_1422,N_220,N_976);
nand U1423 (N_1423,N_856,In_1947);
nand U1424 (N_1424,In_2230,In_1683);
nor U1425 (N_1425,In_329,In_939);
and U1426 (N_1426,N_517,N_277);
nand U1427 (N_1427,In_2584,N_257);
xor U1428 (N_1428,N_178,In_2501);
nand U1429 (N_1429,In_2018,In_1682);
or U1430 (N_1430,In_2568,N_790);
nor U1431 (N_1431,N_771,In_986);
and U1432 (N_1432,In_2757,In_1165);
nand U1433 (N_1433,In_2011,In_1854);
xor U1434 (N_1434,N_95,N_906);
nor U1435 (N_1435,In_521,N_156);
xnor U1436 (N_1436,In_1734,N_590);
xnor U1437 (N_1437,N_184,N_900);
or U1438 (N_1438,In_1706,In_965);
xnor U1439 (N_1439,In_190,In_893);
nor U1440 (N_1440,In_453,N_502);
and U1441 (N_1441,In_1804,In_1378);
nor U1442 (N_1442,In_844,N_671);
nor U1443 (N_1443,N_135,N_737);
and U1444 (N_1444,In_2422,N_853);
or U1445 (N_1445,N_876,N_284);
nand U1446 (N_1446,N_31,In_70);
nand U1447 (N_1447,N_379,N_836);
and U1448 (N_1448,N_904,N_646);
nor U1449 (N_1449,In_684,In_1385);
xnor U1450 (N_1450,In_1939,N_557);
and U1451 (N_1451,In_1785,In_218);
nor U1452 (N_1452,In_2984,In_827);
xnor U1453 (N_1453,In_1752,N_539);
or U1454 (N_1454,In_101,N_684);
nand U1455 (N_1455,In_1689,In_1178);
nor U1456 (N_1456,In_1166,In_1613);
nand U1457 (N_1457,In_2226,In_1564);
nor U1458 (N_1458,N_56,In_2401);
and U1459 (N_1459,N_924,In_1029);
nor U1460 (N_1460,In_1578,N_753);
nor U1461 (N_1461,In_810,N_182);
nor U1462 (N_1462,In_2415,N_944);
nand U1463 (N_1463,N_690,N_456);
xnor U1464 (N_1464,In_1896,In_1217);
and U1465 (N_1465,In_1358,In_917);
nand U1466 (N_1466,N_779,N_722);
nor U1467 (N_1467,In_1437,In_2960);
nand U1468 (N_1468,In_1334,In_2150);
or U1469 (N_1469,In_2627,In_2080);
or U1470 (N_1470,N_744,In_1478);
or U1471 (N_1471,In_1619,N_748);
nor U1472 (N_1472,In_2959,N_86);
xnor U1473 (N_1473,In_1359,N_147);
nor U1474 (N_1474,In_860,In_2114);
nand U1475 (N_1475,N_956,N_279);
or U1476 (N_1476,N_50,N_174);
nand U1477 (N_1477,N_251,In_511);
and U1478 (N_1478,N_888,In_502);
and U1479 (N_1479,In_2365,In_1770);
nand U1480 (N_1480,In_229,In_1907);
nor U1481 (N_1481,N_23,N_928);
nor U1482 (N_1482,In_793,N_937);
and U1483 (N_1483,In_2976,N_362);
nor U1484 (N_1484,N_245,N_983);
and U1485 (N_1485,N_797,N_145);
xor U1486 (N_1486,N_487,In_469);
xor U1487 (N_1487,N_234,In_2168);
or U1488 (N_1488,N_90,In_969);
or U1489 (N_1489,N_259,In_2228);
or U1490 (N_1490,N_466,N_625);
or U1491 (N_1491,In_1649,In_1007);
xor U1492 (N_1492,In_296,In_2734);
or U1493 (N_1493,N_763,N_670);
nor U1494 (N_1494,In_460,In_2549);
and U1495 (N_1495,N_968,N_585);
nand U1496 (N_1496,In_48,In_1585);
or U1497 (N_1497,In_2409,N_584);
or U1498 (N_1498,N_933,In_2910);
or U1499 (N_1499,N_208,N_67);
and U1500 (N_1500,N_695,In_75);
nor U1501 (N_1501,In_45,N_990);
and U1502 (N_1502,N_378,In_1872);
and U1503 (N_1503,In_2660,In_1986);
nor U1504 (N_1504,In_1086,N_402);
nor U1505 (N_1505,N_596,In_1883);
or U1506 (N_1506,In_2107,In_1252);
and U1507 (N_1507,In_2727,In_1117);
nor U1508 (N_1508,N_785,N_155);
or U1509 (N_1509,In_2887,N_162);
or U1510 (N_1510,In_1996,N_749);
and U1511 (N_1511,In_111,N_310);
or U1512 (N_1512,N_462,In_1890);
nor U1513 (N_1513,In_1206,In_736);
nand U1514 (N_1514,In_1349,In_878);
and U1515 (N_1515,In_1697,In_1818);
xnor U1516 (N_1516,N_966,In_1891);
and U1517 (N_1517,In_1338,In_1791);
nand U1518 (N_1518,In_2679,N_495);
xor U1519 (N_1519,In_975,N_951);
nand U1520 (N_1520,N_139,In_1155);
nand U1521 (N_1521,In_540,N_834);
nand U1522 (N_1522,In_2390,In_1130);
nor U1523 (N_1523,In_2122,N_848);
xor U1524 (N_1524,In_2363,N_598);
nor U1525 (N_1525,N_42,In_1128);
and U1526 (N_1526,N_448,N_474);
and U1527 (N_1527,N_92,N_83);
xnor U1528 (N_1528,In_1513,In_2868);
nor U1529 (N_1529,In_230,N_432);
xor U1530 (N_1530,In_217,N_566);
xor U1531 (N_1531,N_504,In_1116);
xor U1532 (N_1532,N_639,In_136);
nor U1533 (N_1533,N_408,In_892);
nand U1534 (N_1534,N_762,N_183);
nor U1535 (N_1535,N_558,N_798);
and U1536 (N_1536,In_16,In_2896);
nand U1537 (N_1537,N_807,N_676);
and U1538 (N_1538,In_1514,In_1503);
nand U1539 (N_1539,N_117,N_942);
nand U1540 (N_1540,N_719,In_1527);
nor U1541 (N_1541,N_576,N_581);
nor U1542 (N_1542,In_2635,In_1240);
and U1543 (N_1543,N_643,N_815);
or U1544 (N_1544,In_338,In_1777);
nor U1545 (N_1545,In_2880,In_2603);
and U1546 (N_1546,In_472,In_1148);
nand U1547 (N_1547,N_709,N_831);
and U1548 (N_1548,N_478,N_297);
and U1549 (N_1549,In_1397,N_740);
and U1550 (N_1550,In_1404,N_282);
or U1551 (N_1551,In_1544,N_96);
or U1552 (N_1552,N_540,N_800);
nand U1553 (N_1553,N_858,N_843);
or U1554 (N_1554,In_2560,N_925);
xnor U1555 (N_1555,In_2351,In_1396);
nand U1556 (N_1556,N_446,In_1724);
xor U1557 (N_1557,N_729,In_618);
xnor U1558 (N_1558,N_910,In_1488);
or U1559 (N_1559,N_13,In_183);
or U1560 (N_1560,In_2081,In_1518);
or U1561 (N_1561,In_1034,In_626);
nand U1562 (N_1562,In_2298,N_743);
nor U1563 (N_1563,In_95,In_2217);
or U1564 (N_1564,In_562,In_1710);
nand U1565 (N_1565,In_2610,In_30);
nand U1566 (N_1566,In_2253,N_919);
nand U1567 (N_1567,N_960,N_621);
xnor U1568 (N_1568,N_213,In_246);
or U1569 (N_1569,N_905,In_1265);
xor U1570 (N_1570,In_2726,N_258);
nand U1571 (N_1571,N_445,In_400);
nor U1572 (N_1572,N_35,N_8);
nand U1573 (N_1573,N_214,N_179);
xnor U1574 (N_1574,N_573,N_318);
or U1575 (N_1575,In_903,In_1408);
nand U1576 (N_1576,N_903,N_322);
and U1577 (N_1577,In_2718,N_793);
and U1578 (N_1578,In_2735,In_1889);
nand U1579 (N_1579,In_1744,N_238);
xor U1580 (N_1580,N_945,In_2451);
nand U1581 (N_1581,In_109,In_2842);
nor U1582 (N_1582,N_833,N_330);
xnor U1583 (N_1583,N_726,N_419);
xor U1584 (N_1584,In_2347,N_593);
nand U1585 (N_1585,N_877,In_1266);
xor U1586 (N_1586,In_2448,In_2475);
nand U1587 (N_1587,In_1802,In_2185);
or U1588 (N_1588,In_1644,In_2094);
xor U1589 (N_1589,N_63,In_1860);
or U1590 (N_1590,N_21,In_385);
xor U1591 (N_1591,N_398,In_1286);
or U1592 (N_1592,N_667,N_62);
or U1593 (N_1593,In_1580,In_1137);
xnor U1594 (N_1594,N_239,In_908);
and U1595 (N_1595,In_1512,In_1158);
or U1596 (N_1596,In_1988,N_376);
and U1597 (N_1597,N_497,In_1698);
and U1598 (N_1598,In_918,In_1764);
nor U1599 (N_1599,N_674,N_469);
nor U1600 (N_1600,N_32,N_403);
nand U1601 (N_1601,In_52,N_759);
nor U1602 (N_1602,In_1732,In_1771);
and U1603 (N_1603,In_513,N_17);
and U1604 (N_1604,In_1063,N_108);
nand U1605 (N_1605,N_476,N_87);
xor U1606 (N_1606,In_2127,In_2458);
and U1607 (N_1607,N_10,N_631);
nand U1608 (N_1608,N_939,In_2694);
and U1609 (N_1609,In_2481,N_522);
and U1610 (N_1610,In_15,In_1688);
and U1611 (N_1611,N_911,N_733);
nand U1612 (N_1612,In_1675,N_543);
nand U1613 (N_1613,N_555,N_312);
xor U1614 (N_1614,In_753,In_991);
nor U1615 (N_1615,N_716,In_1741);
and U1616 (N_1616,N_52,N_879);
and U1617 (N_1617,In_2017,In_492);
xnor U1618 (N_1618,N_589,N_973);
or U1619 (N_1619,In_978,N_943);
or U1620 (N_1620,In_336,In_2361);
xor U1621 (N_1621,N_242,N_657);
xor U1622 (N_1622,In_2302,In_367);
nand U1623 (N_1623,N_623,N_265);
and U1624 (N_1624,In_1058,In_2232);
nor U1625 (N_1625,In_1068,N_321);
or U1626 (N_1626,In_419,N_626);
or U1627 (N_1627,In_393,In_2958);
or U1628 (N_1628,N_846,N_274);
nor U1629 (N_1629,In_2867,In_2121);
xnor U1630 (N_1630,In_735,In_1726);
xnor U1631 (N_1631,N_970,N_611);
nand U1632 (N_1632,In_364,In_1672);
nor U1633 (N_1633,In_647,N_333);
xor U1634 (N_1634,N_936,N_129);
and U1635 (N_1635,N_946,N_48);
nor U1636 (N_1636,N_511,N_751);
xor U1637 (N_1637,N_270,In_588);
xor U1638 (N_1638,N_304,N_199);
nand U1639 (N_1639,In_2690,In_2163);
or U1640 (N_1640,In_1275,N_991);
and U1641 (N_1641,N_809,N_490);
xor U1642 (N_1642,In_2118,N_880);
nand U1643 (N_1643,N_947,N_37);
and U1644 (N_1644,In_2207,In_1961);
nand U1645 (N_1645,N_453,In_757);
nor U1646 (N_1646,In_1964,In_208);
and U1647 (N_1647,N_449,In_814);
or U1648 (N_1648,In_293,N_69);
xor U1649 (N_1649,In_1092,In_2903);
or U1650 (N_1650,In_2159,N_899);
xor U1651 (N_1651,In_2630,In_2881);
xor U1652 (N_1652,N_397,In_1293);
nand U1653 (N_1653,In_287,In_732);
nor U1654 (N_1654,In_2400,N_825);
or U1655 (N_1655,N_176,In_295);
or U1656 (N_1656,In_2663,In_577);
xor U1657 (N_1657,N_114,In_1213);
nand U1658 (N_1658,In_1287,N_981);
nand U1659 (N_1659,N_835,N_221);
xor U1660 (N_1660,In_115,In_1354);
nor U1661 (N_1661,N_754,N_964);
or U1662 (N_1662,N_127,In_187);
xor U1663 (N_1663,N_560,In_1485);
and U1664 (N_1664,N_521,N_159);
or U1665 (N_1665,N_175,N_601);
nor U1666 (N_1666,N_438,In_1878);
nor U1667 (N_1667,N_572,In_1336);
and U1668 (N_1668,N_841,In_1997);
xnor U1669 (N_1669,In_96,N_757);
xnor U1670 (N_1670,N_34,N_891);
nor U1671 (N_1671,In_642,In_291);
xnor U1672 (N_1672,N_603,N_342);
xnor U1673 (N_1673,In_2267,N_428);
xnor U1674 (N_1674,In_2068,In_406);
and U1675 (N_1675,N_972,In_2099);
nand U1676 (N_1676,In_2700,In_93);
xor U1677 (N_1677,N_458,In_2093);
or U1678 (N_1678,N_491,In_1762);
nand U1679 (N_1679,In_2519,In_2297);
nor U1680 (N_1680,N_343,In_1525);
and U1681 (N_1681,In_2240,N_209);
and U1682 (N_1682,In_1797,N_358);
nand U1683 (N_1683,In_1072,N_354);
and U1684 (N_1684,In_2275,N_43);
and U1685 (N_1685,N_637,In_2371);
xnor U1686 (N_1686,In_617,N_482);
nor U1687 (N_1687,In_1078,N_953);
nand U1688 (N_1688,In_673,N_300);
and U1689 (N_1689,N_132,N_422);
xnor U1690 (N_1690,N_832,In_2197);
nor U1691 (N_1691,N_781,N_164);
nor U1692 (N_1692,N_76,In_2352);
nor U1693 (N_1693,In_1283,N_101);
xor U1694 (N_1694,N_587,N_327);
nor U1695 (N_1695,In_2736,In_451);
and U1696 (N_1696,N_393,N_682);
nor U1697 (N_1697,N_166,N_618);
xor U1698 (N_1698,N_546,N_804);
nor U1699 (N_1699,In_2571,N_471);
and U1700 (N_1700,N_396,In_176);
xor U1701 (N_1701,In_2312,N_524);
nand U1702 (N_1702,N_61,In_2946);
nor U1703 (N_1703,N_545,In_235);
nand U1704 (N_1704,N_738,N_194);
or U1705 (N_1705,N_325,In_2339);
or U1706 (N_1706,N_707,N_280);
xnor U1707 (N_1707,In_332,N_85);
nand U1708 (N_1708,In_1568,In_158);
xor U1709 (N_1709,N_200,In_866);
nand U1710 (N_1710,In_2323,N_512);
nand U1711 (N_1711,In_608,In_1628);
nor U1712 (N_1712,In_2015,In_2548);
nand U1713 (N_1713,N_513,In_110);
or U1714 (N_1714,N_746,In_914);
xnor U1715 (N_1715,In_837,N_401);
or U1716 (N_1716,N_91,In_409);
nand U1717 (N_1717,In_539,In_1917);
xor U1718 (N_1718,In_1800,In_1446);
xor U1719 (N_1719,In_2889,N_784);
nand U1720 (N_1720,In_2533,In_2314);
and U1721 (N_1721,N_503,N_849);
xnor U1722 (N_1722,In_1469,In_2758);
nand U1723 (N_1723,In_1347,In_2877);
or U1724 (N_1724,N_439,In_1816);
xor U1725 (N_1725,In_1526,N_662);
nor U1726 (N_1726,In_123,In_1186);
or U1727 (N_1727,In_1235,In_1318);
nor U1728 (N_1728,In_2618,N_496);
or U1729 (N_1729,In_1835,In_1163);
or U1730 (N_1730,In_2774,In_1881);
nand U1731 (N_1731,In_1482,In_504);
nand U1732 (N_1732,In_311,N_551);
or U1733 (N_1733,N_908,N_346);
or U1734 (N_1734,N_814,N_872);
and U1735 (N_1735,In_2382,In_36);
nor U1736 (N_1736,N_860,In_85);
nor U1737 (N_1737,N_45,N_6);
or U1738 (N_1738,N_544,N_806);
nand U1739 (N_1739,In_2449,N_999);
nand U1740 (N_1740,In_553,N_704);
nor U1741 (N_1741,In_1305,N_303);
nor U1742 (N_1742,N_617,N_308);
nand U1743 (N_1743,In_353,In_1416);
or U1744 (N_1744,N_323,N_44);
nor U1745 (N_1745,N_889,In_316);
or U1746 (N_1746,In_559,N_950);
or U1747 (N_1747,In_746,N_177);
nand U1748 (N_1748,In_84,In_308);
or U1749 (N_1749,In_202,In_1490);
xnor U1750 (N_1750,In_1311,In_655);
nand U1751 (N_1751,In_33,In_2191);
nand U1752 (N_1752,N_624,N_222);
xnor U1753 (N_1753,N_326,N_348);
or U1754 (N_1754,N_204,N_196);
nor U1755 (N_1755,N_580,In_2634);
and U1756 (N_1756,In_2599,In_2218);
and U1757 (N_1757,N_616,In_948);
or U1758 (N_1758,In_388,In_2926);
and U1759 (N_1759,N_391,N_661);
nand U1760 (N_1760,N_230,In_152);
nor U1761 (N_1761,N_669,In_2882);
nand U1762 (N_1762,N_752,N_229);
xor U1763 (N_1763,In_1419,N_986);
and U1764 (N_1764,In_654,In_1920);
and U1765 (N_1765,N_72,In_949);
xor U1766 (N_1766,In_2405,N_153);
or U1767 (N_1767,N_731,N_198);
or U1768 (N_1768,N_632,N_187);
xnor U1769 (N_1769,N_640,In_1237);
xnor U1770 (N_1770,N_805,In_2677);
xnor U1771 (N_1771,N_315,In_401);
nand U1772 (N_1772,N_169,N_390);
xor U1773 (N_1773,In_2888,N_732);
or U1774 (N_1774,N_708,N_693);
and U1775 (N_1775,N_27,N_949);
or U1776 (N_1776,N_65,In_2906);
nor U1777 (N_1777,N_605,In_2002);
and U1778 (N_1778,N_577,In_855);
nor U1779 (N_1779,In_1000,N_158);
nor U1780 (N_1780,N_896,N_777);
nand U1781 (N_1781,In_1884,In_838);
and U1782 (N_1782,In_2251,N_356);
xor U1783 (N_1783,N_609,N_847);
nor U1784 (N_1784,In_1256,In_1089);
xor U1785 (N_1785,N_916,In_1074);
or U1786 (N_1786,In_1627,N_11);
and U1787 (N_1787,In_769,In_1010);
and U1788 (N_1788,N_816,In_1278);
or U1789 (N_1789,N_38,In_2457);
nor U1790 (N_1790,In_2629,N_769);
nand U1791 (N_1791,In_2538,In_2370);
xnor U1792 (N_1792,In_1134,In_1573);
or U1793 (N_1793,N_586,N_766);
nor U1794 (N_1794,In_2306,N_718);
xnor U1795 (N_1795,In_718,N_53);
nor U1796 (N_1796,N_437,In_2466);
or U1797 (N_1797,In_1747,In_2504);
nand U1798 (N_1798,In_1703,In_1250);
xor U1799 (N_1799,In_1504,N_772);
and U1800 (N_1800,In_826,N_648);
and U1801 (N_1801,In_2053,N_247);
or U1802 (N_1802,N_519,In_438);
nor U1803 (N_1803,N_113,N_869);
xnor U1804 (N_1804,N_54,In_1202);
and U1805 (N_1805,N_93,N_537);
nand U1806 (N_1806,N_622,In_2071);
or U1807 (N_1807,In_1188,In_1348);
xnor U1808 (N_1808,N_185,In_2137);
nand U1809 (N_1809,In_931,N_137);
and U1810 (N_1810,In_1727,In_213);
or U1811 (N_1811,N_301,In_506);
nor U1812 (N_1812,N_534,N_352);
nand U1813 (N_1813,In_2759,N_614);
or U1814 (N_1814,N_316,In_312);
or U1815 (N_1815,In_638,N_865);
or U1816 (N_1816,N_294,In_2865);
nand U1817 (N_1817,N_33,In_2957);
xnor U1818 (N_1818,N_123,In_1066);
or U1819 (N_1819,N_287,In_1399);
nor U1820 (N_1820,N_427,N_839);
nand U1821 (N_1821,In_214,In_2407);
and U1822 (N_1822,N_211,N_89);
nand U1823 (N_1823,N_459,N_712);
nand U1824 (N_1824,N_570,In_2822);
nand U1825 (N_1825,In_1212,N_485);
xor U1826 (N_1826,N_84,In_2574);
nand U1827 (N_1827,N_16,In_776);
or U1828 (N_1828,In_1289,N_335);
nor U1829 (N_1829,In_1767,In_1193);
and U1830 (N_1830,N_493,N_262);
xor U1831 (N_1831,N_997,N_678);
nor U1832 (N_1832,In_1537,In_2321);
or U1833 (N_1833,In_1429,In_1434);
nand U1834 (N_1834,In_2720,In_1635);
nand U1835 (N_1835,In_442,N_167);
and U1836 (N_1836,In_697,N_163);
xnor U1837 (N_1837,In_2023,In_1326);
nor U1838 (N_1838,N_710,N_386);
nand U1839 (N_1839,In_1855,In_1561);
and U1840 (N_1840,N_768,N_168);
and U1841 (N_1841,N_874,In_1998);
or U1842 (N_1842,In_92,In_1159);
or U1843 (N_1843,In_2214,N_334);
or U1844 (N_1844,N_689,N_472);
xor U1845 (N_1845,In_1065,N_253);
and U1846 (N_1846,In_373,In_578);
nor U1847 (N_1847,N_219,In_1211);
nor U1848 (N_1848,N_538,N_415);
and U1849 (N_1849,In_345,N_205);
nand U1850 (N_1850,N_721,N_808);
xnor U1851 (N_1851,In_1665,In_2258);
nand U1852 (N_1852,N_49,In_1769);
or U1853 (N_1853,In_232,N_223);
and U1854 (N_1854,In_185,N_206);
xor U1855 (N_1855,N_628,N_845);
nor U1856 (N_1856,N_254,N_552);
or U1857 (N_1857,In_4,N_715);
nor U1858 (N_1858,N_736,N_549);
and U1859 (N_1859,N_827,In_138);
and U1860 (N_1860,In_891,N_484);
or U1861 (N_1861,In_2961,In_1622);
nand U1862 (N_1862,N_81,In_537);
xnor U1863 (N_1863,N_591,N_926);
nand U1864 (N_1864,In_1530,N_299);
or U1865 (N_1865,N_278,In_139);
xnor U1866 (N_1866,N_802,N_541);
nor U1867 (N_1867,In_1059,In_6);
nor U1868 (N_1868,N_210,In_637);
nor U1869 (N_1869,N_747,In_2152);
nand U1870 (N_1870,N_530,N_606);
nor U1871 (N_1871,In_1653,N_329);
and U1872 (N_1872,N_927,N_842);
or U1873 (N_1873,In_2341,In_1801);
or U1874 (N_1874,N_232,N_706);
or U1875 (N_1875,N_656,In_184);
nand U1876 (N_1876,N_550,In_1281);
nor U1877 (N_1877,In_1720,N_477);
and U1878 (N_1878,N_140,In_1135);
nand U1879 (N_1879,N_39,N_685);
xor U1880 (N_1880,N_861,N_181);
or U1881 (N_1881,N_126,N_687);
or U1882 (N_1882,N_267,N_499);
and U1883 (N_1883,In_1807,N_241);
nand U1884 (N_1884,N_527,N_2);
nor U1885 (N_1885,N_574,N_840);
nor U1886 (N_1886,In_1586,In_982);
or U1887 (N_1887,In_1466,In_1945);
nand U1888 (N_1888,N_892,N_361);
xnor U1889 (N_1889,N_0,N_604);
and U1890 (N_1890,In_489,N_812);
nor U1891 (N_1891,N_820,In_2428);
xor U1892 (N_1892,N_444,In_1894);
nor U1893 (N_1893,N_41,In_1592);
nand U1894 (N_1894,In_536,N_255);
or U1895 (N_1895,In_1712,N_130);
and U1896 (N_1896,N_659,N_699);
xor U1897 (N_1897,In_2951,In_1975);
and U1898 (N_1898,In_2821,In_2032);
xnor U1899 (N_1899,In_2665,N_149);
nand U1900 (N_1900,In_1239,N_982);
and U1901 (N_1901,In_2044,N_15);
xor U1902 (N_1902,In_907,N_993);
nand U1903 (N_1903,In_1795,In_1455);
xnor U1904 (N_1904,In_276,N_115);
nor U1905 (N_1905,In_2084,In_2219);
and U1906 (N_1906,In_1597,In_1247);
or U1907 (N_1907,N_501,In_714);
and U1908 (N_1908,N_332,N_775);
nand U1909 (N_1909,In_1590,N_418);
nor U1910 (N_1910,N_688,N_47);
xor U1911 (N_1911,N_994,N_696);
xnor U1912 (N_1912,In_2194,N_276);
nor U1913 (N_1913,In_670,In_2525);
or U1914 (N_1914,N_510,N_5);
nand U1915 (N_1915,N_680,N_377);
nand U1916 (N_1916,N_363,N_489);
and U1917 (N_1917,In_2918,N_961);
xor U1918 (N_1918,N_154,N_957);
or U1919 (N_1919,N_9,N_338);
nor U1920 (N_1920,N_429,In_428);
and U1921 (N_1921,N_894,In_993);
and U1922 (N_1922,N_122,N_932);
nor U1923 (N_1923,In_530,In_2973);
or U1924 (N_1924,N_473,In_2944);
or U1925 (N_1925,In_605,In_231);
nand U1926 (N_1926,N_110,N_120);
nand U1927 (N_1927,In_1765,In_156);
or U1928 (N_1928,In_2074,N_547);
and U1929 (N_1929,In_2061,N_88);
and U1930 (N_1930,In_2845,N_460);
xor U1931 (N_1931,N_201,In_681);
xor U1932 (N_1932,In_130,N_778);
nor U1933 (N_1933,N_161,In_2662);
nor U1934 (N_1934,N_58,In_2072);
nand U1935 (N_1935,N_929,N_494);
nand U1936 (N_1936,In_722,N_786);
or U1937 (N_1937,N_405,In_594);
xnor U1938 (N_1938,N_394,N_375);
xor U1939 (N_1939,In_137,N_78);
or U1940 (N_1940,N_269,In_1740);
or U1941 (N_1941,In_2731,N_758);
or U1942 (N_1942,N_959,In_2678);
and U1943 (N_1943,In_1214,In_1614);
and U1944 (N_1944,N_930,N_868);
nor U1945 (N_1945,In_72,In_1716);
nor U1946 (N_1946,N_965,In_1968);
nor U1947 (N_1947,N_828,In_2042);
xnor U1948 (N_1948,N_854,N_486);
and U1949 (N_1949,N_465,In_1032);
xnor U1950 (N_1950,In_2125,N_400);
or U1951 (N_1951,In_634,In_2898);
xnor U1952 (N_1952,N_350,In_1160);
nand U1953 (N_1953,N_532,In_2190);
xnor U1954 (N_1954,N_1,N_60);
nand U1955 (N_1955,N_51,N_3);
nand U1956 (N_1956,N_104,In_1001);
and U1957 (N_1957,N_857,N_148);
xor U1958 (N_1958,In_2578,N_30);
xnor U1959 (N_1959,N_651,In_1445);
nor U1960 (N_1960,In_1529,N_599);
nor U1961 (N_1961,N_288,N_451);
xnor U1962 (N_1962,In_257,N_829);
nor U1963 (N_1963,N_488,In_449);
xnor U1964 (N_1964,In_1659,N_520);
nor U1965 (N_1965,N_203,N_261);
nor U1966 (N_1966,In_2707,In_207);
nand U1967 (N_1967,N_293,N_264);
nand U1968 (N_1968,N_665,In_1129);
xnor U1969 (N_1969,In_2967,N_273);
and U1970 (N_1970,In_1895,N_770);
nor U1971 (N_1971,In_2814,In_1864);
nor U1972 (N_1972,In_2349,N_588);
nand U1973 (N_1973,In_1981,N_14);
or U1974 (N_1974,In_2656,In_2330);
nand U1975 (N_1975,N_500,In_1958);
xor U1976 (N_1976,N_272,In_968);
nand U1977 (N_1977,In_2393,In_1248);
and U1978 (N_1978,In_1829,N_979);
and U1979 (N_1979,N_389,N_357);
and U1980 (N_1980,In_493,In_2055);
or U1981 (N_1981,In_1617,N_381);
nor U1982 (N_1982,N_654,N_664);
or U1983 (N_1983,In_865,N_382);
nor U1984 (N_1984,N_608,In_2128);
xor U1985 (N_1985,N_711,In_1285);
nand U1986 (N_1986,In_1859,In_1821);
and U1987 (N_1987,In_1994,N_116);
nor U1988 (N_1988,In_310,In_1828);
xor U1989 (N_1989,In_2979,N_407);
nand U1990 (N_1990,In_1115,In_1929);
xnor U1991 (N_1991,In_1792,In_82);
or U1992 (N_1992,In_558,N_895);
nor U1993 (N_1993,N_724,N_224);
xnor U1994 (N_1994,In_2453,N_233);
or U1995 (N_1995,N_921,N_915);
and U1996 (N_1996,N_548,N_810);
nor U1997 (N_1997,N_479,In_1731);
xnor U1998 (N_1998,In_1870,In_2052);
nand U1999 (N_1999,In_2904,In_1109);
and U2000 (N_2000,N_1824,N_1063);
or U2001 (N_2001,N_1087,N_1724);
nor U2002 (N_2002,N_1456,N_1714);
xnor U2003 (N_2003,N_1025,N_1305);
or U2004 (N_2004,N_1872,N_1678);
nor U2005 (N_2005,N_1591,N_1895);
and U2006 (N_2006,N_1083,N_1985);
nor U2007 (N_2007,N_1309,N_1925);
nor U2008 (N_2008,N_1915,N_1019);
nand U2009 (N_2009,N_1358,N_1751);
and U2010 (N_2010,N_1891,N_1006);
nand U2011 (N_2011,N_1240,N_1426);
and U2012 (N_2012,N_1058,N_1784);
nand U2013 (N_2013,N_1541,N_1204);
nand U2014 (N_2014,N_1877,N_1203);
nand U2015 (N_2015,N_1804,N_1145);
xor U2016 (N_2016,N_1210,N_1148);
xnor U2017 (N_2017,N_1213,N_1002);
and U2018 (N_2018,N_1064,N_1887);
or U2019 (N_2019,N_1505,N_1435);
nand U2020 (N_2020,N_1289,N_1209);
and U2021 (N_2021,N_1038,N_1229);
and U2022 (N_2022,N_1233,N_1132);
xor U2023 (N_2023,N_1375,N_1901);
or U2024 (N_2024,N_1406,N_1809);
nor U2025 (N_2025,N_1223,N_1042);
xor U2026 (N_2026,N_1394,N_1979);
xnor U2027 (N_2027,N_1323,N_1857);
or U2028 (N_2028,N_1244,N_1712);
nor U2029 (N_2029,N_1753,N_1247);
or U2030 (N_2030,N_1995,N_1922);
xor U2031 (N_2031,N_1629,N_1957);
nand U2032 (N_2032,N_1546,N_1988);
nand U2033 (N_2033,N_1154,N_1592);
or U2034 (N_2034,N_1054,N_1074);
and U2035 (N_2035,N_1357,N_1573);
xnor U2036 (N_2036,N_1873,N_1626);
nor U2037 (N_2037,N_1243,N_1445);
nor U2038 (N_2038,N_1760,N_1013);
and U2039 (N_2039,N_1806,N_1161);
and U2040 (N_2040,N_1056,N_1226);
nor U2041 (N_2041,N_1869,N_1306);
nand U2042 (N_2042,N_1106,N_1333);
nor U2043 (N_2043,N_1321,N_1687);
xnor U2044 (N_2044,N_1397,N_1099);
and U2045 (N_2045,N_1946,N_1920);
nor U2046 (N_2046,N_1744,N_1594);
nand U2047 (N_2047,N_1218,N_1414);
and U2048 (N_2048,N_1647,N_1973);
nor U2049 (N_2049,N_1436,N_1624);
or U2050 (N_2050,N_1476,N_1950);
xnor U2051 (N_2051,N_1715,N_1679);
and U2052 (N_2052,N_1519,N_1819);
and U2053 (N_2053,N_1699,N_1033);
xor U2054 (N_2054,N_1686,N_1384);
nand U2055 (N_2055,N_1266,N_1562);
nor U2056 (N_2056,N_1978,N_1864);
xnor U2057 (N_2057,N_1200,N_1853);
nand U2058 (N_2058,N_1368,N_1367);
nor U2059 (N_2059,N_1708,N_1379);
and U2060 (N_2060,N_1234,N_1997);
or U2061 (N_2061,N_1743,N_1871);
nor U2062 (N_2062,N_1623,N_1655);
and U2063 (N_2063,N_1398,N_1783);
xor U2064 (N_2064,N_1693,N_1727);
nor U2065 (N_2065,N_1944,N_1747);
xnor U2066 (N_2066,N_1604,N_1775);
or U2067 (N_2067,N_1156,N_1822);
nand U2068 (N_2068,N_1577,N_1916);
nor U2069 (N_2069,N_1508,N_1481);
xor U2070 (N_2070,N_1068,N_1958);
and U2071 (N_2071,N_1552,N_1459);
xor U2072 (N_2072,N_1888,N_1188);
nor U2073 (N_2073,N_1745,N_1917);
xnor U2074 (N_2074,N_1475,N_1769);
nand U2075 (N_2075,N_1494,N_1834);
xnor U2076 (N_2076,N_1967,N_1771);
and U2077 (N_2077,N_1963,N_1945);
xor U2078 (N_2078,N_1974,N_1764);
nand U2079 (N_2079,N_1041,N_1903);
xnor U2080 (N_2080,N_1217,N_1731);
nor U2081 (N_2081,N_1503,N_1345);
nand U2082 (N_2082,N_1838,N_1007);
nand U2083 (N_2083,N_1080,N_1166);
nand U2084 (N_2084,N_1449,N_1291);
nor U2085 (N_2085,N_1430,N_1109);
xnor U2086 (N_2086,N_1516,N_1717);
and U2087 (N_2087,N_1488,N_1320);
or U2088 (N_2088,N_1721,N_1311);
or U2089 (N_2089,N_1876,N_1110);
xor U2090 (N_2090,N_1580,N_1868);
nor U2091 (N_2091,N_1421,N_1124);
or U2092 (N_2092,N_1607,N_1990);
nand U2093 (N_2093,N_1105,N_1462);
and U2094 (N_2094,N_1847,N_1911);
and U2095 (N_2095,N_1589,N_1900);
or U2096 (N_2096,N_1179,N_1350);
nor U2097 (N_2097,N_1694,N_1596);
or U2098 (N_2098,N_1278,N_1150);
nand U2099 (N_2099,N_1371,N_1103);
or U2100 (N_2100,N_1720,N_1242);
and U2101 (N_2101,N_1057,N_1996);
nand U2102 (N_2102,N_1411,N_1125);
or U2103 (N_2103,N_1199,N_1685);
and U2104 (N_2104,N_1960,N_1395);
nand U2105 (N_2105,N_1661,N_1961);
and U2106 (N_2106,N_1196,N_1897);
nor U2107 (N_2107,N_1858,N_1739);
or U2108 (N_2108,N_1840,N_1539);
and U2109 (N_2109,N_1113,N_1910);
or U2110 (N_2110,N_1581,N_1785);
or U2111 (N_2111,N_1374,N_1540);
nor U2112 (N_2112,N_1646,N_1018);
and U2113 (N_2113,N_1250,N_1151);
xnor U2114 (N_2114,N_1370,N_1016);
nor U2115 (N_2115,N_1265,N_1768);
nor U2116 (N_2116,N_1931,N_1558);
xnor U2117 (N_2117,N_1641,N_1537);
xnor U2118 (N_2118,N_1183,N_1741);
xor U2119 (N_2119,N_1220,N_1290);
or U2120 (N_2120,N_1376,N_1932);
xnor U2121 (N_2121,N_1228,N_1927);
and U2122 (N_2122,N_1332,N_1193);
and U2123 (N_2123,N_1094,N_1640);
nand U2124 (N_2124,N_1660,N_1093);
or U2125 (N_2125,N_1839,N_1951);
or U2126 (N_2126,N_1575,N_1889);
or U2127 (N_2127,N_1788,N_1606);
nor U2128 (N_2128,N_1984,N_1898);
nor U2129 (N_2129,N_1442,N_1307);
and U2130 (N_2130,N_1935,N_1458);
and U2131 (N_2131,N_1420,N_1830);
and U2132 (N_2132,N_1014,N_1297);
or U2133 (N_2133,N_1500,N_1551);
nor U2134 (N_2134,N_1582,N_1667);
nor U2135 (N_2135,N_1177,N_1614);
and U2136 (N_2136,N_1635,N_1765);
or U2137 (N_2137,N_1652,N_1020);
and U2138 (N_2138,N_1649,N_1850);
xnor U2139 (N_2139,N_1115,N_1104);
and U2140 (N_2140,N_1799,N_1100);
or U2141 (N_2141,N_1918,N_1909);
and U2142 (N_2142,N_1538,N_1464);
and U2143 (N_2143,N_1584,N_1631);
and U2144 (N_2144,N_1095,N_1554);
or U2145 (N_2145,N_1122,N_1031);
nand U2146 (N_2146,N_1969,N_1189);
nor U2147 (N_2147,N_1480,N_1583);
nand U2148 (N_2148,N_1369,N_1719);
and U2149 (N_2149,N_1410,N_1489);
nand U2150 (N_2150,N_1610,N_1860);
nand U2151 (N_2151,N_1102,N_1465);
or U2152 (N_2152,N_1875,N_1593);
xor U2153 (N_2153,N_1281,N_1272);
and U2154 (N_2154,N_1848,N_1062);
and U2155 (N_2155,N_1986,N_1256);
nand U2156 (N_2156,N_1786,N_1515);
nand U2157 (N_2157,N_1224,N_1170);
nand U2158 (N_2158,N_1146,N_1101);
or U2159 (N_2159,N_1619,N_1416);
nand U2160 (N_2160,N_1601,N_1557);
or U2161 (N_2161,N_1767,N_1409);
xnor U2162 (N_2162,N_1510,N_1735);
nor U2163 (N_2163,N_1319,N_1841);
nand U2164 (N_2164,N_1096,N_1527);
and U2165 (N_2165,N_1971,N_1938);
xnor U2166 (N_2166,N_1257,N_1947);
nand U2167 (N_2167,N_1863,N_1136);
nor U2168 (N_2168,N_1908,N_1737);
nand U2169 (N_2169,N_1001,N_1865);
or U2170 (N_2170,N_1457,N_1705);
xnor U2171 (N_2171,N_1674,N_1617);
nor U2172 (N_2172,N_1362,N_1015);
or U2173 (N_2173,N_1817,N_1733);
and U2174 (N_2174,N_1259,N_1455);
xor U2175 (N_2175,N_1241,N_1249);
xor U2176 (N_2176,N_1879,N_1003);
nor U2177 (N_2177,N_1366,N_1301);
or U2178 (N_2178,N_1736,N_1279);
or U2179 (N_2179,N_1588,N_1325);
nor U2180 (N_2180,N_1698,N_1866);
xor U2181 (N_2181,N_1828,N_1123);
xor U2182 (N_2182,N_1522,N_1861);
nor U2183 (N_2183,N_1611,N_1381);
nand U2184 (N_2184,N_1454,N_1388);
nand U2185 (N_2185,N_1514,N_1022);
and U2186 (N_2186,N_1692,N_1178);
xor U2187 (N_2187,N_1341,N_1966);
and U2188 (N_2188,N_1129,N_1077);
nand U2189 (N_2189,N_1339,N_1949);
and U2190 (N_2190,N_1066,N_1560);
or U2191 (N_2191,N_1502,N_1885);
nor U2192 (N_2192,N_1587,N_1498);
nand U2193 (N_2193,N_1772,N_1586);
xnor U2194 (N_2194,N_1347,N_1902);
xor U2195 (N_2195,N_1135,N_1843);
nand U2196 (N_2196,N_1825,N_1884);
nand U2197 (N_2197,N_1127,N_1399);
xnor U2198 (N_2198,N_1725,N_1466);
or U2199 (N_2199,N_1304,N_1616);
and U2200 (N_2200,N_1326,N_1793);
nand U2201 (N_2201,N_1282,N_1982);
nor U2202 (N_2202,N_1331,N_1401);
nor U2203 (N_2203,N_1665,N_1214);
xnor U2204 (N_2204,N_1238,N_1327);
nor U2205 (N_2205,N_1520,N_1254);
xnor U2206 (N_2206,N_1026,N_1980);
or U2207 (N_2207,N_1479,N_1798);
and U2208 (N_2208,N_1695,N_1742);
nand U2209 (N_2209,N_1750,N_1924);
and U2210 (N_2210,N_1048,N_1658);
nand U2211 (N_2211,N_1595,N_1886);
or U2212 (N_2212,N_1726,N_1470);
nor U2213 (N_2213,N_1564,N_1269);
or U2214 (N_2214,N_1656,N_1477);
nor U2215 (N_2215,N_1632,N_1934);
and U2216 (N_2216,N_1512,N_1338);
xnor U2217 (N_2217,N_1299,N_1779);
and U2218 (N_2218,N_1359,N_1088);
and U2219 (N_2219,N_1422,N_1770);
nand U2220 (N_2220,N_1024,N_1073);
nor U2221 (N_2221,N_1992,N_1298);
and U2222 (N_2222,N_1182,N_1471);
xor U2223 (N_2223,N_1496,N_1752);
or U2224 (N_2224,N_1408,N_1482);
nand U2225 (N_2225,N_1757,N_1849);
nor U2226 (N_2226,N_1287,N_1448);
nor U2227 (N_2227,N_1120,N_1152);
nor U2228 (N_2228,N_1981,N_1232);
nand U2229 (N_2229,N_1314,N_1930);
and U2230 (N_2230,N_1463,N_1748);
or U2231 (N_2231,N_1075,N_1942);
and U2232 (N_2232,N_1827,N_1386);
or U2233 (N_2233,N_1570,N_1746);
nand U2234 (N_2234,N_1975,N_1324);
or U2235 (N_2235,N_1427,N_1663);
nor U2236 (N_2236,N_1452,N_1469);
or U2237 (N_2237,N_1219,N_1813);
nor U2238 (N_2238,N_1681,N_1008);
nor U2239 (N_2239,N_1567,N_1991);
nand U2240 (N_2240,N_1518,N_1501);
and U2241 (N_2241,N_1168,N_1603);
nand U2242 (N_2242,N_1155,N_1923);
and U2243 (N_2243,N_1759,N_1716);
or U2244 (N_2244,N_1881,N_1084);
nor U2245 (N_2245,N_1285,N_1977);
nor U2246 (N_2246,N_1485,N_1789);
or U2247 (N_2247,N_1385,N_1237);
and U2248 (N_2248,N_1423,N_1833);
nor U2249 (N_2249,N_1139,N_1212);
and U2250 (N_2250,N_1638,N_1998);
nand U2251 (N_2251,N_1643,N_1569);
nand U2252 (N_2252,N_1650,N_1763);
nand U2253 (N_2253,N_1352,N_1811);
and U2254 (N_2254,N_1533,N_1700);
or U2255 (N_2255,N_1602,N_1317);
xnor U2256 (N_2256,N_1186,N_1164);
and U2257 (N_2257,N_1055,N_1308);
and U2258 (N_2258,N_1052,N_1492);
nor U2259 (N_2259,N_1734,N_1360);
nand U2260 (N_2260,N_1364,N_1790);
and U2261 (N_2261,N_1563,N_1252);
nand U2262 (N_2262,N_1524,N_1070);
or U2263 (N_2263,N_1432,N_1845);
or U2264 (N_2264,N_1114,N_1896);
or U2265 (N_2265,N_1880,N_1085);
and U2266 (N_2266,N_1372,N_1954);
or U2267 (N_2267,N_1439,N_1437);
xor U2268 (N_2268,N_1815,N_1221);
nor U2269 (N_2269,N_1078,N_1277);
nand U2270 (N_2270,N_1802,N_1535);
xor U2271 (N_2271,N_1836,N_1941);
and U2272 (N_2272,N_1044,N_1964);
xor U2273 (N_2273,N_1417,N_1574);
nand U2274 (N_2274,N_1526,N_1709);
or U2275 (N_2275,N_1728,N_1275);
and U2276 (N_2276,N_1994,N_1517);
or U2277 (N_2277,N_1939,N_1671);
and U2278 (N_2278,N_1701,N_1749);
nor U2279 (N_2279,N_1639,N_1870);
or U2280 (N_2280,N_1071,N_1141);
and U2281 (N_2281,N_1316,N_1905);
nor U2282 (N_2282,N_1149,N_1195);
nand U2283 (N_2283,N_1176,N_1559);
nand U2284 (N_2284,N_1491,N_1628);
nand U2285 (N_2285,N_1117,N_1069);
nand U2286 (N_2286,N_1255,N_1805);
nor U2287 (N_2287,N_1555,N_1621);
xor U2288 (N_2288,N_1703,N_1835);
and U2289 (N_2289,N_1782,N_1144);
or U2290 (N_2290,N_1111,N_1549);
and U2291 (N_2291,N_1904,N_1260);
xor U2292 (N_2292,N_1523,N_1756);
nand U2293 (N_2293,N_1021,N_1672);
and U2294 (N_2294,N_1618,N_1206);
xor U2295 (N_2295,N_1017,N_1344);
nor U2296 (N_2296,N_1952,N_1197);
nand U2297 (N_2297,N_1597,N_1133);
xor U2298 (N_2298,N_1882,N_1812);
or U2299 (N_2299,N_1722,N_1440);
nor U2300 (N_2300,N_1590,N_1174);
and U2301 (N_2301,N_1191,N_1528);
and U2302 (N_2302,N_1413,N_1668);
and U2303 (N_2303,N_1867,N_1061);
or U2304 (N_2304,N_1545,N_1684);
or U2305 (N_2305,N_1808,N_1585);
nor U2306 (N_2306,N_1959,N_1509);
and U2307 (N_2307,N_1976,N_1444);
or U2308 (N_2308,N_1207,N_1600);
and U2309 (N_2309,N_1292,N_1576);
or U2310 (N_2310,N_1983,N_1273);
and U2311 (N_2311,N_1940,N_1403);
and U2312 (N_2312,N_1683,N_1023);
and U2313 (N_2313,N_1286,N_1625);
and U2314 (N_2314,N_1513,N_1263);
xor U2315 (N_2315,N_1246,N_1929);
nand U2316 (N_2316,N_1473,N_1082);
nor U2317 (N_2317,N_1697,N_1215);
and U2318 (N_2318,N_1499,N_1377);
nor U2319 (N_2319,N_1556,N_1140);
nor U2320 (N_2320,N_1310,N_1968);
xor U2321 (N_2321,N_1653,N_1644);
nand U2322 (N_2322,N_1211,N_1318);
nand U2323 (N_2323,N_1107,N_1004);
or U2324 (N_2324,N_1495,N_1356);
xnor U2325 (N_2325,N_1418,N_1598);
or U2326 (N_2326,N_1919,N_1890);
nand U2327 (N_2327,N_1451,N_1236);
nand U2328 (N_2328,N_1300,N_1689);
xnor U2329 (N_2329,N_1936,N_1572);
nor U2330 (N_2330,N_1157,N_1067);
nand U2331 (N_2331,N_1258,N_1438);
and U2332 (N_2332,N_1852,N_1086);
nor U2333 (N_2333,N_1312,N_1295);
nand U2334 (N_2334,N_1354,N_1810);
and U2335 (N_2335,N_1682,N_1363);
nand U2336 (N_2336,N_1676,N_1005);
or U2337 (N_2337,N_1637,N_1270);
or U2338 (N_2338,N_1059,N_1134);
or U2339 (N_2339,N_1544,N_1032);
xor U2340 (N_2340,N_1820,N_1566);
nand U2341 (N_2341,N_1844,N_1034);
and U2342 (N_2342,N_1548,N_1579);
and U2343 (N_2343,N_1424,N_1778);
xnor U2344 (N_2344,N_1956,N_1187);
nor U2345 (N_2345,N_1680,N_1267);
xnor U2346 (N_2346,N_1664,N_1340);
and U2347 (N_2347,N_1429,N_1393);
nand U2348 (N_2348,N_1758,N_1669);
xor U2349 (N_2349,N_1239,N_1128);
or U2350 (N_2350,N_1832,N_1511);
nand U2351 (N_2351,N_1821,N_1740);
xnor U2352 (N_2352,N_1999,N_1704);
nand U2353 (N_2353,N_1874,N_1642);
or U2354 (N_2354,N_1543,N_1035);
xor U2355 (N_2355,N_1153,N_1713);
and U2356 (N_2356,N_1796,N_1171);
xnor U2357 (N_2357,N_1612,N_1613);
nand U2358 (N_2358,N_1634,N_1690);
xnor U2359 (N_2359,N_1284,N_1081);
nand U2360 (N_2360,N_1776,N_1400);
or U2361 (N_2361,N_1965,N_1529);
nand U2362 (N_2362,N_1230,N_1172);
or U2363 (N_2363,N_1280,N_1303);
xor U2364 (N_2364,N_1412,N_1264);
and U2365 (N_2365,N_1336,N_1036);
nor U2366 (N_2366,N_1231,N_1090);
xnor U2367 (N_2367,N_1670,N_1355);
nor U2368 (N_2368,N_1648,N_1803);
and U2369 (N_2369,N_1268,N_1862);
nor U2370 (N_2370,N_1142,N_1792);
or U2371 (N_2371,N_1504,N_1245);
nand U2372 (N_2372,N_1723,N_1953);
nand U2373 (N_2373,N_1181,N_1677);
nor U2374 (N_2374,N_1807,N_1630);
or U2375 (N_2375,N_1313,N_1912);
or U2376 (N_2376,N_1027,N_1185);
and U2377 (N_2377,N_1766,N_1497);
or U2378 (N_2378,N_1012,N_1121);
or U2379 (N_2379,N_1274,N_1029);
or U2380 (N_2380,N_1787,N_1390);
or U2381 (N_2381,N_1774,N_1262);
xnor U2382 (N_2382,N_1460,N_1894);
xor U2383 (N_2383,N_1175,N_1955);
nor U2384 (N_2384,N_1706,N_1937);
and U2385 (N_2385,N_1192,N_1119);
or U2386 (N_2386,N_1060,N_1732);
nor U2387 (N_2387,N_1826,N_1553);
nand U2388 (N_2388,N_1165,N_1651);
xnor U2389 (N_2389,N_1450,N_1392);
or U2390 (N_2390,N_1948,N_1261);
and U2391 (N_2391,N_1797,N_1800);
nand U2392 (N_2392,N_1180,N_1046);
xor U2393 (N_2393,N_1160,N_1899);
xor U2394 (N_2394,N_1906,N_1823);
nor U2395 (N_2395,N_1296,N_1216);
xnor U2396 (N_2396,N_1561,N_1235);
or U2397 (N_2397,N_1521,N_1028);
xnor U2398 (N_2398,N_1198,N_1816);
and U2399 (N_2399,N_1348,N_1353);
nor U2400 (N_2400,N_1137,N_1383);
and U2401 (N_2401,N_1831,N_1645);
nand U2402 (N_2402,N_1130,N_1780);
nor U2403 (N_2403,N_1428,N_1098);
nand U2404 (N_2404,N_1707,N_1461);
xnor U2405 (N_2405,N_1138,N_1615);
and U2406 (N_2406,N_1387,N_1525);
and U2407 (N_2407,N_1892,N_1402);
nor U2408 (N_2408,N_1051,N_1037);
xor U2409 (N_2409,N_1484,N_1688);
and U2410 (N_2410,N_1691,N_1933);
or U2411 (N_2411,N_1755,N_1380);
or U2412 (N_2412,N_1378,N_1483);
nor U2413 (N_2413,N_1419,N_1914);
nand U2414 (N_2414,N_1346,N_1711);
nor U2415 (N_2415,N_1550,N_1710);
or U2416 (N_2416,N_1926,N_1116);
xor U2417 (N_2417,N_1335,N_1097);
nor U2418 (N_2418,N_1294,N_1222);
nand U2419 (N_2419,N_1846,N_1276);
nor U2420 (N_2420,N_1030,N_1328);
nand U2421 (N_2421,N_1578,N_1190);
xnor U2422 (N_2422,N_1859,N_1283);
nor U2423 (N_2423,N_1000,N_1605);
nand U2424 (N_2424,N_1043,N_1791);
or U2425 (N_2425,N_1486,N_1507);
and U2426 (N_2426,N_1162,N_1472);
xnor U2427 (N_2427,N_1131,N_1091);
nand U2428 (N_2428,N_1565,N_1718);
xnor U2429 (N_2429,N_1158,N_1329);
xor U2430 (N_2430,N_1928,N_1194);
xor U2431 (N_2431,N_1972,N_1490);
xnor U2432 (N_2432,N_1659,N_1225);
nor U2433 (N_2433,N_1208,N_1673);
or U2434 (N_2434,N_1349,N_1441);
nor U2435 (N_2435,N_1762,N_1163);
nor U2436 (N_2436,N_1468,N_1474);
or U2437 (N_2437,N_1322,N_1993);
and U2438 (N_2438,N_1010,N_1391);
or U2439 (N_2439,N_1729,N_1143);
xor U2440 (N_2440,N_1829,N_1696);
or U2441 (N_2441,N_1365,N_1147);
xnor U2442 (N_2442,N_1907,N_1531);
xor U2443 (N_2443,N_1337,N_1467);
xnor U2444 (N_2444,N_1842,N_1065);
and U2445 (N_2445,N_1666,N_1089);
or U2446 (N_2446,N_1184,N_1288);
nor U2447 (N_2447,N_1506,N_1011);
nand U2448 (N_2448,N_1443,N_1657);
xnor U2449 (N_2449,N_1205,N_1404);
xor U2450 (N_2450,N_1989,N_1818);
and U2451 (N_2451,N_1407,N_1253);
xor U2452 (N_2452,N_1053,N_1636);
or U2453 (N_2453,N_1795,N_1092);
nor U2454 (N_2454,N_1434,N_1921);
xnor U2455 (N_2455,N_1547,N_1302);
and U2456 (N_2456,N_1571,N_1351);
or U2457 (N_2457,N_1389,N_1801);
xnor U2458 (N_2458,N_1987,N_1794);
nand U2459 (N_2459,N_1781,N_1330);
and U2460 (N_2460,N_1493,N_1530);
nand U2461 (N_2461,N_1662,N_1405);
and U2462 (N_2462,N_1738,N_1970);
or U2463 (N_2463,N_1446,N_1761);
and U2464 (N_2464,N_1893,N_1854);
and U2465 (N_2465,N_1169,N_1167);
and U2466 (N_2466,N_1730,N_1248);
nand U2467 (N_2467,N_1754,N_1542);
or U2468 (N_2468,N_1855,N_1201);
xnor U2469 (N_2469,N_1415,N_1361);
nor U2470 (N_2470,N_1396,N_1943);
and U2471 (N_2471,N_1315,N_1009);
and U2472 (N_2472,N_1039,N_1159);
nor U2473 (N_2473,N_1599,N_1654);
nor U2474 (N_2474,N_1568,N_1342);
xnor U2475 (N_2475,N_1433,N_1536);
nor U2476 (N_2476,N_1702,N_1108);
nand U2477 (N_2477,N_1532,N_1072);
nand U2478 (N_2478,N_1622,N_1373);
nand U2479 (N_2479,N_1487,N_1447);
nor U2480 (N_2480,N_1620,N_1126);
or U2481 (N_2481,N_1777,N_1112);
or U2482 (N_2482,N_1050,N_1773);
and U2483 (N_2483,N_1251,N_1627);
nand U2484 (N_2484,N_1675,N_1040);
and U2485 (N_2485,N_1079,N_1878);
and U2486 (N_2486,N_1814,N_1227);
nor U2487 (N_2487,N_1382,N_1856);
and U2488 (N_2488,N_1608,N_1293);
nor U2489 (N_2489,N_1913,N_1271);
xor U2490 (N_2490,N_1425,N_1343);
or U2491 (N_2491,N_1609,N_1049);
nor U2492 (N_2492,N_1851,N_1045);
nor U2493 (N_2493,N_1118,N_1478);
nor U2494 (N_2494,N_1173,N_1334);
or U2495 (N_2495,N_1202,N_1047);
nand U2496 (N_2496,N_1431,N_1076);
or U2497 (N_2497,N_1883,N_1534);
nand U2498 (N_2498,N_1837,N_1633);
xnor U2499 (N_2499,N_1962,N_1453);
or U2500 (N_2500,N_1730,N_1999);
xor U2501 (N_2501,N_1467,N_1008);
xnor U2502 (N_2502,N_1078,N_1297);
nor U2503 (N_2503,N_1775,N_1136);
xor U2504 (N_2504,N_1977,N_1353);
nand U2505 (N_2505,N_1864,N_1777);
and U2506 (N_2506,N_1942,N_1859);
and U2507 (N_2507,N_1826,N_1608);
and U2508 (N_2508,N_1186,N_1257);
nor U2509 (N_2509,N_1899,N_1388);
and U2510 (N_2510,N_1498,N_1364);
nor U2511 (N_2511,N_1318,N_1417);
nand U2512 (N_2512,N_1054,N_1991);
nor U2513 (N_2513,N_1975,N_1346);
and U2514 (N_2514,N_1847,N_1752);
and U2515 (N_2515,N_1434,N_1801);
nor U2516 (N_2516,N_1713,N_1181);
xnor U2517 (N_2517,N_1015,N_1803);
nor U2518 (N_2518,N_1361,N_1903);
or U2519 (N_2519,N_1573,N_1274);
or U2520 (N_2520,N_1859,N_1513);
nor U2521 (N_2521,N_1975,N_1693);
xor U2522 (N_2522,N_1452,N_1111);
or U2523 (N_2523,N_1295,N_1949);
xnor U2524 (N_2524,N_1614,N_1602);
and U2525 (N_2525,N_1337,N_1507);
xor U2526 (N_2526,N_1009,N_1876);
xor U2527 (N_2527,N_1213,N_1572);
nand U2528 (N_2528,N_1785,N_1941);
nor U2529 (N_2529,N_1140,N_1496);
or U2530 (N_2530,N_1395,N_1603);
nor U2531 (N_2531,N_1647,N_1318);
nand U2532 (N_2532,N_1368,N_1949);
nor U2533 (N_2533,N_1282,N_1752);
and U2534 (N_2534,N_1387,N_1497);
nor U2535 (N_2535,N_1145,N_1187);
xor U2536 (N_2536,N_1846,N_1750);
and U2537 (N_2537,N_1905,N_1948);
nand U2538 (N_2538,N_1931,N_1473);
or U2539 (N_2539,N_1680,N_1498);
and U2540 (N_2540,N_1619,N_1926);
and U2541 (N_2541,N_1903,N_1024);
nor U2542 (N_2542,N_1684,N_1732);
or U2543 (N_2543,N_1033,N_1602);
or U2544 (N_2544,N_1239,N_1092);
or U2545 (N_2545,N_1868,N_1118);
xnor U2546 (N_2546,N_1494,N_1370);
nand U2547 (N_2547,N_1401,N_1497);
or U2548 (N_2548,N_1380,N_1611);
or U2549 (N_2549,N_1678,N_1314);
xor U2550 (N_2550,N_1952,N_1127);
and U2551 (N_2551,N_1497,N_1838);
nand U2552 (N_2552,N_1951,N_1108);
nor U2553 (N_2553,N_1710,N_1110);
or U2554 (N_2554,N_1298,N_1973);
xnor U2555 (N_2555,N_1894,N_1194);
nor U2556 (N_2556,N_1462,N_1925);
and U2557 (N_2557,N_1452,N_1342);
nor U2558 (N_2558,N_1970,N_1329);
nor U2559 (N_2559,N_1192,N_1026);
nor U2560 (N_2560,N_1430,N_1564);
and U2561 (N_2561,N_1150,N_1540);
xnor U2562 (N_2562,N_1593,N_1026);
xor U2563 (N_2563,N_1285,N_1184);
or U2564 (N_2564,N_1086,N_1036);
nand U2565 (N_2565,N_1833,N_1377);
or U2566 (N_2566,N_1895,N_1645);
or U2567 (N_2567,N_1314,N_1578);
nand U2568 (N_2568,N_1090,N_1265);
nand U2569 (N_2569,N_1189,N_1147);
xor U2570 (N_2570,N_1919,N_1089);
and U2571 (N_2571,N_1703,N_1377);
and U2572 (N_2572,N_1952,N_1986);
nand U2573 (N_2573,N_1335,N_1410);
or U2574 (N_2574,N_1965,N_1593);
and U2575 (N_2575,N_1013,N_1748);
nand U2576 (N_2576,N_1871,N_1012);
nor U2577 (N_2577,N_1069,N_1245);
or U2578 (N_2578,N_1047,N_1468);
xnor U2579 (N_2579,N_1505,N_1432);
or U2580 (N_2580,N_1884,N_1752);
and U2581 (N_2581,N_1363,N_1704);
xnor U2582 (N_2582,N_1117,N_1701);
and U2583 (N_2583,N_1503,N_1673);
and U2584 (N_2584,N_1697,N_1289);
or U2585 (N_2585,N_1115,N_1264);
xor U2586 (N_2586,N_1503,N_1620);
nand U2587 (N_2587,N_1100,N_1164);
and U2588 (N_2588,N_1982,N_1618);
and U2589 (N_2589,N_1688,N_1597);
or U2590 (N_2590,N_1605,N_1058);
nor U2591 (N_2591,N_1704,N_1769);
or U2592 (N_2592,N_1241,N_1188);
and U2593 (N_2593,N_1555,N_1176);
nor U2594 (N_2594,N_1899,N_1066);
xor U2595 (N_2595,N_1900,N_1220);
nor U2596 (N_2596,N_1985,N_1327);
xnor U2597 (N_2597,N_1351,N_1812);
or U2598 (N_2598,N_1083,N_1281);
nand U2599 (N_2599,N_1484,N_1047);
nor U2600 (N_2600,N_1106,N_1280);
xor U2601 (N_2601,N_1473,N_1209);
nand U2602 (N_2602,N_1600,N_1670);
and U2603 (N_2603,N_1601,N_1672);
and U2604 (N_2604,N_1385,N_1535);
and U2605 (N_2605,N_1157,N_1889);
or U2606 (N_2606,N_1120,N_1555);
and U2607 (N_2607,N_1453,N_1242);
xnor U2608 (N_2608,N_1091,N_1614);
xnor U2609 (N_2609,N_1901,N_1780);
or U2610 (N_2610,N_1991,N_1117);
nor U2611 (N_2611,N_1684,N_1222);
nor U2612 (N_2612,N_1314,N_1544);
or U2613 (N_2613,N_1862,N_1911);
and U2614 (N_2614,N_1334,N_1468);
nor U2615 (N_2615,N_1960,N_1693);
nand U2616 (N_2616,N_1840,N_1745);
and U2617 (N_2617,N_1817,N_1216);
and U2618 (N_2618,N_1037,N_1206);
and U2619 (N_2619,N_1615,N_1791);
and U2620 (N_2620,N_1246,N_1958);
or U2621 (N_2621,N_1912,N_1495);
nand U2622 (N_2622,N_1355,N_1724);
xor U2623 (N_2623,N_1118,N_1205);
or U2624 (N_2624,N_1359,N_1616);
nor U2625 (N_2625,N_1611,N_1835);
nor U2626 (N_2626,N_1065,N_1538);
or U2627 (N_2627,N_1164,N_1389);
nor U2628 (N_2628,N_1732,N_1262);
or U2629 (N_2629,N_1745,N_1018);
or U2630 (N_2630,N_1570,N_1194);
and U2631 (N_2631,N_1093,N_1952);
or U2632 (N_2632,N_1674,N_1347);
nand U2633 (N_2633,N_1461,N_1489);
nor U2634 (N_2634,N_1125,N_1888);
nand U2635 (N_2635,N_1733,N_1913);
xor U2636 (N_2636,N_1894,N_1917);
or U2637 (N_2637,N_1859,N_1565);
and U2638 (N_2638,N_1083,N_1284);
and U2639 (N_2639,N_1543,N_1484);
and U2640 (N_2640,N_1818,N_1218);
and U2641 (N_2641,N_1168,N_1187);
xor U2642 (N_2642,N_1624,N_1892);
or U2643 (N_2643,N_1872,N_1186);
and U2644 (N_2644,N_1629,N_1911);
nand U2645 (N_2645,N_1428,N_1220);
or U2646 (N_2646,N_1749,N_1090);
or U2647 (N_2647,N_1444,N_1264);
or U2648 (N_2648,N_1933,N_1120);
nand U2649 (N_2649,N_1335,N_1415);
and U2650 (N_2650,N_1250,N_1621);
xnor U2651 (N_2651,N_1140,N_1715);
xor U2652 (N_2652,N_1287,N_1951);
xnor U2653 (N_2653,N_1980,N_1462);
and U2654 (N_2654,N_1657,N_1710);
or U2655 (N_2655,N_1330,N_1211);
and U2656 (N_2656,N_1657,N_1681);
or U2657 (N_2657,N_1549,N_1317);
and U2658 (N_2658,N_1808,N_1742);
nand U2659 (N_2659,N_1583,N_1671);
nand U2660 (N_2660,N_1227,N_1872);
and U2661 (N_2661,N_1156,N_1579);
xnor U2662 (N_2662,N_1920,N_1688);
nor U2663 (N_2663,N_1563,N_1870);
nand U2664 (N_2664,N_1873,N_1368);
nor U2665 (N_2665,N_1798,N_1799);
xnor U2666 (N_2666,N_1652,N_1389);
or U2667 (N_2667,N_1183,N_1557);
nor U2668 (N_2668,N_1537,N_1794);
nor U2669 (N_2669,N_1891,N_1893);
and U2670 (N_2670,N_1224,N_1341);
or U2671 (N_2671,N_1621,N_1084);
nand U2672 (N_2672,N_1193,N_1362);
or U2673 (N_2673,N_1347,N_1146);
and U2674 (N_2674,N_1398,N_1163);
and U2675 (N_2675,N_1269,N_1186);
or U2676 (N_2676,N_1942,N_1760);
or U2677 (N_2677,N_1662,N_1169);
xnor U2678 (N_2678,N_1914,N_1358);
nor U2679 (N_2679,N_1373,N_1236);
nand U2680 (N_2680,N_1673,N_1315);
nand U2681 (N_2681,N_1744,N_1803);
or U2682 (N_2682,N_1390,N_1152);
or U2683 (N_2683,N_1951,N_1976);
or U2684 (N_2684,N_1418,N_1855);
and U2685 (N_2685,N_1995,N_1883);
or U2686 (N_2686,N_1111,N_1252);
nor U2687 (N_2687,N_1634,N_1227);
and U2688 (N_2688,N_1238,N_1860);
or U2689 (N_2689,N_1220,N_1746);
or U2690 (N_2690,N_1326,N_1842);
and U2691 (N_2691,N_1617,N_1031);
xnor U2692 (N_2692,N_1534,N_1647);
or U2693 (N_2693,N_1844,N_1671);
nor U2694 (N_2694,N_1218,N_1430);
nor U2695 (N_2695,N_1103,N_1189);
and U2696 (N_2696,N_1057,N_1574);
xor U2697 (N_2697,N_1008,N_1691);
or U2698 (N_2698,N_1563,N_1231);
xnor U2699 (N_2699,N_1323,N_1150);
nor U2700 (N_2700,N_1973,N_1948);
nor U2701 (N_2701,N_1782,N_1722);
nor U2702 (N_2702,N_1961,N_1666);
xor U2703 (N_2703,N_1236,N_1568);
nor U2704 (N_2704,N_1974,N_1116);
nand U2705 (N_2705,N_1048,N_1483);
nand U2706 (N_2706,N_1942,N_1560);
xor U2707 (N_2707,N_1786,N_1133);
nor U2708 (N_2708,N_1274,N_1259);
xor U2709 (N_2709,N_1339,N_1965);
or U2710 (N_2710,N_1893,N_1515);
xnor U2711 (N_2711,N_1297,N_1695);
nand U2712 (N_2712,N_1509,N_1539);
and U2713 (N_2713,N_1789,N_1638);
xor U2714 (N_2714,N_1799,N_1807);
xnor U2715 (N_2715,N_1862,N_1356);
nor U2716 (N_2716,N_1245,N_1261);
and U2717 (N_2717,N_1946,N_1217);
or U2718 (N_2718,N_1595,N_1836);
xor U2719 (N_2719,N_1906,N_1957);
or U2720 (N_2720,N_1046,N_1059);
nand U2721 (N_2721,N_1669,N_1460);
or U2722 (N_2722,N_1740,N_1509);
and U2723 (N_2723,N_1332,N_1050);
or U2724 (N_2724,N_1006,N_1353);
or U2725 (N_2725,N_1261,N_1167);
and U2726 (N_2726,N_1565,N_1583);
or U2727 (N_2727,N_1121,N_1406);
xnor U2728 (N_2728,N_1938,N_1091);
xnor U2729 (N_2729,N_1643,N_1069);
and U2730 (N_2730,N_1125,N_1645);
or U2731 (N_2731,N_1315,N_1713);
nand U2732 (N_2732,N_1082,N_1526);
xor U2733 (N_2733,N_1812,N_1982);
nor U2734 (N_2734,N_1379,N_1321);
nand U2735 (N_2735,N_1417,N_1581);
and U2736 (N_2736,N_1905,N_1427);
or U2737 (N_2737,N_1669,N_1071);
and U2738 (N_2738,N_1115,N_1540);
nor U2739 (N_2739,N_1048,N_1300);
xnor U2740 (N_2740,N_1273,N_1477);
or U2741 (N_2741,N_1073,N_1857);
and U2742 (N_2742,N_1631,N_1202);
and U2743 (N_2743,N_1542,N_1890);
nor U2744 (N_2744,N_1000,N_1715);
nor U2745 (N_2745,N_1933,N_1938);
nand U2746 (N_2746,N_1809,N_1629);
xor U2747 (N_2747,N_1731,N_1123);
and U2748 (N_2748,N_1221,N_1547);
or U2749 (N_2749,N_1783,N_1507);
nor U2750 (N_2750,N_1694,N_1774);
and U2751 (N_2751,N_1824,N_1167);
nor U2752 (N_2752,N_1006,N_1914);
xnor U2753 (N_2753,N_1321,N_1701);
nand U2754 (N_2754,N_1688,N_1835);
nand U2755 (N_2755,N_1088,N_1660);
nand U2756 (N_2756,N_1047,N_1994);
and U2757 (N_2757,N_1335,N_1739);
nor U2758 (N_2758,N_1402,N_1983);
nor U2759 (N_2759,N_1413,N_1096);
or U2760 (N_2760,N_1499,N_1623);
and U2761 (N_2761,N_1064,N_1167);
nor U2762 (N_2762,N_1791,N_1308);
and U2763 (N_2763,N_1127,N_1185);
nand U2764 (N_2764,N_1412,N_1092);
nand U2765 (N_2765,N_1066,N_1303);
nor U2766 (N_2766,N_1058,N_1505);
or U2767 (N_2767,N_1828,N_1270);
or U2768 (N_2768,N_1867,N_1291);
xnor U2769 (N_2769,N_1225,N_1456);
xnor U2770 (N_2770,N_1654,N_1615);
or U2771 (N_2771,N_1139,N_1296);
nand U2772 (N_2772,N_1323,N_1948);
nor U2773 (N_2773,N_1939,N_1995);
nand U2774 (N_2774,N_1740,N_1910);
xor U2775 (N_2775,N_1077,N_1966);
and U2776 (N_2776,N_1610,N_1912);
nor U2777 (N_2777,N_1110,N_1702);
xnor U2778 (N_2778,N_1161,N_1232);
or U2779 (N_2779,N_1685,N_1329);
nand U2780 (N_2780,N_1198,N_1193);
nor U2781 (N_2781,N_1336,N_1629);
nand U2782 (N_2782,N_1386,N_1426);
nor U2783 (N_2783,N_1860,N_1011);
xnor U2784 (N_2784,N_1758,N_1555);
xor U2785 (N_2785,N_1628,N_1869);
xnor U2786 (N_2786,N_1006,N_1855);
and U2787 (N_2787,N_1355,N_1974);
xor U2788 (N_2788,N_1643,N_1013);
or U2789 (N_2789,N_1918,N_1025);
nand U2790 (N_2790,N_1506,N_1748);
xnor U2791 (N_2791,N_1365,N_1557);
nor U2792 (N_2792,N_1883,N_1870);
xnor U2793 (N_2793,N_1127,N_1071);
nor U2794 (N_2794,N_1111,N_1331);
xor U2795 (N_2795,N_1232,N_1679);
and U2796 (N_2796,N_1166,N_1079);
or U2797 (N_2797,N_1883,N_1471);
or U2798 (N_2798,N_1525,N_1474);
or U2799 (N_2799,N_1779,N_1367);
or U2800 (N_2800,N_1273,N_1482);
xor U2801 (N_2801,N_1997,N_1006);
nor U2802 (N_2802,N_1012,N_1680);
nor U2803 (N_2803,N_1451,N_1834);
nand U2804 (N_2804,N_1378,N_1489);
nor U2805 (N_2805,N_1011,N_1869);
or U2806 (N_2806,N_1904,N_1324);
nor U2807 (N_2807,N_1657,N_1164);
xor U2808 (N_2808,N_1897,N_1907);
and U2809 (N_2809,N_1100,N_1905);
or U2810 (N_2810,N_1237,N_1709);
nand U2811 (N_2811,N_1936,N_1586);
nor U2812 (N_2812,N_1971,N_1427);
nor U2813 (N_2813,N_1809,N_1900);
or U2814 (N_2814,N_1175,N_1650);
nor U2815 (N_2815,N_1760,N_1181);
nor U2816 (N_2816,N_1335,N_1466);
or U2817 (N_2817,N_1278,N_1736);
nand U2818 (N_2818,N_1318,N_1065);
xor U2819 (N_2819,N_1381,N_1794);
nand U2820 (N_2820,N_1484,N_1902);
xnor U2821 (N_2821,N_1725,N_1471);
nand U2822 (N_2822,N_1915,N_1330);
nand U2823 (N_2823,N_1259,N_1633);
nand U2824 (N_2824,N_1226,N_1675);
nor U2825 (N_2825,N_1678,N_1048);
or U2826 (N_2826,N_1791,N_1666);
nor U2827 (N_2827,N_1656,N_1662);
and U2828 (N_2828,N_1574,N_1587);
or U2829 (N_2829,N_1028,N_1080);
or U2830 (N_2830,N_1715,N_1698);
xor U2831 (N_2831,N_1875,N_1964);
or U2832 (N_2832,N_1574,N_1324);
or U2833 (N_2833,N_1867,N_1626);
nor U2834 (N_2834,N_1311,N_1567);
or U2835 (N_2835,N_1416,N_1525);
xnor U2836 (N_2836,N_1800,N_1042);
xnor U2837 (N_2837,N_1317,N_1199);
nor U2838 (N_2838,N_1898,N_1221);
or U2839 (N_2839,N_1951,N_1122);
and U2840 (N_2840,N_1052,N_1611);
xnor U2841 (N_2841,N_1850,N_1832);
and U2842 (N_2842,N_1585,N_1642);
or U2843 (N_2843,N_1654,N_1002);
xnor U2844 (N_2844,N_1020,N_1380);
and U2845 (N_2845,N_1569,N_1275);
nand U2846 (N_2846,N_1886,N_1313);
or U2847 (N_2847,N_1256,N_1896);
xor U2848 (N_2848,N_1114,N_1431);
and U2849 (N_2849,N_1518,N_1314);
or U2850 (N_2850,N_1618,N_1606);
nor U2851 (N_2851,N_1294,N_1620);
nor U2852 (N_2852,N_1566,N_1090);
xor U2853 (N_2853,N_1673,N_1185);
and U2854 (N_2854,N_1671,N_1435);
and U2855 (N_2855,N_1279,N_1552);
nor U2856 (N_2856,N_1967,N_1898);
or U2857 (N_2857,N_1088,N_1223);
and U2858 (N_2858,N_1139,N_1519);
nand U2859 (N_2859,N_1397,N_1102);
nand U2860 (N_2860,N_1355,N_1344);
nor U2861 (N_2861,N_1283,N_1498);
xnor U2862 (N_2862,N_1172,N_1697);
or U2863 (N_2863,N_1439,N_1906);
nand U2864 (N_2864,N_1914,N_1075);
and U2865 (N_2865,N_1183,N_1033);
or U2866 (N_2866,N_1180,N_1237);
nand U2867 (N_2867,N_1624,N_1726);
nor U2868 (N_2868,N_1109,N_1790);
or U2869 (N_2869,N_1293,N_1079);
or U2870 (N_2870,N_1368,N_1219);
nand U2871 (N_2871,N_1776,N_1932);
xor U2872 (N_2872,N_1860,N_1883);
or U2873 (N_2873,N_1855,N_1256);
or U2874 (N_2874,N_1756,N_1891);
and U2875 (N_2875,N_1748,N_1349);
and U2876 (N_2876,N_1263,N_1542);
and U2877 (N_2877,N_1016,N_1548);
or U2878 (N_2878,N_1435,N_1271);
nand U2879 (N_2879,N_1408,N_1907);
nand U2880 (N_2880,N_1771,N_1494);
and U2881 (N_2881,N_1546,N_1328);
xnor U2882 (N_2882,N_1904,N_1445);
xor U2883 (N_2883,N_1980,N_1684);
or U2884 (N_2884,N_1080,N_1992);
xnor U2885 (N_2885,N_1456,N_1288);
and U2886 (N_2886,N_1155,N_1931);
or U2887 (N_2887,N_1229,N_1769);
and U2888 (N_2888,N_1670,N_1282);
nand U2889 (N_2889,N_1804,N_1997);
nand U2890 (N_2890,N_1797,N_1230);
nand U2891 (N_2891,N_1984,N_1545);
or U2892 (N_2892,N_1885,N_1751);
nor U2893 (N_2893,N_1026,N_1187);
nor U2894 (N_2894,N_1059,N_1024);
nand U2895 (N_2895,N_1885,N_1081);
or U2896 (N_2896,N_1342,N_1822);
and U2897 (N_2897,N_1667,N_1991);
or U2898 (N_2898,N_1655,N_1675);
or U2899 (N_2899,N_1613,N_1604);
and U2900 (N_2900,N_1102,N_1871);
xor U2901 (N_2901,N_1025,N_1702);
or U2902 (N_2902,N_1710,N_1972);
nor U2903 (N_2903,N_1476,N_1002);
nor U2904 (N_2904,N_1436,N_1170);
and U2905 (N_2905,N_1194,N_1000);
and U2906 (N_2906,N_1590,N_1056);
nor U2907 (N_2907,N_1847,N_1566);
nand U2908 (N_2908,N_1309,N_1976);
or U2909 (N_2909,N_1734,N_1554);
nand U2910 (N_2910,N_1704,N_1811);
or U2911 (N_2911,N_1538,N_1570);
xor U2912 (N_2912,N_1983,N_1070);
nand U2913 (N_2913,N_1661,N_1021);
nand U2914 (N_2914,N_1612,N_1102);
or U2915 (N_2915,N_1561,N_1271);
and U2916 (N_2916,N_1423,N_1172);
nor U2917 (N_2917,N_1486,N_1516);
nor U2918 (N_2918,N_1839,N_1268);
xor U2919 (N_2919,N_1867,N_1751);
xor U2920 (N_2920,N_1610,N_1486);
nand U2921 (N_2921,N_1016,N_1818);
or U2922 (N_2922,N_1788,N_1694);
nand U2923 (N_2923,N_1454,N_1714);
xnor U2924 (N_2924,N_1610,N_1755);
xnor U2925 (N_2925,N_1408,N_1029);
xnor U2926 (N_2926,N_1949,N_1373);
xnor U2927 (N_2927,N_1674,N_1272);
or U2928 (N_2928,N_1975,N_1257);
nand U2929 (N_2929,N_1107,N_1614);
or U2930 (N_2930,N_1923,N_1888);
xnor U2931 (N_2931,N_1202,N_1126);
and U2932 (N_2932,N_1757,N_1487);
xnor U2933 (N_2933,N_1476,N_1708);
nor U2934 (N_2934,N_1572,N_1821);
and U2935 (N_2935,N_1811,N_1281);
and U2936 (N_2936,N_1517,N_1831);
and U2937 (N_2937,N_1082,N_1942);
or U2938 (N_2938,N_1367,N_1182);
nand U2939 (N_2939,N_1069,N_1558);
nor U2940 (N_2940,N_1052,N_1602);
nand U2941 (N_2941,N_1506,N_1742);
nor U2942 (N_2942,N_1959,N_1379);
nor U2943 (N_2943,N_1999,N_1328);
nor U2944 (N_2944,N_1456,N_1619);
and U2945 (N_2945,N_1485,N_1672);
and U2946 (N_2946,N_1557,N_1800);
or U2947 (N_2947,N_1264,N_1420);
nand U2948 (N_2948,N_1424,N_1721);
or U2949 (N_2949,N_1567,N_1141);
or U2950 (N_2950,N_1142,N_1779);
nor U2951 (N_2951,N_1535,N_1267);
xor U2952 (N_2952,N_1389,N_1030);
nand U2953 (N_2953,N_1863,N_1099);
and U2954 (N_2954,N_1880,N_1117);
nand U2955 (N_2955,N_1568,N_1115);
nand U2956 (N_2956,N_1581,N_1810);
or U2957 (N_2957,N_1263,N_1990);
and U2958 (N_2958,N_1748,N_1973);
xor U2959 (N_2959,N_1932,N_1489);
nor U2960 (N_2960,N_1845,N_1693);
nor U2961 (N_2961,N_1713,N_1076);
and U2962 (N_2962,N_1757,N_1730);
nand U2963 (N_2963,N_1887,N_1312);
xor U2964 (N_2964,N_1599,N_1613);
nand U2965 (N_2965,N_1044,N_1118);
nand U2966 (N_2966,N_1297,N_1510);
nor U2967 (N_2967,N_1745,N_1624);
or U2968 (N_2968,N_1964,N_1001);
and U2969 (N_2969,N_1988,N_1314);
xor U2970 (N_2970,N_1789,N_1843);
and U2971 (N_2971,N_1711,N_1752);
nand U2972 (N_2972,N_1666,N_1415);
nand U2973 (N_2973,N_1868,N_1229);
and U2974 (N_2974,N_1224,N_1124);
xor U2975 (N_2975,N_1096,N_1058);
and U2976 (N_2976,N_1442,N_1644);
and U2977 (N_2977,N_1785,N_1269);
nor U2978 (N_2978,N_1692,N_1476);
or U2979 (N_2979,N_1380,N_1155);
or U2980 (N_2980,N_1791,N_1362);
nor U2981 (N_2981,N_1447,N_1912);
xnor U2982 (N_2982,N_1854,N_1739);
xor U2983 (N_2983,N_1623,N_1792);
or U2984 (N_2984,N_1736,N_1524);
or U2985 (N_2985,N_1302,N_1036);
and U2986 (N_2986,N_1480,N_1947);
xor U2987 (N_2987,N_1703,N_1240);
and U2988 (N_2988,N_1211,N_1674);
nand U2989 (N_2989,N_1164,N_1037);
nand U2990 (N_2990,N_1894,N_1215);
nor U2991 (N_2991,N_1148,N_1379);
xnor U2992 (N_2992,N_1847,N_1596);
or U2993 (N_2993,N_1761,N_1999);
or U2994 (N_2994,N_1679,N_1565);
xor U2995 (N_2995,N_1300,N_1049);
nand U2996 (N_2996,N_1633,N_1863);
nor U2997 (N_2997,N_1224,N_1098);
xor U2998 (N_2998,N_1453,N_1039);
xor U2999 (N_2999,N_1139,N_1583);
or U3000 (N_3000,N_2269,N_2327);
and U3001 (N_3001,N_2298,N_2421);
and U3002 (N_3002,N_2429,N_2757);
and U3003 (N_3003,N_2857,N_2897);
and U3004 (N_3004,N_2791,N_2648);
and U3005 (N_3005,N_2081,N_2913);
nand U3006 (N_3006,N_2223,N_2909);
nand U3007 (N_3007,N_2474,N_2052);
nand U3008 (N_3008,N_2307,N_2664);
nand U3009 (N_3009,N_2898,N_2528);
nand U3010 (N_3010,N_2783,N_2501);
or U3011 (N_3011,N_2621,N_2957);
nor U3012 (N_3012,N_2361,N_2236);
nand U3013 (N_3013,N_2690,N_2806);
nor U3014 (N_3014,N_2565,N_2734);
xor U3015 (N_3015,N_2319,N_2162);
xor U3016 (N_3016,N_2753,N_2205);
or U3017 (N_3017,N_2095,N_2656);
xor U3018 (N_3018,N_2695,N_2659);
and U3019 (N_3019,N_2990,N_2500);
nand U3020 (N_3020,N_2297,N_2461);
or U3021 (N_3021,N_2965,N_2493);
xnor U3022 (N_3022,N_2536,N_2330);
nor U3023 (N_3023,N_2449,N_2517);
nor U3024 (N_3024,N_2371,N_2555);
nand U3025 (N_3025,N_2333,N_2038);
or U3026 (N_3026,N_2177,N_2360);
or U3027 (N_3027,N_2788,N_2584);
and U3028 (N_3028,N_2916,N_2434);
nand U3029 (N_3029,N_2132,N_2228);
and U3030 (N_3030,N_2426,N_2168);
nand U3031 (N_3031,N_2787,N_2573);
and U3032 (N_3032,N_2923,N_2586);
nand U3033 (N_3033,N_2531,N_2631);
xnor U3034 (N_3034,N_2422,N_2082);
nand U3035 (N_3035,N_2111,N_2520);
or U3036 (N_3036,N_2894,N_2482);
nand U3037 (N_3037,N_2152,N_2358);
or U3038 (N_3038,N_2660,N_2650);
nor U3039 (N_3039,N_2581,N_2614);
xnor U3040 (N_3040,N_2523,N_2697);
nand U3041 (N_3041,N_2314,N_2532);
nand U3042 (N_3042,N_2993,N_2864);
nand U3043 (N_3043,N_2835,N_2879);
xor U3044 (N_3044,N_2802,N_2811);
or U3045 (N_3045,N_2892,N_2473);
or U3046 (N_3046,N_2272,N_2069);
nor U3047 (N_3047,N_2174,N_2045);
and U3048 (N_3048,N_2277,N_2514);
nor U3049 (N_3049,N_2634,N_2287);
or U3050 (N_3050,N_2369,N_2293);
nor U3051 (N_3051,N_2165,N_2249);
nand U3052 (N_3052,N_2558,N_2605);
xnor U3053 (N_3053,N_2919,N_2109);
or U3054 (N_3054,N_2100,N_2533);
and U3055 (N_3055,N_2642,N_2796);
or U3056 (N_3056,N_2445,N_2946);
or U3057 (N_3057,N_2268,N_2748);
and U3058 (N_3058,N_2112,N_2678);
nand U3059 (N_3059,N_2063,N_2657);
or U3060 (N_3060,N_2896,N_2187);
nor U3061 (N_3061,N_2529,N_2043);
and U3062 (N_3062,N_2732,N_2550);
and U3063 (N_3063,N_2842,N_2543);
and U3064 (N_3064,N_2506,N_2255);
nand U3065 (N_3065,N_2870,N_2556);
nand U3066 (N_3066,N_2023,N_2746);
xor U3067 (N_3067,N_2686,N_2525);
xor U3068 (N_3068,N_2125,N_2803);
nand U3069 (N_3069,N_2188,N_2433);
nor U3070 (N_3070,N_2705,N_2601);
or U3071 (N_3071,N_2206,N_2008);
and U3072 (N_3072,N_2682,N_2486);
nor U3073 (N_3073,N_2831,N_2342);
nand U3074 (N_3074,N_2628,N_2513);
xnor U3075 (N_3075,N_2926,N_2773);
and U3076 (N_3076,N_2325,N_2604);
and U3077 (N_3077,N_2328,N_2074);
or U3078 (N_3078,N_2647,N_2674);
nand U3079 (N_3079,N_2197,N_2385);
and U3080 (N_3080,N_2781,N_2258);
and U3081 (N_3081,N_2457,N_2211);
nor U3082 (N_3082,N_2437,N_2460);
nand U3083 (N_3083,N_2042,N_2282);
or U3084 (N_3084,N_2171,N_2527);
nor U3085 (N_3085,N_2124,N_2175);
xor U3086 (N_3086,N_2311,N_2050);
xor U3087 (N_3087,N_2156,N_2012);
nand U3088 (N_3088,N_2379,N_2858);
nand U3089 (N_3089,N_2497,N_2480);
nand U3090 (N_3090,N_2276,N_2289);
nand U3091 (N_3091,N_2221,N_2538);
nor U3092 (N_3092,N_2088,N_2135);
xnor U3093 (N_3093,N_2428,N_2598);
nand U3094 (N_3094,N_2930,N_2729);
nand U3095 (N_3095,N_2475,N_2562);
xnor U3096 (N_3096,N_2256,N_2723);
nand U3097 (N_3097,N_2855,N_2104);
and U3098 (N_3098,N_2718,N_2530);
nor U3099 (N_3099,N_2317,N_2072);
nor U3100 (N_3100,N_2346,N_2015);
and U3101 (N_3101,N_2917,N_2947);
nand U3102 (N_3102,N_2242,N_2554);
xor U3103 (N_3103,N_2420,N_2488);
nand U3104 (N_3104,N_2900,N_2846);
or U3105 (N_3105,N_2170,N_2180);
xor U3106 (N_3106,N_2464,N_2724);
or U3107 (N_3107,N_2377,N_2058);
xor U3108 (N_3108,N_2146,N_2649);
nor U3109 (N_3109,N_2126,N_2215);
nand U3110 (N_3110,N_2395,N_2364);
xor U3111 (N_3111,N_2114,N_2906);
and U3112 (N_3112,N_2378,N_2545);
nand U3113 (N_3113,N_2003,N_2840);
nand U3114 (N_3114,N_2270,N_2071);
xnor U3115 (N_3115,N_2308,N_2374);
nand U3116 (N_3116,N_2696,N_2386);
nand U3117 (N_3117,N_2925,N_2133);
and U3118 (N_3118,N_2583,N_2606);
nand U3119 (N_3119,N_2341,N_2888);
or U3120 (N_3120,N_2768,N_2630);
nor U3121 (N_3121,N_2334,N_2663);
nor U3122 (N_3122,N_2733,N_2321);
nor U3123 (N_3123,N_2410,N_2243);
nand U3124 (N_3124,N_2975,N_2667);
nand U3125 (N_3125,N_2994,N_2966);
nand U3126 (N_3126,N_2511,N_2079);
and U3127 (N_3127,N_2294,N_2061);
nand U3128 (N_3128,N_2679,N_2713);
xnor U3129 (N_3129,N_2626,N_2116);
and U3130 (N_3130,N_2570,N_2105);
nand U3131 (N_3131,N_2617,N_2343);
or U3132 (N_3132,N_2625,N_2706);
or U3133 (N_3133,N_2235,N_2251);
nor U3134 (N_3134,N_2769,N_2995);
or U3135 (N_3135,N_2394,N_2708);
nor U3136 (N_3136,N_2782,N_2588);
nand U3137 (N_3137,N_2083,N_2406);
xnor U3138 (N_3138,N_2494,N_2024);
or U3139 (N_3139,N_2775,N_2335);
nor U3140 (N_3140,N_2885,N_2728);
nand U3141 (N_3141,N_2551,N_2292);
or U3142 (N_3142,N_2027,N_2914);
nand U3143 (N_3143,N_2717,N_2304);
or U3144 (N_3144,N_2873,N_2837);
xnor U3145 (N_3145,N_2875,N_2978);
and U3146 (N_3146,N_2259,N_2103);
or U3147 (N_3147,N_2026,N_2018);
or U3148 (N_3148,N_2752,N_2131);
nand U3149 (N_3149,N_2792,N_2466);
and U3150 (N_3150,N_2609,N_2329);
xor U3151 (N_3151,N_2789,N_2155);
nor U3152 (N_3152,N_2854,N_2405);
nor U3153 (N_3153,N_2833,N_2350);
or U3154 (N_3154,N_2208,N_2288);
xnor U3155 (N_3155,N_2618,N_2929);
xor U3156 (N_3156,N_2592,N_2407);
nor U3157 (N_3157,N_2381,N_2266);
xor U3158 (N_3158,N_2121,N_2693);
xnor U3159 (N_3159,N_2049,N_2167);
nand U3160 (N_3160,N_2143,N_2546);
nand U3161 (N_3161,N_2683,N_2295);
or U3162 (N_3162,N_2711,N_2987);
and U3163 (N_3163,N_2508,N_2694);
xnor U3164 (N_3164,N_2416,N_2344);
nand U3165 (N_3165,N_2939,N_2349);
or U3166 (N_3166,N_2007,N_2340);
xor U3167 (N_3167,N_2767,N_2560);
xor U3168 (N_3168,N_2305,N_2938);
nor U3169 (N_3169,N_2134,N_2549);
and U3170 (N_3170,N_2799,N_2227);
xnor U3171 (N_3171,N_2274,N_2602);
or U3172 (N_3172,N_2566,N_2302);
xnor U3173 (N_3173,N_2370,N_2563);
nand U3174 (N_3174,N_2337,N_2544);
nand U3175 (N_3175,N_2388,N_2755);
nand U3176 (N_3176,N_2633,N_2816);
nor U3177 (N_3177,N_2366,N_2039);
or U3178 (N_3178,N_2651,N_2323);
xnor U3179 (N_3179,N_2450,N_2593);
or U3180 (N_3180,N_2202,N_2579);
and U3181 (N_3181,N_2456,N_2680);
xor U3182 (N_3182,N_2413,N_2402);
and U3183 (N_3183,N_2964,N_2740);
nor U3184 (N_3184,N_2359,N_2832);
xor U3185 (N_3185,N_2653,N_2192);
and U3186 (N_3186,N_2970,N_2689);
nand U3187 (N_3187,N_2400,N_2285);
nand U3188 (N_3188,N_2485,N_2666);
or U3189 (N_3189,N_2091,N_2320);
xnor U3190 (N_3190,N_2595,N_2036);
nor U3191 (N_3191,N_2076,N_2128);
nor U3192 (N_3192,N_2891,N_2157);
or U3193 (N_3193,N_2830,N_2726);
nor U3194 (N_3194,N_2183,N_2025);
or U3195 (N_3195,N_2749,N_2448);
xor U3196 (N_3196,N_2931,N_2847);
and U3197 (N_3197,N_2950,N_2668);
xor U3198 (N_3198,N_2518,N_2046);
or U3199 (N_3199,N_2415,N_2299);
nand U3200 (N_3200,N_2615,N_2226);
nand U3201 (N_3201,N_2600,N_2438);
nand U3202 (N_3202,N_2179,N_2675);
nand U3203 (N_3203,N_2797,N_2470);
and U3204 (N_3204,N_2639,N_2887);
and U3205 (N_3205,N_2574,N_2540);
nor U3206 (N_3206,N_2213,N_2569);
or U3207 (N_3207,N_2611,N_2060);
xnor U3208 (N_3208,N_2764,N_2252);
and U3209 (N_3209,N_2765,N_2825);
or U3210 (N_3210,N_2159,N_2414);
and U3211 (N_3211,N_2547,N_2557);
or U3212 (N_3212,N_2062,N_2357);
nor U3213 (N_3213,N_2477,N_2827);
nand U3214 (N_3214,N_2120,N_2677);
and U3215 (N_3215,N_2849,N_2160);
nand U3216 (N_3216,N_2199,N_2915);
nand U3217 (N_3217,N_2430,N_2336);
nor U3218 (N_3218,N_2067,N_2890);
nand U3219 (N_3219,N_2954,N_2225);
and U3220 (N_3220,N_2315,N_2099);
xor U3221 (N_3221,N_2725,N_2110);
nor U3222 (N_3222,N_2412,N_2367);
nand U3223 (N_3223,N_2779,N_2844);
xnor U3224 (N_3224,N_2824,N_2423);
and U3225 (N_3225,N_2339,N_2318);
nor U3226 (N_3226,N_2921,N_2204);
nor U3227 (N_3227,N_2309,N_2878);
and U3228 (N_3228,N_2934,N_2087);
nand U3229 (N_3229,N_2130,N_2937);
nand U3230 (N_3230,N_2200,N_2047);
nor U3231 (N_3231,N_2669,N_2608);
nor U3232 (N_3232,N_2392,N_2097);
or U3233 (N_3233,N_2982,N_2056);
xor U3234 (N_3234,N_2471,N_2375);
xnor U3235 (N_3235,N_2229,N_2001);
or U3236 (N_3236,N_2967,N_2637);
or U3237 (N_3237,N_2784,N_2265);
or U3238 (N_3238,N_2214,N_2933);
nor U3239 (N_3239,N_2034,N_2490);
or U3240 (N_3240,N_2823,N_2845);
nor U3241 (N_3241,N_2141,N_2267);
xor U3242 (N_3242,N_2246,N_2762);
nor U3243 (N_3243,N_2670,N_2136);
nand U3244 (N_3244,N_2766,N_2248);
nand U3245 (N_3245,N_2011,N_2090);
nand U3246 (N_3246,N_2568,N_2901);
nand U3247 (N_3247,N_2424,N_2591);
or U3248 (N_3248,N_2075,N_2874);
nor U3249 (N_3249,N_2640,N_2638);
nor U3250 (N_3250,N_2841,N_2055);
or U3251 (N_3251,N_2492,N_2750);
and U3252 (N_3252,N_2498,N_2393);
xnor U3253 (N_3253,N_2941,N_2928);
nor U3254 (N_3254,N_2641,N_2092);
and U3255 (N_3255,N_2122,N_2149);
or U3256 (N_3256,N_2084,N_2190);
nor U3257 (N_3257,N_2869,N_2903);
or U3258 (N_3258,N_2231,N_2040);
nand U3259 (N_3259,N_2665,N_2093);
nor U3260 (N_3260,N_2700,N_2418);
xnor U3261 (N_3261,N_2943,N_2505);
nand U3262 (N_3262,N_2354,N_2240);
nand U3263 (N_3263,N_2247,N_2561);
xnor U3264 (N_3264,N_2409,N_2013);
or U3265 (N_3265,N_2658,N_2376);
or U3266 (N_3266,N_2963,N_2736);
and U3267 (N_3267,N_2113,N_2955);
and U3268 (N_3268,N_2280,N_2193);
nand U3269 (N_3269,N_2217,N_2998);
nand U3270 (N_3270,N_2912,N_2101);
xor U3271 (N_3271,N_2427,N_2182);
and U3272 (N_3272,N_2720,N_2326);
xor U3273 (N_3273,N_2291,N_2312);
nor U3274 (N_3274,N_2580,N_2624);
nand U3275 (N_3275,N_2715,N_2777);
xnor U3276 (N_3276,N_2281,N_2798);
and U3277 (N_3277,N_2189,N_2905);
and U3278 (N_3278,N_2576,N_2447);
xnor U3279 (N_3279,N_2403,N_2707);
nor U3280 (N_3280,N_2810,N_2237);
and U3281 (N_3281,N_2332,N_2463);
and U3282 (N_3282,N_2353,N_2117);
and U3283 (N_3283,N_2851,N_2699);
and U3284 (N_3284,N_2181,N_2028);
nand U3285 (N_3285,N_2852,N_2106);
or U3286 (N_3286,N_2057,N_2219);
nand U3287 (N_3287,N_2623,N_2397);
xnor U3288 (N_3288,N_2552,N_2218);
and U3289 (N_3289,N_2310,N_2861);
nor U3290 (N_3290,N_2949,N_2129);
and U3291 (N_3291,N_2883,N_2599);
and U3292 (N_3292,N_2212,N_2153);
or U3293 (N_3293,N_2942,N_2727);
xor U3294 (N_3294,N_2404,N_2399);
xor U3295 (N_3295,N_2279,N_2661);
nand U3296 (N_3296,N_2644,N_2073);
xnor U3297 (N_3297,N_2244,N_2973);
xor U3298 (N_3298,N_2163,N_2959);
and U3299 (N_3299,N_2991,N_2164);
nand U3300 (N_3300,N_2521,N_2721);
nor U3301 (N_3301,N_2988,N_2037);
or U3302 (N_3302,N_2805,N_2986);
nand U3303 (N_3303,N_2972,N_2968);
nor U3304 (N_3304,N_2564,N_2041);
or U3305 (N_3305,N_2924,N_2610);
or U3306 (N_3306,N_2347,N_2365);
or U3307 (N_3307,N_2989,N_2262);
nor U3308 (N_3308,N_2184,N_2983);
nand U3309 (N_3309,N_2742,N_2597);
nor U3310 (N_3310,N_2691,N_2054);
xor U3311 (N_3311,N_2484,N_2313);
nand U3312 (N_3312,N_2169,N_2085);
xnor U3313 (N_3313,N_2703,N_2822);
or U3314 (N_3314,N_2754,N_2737);
nand U3315 (N_3315,N_2194,N_2853);
xnor U3316 (N_3316,N_2324,N_2389);
nor U3317 (N_3317,N_2222,N_2951);
or U3318 (N_3318,N_2356,N_2716);
or U3319 (N_3319,N_2860,N_2839);
nor U3320 (N_3320,N_2064,N_2185);
nand U3321 (N_3321,N_2515,N_2889);
nand U3322 (N_3322,N_2451,N_2503);
nor U3323 (N_3323,N_2790,N_2144);
nand U3324 (N_3324,N_2303,N_2868);
and U3325 (N_3325,N_2384,N_2431);
and U3326 (N_3326,N_2476,N_2491);
xnor U3327 (N_3327,N_2345,N_2145);
and U3328 (N_3328,N_2077,N_2142);
and U3329 (N_3329,N_2817,N_2107);
xor U3330 (N_3330,N_2616,N_2387);
xnor U3331 (N_3331,N_2462,N_2089);
or U3332 (N_3332,N_2571,N_2301);
or U3333 (N_3333,N_2372,N_2051);
xor U3334 (N_3334,N_2880,N_2006);
nor U3335 (N_3335,N_2622,N_2985);
or U3336 (N_3336,N_2862,N_2760);
xnor U3337 (N_3337,N_2603,N_2070);
nor U3338 (N_3338,N_2710,N_2572);
xnor U3339 (N_3339,N_2390,N_2234);
and U3340 (N_3340,N_2785,N_2866);
or U3341 (N_3341,N_2035,N_2053);
or U3342 (N_3342,N_2882,N_2984);
nor U3343 (N_3343,N_2828,N_2944);
nand U3344 (N_3344,N_2684,N_2148);
or U3345 (N_3345,N_2032,N_2094);
or U3346 (N_3346,N_2322,N_2502);
or U3347 (N_3347,N_2698,N_2867);
nor U3348 (N_3348,N_2758,N_2741);
nor U3349 (N_3349,N_2607,N_2455);
nor U3350 (N_3350,N_2590,N_2865);
nor U3351 (N_3351,N_2818,N_2139);
nand U3352 (N_3352,N_2439,N_2997);
and U3353 (N_3353,N_2098,N_2881);
or U3354 (N_3354,N_2722,N_2958);
nor U3355 (N_3355,N_2363,N_2253);
and U3356 (N_3356,N_2316,N_2196);
or U3357 (N_3357,N_2654,N_2996);
nand U3358 (N_3358,N_2432,N_2468);
xor U3359 (N_3359,N_2065,N_2971);
xnor U3360 (N_3360,N_2102,N_2275);
xor U3361 (N_3361,N_2756,N_2948);
or U3362 (N_3362,N_2000,N_2239);
or U3363 (N_3363,N_2613,N_2636);
xnor U3364 (N_3364,N_2884,N_2738);
nand U3365 (N_3365,N_2059,N_2140);
nand U3366 (N_3366,N_2351,N_2632);
or U3367 (N_3367,N_2922,N_2961);
and U3368 (N_3368,N_2662,N_2022);
or U3369 (N_3369,N_2489,N_2780);
and U3370 (N_3370,N_2553,N_2398);
and U3371 (N_3371,N_2872,N_2735);
nand U3372 (N_3372,N_2453,N_2786);
xor U3373 (N_3373,N_2440,N_2016);
and U3374 (N_3374,N_2976,N_2945);
nor U3375 (N_3375,N_2232,N_2577);
xnor U3376 (N_3376,N_2719,N_2815);
xor U3377 (N_3377,N_2730,N_2701);
and U3378 (N_3378,N_2005,N_2209);
and U3379 (N_3379,N_2655,N_2373);
and U3380 (N_3380,N_2048,N_2210);
xnor U3381 (N_3381,N_2108,N_2150);
nand U3382 (N_3382,N_2794,N_2382);
nor U3383 (N_3383,N_2010,N_2645);
xnor U3384 (N_3384,N_2672,N_2744);
xor U3385 (N_3385,N_2338,N_2178);
or U3386 (N_3386,N_2216,N_2355);
and U3387 (N_3387,N_2688,N_2979);
and U3388 (N_3388,N_2014,N_2425);
and U3389 (N_3389,N_2776,N_2856);
nand U3390 (N_3390,N_2203,N_2250);
xnor U3391 (N_3391,N_2245,N_2257);
or U3392 (N_3392,N_2383,N_2763);
nand U3393 (N_3393,N_2899,N_2459);
nand U3394 (N_3394,N_2516,N_2186);
or U3395 (N_3395,N_2619,N_2368);
or U3396 (N_3396,N_2834,N_2408);
nor U3397 (N_3397,N_2956,N_2031);
nor U3398 (N_3398,N_2800,N_2524);
nand U3399 (N_3399,N_2118,N_2920);
nand U3400 (N_3400,N_2801,N_2522);
and U3401 (N_3401,N_2709,N_2261);
nand U3402 (N_3402,N_2066,N_2138);
nor U3403 (N_3403,N_2458,N_2263);
nand U3404 (N_3404,N_2969,N_2396);
and U3405 (N_3405,N_2286,N_2712);
xnor U3406 (N_3406,N_2620,N_2499);
nand U3407 (N_3407,N_2436,N_2029);
xnor U3408 (N_3408,N_2173,N_2283);
and U3409 (N_3409,N_2172,N_2469);
and U3410 (N_3410,N_2877,N_2567);
xnor U3411 (N_3411,N_2161,N_2578);
nor U3412 (N_3412,N_2539,N_2548);
or U3413 (N_3413,N_2886,N_2962);
nor U3414 (N_3414,N_2331,N_2452);
or U3415 (N_3415,N_2838,N_2770);
xor U3416 (N_3416,N_2936,N_2362);
and U3417 (N_3417,N_2068,N_2575);
and U3418 (N_3418,N_2859,N_2278);
xnor U3419 (N_3419,N_2671,N_2454);
or U3420 (N_3420,N_2465,N_2587);
or U3421 (N_3421,N_2809,N_2086);
or U3422 (N_3422,N_2685,N_2559);
nand U3423 (N_3423,N_2932,N_2443);
nor U3424 (N_3424,N_2017,N_2585);
xor U3425 (N_3425,N_2850,N_2676);
nor U3426 (N_3426,N_2980,N_2201);
nand U3427 (N_3427,N_2537,N_2127);
nand U3428 (N_3428,N_2731,N_2472);
xnor U3429 (N_3429,N_2795,N_2123);
and U3430 (N_3430,N_2198,N_2254);
or U3431 (N_3431,N_2441,N_2444);
or U3432 (N_3432,N_2238,N_2176);
nand U3433 (N_3433,N_2743,N_2927);
or U3434 (N_3434,N_2692,N_2220);
nor U3435 (N_3435,N_2487,N_2166);
and U3436 (N_3436,N_2496,N_2137);
nand U3437 (N_3437,N_2080,N_2774);
and U3438 (N_3438,N_2541,N_2435);
or U3439 (N_3439,N_2004,N_2848);
or U3440 (N_3440,N_2230,N_2296);
nor U3441 (N_3441,N_2195,N_2911);
nor U3442 (N_3442,N_2119,N_2687);
xnor U3443 (N_3443,N_2761,N_2526);
and U3444 (N_3444,N_2977,N_2348);
nand U3445 (N_3445,N_2380,N_2714);
and U3446 (N_3446,N_2030,N_2495);
or U3447 (N_3447,N_2702,N_2273);
nand U3448 (N_3448,N_2417,N_2519);
xnor U3449 (N_3449,N_2271,N_2411);
xor U3450 (N_3450,N_2940,N_2751);
or U3451 (N_3451,N_2509,N_2044);
nand U3452 (N_3452,N_2033,N_2918);
or U3453 (N_3453,N_2871,N_2673);
nor U3454 (N_3454,N_2772,N_2020);
xor U3455 (N_3455,N_2652,N_2306);
and U3456 (N_3456,N_2224,N_2158);
and U3457 (N_3457,N_2813,N_2019);
or U3458 (N_3458,N_2151,N_2808);
nand U3459 (N_3459,N_2935,N_2300);
xor U3460 (N_3460,N_2635,N_2233);
and U3461 (N_3461,N_2907,N_2290);
xor U3462 (N_3462,N_2115,N_2863);
nor U3463 (N_3463,N_2704,N_2612);
xor U3464 (N_3464,N_2895,N_2078);
nor U3465 (N_3465,N_2483,N_2446);
nand U3466 (N_3466,N_2681,N_2419);
xor U3467 (N_3467,N_2542,N_2952);
and U3468 (N_3468,N_2876,N_2627);
nor U3469 (N_3469,N_2260,N_2009);
nor U3470 (N_3470,N_2960,N_2992);
and U3471 (N_3471,N_2771,N_2819);
nand U3472 (N_3472,N_2843,N_2241);
and U3473 (N_3473,N_2504,N_2826);
xnor U3474 (N_3474,N_2154,N_2191);
nand U3475 (N_3475,N_2999,N_2745);
or U3476 (N_3476,N_2804,N_2908);
and U3477 (N_3477,N_2629,N_2442);
and U3478 (N_3478,N_2512,N_2829);
nand U3479 (N_3479,N_2147,N_2535);
or U3480 (N_3480,N_2953,N_2479);
or U3481 (N_3481,N_2739,N_2836);
nand U3482 (N_3482,N_2902,N_2747);
nor U3483 (N_3483,N_2534,N_2352);
or U3484 (N_3484,N_2401,N_2478);
xor U3485 (N_3485,N_2589,N_2778);
nand U3486 (N_3486,N_2643,N_2507);
or U3487 (N_3487,N_2981,N_2910);
and U3488 (N_3488,N_2814,N_2582);
nor U3489 (N_3489,N_2391,N_2021);
xor U3490 (N_3490,N_2759,N_2481);
xnor U3491 (N_3491,N_2793,N_2207);
xnor U3492 (N_3492,N_2646,N_2096);
or U3493 (N_3493,N_2812,N_2821);
and U3494 (N_3494,N_2974,N_2596);
xor U3495 (N_3495,N_2264,N_2820);
nor U3496 (N_3496,N_2467,N_2002);
and U3497 (N_3497,N_2807,N_2594);
and U3498 (N_3498,N_2893,N_2904);
nor U3499 (N_3499,N_2284,N_2510);
nand U3500 (N_3500,N_2852,N_2673);
or U3501 (N_3501,N_2125,N_2312);
xnor U3502 (N_3502,N_2126,N_2869);
and U3503 (N_3503,N_2738,N_2263);
nand U3504 (N_3504,N_2031,N_2477);
xnor U3505 (N_3505,N_2005,N_2327);
nor U3506 (N_3506,N_2818,N_2066);
nor U3507 (N_3507,N_2726,N_2372);
or U3508 (N_3508,N_2999,N_2615);
nand U3509 (N_3509,N_2543,N_2155);
and U3510 (N_3510,N_2721,N_2805);
xor U3511 (N_3511,N_2741,N_2701);
xnor U3512 (N_3512,N_2918,N_2936);
xnor U3513 (N_3513,N_2571,N_2934);
xnor U3514 (N_3514,N_2699,N_2981);
nor U3515 (N_3515,N_2786,N_2924);
nor U3516 (N_3516,N_2231,N_2256);
nand U3517 (N_3517,N_2881,N_2096);
or U3518 (N_3518,N_2723,N_2080);
and U3519 (N_3519,N_2306,N_2653);
nor U3520 (N_3520,N_2940,N_2430);
and U3521 (N_3521,N_2232,N_2520);
nand U3522 (N_3522,N_2507,N_2313);
xnor U3523 (N_3523,N_2251,N_2915);
and U3524 (N_3524,N_2519,N_2211);
nand U3525 (N_3525,N_2678,N_2787);
nand U3526 (N_3526,N_2035,N_2199);
nor U3527 (N_3527,N_2292,N_2801);
or U3528 (N_3528,N_2678,N_2011);
and U3529 (N_3529,N_2520,N_2789);
xnor U3530 (N_3530,N_2068,N_2643);
xor U3531 (N_3531,N_2752,N_2361);
xnor U3532 (N_3532,N_2109,N_2886);
and U3533 (N_3533,N_2614,N_2588);
or U3534 (N_3534,N_2017,N_2851);
or U3535 (N_3535,N_2453,N_2736);
xnor U3536 (N_3536,N_2709,N_2344);
nor U3537 (N_3537,N_2774,N_2815);
or U3538 (N_3538,N_2687,N_2448);
nand U3539 (N_3539,N_2617,N_2601);
or U3540 (N_3540,N_2966,N_2220);
nor U3541 (N_3541,N_2462,N_2203);
nor U3542 (N_3542,N_2194,N_2647);
or U3543 (N_3543,N_2323,N_2836);
or U3544 (N_3544,N_2333,N_2542);
or U3545 (N_3545,N_2764,N_2499);
and U3546 (N_3546,N_2883,N_2580);
xnor U3547 (N_3547,N_2651,N_2373);
nand U3548 (N_3548,N_2866,N_2574);
nor U3549 (N_3549,N_2666,N_2776);
or U3550 (N_3550,N_2930,N_2621);
or U3551 (N_3551,N_2453,N_2258);
nand U3552 (N_3552,N_2355,N_2952);
and U3553 (N_3553,N_2387,N_2684);
and U3554 (N_3554,N_2221,N_2471);
nor U3555 (N_3555,N_2782,N_2338);
or U3556 (N_3556,N_2862,N_2164);
nor U3557 (N_3557,N_2141,N_2982);
xnor U3558 (N_3558,N_2861,N_2549);
nand U3559 (N_3559,N_2383,N_2410);
and U3560 (N_3560,N_2403,N_2103);
nor U3561 (N_3561,N_2545,N_2202);
nand U3562 (N_3562,N_2569,N_2533);
nand U3563 (N_3563,N_2704,N_2732);
and U3564 (N_3564,N_2630,N_2618);
nor U3565 (N_3565,N_2797,N_2012);
xor U3566 (N_3566,N_2567,N_2115);
nor U3567 (N_3567,N_2729,N_2027);
nand U3568 (N_3568,N_2086,N_2427);
or U3569 (N_3569,N_2126,N_2031);
xnor U3570 (N_3570,N_2129,N_2045);
nor U3571 (N_3571,N_2261,N_2859);
xnor U3572 (N_3572,N_2189,N_2650);
xor U3573 (N_3573,N_2502,N_2131);
nor U3574 (N_3574,N_2838,N_2115);
and U3575 (N_3575,N_2292,N_2707);
and U3576 (N_3576,N_2552,N_2548);
and U3577 (N_3577,N_2970,N_2403);
nor U3578 (N_3578,N_2187,N_2038);
and U3579 (N_3579,N_2925,N_2048);
and U3580 (N_3580,N_2775,N_2838);
and U3581 (N_3581,N_2139,N_2808);
or U3582 (N_3582,N_2120,N_2638);
xnor U3583 (N_3583,N_2865,N_2442);
or U3584 (N_3584,N_2468,N_2761);
nand U3585 (N_3585,N_2958,N_2899);
nand U3586 (N_3586,N_2726,N_2086);
nor U3587 (N_3587,N_2916,N_2598);
nand U3588 (N_3588,N_2907,N_2789);
or U3589 (N_3589,N_2431,N_2001);
nand U3590 (N_3590,N_2385,N_2379);
and U3591 (N_3591,N_2562,N_2938);
xor U3592 (N_3592,N_2179,N_2040);
xnor U3593 (N_3593,N_2954,N_2131);
xor U3594 (N_3594,N_2808,N_2747);
or U3595 (N_3595,N_2676,N_2723);
or U3596 (N_3596,N_2172,N_2789);
nand U3597 (N_3597,N_2067,N_2048);
xnor U3598 (N_3598,N_2695,N_2627);
nor U3599 (N_3599,N_2824,N_2269);
xor U3600 (N_3600,N_2591,N_2222);
xnor U3601 (N_3601,N_2900,N_2774);
and U3602 (N_3602,N_2341,N_2189);
or U3603 (N_3603,N_2504,N_2330);
xnor U3604 (N_3604,N_2449,N_2450);
nand U3605 (N_3605,N_2138,N_2831);
xor U3606 (N_3606,N_2071,N_2265);
and U3607 (N_3607,N_2397,N_2385);
xor U3608 (N_3608,N_2366,N_2035);
nor U3609 (N_3609,N_2657,N_2202);
or U3610 (N_3610,N_2866,N_2281);
or U3611 (N_3611,N_2787,N_2057);
xnor U3612 (N_3612,N_2699,N_2826);
xnor U3613 (N_3613,N_2138,N_2140);
and U3614 (N_3614,N_2334,N_2527);
and U3615 (N_3615,N_2780,N_2630);
nor U3616 (N_3616,N_2443,N_2190);
xnor U3617 (N_3617,N_2060,N_2795);
nand U3618 (N_3618,N_2687,N_2856);
and U3619 (N_3619,N_2314,N_2421);
or U3620 (N_3620,N_2681,N_2874);
nor U3621 (N_3621,N_2048,N_2832);
nand U3622 (N_3622,N_2904,N_2922);
and U3623 (N_3623,N_2968,N_2555);
nor U3624 (N_3624,N_2425,N_2192);
or U3625 (N_3625,N_2169,N_2918);
and U3626 (N_3626,N_2301,N_2593);
and U3627 (N_3627,N_2140,N_2697);
nand U3628 (N_3628,N_2935,N_2963);
xnor U3629 (N_3629,N_2688,N_2766);
xor U3630 (N_3630,N_2202,N_2832);
or U3631 (N_3631,N_2117,N_2369);
and U3632 (N_3632,N_2732,N_2768);
xnor U3633 (N_3633,N_2705,N_2027);
or U3634 (N_3634,N_2314,N_2523);
xor U3635 (N_3635,N_2744,N_2901);
or U3636 (N_3636,N_2819,N_2831);
xor U3637 (N_3637,N_2752,N_2074);
or U3638 (N_3638,N_2158,N_2160);
xnor U3639 (N_3639,N_2866,N_2124);
or U3640 (N_3640,N_2093,N_2197);
or U3641 (N_3641,N_2831,N_2188);
xor U3642 (N_3642,N_2192,N_2830);
nand U3643 (N_3643,N_2990,N_2527);
xor U3644 (N_3644,N_2825,N_2513);
and U3645 (N_3645,N_2751,N_2125);
and U3646 (N_3646,N_2962,N_2655);
and U3647 (N_3647,N_2379,N_2619);
or U3648 (N_3648,N_2053,N_2339);
xnor U3649 (N_3649,N_2930,N_2751);
and U3650 (N_3650,N_2077,N_2722);
or U3651 (N_3651,N_2147,N_2386);
nor U3652 (N_3652,N_2598,N_2928);
nand U3653 (N_3653,N_2877,N_2562);
nor U3654 (N_3654,N_2987,N_2593);
nor U3655 (N_3655,N_2988,N_2557);
and U3656 (N_3656,N_2378,N_2918);
and U3657 (N_3657,N_2098,N_2332);
and U3658 (N_3658,N_2306,N_2073);
nand U3659 (N_3659,N_2922,N_2877);
xnor U3660 (N_3660,N_2889,N_2960);
or U3661 (N_3661,N_2125,N_2257);
xnor U3662 (N_3662,N_2522,N_2096);
and U3663 (N_3663,N_2675,N_2338);
and U3664 (N_3664,N_2613,N_2575);
and U3665 (N_3665,N_2908,N_2735);
and U3666 (N_3666,N_2889,N_2548);
or U3667 (N_3667,N_2097,N_2635);
xnor U3668 (N_3668,N_2864,N_2372);
or U3669 (N_3669,N_2855,N_2023);
xnor U3670 (N_3670,N_2723,N_2960);
and U3671 (N_3671,N_2167,N_2600);
nor U3672 (N_3672,N_2448,N_2963);
nor U3673 (N_3673,N_2832,N_2604);
or U3674 (N_3674,N_2633,N_2858);
nor U3675 (N_3675,N_2389,N_2323);
and U3676 (N_3676,N_2215,N_2312);
nand U3677 (N_3677,N_2643,N_2816);
and U3678 (N_3678,N_2892,N_2735);
or U3679 (N_3679,N_2056,N_2079);
nor U3680 (N_3680,N_2675,N_2752);
nand U3681 (N_3681,N_2584,N_2624);
xnor U3682 (N_3682,N_2537,N_2101);
nand U3683 (N_3683,N_2064,N_2563);
nor U3684 (N_3684,N_2527,N_2492);
xnor U3685 (N_3685,N_2023,N_2255);
xor U3686 (N_3686,N_2209,N_2476);
nor U3687 (N_3687,N_2386,N_2638);
or U3688 (N_3688,N_2623,N_2555);
and U3689 (N_3689,N_2228,N_2985);
xnor U3690 (N_3690,N_2190,N_2945);
nor U3691 (N_3691,N_2361,N_2387);
and U3692 (N_3692,N_2940,N_2148);
xor U3693 (N_3693,N_2042,N_2272);
and U3694 (N_3694,N_2200,N_2291);
and U3695 (N_3695,N_2841,N_2019);
xor U3696 (N_3696,N_2828,N_2667);
or U3697 (N_3697,N_2956,N_2903);
and U3698 (N_3698,N_2972,N_2799);
or U3699 (N_3699,N_2563,N_2524);
and U3700 (N_3700,N_2625,N_2596);
nor U3701 (N_3701,N_2498,N_2610);
or U3702 (N_3702,N_2589,N_2265);
xor U3703 (N_3703,N_2358,N_2039);
or U3704 (N_3704,N_2897,N_2565);
xor U3705 (N_3705,N_2941,N_2165);
nor U3706 (N_3706,N_2504,N_2747);
or U3707 (N_3707,N_2031,N_2060);
and U3708 (N_3708,N_2962,N_2305);
and U3709 (N_3709,N_2440,N_2856);
nor U3710 (N_3710,N_2477,N_2469);
xor U3711 (N_3711,N_2548,N_2844);
nand U3712 (N_3712,N_2826,N_2328);
nor U3713 (N_3713,N_2207,N_2409);
or U3714 (N_3714,N_2507,N_2362);
and U3715 (N_3715,N_2984,N_2484);
nand U3716 (N_3716,N_2459,N_2023);
and U3717 (N_3717,N_2047,N_2223);
or U3718 (N_3718,N_2933,N_2468);
and U3719 (N_3719,N_2955,N_2321);
nor U3720 (N_3720,N_2760,N_2903);
nand U3721 (N_3721,N_2129,N_2408);
nand U3722 (N_3722,N_2325,N_2525);
or U3723 (N_3723,N_2087,N_2163);
or U3724 (N_3724,N_2606,N_2338);
or U3725 (N_3725,N_2655,N_2964);
xor U3726 (N_3726,N_2225,N_2059);
or U3727 (N_3727,N_2940,N_2400);
xnor U3728 (N_3728,N_2618,N_2566);
nand U3729 (N_3729,N_2766,N_2203);
nor U3730 (N_3730,N_2782,N_2265);
nand U3731 (N_3731,N_2913,N_2123);
nand U3732 (N_3732,N_2751,N_2484);
nand U3733 (N_3733,N_2985,N_2550);
or U3734 (N_3734,N_2548,N_2908);
xor U3735 (N_3735,N_2410,N_2723);
nor U3736 (N_3736,N_2201,N_2513);
or U3737 (N_3737,N_2884,N_2801);
and U3738 (N_3738,N_2573,N_2690);
nor U3739 (N_3739,N_2401,N_2185);
nand U3740 (N_3740,N_2527,N_2652);
and U3741 (N_3741,N_2024,N_2147);
nand U3742 (N_3742,N_2058,N_2397);
nand U3743 (N_3743,N_2008,N_2542);
xnor U3744 (N_3744,N_2704,N_2200);
nor U3745 (N_3745,N_2533,N_2064);
nor U3746 (N_3746,N_2959,N_2604);
nand U3747 (N_3747,N_2318,N_2951);
nand U3748 (N_3748,N_2920,N_2361);
nand U3749 (N_3749,N_2394,N_2896);
nand U3750 (N_3750,N_2674,N_2404);
nand U3751 (N_3751,N_2770,N_2855);
and U3752 (N_3752,N_2499,N_2993);
nand U3753 (N_3753,N_2200,N_2057);
xnor U3754 (N_3754,N_2883,N_2328);
or U3755 (N_3755,N_2377,N_2351);
nor U3756 (N_3756,N_2187,N_2380);
and U3757 (N_3757,N_2153,N_2179);
nor U3758 (N_3758,N_2326,N_2565);
xor U3759 (N_3759,N_2486,N_2513);
nor U3760 (N_3760,N_2636,N_2024);
nand U3761 (N_3761,N_2749,N_2775);
xnor U3762 (N_3762,N_2610,N_2385);
and U3763 (N_3763,N_2972,N_2219);
nor U3764 (N_3764,N_2323,N_2149);
or U3765 (N_3765,N_2272,N_2304);
nor U3766 (N_3766,N_2885,N_2480);
nor U3767 (N_3767,N_2813,N_2117);
nor U3768 (N_3768,N_2362,N_2150);
xor U3769 (N_3769,N_2922,N_2569);
nand U3770 (N_3770,N_2740,N_2709);
or U3771 (N_3771,N_2770,N_2651);
nor U3772 (N_3772,N_2119,N_2680);
nand U3773 (N_3773,N_2708,N_2528);
nand U3774 (N_3774,N_2633,N_2483);
nor U3775 (N_3775,N_2098,N_2397);
xnor U3776 (N_3776,N_2010,N_2950);
xor U3777 (N_3777,N_2284,N_2088);
xnor U3778 (N_3778,N_2219,N_2258);
nor U3779 (N_3779,N_2008,N_2217);
or U3780 (N_3780,N_2312,N_2289);
nand U3781 (N_3781,N_2942,N_2598);
nor U3782 (N_3782,N_2247,N_2845);
nor U3783 (N_3783,N_2356,N_2123);
and U3784 (N_3784,N_2392,N_2203);
nand U3785 (N_3785,N_2766,N_2675);
and U3786 (N_3786,N_2907,N_2520);
and U3787 (N_3787,N_2403,N_2162);
xor U3788 (N_3788,N_2799,N_2291);
nor U3789 (N_3789,N_2818,N_2172);
nor U3790 (N_3790,N_2703,N_2951);
xnor U3791 (N_3791,N_2930,N_2259);
nor U3792 (N_3792,N_2721,N_2698);
and U3793 (N_3793,N_2874,N_2483);
nor U3794 (N_3794,N_2797,N_2269);
or U3795 (N_3795,N_2023,N_2021);
and U3796 (N_3796,N_2935,N_2942);
and U3797 (N_3797,N_2620,N_2887);
nand U3798 (N_3798,N_2893,N_2199);
and U3799 (N_3799,N_2726,N_2275);
or U3800 (N_3800,N_2586,N_2200);
or U3801 (N_3801,N_2152,N_2108);
or U3802 (N_3802,N_2348,N_2673);
nor U3803 (N_3803,N_2097,N_2206);
xor U3804 (N_3804,N_2162,N_2990);
or U3805 (N_3805,N_2072,N_2670);
nand U3806 (N_3806,N_2767,N_2327);
xnor U3807 (N_3807,N_2870,N_2140);
or U3808 (N_3808,N_2550,N_2556);
and U3809 (N_3809,N_2312,N_2418);
xnor U3810 (N_3810,N_2767,N_2858);
nand U3811 (N_3811,N_2726,N_2923);
xnor U3812 (N_3812,N_2149,N_2555);
nand U3813 (N_3813,N_2418,N_2609);
and U3814 (N_3814,N_2458,N_2676);
nand U3815 (N_3815,N_2061,N_2245);
xnor U3816 (N_3816,N_2288,N_2648);
nor U3817 (N_3817,N_2573,N_2665);
xor U3818 (N_3818,N_2482,N_2869);
nor U3819 (N_3819,N_2914,N_2829);
nor U3820 (N_3820,N_2922,N_2522);
and U3821 (N_3821,N_2179,N_2583);
nor U3822 (N_3822,N_2897,N_2915);
or U3823 (N_3823,N_2540,N_2227);
nand U3824 (N_3824,N_2504,N_2890);
nor U3825 (N_3825,N_2960,N_2464);
nand U3826 (N_3826,N_2850,N_2841);
and U3827 (N_3827,N_2888,N_2747);
nand U3828 (N_3828,N_2310,N_2441);
nand U3829 (N_3829,N_2312,N_2879);
nand U3830 (N_3830,N_2364,N_2343);
or U3831 (N_3831,N_2430,N_2497);
or U3832 (N_3832,N_2215,N_2885);
xor U3833 (N_3833,N_2776,N_2379);
and U3834 (N_3834,N_2700,N_2424);
nand U3835 (N_3835,N_2103,N_2211);
or U3836 (N_3836,N_2964,N_2221);
or U3837 (N_3837,N_2685,N_2449);
xor U3838 (N_3838,N_2195,N_2581);
nand U3839 (N_3839,N_2511,N_2833);
nand U3840 (N_3840,N_2974,N_2186);
and U3841 (N_3841,N_2689,N_2218);
and U3842 (N_3842,N_2267,N_2281);
nor U3843 (N_3843,N_2258,N_2373);
xor U3844 (N_3844,N_2093,N_2354);
nand U3845 (N_3845,N_2942,N_2934);
and U3846 (N_3846,N_2344,N_2222);
and U3847 (N_3847,N_2802,N_2052);
nor U3848 (N_3848,N_2612,N_2289);
nand U3849 (N_3849,N_2432,N_2725);
nand U3850 (N_3850,N_2655,N_2255);
nand U3851 (N_3851,N_2610,N_2702);
and U3852 (N_3852,N_2186,N_2600);
nand U3853 (N_3853,N_2468,N_2993);
xor U3854 (N_3854,N_2981,N_2627);
nor U3855 (N_3855,N_2922,N_2114);
and U3856 (N_3856,N_2999,N_2698);
and U3857 (N_3857,N_2614,N_2044);
nor U3858 (N_3858,N_2457,N_2112);
nand U3859 (N_3859,N_2256,N_2852);
and U3860 (N_3860,N_2470,N_2835);
and U3861 (N_3861,N_2999,N_2012);
and U3862 (N_3862,N_2544,N_2813);
and U3863 (N_3863,N_2673,N_2914);
nand U3864 (N_3864,N_2067,N_2515);
and U3865 (N_3865,N_2227,N_2834);
xor U3866 (N_3866,N_2623,N_2347);
nand U3867 (N_3867,N_2639,N_2917);
or U3868 (N_3868,N_2147,N_2787);
xor U3869 (N_3869,N_2941,N_2890);
xor U3870 (N_3870,N_2694,N_2306);
xnor U3871 (N_3871,N_2178,N_2656);
and U3872 (N_3872,N_2100,N_2087);
or U3873 (N_3873,N_2575,N_2151);
nor U3874 (N_3874,N_2835,N_2786);
or U3875 (N_3875,N_2729,N_2755);
and U3876 (N_3876,N_2531,N_2836);
nand U3877 (N_3877,N_2707,N_2723);
and U3878 (N_3878,N_2184,N_2262);
or U3879 (N_3879,N_2830,N_2686);
or U3880 (N_3880,N_2033,N_2736);
or U3881 (N_3881,N_2244,N_2448);
nor U3882 (N_3882,N_2785,N_2804);
nand U3883 (N_3883,N_2679,N_2816);
or U3884 (N_3884,N_2239,N_2245);
and U3885 (N_3885,N_2309,N_2332);
nor U3886 (N_3886,N_2749,N_2886);
nand U3887 (N_3887,N_2892,N_2484);
or U3888 (N_3888,N_2326,N_2736);
and U3889 (N_3889,N_2258,N_2290);
nand U3890 (N_3890,N_2564,N_2408);
or U3891 (N_3891,N_2376,N_2178);
nor U3892 (N_3892,N_2745,N_2574);
xor U3893 (N_3893,N_2936,N_2197);
and U3894 (N_3894,N_2040,N_2793);
nor U3895 (N_3895,N_2217,N_2530);
nand U3896 (N_3896,N_2531,N_2162);
nor U3897 (N_3897,N_2864,N_2639);
and U3898 (N_3898,N_2666,N_2723);
and U3899 (N_3899,N_2052,N_2767);
nand U3900 (N_3900,N_2777,N_2727);
or U3901 (N_3901,N_2957,N_2260);
or U3902 (N_3902,N_2389,N_2478);
nor U3903 (N_3903,N_2454,N_2473);
or U3904 (N_3904,N_2004,N_2068);
nor U3905 (N_3905,N_2556,N_2387);
xnor U3906 (N_3906,N_2954,N_2632);
and U3907 (N_3907,N_2411,N_2218);
or U3908 (N_3908,N_2214,N_2316);
nand U3909 (N_3909,N_2427,N_2586);
xnor U3910 (N_3910,N_2212,N_2407);
nor U3911 (N_3911,N_2999,N_2924);
nand U3912 (N_3912,N_2740,N_2913);
nor U3913 (N_3913,N_2984,N_2226);
and U3914 (N_3914,N_2761,N_2127);
xor U3915 (N_3915,N_2548,N_2886);
nand U3916 (N_3916,N_2291,N_2678);
xnor U3917 (N_3917,N_2993,N_2605);
or U3918 (N_3918,N_2936,N_2919);
xor U3919 (N_3919,N_2271,N_2902);
and U3920 (N_3920,N_2465,N_2383);
xor U3921 (N_3921,N_2425,N_2688);
or U3922 (N_3922,N_2197,N_2199);
nand U3923 (N_3923,N_2989,N_2357);
xor U3924 (N_3924,N_2081,N_2393);
nand U3925 (N_3925,N_2639,N_2621);
and U3926 (N_3926,N_2492,N_2967);
or U3927 (N_3927,N_2889,N_2147);
xor U3928 (N_3928,N_2585,N_2295);
and U3929 (N_3929,N_2157,N_2469);
and U3930 (N_3930,N_2186,N_2114);
or U3931 (N_3931,N_2368,N_2479);
or U3932 (N_3932,N_2340,N_2847);
or U3933 (N_3933,N_2169,N_2495);
and U3934 (N_3934,N_2606,N_2683);
xnor U3935 (N_3935,N_2573,N_2033);
xnor U3936 (N_3936,N_2269,N_2657);
xnor U3937 (N_3937,N_2090,N_2585);
and U3938 (N_3938,N_2265,N_2561);
nand U3939 (N_3939,N_2764,N_2843);
xnor U3940 (N_3940,N_2627,N_2494);
and U3941 (N_3941,N_2206,N_2708);
xnor U3942 (N_3942,N_2337,N_2352);
or U3943 (N_3943,N_2673,N_2932);
nor U3944 (N_3944,N_2228,N_2773);
and U3945 (N_3945,N_2357,N_2129);
nor U3946 (N_3946,N_2896,N_2784);
and U3947 (N_3947,N_2161,N_2000);
nor U3948 (N_3948,N_2414,N_2993);
xor U3949 (N_3949,N_2493,N_2721);
and U3950 (N_3950,N_2165,N_2595);
or U3951 (N_3951,N_2002,N_2299);
or U3952 (N_3952,N_2140,N_2428);
and U3953 (N_3953,N_2170,N_2321);
or U3954 (N_3954,N_2742,N_2889);
nor U3955 (N_3955,N_2148,N_2036);
and U3956 (N_3956,N_2281,N_2202);
xor U3957 (N_3957,N_2780,N_2535);
nand U3958 (N_3958,N_2454,N_2525);
nor U3959 (N_3959,N_2081,N_2621);
xnor U3960 (N_3960,N_2074,N_2639);
or U3961 (N_3961,N_2351,N_2234);
or U3962 (N_3962,N_2724,N_2125);
and U3963 (N_3963,N_2598,N_2589);
xor U3964 (N_3964,N_2219,N_2550);
xnor U3965 (N_3965,N_2066,N_2630);
or U3966 (N_3966,N_2276,N_2609);
nor U3967 (N_3967,N_2622,N_2087);
nand U3968 (N_3968,N_2107,N_2385);
nor U3969 (N_3969,N_2363,N_2023);
or U3970 (N_3970,N_2440,N_2366);
nor U3971 (N_3971,N_2951,N_2548);
and U3972 (N_3972,N_2751,N_2981);
or U3973 (N_3973,N_2913,N_2577);
nand U3974 (N_3974,N_2744,N_2524);
xor U3975 (N_3975,N_2140,N_2698);
nor U3976 (N_3976,N_2603,N_2920);
or U3977 (N_3977,N_2257,N_2011);
and U3978 (N_3978,N_2474,N_2196);
nor U3979 (N_3979,N_2843,N_2716);
or U3980 (N_3980,N_2661,N_2540);
and U3981 (N_3981,N_2189,N_2906);
xnor U3982 (N_3982,N_2143,N_2463);
and U3983 (N_3983,N_2923,N_2076);
nor U3984 (N_3984,N_2957,N_2375);
xnor U3985 (N_3985,N_2161,N_2272);
nor U3986 (N_3986,N_2210,N_2995);
nor U3987 (N_3987,N_2722,N_2325);
nor U3988 (N_3988,N_2151,N_2073);
or U3989 (N_3989,N_2354,N_2148);
or U3990 (N_3990,N_2844,N_2300);
and U3991 (N_3991,N_2380,N_2807);
xnor U3992 (N_3992,N_2627,N_2587);
nor U3993 (N_3993,N_2601,N_2472);
xnor U3994 (N_3994,N_2251,N_2132);
nand U3995 (N_3995,N_2080,N_2433);
or U3996 (N_3996,N_2661,N_2352);
xor U3997 (N_3997,N_2844,N_2346);
nand U3998 (N_3998,N_2051,N_2332);
and U3999 (N_3999,N_2716,N_2861);
nor U4000 (N_4000,N_3108,N_3694);
xor U4001 (N_4001,N_3501,N_3855);
nor U4002 (N_4002,N_3093,N_3460);
nand U4003 (N_4003,N_3056,N_3813);
or U4004 (N_4004,N_3780,N_3662);
nand U4005 (N_4005,N_3628,N_3533);
nor U4006 (N_4006,N_3920,N_3812);
nor U4007 (N_4007,N_3912,N_3410);
nand U4008 (N_4008,N_3206,N_3217);
and U4009 (N_4009,N_3610,N_3753);
nor U4010 (N_4010,N_3637,N_3591);
and U4011 (N_4011,N_3403,N_3671);
nand U4012 (N_4012,N_3595,N_3751);
xor U4013 (N_4013,N_3193,N_3394);
nor U4014 (N_4014,N_3650,N_3622);
and U4015 (N_4015,N_3534,N_3292);
xnor U4016 (N_4016,N_3042,N_3086);
nor U4017 (N_4017,N_3377,N_3679);
nor U4018 (N_4018,N_3287,N_3604);
or U4019 (N_4019,N_3562,N_3878);
xor U4020 (N_4020,N_3357,N_3575);
xnor U4021 (N_4021,N_3366,N_3259);
xnor U4022 (N_4022,N_3865,N_3379);
nor U4023 (N_4023,N_3049,N_3654);
and U4024 (N_4024,N_3787,N_3888);
nand U4025 (N_4025,N_3022,N_3491);
and U4026 (N_4026,N_3640,N_3487);
nor U4027 (N_4027,N_3015,N_3757);
xor U4028 (N_4028,N_3051,N_3105);
nand U4029 (N_4029,N_3556,N_3370);
or U4030 (N_4030,N_3153,N_3758);
or U4031 (N_4031,N_3311,N_3331);
nand U4032 (N_4032,N_3378,N_3882);
or U4033 (N_4033,N_3162,N_3172);
nand U4034 (N_4034,N_3146,N_3877);
nand U4035 (N_4035,N_3045,N_3012);
nand U4036 (N_4036,N_3037,N_3858);
nor U4037 (N_4037,N_3148,N_3618);
xor U4038 (N_4038,N_3356,N_3034);
or U4039 (N_4039,N_3171,N_3299);
or U4040 (N_4040,N_3922,N_3669);
nand U4041 (N_4041,N_3164,N_3623);
and U4042 (N_4042,N_3973,N_3434);
and U4043 (N_4043,N_3512,N_3866);
and U4044 (N_4044,N_3317,N_3999);
or U4045 (N_4045,N_3754,N_3004);
nor U4046 (N_4046,N_3278,N_3030);
nor U4047 (N_4047,N_3002,N_3509);
nand U4048 (N_4048,N_3833,N_3660);
and U4049 (N_4049,N_3426,N_3756);
or U4050 (N_4050,N_3282,N_3231);
and U4051 (N_4051,N_3074,N_3306);
and U4052 (N_4052,N_3747,N_3627);
xor U4053 (N_4053,N_3392,N_3427);
and U4054 (N_4054,N_3061,N_3048);
or U4055 (N_4055,N_3670,N_3547);
and U4056 (N_4056,N_3233,N_3986);
nor U4057 (N_4057,N_3507,N_3988);
xor U4058 (N_4058,N_3302,N_3658);
nor U4059 (N_4059,N_3177,N_3797);
nor U4060 (N_4060,N_3943,N_3273);
nand U4061 (N_4061,N_3429,N_3358);
or U4062 (N_4062,N_3836,N_3350);
nor U4063 (N_4063,N_3175,N_3774);
or U4064 (N_4064,N_3652,N_3038);
or U4065 (N_4065,N_3886,N_3214);
and U4066 (N_4066,N_3527,N_3284);
nand U4067 (N_4067,N_3021,N_3188);
nand U4068 (N_4068,N_3016,N_3160);
and U4069 (N_4069,N_3708,N_3229);
or U4070 (N_4070,N_3389,N_3340);
or U4071 (N_4071,N_3723,N_3421);
and U4072 (N_4072,N_3211,N_3228);
nand U4073 (N_4073,N_3207,N_3482);
or U4074 (N_4074,N_3448,N_3535);
xnor U4075 (N_4075,N_3847,N_3589);
xor U4076 (N_4076,N_3123,N_3449);
and U4077 (N_4077,N_3614,N_3314);
xor U4078 (N_4078,N_3274,N_3083);
nand U4079 (N_4079,N_3245,N_3498);
and U4080 (N_4080,N_3633,N_3140);
and U4081 (N_4081,N_3731,N_3312);
nor U4082 (N_4082,N_3839,N_3446);
or U4083 (N_4083,N_3985,N_3892);
xor U4084 (N_4084,N_3133,N_3323);
xor U4085 (N_4085,N_3997,N_3316);
nor U4086 (N_4086,N_3280,N_3683);
nor U4087 (N_4087,N_3542,N_3066);
or U4088 (N_4088,N_3386,N_3064);
nand U4089 (N_4089,N_3802,N_3435);
nor U4090 (N_4090,N_3856,N_3724);
nor U4091 (N_4091,N_3383,N_3117);
or U4092 (N_4092,N_3649,N_3818);
or U4093 (N_4093,N_3032,N_3529);
and U4094 (N_4094,N_3848,N_3684);
xnor U4095 (N_4095,N_3772,N_3979);
xnor U4096 (N_4096,N_3354,N_3289);
or U4097 (N_4097,N_3700,N_3104);
and U4098 (N_4098,N_3578,N_3178);
nor U4099 (N_4099,N_3009,N_3863);
nand U4100 (N_4100,N_3442,N_3933);
nor U4101 (N_4101,N_3272,N_3809);
and U4102 (N_4102,N_3906,N_3225);
xor U4103 (N_4103,N_3510,N_3664);
nand U4104 (N_4104,N_3202,N_3293);
nand U4105 (N_4105,N_3439,N_3007);
and U4106 (N_4106,N_3805,N_3408);
nor U4107 (N_4107,N_3275,N_3308);
and U4108 (N_4108,N_3918,N_3931);
and U4109 (N_4109,N_3381,N_3976);
and U4110 (N_4110,N_3062,N_3196);
or U4111 (N_4111,N_3174,N_3387);
or U4112 (N_4112,N_3041,N_3619);
nand U4113 (N_4113,N_3859,N_3644);
or U4114 (N_4114,N_3363,N_3224);
or U4115 (N_4115,N_3817,N_3852);
and U4116 (N_4116,N_3279,N_3755);
xnor U4117 (N_4117,N_3219,N_3617);
and U4118 (N_4118,N_3063,N_3554);
xnor U4119 (N_4119,N_3666,N_3341);
xor U4120 (N_4120,N_3629,N_3096);
and U4121 (N_4121,N_3409,N_3053);
or U4122 (N_4122,N_3201,N_3348);
nor U4123 (N_4123,N_3549,N_3396);
or U4124 (N_4124,N_3620,N_3268);
nor U4125 (N_4125,N_3538,N_3420);
nand U4126 (N_4126,N_3098,N_3422);
and U4127 (N_4127,N_3028,N_3101);
nor U4128 (N_4128,N_3067,N_3154);
or U4129 (N_4129,N_3929,N_3398);
xor U4130 (N_4130,N_3630,N_3641);
nand U4131 (N_4131,N_3825,N_3784);
xnor U4132 (N_4132,N_3965,N_3087);
or U4133 (N_4133,N_3406,N_3827);
nand U4134 (N_4134,N_3415,N_3967);
nor U4135 (N_4135,N_3466,N_3186);
nand U4136 (N_4136,N_3657,N_3078);
nand U4137 (N_4137,N_3260,N_3786);
and U4138 (N_4138,N_3710,N_3467);
nor U4139 (N_4139,N_3646,N_3743);
nand U4140 (N_4140,N_3477,N_3371);
xor U4141 (N_4141,N_3709,N_3514);
nor U4142 (N_4142,N_3001,N_3438);
nor U4143 (N_4143,N_3904,N_3185);
nand U4144 (N_4144,N_3076,N_3795);
xor U4145 (N_4145,N_3800,N_3347);
xnor U4146 (N_4146,N_3271,N_3842);
or U4147 (N_4147,N_3879,N_3187);
and U4148 (N_4148,N_3740,N_3447);
nand U4149 (N_4149,N_3638,N_3073);
nand U4150 (N_4150,N_3494,N_3111);
or U4151 (N_4151,N_3632,N_3414);
xor U4152 (N_4152,N_3497,N_3254);
xnor U4153 (N_4153,N_3601,N_3876);
nand U4154 (N_4154,N_3526,N_3496);
and U4155 (N_4155,N_3677,N_3785);
nand U4156 (N_4156,N_3959,N_3136);
or U4157 (N_4157,N_3499,N_3080);
nand U4158 (N_4158,N_3465,N_3916);
and U4159 (N_4159,N_3360,N_3635);
and U4160 (N_4160,N_3712,N_3995);
nand U4161 (N_4161,N_3424,N_3144);
xor U4162 (N_4162,N_3897,N_3303);
xnor U4163 (N_4163,N_3744,N_3141);
nand U4164 (N_4164,N_3810,N_3791);
nor U4165 (N_4165,N_3163,N_3269);
nor U4166 (N_4166,N_3513,N_3701);
nor U4167 (N_4167,N_3645,N_3900);
or U4168 (N_4168,N_3052,N_3546);
xor U4169 (N_4169,N_3721,N_3972);
and U4170 (N_4170,N_3213,N_3147);
and U4171 (N_4171,N_3905,N_3811);
or U4172 (N_4172,N_3692,N_3412);
or U4173 (N_4173,N_3031,N_3992);
and U4174 (N_4174,N_3796,N_3395);
and U4175 (N_4175,N_3486,N_3806);
xor U4176 (N_4176,N_3966,N_3816);
nand U4177 (N_4177,N_3521,N_3661);
xnor U4178 (N_4178,N_3713,N_3763);
xor U4179 (N_4179,N_3215,N_3720);
nor U4180 (N_4180,N_3871,N_3019);
or U4181 (N_4181,N_3516,N_3330);
or U4182 (N_4182,N_3814,N_3932);
nor U4183 (N_4183,N_3776,N_3176);
or U4184 (N_4184,N_3565,N_3574);
nor U4185 (N_4185,N_3699,N_3653);
nor U4186 (N_4186,N_3599,N_3373);
nor U4187 (N_4187,N_3896,N_3968);
or U4188 (N_4188,N_3334,N_3958);
nor U4189 (N_4189,N_3735,N_3327);
nor U4190 (N_4190,N_3286,N_3949);
or U4191 (N_4191,N_3970,N_3010);
nor U4192 (N_4192,N_3425,N_3975);
xnor U4193 (N_4193,N_3479,N_3613);
or U4194 (N_4194,N_3831,N_3138);
nor U4195 (N_4195,N_3539,N_3401);
or U4196 (N_4196,N_3634,N_3707);
and U4197 (N_4197,N_3075,N_3911);
nand U4198 (N_4198,N_3752,N_3790);
or U4199 (N_4199,N_3974,N_3393);
nand U4200 (N_4200,N_3902,N_3663);
or U4201 (N_4201,N_3026,N_3440);
and U4202 (N_4202,N_3167,N_3265);
nand U4203 (N_4203,N_3946,N_3359);
and U4204 (N_4204,N_3291,N_3263);
and U4205 (N_4205,N_3184,N_3113);
xor U4206 (N_4206,N_3977,N_3616);
nor U4207 (N_4207,N_3005,N_3500);
nand U4208 (N_4208,N_3470,N_3696);
xor U4209 (N_4209,N_3339,N_3255);
xnor U4210 (N_4210,N_3605,N_3698);
nor U4211 (N_4211,N_3018,N_3251);
and U4212 (N_4212,N_3901,N_3475);
xor U4213 (N_4213,N_3261,N_3917);
nor U4214 (N_4214,N_3055,N_3264);
and U4215 (N_4215,N_3304,N_3192);
nand U4216 (N_4216,N_3557,N_3262);
and U4217 (N_4217,N_3913,N_3947);
and U4218 (N_4218,N_3782,N_3281);
nand U4219 (N_4219,N_3384,N_3132);
xor U4220 (N_4220,N_3603,N_3155);
nor U4221 (N_4221,N_3563,N_3365);
or U4222 (N_4222,N_3399,N_3194);
and U4223 (N_4223,N_3687,N_3071);
and U4224 (N_4224,N_3189,N_3530);
or U4225 (N_4225,N_3079,N_3585);
or U4226 (N_4226,N_3006,N_3511);
nand U4227 (N_4227,N_3523,N_3860);
and U4228 (N_4228,N_3870,N_3220);
nor U4229 (N_4229,N_3114,N_3702);
xnor U4230 (N_4230,N_3173,N_3586);
nand U4231 (N_4231,N_3550,N_3191);
nand U4232 (N_4232,N_3775,N_3333);
and U4233 (N_4233,N_3161,N_3919);
nand U4234 (N_4234,N_3077,N_3602);
and U4235 (N_4235,N_3741,N_3119);
and U4236 (N_4236,N_3808,N_3573);
or U4237 (N_4237,N_3584,N_3714);
and U4238 (N_4238,N_3715,N_3989);
xnor U4239 (N_4239,N_3954,N_3216);
nand U4240 (N_4240,N_3835,N_3935);
or U4241 (N_4241,N_3070,N_3013);
nand U4242 (N_4242,N_3490,N_3792);
nor U4243 (N_4243,N_3941,N_3374);
xnor U4244 (N_4244,N_3828,N_3205);
xnor U4245 (N_4245,N_3506,N_3115);
xnor U4246 (N_4246,N_3168,N_3971);
nor U4247 (N_4247,N_3643,N_3054);
nor U4248 (N_4248,N_3993,N_3481);
nor U4249 (N_4249,N_3517,N_3588);
nand U4250 (N_4250,N_3221,N_3571);
or U4251 (N_4251,N_3801,N_3624);
nor U4252 (N_4252,N_3493,N_3914);
nand U4253 (N_4253,N_3469,N_3139);
xor U4254 (N_4254,N_3594,N_3937);
or U4255 (N_4255,N_3346,N_3771);
nor U4256 (N_4256,N_3718,N_3572);
nor U4257 (N_4257,N_3407,N_3452);
xnor U4258 (N_4258,N_3459,N_3208);
nand U4259 (N_4259,N_3738,N_3222);
and U4260 (N_4260,N_3344,N_3597);
nor U4261 (N_4261,N_3058,N_3727);
nand U4262 (N_4262,N_3829,N_3120);
and U4263 (N_4263,N_3088,N_3711);
nand U4264 (N_4264,N_3717,N_3248);
xnor U4265 (N_4265,N_3226,N_3823);
nor U4266 (N_4266,N_3300,N_3890);
xnor U4267 (N_4267,N_3545,N_3118);
or U4268 (N_4268,N_3925,N_3256);
xor U4269 (N_4269,N_3781,N_3861);
xnor U4270 (N_4270,N_3250,N_3242);
nand U4271 (N_4271,N_3561,N_3124);
or U4272 (N_4272,N_3068,N_3143);
and U4273 (N_4273,N_3478,N_3209);
nand U4274 (N_4274,N_3899,N_3129);
or U4275 (N_4275,N_3704,N_3235);
nand U4276 (N_4276,N_3152,N_3779);
xor U4277 (N_4277,N_3642,N_3474);
or U4278 (N_4278,N_3874,N_3742);
or U4279 (N_4279,N_3458,N_3036);
or U4280 (N_4280,N_3020,N_3868);
xnor U4281 (N_4281,N_3765,N_3569);
nand U4282 (N_4282,N_3468,N_3000);
xor U4283 (N_4283,N_3655,N_3889);
nand U4284 (N_4284,N_3609,N_3705);
or U4285 (N_4285,N_3277,N_3921);
xor U4286 (N_4286,N_3598,N_3955);
xor U4287 (N_4287,N_3008,N_3390);
or U4288 (N_4288,N_3587,N_3212);
and U4289 (N_4289,N_3957,N_3436);
nand U4290 (N_4290,N_3544,N_3450);
or U4291 (N_4291,N_3247,N_3950);
nand U4292 (N_4292,N_3626,N_3532);
or U4293 (N_4293,N_3046,N_3841);
or U4294 (N_4294,N_3788,N_3252);
nand U4295 (N_4295,N_3908,N_3157);
xor U4296 (N_4296,N_3431,N_3887);
nor U4297 (N_4297,N_3417,N_3762);
and U4298 (N_4298,N_3543,N_3290);
xnor U4299 (N_4299,N_3749,N_3745);
and U4300 (N_4300,N_3990,N_3336);
nor U4301 (N_4301,N_3319,N_3996);
nand U4302 (N_4302,N_3199,N_3433);
xnor U4303 (N_4303,N_3862,N_3822);
nand U4304 (N_4304,N_3726,N_3159);
and U4305 (N_4305,N_3195,N_3730);
and U4306 (N_4306,N_3349,N_3611);
or U4307 (N_4307,N_3940,N_3703);
or U4308 (N_4308,N_3737,N_3555);
or U4309 (N_4309,N_3551,N_3190);
or U4310 (N_4310,N_3137,N_3276);
xnor U4311 (N_4311,N_3566,N_3150);
nand U4312 (N_4312,N_3799,N_3069);
xor U4313 (N_4313,N_3930,N_3678);
or U4314 (N_4314,N_3991,N_3179);
xor U4315 (N_4315,N_3027,N_3983);
xor U4316 (N_4316,N_3218,N_3361);
nor U4317 (N_4317,N_3368,N_3576);
nor U4318 (N_4318,N_3608,N_3335);
or U4319 (N_4319,N_3091,N_3739);
or U4320 (N_4320,N_3044,N_3085);
xor U4321 (N_4321,N_3722,N_3345);
and U4322 (N_4322,N_3103,N_3040);
nand U4323 (N_4323,N_3230,N_3454);
nand U4324 (N_4324,N_3909,N_3948);
or U4325 (N_4325,N_3382,N_3102);
nand U4326 (N_4326,N_3736,N_3553);
and U4327 (N_4327,N_3668,N_3488);
nand U4328 (N_4328,N_3364,N_3156);
or U4329 (N_4329,N_3234,N_3732);
or U4330 (N_4330,N_3107,N_3047);
nor U4331 (N_4331,N_3244,N_3112);
or U4332 (N_4332,N_3307,N_3166);
or U4333 (N_4333,N_3158,N_3821);
and U4334 (N_4334,N_3794,N_3980);
xor U4335 (N_4335,N_3489,N_3203);
or U4336 (N_4336,N_3528,N_3180);
nand U4337 (N_4337,N_3391,N_3938);
nand U4338 (N_4338,N_3223,N_3548);
or U4339 (N_4339,N_3778,N_3524);
nor U4340 (N_4340,N_3734,N_3116);
nand U4341 (N_4341,N_3332,N_3135);
nor U4342 (N_4342,N_3964,N_3639);
and U4343 (N_4343,N_3615,N_3880);
and U4344 (N_4344,N_3819,N_3039);
nand U4345 (N_4345,N_3232,N_3035);
nand U4346 (N_4346,N_3301,N_3266);
xnor U4347 (N_4347,N_3537,N_3324);
and U4348 (N_4348,N_3981,N_3681);
nor U4349 (N_4349,N_3552,N_3325);
nor U4350 (N_4350,N_3200,N_3559);
nand U4351 (N_4351,N_3456,N_3854);
xnor U4352 (N_4352,N_3881,N_3636);
nor U4353 (N_4353,N_3437,N_3680);
nor U4354 (N_4354,N_3525,N_3834);
and U4355 (N_4355,N_3952,N_3750);
and U4356 (N_4356,N_3607,N_3893);
or U4357 (N_4357,N_3285,N_3376);
and U4358 (N_4358,N_3313,N_3830);
nor U4359 (N_4359,N_3181,N_3928);
xor U4360 (N_4360,N_3891,N_3170);
and U4361 (N_4361,N_3518,N_3564);
nand U4362 (N_4362,N_3612,N_3142);
nand U4363 (N_4363,N_3850,N_3237);
xnor U4364 (N_4364,N_3998,N_3025);
nand U4365 (N_4365,N_3693,N_3227);
nor U4366 (N_4366,N_3318,N_3322);
nand U4367 (N_4367,N_3789,N_3939);
or U4368 (N_4368,N_3283,N_3631);
nand U4369 (N_4369,N_3471,N_3826);
and U4370 (N_4370,N_3926,N_3923);
or U4371 (N_4371,N_3131,N_3577);
and U4372 (N_4372,N_3725,N_3023);
nand U4373 (N_4373,N_3298,N_3984);
xnor U4374 (N_4374,N_3793,N_3804);
xor U4375 (N_4375,N_3461,N_3445);
xor U4376 (N_4376,N_3296,N_3873);
nor U4377 (N_4377,N_3502,N_3648);
nor U4378 (N_4378,N_3903,N_3457);
nand U4379 (N_4379,N_3149,N_3803);
and U4380 (N_4380,N_3894,N_3978);
xor U4381 (N_4381,N_3110,N_3090);
nand U4382 (N_4382,N_3536,N_3695);
nor U4383 (N_4383,N_3570,N_3483);
nor U4384 (N_4384,N_3329,N_3197);
xnor U4385 (N_4385,N_3851,N_3883);
nand U4386 (N_4386,N_3128,N_3484);
or U4387 (N_4387,N_3432,N_3081);
xnor U4388 (N_4388,N_3682,N_3443);
or U4389 (N_4389,N_3253,N_3838);
and U4390 (N_4390,N_3647,N_3092);
and U4391 (N_4391,N_3568,N_3961);
nand U4392 (N_4392,N_3485,N_3441);
xor U4393 (N_4393,N_3685,N_3369);
and U4394 (N_4394,N_3910,N_3134);
nor U4395 (N_4395,N_3151,N_3656);
and U4396 (N_4396,N_3690,N_3849);
nor U4397 (N_4397,N_3689,N_3853);
nand U4398 (N_4398,N_3728,N_3582);
and U4399 (N_4399,N_3515,N_3082);
nand U4400 (N_4400,N_3473,N_3326);
nor U4401 (N_4401,N_3321,N_3464);
nor U4402 (N_4402,N_3182,N_3686);
nand U4403 (N_4403,N_3867,N_3342);
or U4404 (N_4404,N_3519,N_3934);
and U4405 (N_4405,N_3258,N_3915);
and U4406 (N_4406,N_3592,N_3352);
and U4407 (N_4407,N_3017,N_3210);
nand U4408 (N_4408,N_3444,N_3746);
and U4409 (N_4409,N_3011,N_3305);
and U4410 (N_4410,N_3807,N_3820);
xor U4411 (N_4411,N_3982,N_3463);
nor U4412 (N_4412,N_3541,N_3243);
nor U4413 (N_4413,N_3504,N_3845);
nor U4414 (N_4414,N_3885,N_3675);
and U4415 (N_4415,N_3315,N_3249);
nor U4416 (N_4416,N_3770,N_3560);
and U4417 (N_4417,N_3697,N_3783);
xor U4418 (N_4418,N_3625,N_3462);
nand U4419 (N_4419,N_3130,N_3204);
xor U4420 (N_4420,N_3288,N_3404);
and U4421 (N_4421,N_3580,N_3430);
xor U4422 (N_4422,N_3798,N_3169);
and U4423 (N_4423,N_3418,N_3773);
nor U4424 (N_4424,N_3667,N_3372);
and U4425 (N_4425,N_3651,N_3531);
and U4426 (N_4426,N_3583,N_3413);
nor U4427 (N_4427,N_3428,N_3869);
and U4428 (N_4428,N_3072,N_3385);
nand U4429 (N_4429,N_3942,N_3065);
or U4430 (N_4430,N_3472,N_3127);
and U4431 (N_4431,N_3884,N_3691);
nor U4432 (N_4432,N_3864,N_3050);
xnor U4433 (N_4433,N_3857,N_3522);
xnor U4434 (N_4434,N_3099,N_3380);
or U4435 (N_4435,N_3846,N_3665);
and U4436 (N_4436,N_3719,N_3875);
and U4437 (N_4437,N_3238,N_3060);
nand U4438 (N_4438,N_3520,N_3402);
nor U4439 (N_4439,N_3672,N_3767);
nor U4440 (N_4440,N_3844,N_3239);
nor U4441 (N_4441,N_3907,N_3236);
xnor U4442 (N_4442,N_3343,N_3014);
and U4443 (N_4443,N_3729,N_3351);
nor U4444 (N_4444,N_3963,N_3590);
nor U4445 (N_4445,N_3411,N_3927);
nand U4446 (N_4446,N_3621,N_3503);
and U4447 (N_4447,N_3320,N_3059);
xnor U4448 (N_4448,N_3097,N_3145);
xor U4449 (N_4449,N_3688,N_3768);
xor U4450 (N_4450,N_3453,N_3766);
xor U4451 (N_4451,N_3924,N_3898);
nor U4452 (N_4452,N_3843,N_3126);
nor U4453 (N_4453,N_3043,N_3270);
xor U4454 (N_4454,N_3673,N_3125);
or U4455 (N_4455,N_3960,N_3581);
nor U4456 (N_4456,N_3183,N_3777);
and U4457 (N_4457,N_3944,N_3659);
and U4458 (N_4458,N_3338,N_3540);
nand U4459 (N_4459,N_3257,N_3375);
nand U4460 (N_4460,N_3337,N_3423);
nor U4461 (N_4461,N_3769,N_3815);
nand U4462 (N_4462,N_3676,N_3109);
nand U4463 (N_4463,N_3951,N_3451);
and U4464 (N_4464,N_3600,N_3953);
nor U4465 (N_4465,N_3733,N_3241);
xor U4466 (N_4466,N_3716,N_3084);
xor U4467 (N_4467,N_3095,N_3759);
and U4468 (N_4468,N_3106,N_3033);
and U4469 (N_4469,N_3760,N_3416);
or U4470 (N_4470,N_3198,N_3495);
nand U4471 (N_4471,N_3872,N_3094);
and U4472 (N_4472,N_3367,N_3400);
or U4473 (N_4473,N_3579,N_3328);
nor U4474 (N_4474,N_3505,N_3962);
or U4475 (N_4475,N_3294,N_3246);
nand U4476 (N_4476,N_3362,N_3748);
xor U4477 (N_4477,N_3057,N_3558);
and U4478 (N_4478,N_3764,N_3003);
nor U4479 (N_4479,N_3353,N_3405);
and U4480 (N_4480,N_3240,N_3100);
or U4481 (N_4481,N_3832,N_3310);
xnor U4482 (N_4482,N_3936,N_3945);
nor U4483 (N_4483,N_3355,N_3267);
and U4484 (N_4484,N_3419,N_3596);
nor U4485 (N_4485,N_3840,N_3121);
and U4486 (N_4486,N_3309,N_3706);
nor U4487 (N_4487,N_3165,N_3029);
nand U4488 (N_4488,N_3508,N_3593);
nor U4489 (N_4489,N_3492,N_3761);
nand U4490 (N_4490,N_3994,N_3122);
or U4491 (N_4491,N_3388,N_3956);
and U4492 (N_4492,N_3824,N_3606);
nor U4493 (N_4493,N_3969,N_3476);
or U4494 (N_4494,N_3089,N_3480);
and U4495 (N_4495,N_3674,N_3455);
nand U4496 (N_4496,N_3567,N_3295);
nor U4497 (N_4497,N_3837,N_3024);
or U4498 (N_4498,N_3895,N_3397);
nand U4499 (N_4499,N_3297,N_3987);
or U4500 (N_4500,N_3859,N_3935);
and U4501 (N_4501,N_3712,N_3278);
and U4502 (N_4502,N_3829,N_3557);
or U4503 (N_4503,N_3750,N_3916);
or U4504 (N_4504,N_3762,N_3437);
and U4505 (N_4505,N_3558,N_3314);
xor U4506 (N_4506,N_3517,N_3539);
nor U4507 (N_4507,N_3056,N_3224);
nand U4508 (N_4508,N_3091,N_3883);
and U4509 (N_4509,N_3621,N_3081);
and U4510 (N_4510,N_3640,N_3358);
nor U4511 (N_4511,N_3416,N_3354);
nand U4512 (N_4512,N_3565,N_3088);
and U4513 (N_4513,N_3452,N_3619);
nand U4514 (N_4514,N_3083,N_3258);
xnor U4515 (N_4515,N_3075,N_3835);
or U4516 (N_4516,N_3507,N_3471);
or U4517 (N_4517,N_3222,N_3113);
xnor U4518 (N_4518,N_3708,N_3839);
and U4519 (N_4519,N_3164,N_3707);
xnor U4520 (N_4520,N_3263,N_3839);
or U4521 (N_4521,N_3379,N_3099);
nand U4522 (N_4522,N_3288,N_3959);
nor U4523 (N_4523,N_3999,N_3158);
or U4524 (N_4524,N_3008,N_3161);
xnor U4525 (N_4525,N_3900,N_3971);
and U4526 (N_4526,N_3773,N_3360);
xnor U4527 (N_4527,N_3417,N_3788);
nor U4528 (N_4528,N_3608,N_3349);
xnor U4529 (N_4529,N_3211,N_3976);
xor U4530 (N_4530,N_3426,N_3408);
nor U4531 (N_4531,N_3169,N_3830);
nand U4532 (N_4532,N_3019,N_3504);
nor U4533 (N_4533,N_3542,N_3109);
nor U4534 (N_4534,N_3825,N_3864);
nand U4535 (N_4535,N_3138,N_3952);
nand U4536 (N_4536,N_3262,N_3547);
nand U4537 (N_4537,N_3239,N_3628);
xnor U4538 (N_4538,N_3906,N_3155);
nand U4539 (N_4539,N_3794,N_3598);
and U4540 (N_4540,N_3910,N_3829);
xnor U4541 (N_4541,N_3677,N_3097);
nand U4542 (N_4542,N_3198,N_3700);
nand U4543 (N_4543,N_3782,N_3794);
xnor U4544 (N_4544,N_3538,N_3738);
and U4545 (N_4545,N_3143,N_3423);
nor U4546 (N_4546,N_3995,N_3986);
nor U4547 (N_4547,N_3727,N_3234);
and U4548 (N_4548,N_3520,N_3351);
nand U4549 (N_4549,N_3376,N_3138);
xor U4550 (N_4550,N_3885,N_3476);
nand U4551 (N_4551,N_3371,N_3431);
or U4552 (N_4552,N_3690,N_3596);
or U4553 (N_4553,N_3556,N_3844);
xor U4554 (N_4554,N_3397,N_3781);
nand U4555 (N_4555,N_3129,N_3994);
or U4556 (N_4556,N_3089,N_3066);
or U4557 (N_4557,N_3809,N_3908);
or U4558 (N_4558,N_3975,N_3564);
or U4559 (N_4559,N_3985,N_3604);
and U4560 (N_4560,N_3150,N_3171);
xor U4561 (N_4561,N_3862,N_3804);
or U4562 (N_4562,N_3634,N_3665);
or U4563 (N_4563,N_3932,N_3595);
nand U4564 (N_4564,N_3125,N_3518);
or U4565 (N_4565,N_3650,N_3781);
xor U4566 (N_4566,N_3689,N_3785);
and U4567 (N_4567,N_3435,N_3807);
nand U4568 (N_4568,N_3212,N_3288);
nor U4569 (N_4569,N_3908,N_3862);
xnor U4570 (N_4570,N_3859,N_3940);
or U4571 (N_4571,N_3499,N_3064);
or U4572 (N_4572,N_3668,N_3148);
nor U4573 (N_4573,N_3280,N_3586);
nor U4574 (N_4574,N_3336,N_3070);
nor U4575 (N_4575,N_3404,N_3717);
or U4576 (N_4576,N_3318,N_3374);
and U4577 (N_4577,N_3609,N_3787);
nor U4578 (N_4578,N_3657,N_3714);
nor U4579 (N_4579,N_3787,N_3386);
xnor U4580 (N_4580,N_3712,N_3392);
nand U4581 (N_4581,N_3892,N_3553);
xor U4582 (N_4582,N_3730,N_3137);
and U4583 (N_4583,N_3960,N_3692);
nand U4584 (N_4584,N_3962,N_3543);
nand U4585 (N_4585,N_3685,N_3752);
nand U4586 (N_4586,N_3055,N_3132);
and U4587 (N_4587,N_3943,N_3652);
nor U4588 (N_4588,N_3402,N_3374);
xor U4589 (N_4589,N_3346,N_3937);
xor U4590 (N_4590,N_3753,N_3097);
or U4591 (N_4591,N_3022,N_3389);
nand U4592 (N_4592,N_3174,N_3508);
nor U4593 (N_4593,N_3681,N_3717);
or U4594 (N_4594,N_3060,N_3842);
nor U4595 (N_4595,N_3956,N_3128);
xor U4596 (N_4596,N_3193,N_3896);
or U4597 (N_4597,N_3764,N_3324);
and U4598 (N_4598,N_3648,N_3318);
nand U4599 (N_4599,N_3124,N_3274);
xor U4600 (N_4600,N_3805,N_3385);
nor U4601 (N_4601,N_3431,N_3645);
nand U4602 (N_4602,N_3259,N_3776);
nor U4603 (N_4603,N_3894,N_3202);
nand U4604 (N_4604,N_3853,N_3935);
and U4605 (N_4605,N_3016,N_3041);
xnor U4606 (N_4606,N_3935,N_3467);
or U4607 (N_4607,N_3163,N_3589);
xnor U4608 (N_4608,N_3198,N_3467);
and U4609 (N_4609,N_3994,N_3482);
and U4610 (N_4610,N_3319,N_3074);
nor U4611 (N_4611,N_3494,N_3722);
nand U4612 (N_4612,N_3641,N_3646);
nand U4613 (N_4613,N_3575,N_3895);
xnor U4614 (N_4614,N_3350,N_3716);
nand U4615 (N_4615,N_3257,N_3211);
nor U4616 (N_4616,N_3289,N_3819);
xor U4617 (N_4617,N_3586,N_3882);
and U4618 (N_4618,N_3852,N_3722);
nor U4619 (N_4619,N_3455,N_3540);
and U4620 (N_4620,N_3399,N_3914);
and U4621 (N_4621,N_3350,N_3949);
nor U4622 (N_4622,N_3257,N_3298);
xnor U4623 (N_4623,N_3660,N_3000);
and U4624 (N_4624,N_3535,N_3288);
xnor U4625 (N_4625,N_3859,N_3019);
and U4626 (N_4626,N_3008,N_3876);
or U4627 (N_4627,N_3371,N_3430);
nor U4628 (N_4628,N_3613,N_3684);
and U4629 (N_4629,N_3957,N_3715);
and U4630 (N_4630,N_3395,N_3834);
or U4631 (N_4631,N_3655,N_3075);
nor U4632 (N_4632,N_3496,N_3491);
or U4633 (N_4633,N_3516,N_3867);
nor U4634 (N_4634,N_3096,N_3908);
and U4635 (N_4635,N_3569,N_3135);
nor U4636 (N_4636,N_3516,N_3974);
or U4637 (N_4637,N_3134,N_3240);
xnor U4638 (N_4638,N_3773,N_3239);
and U4639 (N_4639,N_3116,N_3855);
or U4640 (N_4640,N_3379,N_3074);
or U4641 (N_4641,N_3063,N_3986);
and U4642 (N_4642,N_3193,N_3842);
and U4643 (N_4643,N_3101,N_3322);
and U4644 (N_4644,N_3060,N_3190);
and U4645 (N_4645,N_3031,N_3004);
nor U4646 (N_4646,N_3855,N_3253);
xnor U4647 (N_4647,N_3200,N_3702);
and U4648 (N_4648,N_3008,N_3856);
nor U4649 (N_4649,N_3405,N_3031);
or U4650 (N_4650,N_3034,N_3606);
or U4651 (N_4651,N_3525,N_3373);
nor U4652 (N_4652,N_3168,N_3745);
and U4653 (N_4653,N_3973,N_3513);
nand U4654 (N_4654,N_3068,N_3727);
nor U4655 (N_4655,N_3450,N_3335);
nor U4656 (N_4656,N_3719,N_3880);
nand U4657 (N_4657,N_3482,N_3156);
nor U4658 (N_4658,N_3649,N_3542);
nand U4659 (N_4659,N_3640,N_3277);
nor U4660 (N_4660,N_3489,N_3323);
and U4661 (N_4661,N_3533,N_3123);
xnor U4662 (N_4662,N_3566,N_3880);
or U4663 (N_4663,N_3100,N_3550);
xnor U4664 (N_4664,N_3718,N_3008);
nand U4665 (N_4665,N_3913,N_3332);
nor U4666 (N_4666,N_3490,N_3435);
nor U4667 (N_4667,N_3741,N_3667);
or U4668 (N_4668,N_3718,N_3845);
and U4669 (N_4669,N_3457,N_3846);
xnor U4670 (N_4670,N_3106,N_3149);
xor U4671 (N_4671,N_3344,N_3654);
xor U4672 (N_4672,N_3444,N_3555);
nor U4673 (N_4673,N_3318,N_3436);
nor U4674 (N_4674,N_3139,N_3417);
and U4675 (N_4675,N_3536,N_3385);
xnor U4676 (N_4676,N_3291,N_3127);
and U4677 (N_4677,N_3814,N_3188);
xnor U4678 (N_4678,N_3356,N_3803);
xnor U4679 (N_4679,N_3836,N_3302);
nor U4680 (N_4680,N_3516,N_3042);
or U4681 (N_4681,N_3180,N_3899);
nand U4682 (N_4682,N_3044,N_3822);
and U4683 (N_4683,N_3277,N_3393);
nand U4684 (N_4684,N_3188,N_3747);
or U4685 (N_4685,N_3997,N_3393);
or U4686 (N_4686,N_3502,N_3059);
xor U4687 (N_4687,N_3624,N_3802);
xnor U4688 (N_4688,N_3590,N_3131);
and U4689 (N_4689,N_3086,N_3309);
nor U4690 (N_4690,N_3642,N_3291);
nor U4691 (N_4691,N_3902,N_3343);
or U4692 (N_4692,N_3143,N_3080);
nand U4693 (N_4693,N_3909,N_3862);
or U4694 (N_4694,N_3856,N_3187);
or U4695 (N_4695,N_3832,N_3292);
or U4696 (N_4696,N_3719,N_3991);
xor U4697 (N_4697,N_3086,N_3114);
and U4698 (N_4698,N_3257,N_3333);
and U4699 (N_4699,N_3119,N_3327);
xnor U4700 (N_4700,N_3936,N_3214);
nor U4701 (N_4701,N_3034,N_3345);
xnor U4702 (N_4702,N_3684,N_3310);
and U4703 (N_4703,N_3878,N_3772);
xor U4704 (N_4704,N_3408,N_3661);
nor U4705 (N_4705,N_3994,N_3035);
or U4706 (N_4706,N_3946,N_3973);
or U4707 (N_4707,N_3845,N_3147);
nor U4708 (N_4708,N_3318,N_3813);
or U4709 (N_4709,N_3211,N_3237);
nor U4710 (N_4710,N_3628,N_3727);
and U4711 (N_4711,N_3646,N_3205);
nand U4712 (N_4712,N_3222,N_3083);
or U4713 (N_4713,N_3331,N_3870);
nor U4714 (N_4714,N_3601,N_3703);
nand U4715 (N_4715,N_3770,N_3454);
and U4716 (N_4716,N_3575,N_3137);
or U4717 (N_4717,N_3098,N_3807);
nor U4718 (N_4718,N_3252,N_3699);
and U4719 (N_4719,N_3561,N_3805);
nor U4720 (N_4720,N_3761,N_3302);
nand U4721 (N_4721,N_3238,N_3729);
xor U4722 (N_4722,N_3763,N_3352);
and U4723 (N_4723,N_3241,N_3655);
nor U4724 (N_4724,N_3427,N_3618);
nor U4725 (N_4725,N_3673,N_3014);
xor U4726 (N_4726,N_3723,N_3904);
or U4727 (N_4727,N_3659,N_3435);
nand U4728 (N_4728,N_3345,N_3462);
or U4729 (N_4729,N_3682,N_3548);
and U4730 (N_4730,N_3011,N_3633);
and U4731 (N_4731,N_3322,N_3821);
and U4732 (N_4732,N_3442,N_3849);
nand U4733 (N_4733,N_3078,N_3496);
and U4734 (N_4734,N_3906,N_3437);
and U4735 (N_4735,N_3812,N_3217);
xnor U4736 (N_4736,N_3442,N_3172);
nor U4737 (N_4737,N_3548,N_3779);
xor U4738 (N_4738,N_3181,N_3579);
nand U4739 (N_4739,N_3115,N_3250);
nand U4740 (N_4740,N_3766,N_3187);
or U4741 (N_4741,N_3567,N_3900);
or U4742 (N_4742,N_3921,N_3292);
and U4743 (N_4743,N_3805,N_3982);
xor U4744 (N_4744,N_3015,N_3297);
nand U4745 (N_4745,N_3847,N_3169);
and U4746 (N_4746,N_3443,N_3489);
xor U4747 (N_4747,N_3458,N_3347);
nand U4748 (N_4748,N_3291,N_3297);
and U4749 (N_4749,N_3183,N_3412);
nand U4750 (N_4750,N_3186,N_3862);
or U4751 (N_4751,N_3403,N_3747);
xor U4752 (N_4752,N_3415,N_3258);
xnor U4753 (N_4753,N_3954,N_3233);
nor U4754 (N_4754,N_3364,N_3110);
or U4755 (N_4755,N_3339,N_3416);
nor U4756 (N_4756,N_3373,N_3801);
xnor U4757 (N_4757,N_3324,N_3189);
nor U4758 (N_4758,N_3990,N_3621);
nor U4759 (N_4759,N_3468,N_3463);
nand U4760 (N_4760,N_3148,N_3385);
nor U4761 (N_4761,N_3131,N_3955);
or U4762 (N_4762,N_3179,N_3129);
or U4763 (N_4763,N_3395,N_3976);
xor U4764 (N_4764,N_3302,N_3196);
or U4765 (N_4765,N_3450,N_3349);
and U4766 (N_4766,N_3071,N_3532);
xnor U4767 (N_4767,N_3391,N_3825);
xnor U4768 (N_4768,N_3372,N_3544);
or U4769 (N_4769,N_3688,N_3306);
xor U4770 (N_4770,N_3437,N_3922);
or U4771 (N_4771,N_3703,N_3654);
nor U4772 (N_4772,N_3797,N_3511);
nand U4773 (N_4773,N_3996,N_3864);
and U4774 (N_4774,N_3416,N_3361);
nor U4775 (N_4775,N_3052,N_3305);
xor U4776 (N_4776,N_3517,N_3026);
xor U4777 (N_4777,N_3095,N_3297);
xnor U4778 (N_4778,N_3269,N_3828);
xnor U4779 (N_4779,N_3232,N_3515);
and U4780 (N_4780,N_3575,N_3813);
or U4781 (N_4781,N_3811,N_3437);
xor U4782 (N_4782,N_3279,N_3717);
or U4783 (N_4783,N_3092,N_3631);
and U4784 (N_4784,N_3047,N_3753);
or U4785 (N_4785,N_3440,N_3443);
and U4786 (N_4786,N_3822,N_3801);
nand U4787 (N_4787,N_3319,N_3894);
nand U4788 (N_4788,N_3802,N_3895);
or U4789 (N_4789,N_3148,N_3124);
nor U4790 (N_4790,N_3652,N_3317);
nand U4791 (N_4791,N_3945,N_3439);
and U4792 (N_4792,N_3583,N_3079);
nand U4793 (N_4793,N_3946,N_3075);
and U4794 (N_4794,N_3127,N_3263);
and U4795 (N_4795,N_3850,N_3408);
nor U4796 (N_4796,N_3779,N_3627);
nor U4797 (N_4797,N_3618,N_3084);
nand U4798 (N_4798,N_3266,N_3752);
xnor U4799 (N_4799,N_3863,N_3986);
and U4800 (N_4800,N_3230,N_3895);
nand U4801 (N_4801,N_3096,N_3776);
or U4802 (N_4802,N_3615,N_3398);
xor U4803 (N_4803,N_3498,N_3198);
and U4804 (N_4804,N_3298,N_3003);
or U4805 (N_4805,N_3797,N_3317);
nand U4806 (N_4806,N_3737,N_3062);
nor U4807 (N_4807,N_3517,N_3357);
nand U4808 (N_4808,N_3265,N_3852);
xnor U4809 (N_4809,N_3600,N_3386);
and U4810 (N_4810,N_3134,N_3964);
or U4811 (N_4811,N_3475,N_3626);
xnor U4812 (N_4812,N_3169,N_3875);
nand U4813 (N_4813,N_3004,N_3118);
nand U4814 (N_4814,N_3339,N_3061);
nand U4815 (N_4815,N_3407,N_3757);
nand U4816 (N_4816,N_3930,N_3843);
nor U4817 (N_4817,N_3503,N_3252);
or U4818 (N_4818,N_3989,N_3223);
xor U4819 (N_4819,N_3225,N_3681);
nor U4820 (N_4820,N_3407,N_3345);
or U4821 (N_4821,N_3117,N_3269);
nand U4822 (N_4822,N_3952,N_3022);
xnor U4823 (N_4823,N_3221,N_3000);
nor U4824 (N_4824,N_3361,N_3086);
nand U4825 (N_4825,N_3112,N_3062);
nor U4826 (N_4826,N_3464,N_3809);
or U4827 (N_4827,N_3536,N_3935);
and U4828 (N_4828,N_3033,N_3946);
nand U4829 (N_4829,N_3202,N_3612);
xnor U4830 (N_4830,N_3809,N_3084);
or U4831 (N_4831,N_3713,N_3196);
nand U4832 (N_4832,N_3332,N_3578);
and U4833 (N_4833,N_3507,N_3572);
nand U4834 (N_4834,N_3872,N_3090);
nand U4835 (N_4835,N_3244,N_3606);
nor U4836 (N_4836,N_3676,N_3001);
and U4837 (N_4837,N_3232,N_3973);
nor U4838 (N_4838,N_3935,N_3772);
nor U4839 (N_4839,N_3231,N_3827);
or U4840 (N_4840,N_3158,N_3638);
nor U4841 (N_4841,N_3454,N_3289);
nor U4842 (N_4842,N_3315,N_3790);
xor U4843 (N_4843,N_3994,N_3897);
and U4844 (N_4844,N_3901,N_3734);
nand U4845 (N_4845,N_3774,N_3936);
and U4846 (N_4846,N_3433,N_3924);
xor U4847 (N_4847,N_3141,N_3580);
nand U4848 (N_4848,N_3567,N_3229);
or U4849 (N_4849,N_3512,N_3802);
and U4850 (N_4850,N_3884,N_3666);
or U4851 (N_4851,N_3539,N_3174);
or U4852 (N_4852,N_3269,N_3835);
or U4853 (N_4853,N_3361,N_3060);
and U4854 (N_4854,N_3223,N_3263);
xnor U4855 (N_4855,N_3870,N_3979);
and U4856 (N_4856,N_3598,N_3072);
xor U4857 (N_4857,N_3328,N_3524);
nand U4858 (N_4858,N_3960,N_3945);
or U4859 (N_4859,N_3407,N_3546);
or U4860 (N_4860,N_3045,N_3092);
xnor U4861 (N_4861,N_3611,N_3571);
nor U4862 (N_4862,N_3127,N_3881);
nand U4863 (N_4863,N_3818,N_3127);
xnor U4864 (N_4864,N_3780,N_3618);
nand U4865 (N_4865,N_3539,N_3614);
nor U4866 (N_4866,N_3987,N_3517);
or U4867 (N_4867,N_3990,N_3612);
nand U4868 (N_4868,N_3424,N_3056);
or U4869 (N_4869,N_3575,N_3069);
nor U4870 (N_4870,N_3813,N_3312);
xnor U4871 (N_4871,N_3675,N_3406);
or U4872 (N_4872,N_3392,N_3849);
or U4873 (N_4873,N_3430,N_3842);
or U4874 (N_4874,N_3865,N_3524);
xor U4875 (N_4875,N_3121,N_3110);
and U4876 (N_4876,N_3718,N_3214);
nand U4877 (N_4877,N_3655,N_3173);
xnor U4878 (N_4878,N_3560,N_3711);
xor U4879 (N_4879,N_3270,N_3661);
xnor U4880 (N_4880,N_3024,N_3537);
nor U4881 (N_4881,N_3011,N_3687);
xor U4882 (N_4882,N_3259,N_3434);
and U4883 (N_4883,N_3475,N_3944);
nand U4884 (N_4884,N_3874,N_3885);
or U4885 (N_4885,N_3100,N_3884);
and U4886 (N_4886,N_3209,N_3431);
and U4887 (N_4887,N_3516,N_3935);
and U4888 (N_4888,N_3462,N_3368);
or U4889 (N_4889,N_3370,N_3175);
and U4890 (N_4890,N_3044,N_3259);
xor U4891 (N_4891,N_3717,N_3007);
nand U4892 (N_4892,N_3704,N_3499);
nand U4893 (N_4893,N_3917,N_3287);
nand U4894 (N_4894,N_3706,N_3570);
and U4895 (N_4895,N_3879,N_3623);
nand U4896 (N_4896,N_3233,N_3482);
nand U4897 (N_4897,N_3403,N_3835);
or U4898 (N_4898,N_3362,N_3777);
nor U4899 (N_4899,N_3384,N_3559);
nor U4900 (N_4900,N_3685,N_3882);
and U4901 (N_4901,N_3244,N_3375);
nand U4902 (N_4902,N_3299,N_3970);
xor U4903 (N_4903,N_3036,N_3590);
nor U4904 (N_4904,N_3639,N_3980);
nor U4905 (N_4905,N_3449,N_3492);
and U4906 (N_4906,N_3004,N_3251);
nor U4907 (N_4907,N_3317,N_3565);
nor U4908 (N_4908,N_3462,N_3957);
nand U4909 (N_4909,N_3608,N_3297);
xnor U4910 (N_4910,N_3105,N_3632);
and U4911 (N_4911,N_3269,N_3182);
xnor U4912 (N_4912,N_3651,N_3791);
nand U4913 (N_4913,N_3468,N_3461);
and U4914 (N_4914,N_3154,N_3571);
or U4915 (N_4915,N_3008,N_3416);
nor U4916 (N_4916,N_3243,N_3972);
nand U4917 (N_4917,N_3247,N_3155);
or U4918 (N_4918,N_3364,N_3907);
nand U4919 (N_4919,N_3948,N_3224);
and U4920 (N_4920,N_3271,N_3689);
and U4921 (N_4921,N_3112,N_3312);
and U4922 (N_4922,N_3009,N_3343);
nand U4923 (N_4923,N_3716,N_3199);
and U4924 (N_4924,N_3795,N_3897);
and U4925 (N_4925,N_3970,N_3666);
and U4926 (N_4926,N_3014,N_3417);
nor U4927 (N_4927,N_3939,N_3027);
nor U4928 (N_4928,N_3490,N_3222);
nand U4929 (N_4929,N_3177,N_3075);
nor U4930 (N_4930,N_3658,N_3604);
nand U4931 (N_4931,N_3268,N_3575);
nor U4932 (N_4932,N_3935,N_3993);
or U4933 (N_4933,N_3221,N_3377);
nand U4934 (N_4934,N_3440,N_3967);
nor U4935 (N_4935,N_3372,N_3183);
nor U4936 (N_4936,N_3449,N_3563);
xnor U4937 (N_4937,N_3316,N_3496);
or U4938 (N_4938,N_3474,N_3452);
nand U4939 (N_4939,N_3385,N_3909);
or U4940 (N_4940,N_3585,N_3908);
xor U4941 (N_4941,N_3084,N_3571);
xor U4942 (N_4942,N_3181,N_3376);
nor U4943 (N_4943,N_3441,N_3124);
and U4944 (N_4944,N_3910,N_3953);
nor U4945 (N_4945,N_3594,N_3917);
and U4946 (N_4946,N_3456,N_3390);
and U4947 (N_4947,N_3619,N_3818);
or U4948 (N_4948,N_3664,N_3958);
or U4949 (N_4949,N_3888,N_3856);
and U4950 (N_4950,N_3313,N_3432);
nand U4951 (N_4951,N_3997,N_3517);
xor U4952 (N_4952,N_3239,N_3789);
xnor U4953 (N_4953,N_3937,N_3487);
nor U4954 (N_4954,N_3809,N_3179);
xnor U4955 (N_4955,N_3548,N_3738);
nand U4956 (N_4956,N_3520,N_3261);
and U4957 (N_4957,N_3875,N_3637);
or U4958 (N_4958,N_3134,N_3475);
nand U4959 (N_4959,N_3438,N_3279);
and U4960 (N_4960,N_3188,N_3812);
and U4961 (N_4961,N_3907,N_3947);
nor U4962 (N_4962,N_3650,N_3746);
nor U4963 (N_4963,N_3955,N_3567);
nand U4964 (N_4964,N_3826,N_3429);
and U4965 (N_4965,N_3959,N_3994);
xnor U4966 (N_4966,N_3798,N_3519);
or U4967 (N_4967,N_3178,N_3859);
xnor U4968 (N_4968,N_3840,N_3790);
and U4969 (N_4969,N_3979,N_3207);
or U4970 (N_4970,N_3901,N_3919);
xnor U4971 (N_4971,N_3834,N_3668);
and U4972 (N_4972,N_3083,N_3061);
or U4973 (N_4973,N_3930,N_3698);
xor U4974 (N_4974,N_3823,N_3754);
xnor U4975 (N_4975,N_3021,N_3543);
nor U4976 (N_4976,N_3784,N_3383);
xor U4977 (N_4977,N_3533,N_3144);
nand U4978 (N_4978,N_3629,N_3747);
or U4979 (N_4979,N_3231,N_3702);
nand U4980 (N_4980,N_3306,N_3873);
xor U4981 (N_4981,N_3163,N_3987);
xnor U4982 (N_4982,N_3744,N_3578);
or U4983 (N_4983,N_3104,N_3919);
nand U4984 (N_4984,N_3632,N_3389);
xor U4985 (N_4985,N_3846,N_3766);
and U4986 (N_4986,N_3264,N_3393);
nor U4987 (N_4987,N_3725,N_3316);
nand U4988 (N_4988,N_3358,N_3528);
and U4989 (N_4989,N_3988,N_3929);
nand U4990 (N_4990,N_3128,N_3633);
or U4991 (N_4991,N_3036,N_3298);
and U4992 (N_4992,N_3784,N_3886);
nand U4993 (N_4993,N_3719,N_3001);
nand U4994 (N_4994,N_3705,N_3924);
xnor U4995 (N_4995,N_3014,N_3073);
and U4996 (N_4996,N_3540,N_3731);
or U4997 (N_4997,N_3645,N_3558);
nand U4998 (N_4998,N_3831,N_3167);
nor U4999 (N_4999,N_3804,N_3683);
and U5000 (N_5000,N_4196,N_4376);
or U5001 (N_5001,N_4882,N_4440);
and U5002 (N_5002,N_4582,N_4037);
nor U5003 (N_5003,N_4746,N_4971);
nand U5004 (N_5004,N_4891,N_4159);
xor U5005 (N_5005,N_4980,N_4304);
or U5006 (N_5006,N_4783,N_4527);
nand U5007 (N_5007,N_4325,N_4343);
nand U5008 (N_5008,N_4931,N_4132);
xnor U5009 (N_5009,N_4847,N_4243);
and U5010 (N_5010,N_4462,N_4775);
and U5011 (N_5011,N_4811,N_4076);
and U5012 (N_5012,N_4475,N_4898);
xor U5013 (N_5013,N_4581,N_4574);
or U5014 (N_5014,N_4083,N_4285);
and U5015 (N_5015,N_4602,N_4727);
nor U5016 (N_5016,N_4853,N_4705);
xnor U5017 (N_5017,N_4826,N_4820);
nor U5018 (N_5018,N_4194,N_4982);
nand U5019 (N_5019,N_4320,N_4839);
and U5020 (N_5020,N_4500,N_4695);
xnor U5021 (N_5021,N_4352,N_4426);
nor U5022 (N_5022,N_4437,N_4934);
and U5023 (N_5023,N_4019,N_4796);
or U5024 (N_5024,N_4688,N_4664);
nor U5025 (N_5025,N_4832,N_4039);
and U5026 (N_5026,N_4863,N_4303);
xor U5027 (N_5027,N_4093,N_4556);
nor U5028 (N_5028,N_4924,N_4279);
and U5029 (N_5029,N_4702,N_4254);
nand U5030 (N_5030,N_4234,N_4072);
or U5031 (N_5031,N_4785,N_4681);
and U5032 (N_5032,N_4311,N_4309);
or U5033 (N_5033,N_4950,N_4275);
and U5034 (N_5034,N_4897,N_4703);
nand U5035 (N_5035,N_4116,N_4096);
nand U5036 (N_5036,N_4400,N_4937);
or U5037 (N_5037,N_4877,N_4424);
nor U5038 (N_5038,N_4158,N_4386);
and U5039 (N_5039,N_4113,N_4719);
nand U5040 (N_5040,N_4317,N_4517);
and U5041 (N_5041,N_4207,N_4585);
nand U5042 (N_5042,N_4562,N_4224);
nand U5043 (N_5043,N_4564,N_4095);
and U5044 (N_5044,N_4444,N_4846);
nor U5045 (N_5045,N_4187,N_4670);
or U5046 (N_5046,N_4617,N_4354);
and U5047 (N_5047,N_4435,N_4868);
or U5048 (N_5048,N_4294,N_4412);
nor U5049 (N_5049,N_4876,N_4115);
xnor U5050 (N_5050,N_4804,N_4150);
nand U5051 (N_5051,N_4481,N_4666);
xnor U5052 (N_5052,N_4422,N_4431);
or U5053 (N_5053,N_4884,N_4256);
and U5054 (N_5054,N_4121,N_4339);
and U5055 (N_5055,N_4735,N_4633);
nand U5056 (N_5056,N_4896,N_4554);
xnor U5057 (N_5057,N_4102,N_4053);
xor U5058 (N_5058,N_4949,N_4913);
or U5059 (N_5059,N_4786,N_4830);
and U5060 (N_5060,N_4933,N_4993);
xor U5061 (N_5061,N_4887,N_4097);
and U5062 (N_5062,N_4940,N_4511);
nand U5063 (N_5063,N_4689,N_4212);
nor U5064 (N_5064,N_4484,N_4960);
xnor U5065 (N_5065,N_4507,N_4200);
and U5066 (N_5066,N_4349,N_4359);
xor U5067 (N_5067,N_4405,N_4985);
and U5068 (N_5068,N_4333,N_4394);
nor U5069 (N_5069,N_4206,N_4434);
or U5070 (N_5070,N_4945,N_4742);
nand U5071 (N_5071,N_4432,N_4717);
nor U5072 (N_5072,N_4506,N_4344);
or U5073 (N_5073,N_4061,N_4122);
nor U5074 (N_5074,N_4608,N_4908);
and U5075 (N_5075,N_4370,N_4018);
or U5076 (N_5076,N_4546,N_4544);
xor U5077 (N_5077,N_4246,N_4458);
nand U5078 (N_5078,N_4883,N_4998);
or U5079 (N_5079,N_4621,N_4218);
nand U5080 (N_5080,N_4932,N_4560);
nand U5081 (N_5081,N_4180,N_4542);
nand U5082 (N_5082,N_4916,N_4117);
xnor U5083 (N_5083,N_4084,N_4973);
xor U5084 (N_5084,N_4657,N_4718);
and U5085 (N_5085,N_4905,N_4163);
and U5086 (N_5086,N_4014,N_4690);
nor U5087 (N_5087,N_4185,N_4227);
or U5088 (N_5088,N_4655,N_4318);
and U5089 (N_5089,N_4966,N_4013);
xor U5090 (N_5090,N_4989,N_4332);
and U5091 (N_5091,N_4611,N_4824);
xor U5092 (N_5092,N_4189,N_4045);
nor U5093 (N_5093,N_4699,N_4160);
and U5094 (N_5094,N_4192,N_4648);
or U5095 (N_5095,N_4263,N_4062);
or U5096 (N_5096,N_4360,N_4799);
and U5097 (N_5097,N_4134,N_4576);
nor U5098 (N_5098,N_4645,N_4442);
xor U5099 (N_5099,N_4268,N_4502);
nand U5100 (N_5100,N_4274,N_4569);
nor U5101 (N_5101,N_4822,N_4551);
xnor U5102 (N_5102,N_4384,N_4741);
or U5103 (N_5103,N_4111,N_4030);
nor U5104 (N_5104,N_4778,N_4600);
xnor U5105 (N_5105,N_4629,N_4635);
nor U5106 (N_5106,N_4472,N_4092);
xnor U5107 (N_5107,N_4114,N_4978);
and U5108 (N_5108,N_4235,N_4052);
and U5109 (N_5109,N_4854,N_4994);
nor U5110 (N_5110,N_4406,N_4747);
nand U5111 (N_5111,N_4892,N_4033);
xor U5112 (N_5112,N_4990,N_4557);
or U5113 (N_5113,N_4380,N_4436);
or U5114 (N_5114,N_4547,N_4043);
xor U5115 (N_5115,N_4504,N_4141);
or U5116 (N_5116,N_4772,N_4918);
or U5117 (N_5117,N_4120,N_4181);
or U5118 (N_5118,N_4445,N_4687);
xor U5119 (N_5119,N_4031,N_4907);
nand U5120 (N_5120,N_4813,N_4829);
nor U5121 (N_5121,N_4347,N_4787);
or U5122 (N_5122,N_4425,N_4647);
nand U5123 (N_5123,N_4081,N_4968);
nor U5124 (N_5124,N_4650,N_4776);
and U5125 (N_5125,N_4566,N_4027);
nor U5126 (N_5126,N_4708,N_4129);
nand U5127 (N_5127,N_4329,N_4821);
or U5128 (N_5128,N_4496,N_4624);
or U5129 (N_5129,N_4165,N_4515);
xnor U5130 (N_5130,N_4914,N_4237);
or U5131 (N_5131,N_4010,N_4798);
or U5132 (N_5132,N_4397,N_4872);
or U5133 (N_5133,N_4692,N_4125);
or U5134 (N_5134,N_4273,N_4691);
nand U5135 (N_5135,N_4002,N_4245);
nor U5136 (N_5136,N_4086,N_4539);
and U5137 (N_5137,N_4730,N_4952);
nand U5138 (N_5138,N_4459,N_4886);
xnor U5139 (N_5139,N_4720,N_4843);
nor U5140 (N_5140,N_4963,N_4365);
nand U5141 (N_5141,N_4548,N_4806);
nor U5142 (N_5142,N_4885,N_4499);
or U5143 (N_5143,N_4240,N_4755);
xor U5144 (N_5144,N_4005,N_4056);
xnor U5145 (N_5145,N_4108,N_4906);
nand U5146 (N_5146,N_4172,N_4494);
nor U5147 (N_5147,N_4922,N_4618);
and U5148 (N_5148,N_4954,N_4251);
or U5149 (N_5149,N_4613,N_4233);
or U5150 (N_5150,N_4135,N_4654);
and U5151 (N_5151,N_4679,N_4764);
nor U5152 (N_5152,N_4610,N_4464);
nand U5153 (N_5153,N_4865,N_4797);
or U5154 (N_5154,N_4174,N_4216);
xor U5155 (N_5155,N_4580,N_4751);
and U5156 (N_5156,N_4525,N_4759);
nor U5157 (N_5157,N_4939,N_4678);
xor U5158 (N_5158,N_4082,N_4368);
xnor U5159 (N_5159,N_4300,N_4131);
nor U5160 (N_5160,N_4202,N_4947);
nor U5161 (N_5161,N_4930,N_4659);
nor U5162 (N_5162,N_4941,N_4632);
xor U5163 (N_5163,N_4995,N_4833);
xnor U5164 (N_5164,N_4901,N_4622);
and U5165 (N_5165,N_4334,N_4259);
nor U5166 (N_5166,N_4697,N_4297);
xnor U5167 (N_5167,N_4593,N_4350);
nor U5168 (N_5168,N_4029,N_4249);
or U5169 (N_5169,N_4616,N_4549);
or U5170 (N_5170,N_4091,N_4408);
nand U5171 (N_5171,N_4669,N_4649);
nor U5172 (N_5172,N_4371,N_4565);
xor U5173 (N_5173,N_4143,N_4737);
xnor U5174 (N_5174,N_4501,N_4016);
nor U5175 (N_5175,N_4430,N_4416);
or U5176 (N_5176,N_4676,N_4677);
xor U5177 (N_5177,N_4302,N_4603);
xor U5178 (N_5178,N_4849,N_4178);
nor U5179 (N_5179,N_4470,N_4348);
nor U5180 (N_5180,N_4269,N_4844);
nor U5181 (N_5181,N_4726,N_4293);
xnor U5182 (N_5182,N_4401,N_4402);
nand U5183 (N_5183,N_4861,N_4773);
xor U5184 (N_5184,N_4684,N_4340);
nor U5185 (N_5185,N_4152,N_4673);
and U5186 (N_5186,N_4761,N_4035);
and U5187 (N_5187,N_4623,N_4310);
nor U5188 (N_5188,N_4698,N_4197);
or U5189 (N_5189,N_4722,N_4510);
or U5190 (N_5190,N_4656,N_4837);
nor U5191 (N_5191,N_4757,N_4041);
or U5192 (N_5192,N_4301,N_4578);
or U5193 (N_5193,N_4651,N_4403);
or U5194 (N_5194,N_4970,N_4858);
and U5195 (N_5195,N_4307,N_4848);
nor U5196 (N_5196,N_4381,N_4721);
nor U5197 (N_5197,N_4055,N_4771);
or U5198 (N_5198,N_4419,N_4996);
xor U5199 (N_5199,N_4860,N_4740);
and U5200 (N_5200,N_4377,N_4149);
nand U5201 (N_5201,N_4473,N_4463);
or U5202 (N_5202,N_4151,N_4754);
or U5203 (N_5203,N_4211,N_4864);
and U5204 (N_5204,N_4592,N_4157);
nor U5205 (N_5205,N_4059,N_4079);
xor U5206 (N_5206,N_4888,N_4553);
xor U5207 (N_5207,N_4587,N_4766);
nor U5208 (N_5208,N_4760,N_4792);
and U5209 (N_5209,N_4044,N_4241);
xnor U5210 (N_5210,N_4193,N_4460);
nand U5211 (N_5211,N_4457,N_4714);
nand U5212 (N_5212,N_4953,N_4015);
nor U5213 (N_5213,N_4204,N_4260);
or U5214 (N_5214,N_4244,N_4369);
nand U5215 (N_5215,N_4447,N_4784);
nand U5216 (N_5216,N_4836,N_4733);
nand U5217 (N_5217,N_4319,N_4186);
nor U5218 (N_5218,N_4644,N_4372);
and U5219 (N_5219,N_4599,N_4713);
xor U5220 (N_5220,N_4471,N_4063);
nand U5221 (N_5221,N_4983,N_4028);
and U5222 (N_5222,N_4258,N_4284);
or U5223 (N_5223,N_4628,N_4667);
and U5224 (N_5224,N_4336,N_4351);
and U5225 (N_5225,N_4728,N_4098);
or U5226 (N_5226,N_4382,N_4909);
nand U5227 (N_5227,N_4314,N_4774);
xnor U5228 (N_5228,N_4414,N_4346);
nand U5229 (N_5229,N_4326,N_4630);
nor U5230 (N_5230,N_4631,N_4146);
and U5231 (N_5231,N_4281,N_4040);
nand U5232 (N_5232,N_4429,N_4085);
nand U5233 (N_5233,N_4000,N_4903);
and U5234 (N_5234,N_4110,N_4461);
or U5235 (N_5235,N_4374,N_4021);
and U5236 (N_5236,N_4961,N_4609);
xor U5237 (N_5237,N_4385,N_4127);
or U5238 (N_5238,N_4391,N_4859);
nor U5239 (N_5239,N_4242,N_4208);
nand U5240 (N_5240,N_4105,N_4809);
nor U5241 (N_5241,N_4946,N_4944);
xnor U5242 (N_5242,N_4130,N_4731);
or U5243 (N_5243,N_4800,N_4768);
or U5244 (N_5244,N_4817,N_4514);
and U5245 (N_5245,N_4753,N_4591);
nand U5246 (N_5246,N_4586,N_4841);
and U5247 (N_5247,N_4270,N_4604);
nand U5248 (N_5248,N_4987,N_4283);
and U5249 (N_5249,N_4577,N_4590);
or U5250 (N_5250,N_4606,N_4873);
or U5251 (N_5251,N_4803,N_4453);
nor U5252 (N_5252,N_4355,N_4739);
and U5253 (N_5253,N_4917,N_4605);
nand U5254 (N_5254,N_4915,N_4723);
or U5255 (N_5255,N_4818,N_4221);
nand U5256 (N_5256,N_4926,N_4036);
and U5257 (N_5257,N_4451,N_4477);
nand U5258 (N_5258,N_4520,N_4812);
nand U5259 (N_5259,N_4526,N_4353);
or U5260 (N_5260,N_4571,N_4356);
and U5261 (N_5261,N_4533,N_4443);
xor U5262 (N_5262,N_4674,N_4831);
and U5263 (N_5263,N_4298,N_4265);
or U5264 (N_5264,N_4750,N_4835);
nand U5265 (N_5265,N_4900,N_4073);
xnor U5266 (N_5266,N_4308,N_4252);
or U5267 (N_5267,N_4358,N_4389);
xor U5268 (N_5268,N_4025,N_4049);
or U5269 (N_5269,N_4199,N_4070);
nor U5270 (N_5270,N_4572,N_4749);
or U5271 (N_5271,N_4008,N_4064);
nand U5272 (N_5272,N_4312,N_4524);
nand U5273 (N_5273,N_4153,N_4716);
xor U5274 (N_5274,N_4991,N_4065);
or U5275 (N_5275,N_4663,N_4827);
nand U5276 (N_5276,N_4540,N_4942);
and U5277 (N_5277,N_4438,N_4051);
nor U5278 (N_5278,N_4390,N_4573);
xor U5279 (N_5279,N_4267,N_4485);
and U5280 (N_5280,N_4893,N_4852);
nand U5281 (N_5281,N_4048,N_4230);
and U5282 (N_5282,N_4266,N_4951);
or U5283 (N_5283,N_4902,N_4646);
or U5284 (N_5284,N_4017,N_4675);
nor U5285 (N_5285,N_4929,N_4541);
xor U5286 (N_5286,N_4579,N_4291);
and U5287 (N_5287,N_4958,N_4808);
or U5288 (N_5288,N_4338,N_4222);
nand U5289 (N_5289,N_4815,N_4306);
and U5290 (N_5290,N_4155,N_4142);
nor U5291 (N_5291,N_4228,N_4752);
or U5292 (N_5292,N_4090,N_4099);
xnor U5293 (N_5293,N_4439,N_4450);
xor U5294 (N_5294,N_4066,N_4182);
nor U5295 (N_5295,N_4103,N_4088);
or U5296 (N_5296,N_4870,N_4530);
nand U5297 (N_5297,N_4781,N_4089);
xor U5298 (N_5298,N_4177,N_4253);
and U5299 (N_5299,N_4466,N_4706);
nor U5300 (N_5300,N_4977,N_4169);
and U5301 (N_5301,N_4957,N_4156);
and U5302 (N_5302,N_4383,N_4054);
and U5303 (N_5303,N_4851,N_4094);
xor U5304 (N_5304,N_4660,N_4226);
xor U5305 (N_5305,N_4936,N_4503);
xnor U5306 (N_5306,N_4855,N_4642);
and U5307 (N_5307,N_4173,N_4805);
nand U5308 (N_5308,N_4825,N_4563);
nor U5309 (N_5309,N_4058,N_4528);
nand U5310 (N_5310,N_4175,N_4967);
xnor U5311 (N_5311,N_4545,N_4683);
or U5312 (N_5312,N_4456,N_4509);
xnor U5313 (N_5313,N_4662,N_4489);
nand U5314 (N_5314,N_4838,N_4136);
and U5315 (N_5315,N_4255,N_4060);
nand U5316 (N_5316,N_4984,N_4261);
xnor U5317 (N_5317,N_4550,N_4395);
nand U5318 (N_5318,N_4184,N_4620);
and U5319 (N_5319,N_4535,N_4857);
and U5320 (N_5320,N_4195,N_4583);
nor U5321 (N_5321,N_4322,N_4516);
and U5322 (N_5322,N_4387,N_4328);
and U5323 (N_5323,N_4124,N_4938);
xnor U5324 (N_5324,N_4139,N_4123);
nor U5325 (N_5325,N_4075,N_4828);
nor U5326 (N_5326,N_4441,N_4842);
xnor U5327 (N_5327,N_4162,N_4331);
or U5328 (N_5328,N_4878,N_4508);
xor U5329 (N_5329,N_4969,N_4209);
nor U5330 (N_5330,N_4974,N_4363);
and U5331 (N_5331,N_4100,N_4671);
and U5332 (N_5332,N_4128,N_4046);
nor U5333 (N_5333,N_4479,N_4396);
nand U5334 (N_5334,N_4126,N_4203);
nor U5335 (N_5335,N_4513,N_4619);
and U5336 (N_5336,N_4536,N_4834);
nor U5337 (N_5337,N_4410,N_4788);
and U5338 (N_5338,N_4736,N_4956);
or U5339 (N_5339,N_4379,N_4819);
xor U5340 (N_5340,N_4170,N_4264);
xor U5341 (N_5341,N_4641,N_4715);
or U5342 (N_5342,N_4814,N_4866);
and U5343 (N_5343,N_4552,N_4236);
and U5344 (N_5344,N_4899,N_4250);
and U5345 (N_5345,N_4867,N_4247);
nor U5346 (N_5346,N_4532,N_4191);
xnor U5347 (N_5347,N_4393,N_4487);
nand U5348 (N_5348,N_4006,N_4694);
and U5349 (N_5349,N_4341,N_4042);
nand U5350 (N_5350,N_4313,N_4357);
nand U5351 (N_5351,N_4789,N_4217);
xnor U5352 (N_5352,N_4894,N_4337);
or U5353 (N_5353,N_4965,N_4589);
nor U5354 (N_5354,N_4286,N_4057);
and U5355 (N_5355,N_4144,N_4315);
and U5356 (N_5356,N_4292,N_4032);
and U5357 (N_5357,N_4280,N_4433);
xor U5358 (N_5358,N_4748,N_4067);
and U5359 (N_5359,N_4491,N_4107);
xor U5360 (N_5360,N_4874,N_4568);
or U5361 (N_5361,N_4483,N_4597);
or U5362 (N_5362,N_4047,N_4271);
nand U5363 (N_5363,N_4069,N_4935);
or U5364 (N_5364,N_4188,N_4596);
and U5365 (N_5365,N_4345,N_4215);
or U5366 (N_5366,N_4038,N_4148);
xor U5367 (N_5367,N_4003,N_4004);
xor U5368 (N_5368,N_4278,N_4665);
nand U5369 (N_5369,N_4823,N_4495);
or U5370 (N_5370,N_4588,N_4810);
and U5371 (N_5371,N_4988,N_4636);
or U5372 (N_5372,N_4167,N_4482);
xor U5373 (N_5373,N_4943,N_4637);
or U5374 (N_5374,N_4512,N_4895);
and U5375 (N_5375,N_4871,N_4104);
nor U5376 (N_5376,N_4407,N_4879);
xnor U5377 (N_5377,N_4529,N_4537);
and U5378 (N_5378,N_4734,N_4612);
and U5379 (N_5379,N_4364,N_4106);
and U5380 (N_5380,N_4201,N_4880);
nand U5381 (N_5381,N_4779,N_4680);
nand U5382 (N_5382,N_4919,N_4168);
or U5383 (N_5383,N_4685,N_4986);
xnor U5384 (N_5384,N_4220,N_4962);
nand U5385 (N_5385,N_4179,N_4782);
or U5386 (N_5386,N_4225,N_4904);
or U5387 (N_5387,N_4133,N_4518);
nor U5388 (N_5388,N_4468,N_4321);
or U5389 (N_5389,N_4729,N_4421);
xnor U5390 (N_5390,N_4476,N_4816);
xnor U5391 (N_5391,N_4229,N_4558);
nand U5392 (N_5392,N_4745,N_4166);
xor U5393 (N_5393,N_4519,N_4658);
and U5394 (N_5394,N_4068,N_4807);
nand U5395 (N_5395,N_4087,N_4700);
and U5396 (N_5396,N_4875,N_4210);
xnor U5397 (N_5397,N_4570,N_4625);
or U5398 (N_5398,N_4561,N_4001);
xnor U5399 (N_5399,N_4790,N_4299);
or U5400 (N_5400,N_4454,N_4296);
xnor U5401 (N_5401,N_4335,N_4701);
nand U5402 (N_5402,N_4738,N_4682);
nor U5403 (N_5403,N_4765,N_4626);
or U5404 (N_5404,N_4594,N_4712);
or U5405 (N_5405,N_4493,N_4881);
nor U5406 (N_5406,N_4534,N_4011);
xor U5407 (N_5407,N_4707,N_4955);
xor U5408 (N_5408,N_4007,N_4638);
nor U5409 (N_5409,N_4295,N_4050);
xor U5410 (N_5410,N_4147,N_4024);
nor U5411 (N_5411,N_4672,N_4497);
xnor U5412 (N_5412,N_4762,N_4743);
or U5413 (N_5413,N_4923,N_4595);
nor U5414 (N_5414,N_4975,N_4999);
nor U5415 (N_5415,N_4490,N_4869);
nor U5416 (N_5416,N_4711,N_4219);
or U5417 (N_5417,N_4639,N_4118);
and U5418 (N_5418,N_4492,N_4288);
nand U5419 (N_5419,N_4911,N_4979);
or U5420 (N_5420,N_4465,N_4981);
nand U5421 (N_5421,N_4710,N_4138);
nor U5422 (N_5422,N_4538,N_4272);
xnor U5423 (N_5423,N_4584,N_4290);
nand U5424 (N_5424,N_4119,N_4446);
nor U5425 (N_5425,N_4480,N_4972);
nor U5426 (N_5426,N_4693,N_4257);
nand U5427 (N_5427,N_4388,N_4342);
and U5428 (N_5428,N_4238,N_4959);
or U5429 (N_5429,N_4282,N_4327);
or U5430 (N_5430,N_4398,N_4777);
or U5431 (N_5431,N_4223,N_4575);
or U5432 (N_5432,N_4668,N_4078);
or U5433 (N_5433,N_4474,N_4467);
xor U5434 (N_5434,N_4276,N_4652);
and U5435 (N_5435,N_4022,N_4627);
nor U5436 (N_5436,N_4176,N_4109);
nor U5437 (N_5437,N_4080,N_4140);
or U5438 (N_5438,N_4505,N_4890);
xor U5439 (N_5439,N_4724,N_4420);
or U5440 (N_5440,N_4330,N_4469);
nand U5441 (N_5441,N_4183,N_4034);
nand U5442 (N_5442,N_4361,N_4567);
or U5443 (N_5443,N_4077,N_4411);
nand U5444 (N_5444,N_4417,N_4316);
or U5445 (N_5445,N_4486,N_4262);
nor U5446 (N_5446,N_4927,N_4289);
and U5447 (N_5447,N_4232,N_4696);
nor U5448 (N_5448,N_4850,N_4101);
and U5449 (N_5449,N_4862,N_4964);
xor U5450 (N_5450,N_4427,N_4607);
and U5451 (N_5451,N_4921,N_4305);
nor U5452 (N_5452,N_4794,N_4521);
xnor U5453 (N_5453,N_4231,N_4449);
xnor U5454 (N_5454,N_4171,N_4889);
nor U5455 (N_5455,N_4362,N_4409);
xor U5456 (N_5456,N_4378,N_4023);
or U5457 (N_5457,N_4367,N_4634);
or U5458 (N_5458,N_4423,N_4366);
nand U5459 (N_5459,N_4770,N_4012);
xnor U5460 (N_5460,N_4601,N_4744);
and U5461 (N_5461,N_4428,N_4997);
or U5462 (N_5462,N_4026,N_4455);
and U5463 (N_5463,N_4287,N_4145);
xnor U5464 (N_5464,N_4478,N_4614);
and U5465 (N_5465,N_4543,N_4948);
nor U5466 (N_5466,N_4373,N_4976);
nand U5467 (N_5467,N_4653,N_4112);
nor U5468 (N_5468,N_4615,N_4452);
xor U5469 (N_5469,N_4767,N_4769);
xor U5470 (N_5470,N_4531,N_4074);
or U5471 (N_5471,N_4161,N_4840);
nand U5472 (N_5472,N_4448,N_4732);
nand U5473 (N_5473,N_4845,N_4912);
or U5474 (N_5474,N_4756,N_4137);
nor U5475 (N_5475,N_4928,N_4498);
and U5476 (N_5476,N_4239,N_4214);
nand U5477 (N_5477,N_4780,N_4910);
xnor U5478 (N_5478,N_4791,N_4248);
or U5479 (N_5479,N_4686,N_4375);
and U5480 (N_5480,N_4198,N_4640);
nand U5481 (N_5481,N_4801,N_4071);
or U5482 (N_5482,N_4559,N_4205);
or U5483 (N_5483,N_4522,N_4598);
or U5484 (N_5484,N_4213,N_4793);
nor U5485 (N_5485,N_4392,N_4324);
nor U5486 (N_5486,N_4856,N_4992);
nand U5487 (N_5487,N_4661,N_4758);
xnor U5488 (N_5488,N_4413,N_4418);
nand U5489 (N_5489,N_4523,N_4009);
nand U5490 (N_5490,N_4704,N_4643);
xnor U5491 (N_5491,N_4488,N_4555);
xnor U5492 (N_5492,N_4404,N_4190);
and U5493 (N_5493,N_4795,N_4763);
and U5494 (N_5494,N_4925,N_4920);
nor U5495 (N_5495,N_4164,N_4709);
xnor U5496 (N_5496,N_4020,N_4399);
or U5497 (N_5497,N_4277,N_4415);
xnor U5498 (N_5498,N_4725,N_4323);
xnor U5499 (N_5499,N_4802,N_4154);
xor U5500 (N_5500,N_4473,N_4055);
nor U5501 (N_5501,N_4205,N_4073);
and U5502 (N_5502,N_4441,N_4071);
or U5503 (N_5503,N_4277,N_4740);
nand U5504 (N_5504,N_4213,N_4206);
or U5505 (N_5505,N_4208,N_4423);
and U5506 (N_5506,N_4013,N_4425);
xor U5507 (N_5507,N_4674,N_4020);
nand U5508 (N_5508,N_4185,N_4509);
nor U5509 (N_5509,N_4966,N_4938);
nand U5510 (N_5510,N_4119,N_4359);
or U5511 (N_5511,N_4777,N_4005);
nor U5512 (N_5512,N_4343,N_4489);
or U5513 (N_5513,N_4965,N_4851);
and U5514 (N_5514,N_4050,N_4771);
nand U5515 (N_5515,N_4706,N_4061);
or U5516 (N_5516,N_4742,N_4766);
nor U5517 (N_5517,N_4538,N_4263);
xor U5518 (N_5518,N_4766,N_4554);
and U5519 (N_5519,N_4772,N_4708);
or U5520 (N_5520,N_4026,N_4395);
nor U5521 (N_5521,N_4084,N_4891);
nor U5522 (N_5522,N_4035,N_4598);
and U5523 (N_5523,N_4089,N_4688);
xor U5524 (N_5524,N_4135,N_4929);
or U5525 (N_5525,N_4030,N_4264);
xor U5526 (N_5526,N_4169,N_4096);
xor U5527 (N_5527,N_4061,N_4782);
xnor U5528 (N_5528,N_4707,N_4471);
or U5529 (N_5529,N_4960,N_4229);
xor U5530 (N_5530,N_4093,N_4478);
nor U5531 (N_5531,N_4051,N_4526);
nor U5532 (N_5532,N_4228,N_4041);
and U5533 (N_5533,N_4652,N_4406);
nand U5534 (N_5534,N_4663,N_4600);
and U5535 (N_5535,N_4778,N_4032);
nand U5536 (N_5536,N_4310,N_4973);
xnor U5537 (N_5537,N_4869,N_4275);
and U5538 (N_5538,N_4727,N_4358);
nor U5539 (N_5539,N_4904,N_4161);
nand U5540 (N_5540,N_4833,N_4411);
and U5541 (N_5541,N_4543,N_4548);
nor U5542 (N_5542,N_4425,N_4824);
or U5543 (N_5543,N_4287,N_4582);
xor U5544 (N_5544,N_4100,N_4645);
nor U5545 (N_5545,N_4238,N_4727);
xnor U5546 (N_5546,N_4282,N_4520);
and U5547 (N_5547,N_4238,N_4151);
and U5548 (N_5548,N_4424,N_4911);
nand U5549 (N_5549,N_4640,N_4867);
xor U5550 (N_5550,N_4901,N_4777);
or U5551 (N_5551,N_4196,N_4962);
xor U5552 (N_5552,N_4500,N_4342);
or U5553 (N_5553,N_4542,N_4596);
xnor U5554 (N_5554,N_4486,N_4391);
and U5555 (N_5555,N_4770,N_4112);
nor U5556 (N_5556,N_4201,N_4227);
nand U5557 (N_5557,N_4947,N_4440);
xor U5558 (N_5558,N_4889,N_4656);
and U5559 (N_5559,N_4138,N_4330);
nand U5560 (N_5560,N_4761,N_4398);
nor U5561 (N_5561,N_4410,N_4075);
and U5562 (N_5562,N_4567,N_4045);
or U5563 (N_5563,N_4408,N_4207);
and U5564 (N_5564,N_4688,N_4599);
nand U5565 (N_5565,N_4415,N_4037);
nand U5566 (N_5566,N_4939,N_4938);
nand U5567 (N_5567,N_4079,N_4739);
and U5568 (N_5568,N_4892,N_4160);
nor U5569 (N_5569,N_4862,N_4143);
nand U5570 (N_5570,N_4189,N_4199);
nand U5571 (N_5571,N_4346,N_4221);
xor U5572 (N_5572,N_4808,N_4522);
and U5573 (N_5573,N_4676,N_4942);
xor U5574 (N_5574,N_4194,N_4246);
nand U5575 (N_5575,N_4512,N_4504);
nor U5576 (N_5576,N_4159,N_4314);
nor U5577 (N_5577,N_4891,N_4401);
or U5578 (N_5578,N_4268,N_4636);
nor U5579 (N_5579,N_4561,N_4041);
nand U5580 (N_5580,N_4421,N_4174);
and U5581 (N_5581,N_4635,N_4798);
and U5582 (N_5582,N_4942,N_4971);
or U5583 (N_5583,N_4146,N_4410);
or U5584 (N_5584,N_4479,N_4160);
and U5585 (N_5585,N_4533,N_4422);
nand U5586 (N_5586,N_4814,N_4992);
and U5587 (N_5587,N_4918,N_4745);
xor U5588 (N_5588,N_4234,N_4706);
nor U5589 (N_5589,N_4142,N_4531);
or U5590 (N_5590,N_4039,N_4883);
nor U5591 (N_5591,N_4012,N_4088);
nand U5592 (N_5592,N_4307,N_4280);
nand U5593 (N_5593,N_4254,N_4759);
or U5594 (N_5594,N_4980,N_4667);
and U5595 (N_5595,N_4807,N_4318);
or U5596 (N_5596,N_4615,N_4329);
nor U5597 (N_5597,N_4391,N_4823);
nand U5598 (N_5598,N_4866,N_4628);
xor U5599 (N_5599,N_4084,N_4201);
nand U5600 (N_5600,N_4309,N_4668);
nor U5601 (N_5601,N_4488,N_4061);
and U5602 (N_5602,N_4307,N_4876);
nor U5603 (N_5603,N_4062,N_4704);
nand U5604 (N_5604,N_4078,N_4152);
nand U5605 (N_5605,N_4525,N_4794);
nand U5606 (N_5606,N_4397,N_4172);
nand U5607 (N_5607,N_4157,N_4401);
xnor U5608 (N_5608,N_4807,N_4500);
or U5609 (N_5609,N_4410,N_4175);
nand U5610 (N_5610,N_4272,N_4329);
and U5611 (N_5611,N_4594,N_4387);
or U5612 (N_5612,N_4216,N_4926);
or U5613 (N_5613,N_4959,N_4216);
xor U5614 (N_5614,N_4143,N_4017);
nor U5615 (N_5615,N_4470,N_4046);
and U5616 (N_5616,N_4437,N_4391);
nor U5617 (N_5617,N_4894,N_4755);
nor U5618 (N_5618,N_4900,N_4755);
and U5619 (N_5619,N_4997,N_4599);
nor U5620 (N_5620,N_4932,N_4187);
and U5621 (N_5621,N_4434,N_4615);
nor U5622 (N_5622,N_4385,N_4932);
nand U5623 (N_5623,N_4162,N_4336);
nor U5624 (N_5624,N_4154,N_4844);
or U5625 (N_5625,N_4009,N_4056);
and U5626 (N_5626,N_4228,N_4925);
and U5627 (N_5627,N_4761,N_4413);
xor U5628 (N_5628,N_4076,N_4676);
xor U5629 (N_5629,N_4054,N_4353);
nand U5630 (N_5630,N_4980,N_4391);
nor U5631 (N_5631,N_4444,N_4966);
and U5632 (N_5632,N_4818,N_4751);
xnor U5633 (N_5633,N_4631,N_4010);
or U5634 (N_5634,N_4928,N_4426);
nor U5635 (N_5635,N_4292,N_4604);
nor U5636 (N_5636,N_4409,N_4697);
nor U5637 (N_5637,N_4086,N_4887);
nand U5638 (N_5638,N_4436,N_4682);
nand U5639 (N_5639,N_4449,N_4844);
or U5640 (N_5640,N_4629,N_4158);
or U5641 (N_5641,N_4110,N_4701);
or U5642 (N_5642,N_4448,N_4760);
or U5643 (N_5643,N_4826,N_4372);
nor U5644 (N_5644,N_4355,N_4041);
xor U5645 (N_5645,N_4502,N_4289);
or U5646 (N_5646,N_4830,N_4774);
or U5647 (N_5647,N_4182,N_4578);
nand U5648 (N_5648,N_4930,N_4707);
nor U5649 (N_5649,N_4892,N_4084);
nand U5650 (N_5650,N_4984,N_4773);
xnor U5651 (N_5651,N_4303,N_4104);
xnor U5652 (N_5652,N_4971,N_4671);
or U5653 (N_5653,N_4342,N_4464);
nand U5654 (N_5654,N_4764,N_4211);
nor U5655 (N_5655,N_4413,N_4736);
nand U5656 (N_5656,N_4376,N_4480);
and U5657 (N_5657,N_4360,N_4364);
or U5658 (N_5658,N_4163,N_4618);
xnor U5659 (N_5659,N_4719,N_4604);
xnor U5660 (N_5660,N_4507,N_4616);
nand U5661 (N_5661,N_4732,N_4017);
or U5662 (N_5662,N_4523,N_4324);
nor U5663 (N_5663,N_4257,N_4413);
xor U5664 (N_5664,N_4985,N_4078);
nor U5665 (N_5665,N_4616,N_4270);
xnor U5666 (N_5666,N_4079,N_4125);
or U5667 (N_5667,N_4277,N_4410);
nand U5668 (N_5668,N_4674,N_4373);
nor U5669 (N_5669,N_4352,N_4027);
or U5670 (N_5670,N_4918,N_4570);
and U5671 (N_5671,N_4688,N_4873);
nand U5672 (N_5672,N_4621,N_4099);
nor U5673 (N_5673,N_4739,N_4149);
and U5674 (N_5674,N_4259,N_4843);
and U5675 (N_5675,N_4099,N_4135);
nand U5676 (N_5676,N_4255,N_4581);
or U5677 (N_5677,N_4441,N_4133);
xor U5678 (N_5678,N_4640,N_4902);
or U5679 (N_5679,N_4641,N_4681);
or U5680 (N_5680,N_4673,N_4068);
nor U5681 (N_5681,N_4247,N_4173);
xnor U5682 (N_5682,N_4504,N_4449);
xor U5683 (N_5683,N_4047,N_4286);
and U5684 (N_5684,N_4273,N_4624);
or U5685 (N_5685,N_4519,N_4986);
and U5686 (N_5686,N_4139,N_4605);
or U5687 (N_5687,N_4530,N_4116);
nor U5688 (N_5688,N_4576,N_4099);
nor U5689 (N_5689,N_4460,N_4771);
or U5690 (N_5690,N_4334,N_4903);
nand U5691 (N_5691,N_4325,N_4540);
nand U5692 (N_5692,N_4641,N_4813);
nor U5693 (N_5693,N_4672,N_4358);
or U5694 (N_5694,N_4578,N_4631);
nor U5695 (N_5695,N_4709,N_4613);
nor U5696 (N_5696,N_4467,N_4079);
and U5697 (N_5697,N_4437,N_4450);
nand U5698 (N_5698,N_4318,N_4360);
and U5699 (N_5699,N_4347,N_4699);
nand U5700 (N_5700,N_4902,N_4278);
nor U5701 (N_5701,N_4463,N_4173);
xnor U5702 (N_5702,N_4713,N_4747);
nand U5703 (N_5703,N_4924,N_4881);
and U5704 (N_5704,N_4520,N_4182);
or U5705 (N_5705,N_4267,N_4828);
or U5706 (N_5706,N_4449,N_4670);
and U5707 (N_5707,N_4401,N_4907);
xnor U5708 (N_5708,N_4675,N_4003);
and U5709 (N_5709,N_4755,N_4061);
and U5710 (N_5710,N_4186,N_4333);
nor U5711 (N_5711,N_4485,N_4412);
xnor U5712 (N_5712,N_4796,N_4466);
or U5713 (N_5713,N_4177,N_4833);
or U5714 (N_5714,N_4556,N_4538);
or U5715 (N_5715,N_4714,N_4799);
xnor U5716 (N_5716,N_4572,N_4963);
or U5717 (N_5717,N_4065,N_4144);
nor U5718 (N_5718,N_4224,N_4803);
nor U5719 (N_5719,N_4261,N_4578);
or U5720 (N_5720,N_4385,N_4461);
nor U5721 (N_5721,N_4598,N_4247);
or U5722 (N_5722,N_4899,N_4721);
nor U5723 (N_5723,N_4170,N_4830);
nand U5724 (N_5724,N_4436,N_4690);
or U5725 (N_5725,N_4465,N_4184);
or U5726 (N_5726,N_4457,N_4301);
or U5727 (N_5727,N_4891,N_4886);
or U5728 (N_5728,N_4702,N_4492);
xnor U5729 (N_5729,N_4669,N_4015);
nor U5730 (N_5730,N_4732,N_4961);
xnor U5731 (N_5731,N_4786,N_4555);
xor U5732 (N_5732,N_4279,N_4227);
xnor U5733 (N_5733,N_4752,N_4479);
xnor U5734 (N_5734,N_4097,N_4479);
or U5735 (N_5735,N_4998,N_4121);
nor U5736 (N_5736,N_4837,N_4044);
nor U5737 (N_5737,N_4419,N_4732);
nor U5738 (N_5738,N_4097,N_4752);
xor U5739 (N_5739,N_4246,N_4668);
nand U5740 (N_5740,N_4537,N_4823);
xor U5741 (N_5741,N_4951,N_4615);
xnor U5742 (N_5742,N_4052,N_4786);
xor U5743 (N_5743,N_4265,N_4254);
nand U5744 (N_5744,N_4190,N_4358);
nand U5745 (N_5745,N_4088,N_4907);
xor U5746 (N_5746,N_4499,N_4428);
nor U5747 (N_5747,N_4911,N_4767);
nand U5748 (N_5748,N_4191,N_4645);
or U5749 (N_5749,N_4929,N_4409);
or U5750 (N_5750,N_4077,N_4176);
nand U5751 (N_5751,N_4979,N_4962);
or U5752 (N_5752,N_4845,N_4755);
nor U5753 (N_5753,N_4254,N_4427);
xnor U5754 (N_5754,N_4563,N_4081);
xnor U5755 (N_5755,N_4227,N_4014);
nor U5756 (N_5756,N_4585,N_4223);
and U5757 (N_5757,N_4693,N_4964);
nor U5758 (N_5758,N_4938,N_4540);
xnor U5759 (N_5759,N_4546,N_4585);
nand U5760 (N_5760,N_4317,N_4688);
and U5761 (N_5761,N_4035,N_4497);
and U5762 (N_5762,N_4018,N_4761);
or U5763 (N_5763,N_4652,N_4358);
nor U5764 (N_5764,N_4722,N_4229);
nand U5765 (N_5765,N_4251,N_4608);
or U5766 (N_5766,N_4244,N_4248);
nor U5767 (N_5767,N_4210,N_4174);
xor U5768 (N_5768,N_4099,N_4906);
or U5769 (N_5769,N_4402,N_4717);
and U5770 (N_5770,N_4932,N_4076);
and U5771 (N_5771,N_4153,N_4346);
or U5772 (N_5772,N_4308,N_4213);
and U5773 (N_5773,N_4502,N_4916);
nand U5774 (N_5774,N_4354,N_4232);
or U5775 (N_5775,N_4929,N_4455);
or U5776 (N_5776,N_4793,N_4331);
or U5777 (N_5777,N_4439,N_4775);
or U5778 (N_5778,N_4583,N_4270);
xnor U5779 (N_5779,N_4745,N_4461);
nor U5780 (N_5780,N_4045,N_4820);
or U5781 (N_5781,N_4132,N_4516);
nand U5782 (N_5782,N_4177,N_4436);
xnor U5783 (N_5783,N_4527,N_4060);
and U5784 (N_5784,N_4470,N_4178);
xnor U5785 (N_5785,N_4739,N_4281);
and U5786 (N_5786,N_4365,N_4498);
or U5787 (N_5787,N_4177,N_4196);
and U5788 (N_5788,N_4396,N_4653);
nand U5789 (N_5789,N_4049,N_4398);
nand U5790 (N_5790,N_4598,N_4300);
and U5791 (N_5791,N_4337,N_4311);
nand U5792 (N_5792,N_4226,N_4737);
nor U5793 (N_5793,N_4195,N_4630);
xor U5794 (N_5794,N_4193,N_4793);
and U5795 (N_5795,N_4219,N_4016);
and U5796 (N_5796,N_4374,N_4251);
and U5797 (N_5797,N_4142,N_4965);
or U5798 (N_5798,N_4159,N_4234);
nor U5799 (N_5799,N_4173,N_4578);
or U5800 (N_5800,N_4719,N_4418);
nor U5801 (N_5801,N_4361,N_4250);
xnor U5802 (N_5802,N_4933,N_4065);
xor U5803 (N_5803,N_4643,N_4200);
xor U5804 (N_5804,N_4504,N_4845);
nand U5805 (N_5805,N_4145,N_4040);
nor U5806 (N_5806,N_4188,N_4170);
or U5807 (N_5807,N_4138,N_4683);
xor U5808 (N_5808,N_4919,N_4612);
and U5809 (N_5809,N_4125,N_4080);
nor U5810 (N_5810,N_4732,N_4739);
xnor U5811 (N_5811,N_4633,N_4889);
and U5812 (N_5812,N_4989,N_4626);
nand U5813 (N_5813,N_4374,N_4925);
or U5814 (N_5814,N_4492,N_4084);
nor U5815 (N_5815,N_4343,N_4665);
or U5816 (N_5816,N_4913,N_4851);
nor U5817 (N_5817,N_4181,N_4970);
nor U5818 (N_5818,N_4417,N_4653);
nand U5819 (N_5819,N_4978,N_4919);
nor U5820 (N_5820,N_4236,N_4229);
nor U5821 (N_5821,N_4100,N_4447);
xor U5822 (N_5822,N_4026,N_4607);
nor U5823 (N_5823,N_4335,N_4502);
or U5824 (N_5824,N_4571,N_4597);
nor U5825 (N_5825,N_4949,N_4515);
nor U5826 (N_5826,N_4747,N_4184);
xor U5827 (N_5827,N_4542,N_4647);
nor U5828 (N_5828,N_4851,N_4138);
nand U5829 (N_5829,N_4718,N_4069);
xnor U5830 (N_5830,N_4453,N_4079);
xnor U5831 (N_5831,N_4922,N_4256);
or U5832 (N_5832,N_4936,N_4008);
xnor U5833 (N_5833,N_4650,N_4218);
or U5834 (N_5834,N_4117,N_4368);
or U5835 (N_5835,N_4193,N_4673);
and U5836 (N_5836,N_4522,N_4765);
nor U5837 (N_5837,N_4654,N_4334);
nand U5838 (N_5838,N_4381,N_4643);
xor U5839 (N_5839,N_4110,N_4059);
or U5840 (N_5840,N_4436,N_4515);
nor U5841 (N_5841,N_4723,N_4622);
nor U5842 (N_5842,N_4453,N_4181);
or U5843 (N_5843,N_4235,N_4263);
nor U5844 (N_5844,N_4218,N_4628);
nor U5845 (N_5845,N_4512,N_4536);
or U5846 (N_5846,N_4389,N_4266);
or U5847 (N_5847,N_4643,N_4763);
or U5848 (N_5848,N_4022,N_4147);
xnor U5849 (N_5849,N_4264,N_4125);
nand U5850 (N_5850,N_4970,N_4646);
nand U5851 (N_5851,N_4120,N_4219);
or U5852 (N_5852,N_4354,N_4694);
nand U5853 (N_5853,N_4436,N_4256);
xnor U5854 (N_5854,N_4605,N_4550);
and U5855 (N_5855,N_4024,N_4805);
nor U5856 (N_5856,N_4492,N_4528);
and U5857 (N_5857,N_4236,N_4971);
xor U5858 (N_5858,N_4743,N_4925);
or U5859 (N_5859,N_4748,N_4394);
and U5860 (N_5860,N_4563,N_4354);
and U5861 (N_5861,N_4838,N_4103);
and U5862 (N_5862,N_4496,N_4044);
nor U5863 (N_5863,N_4067,N_4354);
and U5864 (N_5864,N_4704,N_4867);
and U5865 (N_5865,N_4819,N_4822);
or U5866 (N_5866,N_4917,N_4010);
nand U5867 (N_5867,N_4449,N_4589);
xnor U5868 (N_5868,N_4622,N_4107);
nand U5869 (N_5869,N_4701,N_4642);
and U5870 (N_5870,N_4323,N_4825);
nor U5871 (N_5871,N_4144,N_4617);
nor U5872 (N_5872,N_4372,N_4085);
or U5873 (N_5873,N_4727,N_4662);
and U5874 (N_5874,N_4083,N_4018);
nor U5875 (N_5875,N_4084,N_4400);
xnor U5876 (N_5876,N_4421,N_4911);
and U5877 (N_5877,N_4410,N_4178);
nor U5878 (N_5878,N_4926,N_4800);
xor U5879 (N_5879,N_4820,N_4394);
xnor U5880 (N_5880,N_4914,N_4538);
xnor U5881 (N_5881,N_4742,N_4162);
xnor U5882 (N_5882,N_4038,N_4232);
or U5883 (N_5883,N_4690,N_4099);
nand U5884 (N_5884,N_4724,N_4923);
nor U5885 (N_5885,N_4374,N_4247);
nor U5886 (N_5886,N_4306,N_4750);
nor U5887 (N_5887,N_4948,N_4113);
xor U5888 (N_5888,N_4023,N_4019);
xnor U5889 (N_5889,N_4263,N_4786);
or U5890 (N_5890,N_4160,N_4626);
xor U5891 (N_5891,N_4633,N_4038);
and U5892 (N_5892,N_4834,N_4959);
nand U5893 (N_5893,N_4450,N_4765);
nor U5894 (N_5894,N_4041,N_4800);
and U5895 (N_5895,N_4698,N_4979);
or U5896 (N_5896,N_4038,N_4412);
and U5897 (N_5897,N_4846,N_4756);
and U5898 (N_5898,N_4510,N_4484);
and U5899 (N_5899,N_4268,N_4021);
or U5900 (N_5900,N_4142,N_4330);
xor U5901 (N_5901,N_4079,N_4593);
and U5902 (N_5902,N_4672,N_4885);
nand U5903 (N_5903,N_4342,N_4365);
nand U5904 (N_5904,N_4205,N_4245);
or U5905 (N_5905,N_4158,N_4773);
nand U5906 (N_5906,N_4072,N_4573);
and U5907 (N_5907,N_4706,N_4179);
xor U5908 (N_5908,N_4806,N_4069);
nor U5909 (N_5909,N_4048,N_4868);
nor U5910 (N_5910,N_4662,N_4397);
xnor U5911 (N_5911,N_4334,N_4046);
xnor U5912 (N_5912,N_4275,N_4141);
nand U5913 (N_5913,N_4006,N_4600);
xor U5914 (N_5914,N_4161,N_4458);
nand U5915 (N_5915,N_4596,N_4964);
nand U5916 (N_5916,N_4540,N_4171);
xnor U5917 (N_5917,N_4339,N_4074);
nor U5918 (N_5918,N_4792,N_4945);
xnor U5919 (N_5919,N_4405,N_4072);
nand U5920 (N_5920,N_4156,N_4393);
nor U5921 (N_5921,N_4744,N_4532);
and U5922 (N_5922,N_4898,N_4022);
and U5923 (N_5923,N_4826,N_4211);
and U5924 (N_5924,N_4424,N_4727);
and U5925 (N_5925,N_4209,N_4755);
nand U5926 (N_5926,N_4471,N_4649);
xor U5927 (N_5927,N_4306,N_4754);
nand U5928 (N_5928,N_4075,N_4841);
nor U5929 (N_5929,N_4218,N_4036);
nand U5930 (N_5930,N_4752,N_4976);
nand U5931 (N_5931,N_4383,N_4491);
nand U5932 (N_5932,N_4226,N_4083);
nor U5933 (N_5933,N_4456,N_4123);
nor U5934 (N_5934,N_4416,N_4925);
nor U5935 (N_5935,N_4284,N_4834);
and U5936 (N_5936,N_4202,N_4854);
and U5937 (N_5937,N_4091,N_4192);
nand U5938 (N_5938,N_4403,N_4875);
nor U5939 (N_5939,N_4047,N_4863);
nand U5940 (N_5940,N_4652,N_4797);
nand U5941 (N_5941,N_4693,N_4797);
and U5942 (N_5942,N_4464,N_4537);
nor U5943 (N_5943,N_4291,N_4016);
nand U5944 (N_5944,N_4036,N_4906);
and U5945 (N_5945,N_4333,N_4087);
or U5946 (N_5946,N_4500,N_4885);
or U5947 (N_5947,N_4669,N_4986);
or U5948 (N_5948,N_4758,N_4577);
nor U5949 (N_5949,N_4606,N_4226);
or U5950 (N_5950,N_4133,N_4804);
and U5951 (N_5951,N_4740,N_4800);
and U5952 (N_5952,N_4936,N_4840);
nand U5953 (N_5953,N_4952,N_4097);
xor U5954 (N_5954,N_4489,N_4236);
nor U5955 (N_5955,N_4563,N_4341);
xor U5956 (N_5956,N_4610,N_4843);
or U5957 (N_5957,N_4095,N_4182);
nand U5958 (N_5958,N_4983,N_4777);
or U5959 (N_5959,N_4190,N_4749);
nand U5960 (N_5960,N_4645,N_4246);
or U5961 (N_5961,N_4331,N_4981);
nor U5962 (N_5962,N_4134,N_4739);
and U5963 (N_5963,N_4615,N_4212);
and U5964 (N_5964,N_4193,N_4117);
xnor U5965 (N_5965,N_4574,N_4514);
or U5966 (N_5966,N_4212,N_4908);
nor U5967 (N_5967,N_4324,N_4186);
nand U5968 (N_5968,N_4858,N_4415);
nand U5969 (N_5969,N_4621,N_4659);
xor U5970 (N_5970,N_4498,N_4216);
nor U5971 (N_5971,N_4589,N_4486);
nor U5972 (N_5972,N_4099,N_4509);
and U5973 (N_5973,N_4943,N_4119);
nand U5974 (N_5974,N_4870,N_4816);
xnor U5975 (N_5975,N_4307,N_4469);
xor U5976 (N_5976,N_4867,N_4716);
nor U5977 (N_5977,N_4551,N_4960);
xnor U5978 (N_5978,N_4852,N_4206);
nand U5979 (N_5979,N_4965,N_4565);
nand U5980 (N_5980,N_4010,N_4147);
and U5981 (N_5981,N_4970,N_4891);
xor U5982 (N_5982,N_4997,N_4585);
or U5983 (N_5983,N_4989,N_4170);
and U5984 (N_5984,N_4143,N_4482);
nor U5985 (N_5985,N_4110,N_4463);
and U5986 (N_5986,N_4558,N_4451);
xnor U5987 (N_5987,N_4606,N_4403);
nand U5988 (N_5988,N_4809,N_4403);
nor U5989 (N_5989,N_4737,N_4889);
nor U5990 (N_5990,N_4781,N_4380);
or U5991 (N_5991,N_4690,N_4837);
nor U5992 (N_5992,N_4170,N_4557);
nor U5993 (N_5993,N_4192,N_4049);
nor U5994 (N_5994,N_4278,N_4416);
and U5995 (N_5995,N_4648,N_4690);
xnor U5996 (N_5996,N_4816,N_4379);
and U5997 (N_5997,N_4979,N_4130);
xnor U5998 (N_5998,N_4736,N_4054);
nor U5999 (N_5999,N_4144,N_4847);
xor U6000 (N_6000,N_5888,N_5697);
or U6001 (N_6001,N_5304,N_5122);
xnor U6002 (N_6002,N_5693,N_5193);
xor U6003 (N_6003,N_5300,N_5802);
nand U6004 (N_6004,N_5833,N_5967);
nand U6005 (N_6005,N_5924,N_5238);
or U6006 (N_6006,N_5762,N_5814);
nand U6007 (N_6007,N_5652,N_5959);
nor U6008 (N_6008,N_5824,N_5742);
xnor U6009 (N_6009,N_5582,N_5889);
nand U6010 (N_6010,N_5328,N_5326);
nand U6011 (N_6011,N_5230,N_5963);
nand U6012 (N_6012,N_5797,N_5110);
xor U6013 (N_6013,N_5738,N_5320);
nand U6014 (N_6014,N_5472,N_5624);
and U6015 (N_6015,N_5861,N_5043);
xnor U6016 (N_6016,N_5605,N_5313);
nand U6017 (N_6017,N_5239,N_5447);
and U6018 (N_6018,N_5126,N_5836);
nand U6019 (N_6019,N_5612,N_5021);
nand U6020 (N_6020,N_5030,N_5800);
nand U6021 (N_6021,N_5529,N_5808);
or U6022 (N_6022,N_5669,N_5278);
nor U6023 (N_6023,N_5898,N_5567);
nor U6024 (N_6024,N_5639,N_5465);
nand U6025 (N_6025,N_5779,N_5407);
or U6026 (N_6026,N_5773,N_5466);
nand U6027 (N_6027,N_5401,N_5424);
or U6028 (N_6028,N_5728,N_5191);
or U6029 (N_6029,N_5558,N_5753);
xor U6030 (N_6030,N_5720,N_5055);
nand U6031 (N_6031,N_5442,N_5537);
nor U6032 (N_6032,N_5458,N_5976);
or U6033 (N_6033,N_5283,N_5526);
nor U6034 (N_6034,N_5091,N_5979);
nand U6035 (N_6035,N_5205,N_5410);
and U6036 (N_6036,N_5020,N_5332);
and U6037 (N_6037,N_5569,N_5983);
xnor U6038 (N_6038,N_5518,N_5668);
and U6039 (N_6039,N_5513,N_5766);
or U6040 (N_6040,N_5843,N_5428);
nand U6041 (N_6041,N_5207,N_5658);
xnor U6042 (N_6042,N_5461,N_5974);
xnor U6043 (N_6043,N_5370,N_5094);
nand U6044 (N_6044,N_5900,N_5998);
nor U6045 (N_6045,N_5684,N_5689);
or U6046 (N_6046,N_5215,N_5895);
nand U6047 (N_6047,N_5835,N_5904);
nor U6048 (N_6048,N_5760,N_5830);
xor U6049 (N_6049,N_5681,N_5040);
nor U6050 (N_6050,N_5364,N_5457);
nand U6051 (N_6051,N_5573,N_5908);
and U6052 (N_6052,N_5548,N_5295);
or U6053 (N_6053,N_5910,N_5726);
or U6054 (N_6054,N_5148,N_5616);
nand U6055 (N_6055,N_5003,N_5377);
and U6056 (N_6056,N_5663,N_5670);
nand U6057 (N_6057,N_5919,N_5866);
nand U6058 (N_6058,N_5378,N_5108);
nor U6059 (N_6059,N_5783,N_5851);
xor U6060 (N_6060,N_5539,N_5488);
and U6061 (N_6061,N_5957,N_5025);
and U6062 (N_6062,N_5072,N_5867);
xor U6063 (N_6063,N_5449,N_5599);
xnor U6064 (N_6064,N_5228,N_5109);
nand U6065 (N_6065,N_5994,N_5568);
nand U6066 (N_6066,N_5501,N_5206);
xor U6067 (N_6067,N_5199,N_5279);
or U6068 (N_6068,N_5677,N_5293);
nor U6069 (N_6069,N_5188,N_5388);
xor U6070 (N_6070,N_5446,N_5035);
nor U6071 (N_6071,N_5099,N_5724);
xnor U6072 (N_6072,N_5009,N_5068);
xor U6073 (N_6073,N_5982,N_5112);
and U6074 (N_6074,N_5267,N_5318);
xnor U6075 (N_6075,N_5225,N_5392);
nand U6076 (N_6076,N_5553,N_5417);
or U6077 (N_6077,N_5528,N_5981);
and U6078 (N_6078,N_5700,N_5602);
xor U6079 (N_6079,N_5273,N_5234);
nor U6080 (N_6080,N_5036,N_5868);
nor U6081 (N_6081,N_5923,N_5419);
nor U6082 (N_6082,N_5363,N_5477);
xnor U6083 (N_6083,N_5949,N_5022);
nand U6084 (N_6084,N_5512,N_5141);
xnor U6085 (N_6085,N_5819,N_5823);
or U6086 (N_6086,N_5408,N_5792);
or U6087 (N_6087,N_5996,N_5758);
nor U6088 (N_6088,N_5805,N_5849);
and U6089 (N_6089,N_5655,N_5717);
xor U6090 (N_6090,N_5361,N_5033);
nor U6091 (N_6091,N_5761,N_5358);
and U6092 (N_6092,N_5649,N_5827);
and U6093 (N_6093,N_5777,N_5789);
nor U6094 (N_6094,N_5166,N_5445);
nor U6095 (N_6095,N_5044,N_5479);
or U6096 (N_6096,N_5354,N_5365);
xnor U6097 (N_6097,N_5591,N_5580);
nand U6098 (N_6098,N_5715,N_5351);
nand U6099 (N_6099,N_5990,N_5067);
nor U6100 (N_6100,N_5809,N_5653);
nand U6101 (N_6101,N_5610,N_5414);
or U6102 (N_6102,N_5375,N_5884);
and U6103 (N_6103,N_5379,N_5810);
nand U6104 (N_6104,N_5050,N_5588);
xnor U6105 (N_6105,N_5498,N_5947);
nor U6106 (N_6106,N_5807,N_5570);
or U6107 (N_6107,N_5221,N_5916);
xor U6108 (N_6108,N_5418,N_5864);
xnor U6109 (N_6109,N_5015,N_5059);
and U6110 (N_6110,N_5984,N_5355);
or U6111 (N_6111,N_5285,N_5121);
and U6112 (N_6112,N_5821,N_5942);
and U6113 (N_6113,N_5662,N_5995);
or U6114 (N_6114,N_5000,N_5269);
and U6115 (N_6115,N_5493,N_5989);
nand U6116 (N_6116,N_5322,N_5846);
or U6117 (N_6117,N_5891,N_5048);
or U6118 (N_6118,N_5063,N_5312);
xor U6119 (N_6119,N_5769,N_5552);
and U6120 (N_6120,N_5422,N_5385);
or U6121 (N_6121,N_5775,N_5223);
nand U6122 (N_6122,N_5075,N_5511);
xnor U6123 (N_6123,N_5741,N_5400);
nand U6124 (N_6124,N_5540,N_5462);
or U6125 (N_6125,N_5444,N_5659);
xnor U6126 (N_6126,N_5265,N_5464);
or U6127 (N_6127,N_5127,N_5887);
nand U6128 (N_6128,N_5679,N_5186);
or U6129 (N_6129,N_5058,N_5394);
nor U6130 (N_6130,N_5382,N_5832);
or U6131 (N_6131,N_5787,N_5443);
and U6132 (N_6132,N_5842,N_5156);
nand U6133 (N_6133,N_5712,N_5826);
nand U6134 (N_6134,N_5794,N_5241);
nand U6135 (N_6135,N_5502,N_5747);
nor U6136 (N_6136,N_5018,N_5237);
xnor U6137 (N_6137,N_5470,N_5771);
or U6138 (N_6138,N_5294,N_5426);
nand U6139 (N_6139,N_5157,N_5521);
and U6140 (N_6140,N_5271,N_5071);
or U6141 (N_6141,N_5115,N_5510);
xor U6142 (N_6142,N_5371,N_5671);
or U6143 (N_6143,N_5686,N_5813);
nor U6144 (N_6144,N_5154,N_5913);
nand U6145 (N_6145,N_5803,N_5985);
nor U6146 (N_6146,N_5174,N_5874);
xor U6147 (N_6147,N_5841,N_5829);
or U6148 (N_6148,N_5232,N_5324);
xor U6149 (N_6149,N_5703,N_5111);
nor U6150 (N_6150,N_5434,N_5439);
nor U6151 (N_6151,N_5594,N_5423);
and U6152 (N_6152,N_5343,N_5336);
xor U6153 (N_6153,N_5459,N_5116);
nand U6154 (N_6154,N_5276,N_5845);
nand U6155 (N_6155,N_5871,N_5574);
and U6156 (N_6156,N_5484,N_5218);
xor U6157 (N_6157,N_5604,N_5413);
xnor U6158 (N_6158,N_5956,N_5796);
or U6159 (N_6159,N_5878,N_5245);
xor U6160 (N_6160,N_5455,N_5136);
nor U6161 (N_6161,N_5759,N_5585);
nand U6162 (N_6162,N_5212,N_5793);
nor U6163 (N_6163,N_5259,N_5281);
or U6164 (N_6164,N_5630,N_5219);
and U6165 (N_6165,N_5691,N_5535);
or U6166 (N_6166,N_5905,N_5161);
and U6167 (N_6167,N_5032,N_5646);
and U6168 (N_6168,N_5229,N_5028);
and U6169 (N_6169,N_5600,N_5523);
nand U6170 (N_6170,N_5804,N_5678);
or U6171 (N_6171,N_5782,N_5489);
or U6172 (N_6172,N_5119,N_5708);
or U6173 (N_6173,N_5150,N_5965);
and U6174 (N_6174,N_5093,N_5914);
and U6175 (N_6175,N_5881,N_5969);
xor U6176 (N_6176,N_5356,N_5638);
nand U6177 (N_6177,N_5690,N_5216);
nand U6178 (N_6178,N_5897,N_5946);
or U6179 (N_6179,N_5516,N_5393);
and U6180 (N_6180,N_5340,N_5374);
nand U6181 (N_6181,N_5549,N_5896);
and U6182 (N_6182,N_5123,N_5860);
or U6183 (N_6183,N_5714,N_5817);
or U6184 (N_6184,N_5270,N_5938);
nor U6185 (N_6185,N_5926,N_5197);
and U6186 (N_6186,N_5873,N_5791);
nand U6187 (N_6187,N_5673,N_5146);
nor U6188 (N_6188,N_5389,N_5348);
xnor U6189 (N_6189,N_5980,N_5233);
nor U6190 (N_6190,N_5615,N_5092);
nand U6191 (N_6191,N_5756,N_5785);
nor U6192 (N_6192,N_5001,N_5194);
or U6193 (N_6193,N_5383,N_5576);
or U6194 (N_6194,N_5227,N_5149);
or U6195 (N_6195,N_5460,N_5357);
xnor U6196 (N_6196,N_5587,N_5837);
or U6197 (N_6197,N_5920,N_5718);
nor U6198 (N_6198,N_5192,N_5883);
and U6199 (N_6199,N_5546,N_5262);
or U6200 (N_6200,N_5258,N_5080);
and U6201 (N_6201,N_5902,N_5491);
and U6202 (N_6202,N_5748,N_5554);
xor U6203 (N_6203,N_5261,N_5704);
nand U6204 (N_6204,N_5863,N_5153);
nand U6205 (N_6205,N_5972,N_5171);
xnor U6206 (N_6206,N_5243,N_5432);
nor U6207 (N_6207,N_5142,N_5155);
nand U6208 (N_6208,N_5289,N_5143);
and U6209 (N_6209,N_5534,N_5515);
nand U6210 (N_6210,N_5006,N_5654);
or U6211 (N_6211,N_5330,N_5812);
nand U6212 (N_6212,N_5179,N_5625);
xnor U6213 (N_6213,N_5073,N_5606);
nand U6214 (N_6214,N_5007,N_5945);
nor U6215 (N_6215,N_5104,N_5672);
nand U6216 (N_6216,N_5359,N_5505);
and U6217 (N_6217,N_5380,N_5381);
or U6218 (N_6218,N_5869,N_5931);
or U6219 (N_6219,N_5211,N_5027);
or U6220 (N_6220,N_5165,N_5590);
nand U6221 (N_6221,N_5469,N_5577);
nor U6222 (N_6222,N_5209,N_5189);
nand U6223 (N_6223,N_5347,N_5848);
nand U6224 (N_6224,N_5463,N_5499);
xor U6225 (N_6225,N_5744,N_5079);
nand U6226 (N_6226,N_5288,N_5768);
nand U6227 (N_6227,N_5362,N_5941);
nand U6228 (N_6228,N_5065,N_5120);
xnor U6229 (N_6229,N_5066,N_5522);
nand U6230 (N_6230,N_5632,N_5396);
and U6231 (N_6231,N_5251,N_5917);
nor U6232 (N_6232,N_5042,N_5431);
nand U6233 (N_6233,N_5964,N_5342);
xnor U6234 (N_6234,N_5729,N_5406);
nand U6235 (N_6235,N_5618,N_5029);
or U6236 (N_6236,N_5563,N_5436);
and U6237 (N_6237,N_5933,N_5547);
nand U6238 (N_6238,N_5482,N_5593);
nand U6239 (N_6239,N_5685,N_5627);
and U6240 (N_6240,N_5709,N_5629);
nand U6241 (N_6241,N_5263,N_5088);
nand U6242 (N_6242,N_5564,N_5101);
nor U6243 (N_6243,N_5244,N_5628);
and U6244 (N_6244,N_5187,N_5642);
xnor U6245 (N_6245,N_5531,N_5064);
nor U6246 (N_6246,N_5087,N_5640);
xor U6247 (N_6247,N_5719,N_5822);
or U6248 (N_6248,N_5305,N_5085);
xor U6249 (N_6249,N_5614,N_5453);
xnor U6250 (N_6250,N_5284,N_5977);
or U6251 (N_6251,N_5702,N_5637);
nand U6252 (N_6252,N_5114,N_5317);
and U6253 (N_6253,N_5710,N_5158);
and U6254 (N_6254,N_5429,N_5550);
or U6255 (N_6255,N_5277,N_5944);
or U6256 (N_6256,N_5954,N_5476);
nand U6257 (N_6257,N_5858,N_5788);
nand U6258 (N_6258,N_5175,N_5506);
or U6259 (N_6259,N_5831,N_5196);
nor U6260 (N_6260,N_5152,N_5943);
nor U6261 (N_6261,N_5303,N_5405);
and U6262 (N_6262,N_5057,N_5236);
nand U6263 (N_6263,N_5090,N_5774);
and U6264 (N_6264,N_5598,N_5930);
xnor U6265 (N_6265,N_5815,N_5879);
nand U6266 (N_6266,N_5096,N_5200);
nand U6267 (N_6267,N_5584,N_5222);
and U6268 (N_6268,N_5765,N_5260);
nand U6269 (N_6269,N_5369,N_5940);
nand U6270 (N_6270,N_5409,N_5387);
and U6271 (N_6271,N_5695,N_5743);
nand U6272 (N_6272,N_5854,N_5880);
or U6273 (N_6273,N_5333,N_5705);
nand U6274 (N_6274,N_5853,N_5133);
xor U6275 (N_6275,N_5301,N_5611);
nor U6276 (N_6276,N_5666,N_5339);
xor U6277 (N_6277,N_5648,N_5935);
and U6278 (N_6278,N_5008,N_5195);
and U6279 (N_6279,N_5962,N_5562);
nor U6280 (N_6280,N_5046,N_5780);
xor U6281 (N_6281,N_5970,N_5083);
and U6282 (N_6282,N_5772,N_5138);
and U6283 (N_6283,N_5275,N_5524);
and U6284 (N_6284,N_5737,N_5013);
nor U6285 (N_6285,N_5635,N_5016);
nand U6286 (N_6286,N_5183,N_5975);
xor U6287 (N_6287,N_5286,N_5352);
nor U6288 (N_6288,N_5082,N_5816);
and U6289 (N_6289,N_5078,N_5253);
nor U6290 (N_6290,N_5494,N_5680);
or U6291 (N_6291,N_5918,N_5372);
nor U6292 (N_6292,N_5621,N_5037);
nand U6293 (N_6293,N_5163,N_5958);
or U6294 (N_6294,N_5725,N_5100);
xnor U6295 (N_6295,N_5017,N_5749);
nand U6296 (N_6296,N_5107,N_5168);
and U6297 (N_6297,N_5485,N_5315);
and U6298 (N_6298,N_5214,N_5852);
and U6299 (N_6299,N_5692,N_5948);
nor U6300 (N_6300,N_5732,N_5438);
xnor U6301 (N_6301,N_5840,N_5925);
xnor U6302 (N_6302,N_5665,N_5583);
xor U6303 (N_6303,N_5242,N_5473);
nor U6304 (N_6304,N_5292,N_5249);
nor U6305 (N_6305,N_5899,N_5723);
and U6306 (N_6306,N_5177,N_5592);
nor U6307 (N_6307,N_5151,N_5565);
nor U6308 (N_6308,N_5901,N_5280);
and U6309 (N_6309,N_5538,N_5204);
xor U6310 (N_6310,N_5145,N_5575);
xor U6311 (N_6311,N_5329,N_5937);
and U6312 (N_6312,N_5581,N_5254);
nand U6313 (N_6313,N_5334,N_5450);
xor U6314 (N_6314,N_5213,N_5299);
nor U6315 (N_6315,N_5801,N_5694);
nand U6316 (N_6316,N_5993,N_5014);
and U6317 (N_6317,N_5164,N_5786);
xnor U6318 (N_6318,N_5492,N_5520);
xnor U6319 (N_6319,N_5291,N_5951);
xnor U6320 (N_6320,N_5038,N_5160);
nor U6321 (N_6321,N_5266,N_5248);
xor U6322 (N_6322,N_5256,N_5857);
nor U6323 (N_6323,N_5129,N_5561);
nor U6324 (N_6324,N_5325,N_5246);
nand U6325 (N_6325,N_5620,N_5026);
or U6326 (N_6326,N_5345,N_5113);
nor U6327 (N_6327,N_5566,N_5571);
or U6328 (N_6328,N_5471,N_5437);
nor U6329 (N_6329,N_5316,N_5024);
xnor U6330 (N_6330,N_5707,N_5346);
xnor U6331 (N_6331,N_5882,N_5435);
xor U6332 (N_6332,N_5847,N_5201);
and U6333 (N_6333,N_5595,N_5532);
nand U6334 (N_6334,N_5274,N_5674);
or U6335 (N_6335,N_5327,N_5736);
nand U6336 (N_6336,N_5631,N_5391);
or U6337 (N_6337,N_5433,N_5536);
and U6338 (N_6338,N_5739,N_5384);
or U6339 (N_6339,N_5496,N_5420);
nand U6340 (N_6340,N_5118,N_5633);
or U6341 (N_6341,N_5481,N_5335);
nand U6342 (N_6342,N_5162,N_5130);
nor U6343 (N_6343,N_5416,N_5656);
xor U6344 (N_6344,N_5172,N_5876);
xor U6345 (N_6345,N_5667,N_5607);
xor U6346 (N_6346,N_5608,N_5514);
xor U6347 (N_6347,N_5039,N_5240);
nor U6348 (N_6348,N_5440,N_5184);
nor U6349 (N_6349,N_5906,N_5302);
and U6350 (N_6350,N_5235,N_5395);
xor U6351 (N_6351,N_5820,N_5634);
or U6352 (N_6352,N_5102,N_5504);
and U6353 (N_6353,N_5456,N_5031);
nand U6354 (N_6354,N_5750,N_5745);
and U6355 (N_6355,N_5997,N_5799);
and U6356 (N_6356,N_5675,N_5004);
or U6357 (N_6357,N_5323,N_5311);
or U6358 (N_6358,N_5106,N_5716);
xor U6359 (N_6359,N_5202,N_5170);
or U6360 (N_6360,N_5856,N_5427);
or U6361 (N_6361,N_5641,N_5727);
nor U6362 (N_6362,N_5041,N_5986);
nand U6363 (N_6363,N_5936,N_5603);
nor U6364 (N_6364,N_5002,N_5005);
xnor U6365 (N_6365,N_5934,N_5870);
or U6366 (N_6366,N_5733,N_5203);
nand U6367 (N_6367,N_5134,N_5398);
xnor U6368 (N_6368,N_5688,N_5746);
and U6369 (N_6369,N_5023,N_5767);
nand U6370 (N_6370,N_5754,N_5474);
nand U6371 (N_6371,N_5706,N_5660);
or U6372 (N_6372,N_5875,N_5676);
nor U6373 (N_6373,N_5084,N_5525);
and U6374 (N_6374,N_5403,N_5839);
and U6375 (N_6375,N_5250,N_5507);
nor U6376 (N_6376,N_5045,N_5623);
and U6377 (N_6377,N_5337,N_5198);
nor U6378 (N_6378,N_5467,N_5838);
nand U6379 (N_6379,N_5661,N_5541);
nor U6380 (N_6380,N_5220,N_5950);
or U6381 (N_6381,N_5349,N_5907);
or U6382 (N_6382,N_5415,N_5784);
or U6383 (N_6383,N_5763,N_5961);
and U6384 (N_6384,N_5644,N_5180);
or U6385 (N_6385,N_5117,N_5555);
nor U6386 (N_6386,N_5651,N_5734);
nor U6387 (N_6387,N_5069,N_5139);
xor U6388 (N_6388,N_5721,N_5911);
nor U6389 (N_6389,N_5287,N_5297);
and U6390 (N_6390,N_5308,N_5696);
nand U6391 (N_6391,N_5862,N_5097);
or U6392 (N_6392,N_5664,N_5503);
xor U6393 (N_6393,N_5795,N_5764);
and U6394 (N_6394,N_5572,N_5076);
or U6395 (N_6395,N_5527,N_5210);
nand U6396 (N_6396,N_5892,N_5735);
xnor U6397 (N_6397,N_5144,N_5955);
nand U6398 (N_6398,N_5617,N_5991);
xor U6399 (N_6399,N_5921,N_5190);
or U6400 (N_6400,N_5077,N_5790);
and U6401 (N_6401,N_5257,N_5579);
and U6402 (N_6402,N_5089,N_5519);
xor U6403 (N_6403,N_5647,N_5886);
xor U6404 (N_6404,N_5178,N_5098);
nand U6405 (N_6405,N_5844,N_5103);
or U6406 (N_6406,N_5645,N_5282);
or U6407 (N_6407,N_5344,N_5255);
and U6408 (N_6408,N_5953,N_5601);
nand U6409 (N_6409,N_5074,N_5131);
and U6410 (N_6410,N_5971,N_5751);
or U6411 (N_6411,N_5872,N_5885);
nor U6412 (N_6412,N_5051,N_5508);
and U6413 (N_6413,N_5912,N_5966);
nor U6414 (N_6414,N_5855,N_5341);
or U6415 (N_6415,N_5061,N_5557);
xor U6416 (N_6416,N_5530,N_5310);
nor U6417 (N_6417,N_5386,N_5441);
or U6418 (N_6418,N_5988,N_5894);
nand U6419 (N_6419,N_5338,N_5306);
nand U6420 (N_6420,N_5877,N_5296);
or U6421 (N_6421,N_5560,N_5366);
nand U6422 (N_6422,N_5825,N_5740);
and U6423 (N_6423,N_5321,N_5181);
nor U6424 (N_6424,N_5682,N_5609);
xor U6425 (N_6425,N_5319,N_5722);
or U6426 (N_6426,N_5404,N_5757);
or U6427 (N_6427,N_5095,N_5999);
and U6428 (N_6428,N_5368,N_5711);
nor U6429 (N_6429,N_5376,N_5486);
and U6430 (N_6430,N_5132,N_5425);
nor U6431 (N_6431,N_5834,N_5657);
nor U6432 (N_6432,N_5701,N_5052);
nor U6433 (N_6433,N_5487,N_5865);
and U6434 (N_6434,N_5411,N_5850);
or U6435 (N_6435,N_5056,N_5643);
and U6436 (N_6436,N_5909,N_5053);
and U6437 (N_6437,N_5176,N_5596);
nand U6438 (N_6438,N_5147,N_5252);
nand U6439 (N_6439,N_5698,N_5890);
xor U6440 (N_6440,N_5070,N_5928);
or U6441 (N_6441,N_5360,N_5208);
and U6442 (N_6442,N_5770,N_5622);
nor U6443 (N_6443,N_5135,N_5390);
xor U6444 (N_6444,N_5011,N_5290);
nand U6445 (N_6445,N_5128,N_5500);
xor U6446 (N_6446,N_5903,N_5012);
or U6447 (N_6447,N_5929,N_5086);
nand U6448 (N_6448,N_5034,N_5922);
xnor U6449 (N_6449,N_5586,N_5397);
nand U6450 (N_6450,N_5798,N_5185);
xor U6451 (N_6451,N_5992,N_5893);
nand U6452 (N_6452,N_5543,N_5578);
nor U6453 (N_6453,N_5452,N_5224);
nand U6454 (N_6454,N_5960,N_5402);
xor U6455 (N_6455,N_5619,N_5399);
or U6456 (N_6456,N_5968,N_5687);
or U6457 (N_6457,N_5478,N_5331);
nand U6458 (N_6458,N_5987,N_5019);
nor U6459 (N_6459,N_5730,N_5373);
nor U6460 (N_6460,N_5081,N_5495);
or U6461 (N_6461,N_5350,N_5060);
nor U6462 (N_6462,N_5613,N_5713);
and U6463 (N_6463,N_5353,N_5451);
and U6464 (N_6464,N_5159,N_5781);
or U6465 (N_6465,N_5231,N_5309);
nor U6466 (N_6466,N_5533,N_5626);
xor U6467 (N_6467,N_5226,N_5927);
xnor U6468 (N_6468,N_5752,N_5448);
nand U6469 (N_6469,N_5828,N_5054);
nand U6470 (N_6470,N_5182,N_5264);
xor U6471 (N_6471,N_5509,N_5137);
nor U6472 (N_6472,N_5811,N_5699);
xor U6473 (N_6473,N_5272,N_5973);
and U6474 (N_6474,N_5490,N_5217);
nand U6475 (N_6475,N_5544,N_5683);
xnor U6476 (N_6476,N_5545,N_5047);
nand U6477 (N_6477,N_5468,N_5542);
nor U6478 (N_6478,N_5454,N_5932);
or U6479 (N_6479,N_5650,N_5167);
nor U6480 (N_6480,N_5939,N_5755);
xnor U6481 (N_6481,N_5475,N_5298);
and U6482 (N_6482,N_5049,N_5952);
and U6483 (N_6483,N_5367,N_5589);
xnor U6484 (N_6484,N_5307,N_5806);
xnor U6485 (N_6485,N_5731,N_5597);
nor U6486 (N_6486,N_5105,N_5497);
nand U6487 (N_6487,N_5268,N_5776);
and U6488 (N_6488,N_5483,N_5140);
xnor U6489 (N_6489,N_5859,N_5480);
nand U6490 (N_6490,N_5978,N_5314);
xor U6491 (N_6491,N_5517,N_5915);
nor U6492 (N_6492,N_5778,N_5247);
nor U6493 (N_6493,N_5421,N_5412);
or U6494 (N_6494,N_5636,N_5124);
nor U6495 (N_6495,N_5551,N_5430);
and U6496 (N_6496,N_5010,N_5173);
xor U6497 (N_6497,N_5062,N_5559);
and U6498 (N_6498,N_5818,N_5169);
xnor U6499 (N_6499,N_5556,N_5125);
and U6500 (N_6500,N_5528,N_5997);
xnor U6501 (N_6501,N_5257,N_5035);
or U6502 (N_6502,N_5688,N_5830);
xnor U6503 (N_6503,N_5487,N_5662);
nor U6504 (N_6504,N_5628,N_5003);
and U6505 (N_6505,N_5293,N_5965);
xnor U6506 (N_6506,N_5294,N_5366);
xor U6507 (N_6507,N_5168,N_5824);
or U6508 (N_6508,N_5371,N_5546);
nor U6509 (N_6509,N_5102,N_5075);
or U6510 (N_6510,N_5460,N_5184);
or U6511 (N_6511,N_5028,N_5623);
nand U6512 (N_6512,N_5507,N_5832);
and U6513 (N_6513,N_5861,N_5649);
xor U6514 (N_6514,N_5121,N_5598);
and U6515 (N_6515,N_5912,N_5108);
and U6516 (N_6516,N_5767,N_5236);
nor U6517 (N_6517,N_5921,N_5868);
and U6518 (N_6518,N_5638,N_5015);
and U6519 (N_6519,N_5839,N_5149);
and U6520 (N_6520,N_5620,N_5559);
or U6521 (N_6521,N_5578,N_5488);
or U6522 (N_6522,N_5068,N_5082);
and U6523 (N_6523,N_5726,N_5148);
nand U6524 (N_6524,N_5502,N_5535);
nor U6525 (N_6525,N_5781,N_5042);
or U6526 (N_6526,N_5869,N_5087);
xor U6527 (N_6527,N_5949,N_5786);
and U6528 (N_6528,N_5232,N_5154);
nand U6529 (N_6529,N_5228,N_5238);
nand U6530 (N_6530,N_5641,N_5048);
or U6531 (N_6531,N_5738,N_5132);
or U6532 (N_6532,N_5966,N_5312);
and U6533 (N_6533,N_5748,N_5385);
xnor U6534 (N_6534,N_5876,N_5786);
and U6535 (N_6535,N_5561,N_5921);
xor U6536 (N_6536,N_5673,N_5713);
nor U6537 (N_6537,N_5193,N_5127);
xnor U6538 (N_6538,N_5816,N_5307);
or U6539 (N_6539,N_5799,N_5605);
nor U6540 (N_6540,N_5002,N_5747);
or U6541 (N_6541,N_5118,N_5782);
nand U6542 (N_6542,N_5774,N_5288);
xor U6543 (N_6543,N_5646,N_5288);
and U6544 (N_6544,N_5023,N_5852);
and U6545 (N_6545,N_5730,N_5238);
or U6546 (N_6546,N_5876,N_5308);
nand U6547 (N_6547,N_5210,N_5579);
nor U6548 (N_6548,N_5450,N_5960);
nor U6549 (N_6549,N_5310,N_5116);
nor U6550 (N_6550,N_5777,N_5702);
xor U6551 (N_6551,N_5476,N_5461);
xor U6552 (N_6552,N_5385,N_5090);
xor U6553 (N_6553,N_5878,N_5064);
or U6554 (N_6554,N_5013,N_5114);
xor U6555 (N_6555,N_5525,N_5512);
nor U6556 (N_6556,N_5323,N_5355);
and U6557 (N_6557,N_5954,N_5579);
and U6558 (N_6558,N_5344,N_5917);
and U6559 (N_6559,N_5016,N_5931);
or U6560 (N_6560,N_5804,N_5336);
nand U6561 (N_6561,N_5955,N_5245);
nor U6562 (N_6562,N_5143,N_5261);
and U6563 (N_6563,N_5620,N_5386);
nand U6564 (N_6564,N_5493,N_5015);
nand U6565 (N_6565,N_5696,N_5379);
nor U6566 (N_6566,N_5118,N_5595);
or U6567 (N_6567,N_5047,N_5249);
and U6568 (N_6568,N_5122,N_5650);
xnor U6569 (N_6569,N_5912,N_5761);
xnor U6570 (N_6570,N_5140,N_5237);
or U6571 (N_6571,N_5015,N_5473);
nor U6572 (N_6572,N_5430,N_5122);
nand U6573 (N_6573,N_5137,N_5606);
nor U6574 (N_6574,N_5914,N_5571);
and U6575 (N_6575,N_5405,N_5433);
nand U6576 (N_6576,N_5872,N_5823);
and U6577 (N_6577,N_5017,N_5866);
nor U6578 (N_6578,N_5651,N_5521);
nor U6579 (N_6579,N_5556,N_5893);
nand U6580 (N_6580,N_5704,N_5194);
xor U6581 (N_6581,N_5161,N_5336);
and U6582 (N_6582,N_5049,N_5285);
or U6583 (N_6583,N_5883,N_5549);
or U6584 (N_6584,N_5191,N_5748);
or U6585 (N_6585,N_5229,N_5074);
nand U6586 (N_6586,N_5964,N_5990);
xor U6587 (N_6587,N_5001,N_5963);
and U6588 (N_6588,N_5182,N_5282);
or U6589 (N_6589,N_5705,N_5638);
nand U6590 (N_6590,N_5574,N_5676);
nand U6591 (N_6591,N_5468,N_5404);
nor U6592 (N_6592,N_5730,N_5107);
or U6593 (N_6593,N_5626,N_5177);
nand U6594 (N_6594,N_5625,N_5297);
and U6595 (N_6595,N_5911,N_5930);
and U6596 (N_6596,N_5492,N_5592);
xnor U6597 (N_6597,N_5703,N_5676);
xnor U6598 (N_6598,N_5612,N_5510);
nand U6599 (N_6599,N_5662,N_5464);
or U6600 (N_6600,N_5984,N_5180);
xnor U6601 (N_6601,N_5631,N_5687);
nor U6602 (N_6602,N_5502,N_5792);
xor U6603 (N_6603,N_5457,N_5362);
or U6604 (N_6604,N_5646,N_5403);
or U6605 (N_6605,N_5820,N_5747);
nor U6606 (N_6606,N_5924,N_5100);
and U6607 (N_6607,N_5880,N_5777);
nor U6608 (N_6608,N_5006,N_5960);
or U6609 (N_6609,N_5938,N_5985);
and U6610 (N_6610,N_5489,N_5108);
or U6611 (N_6611,N_5239,N_5281);
and U6612 (N_6612,N_5473,N_5415);
or U6613 (N_6613,N_5634,N_5092);
xor U6614 (N_6614,N_5924,N_5819);
nand U6615 (N_6615,N_5853,N_5653);
nor U6616 (N_6616,N_5986,N_5618);
xnor U6617 (N_6617,N_5122,N_5395);
nor U6618 (N_6618,N_5187,N_5122);
nor U6619 (N_6619,N_5478,N_5831);
xor U6620 (N_6620,N_5131,N_5442);
and U6621 (N_6621,N_5729,N_5754);
nor U6622 (N_6622,N_5142,N_5856);
and U6623 (N_6623,N_5913,N_5162);
nor U6624 (N_6624,N_5029,N_5487);
nor U6625 (N_6625,N_5555,N_5393);
xor U6626 (N_6626,N_5660,N_5308);
nor U6627 (N_6627,N_5729,N_5675);
and U6628 (N_6628,N_5211,N_5380);
xnor U6629 (N_6629,N_5169,N_5518);
and U6630 (N_6630,N_5919,N_5604);
nand U6631 (N_6631,N_5284,N_5843);
nand U6632 (N_6632,N_5519,N_5980);
and U6633 (N_6633,N_5946,N_5580);
and U6634 (N_6634,N_5013,N_5792);
nand U6635 (N_6635,N_5538,N_5296);
nor U6636 (N_6636,N_5285,N_5522);
and U6637 (N_6637,N_5027,N_5729);
nor U6638 (N_6638,N_5540,N_5611);
or U6639 (N_6639,N_5935,N_5191);
or U6640 (N_6640,N_5021,N_5589);
xnor U6641 (N_6641,N_5739,N_5816);
xor U6642 (N_6642,N_5512,N_5523);
xnor U6643 (N_6643,N_5627,N_5471);
and U6644 (N_6644,N_5979,N_5709);
and U6645 (N_6645,N_5592,N_5451);
nor U6646 (N_6646,N_5606,N_5009);
or U6647 (N_6647,N_5291,N_5789);
nor U6648 (N_6648,N_5294,N_5121);
nand U6649 (N_6649,N_5504,N_5482);
or U6650 (N_6650,N_5051,N_5337);
nand U6651 (N_6651,N_5371,N_5813);
nor U6652 (N_6652,N_5415,N_5374);
and U6653 (N_6653,N_5876,N_5393);
xnor U6654 (N_6654,N_5535,N_5861);
xor U6655 (N_6655,N_5673,N_5261);
and U6656 (N_6656,N_5991,N_5883);
and U6657 (N_6657,N_5797,N_5552);
nand U6658 (N_6658,N_5459,N_5617);
or U6659 (N_6659,N_5342,N_5249);
or U6660 (N_6660,N_5865,N_5800);
nand U6661 (N_6661,N_5126,N_5602);
or U6662 (N_6662,N_5500,N_5740);
xor U6663 (N_6663,N_5266,N_5009);
or U6664 (N_6664,N_5084,N_5436);
and U6665 (N_6665,N_5803,N_5585);
xor U6666 (N_6666,N_5485,N_5183);
nor U6667 (N_6667,N_5880,N_5267);
nor U6668 (N_6668,N_5349,N_5187);
or U6669 (N_6669,N_5448,N_5298);
xnor U6670 (N_6670,N_5391,N_5948);
nor U6671 (N_6671,N_5619,N_5426);
nor U6672 (N_6672,N_5645,N_5788);
or U6673 (N_6673,N_5895,N_5521);
and U6674 (N_6674,N_5114,N_5294);
xnor U6675 (N_6675,N_5671,N_5417);
nand U6676 (N_6676,N_5979,N_5007);
and U6677 (N_6677,N_5340,N_5134);
nor U6678 (N_6678,N_5149,N_5465);
and U6679 (N_6679,N_5869,N_5459);
nor U6680 (N_6680,N_5113,N_5332);
and U6681 (N_6681,N_5761,N_5851);
or U6682 (N_6682,N_5154,N_5672);
or U6683 (N_6683,N_5907,N_5790);
nor U6684 (N_6684,N_5022,N_5819);
and U6685 (N_6685,N_5537,N_5196);
xnor U6686 (N_6686,N_5573,N_5729);
and U6687 (N_6687,N_5865,N_5459);
nor U6688 (N_6688,N_5829,N_5099);
nor U6689 (N_6689,N_5731,N_5239);
or U6690 (N_6690,N_5805,N_5025);
or U6691 (N_6691,N_5894,N_5423);
and U6692 (N_6692,N_5870,N_5894);
xor U6693 (N_6693,N_5676,N_5031);
nand U6694 (N_6694,N_5159,N_5192);
nor U6695 (N_6695,N_5797,N_5360);
and U6696 (N_6696,N_5808,N_5978);
xnor U6697 (N_6697,N_5213,N_5000);
and U6698 (N_6698,N_5301,N_5134);
xnor U6699 (N_6699,N_5456,N_5807);
or U6700 (N_6700,N_5979,N_5240);
or U6701 (N_6701,N_5707,N_5383);
xnor U6702 (N_6702,N_5969,N_5216);
and U6703 (N_6703,N_5121,N_5316);
nor U6704 (N_6704,N_5385,N_5998);
or U6705 (N_6705,N_5141,N_5572);
and U6706 (N_6706,N_5486,N_5671);
and U6707 (N_6707,N_5518,N_5038);
nor U6708 (N_6708,N_5932,N_5437);
xnor U6709 (N_6709,N_5083,N_5268);
xor U6710 (N_6710,N_5312,N_5511);
or U6711 (N_6711,N_5726,N_5095);
and U6712 (N_6712,N_5473,N_5046);
nand U6713 (N_6713,N_5034,N_5799);
nand U6714 (N_6714,N_5126,N_5296);
nor U6715 (N_6715,N_5030,N_5876);
xnor U6716 (N_6716,N_5289,N_5347);
nor U6717 (N_6717,N_5326,N_5559);
nor U6718 (N_6718,N_5013,N_5952);
nand U6719 (N_6719,N_5912,N_5194);
nand U6720 (N_6720,N_5273,N_5952);
xor U6721 (N_6721,N_5667,N_5911);
xor U6722 (N_6722,N_5493,N_5342);
nand U6723 (N_6723,N_5724,N_5972);
and U6724 (N_6724,N_5699,N_5797);
and U6725 (N_6725,N_5387,N_5428);
or U6726 (N_6726,N_5953,N_5966);
or U6727 (N_6727,N_5592,N_5652);
or U6728 (N_6728,N_5585,N_5120);
or U6729 (N_6729,N_5284,N_5224);
and U6730 (N_6730,N_5437,N_5912);
xor U6731 (N_6731,N_5239,N_5070);
nand U6732 (N_6732,N_5101,N_5770);
or U6733 (N_6733,N_5103,N_5676);
nor U6734 (N_6734,N_5490,N_5864);
xnor U6735 (N_6735,N_5720,N_5820);
nor U6736 (N_6736,N_5943,N_5849);
nor U6737 (N_6737,N_5341,N_5907);
or U6738 (N_6738,N_5813,N_5118);
xor U6739 (N_6739,N_5659,N_5276);
or U6740 (N_6740,N_5489,N_5989);
nor U6741 (N_6741,N_5884,N_5048);
nand U6742 (N_6742,N_5665,N_5018);
nor U6743 (N_6743,N_5579,N_5093);
nor U6744 (N_6744,N_5519,N_5082);
and U6745 (N_6745,N_5075,N_5671);
or U6746 (N_6746,N_5929,N_5397);
nor U6747 (N_6747,N_5457,N_5623);
xnor U6748 (N_6748,N_5786,N_5306);
and U6749 (N_6749,N_5223,N_5938);
nand U6750 (N_6750,N_5160,N_5718);
nor U6751 (N_6751,N_5525,N_5288);
and U6752 (N_6752,N_5733,N_5480);
nor U6753 (N_6753,N_5402,N_5673);
nor U6754 (N_6754,N_5967,N_5460);
nand U6755 (N_6755,N_5018,N_5682);
and U6756 (N_6756,N_5830,N_5295);
nand U6757 (N_6757,N_5548,N_5072);
nand U6758 (N_6758,N_5757,N_5308);
nand U6759 (N_6759,N_5037,N_5398);
or U6760 (N_6760,N_5465,N_5794);
nand U6761 (N_6761,N_5415,N_5576);
or U6762 (N_6762,N_5654,N_5829);
or U6763 (N_6763,N_5501,N_5296);
nor U6764 (N_6764,N_5830,N_5885);
nand U6765 (N_6765,N_5326,N_5166);
nor U6766 (N_6766,N_5467,N_5272);
nand U6767 (N_6767,N_5147,N_5638);
and U6768 (N_6768,N_5401,N_5834);
and U6769 (N_6769,N_5709,N_5159);
nand U6770 (N_6770,N_5606,N_5551);
or U6771 (N_6771,N_5117,N_5668);
and U6772 (N_6772,N_5968,N_5460);
or U6773 (N_6773,N_5634,N_5894);
nand U6774 (N_6774,N_5837,N_5808);
nand U6775 (N_6775,N_5261,N_5626);
and U6776 (N_6776,N_5897,N_5156);
xor U6777 (N_6777,N_5770,N_5277);
or U6778 (N_6778,N_5393,N_5927);
nor U6779 (N_6779,N_5390,N_5629);
or U6780 (N_6780,N_5438,N_5607);
nor U6781 (N_6781,N_5010,N_5342);
xnor U6782 (N_6782,N_5839,N_5473);
or U6783 (N_6783,N_5442,N_5677);
xnor U6784 (N_6784,N_5817,N_5975);
xor U6785 (N_6785,N_5370,N_5452);
and U6786 (N_6786,N_5511,N_5894);
or U6787 (N_6787,N_5235,N_5982);
nand U6788 (N_6788,N_5295,N_5238);
nor U6789 (N_6789,N_5357,N_5349);
and U6790 (N_6790,N_5665,N_5556);
nor U6791 (N_6791,N_5417,N_5048);
or U6792 (N_6792,N_5201,N_5484);
and U6793 (N_6793,N_5926,N_5443);
nor U6794 (N_6794,N_5227,N_5486);
nor U6795 (N_6795,N_5446,N_5423);
and U6796 (N_6796,N_5063,N_5867);
or U6797 (N_6797,N_5150,N_5905);
xnor U6798 (N_6798,N_5855,N_5378);
nor U6799 (N_6799,N_5974,N_5291);
or U6800 (N_6800,N_5199,N_5996);
and U6801 (N_6801,N_5598,N_5313);
and U6802 (N_6802,N_5423,N_5553);
or U6803 (N_6803,N_5275,N_5950);
and U6804 (N_6804,N_5104,N_5649);
and U6805 (N_6805,N_5769,N_5497);
xnor U6806 (N_6806,N_5867,N_5706);
and U6807 (N_6807,N_5961,N_5881);
and U6808 (N_6808,N_5735,N_5393);
and U6809 (N_6809,N_5304,N_5836);
xnor U6810 (N_6810,N_5538,N_5058);
or U6811 (N_6811,N_5500,N_5743);
nor U6812 (N_6812,N_5422,N_5236);
xnor U6813 (N_6813,N_5811,N_5059);
xnor U6814 (N_6814,N_5304,N_5380);
and U6815 (N_6815,N_5147,N_5419);
nand U6816 (N_6816,N_5599,N_5611);
nor U6817 (N_6817,N_5874,N_5796);
and U6818 (N_6818,N_5708,N_5896);
and U6819 (N_6819,N_5439,N_5632);
nand U6820 (N_6820,N_5749,N_5383);
nor U6821 (N_6821,N_5782,N_5186);
or U6822 (N_6822,N_5126,N_5133);
nand U6823 (N_6823,N_5335,N_5184);
nand U6824 (N_6824,N_5081,N_5992);
or U6825 (N_6825,N_5524,N_5240);
nand U6826 (N_6826,N_5465,N_5260);
or U6827 (N_6827,N_5537,N_5143);
nand U6828 (N_6828,N_5365,N_5568);
nor U6829 (N_6829,N_5234,N_5823);
xnor U6830 (N_6830,N_5331,N_5134);
or U6831 (N_6831,N_5386,N_5076);
nand U6832 (N_6832,N_5070,N_5858);
nand U6833 (N_6833,N_5183,N_5788);
or U6834 (N_6834,N_5840,N_5145);
nor U6835 (N_6835,N_5013,N_5958);
xnor U6836 (N_6836,N_5181,N_5232);
xor U6837 (N_6837,N_5371,N_5996);
and U6838 (N_6838,N_5142,N_5259);
or U6839 (N_6839,N_5965,N_5544);
nand U6840 (N_6840,N_5264,N_5874);
and U6841 (N_6841,N_5028,N_5820);
and U6842 (N_6842,N_5123,N_5275);
xnor U6843 (N_6843,N_5929,N_5131);
or U6844 (N_6844,N_5622,N_5683);
xor U6845 (N_6845,N_5543,N_5831);
and U6846 (N_6846,N_5335,N_5669);
xor U6847 (N_6847,N_5394,N_5772);
nor U6848 (N_6848,N_5726,N_5944);
xnor U6849 (N_6849,N_5332,N_5844);
nand U6850 (N_6850,N_5950,N_5816);
and U6851 (N_6851,N_5890,N_5068);
nor U6852 (N_6852,N_5595,N_5589);
nand U6853 (N_6853,N_5895,N_5896);
nand U6854 (N_6854,N_5406,N_5652);
or U6855 (N_6855,N_5343,N_5628);
and U6856 (N_6856,N_5973,N_5783);
xor U6857 (N_6857,N_5735,N_5291);
and U6858 (N_6858,N_5491,N_5485);
xor U6859 (N_6859,N_5106,N_5509);
nor U6860 (N_6860,N_5979,N_5158);
and U6861 (N_6861,N_5475,N_5972);
and U6862 (N_6862,N_5573,N_5915);
nor U6863 (N_6863,N_5958,N_5621);
nor U6864 (N_6864,N_5599,N_5134);
xnor U6865 (N_6865,N_5642,N_5923);
nand U6866 (N_6866,N_5468,N_5375);
nor U6867 (N_6867,N_5511,N_5399);
nand U6868 (N_6868,N_5749,N_5350);
nor U6869 (N_6869,N_5661,N_5907);
or U6870 (N_6870,N_5756,N_5903);
nor U6871 (N_6871,N_5607,N_5909);
nor U6872 (N_6872,N_5588,N_5023);
xor U6873 (N_6873,N_5402,N_5366);
and U6874 (N_6874,N_5576,N_5568);
nand U6875 (N_6875,N_5312,N_5415);
xor U6876 (N_6876,N_5827,N_5083);
or U6877 (N_6877,N_5544,N_5773);
and U6878 (N_6878,N_5055,N_5743);
nand U6879 (N_6879,N_5173,N_5728);
or U6880 (N_6880,N_5821,N_5913);
nor U6881 (N_6881,N_5392,N_5496);
or U6882 (N_6882,N_5254,N_5603);
or U6883 (N_6883,N_5870,N_5546);
nor U6884 (N_6884,N_5252,N_5677);
nand U6885 (N_6885,N_5787,N_5335);
xnor U6886 (N_6886,N_5225,N_5559);
or U6887 (N_6887,N_5004,N_5910);
nor U6888 (N_6888,N_5782,N_5729);
nand U6889 (N_6889,N_5175,N_5622);
nor U6890 (N_6890,N_5938,N_5628);
or U6891 (N_6891,N_5979,N_5449);
xnor U6892 (N_6892,N_5803,N_5116);
xor U6893 (N_6893,N_5399,N_5515);
nor U6894 (N_6894,N_5691,N_5283);
xnor U6895 (N_6895,N_5715,N_5287);
or U6896 (N_6896,N_5375,N_5568);
or U6897 (N_6897,N_5839,N_5968);
nand U6898 (N_6898,N_5749,N_5853);
and U6899 (N_6899,N_5841,N_5234);
and U6900 (N_6900,N_5655,N_5400);
and U6901 (N_6901,N_5006,N_5368);
nor U6902 (N_6902,N_5819,N_5455);
nand U6903 (N_6903,N_5543,N_5963);
or U6904 (N_6904,N_5341,N_5964);
xnor U6905 (N_6905,N_5662,N_5039);
nor U6906 (N_6906,N_5296,N_5268);
and U6907 (N_6907,N_5893,N_5832);
xor U6908 (N_6908,N_5975,N_5368);
xnor U6909 (N_6909,N_5193,N_5660);
nand U6910 (N_6910,N_5971,N_5668);
and U6911 (N_6911,N_5283,N_5429);
nor U6912 (N_6912,N_5419,N_5468);
nor U6913 (N_6913,N_5852,N_5482);
and U6914 (N_6914,N_5275,N_5287);
xnor U6915 (N_6915,N_5399,N_5698);
xor U6916 (N_6916,N_5464,N_5419);
and U6917 (N_6917,N_5612,N_5702);
nor U6918 (N_6918,N_5666,N_5419);
nor U6919 (N_6919,N_5856,N_5897);
or U6920 (N_6920,N_5509,N_5942);
nor U6921 (N_6921,N_5419,N_5390);
nor U6922 (N_6922,N_5870,N_5823);
and U6923 (N_6923,N_5780,N_5382);
nand U6924 (N_6924,N_5523,N_5070);
or U6925 (N_6925,N_5883,N_5908);
nand U6926 (N_6926,N_5422,N_5026);
nand U6927 (N_6927,N_5457,N_5870);
and U6928 (N_6928,N_5742,N_5474);
nand U6929 (N_6929,N_5286,N_5491);
xor U6930 (N_6930,N_5374,N_5669);
and U6931 (N_6931,N_5583,N_5150);
or U6932 (N_6932,N_5753,N_5590);
nand U6933 (N_6933,N_5801,N_5546);
nand U6934 (N_6934,N_5083,N_5426);
or U6935 (N_6935,N_5917,N_5706);
nor U6936 (N_6936,N_5507,N_5750);
xnor U6937 (N_6937,N_5079,N_5407);
nor U6938 (N_6938,N_5789,N_5127);
nor U6939 (N_6939,N_5655,N_5318);
nand U6940 (N_6940,N_5739,N_5770);
or U6941 (N_6941,N_5184,N_5960);
and U6942 (N_6942,N_5604,N_5940);
or U6943 (N_6943,N_5871,N_5876);
xnor U6944 (N_6944,N_5789,N_5152);
and U6945 (N_6945,N_5543,N_5172);
nand U6946 (N_6946,N_5786,N_5765);
nand U6947 (N_6947,N_5567,N_5127);
xnor U6948 (N_6948,N_5276,N_5985);
nand U6949 (N_6949,N_5979,N_5575);
or U6950 (N_6950,N_5784,N_5557);
xor U6951 (N_6951,N_5572,N_5254);
and U6952 (N_6952,N_5944,N_5577);
or U6953 (N_6953,N_5330,N_5022);
or U6954 (N_6954,N_5244,N_5783);
and U6955 (N_6955,N_5055,N_5999);
xor U6956 (N_6956,N_5946,N_5300);
nor U6957 (N_6957,N_5840,N_5539);
nand U6958 (N_6958,N_5502,N_5198);
xor U6959 (N_6959,N_5436,N_5991);
and U6960 (N_6960,N_5218,N_5897);
or U6961 (N_6961,N_5596,N_5653);
xnor U6962 (N_6962,N_5956,N_5471);
nand U6963 (N_6963,N_5235,N_5699);
nand U6964 (N_6964,N_5357,N_5841);
nand U6965 (N_6965,N_5386,N_5264);
xnor U6966 (N_6966,N_5278,N_5898);
nor U6967 (N_6967,N_5430,N_5137);
or U6968 (N_6968,N_5548,N_5486);
xnor U6969 (N_6969,N_5364,N_5837);
or U6970 (N_6970,N_5575,N_5655);
or U6971 (N_6971,N_5737,N_5578);
or U6972 (N_6972,N_5827,N_5926);
or U6973 (N_6973,N_5569,N_5104);
nor U6974 (N_6974,N_5511,N_5143);
nor U6975 (N_6975,N_5798,N_5324);
or U6976 (N_6976,N_5092,N_5028);
or U6977 (N_6977,N_5480,N_5039);
or U6978 (N_6978,N_5217,N_5023);
nor U6979 (N_6979,N_5779,N_5556);
and U6980 (N_6980,N_5434,N_5148);
nand U6981 (N_6981,N_5350,N_5440);
nand U6982 (N_6982,N_5932,N_5366);
nand U6983 (N_6983,N_5272,N_5045);
xnor U6984 (N_6984,N_5541,N_5278);
or U6985 (N_6985,N_5127,N_5436);
and U6986 (N_6986,N_5566,N_5632);
xnor U6987 (N_6987,N_5489,N_5062);
xor U6988 (N_6988,N_5461,N_5622);
nand U6989 (N_6989,N_5407,N_5134);
or U6990 (N_6990,N_5784,N_5695);
nand U6991 (N_6991,N_5116,N_5671);
nor U6992 (N_6992,N_5915,N_5364);
and U6993 (N_6993,N_5962,N_5673);
nor U6994 (N_6994,N_5537,N_5504);
xnor U6995 (N_6995,N_5137,N_5251);
and U6996 (N_6996,N_5939,N_5743);
xnor U6997 (N_6997,N_5881,N_5365);
and U6998 (N_6998,N_5177,N_5554);
nand U6999 (N_6999,N_5370,N_5754);
nor U7000 (N_7000,N_6638,N_6324);
and U7001 (N_7001,N_6276,N_6826);
and U7002 (N_7002,N_6146,N_6740);
nand U7003 (N_7003,N_6603,N_6992);
nand U7004 (N_7004,N_6148,N_6670);
or U7005 (N_7005,N_6341,N_6389);
nand U7006 (N_7006,N_6084,N_6766);
xnor U7007 (N_7007,N_6073,N_6683);
nor U7008 (N_7008,N_6125,N_6921);
nand U7009 (N_7009,N_6449,N_6380);
xnor U7010 (N_7010,N_6281,N_6506);
nand U7011 (N_7011,N_6106,N_6785);
xor U7012 (N_7012,N_6623,N_6953);
or U7013 (N_7013,N_6120,N_6864);
and U7014 (N_7014,N_6450,N_6868);
and U7015 (N_7015,N_6107,N_6536);
or U7016 (N_7016,N_6489,N_6105);
nand U7017 (N_7017,N_6233,N_6198);
or U7018 (N_7018,N_6734,N_6203);
nand U7019 (N_7019,N_6156,N_6566);
and U7020 (N_7020,N_6798,N_6141);
nor U7021 (N_7021,N_6033,N_6978);
and U7022 (N_7022,N_6304,N_6279);
and U7023 (N_7023,N_6849,N_6537);
nor U7024 (N_7024,N_6460,N_6250);
nor U7025 (N_7025,N_6297,N_6760);
and U7026 (N_7026,N_6694,N_6583);
or U7027 (N_7027,N_6815,N_6201);
nor U7028 (N_7028,N_6699,N_6172);
and U7029 (N_7029,N_6104,N_6322);
nand U7030 (N_7030,N_6021,N_6923);
and U7031 (N_7031,N_6856,N_6754);
nand U7032 (N_7032,N_6966,N_6695);
or U7033 (N_7033,N_6735,N_6876);
xor U7034 (N_7034,N_6432,N_6543);
nor U7035 (N_7035,N_6689,N_6692);
and U7036 (N_7036,N_6265,N_6729);
xor U7037 (N_7037,N_6244,N_6257);
xnor U7038 (N_7038,N_6679,N_6716);
or U7039 (N_7039,N_6581,N_6578);
nor U7040 (N_7040,N_6420,N_6762);
and U7041 (N_7041,N_6841,N_6122);
or U7042 (N_7042,N_6743,N_6527);
nand U7043 (N_7043,N_6775,N_6852);
and U7044 (N_7044,N_6645,N_6666);
xor U7045 (N_7045,N_6379,N_6182);
nand U7046 (N_7046,N_6837,N_6941);
xnor U7047 (N_7047,N_6544,N_6491);
xnor U7048 (N_7048,N_6660,N_6056);
and U7049 (N_7049,N_6354,N_6686);
nor U7050 (N_7050,N_6626,N_6300);
or U7051 (N_7051,N_6569,N_6005);
or U7052 (N_7052,N_6907,N_6671);
and U7053 (N_7053,N_6816,N_6616);
nand U7054 (N_7054,N_6091,N_6865);
xor U7055 (N_7055,N_6863,N_6443);
and U7056 (N_7056,N_6565,N_6522);
and U7057 (N_7057,N_6222,N_6625);
nor U7058 (N_7058,N_6412,N_6903);
nand U7059 (N_7059,N_6758,N_6594);
and U7060 (N_7060,N_6405,N_6121);
or U7061 (N_7061,N_6805,N_6790);
nand U7062 (N_7062,N_6756,N_6060);
and U7063 (N_7063,N_6009,N_6458);
nand U7064 (N_7064,N_6482,N_6969);
and U7065 (N_7065,N_6211,N_6497);
nand U7066 (N_7066,N_6045,N_6847);
and U7067 (N_7067,N_6440,N_6610);
nor U7068 (N_7068,N_6368,N_6499);
nor U7069 (N_7069,N_6183,N_6696);
and U7070 (N_7070,N_6930,N_6363);
xor U7071 (N_7071,N_6472,N_6398);
nand U7072 (N_7072,N_6212,N_6653);
nand U7073 (N_7073,N_6526,N_6076);
nand U7074 (N_7074,N_6051,N_6628);
xor U7075 (N_7075,N_6905,N_6476);
nor U7076 (N_7076,N_6285,N_6874);
nand U7077 (N_7077,N_6192,N_6587);
nand U7078 (N_7078,N_6187,N_6232);
nand U7079 (N_7079,N_6801,N_6913);
nand U7080 (N_7080,N_6654,N_6888);
or U7081 (N_7081,N_6908,N_6361);
nor U7082 (N_7082,N_6596,N_6438);
and U7083 (N_7083,N_6977,N_6800);
nor U7084 (N_7084,N_6755,N_6474);
or U7085 (N_7085,N_6889,N_6316);
xor U7086 (N_7086,N_6485,N_6226);
nand U7087 (N_7087,N_6242,N_6964);
xnor U7088 (N_7088,N_6131,N_6000);
nor U7089 (N_7089,N_6306,N_6983);
and U7090 (N_7090,N_6809,N_6554);
and U7091 (N_7091,N_6912,N_6077);
xnor U7092 (N_7092,N_6325,N_6965);
nand U7093 (N_7093,N_6159,N_6832);
or U7094 (N_7094,N_6987,N_6188);
xnor U7095 (N_7095,N_6402,N_6821);
xnor U7096 (N_7096,N_6410,N_6417);
or U7097 (N_7097,N_6378,N_6372);
or U7098 (N_7098,N_6280,N_6083);
or U7099 (N_7099,N_6600,N_6627);
and U7100 (N_7100,N_6041,N_6990);
xor U7101 (N_7101,N_6003,N_6513);
nor U7102 (N_7102,N_6687,N_6020);
xor U7103 (N_7103,N_6524,N_6481);
or U7104 (N_7104,N_6910,N_6066);
or U7105 (N_7105,N_6563,N_6215);
and U7106 (N_7106,N_6100,N_6980);
nand U7107 (N_7107,N_6911,N_6113);
nand U7108 (N_7108,N_6640,N_6011);
nand U7109 (N_7109,N_6468,N_6328);
or U7110 (N_7110,N_6291,N_6124);
nand U7111 (N_7111,N_6437,N_6512);
or U7112 (N_7112,N_6193,N_6168);
and U7113 (N_7113,N_6480,N_6646);
and U7114 (N_7114,N_6312,N_6181);
nor U7115 (N_7115,N_6890,N_6311);
nor U7116 (N_7116,N_6882,N_6757);
nor U7117 (N_7117,N_6797,N_6326);
and U7118 (N_7118,N_6254,N_6031);
nor U7119 (N_7119,N_6200,N_6597);
and U7120 (N_7120,N_6961,N_6118);
or U7121 (N_7121,N_6715,N_6099);
and U7122 (N_7122,N_6338,N_6278);
or U7123 (N_7123,N_6949,N_6299);
nand U7124 (N_7124,N_6724,N_6958);
or U7125 (N_7125,N_6772,N_6708);
or U7126 (N_7126,N_6477,N_6598);
nor U7127 (N_7127,N_6317,N_6516);
and U7128 (N_7128,N_6137,N_6605);
xnor U7129 (N_7129,N_6142,N_6749);
and U7130 (N_7130,N_6658,N_6162);
or U7131 (N_7131,N_6768,N_6942);
nor U7132 (N_7132,N_6274,N_6109);
and U7133 (N_7133,N_6843,N_6639);
or U7134 (N_7134,N_6602,N_6519);
and U7135 (N_7135,N_6424,N_6469);
or U7136 (N_7136,N_6520,N_6415);
or U7137 (N_7137,N_6404,N_6675);
nor U7138 (N_7138,N_6691,N_6240);
or U7139 (N_7139,N_6582,N_6238);
and U7140 (N_7140,N_6834,N_6272);
nor U7141 (N_7141,N_6169,N_6887);
nor U7142 (N_7142,N_6089,N_6848);
and U7143 (N_7143,N_6585,N_6776);
nand U7144 (N_7144,N_6221,N_6838);
and U7145 (N_7145,N_6777,N_6769);
nor U7146 (N_7146,N_6062,N_6705);
and U7147 (N_7147,N_6688,N_6016);
nand U7148 (N_7148,N_6057,N_6343);
nor U7149 (N_7149,N_6008,N_6642);
xnor U7150 (N_7150,N_6262,N_6377);
or U7151 (N_7151,N_6013,N_6676);
xor U7152 (N_7152,N_6258,N_6134);
or U7153 (N_7153,N_6737,N_6150);
or U7154 (N_7154,N_6473,N_6032);
or U7155 (N_7155,N_6668,N_6487);
or U7156 (N_7156,N_6984,N_6535);
or U7157 (N_7157,N_6557,N_6534);
nor U7158 (N_7158,N_6080,N_6919);
or U7159 (N_7159,N_6929,N_6701);
nand U7160 (N_7160,N_6647,N_6508);
xor U7161 (N_7161,N_6390,N_6173);
or U7162 (N_7162,N_6738,N_6770);
nand U7163 (N_7163,N_6560,N_6962);
nor U7164 (N_7164,N_6446,N_6661);
or U7165 (N_7165,N_6822,N_6096);
nand U7166 (N_7166,N_6103,N_6733);
xnor U7167 (N_7167,N_6224,N_6877);
or U7168 (N_7168,N_6589,N_6902);
nand U7169 (N_7169,N_6720,N_6901);
xnor U7170 (N_7170,N_6808,N_6176);
xnor U7171 (N_7171,N_6622,N_6027);
or U7172 (N_7172,N_6464,N_6972);
nand U7173 (N_7173,N_6550,N_6213);
nand U7174 (N_7174,N_6664,N_6730);
and U7175 (N_7175,N_6164,N_6988);
nor U7176 (N_7176,N_6175,N_6456);
xnor U7177 (N_7177,N_6936,N_6995);
nand U7178 (N_7178,N_6548,N_6712);
nor U7179 (N_7179,N_6028,N_6145);
xor U7180 (N_7180,N_6951,N_6305);
or U7181 (N_7181,N_6358,N_6985);
nand U7182 (N_7182,N_6086,N_6523);
nand U7183 (N_7183,N_6078,N_6861);
xnor U7184 (N_7184,N_6117,N_6154);
and U7185 (N_7185,N_6531,N_6742);
and U7186 (N_7186,N_6619,N_6228);
xor U7187 (N_7187,N_6167,N_6196);
nand U7188 (N_7188,N_6891,N_6039);
or U7189 (N_7189,N_6824,N_6851);
nand U7190 (N_7190,N_6401,N_6067);
nor U7191 (N_7191,N_6759,N_6894);
nor U7192 (N_7192,N_6436,N_6165);
or U7193 (N_7193,N_6806,N_6239);
or U7194 (N_7194,N_6726,N_6747);
and U7195 (N_7195,N_6095,N_6636);
nand U7196 (N_7196,N_6088,N_6723);
xnor U7197 (N_7197,N_6502,N_6204);
or U7198 (N_7198,N_6765,N_6553);
and U7199 (N_7199,N_6425,N_6518);
nor U7200 (N_7200,N_6706,N_6914);
and U7201 (N_7201,N_6385,N_6267);
xnor U7202 (N_7202,N_6624,N_6371);
or U7203 (N_7203,N_6273,N_6245);
nand U7204 (N_7204,N_6799,N_6116);
nor U7205 (N_7205,N_6320,N_6064);
nor U7206 (N_7206,N_6043,N_6703);
xor U7207 (N_7207,N_6321,N_6471);
nand U7208 (N_7208,N_6023,N_6869);
and U7209 (N_7209,N_6549,N_6875);
or U7210 (N_7210,N_6132,N_6042);
nor U7211 (N_7211,N_6301,N_6793);
or U7212 (N_7212,N_6677,N_6879);
nor U7213 (N_7213,N_6383,N_6633);
nand U7214 (N_7214,N_6270,N_6794);
and U7215 (N_7215,N_6422,N_6959);
and U7216 (N_7216,N_6917,N_6922);
xnor U7217 (N_7217,N_6857,N_6573);
nor U7218 (N_7218,N_6050,N_6135);
and U7219 (N_7219,N_6955,N_6202);
and U7220 (N_7220,N_6909,N_6867);
xnor U7221 (N_7221,N_6503,N_6199);
nand U7222 (N_7222,N_6058,N_6356);
nand U7223 (N_7223,N_6157,N_6496);
and U7224 (N_7224,N_6982,N_6463);
and U7225 (N_7225,N_6210,N_6128);
nor U7226 (N_7226,N_6556,N_6219);
or U7227 (N_7227,N_6376,N_6344);
nand U7228 (N_7228,N_6810,N_6348);
xor U7229 (N_7229,N_6457,N_6746);
or U7230 (N_7230,N_6085,N_6813);
nand U7231 (N_7231,N_6916,N_6643);
xor U7232 (N_7232,N_6564,N_6359);
nor U7233 (N_7233,N_6830,N_6880);
nand U7234 (N_7234,N_6214,N_6467);
or U7235 (N_7235,N_6858,N_6697);
nor U7236 (N_7236,N_6353,N_6030);
and U7237 (N_7237,N_6840,N_6260);
or U7238 (N_7238,N_6571,N_6345);
xor U7239 (N_7239,N_6026,N_6998);
or U7240 (N_7240,N_6352,N_6391);
xor U7241 (N_7241,N_6652,N_6539);
xnor U7242 (N_7242,N_6483,N_6786);
and U7243 (N_7243,N_6866,N_6490);
and U7244 (N_7244,N_6022,N_6119);
and U7245 (N_7245,N_6590,N_6528);
nand U7246 (N_7246,N_6933,N_6433);
or U7247 (N_7247,N_6246,N_6349);
xor U7248 (N_7248,N_6384,N_6374);
or U7249 (N_7249,N_6362,N_6814);
or U7250 (N_7250,N_6938,N_6672);
nand U7251 (N_7251,N_6466,N_6323);
nor U7252 (N_7252,N_6409,N_6659);
nand U7253 (N_7253,N_6403,N_6006);
or U7254 (N_7254,N_6515,N_6546);
xnor U7255 (N_7255,N_6632,N_6991);
and U7256 (N_7256,N_6595,N_6063);
and U7257 (N_7257,N_6835,N_6782);
xor U7258 (N_7258,N_6225,N_6993);
nand U7259 (N_7259,N_6753,N_6558);
nor U7260 (N_7260,N_6130,N_6140);
or U7261 (N_7261,N_6504,N_6327);
or U7262 (N_7262,N_6094,N_6828);
nand U7263 (N_7263,N_6126,N_6494);
or U7264 (N_7264,N_6829,N_6388);
or U7265 (N_7265,N_6657,N_6495);
nor U7266 (N_7266,N_6364,N_6722);
xnor U7267 (N_7267,N_6484,N_6637);
nor U7268 (N_7268,N_6997,N_6387);
nand U7269 (N_7269,N_6873,N_6714);
or U7270 (N_7270,N_6631,N_6400);
or U7271 (N_7271,N_6307,N_6957);
and U7272 (N_7272,N_6186,N_6773);
and U7273 (N_7273,N_6313,N_6570);
nor U7274 (N_7274,N_6802,N_6396);
and U7275 (N_7275,N_6920,N_6408);
and U7276 (N_7276,N_6360,N_6454);
and U7277 (N_7277,N_6872,N_6711);
and U7278 (N_7278,N_6673,N_6897);
and U7279 (N_7279,N_6634,N_6071);
nor U7280 (N_7280,N_6110,N_6399);
nand U7281 (N_7281,N_6207,N_6842);
and U7282 (N_7282,N_6330,N_6604);
xor U7283 (N_7283,N_6470,N_6235);
xor U7284 (N_7284,N_6255,N_6540);
nand U7285 (N_7285,N_6833,N_6347);
nand U7286 (N_7286,N_6074,N_6034);
nand U7287 (N_7287,N_6994,N_6611);
and U7288 (N_7288,N_6937,N_6092);
and U7289 (N_7289,N_6309,N_6895);
nor U7290 (N_7290,N_6139,N_6748);
and U7291 (N_7291,N_6771,N_6745);
xnor U7292 (N_7292,N_6217,N_6445);
and U7293 (N_7293,N_6447,N_6068);
nand U7294 (N_7294,N_6241,N_6599);
xor U7295 (N_7295,N_6789,N_6684);
nor U7296 (N_7296,N_6682,N_6788);
or U7297 (N_7297,N_6944,N_6236);
and U7298 (N_7298,N_6151,N_6451);
or U7299 (N_7299,N_6514,N_6606);
or U7300 (N_7300,N_6205,N_6819);
or U7301 (N_7301,N_6946,N_6862);
or U7302 (N_7302,N_6049,N_6690);
or U7303 (N_7303,N_6663,N_6114);
xnor U7304 (N_7304,N_6845,N_6259);
or U7305 (N_7305,N_6886,N_6541);
or U7306 (N_7306,N_6855,N_6780);
xor U7307 (N_7307,N_6973,N_6426);
or U7308 (N_7308,N_6906,N_6488);
xor U7309 (N_7309,N_6700,N_6040);
or U7310 (N_7310,N_6635,N_6532);
xor U7311 (N_7311,N_6138,N_6655);
or U7312 (N_7312,N_6918,N_6015);
nand U7313 (N_7313,N_6956,N_6069);
nor U7314 (N_7314,N_6898,N_6542);
xnor U7315 (N_7315,N_6266,N_6435);
and U7316 (N_7316,N_6282,N_6791);
or U7317 (N_7317,N_6601,N_6588);
nor U7318 (N_7318,N_6247,N_6029);
nor U7319 (N_7319,N_6072,N_6248);
nand U7320 (N_7320,N_6044,N_6434);
and U7321 (N_7321,N_6174,N_6112);
or U7322 (N_7322,N_6333,N_6620);
nand U7323 (N_7323,N_6665,N_6795);
nand U7324 (N_7324,N_6413,N_6237);
nand U7325 (N_7325,N_6047,N_6098);
nor U7326 (N_7326,N_6761,N_6899);
and U7327 (N_7327,N_6411,N_6195);
and U7328 (N_7328,N_6284,N_6249);
and U7329 (N_7329,N_6290,N_6739);
xor U7330 (N_7330,N_6394,N_6303);
or U7331 (N_7331,N_6613,N_6179);
nand U7332 (N_7332,N_6346,N_6271);
and U7333 (N_7333,N_6498,N_6896);
nor U7334 (N_7334,N_6302,N_6319);
and U7335 (N_7335,N_6155,N_6289);
nor U7336 (N_7336,N_6823,N_6976);
xnor U7337 (N_7337,N_6669,N_6817);
xor U7338 (N_7338,N_6461,N_6406);
or U7339 (N_7339,N_6101,N_6996);
nor U7340 (N_7340,N_6693,N_6803);
nor U7341 (N_7341,N_6885,N_6779);
and U7342 (N_7342,N_6732,N_6521);
or U7343 (N_7343,N_6243,N_6418);
and U7344 (N_7344,N_6967,N_6392);
and U7345 (N_7345,N_6763,N_6796);
xor U7346 (N_7346,N_6059,N_6648);
or U7347 (N_7347,N_6630,N_6629);
nor U7348 (N_7348,N_6681,N_6575);
nor U7349 (N_7349,N_6475,N_6315);
nand U7350 (N_7350,N_6427,N_6012);
or U7351 (N_7351,N_6999,N_6048);
xnor U7352 (N_7352,N_6678,N_6430);
nor U7353 (N_7353,N_6053,N_6839);
xnor U7354 (N_7354,N_6736,N_6334);
and U7355 (N_7355,N_6925,N_6774);
nor U7356 (N_7356,N_6781,N_6052);
and U7357 (N_7357,N_6416,N_6778);
or U7358 (N_7358,N_6455,N_6567);
nor U7359 (N_7359,N_6293,N_6509);
or U7360 (N_7360,N_6511,N_6900);
nand U7361 (N_7361,N_6127,N_6337);
nor U7362 (N_7362,N_6807,N_6717);
nand U7363 (N_7363,N_6952,N_6492);
or U7364 (N_7364,N_6728,N_6707);
or U7365 (N_7365,N_6950,N_6428);
xor U7366 (N_7366,N_6336,N_6024);
xor U7367 (N_7367,N_6442,N_6256);
and U7368 (N_7368,N_6342,N_6375);
nand U7369 (N_7369,N_6892,N_6986);
xor U7370 (N_7370,N_6932,N_6178);
and U7371 (N_7371,N_6097,N_6915);
or U7372 (N_7372,N_6552,N_6340);
and U7373 (N_7373,N_6584,N_6180);
nor U7374 (N_7374,N_6161,N_6968);
nor U7375 (N_7375,N_6268,N_6357);
or U7376 (N_7376,N_6517,N_6505);
or U7377 (N_7377,N_6818,N_6975);
nand U7378 (N_7378,N_6081,N_6744);
or U7379 (N_7379,N_6355,N_6854);
nand U7380 (N_7380,N_6439,N_6870);
and U7381 (N_7381,N_6820,N_6393);
xor U7382 (N_7382,N_6721,N_6727);
or U7383 (N_7383,N_6928,N_6981);
xnor U7384 (N_7384,N_6018,N_6478);
xor U7385 (N_7385,N_6331,N_6314);
and U7386 (N_7386,N_6787,N_6251);
and U7387 (N_7387,N_6339,N_6662);
and U7388 (N_7388,N_6644,N_6264);
nand U7389 (N_7389,N_6926,N_6287);
xor U7390 (N_7390,N_6545,N_6871);
nor U7391 (N_7391,N_6153,N_6351);
nor U7392 (N_7392,N_6783,N_6037);
and U7393 (N_7393,N_6194,N_6252);
and U7394 (N_7394,N_6764,N_6054);
nand U7395 (N_7395,N_6017,N_6452);
and U7396 (N_7396,N_6366,N_6963);
xnor U7397 (N_7397,N_6883,N_6007);
nand U7398 (N_7398,N_6079,N_6158);
or U7399 (N_7399,N_6844,N_6853);
nor U7400 (N_7400,N_6332,N_6102);
and U7401 (N_7401,N_6935,N_6429);
and U7402 (N_7402,N_6507,N_6036);
nor U7403 (N_7403,N_6136,N_6465);
xor U7404 (N_7404,N_6070,N_6189);
xnor U7405 (N_7405,N_6989,N_6350);
nor U7406 (N_7406,N_6329,N_6580);
nand U7407 (N_7407,N_6574,N_6612);
nand U7408 (N_7408,N_6444,N_6731);
xnor U7409 (N_7409,N_6709,N_6904);
and U7410 (N_7410,N_6698,N_6253);
nor U7411 (N_7411,N_6209,N_6230);
xnor U7412 (N_7412,N_6831,N_6493);
xor U7413 (N_7413,N_6547,N_6190);
or U7414 (N_7414,N_6133,N_6974);
nor U7415 (N_7415,N_6218,N_6621);
nand U7416 (N_7416,N_6586,N_6529);
nand U7417 (N_7417,N_6934,N_6382);
nor U7418 (N_7418,N_6144,N_6884);
or U7419 (N_7419,N_6421,N_6649);
and U7420 (N_7420,N_6191,N_6533);
nor U7421 (N_7421,N_6093,N_6227);
nor U7422 (N_7422,N_6229,N_6123);
nor U7423 (N_7423,N_6500,N_6954);
nand U7424 (N_7424,N_6082,N_6607);
nand U7425 (N_7425,N_6577,N_6859);
nand U7426 (N_7426,N_6713,N_6367);
xnor U7427 (N_7427,N_6170,N_6335);
xor U7428 (N_7428,N_6943,N_6220);
xnor U7429 (N_7429,N_6010,N_6931);
xor U7430 (N_7430,N_6397,N_6294);
and U7431 (N_7431,N_6001,N_6559);
nand U7432 (N_7432,N_6035,N_6171);
and U7433 (N_7433,N_6295,N_6970);
or U7434 (N_7434,N_6166,N_6046);
nand U7435 (N_7435,N_6555,N_6308);
xor U7436 (N_7436,N_6292,N_6090);
nor U7437 (N_7437,N_6751,N_6231);
or U7438 (N_7438,N_6572,N_6836);
or U7439 (N_7439,N_6741,N_6061);
xnor U7440 (N_7440,N_6592,N_6680);
nand U7441 (N_7441,N_6479,N_6927);
nor U7442 (N_7442,N_6111,N_6811);
xnor U7443 (N_7443,N_6275,N_6462);
nor U7444 (N_7444,N_6004,N_6685);
xnor U7445 (N_7445,N_6945,N_6579);
xnor U7446 (N_7446,N_6827,N_6152);
nand U7447 (N_7447,N_6108,N_6160);
or U7448 (N_7448,N_6441,N_6947);
xor U7449 (N_7449,N_6370,N_6752);
xnor U7450 (N_7450,N_6407,N_6269);
or U7451 (N_7451,N_6538,N_6561);
nor U7452 (N_7452,N_6924,N_6725);
xor U7453 (N_7453,N_6197,N_6065);
or U7454 (N_7454,N_6767,N_6719);
xor U7455 (N_7455,N_6702,N_6710);
and U7456 (N_7456,N_6940,N_6277);
xor U7457 (N_7457,N_6459,N_6878);
nand U7458 (N_7458,N_6381,N_6656);
or U7459 (N_7459,N_6087,N_6674);
and U7460 (N_7460,N_6667,N_6185);
nand U7461 (N_7461,N_6234,N_6149);
or U7462 (N_7462,N_6115,N_6025);
xnor U7463 (N_7463,N_6419,N_6019);
and U7464 (N_7464,N_6453,N_6386);
nor U7465 (N_7465,N_6288,N_6263);
nor U7466 (N_7466,N_6373,N_6860);
nand U7467 (N_7467,N_6615,N_6960);
and U7468 (N_7468,N_6147,N_6641);
and U7469 (N_7469,N_6593,N_6223);
xnor U7470 (N_7470,N_6395,N_6163);
nand U7471 (N_7471,N_6501,N_6530);
or U7472 (N_7472,N_6014,N_6562);
or U7473 (N_7473,N_6486,N_6591);
and U7474 (N_7474,N_6881,N_6296);
and U7475 (N_7475,N_6618,N_6614);
nand U7476 (N_7476,N_6979,N_6525);
nor U7477 (N_7477,N_6608,N_6369);
and U7478 (N_7478,N_6850,N_6206);
xor U7479 (N_7479,N_6812,N_6002);
nand U7480 (N_7480,N_6143,N_6568);
xor U7481 (N_7481,N_6718,N_6704);
xnor U7482 (N_7482,N_6365,N_6283);
or U7483 (N_7483,N_6216,N_6208);
and U7484 (N_7484,N_6423,N_6825);
xnor U7485 (N_7485,N_6551,N_6971);
xor U7486 (N_7486,N_6177,N_6318);
xnor U7487 (N_7487,N_6650,N_6948);
nand U7488 (N_7488,N_6893,N_6750);
nand U7489 (N_7489,N_6792,N_6448);
or U7490 (N_7490,N_6576,N_6784);
or U7491 (N_7491,N_6038,N_6298);
nand U7492 (N_7492,N_6414,N_6129);
xor U7493 (N_7493,N_6804,N_6651);
and U7494 (N_7494,N_6617,N_6075);
nor U7495 (N_7495,N_6846,N_6261);
and U7496 (N_7496,N_6609,N_6431);
xnor U7497 (N_7497,N_6310,N_6184);
or U7498 (N_7498,N_6939,N_6510);
or U7499 (N_7499,N_6055,N_6286);
xnor U7500 (N_7500,N_6160,N_6912);
nand U7501 (N_7501,N_6501,N_6054);
nand U7502 (N_7502,N_6519,N_6612);
and U7503 (N_7503,N_6618,N_6995);
or U7504 (N_7504,N_6563,N_6585);
xnor U7505 (N_7505,N_6933,N_6466);
xnor U7506 (N_7506,N_6355,N_6880);
nor U7507 (N_7507,N_6037,N_6770);
nor U7508 (N_7508,N_6519,N_6940);
and U7509 (N_7509,N_6844,N_6148);
xnor U7510 (N_7510,N_6019,N_6985);
nand U7511 (N_7511,N_6465,N_6346);
xnor U7512 (N_7512,N_6738,N_6989);
or U7513 (N_7513,N_6555,N_6961);
or U7514 (N_7514,N_6658,N_6184);
nor U7515 (N_7515,N_6578,N_6585);
nor U7516 (N_7516,N_6477,N_6384);
or U7517 (N_7517,N_6315,N_6988);
or U7518 (N_7518,N_6439,N_6542);
nand U7519 (N_7519,N_6320,N_6561);
nand U7520 (N_7520,N_6243,N_6951);
nand U7521 (N_7521,N_6459,N_6296);
nor U7522 (N_7522,N_6794,N_6519);
or U7523 (N_7523,N_6941,N_6856);
and U7524 (N_7524,N_6838,N_6153);
and U7525 (N_7525,N_6423,N_6812);
nor U7526 (N_7526,N_6957,N_6552);
and U7527 (N_7527,N_6163,N_6741);
nand U7528 (N_7528,N_6095,N_6078);
nand U7529 (N_7529,N_6177,N_6918);
and U7530 (N_7530,N_6791,N_6430);
xnor U7531 (N_7531,N_6345,N_6945);
nand U7532 (N_7532,N_6436,N_6929);
xor U7533 (N_7533,N_6073,N_6668);
or U7534 (N_7534,N_6237,N_6428);
and U7535 (N_7535,N_6966,N_6773);
nor U7536 (N_7536,N_6069,N_6670);
and U7537 (N_7537,N_6727,N_6912);
nand U7538 (N_7538,N_6428,N_6944);
or U7539 (N_7539,N_6686,N_6513);
xnor U7540 (N_7540,N_6520,N_6349);
nand U7541 (N_7541,N_6298,N_6326);
and U7542 (N_7542,N_6957,N_6788);
nor U7543 (N_7543,N_6416,N_6136);
xor U7544 (N_7544,N_6871,N_6612);
nor U7545 (N_7545,N_6571,N_6262);
nand U7546 (N_7546,N_6785,N_6510);
nand U7547 (N_7547,N_6135,N_6955);
or U7548 (N_7548,N_6431,N_6935);
nand U7549 (N_7549,N_6473,N_6006);
nand U7550 (N_7550,N_6579,N_6138);
or U7551 (N_7551,N_6772,N_6414);
and U7552 (N_7552,N_6773,N_6257);
xor U7553 (N_7553,N_6341,N_6601);
nor U7554 (N_7554,N_6494,N_6967);
nor U7555 (N_7555,N_6630,N_6272);
nor U7556 (N_7556,N_6949,N_6483);
or U7557 (N_7557,N_6866,N_6110);
xor U7558 (N_7558,N_6278,N_6419);
xnor U7559 (N_7559,N_6302,N_6163);
nand U7560 (N_7560,N_6549,N_6565);
nand U7561 (N_7561,N_6037,N_6638);
nand U7562 (N_7562,N_6413,N_6776);
and U7563 (N_7563,N_6327,N_6446);
or U7564 (N_7564,N_6613,N_6542);
xnor U7565 (N_7565,N_6358,N_6125);
and U7566 (N_7566,N_6690,N_6827);
or U7567 (N_7567,N_6912,N_6907);
xnor U7568 (N_7568,N_6674,N_6411);
nand U7569 (N_7569,N_6944,N_6376);
nor U7570 (N_7570,N_6701,N_6705);
nand U7571 (N_7571,N_6890,N_6797);
nand U7572 (N_7572,N_6813,N_6097);
or U7573 (N_7573,N_6089,N_6228);
nor U7574 (N_7574,N_6287,N_6202);
xnor U7575 (N_7575,N_6382,N_6026);
xnor U7576 (N_7576,N_6825,N_6968);
nand U7577 (N_7577,N_6290,N_6882);
and U7578 (N_7578,N_6370,N_6555);
nand U7579 (N_7579,N_6960,N_6029);
nor U7580 (N_7580,N_6558,N_6447);
nand U7581 (N_7581,N_6970,N_6041);
and U7582 (N_7582,N_6495,N_6650);
and U7583 (N_7583,N_6799,N_6859);
nor U7584 (N_7584,N_6154,N_6109);
and U7585 (N_7585,N_6006,N_6632);
nor U7586 (N_7586,N_6776,N_6302);
xnor U7587 (N_7587,N_6318,N_6223);
nor U7588 (N_7588,N_6462,N_6915);
nor U7589 (N_7589,N_6733,N_6243);
nor U7590 (N_7590,N_6618,N_6154);
or U7591 (N_7591,N_6667,N_6499);
xor U7592 (N_7592,N_6485,N_6777);
nand U7593 (N_7593,N_6369,N_6542);
nand U7594 (N_7594,N_6636,N_6873);
nand U7595 (N_7595,N_6490,N_6378);
nor U7596 (N_7596,N_6024,N_6285);
nor U7597 (N_7597,N_6444,N_6235);
xor U7598 (N_7598,N_6051,N_6175);
and U7599 (N_7599,N_6172,N_6784);
or U7600 (N_7600,N_6700,N_6148);
nand U7601 (N_7601,N_6489,N_6961);
or U7602 (N_7602,N_6018,N_6258);
xnor U7603 (N_7603,N_6755,N_6524);
or U7604 (N_7604,N_6383,N_6263);
nor U7605 (N_7605,N_6955,N_6642);
nand U7606 (N_7606,N_6071,N_6419);
nor U7607 (N_7607,N_6429,N_6395);
or U7608 (N_7608,N_6411,N_6244);
and U7609 (N_7609,N_6188,N_6601);
nor U7610 (N_7610,N_6949,N_6027);
or U7611 (N_7611,N_6386,N_6373);
nor U7612 (N_7612,N_6982,N_6578);
nand U7613 (N_7613,N_6983,N_6376);
xor U7614 (N_7614,N_6588,N_6879);
nor U7615 (N_7615,N_6496,N_6331);
xor U7616 (N_7616,N_6485,N_6407);
xnor U7617 (N_7617,N_6357,N_6413);
nand U7618 (N_7618,N_6089,N_6352);
nand U7619 (N_7619,N_6682,N_6985);
xor U7620 (N_7620,N_6453,N_6162);
nand U7621 (N_7621,N_6861,N_6739);
xor U7622 (N_7622,N_6244,N_6746);
or U7623 (N_7623,N_6825,N_6767);
or U7624 (N_7624,N_6460,N_6393);
and U7625 (N_7625,N_6175,N_6285);
nand U7626 (N_7626,N_6721,N_6679);
xnor U7627 (N_7627,N_6330,N_6948);
xnor U7628 (N_7628,N_6149,N_6959);
and U7629 (N_7629,N_6818,N_6064);
or U7630 (N_7630,N_6205,N_6212);
or U7631 (N_7631,N_6710,N_6557);
nor U7632 (N_7632,N_6117,N_6459);
xor U7633 (N_7633,N_6853,N_6004);
xnor U7634 (N_7634,N_6195,N_6619);
xor U7635 (N_7635,N_6203,N_6021);
or U7636 (N_7636,N_6601,N_6312);
or U7637 (N_7637,N_6877,N_6842);
or U7638 (N_7638,N_6031,N_6316);
nor U7639 (N_7639,N_6222,N_6691);
and U7640 (N_7640,N_6181,N_6314);
xnor U7641 (N_7641,N_6905,N_6480);
or U7642 (N_7642,N_6930,N_6345);
nor U7643 (N_7643,N_6335,N_6512);
xor U7644 (N_7644,N_6444,N_6322);
or U7645 (N_7645,N_6450,N_6007);
nor U7646 (N_7646,N_6765,N_6634);
nand U7647 (N_7647,N_6029,N_6512);
or U7648 (N_7648,N_6741,N_6416);
xor U7649 (N_7649,N_6408,N_6305);
nor U7650 (N_7650,N_6976,N_6799);
nor U7651 (N_7651,N_6689,N_6378);
and U7652 (N_7652,N_6016,N_6542);
nand U7653 (N_7653,N_6798,N_6975);
xnor U7654 (N_7654,N_6717,N_6675);
xnor U7655 (N_7655,N_6419,N_6907);
or U7656 (N_7656,N_6551,N_6095);
nand U7657 (N_7657,N_6547,N_6178);
nor U7658 (N_7658,N_6713,N_6120);
nor U7659 (N_7659,N_6194,N_6213);
and U7660 (N_7660,N_6805,N_6007);
or U7661 (N_7661,N_6370,N_6649);
xor U7662 (N_7662,N_6292,N_6227);
and U7663 (N_7663,N_6403,N_6372);
and U7664 (N_7664,N_6019,N_6362);
nor U7665 (N_7665,N_6462,N_6027);
and U7666 (N_7666,N_6730,N_6891);
nand U7667 (N_7667,N_6438,N_6489);
nand U7668 (N_7668,N_6411,N_6217);
nor U7669 (N_7669,N_6699,N_6161);
or U7670 (N_7670,N_6107,N_6466);
nand U7671 (N_7671,N_6534,N_6494);
nor U7672 (N_7672,N_6860,N_6063);
and U7673 (N_7673,N_6931,N_6105);
xor U7674 (N_7674,N_6344,N_6868);
nand U7675 (N_7675,N_6318,N_6033);
xor U7676 (N_7676,N_6792,N_6765);
xor U7677 (N_7677,N_6325,N_6903);
xnor U7678 (N_7678,N_6970,N_6280);
nand U7679 (N_7679,N_6582,N_6949);
or U7680 (N_7680,N_6297,N_6975);
nor U7681 (N_7681,N_6528,N_6422);
nand U7682 (N_7682,N_6838,N_6077);
xnor U7683 (N_7683,N_6500,N_6270);
or U7684 (N_7684,N_6825,N_6820);
and U7685 (N_7685,N_6906,N_6450);
xnor U7686 (N_7686,N_6603,N_6995);
and U7687 (N_7687,N_6747,N_6640);
and U7688 (N_7688,N_6190,N_6766);
and U7689 (N_7689,N_6802,N_6961);
nor U7690 (N_7690,N_6105,N_6711);
and U7691 (N_7691,N_6613,N_6559);
and U7692 (N_7692,N_6715,N_6649);
and U7693 (N_7693,N_6647,N_6862);
or U7694 (N_7694,N_6719,N_6062);
nor U7695 (N_7695,N_6811,N_6405);
nor U7696 (N_7696,N_6654,N_6463);
xnor U7697 (N_7697,N_6527,N_6118);
xor U7698 (N_7698,N_6846,N_6926);
nor U7699 (N_7699,N_6600,N_6760);
nand U7700 (N_7700,N_6260,N_6293);
or U7701 (N_7701,N_6432,N_6727);
nor U7702 (N_7702,N_6065,N_6925);
and U7703 (N_7703,N_6846,N_6012);
nand U7704 (N_7704,N_6127,N_6184);
or U7705 (N_7705,N_6463,N_6369);
or U7706 (N_7706,N_6503,N_6384);
nand U7707 (N_7707,N_6935,N_6287);
or U7708 (N_7708,N_6500,N_6058);
nor U7709 (N_7709,N_6607,N_6070);
nor U7710 (N_7710,N_6591,N_6069);
or U7711 (N_7711,N_6873,N_6218);
nor U7712 (N_7712,N_6337,N_6064);
nand U7713 (N_7713,N_6798,N_6339);
nor U7714 (N_7714,N_6018,N_6255);
xor U7715 (N_7715,N_6539,N_6210);
nor U7716 (N_7716,N_6975,N_6075);
nor U7717 (N_7717,N_6001,N_6020);
nor U7718 (N_7718,N_6028,N_6308);
xor U7719 (N_7719,N_6517,N_6113);
and U7720 (N_7720,N_6774,N_6031);
nand U7721 (N_7721,N_6481,N_6629);
xnor U7722 (N_7722,N_6133,N_6584);
nor U7723 (N_7723,N_6735,N_6553);
nor U7724 (N_7724,N_6801,N_6706);
xor U7725 (N_7725,N_6482,N_6462);
and U7726 (N_7726,N_6217,N_6295);
and U7727 (N_7727,N_6560,N_6538);
and U7728 (N_7728,N_6319,N_6316);
or U7729 (N_7729,N_6946,N_6013);
xor U7730 (N_7730,N_6184,N_6837);
and U7731 (N_7731,N_6374,N_6158);
and U7732 (N_7732,N_6972,N_6583);
or U7733 (N_7733,N_6038,N_6879);
and U7734 (N_7734,N_6349,N_6370);
nor U7735 (N_7735,N_6272,N_6406);
or U7736 (N_7736,N_6250,N_6776);
nand U7737 (N_7737,N_6059,N_6136);
nand U7738 (N_7738,N_6329,N_6096);
or U7739 (N_7739,N_6060,N_6516);
nor U7740 (N_7740,N_6680,N_6270);
xnor U7741 (N_7741,N_6082,N_6887);
and U7742 (N_7742,N_6986,N_6680);
xor U7743 (N_7743,N_6735,N_6613);
and U7744 (N_7744,N_6055,N_6971);
and U7745 (N_7745,N_6357,N_6625);
and U7746 (N_7746,N_6937,N_6373);
nor U7747 (N_7747,N_6127,N_6340);
nor U7748 (N_7748,N_6244,N_6154);
or U7749 (N_7749,N_6672,N_6376);
nor U7750 (N_7750,N_6747,N_6589);
or U7751 (N_7751,N_6133,N_6490);
or U7752 (N_7752,N_6660,N_6891);
xor U7753 (N_7753,N_6511,N_6867);
nand U7754 (N_7754,N_6954,N_6415);
and U7755 (N_7755,N_6599,N_6852);
nand U7756 (N_7756,N_6856,N_6547);
xnor U7757 (N_7757,N_6141,N_6739);
nor U7758 (N_7758,N_6152,N_6072);
xor U7759 (N_7759,N_6565,N_6641);
and U7760 (N_7760,N_6231,N_6926);
nor U7761 (N_7761,N_6895,N_6291);
nand U7762 (N_7762,N_6604,N_6833);
or U7763 (N_7763,N_6304,N_6163);
nor U7764 (N_7764,N_6157,N_6430);
xnor U7765 (N_7765,N_6798,N_6309);
or U7766 (N_7766,N_6869,N_6399);
xor U7767 (N_7767,N_6681,N_6002);
nor U7768 (N_7768,N_6683,N_6452);
xor U7769 (N_7769,N_6306,N_6038);
xnor U7770 (N_7770,N_6554,N_6317);
or U7771 (N_7771,N_6858,N_6339);
nor U7772 (N_7772,N_6274,N_6524);
nor U7773 (N_7773,N_6897,N_6162);
nand U7774 (N_7774,N_6918,N_6764);
nor U7775 (N_7775,N_6917,N_6470);
nand U7776 (N_7776,N_6588,N_6781);
or U7777 (N_7777,N_6570,N_6254);
xor U7778 (N_7778,N_6232,N_6108);
or U7779 (N_7779,N_6353,N_6789);
nand U7780 (N_7780,N_6791,N_6375);
xnor U7781 (N_7781,N_6827,N_6771);
nand U7782 (N_7782,N_6898,N_6926);
xor U7783 (N_7783,N_6185,N_6482);
and U7784 (N_7784,N_6219,N_6881);
or U7785 (N_7785,N_6447,N_6336);
nor U7786 (N_7786,N_6922,N_6607);
nor U7787 (N_7787,N_6150,N_6320);
nor U7788 (N_7788,N_6676,N_6105);
and U7789 (N_7789,N_6649,N_6546);
or U7790 (N_7790,N_6132,N_6087);
xnor U7791 (N_7791,N_6943,N_6672);
and U7792 (N_7792,N_6818,N_6259);
and U7793 (N_7793,N_6518,N_6067);
nor U7794 (N_7794,N_6772,N_6331);
xor U7795 (N_7795,N_6829,N_6436);
nand U7796 (N_7796,N_6415,N_6983);
nor U7797 (N_7797,N_6094,N_6847);
and U7798 (N_7798,N_6718,N_6973);
and U7799 (N_7799,N_6636,N_6966);
or U7800 (N_7800,N_6386,N_6116);
nand U7801 (N_7801,N_6717,N_6193);
or U7802 (N_7802,N_6712,N_6715);
and U7803 (N_7803,N_6833,N_6664);
nor U7804 (N_7804,N_6373,N_6458);
nor U7805 (N_7805,N_6511,N_6231);
nor U7806 (N_7806,N_6289,N_6427);
and U7807 (N_7807,N_6827,N_6658);
and U7808 (N_7808,N_6006,N_6551);
nand U7809 (N_7809,N_6733,N_6669);
and U7810 (N_7810,N_6479,N_6149);
xor U7811 (N_7811,N_6623,N_6509);
or U7812 (N_7812,N_6661,N_6148);
xnor U7813 (N_7813,N_6890,N_6127);
xor U7814 (N_7814,N_6201,N_6385);
or U7815 (N_7815,N_6099,N_6918);
nand U7816 (N_7816,N_6008,N_6963);
and U7817 (N_7817,N_6920,N_6170);
xnor U7818 (N_7818,N_6670,N_6296);
nand U7819 (N_7819,N_6714,N_6997);
nor U7820 (N_7820,N_6277,N_6863);
nand U7821 (N_7821,N_6544,N_6421);
nor U7822 (N_7822,N_6433,N_6082);
xor U7823 (N_7823,N_6720,N_6763);
or U7824 (N_7824,N_6103,N_6859);
xnor U7825 (N_7825,N_6391,N_6284);
nand U7826 (N_7826,N_6139,N_6179);
or U7827 (N_7827,N_6858,N_6177);
nand U7828 (N_7828,N_6853,N_6669);
nand U7829 (N_7829,N_6837,N_6323);
xnor U7830 (N_7830,N_6148,N_6598);
nand U7831 (N_7831,N_6419,N_6477);
nor U7832 (N_7832,N_6041,N_6134);
xnor U7833 (N_7833,N_6628,N_6012);
nor U7834 (N_7834,N_6332,N_6505);
xnor U7835 (N_7835,N_6819,N_6185);
or U7836 (N_7836,N_6925,N_6497);
or U7837 (N_7837,N_6780,N_6523);
nand U7838 (N_7838,N_6865,N_6528);
and U7839 (N_7839,N_6871,N_6784);
nand U7840 (N_7840,N_6657,N_6760);
and U7841 (N_7841,N_6171,N_6239);
nand U7842 (N_7842,N_6826,N_6968);
xnor U7843 (N_7843,N_6009,N_6858);
nor U7844 (N_7844,N_6063,N_6199);
nand U7845 (N_7845,N_6804,N_6904);
xor U7846 (N_7846,N_6656,N_6340);
or U7847 (N_7847,N_6184,N_6569);
or U7848 (N_7848,N_6249,N_6179);
nand U7849 (N_7849,N_6833,N_6687);
xnor U7850 (N_7850,N_6263,N_6243);
or U7851 (N_7851,N_6812,N_6059);
nor U7852 (N_7852,N_6972,N_6238);
xnor U7853 (N_7853,N_6146,N_6665);
nand U7854 (N_7854,N_6214,N_6853);
or U7855 (N_7855,N_6939,N_6802);
and U7856 (N_7856,N_6921,N_6502);
nand U7857 (N_7857,N_6531,N_6201);
xnor U7858 (N_7858,N_6830,N_6653);
nand U7859 (N_7859,N_6036,N_6220);
nand U7860 (N_7860,N_6348,N_6479);
or U7861 (N_7861,N_6537,N_6934);
nor U7862 (N_7862,N_6629,N_6746);
and U7863 (N_7863,N_6925,N_6835);
and U7864 (N_7864,N_6205,N_6525);
and U7865 (N_7865,N_6442,N_6445);
xor U7866 (N_7866,N_6409,N_6922);
nand U7867 (N_7867,N_6478,N_6720);
nor U7868 (N_7868,N_6492,N_6665);
nand U7869 (N_7869,N_6234,N_6702);
nor U7870 (N_7870,N_6954,N_6115);
xor U7871 (N_7871,N_6450,N_6683);
xnor U7872 (N_7872,N_6517,N_6038);
nand U7873 (N_7873,N_6667,N_6267);
nor U7874 (N_7874,N_6420,N_6289);
nand U7875 (N_7875,N_6274,N_6005);
xor U7876 (N_7876,N_6074,N_6875);
nand U7877 (N_7877,N_6855,N_6630);
nand U7878 (N_7878,N_6974,N_6863);
or U7879 (N_7879,N_6824,N_6409);
xor U7880 (N_7880,N_6719,N_6979);
and U7881 (N_7881,N_6357,N_6572);
and U7882 (N_7882,N_6559,N_6072);
nor U7883 (N_7883,N_6479,N_6712);
xnor U7884 (N_7884,N_6254,N_6763);
or U7885 (N_7885,N_6325,N_6895);
xnor U7886 (N_7886,N_6923,N_6562);
nand U7887 (N_7887,N_6618,N_6344);
and U7888 (N_7888,N_6050,N_6537);
nand U7889 (N_7889,N_6788,N_6022);
nor U7890 (N_7890,N_6915,N_6222);
xor U7891 (N_7891,N_6232,N_6754);
xor U7892 (N_7892,N_6294,N_6576);
nor U7893 (N_7893,N_6464,N_6171);
or U7894 (N_7894,N_6542,N_6193);
xnor U7895 (N_7895,N_6869,N_6521);
or U7896 (N_7896,N_6433,N_6834);
nor U7897 (N_7897,N_6708,N_6142);
xor U7898 (N_7898,N_6569,N_6204);
nand U7899 (N_7899,N_6800,N_6549);
or U7900 (N_7900,N_6114,N_6517);
nor U7901 (N_7901,N_6739,N_6695);
nor U7902 (N_7902,N_6353,N_6149);
nor U7903 (N_7903,N_6206,N_6113);
and U7904 (N_7904,N_6774,N_6009);
and U7905 (N_7905,N_6113,N_6501);
nor U7906 (N_7906,N_6777,N_6043);
nor U7907 (N_7907,N_6636,N_6408);
nand U7908 (N_7908,N_6659,N_6854);
nand U7909 (N_7909,N_6660,N_6453);
and U7910 (N_7910,N_6247,N_6023);
xnor U7911 (N_7911,N_6577,N_6436);
or U7912 (N_7912,N_6209,N_6468);
nor U7913 (N_7913,N_6988,N_6515);
and U7914 (N_7914,N_6980,N_6609);
xnor U7915 (N_7915,N_6949,N_6630);
xor U7916 (N_7916,N_6740,N_6484);
nor U7917 (N_7917,N_6807,N_6961);
xnor U7918 (N_7918,N_6052,N_6169);
or U7919 (N_7919,N_6040,N_6079);
and U7920 (N_7920,N_6589,N_6247);
or U7921 (N_7921,N_6987,N_6189);
and U7922 (N_7922,N_6051,N_6329);
nor U7923 (N_7923,N_6877,N_6561);
and U7924 (N_7924,N_6951,N_6210);
nor U7925 (N_7925,N_6117,N_6166);
xnor U7926 (N_7926,N_6988,N_6662);
xnor U7927 (N_7927,N_6811,N_6687);
and U7928 (N_7928,N_6680,N_6107);
or U7929 (N_7929,N_6082,N_6027);
xor U7930 (N_7930,N_6765,N_6313);
nand U7931 (N_7931,N_6684,N_6299);
xor U7932 (N_7932,N_6599,N_6813);
or U7933 (N_7933,N_6158,N_6062);
and U7934 (N_7934,N_6298,N_6523);
xor U7935 (N_7935,N_6315,N_6461);
nor U7936 (N_7936,N_6938,N_6376);
nor U7937 (N_7937,N_6980,N_6492);
xor U7938 (N_7938,N_6495,N_6215);
and U7939 (N_7939,N_6208,N_6167);
xnor U7940 (N_7940,N_6762,N_6781);
nand U7941 (N_7941,N_6934,N_6170);
nor U7942 (N_7942,N_6213,N_6452);
nor U7943 (N_7943,N_6905,N_6797);
nand U7944 (N_7944,N_6370,N_6482);
xor U7945 (N_7945,N_6017,N_6662);
and U7946 (N_7946,N_6219,N_6463);
nand U7947 (N_7947,N_6774,N_6763);
or U7948 (N_7948,N_6279,N_6895);
xor U7949 (N_7949,N_6562,N_6698);
nor U7950 (N_7950,N_6017,N_6390);
xor U7951 (N_7951,N_6151,N_6996);
nor U7952 (N_7952,N_6012,N_6094);
nor U7953 (N_7953,N_6947,N_6922);
nor U7954 (N_7954,N_6997,N_6933);
or U7955 (N_7955,N_6238,N_6420);
or U7956 (N_7956,N_6380,N_6822);
or U7957 (N_7957,N_6910,N_6756);
or U7958 (N_7958,N_6580,N_6408);
xnor U7959 (N_7959,N_6723,N_6690);
or U7960 (N_7960,N_6593,N_6897);
xnor U7961 (N_7961,N_6779,N_6108);
nand U7962 (N_7962,N_6789,N_6942);
nand U7963 (N_7963,N_6055,N_6169);
nor U7964 (N_7964,N_6255,N_6823);
nand U7965 (N_7965,N_6961,N_6213);
and U7966 (N_7966,N_6916,N_6874);
and U7967 (N_7967,N_6665,N_6334);
xor U7968 (N_7968,N_6664,N_6506);
or U7969 (N_7969,N_6071,N_6561);
nand U7970 (N_7970,N_6560,N_6524);
and U7971 (N_7971,N_6179,N_6338);
and U7972 (N_7972,N_6518,N_6879);
nand U7973 (N_7973,N_6899,N_6354);
nand U7974 (N_7974,N_6204,N_6149);
or U7975 (N_7975,N_6880,N_6520);
nand U7976 (N_7976,N_6445,N_6433);
nand U7977 (N_7977,N_6896,N_6455);
or U7978 (N_7978,N_6043,N_6899);
or U7979 (N_7979,N_6058,N_6847);
or U7980 (N_7980,N_6138,N_6673);
nor U7981 (N_7981,N_6845,N_6529);
or U7982 (N_7982,N_6536,N_6197);
and U7983 (N_7983,N_6639,N_6752);
nor U7984 (N_7984,N_6654,N_6424);
xnor U7985 (N_7985,N_6060,N_6589);
nand U7986 (N_7986,N_6613,N_6885);
nand U7987 (N_7987,N_6734,N_6108);
or U7988 (N_7988,N_6315,N_6459);
nor U7989 (N_7989,N_6533,N_6970);
xnor U7990 (N_7990,N_6055,N_6440);
and U7991 (N_7991,N_6085,N_6799);
nand U7992 (N_7992,N_6374,N_6798);
and U7993 (N_7993,N_6042,N_6238);
and U7994 (N_7994,N_6711,N_6987);
nand U7995 (N_7995,N_6373,N_6415);
xor U7996 (N_7996,N_6075,N_6679);
nand U7997 (N_7997,N_6610,N_6285);
xnor U7998 (N_7998,N_6322,N_6094);
nand U7999 (N_7999,N_6498,N_6929);
and U8000 (N_8000,N_7639,N_7445);
xor U8001 (N_8001,N_7843,N_7151);
xor U8002 (N_8002,N_7520,N_7970);
nor U8003 (N_8003,N_7072,N_7273);
and U8004 (N_8004,N_7663,N_7534);
nor U8005 (N_8005,N_7932,N_7923);
or U8006 (N_8006,N_7166,N_7360);
nor U8007 (N_8007,N_7288,N_7752);
and U8008 (N_8008,N_7801,N_7355);
xor U8009 (N_8009,N_7007,N_7759);
nor U8010 (N_8010,N_7548,N_7928);
or U8011 (N_8011,N_7834,N_7430);
xnor U8012 (N_8012,N_7758,N_7167);
nand U8013 (N_8013,N_7260,N_7099);
nor U8014 (N_8014,N_7746,N_7233);
xnor U8015 (N_8015,N_7016,N_7366);
nand U8016 (N_8016,N_7154,N_7836);
or U8017 (N_8017,N_7473,N_7209);
xnor U8018 (N_8018,N_7344,N_7175);
xnor U8019 (N_8019,N_7791,N_7503);
nor U8020 (N_8020,N_7434,N_7457);
or U8021 (N_8021,N_7677,N_7950);
nand U8022 (N_8022,N_7346,N_7227);
nand U8023 (N_8023,N_7308,N_7540);
or U8024 (N_8024,N_7743,N_7010);
or U8025 (N_8025,N_7555,N_7044);
xnor U8026 (N_8026,N_7341,N_7157);
or U8027 (N_8027,N_7423,N_7414);
nor U8028 (N_8028,N_7169,N_7625);
and U8029 (N_8029,N_7137,N_7692);
nor U8030 (N_8030,N_7714,N_7249);
and U8031 (N_8031,N_7148,N_7394);
or U8032 (N_8032,N_7664,N_7674);
or U8033 (N_8033,N_7488,N_7860);
xnor U8034 (N_8034,N_7586,N_7588);
and U8035 (N_8035,N_7571,N_7969);
xnor U8036 (N_8036,N_7324,N_7163);
nand U8037 (N_8037,N_7785,N_7908);
and U8038 (N_8038,N_7081,N_7601);
xor U8039 (N_8039,N_7297,N_7237);
and U8040 (N_8040,N_7626,N_7257);
or U8041 (N_8041,N_7740,N_7840);
xor U8042 (N_8042,N_7939,N_7609);
or U8043 (N_8043,N_7802,N_7196);
nor U8044 (N_8044,N_7915,N_7943);
nand U8045 (N_8045,N_7831,N_7634);
nand U8046 (N_8046,N_7242,N_7245);
nor U8047 (N_8047,N_7486,N_7980);
or U8048 (N_8048,N_7188,N_7968);
nor U8049 (N_8049,N_7522,N_7628);
nor U8050 (N_8050,N_7333,N_7780);
and U8051 (N_8051,N_7418,N_7938);
xor U8052 (N_8052,N_7795,N_7222);
xnor U8053 (N_8053,N_7413,N_7589);
xnor U8054 (N_8054,N_7976,N_7567);
and U8055 (N_8055,N_7104,N_7255);
nand U8056 (N_8056,N_7431,N_7761);
and U8057 (N_8057,N_7496,N_7158);
nor U8058 (N_8058,N_7213,N_7367);
or U8059 (N_8059,N_7595,N_7047);
or U8060 (N_8060,N_7129,N_7974);
and U8061 (N_8061,N_7028,N_7807);
or U8062 (N_8062,N_7830,N_7820);
nand U8063 (N_8063,N_7614,N_7141);
nor U8064 (N_8064,N_7187,N_7191);
xor U8065 (N_8065,N_7093,N_7608);
nand U8066 (N_8066,N_7882,N_7310);
and U8067 (N_8067,N_7847,N_7858);
nand U8068 (N_8068,N_7754,N_7916);
and U8069 (N_8069,N_7929,N_7417);
xnor U8070 (N_8070,N_7981,N_7318);
and U8071 (N_8071,N_7100,N_7616);
nor U8072 (N_8072,N_7685,N_7914);
nor U8073 (N_8073,N_7862,N_7621);
nor U8074 (N_8074,N_7507,N_7777);
and U8075 (N_8075,N_7591,N_7700);
or U8076 (N_8076,N_7605,N_7892);
and U8077 (N_8077,N_7117,N_7263);
nor U8078 (N_8078,N_7879,N_7361);
or U8079 (N_8079,N_7181,N_7881);
nand U8080 (N_8080,N_7236,N_7271);
xnor U8081 (N_8081,N_7744,N_7107);
nor U8082 (N_8082,N_7941,N_7889);
nand U8083 (N_8083,N_7088,N_7230);
xor U8084 (N_8084,N_7190,N_7715);
or U8085 (N_8085,N_7265,N_7364);
nor U8086 (N_8086,N_7436,N_7351);
or U8087 (N_8087,N_7471,N_7839);
or U8088 (N_8088,N_7809,N_7682);
nor U8089 (N_8089,N_7327,N_7816);
and U8090 (N_8090,N_7304,N_7590);
xnor U8091 (N_8091,N_7670,N_7138);
or U8092 (N_8092,N_7145,N_7221);
and U8093 (N_8093,N_7096,N_7641);
nor U8094 (N_8094,N_7109,N_7579);
and U8095 (N_8095,N_7289,N_7199);
nand U8096 (N_8096,N_7875,N_7426);
xnor U8097 (N_8097,N_7212,N_7671);
nor U8098 (N_8098,N_7721,N_7565);
nand U8099 (N_8099,N_7983,N_7440);
nor U8100 (N_8100,N_7246,N_7127);
xnor U8101 (N_8101,N_7935,N_7610);
or U8102 (N_8102,N_7143,N_7400);
nand U8103 (N_8103,N_7893,N_7907);
nand U8104 (N_8104,N_7696,N_7959);
or U8105 (N_8105,N_7624,N_7676);
nor U8106 (N_8106,N_7003,N_7660);
nor U8107 (N_8107,N_7703,N_7032);
nor U8108 (N_8108,N_7656,N_7755);
nand U8109 (N_8109,N_7511,N_7593);
nor U8110 (N_8110,N_7992,N_7038);
or U8111 (N_8111,N_7015,N_7200);
or U8112 (N_8112,N_7712,N_7899);
nor U8113 (N_8113,N_7517,N_7902);
or U8114 (N_8114,N_7215,N_7037);
and U8115 (N_8115,N_7244,N_7460);
or U8116 (N_8116,N_7543,N_7863);
nor U8117 (N_8117,N_7528,N_7080);
and U8118 (N_8118,N_7856,N_7410);
or U8119 (N_8119,N_7266,N_7612);
or U8120 (N_8120,N_7203,N_7006);
nor U8121 (N_8121,N_7570,N_7115);
and U8122 (N_8122,N_7510,N_7325);
nor U8123 (N_8123,N_7458,N_7197);
and U8124 (N_8124,N_7066,N_7312);
or U8125 (N_8125,N_7952,N_7264);
xnor U8126 (N_8126,N_7763,N_7002);
xnor U8127 (N_8127,N_7438,N_7290);
xor U8128 (N_8128,N_7786,N_7388);
and U8129 (N_8129,N_7111,N_7599);
nand U8130 (N_8130,N_7352,N_7741);
nand U8131 (N_8131,N_7173,N_7894);
or U8132 (N_8132,N_7492,N_7408);
nand U8133 (N_8133,N_7320,N_7615);
xor U8134 (N_8134,N_7424,N_7076);
and U8135 (N_8135,N_7461,N_7018);
nand U8136 (N_8136,N_7219,N_7800);
nand U8137 (N_8137,N_7949,N_7027);
and U8138 (N_8138,N_7268,N_7794);
xor U8139 (N_8139,N_7594,N_7049);
xor U8140 (N_8140,N_7961,N_7299);
xnor U8141 (N_8141,N_7709,N_7449);
nand U8142 (N_8142,N_7720,N_7295);
xnor U8143 (N_8143,N_7033,N_7105);
xnor U8144 (N_8144,N_7012,N_7229);
xor U8145 (N_8145,N_7724,N_7201);
nor U8146 (N_8146,N_7654,N_7505);
xor U8147 (N_8147,N_7706,N_7334);
and U8148 (N_8148,N_7155,N_7963);
nor U8149 (N_8149,N_7697,N_7409);
and U8150 (N_8150,N_7905,N_7693);
xnor U8151 (N_8151,N_7011,N_7087);
xnor U8152 (N_8152,N_7067,N_7330);
xor U8153 (N_8153,N_7705,N_7848);
nand U8154 (N_8154,N_7845,N_7885);
xor U8155 (N_8155,N_7910,N_7248);
xor U8156 (N_8156,N_7851,N_7871);
nor U8157 (N_8157,N_7735,N_7887);
nor U8158 (N_8158,N_7835,N_7787);
nand U8159 (N_8159,N_7844,N_7582);
xor U8160 (N_8160,N_7165,N_7643);
nor U8161 (N_8161,N_7162,N_7640);
or U8162 (N_8162,N_7874,N_7554);
and U8163 (N_8163,N_7279,N_7782);
or U8164 (N_8164,N_7546,N_7526);
nand U8165 (N_8165,N_7684,N_7549);
and U8166 (N_8166,N_7827,N_7149);
nand U8167 (N_8167,N_7506,N_7210);
or U8168 (N_8168,N_7922,N_7962);
xnor U8169 (N_8169,N_7252,N_7756);
nor U8170 (N_8170,N_7134,N_7369);
or U8171 (N_8171,N_7285,N_7850);
and U8172 (N_8172,N_7281,N_7926);
nand U8173 (N_8173,N_7828,N_7483);
nand U8174 (N_8174,N_7957,N_7411);
or U8175 (N_8175,N_7432,N_7017);
or U8176 (N_8176,N_7421,N_7023);
nand U8177 (N_8177,N_7493,N_7365);
nand U8178 (N_8178,N_7177,N_7945);
and U8179 (N_8179,N_7372,N_7514);
or U8180 (N_8180,N_7467,N_7931);
and U8181 (N_8181,N_7453,N_7204);
nor U8182 (N_8182,N_7533,N_7869);
nor U8183 (N_8183,N_7123,N_7283);
or U8184 (N_8184,N_7420,N_7909);
xor U8185 (N_8185,N_7995,N_7933);
xnor U8186 (N_8186,N_7478,N_7098);
and U8187 (N_8187,N_7393,N_7357);
and U8188 (N_8188,N_7536,N_7342);
nand U8189 (N_8189,N_7597,N_7370);
xnor U8190 (N_8190,N_7443,N_7852);
or U8191 (N_8191,N_7773,N_7658);
and U8192 (N_8192,N_7532,N_7259);
and U8193 (N_8193,N_7707,N_7620);
nand U8194 (N_8194,N_7223,N_7888);
nor U8195 (N_8195,N_7508,N_7525);
and U8196 (N_8196,N_7619,N_7766);
xor U8197 (N_8197,N_7822,N_7803);
xnor U8198 (N_8198,N_7328,N_7025);
and U8199 (N_8199,N_7194,N_7000);
nand U8200 (N_8200,N_7812,N_7530);
and U8201 (N_8201,N_7632,N_7054);
and U8202 (N_8202,N_7673,N_7477);
nor U8203 (N_8203,N_7435,N_7195);
or U8204 (N_8204,N_7119,N_7031);
and U8205 (N_8205,N_7009,N_7069);
nand U8206 (N_8206,N_7234,N_7253);
or U8207 (N_8207,N_7552,N_7384);
xor U8208 (N_8208,N_7723,N_7153);
xnor U8209 (N_8209,N_7985,N_7518);
or U8210 (N_8210,N_7247,N_7326);
nor U8211 (N_8211,N_7060,N_7651);
and U8212 (N_8212,N_7359,N_7183);
nand U8213 (N_8213,N_7866,N_7984);
nand U8214 (N_8214,N_7070,N_7005);
nor U8215 (N_8215,N_7332,N_7250);
or U8216 (N_8216,N_7897,N_7272);
nor U8217 (N_8217,N_7085,N_7704);
nand U8218 (N_8218,N_7077,N_7428);
and U8219 (N_8219,N_7282,N_7427);
xor U8220 (N_8220,N_7655,N_7258);
nand U8221 (N_8221,N_7316,N_7113);
xor U8222 (N_8222,N_7627,N_7065);
nor U8223 (N_8223,N_7808,N_7490);
or U8224 (N_8224,N_7819,N_7485);
xor U8225 (N_8225,N_7404,N_7292);
or U8226 (N_8226,N_7736,N_7924);
nand U8227 (N_8227,N_7321,N_7966);
xnor U8228 (N_8228,N_7128,N_7030);
nand U8229 (N_8229,N_7561,N_7405);
xor U8230 (N_8230,N_7563,N_7806);
nand U8231 (N_8231,N_7967,N_7675);
nand U8232 (N_8232,N_7479,N_7583);
nand U8233 (N_8233,N_7878,N_7515);
xnor U8234 (N_8234,N_7101,N_7097);
or U8235 (N_8235,N_7934,N_7550);
and U8236 (N_8236,N_7979,N_7661);
or U8237 (N_8237,N_7564,N_7544);
and U8238 (N_8238,N_7121,N_7398);
and U8239 (N_8239,N_7379,N_7455);
or U8240 (N_8240,N_7577,N_7513);
and U8241 (N_8241,N_7810,N_7349);
xor U8242 (N_8242,N_7650,N_7855);
nor U8243 (N_8243,N_7013,N_7781);
xor U8244 (N_8244,N_7132,N_7681);
nand U8245 (N_8245,N_7226,N_7337);
nand U8246 (N_8246,N_7462,N_7406);
or U8247 (N_8247,N_7059,N_7116);
nor U8248 (N_8248,N_7319,N_7068);
or U8249 (N_8249,N_7383,N_7896);
xor U8250 (N_8250,N_7192,N_7558);
nor U8251 (N_8251,N_7906,N_7779);
xor U8252 (N_8252,N_7161,N_7433);
or U8253 (N_8253,N_7464,N_7380);
or U8254 (N_8254,N_7039,N_7989);
or U8255 (N_8255,N_7416,N_7662);
nor U8256 (N_8256,N_7886,N_7238);
nor U8257 (N_8257,N_7498,N_7322);
nand U8258 (N_8258,N_7374,N_7870);
and U8259 (N_8259,N_7336,N_7140);
xor U8260 (N_8260,N_7106,N_7760);
nand U8261 (N_8261,N_7277,N_7725);
xnor U8262 (N_8262,N_7542,N_7557);
nand U8263 (N_8263,N_7126,N_7958);
and U8264 (N_8264,N_7206,N_7824);
nand U8265 (N_8265,N_7680,N_7559);
or U8266 (N_8266,N_7647,N_7178);
xnor U8267 (N_8267,N_7446,N_7999);
nor U8268 (N_8268,N_7082,N_7971);
nand U8269 (N_8269,N_7224,N_7450);
nor U8270 (N_8270,N_7672,N_7991);
or U8271 (N_8271,N_7338,N_7056);
nor U8272 (N_8272,N_7090,N_7275);
or U8273 (N_8273,N_7302,N_7857);
nand U8274 (N_8274,N_7306,N_7474);
nor U8275 (N_8275,N_7553,N_7377);
xor U8276 (N_8276,N_7294,N_7644);
nand U8277 (N_8277,N_7683,N_7489);
nor U8278 (N_8278,N_7103,N_7347);
xor U8279 (N_8279,N_7978,N_7666);
nand U8280 (N_8280,N_7083,N_7646);
nand U8281 (N_8281,N_7497,N_7502);
or U8282 (N_8282,N_7243,N_7074);
xnor U8283 (N_8283,N_7538,N_7964);
xnor U8284 (N_8284,N_7982,N_7241);
and U8285 (N_8285,N_7535,N_7459);
and U8286 (N_8286,N_7749,N_7118);
and U8287 (N_8287,N_7186,N_7391);
and U8288 (N_8288,N_7251,N_7147);
nor U8289 (N_8289,N_7220,N_7491);
or U8290 (N_8290,N_7667,N_7062);
xnor U8291 (N_8291,N_7466,N_7600);
nand U8292 (N_8292,N_7125,N_7815);
and U8293 (N_8293,N_7362,N_7208);
nor U8294 (N_8294,N_7176,N_7798);
or U8295 (N_8295,N_7311,N_7396);
xor U8296 (N_8296,N_7955,N_7771);
xor U8297 (N_8297,N_7231,N_7114);
nor U8298 (N_8298,N_7737,N_7371);
and U8299 (N_8299,N_7254,N_7678);
or U8300 (N_8300,N_7164,N_7545);
nor U8301 (N_8301,N_7774,N_7642);
or U8302 (N_8302,N_7596,N_7694);
nor U8303 (N_8303,N_7776,N_7136);
and U8304 (N_8304,N_7734,N_7531);
nor U8305 (N_8305,N_7986,N_7783);
and U8306 (N_8306,N_7637,N_7829);
or U8307 (N_8307,N_7811,N_7159);
nor U8308 (N_8308,N_7315,N_7052);
nand U8309 (N_8309,N_7020,N_7732);
nand U8310 (N_8310,N_7339,N_7818);
nand U8311 (N_8311,N_7193,N_7180);
xor U8312 (N_8312,N_7269,N_7718);
xnor U8313 (N_8313,N_7940,N_7444);
nor U8314 (N_8314,N_7956,N_7742);
nand U8315 (N_8315,N_7021,N_7690);
nor U8316 (N_8316,N_7919,N_7392);
or U8317 (N_8317,N_7842,N_7521);
nor U8318 (N_8318,N_7973,N_7185);
nor U8319 (N_8319,N_7035,N_7805);
or U8320 (N_8320,N_7613,N_7838);
nor U8321 (N_8321,N_7198,N_7580);
or U8322 (N_8322,N_7356,N_7454);
and U8323 (N_8323,N_7468,N_7975);
xnor U8324 (N_8324,N_7512,N_7399);
nand U8325 (N_8325,N_7699,N_7131);
or U8326 (N_8326,N_7872,N_7764);
or U8327 (N_8327,N_7301,N_7041);
and U8328 (N_8328,N_7340,N_7849);
or U8329 (N_8329,N_7071,N_7772);
xor U8330 (N_8330,N_7348,N_7469);
nand U8331 (N_8331,N_7280,N_7293);
nor U8332 (N_8332,N_7635,N_7837);
xnor U8333 (N_8333,N_7439,N_7636);
nand U8334 (N_8334,N_7733,N_7951);
nor U8335 (N_8335,N_7930,N_7256);
and U8336 (N_8336,N_7343,N_7451);
and U8337 (N_8337,N_7086,N_7948);
nand U8338 (N_8338,N_7079,N_7726);
nor U8339 (N_8339,N_7972,N_7904);
xnor U8340 (N_8340,N_7821,N_7207);
xnor U8341 (N_8341,N_7403,N_7584);
or U8342 (N_8342,N_7711,N_7412);
nand U8343 (N_8343,N_7305,N_7397);
and U8344 (N_8344,N_7911,N_7817);
and U8345 (N_8345,N_7622,N_7051);
or U8346 (N_8346,N_7823,N_7730);
nand U8347 (N_8347,N_7789,N_7329);
and U8348 (N_8348,N_7437,N_7386);
nor U8349 (N_8349,N_7040,N_7572);
or U8350 (N_8350,N_7876,N_7345);
nor U8351 (N_8351,N_7481,N_7381);
nor U8352 (N_8352,N_7019,N_7058);
and U8353 (N_8353,N_7063,N_7576);
nor U8354 (N_8354,N_7873,N_7470);
nor U8355 (N_8355,N_7566,N_7202);
nor U8356 (N_8356,N_7323,N_7793);
nor U8357 (N_8357,N_7084,N_7859);
xor U8358 (N_8358,N_7687,N_7078);
xnor U8359 (N_8359,N_7053,N_7698);
nand U8360 (N_8360,N_7465,N_7146);
or U8361 (N_8361,N_7547,N_7092);
and U8362 (N_8362,N_7602,N_7900);
xor U8363 (N_8363,N_7638,N_7977);
xor U8364 (N_8364,N_7592,N_7997);
nand U8365 (N_8365,N_7965,N_7569);
nor U8366 (N_8366,N_7927,N_7133);
and U8367 (N_8367,N_7659,N_7944);
nand U8368 (N_8368,N_7335,N_7182);
xor U8369 (N_8369,N_7757,N_7797);
nand U8370 (N_8370,N_7790,N_7738);
and U8371 (N_8371,N_7150,N_7708);
nor U8372 (N_8372,N_7286,N_7937);
or U8373 (N_8373,N_7633,N_7029);
or U8374 (N_8374,N_7441,N_7172);
nor U8375 (N_8375,N_7649,N_7274);
nor U8376 (N_8376,N_7014,N_7987);
or U8377 (N_8377,N_7679,N_7731);
nor U8378 (N_8378,N_7363,N_7036);
or U8379 (N_8379,N_7373,N_7240);
and U8380 (N_8380,N_7917,N_7719);
or U8381 (N_8381,N_7753,N_7314);
or U8382 (N_8382,N_7799,N_7890);
nand U8383 (N_8383,N_7389,N_7217);
nand U8384 (N_8384,N_7205,N_7826);
nor U8385 (N_8385,N_7108,N_7270);
and U8386 (N_8386,N_7287,N_7901);
xor U8387 (N_8387,N_7232,N_7990);
xor U8388 (N_8388,N_7750,N_7551);
xor U8389 (N_8389,N_7401,N_7560);
or U8390 (N_8390,N_7390,N_7832);
or U8391 (N_8391,N_7568,N_7225);
nor U8392 (N_8392,N_7804,N_7387);
or U8393 (N_8393,N_7276,N_7144);
nor U8394 (N_8394,N_7695,N_7218);
and U8395 (N_8395,N_7745,N_7523);
nor U8396 (N_8396,N_7152,N_7214);
or U8397 (N_8397,N_7668,N_7607);
nand U8398 (N_8398,N_7026,N_7122);
or U8399 (N_8399,N_7598,N_7701);
nor U8400 (N_8400,N_7618,N_7717);
and U8401 (N_8401,N_7500,N_7884);
nor U8402 (N_8402,N_7606,N_7994);
and U8403 (N_8403,N_7385,N_7456);
nor U8404 (N_8404,N_7880,N_7284);
or U8405 (N_8405,N_7947,N_7216);
and U8406 (N_8406,N_7509,N_7050);
nor U8407 (N_8407,N_7350,N_7475);
nor U8408 (N_8408,N_7094,N_7556);
and U8409 (N_8409,N_7075,N_7189);
nand U8410 (N_8410,N_7912,N_7448);
nand U8411 (N_8411,N_7537,N_7494);
nor U8412 (N_8412,N_7630,N_7024);
nand U8413 (N_8413,N_7993,N_7665);
or U8414 (N_8414,N_7042,N_7541);
xor U8415 (N_8415,N_7317,N_7747);
and U8416 (N_8416,N_7891,N_7688);
or U8417 (N_8417,N_7110,N_7629);
nand U8418 (N_8418,N_7046,N_7846);
or U8419 (N_8419,N_7702,N_7689);
xnor U8420 (N_8420,N_7686,N_7788);
and U8421 (N_8421,N_7472,N_7102);
nand U8422 (N_8422,N_7442,N_7358);
xnor U8423 (N_8423,N_7727,N_7942);
nor U8424 (N_8424,N_7796,N_7353);
nand U8425 (N_8425,N_7867,N_7235);
nand U8426 (N_8426,N_7331,N_7422);
xnor U8427 (N_8427,N_7861,N_7061);
or U8428 (N_8428,N_7179,N_7996);
nand U8429 (N_8429,N_7657,N_7376);
nor U8430 (N_8430,N_7171,N_7691);
xnor U8431 (N_8431,N_7073,N_7415);
xnor U8432 (N_8432,N_7001,N_7669);
or U8433 (N_8433,N_7055,N_7645);
nor U8434 (N_8434,N_7278,N_7617);
and U8435 (N_8435,N_7921,N_7913);
xor U8436 (N_8436,N_7419,N_7382);
nand U8437 (N_8437,N_7853,N_7184);
and U8438 (N_8438,N_7562,N_7407);
xor U8439 (N_8439,N_7499,N_7769);
nor U8440 (N_8440,N_7877,N_7452);
nor U8441 (N_8441,N_7784,N_7048);
or U8442 (N_8442,N_7713,N_7895);
xor U8443 (N_8443,N_7211,N_7585);
and U8444 (N_8444,N_7775,N_7261);
or U8445 (N_8445,N_7168,N_7988);
or U8446 (N_8446,N_7296,N_7573);
nor U8447 (N_8447,N_7751,N_7124);
xnor U8448 (N_8448,N_7008,N_7375);
or U8449 (N_8449,N_7920,N_7710);
and U8450 (N_8450,N_7918,N_7501);
or U8451 (N_8451,N_7395,N_7034);
or U8452 (N_8452,N_7174,N_7298);
or U8453 (N_8453,N_7765,N_7529);
nor U8454 (N_8454,N_7043,N_7262);
or U8455 (N_8455,N_7524,N_7045);
or U8456 (N_8456,N_7611,N_7504);
nand U8457 (N_8457,N_7604,N_7463);
nor U8458 (N_8458,N_7156,N_7378);
or U8459 (N_8459,N_7623,N_7739);
nand U8460 (N_8460,N_7309,N_7307);
nor U8461 (N_8461,N_7354,N_7716);
nor U8462 (N_8462,N_7057,N_7768);
nor U8463 (N_8463,N_7903,N_7303);
xor U8464 (N_8464,N_7095,N_7631);
nor U8465 (N_8465,N_7527,N_7004);
and U8466 (N_8466,N_7135,N_7729);
nor U8467 (N_8467,N_7447,N_7841);
nand U8468 (N_8468,N_7898,N_7574);
nand U8469 (N_8469,N_7762,N_7228);
and U8470 (N_8470,N_7814,N_7425);
or U8471 (N_8471,N_7722,N_7022);
and U8472 (N_8472,N_7936,N_7946);
xor U8473 (N_8473,N_7291,N_7603);
xnor U8474 (N_8474,N_7495,N_7587);
xnor U8475 (N_8475,N_7833,N_7482);
or U8476 (N_8476,N_7300,N_7770);
and U8477 (N_8477,N_7130,N_7170);
nor U8478 (N_8478,N_7239,N_7953);
nand U8479 (N_8479,N_7648,N_7960);
nor U8480 (N_8480,N_7313,N_7064);
xnor U8481 (N_8481,N_7112,N_7653);
nor U8482 (N_8482,N_7142,N_7368);
xnor U8483 (N_8483,N_7120,N_7429);
xnor U8484 (N_8484,N_7767,N_7883);
xnor U8485 (N_8485,N_7728,N_7519);
and U8486 (N_8486,N_7487,N_7476);
and U8487 (N_8487,N_7575,N_7484);
nor U8488 (N_8488,N_7480,N_7402);
and U8489 (N_8489,N_7864,N_7792);
nand U8490 (N_8490,N_7160,N_7925);
and U8491 (N_8491,N_7578,N_7868);
and U8492 (N_8492,N_7139,N_7778);
nor U8493 (N_8493,N_7998,N_7089);
and U8494 (N_8494,N_7748,N_7954);
or U8495 (N_8495,N_7854,N_7813);
nand U8496 (N_8496,N_7581,N_7825);
or U8497 (N_8497,N_7865,N_7091);
or U8498 (N_8498,N_7539,N_7516);
nand U8499 (N_8499,N_7267,N_7652);
nand U8500 (N_8500,N_7076,N_7035);
and U8501 (N_8501,N_7150,N_7200);
nor U8502 (N_8502,N_7766,N_7811);
or U8503 (N_8503,N_7488,N_7502);
xor U8504 (N_8504,N_7007,N_7293);
nand U8505 (N_8505,N_7159,N_7945);
or U8506 (N_8506,N_7140,N_7318);
xor U8507 (N_8507,N_7354,N_7534);
or U8508 (N_8508,N_7004,N_7777);
or U8509 (N_8509,N_7969,N_7027);
nor U8510 (N_8510,N_7275,N_7813);
or U8511 (N_8511,N_7721,N_7864);
and U8512 (N_8512,N_7761,N_7736);
nand U8513 (N_8513,N_7689,N_7959);
xnor U8514 (N_8514,N_7233,N_7941);
nor U8515 (N_8515,N_7920,N_7358);
nand U8516 (N_8516,N_7568,N_7091);
nor U8517 (N_8517,N_7618,N_7152);
and U8518 (N_8518,N_7210,N_7654);
or U8519 (N_8519,N_7352,N_7112);
xor U8520 (N_8520,N_7993,N_7667);
xor U8521 (N_8521,N_7674,N_7399);
nor U8522 (N_8522,N_7224,N_7691);
or U8523 (N_8523,N_7157,N_7867);
nand U8524 (N_8524,N_7988,N_7115);
nand U8525 (N_8525,N_7091,N_7394);
xor U8526 (N_8526,N_7574,N_7448);
or U8527 (N_8527,N_7658,N_7004);
and U8528 (N_8528,N_7191,N_7259);
xor U8529 (N_8529,N_7076,N_7752);
or U8530 (N_8530,N_7314,N_7385);
xnor U8531 (N_8531,N_7882,N_7879);
or U8532 (N_8532,N_7908,N_7040);
xnor U8533 (N_8533,N_7197,N_7435);
nor U8534 (N_8534,N_7494,N_7540);
nand U8535 (N_8535,N_7419,N_7708);
xnor U8536 (N_8536,N_7229,N_7525);
xnor U8537 (N_8537,N_7448,N_7038);
or U8538 (N_8538,N_7739,N_7213);
nand U8539 (N_8539,N_7107,N_7899);
xnor U8540 (N_8540,N_7367,N_7675);
and U8541 (N_8541,N_7692,N_7245);
xnor U8542 (N_8542,N_7730,N_7244);
and U8543 (N_8543,N_7909,N_7894);
nand U8544 (N_8544,N_7060,N_7831);
or U8545 (N_8545,N_7020,N_7463);
or U8546 (N_8546,N_7824,N_7243);
or U8547 (N_8547,N_7480,N_7772);
and U8548 (N_8548,N_7178,N_7629);
or U8549 (N_8549,N_7679,N_7036);
nor U8550 (N_8550,N_7993,N_7182);
nor U8551 (N_8551,N_7766,N_7441);
xnor U8552 (N_8552,N_7975,N_7230);
xnor U8553 (N_8553,N_7462,N_7021);
and U8554 (N_8554,N_7659,N_7648);
nand U8555 (N_8555,N_7351,N_7862);
and U8556 (N_8556,N_7257,N_7689);
and U8557 (N_8557,N_7618,N_7586);
nand U8558 (N_8558,N_7587,N_7217);
xor U8559 (N_8559,N_7550,N_7444);
nand U8560 (N_8560,N_7278,N_7079);
xor U8561 (N_8561,N_7635,N_7530);
and U8562 (N_8562,N_7977,N_7747);
nand U8563 (N_8563,N_7175,N_7089);
nor U8564 (N_8564,N_7152,N_7603);
xor U8565 (N_8565,N_7368,N_7930);
nor U8566 (N_8566,N_7766,N_7366);
nor U8567 (N_8567,N_7604,N_7205);
nor U8568 (N_8568,N_7457,N_7109);
or U8569 (N_8569,N_7245,N_7341);
and U8570 (N_8570,N_7837,N_7788);
nand U8571 (N_8571,N_7921,N_7455);
xnor U8572 (N_8572,N_7392,N_7290);
nor U8573 (N_8573,N_7118,N_7064);
nor U8574 (N_8574,N_7780,N_7311);
or U8575 (N_8575,N_7966,N_7311);
and U8576 (N_8576,N_7561,N_7944);
nor U8577 (N_8577,N_7372,N_7792);
or U8578 (N_8578,N_7220,N_7955);
nor U8579 (N_8579,N_7429,N_7662);
or U8580 (N_8580,N_7228,N_7103);
or U8581 (N_8581,N_7701,N_7594);
or U8582 (N_8582,N_7261,N_7065);
and U8583 (N_8583,N_7823,N_7988);
xnor U8584 (N_8584,N_7753,N_7935);
or U8585 (N_8585,N_7262,N_7089);
and U8586 (N_8586,N_7956,N_7857);
nor U8587 (N_8587,N_7056,N_7525);
and U8588 (N_8588,N_7942,N_7640);
xor U8589 (N_8589,N_7311,N_7118);
and U8590 (N_8590,N_7115,N_7420);
and U8591 (N_8591,N_7818,N_7844);
nor U8592 (N_8592,N_7949,N_7078);
or U8593 (N_8593,N_7508,N_7821);
or U8594 (N_8594,N_7555,N_7791);
nand U8595 (N_8595,N_7825,N_7491);
nor U8596 (N_8596,N_7490,N_7272);
nand U8597 (N_8597,N_7524,N_7921);
xor U8598 (N_8598,N_7852,N_7479);
or U8599 (N_8599,N_7207,N_7772);
nor U8600 (N_8600,N_7022,N_7796);
xor U8601 (N_8601,N_7614,N_7685);
and U8602 (N_8602,N_7693,N_7313);
xor U8603 (N_8603,N_7408,N_7299);
nor U8604 (N_8604,N_7500,N_7038);
xor U8605 (N_8605,N_7541,N_7253);
or U8606 (N_8606,N_7630,N_7978);
nor U8607 (N_8607,N_7877,N_7260);
nor U8608 (N_8608,N_7211,N_7489);
nor U8609 (N_8609,N_7599,N_7059);
nor U8610 (N_8610,N_7801,N_7984);
or U8611 (N_8611,N_7653,N_7149);
xnor U8612 (N_8612,N_7690,N_7654);
and U8613 (N_8613,N_7394,N_7465);
nor U8614 (N_8614,N_7792,N_7514);
xnor U8615 (N_8615,N_7086,N_7905);
nor U8616 (N_8616,N_7490,N_7348);
xnor U8617 (N_8617,N_7486,N_7947);
or U8618 (N_8618,N_7399,N_7097);
xor U8619 (N_8619,N_7305,N_7533);
nand U8620 (N_8620,N_7720,N_7204);
xor U8621 (N_8621,N_7716,N_7195);
xnor U8622 (N_8622,N_7569,N_7732);
and U8623 (N_8623,N_7868,N_7648);
nor U8624 (N_8624,N_7246,N_7124);
and U8625 (N_8625,N_7524,N_7943);
xor U8626 (N_8626,N_7894,N_7585);
or U8627 (N_8627,N_7199,N_7619);
nor U8628 (N_8628,N_7964,N_7228);
nand U8629 (N_8629,N_7554,N_7771);
and U8630 (N_8630,N_7314,N_7347);
nand U8631 (N_8631,N_7019,N_7579);
nor U8632 (N_8632,N_7208,N_7729);
and U8633 (N_8633,N_7166,N_7764);
xor U8634 (N_8634,N_7934,N_7754);
xnor U8635 (N_8635,N_7832,N_7239);
nor U8636 (N_8636,N_7016,N_7747);
xnor U8637 (N_8637,N_7866,N_7159);
nand U8638 (N_8638,N_7224,N_7934);
nand U8639 (N_8639,N_7431,N_7193);
and U8640 (N_8640,N_7413,N_7328);
nand U8641 (N_8641,N_7719,N_7055);
nand U8642 (N_8642,N_7317,N_7573);
and U8643 (N_8643,N_7546,N_7687);
xnor U8644 (N_8644,N_7909,N_7248);
xnor U8645 (N_8645,N_7662,N_7780);
or U8646 (N_8646,N_7603,N_7912);
nand U8647 (N_8647,N_7082,N_7438);
and U8648 (N_8648,N_7243,N_7269);
nor U8649 (N_8649,N_7867,N_7036);
nor U8650 (N_8650,N_7216,N_7150);
nor U8651 (N_8651,N_7823,N_7484);
and U8652 (N_8652,N_7880,N_7915);
and U8653 (N_8653,N_7077,N_7934);
nand U8654 (N_8654,N_7992,N_7115);
or U8655 (N_8655,N_7482,N_7780);
nand U8656 (N_8656,N_7072,N_7982);
xnor U8657 (N_8657,N_7124,N_7452);
nor U8658 (N_8658,N_7420,N_7369);
nor U8659 (N_8659,N_7001,N_7744);
xnor U8660 (N_8660,N_7985,N_7683);
and U8661 (N_8661,N_7525,N_7624);
nand U8662 (N_8662,N_7484,N_7396);
nand U8663 (N_8663,N_7645,N_7509);
xnor U8664 (N_8664,N_7969,N_7086);
nor U8665 (N_8665,N_7032,N_7731);
nor U8666 (N_8666,N_7404,N_7291);
xor U8667 (N_8667,N_7733,N_7993);
nand U8668 (N_8668,N_7245,N_7496);
xnor U8669 (N_8669,N_7910,N_7842);
nor U8670 (N_8670,N_7459,N_7516);
nand U8671 (N_8671,N_7390,N_7291);
xor U8672 (N_8672,N_7767,N_7612);
nand U8673 (N_8673,N_7522,N_7687);
and U8674 (N_8674,N_7430,N_7937);
nor U8675 (N_8675,N_7630,N_7400);
and U8676 (N_8676,N_7788,N_7747);
or U8677 (N_8677,N_7069,N_7997);
xnor U8678 (N_8678,N_7652,N_7633);
nor U8679 (N_8679,N_7238,N_7830);
nor U8680 (N_8680,N_7094,N_7633);
and U8681 (N_8681,N_7105,N_7094);
or U8682 (N_8682,N_7082,N_7348);
xor U8683 (N_8683,N_7761,N_7886);
nor U8684 (N_8684,N_7523,N_7582);
nand U8685 (N_8685,N_7068,N_7428);
or U8686 (N_8686,N_7328,N_7392);
or U8687 (N_8687,N_7321,N_7209);
and U8688 (N_8688,N_7366,N_7906);
or U8689 (N_8689,N_7946,N_7679);
nor U8690 (N_8690,N_7388,N_7197);
xor U8691 (N_8691,N_7879,N_7363);
nor U8692 (N_8692,N_7182,N_7553);
xor U8693 (N_8693,N_7713,N_7068);
xor U8694 (N_8694,N_7483,N_7004);
xnor U8695 (N_8695,N_7530,N_7332);
or U8696 (N_8696,N_7911,N_7846);
nand U8697 (N_8697,N_7561,N_7623);
and U8698 (N_8698,N_7988,N_7465);
nor U8699 (N_8699,N_7985,N_7087);
and U8700 (N_8700,N_7028,N_7529);
nor U8701 (N_8701,N_7561,N_7376);
nand U8702 (N_8702,N_7507,N_7684);
and U8703 (N_8703,N_7075,N_7085);
nor U8704 (N_8704,N_7002,N_7689);
nor U8705 (N_8705,N_7634,N_7494);
or U8706 (N_8706,N_7397,N_7280);
xor U8707 (N_8707,N_7046,N_7708);
nor U8708 (N_8708,N_7227,N_7146);
and U8709 (N_8709,N_7707,N_7185);
and U8710 (N_8710,N_7965,N_7332);
nand U8711 (N_8711,N_7318,N_7685);
and U8712 (N_8712,N_7349,N_7644);
or U8713 (N_8713,N_7642,N_7582);
nand U8714 (N_8714,N_7907,N_7508);
and U8715 (N_8715,N_7649,N_7826);
and U8716 (N_8716,N_7095,N_7385);
and U8717 (N_8717,N_7922,N_7622);
or U8718 (N_8718,N_7130,N_7214);
nand U8719 (N_8719,N_7398,N_7373);
and U8720 (N_8720,N_7950,N_7601);
nand U8721 (N_8721,N_7780,N_7964);
nor U8722 (N_8722,N_7391,N_7433);
nand U8723 (N_8723,N_7398,N_7191);
nor U8724 (N_8724,N_7838,N_7305);
nand U8725 (N_8725,N_7505,N_7564);
nand U8726 (N_8726,N_7694,N_7289);
and U8727 (N_8727,N_7295,N_7660);
xor U8728 (N_8728,N_7944,N_7026);
xor U8729 (N_8729,N_7948,N_7627);
nand U8730 (N_8730,N_7150,N_7605);
xor U8731 (N_8731,N_7732,N_7683);
xnor U8732 (N_8732,N_7041,N_7556);
and U8733 (N_8733,N_7306,N_7764);
nor U8734 (N_8734,N_7342,N_7654);
nor U8735 (N_8735,N_7823,N_7631);
xnor U8736 (N_8736,N_7268,N_7784);
nand U8737 (N_8737,N_7500,N_7098);
nand U8738 (N_8738,N_7437,N_7124);
xor U8739 (N_8739,N_7885,N_7214);
and U8740 (N_8740,N_7989,N_7831);
nand U8741 (N_8741,N_7434,N_7430);
nor U8742 (N_8742,N_7921,N_7795);
nand U8743 (N_8743,N_7562,N_7577);
nor U8744 (N_8744,N_7689,N_7648);
xor U8745 (N_8745,N_7552,N_7049);
or U8746 (N_8746,N_7319,N_7301);
xor U8747 (N_8747,N_7284,N_7401);
or U8748 (N_8748,N_7240,N_7867);
nand U8749 (N_8749,N_7819,N_7708);
or U8750 (N_8750,N_7333,N_7776);
nor U8751 (N_8751,N_7619,N_7110);
nor U8752 (N_8752,N_7559,N_7304);
nor U8753 (N_8753,N_7637,N_7483);
and U8754 (N_8754,N_7930,N_7523);
nand U8755 (N_8755,N_7704,N_7631);
xnor U8756 (N_8756,N_7709,N_7873);
xnor U8757 (N_8757,N_7288,N_7296);
or U8758 (N_8758,N_7174,N_7878);
nor U8759 (N_8759,N_7418,N_7417);
or U8760 (N_8760,N_7982,N_7642);
xnor U8761 (N_8761,N_7504,N_7663);
nor U8762 (N_8762,N_7933,N_7529);
nor U8763 (N_8763,N_7676,N_7228);
or U8764 (N_8764,N_7605,N_7485);
nor U8765 (N_8765,N_7058,N_7863);
and U8766 (N_8766,N_7601,N_7013);
nand U8767 (N_8767,N_7110,N_7596);
nor U8768 (N_8768,N_7923,N_7744);
nand U8769 (N_8769,N_7327,N_7713);
or U8770 (N_8770,N_7659,N_7307);
or U8771 (N_8771,N_7266,N_7033);
xor U8772 (N_8772,N_7423,N_7607);
and U8773 (N_8773,N_7382,N_7876);
nor U8774 (N_8774,N_7320,N_7522);
xor U8775 (N_8775,N_7073,N_7244);
or U8776 (N_8776,N_7425,N_7180);
or U8777 (N_8777,N_7999,N_7167);
or U8778 (N_8778,N_7999,N_7633);
xnor U8779 (N_8779,N_7705,N_7563);
nand U8780 (N_8780,N_7452,N_7139);
xnor U8781 (N_8781,N_7979,N_7859);
xor U8782 (N_8782,N_7041,N_7088);
xnor U8783 (N_8783,N_7914,N_7810);
and U8784 (N_8784,N_7702,N_7158);
or U8785 (N_8785,N_7066,N_7832);
or U8786 (N_8786,N_7367,N_7402);
nor U8787 (N_8787,N_7637,N_7189);
xor U8788 (N_8788,N_7058,N_7013);
or U8789 (N_8789,N_7666,N_7902);
or U8790 (N_8790,N_7627,N_7380);
xor U8791 (N_8791,N_7615,N_7287);
xnor U8792 (N_8792,N_7578,N_7437);
or U8793 (N_8793,N_7786,N_7616);
and U8794 (N_8794,N_7051,N_7638);
or U8795 (N_8795,N_7730,N_7917);
or U8796 (N_8796,N_7866,N_7450);
nand U8797 (N_8797,N_7803,N_7683);
nand U8798 (N_8798,N_7566,N_7327);
nor U8799 (N_8799,N_7438,N_7143);
nand U8800 (N_8800,N_7128,N_7855);
nor U8801 (N_8801,N_7137,N_7218);
nor U8802 (N_8802,N_7489,N_7770);
nand U8803 (N_8803,N_7223,N_7126);
nand U8804 (N_8804,N_7646,N_7824);
xnor U8805 (N_8805,N_7815,N_7247);
and U8806 (N_8806,N_7365,N_7366);
nand U8807 (N_8807,N_7741,N_7359);
and U8808 (N_8808,N_7875,N_7530);
nor U8809 (N_8809,N_7030,N_7999);
nand U8810 (N_8810,N_7696,N_7225);
nor U8811 (N_8811,N_7827,N_7321);
or U8812 (N_8812,N_7687,N_7353);
xnor U8813 (N_8813,N_7609,N_7703);
xor U8814 (N_8814,N_7318,N_7248);
nand U8815 (N_8815,N_7454,N_7139);
and U8816 (N_8816,N_7963,N_7824);
xor U8817 (N_8817,N_7391,N_7987);
xnor U8818 (N_8818,N_7529,N_7037);
and U8819 (N_8819,N_7875,N_7865);
nor U8820 (N_8820,N_7010,N_7400);
or U8821 (N_8821,N_7071,N_7063);
xor U8822 (N_8822,N_7269,N_7290);
or U8823 (N_8823,N_7936,N_7299);
or U8824 (N_8824,N_7808,N_7566);
xor U8825 (N_8825,N_7174,N_7385);
and U8826 (N_8826,N_7546,N_7376);
or U8827 (N_8827,N_7932,N_7909);
nor U8828 (N_8828,N_7188,N_7234);
nor U8829 (N_8829,N_7856,N_7450);
xor U8830 (N_8830,N_7731,N_7705);
nand U8831 (N_8831,N_7304,N_7139);
xnor U8832 (N_8832,N_7798,N_7587);
xor U8833 (N_8833,N_7200,N_7484);
and U8834 (N_8834,N_7673,N_7334);
nand U8835 (N_8835,N_7728,N_7722);
xnor U8836 (N_8836,N_7867,N_7736);
nand U8837 (N_8837,N_7618,N_7300);
xor U8838 (N_8838,N_7196,N_7729);
nor U8839 (N_8839,N_7261,N_7401);
xnor U8840 (N_8840,N_7822,N_7724);
and U8841 (N_8841,N_7238,N_7506);
or U8842 (N_8842,N_7597,N_7385);
or U8843 (N_8843,N_7030,N_7474);
and U8844 (N_8844,N_7054,N_7201);
xnor U8845 (N_8845,N_7779,N_7305);
xor U8846 (N_8846,N_7531,N_7298);
nor U8847 (N_8847,N_7684,N_7233);
or U8848 (N_8848,N_7251,N_7686);
nand U8849 (N_8849,N_7192,N_7959);
xnor U8850 (N_8850,N_7401,N_7391);
nand U8851 (N_8851,N_7895,N_7992);
xor U8852 (N_8852,N_7817,N_7842);
and U8853 (N_8853,N_7145,N_7425);
xor U8854 (N_8854,N_7468,N_7608);
and U8855 (N_8855,N_7001,N_7385);
xnor U8856 (N_8856,N_7458,N_7170);
nor U8857 (N_8857,N_7393,N_7948);
nor U8858 (N_8858,N_7036,N_7983);
nand U8859 (N_8859,N_7331,N_7410);
or U8860 (N_8860,N_7752,N_7721);
xor U8861 (N_8861,N_7259,N_7031);
nand U8862 (N_8862,N_7848,N_7562);
and U8863 (N_8863,N_7225,N_7727);
xor U8864 (N_8864,N_7577,N_7922);
nor U8865 (N_8865,N_7064,N_7285);
nor U8866 (N_8866,N_7304,N_7719);
nand U8867 (N_8867,N_7869,N_7072);
nand U8868 (N_8868,N_7909,N_7035);
or U8869 (N_8869,N_7003,N_7585);
nand U8870 (N_8870,N_7695,N_7286);
nor U8871 (N_8871,N_7023,N_7299);
nand U8872 (N_8872,N_7897,N_7370);
and U8873 (N_8873,N_7063,N_7029);
and U8874 (N_8874,N_7164,N_7713);
or U8875 (N_8875,N_7071,N_7094);
nand U8876 (N_8876,N_7470,N_7848);
xor U8877 (N_8877,N_7317,N_7248);
xor U8878 (N_8878,N_7724,N_7787);
and U8879 (N_8879,N_7353,N_7069);
and U8880 (N_8880,N_7605,N_7555);
xor U8881 (N_8881,N_7829,N_7978);
xor U8882 (N_8882,N_7245,N_7911);
or U8883 (N_8883,N_7099,N_7609);
and U8884 (N_8884,N_7842,N_7632);
and U8885 (N_8885,N_7136,N_7893);
nand U8886 (N_8886,N_7663,N_7002);
nand U8887 (N_8887,N_7451,N_7705);
xor U8888 (N_8888,N_7245,N_7012);
nor U8889 (N_8889,N_7558,N_7541);
or U8890 (N_8890,N_7951,N_7900);
xor U8891 (N_8891,N_7214,N_7633);
nor U8892 (N_8892,N_7905,N_7068);
nor U8893 (N_8893,N_7505,N_7550);
xor U8894 (N_8894,N_7642,N_7649);
nand U8895 (N_8895,N_7366,N_7521);
or U8896 (N_8896,N_7984,N_7528);
and U8897 (N_8897,N_7452,N_7426);
or U8898 (N_8898,N_7623,N_7997);
xor U8899 (N_8899,N_7322,N_7395);
and U8900 (N_8900,N_7865,N_7467);
and U8901 (N_8901,N_7571,N_7995);
nand U8902 (N_8902,N_7779,N_7762);
xnor U8903 (N_8903,N_7107,N_7437);
nor U8904 (N_8904,N_7899,N_7763);
or U8905 (N_8905,N_7084,N_7525);
xor U8906 (N_8906,N_7533,N_7766);
or U8907 (N_8907,N_7957,N_7145);
xor U8908 (N_8908,N_7395,N_7229);
xor U8909 (N_8909,N_7400,N_7153);
or U8910 (N_8910,N_7313,N_7221);
nand U8911 (N_8911,N_7494,N_7826);
nand U8912 (N_8912,N_7708,N_7570);
nor U8913 (N_8913,N_7453,N_7854);
or U8914 (N_8914,N_7548,N_7202);
nand U8915 (N_8915,N_7785,N_7649);
and U8916 (N_8916,N_7686,N_7227);
nor U8917 (N_8917,N_7093,N_7465);
xor U8918 (N_8918,N_7573,N_7128);
nor U8919 (N_8919,N_7571,N_7717);
and U8920 (N_8920,N_7415,N_7041);
and U8921 (N_8921,N_7326,N_7036);
and U8922 (N_8922,N_7258,N_7335);
and U8923 (N_8923,N_7991,N_7781);
xor U8924 (N_8924,N_7332,N_7128);
nor U8925 (N_8925,N_7088,N_7492);
nor U8926 (N_8926,N_7044,N_7850);
nor U8927 (N_8927,N_7058,N_7304);
or U8928 (N_8928,N_7970,N_7131);
or U8929 (N_8929,N_7197,N_7427);
nand U8930 (N_8930,N_7110,N_7389);
and U8931 (N_8931,N_7709,N_7316);
nand U8932 (N_8932,N_7307,N_7065);
and U8933 (N_8933,N_7223,N_7801);
and U8934 (N_8934,N_7774,N_7620);
and U8935 (N_8935,N_7861,N_7704);
and U8936 (N_8936,N_7546,N_7955);
nor U8937 (N_8937,N_7493,N_7826);
or U8938 (N_8938,N_7733,N_7360);
nand U8939 (N_8939,N_7850,N_7827);
xor U8940 (N_8940,N_7139,N_7893);
nor U8941 (N_8941,N_7616,N_7611);
or U8942 (N_8942,N_7984,N_7922);
and U8943 (N_8943,N_7131,N_7754);
xnor U8944 (N_8944,N_7619,N_7174);
xor U8945 (N_8945,N_7642,N_7097);
nand U8946 (N_8946,N_7765,N_7485);
and U8947 (N_8947,N_7834,N_7630);
nand U8948 (N_8948,N_7626,N_7237);
and U8949 (N_8949,N_7621,N_7305);
nand U8950 (N_8950,N_7823,N_7764);
and U8951 (N_8951,N_7908,N_7412);
nand U8952 (N_8952,N_7232,N_7776);
or U8953 (N_8953,N_7472,N_7812);
xnor U8954 (N_8954,N_7212,N_7161);
and U8955 (N_8955,N_7789,N_7315);
or U8956 (N_8956,N_7154,N_7058);
xnor U8957 (N_8957,N_7444,N_7481);
and U8958 (N_8958,N_7515,N_7686);
or U8959 (N_8959,N_7163,N_7159);
xnor U8960 (N_8960,N_7263,N_7991);
or U8961 (N_8961,N_7072,N_7319);
nor U8962 (N_8962,N_7025,N_7803);
nor U8963 (N_8963,N_7659,N_7622);
or U8964 (N_8964,N_7158,N_7220);
xnor U8965 (N_8965,N_7179,N_7328);
xor U8966 (N_8966,N_7583,N_7370);
or U8967 (N_8967,N_7023,N_7566);
and U8968 (N_8968,N_7599,N_7893);
nand U8969 (N_8969,N_7885,N_7537);
and U8970 (N_8970,N_7683,N_7418);
and U8971 (N_8971,N_7882,N_7324);
or U8972 (N_8972,N_7359,N_7976);
xnor U8973 (N_8973,N_7032,N_7818);
xnor U8974 (N_8974,N_7674,N_7684);
or U8975 (N_8975,N_7816,N_7681);
nor U8976 (N_8976,N_7848,N_7315);
or U8977 (N_8977,N_7094,N_7313);
xnor U8978 (N_8978,N_7057,N_7506);
nor U8979 (N_8979,N_7223,N_7808);
nor U8980 (N_8980,N_7219,N_7269);
nand U8981 (N_8981,N_7466,N_7986);
nand U8982 (N_8982,N_7854,N_7647);
nand U8983 (N_8983,N_7108,N_7365);
or U8984 (N_8984,N_7047,N_7924);
nand U8985 (N_8985,N_7360,N_7722);
nor U8986 (N_8986,N_7372,N_7064);
and U8987 (N_8987,N_7984,N_7354);
nand U8988 (N_8988,N_7238,N_7106);
nor U8989 (N_8989,N_7163,N_7617);
and U8990 (N_8990,N_7407,N_7624);
nand U8991 (N_8991,N_7182,N_7831);
or U8992 (N_8992,N_7364,N_7314);
nor U8993 (N_8993,N_7995,N_7858);
nand U8994 (N_8994,N_7979,N_7134);
nor U8995 (N_8995,N_7574,N_7473);
or U8996 (N_8996,N_7954,N_7176);
nand U8997 (N_8997,N_7143,N_7140);
and U8998 (N_8998,N_7584,N_7961);
and U8999 (N_8999,N_7453,N_7812);
and U9000 (N_9000,N_8763,N_8465);
xnor U9001 (N_9001,N_8463,N_8908);
xnor U9002 (N_9002,N_8687,N_8565);
and U9003 (N_9003,N_8830,N_8601);
nand U9004 (N_9004,N_8958,N_8878);
or U9005 (N_9005,N_8652,N_8794);
and U9006 (N_9006,N_8433,N_8105);
or U9007 (N_9007,N_8654,N_8029);
or U9008 (N_9008,N_8183,N_8828);
xnor U9009 (N_9009,N_8765,N_8408);
nor U9010 (N_9010,N_8849,N_8955);
nor U9011 (N_9011,N_8422,N_8936);
xor U9012 (N_9012,N_8998,N_8815);
nor U9013 (N_9013,N_8742,N_8527);
nand U9014 (N_9014,N_8203,N_8412);
nand U9015 (N_9015,N_8109,N_8483);
or U9016 (N_9016,N_8631,N_8043);
and U9017 (N_9017,N_8773,N_8918);
nor U9018 (N_9018,N_8536,N_8666);
nor U9019 (N_9019,N_8395,N_8805);
nand U9020 (N_9020,N_8385,N_8801);
nor U9021 (N_9021,N_8197,N_8092);
nand U9022 (N_9022,N_8939,N_8295);
and U9023 (N_9023,N_8838,N_8270);
nor U9024 (N_9024,N_8829,N_8747);
nand U9025 (N_9025,N_8680,N_8358);
nand U9026 (N_9026,N_8056,N_8006);
xnor U9027 (N_9027,N_8480,N_8038);
and U9028 (N_9028,N_8702,N_8416);
or U9029 (N_9029,N_8984,N_8360);
nor U9030 (N_9030,N_8477,N_8079);
and U9031 (N_9031,N_8276,N_8032);
and U9032 (N_9032,N_8299,N_8825);
and U9033 (N_9033,N_8751,N_8640);
nor U9034 (N_9034,N_8639,N_8369);
xnor U9035 (N_9035,N_8133,N_8693);
and U9036 (N_9036,N_8629,N_8841);
and U9037 (N_9037,N_8608,N_8003);
and U9038 (N_9038,N_8610,N_8023);
nor U9039 (N_9039,N_8326,N_8641);
xnor U9040 (N_9040,N_8205,N_8852);
xnor U9041 (N_9041,N_8909,N_8864);
nand U9042 (N_9042,N_8267,N_8789);
xnor U9043 (N_9043,N_8835,N_8745);
nand U9044 (N_9044,N_8219,N_8040);
nand U9045 (N_9045,N_8668,N_8365);
xor U9046 (N_9046,N_8274,N_8927);
xor U9047 (N_9047,N_8869,N_8871);
and U9048 (N_9048,N_8158,N_8701);
nand U9049 (N_9049,N_8099,N_8401);
nor U9050 (N_9050,N_8308,N_8647);
and U9051 (N_9051,N_8978,N_8350);
xor U9052 (N_9052,N_8713,N_8626);
and U9053 (N_9053,N_8086,N_8009);
nand U9054 (N_9054,N_8265,N_8620);
xor U9055 (N_9055,N_8728,N_8923);
and U9056 (N_9056,N_8389,N_8275);
nand U9057 (N_9057,N_8934,N_8893);
and U9058 (N_9058,N_8147,N_8288);
and U9059 (N_9059,N_8272,N_8904);
xnor U9060 (N_9060,N_8187,N_8305);
or U9061 (N_9061,N_8714,N_8840);
or U9062 (N_9062,N_8195,N_8814);
nor U9063 (N_9063,N_8162,N_8069);
nor U9064 (N_9064,N_8057,N_8819);
or U9065 (N_9065,N_8129,N_8266);
and U9066 (N_9066,N_8026,N_8543);
and U9067 (N_9067,N_8286,N_8220);
nor U9068 (N_9068,N_8740,N_8769);
nor U9069 (N_9069,N_8222,N_8906);
or U9070 (N_9070,N_8604,N_8074);
nand U9071 (N_9071,N_8883,N_8607);
nand U9072 (N_9072,N_8466,N_8375);
nor U9073 (N_9073,N_8571,N_8336);
xor U9074 (N_9074,N_8039,N_8446);
xor U9075 (N_9075,N_8552,N_8068);
and U9076 (N_9076,N_8468,N_8847);
and U9077 (N_9077,N_8420,N_8432);
nor U9078 (N_9078,N_8021,N_8627);
nor U9079 (N_9079,N_8882,N_8381);
or U9080 (N_9080,N_8752,N_8064);
and U9081 (N_9081,N_8228,N_8212);
nand U9082 (N_9082,N_8171,N_8355);
and U9083 (N_9083,N_8614,N_8999);
nor U9084 (N_9084,N_8262,N_8083);
or U9085 (N_9085,N_8261,N_8136);
nor U9086 (N_9086,N_8470,N_8001);
nand U9087 (N_9087,N_8234,N_8844);
nor U9088 (N_9088,N_8020,N_8865);
and U9089 (N_9089,N_8863,N_8623);
xor U9090 (N_9090,N_8076,N_8634);
or U9091 (N_9091,N_8135,N_8758);
nand U9092 (N_9092,N_8502,N_8066);
xor U9093 (N_9093,N_8550,N_8532);
nor U9094 (N_9094,N_8720,N_8755);
xnor U9095 (N_9095,N_8901,N_8428);
or U9096 (N_9096,N_8448,N_8493);
and U9097 (N_9097,N_8596,N_8278);
or U9098 (N_9098,N_8160,N_8948);
nor U9099 (N_9099,N_8733,N_8012);
nor U9100 (N_9100,N_8979,N_8277);
and U9101 (N_9101,N_8941,N_8318);
nor U9102 (N_9102,N_8496,N_8748);
nor U9103 (N_9103,N_8879,N_8184);
nand U9104 (N_9104,N_8150,N_8762);
nand U9105 (N_9105,N_8264,N_8584);
and U9106 (N_9106,N_8378,N_8097);
and U9107 (N_9107,N_8132,N_8925);
nand U9108 (N_9108,N_8689,N_8174);
and U9109 (N_9109,N_8319,N_8642);
or U9110 (N_9110,N_8104,N_8866);
xor U9111 (N_9111,N_8192,N_8254);
nor U9112 (N_9112,N_8191,N_8089);
nand U9113 (N_9113,N_8581,N_8303);
nor U9114 (N_9114,N_8398,N_8250);
or U9115 (N_9115,N_8935,N_8000);
or U9116 (N_9116,N_8910,N_8294);
xnor U9117 (N_9117,N_8945,N_8157);
xor U9118 (N_9118,N_8193,N_8090);
and U9119 (N_9119,N_8972,N_8232);
and U9120 (N_9120,N_8479,N_8669);
or U9121 (N_9121,N_8062,N_8309);
nor U9122 (N_9122,N_8684,N_8874);
xor U9123 (N_9123,N_8506,N_8903);
and U9124 (N_9124,N_8795,N_8928);
nand U9125 (N_9125,N_8746,N_8737);
xor U9126 (N_9126,N_8558,N_8400);
xnor U9127 (N_9127,N_8321,N_8142);
xnor U9128 (N_9128,N_8427,N_8575);
nor U9129 (N_9129,N_8167,N_8644);
nand U9130 (N_9130,N_8606,N_8329);
and U9131 (N_9131,N_8987,N_8842);
nand U9132 (N_9132,N_8402,N_8813);
nand U9133 (N_9133,N_8512,N_8573);
and U9134 (N_9134,N_8485,N_8559);
xor U9135 (N_9135,N_8504,N_8215);
and U9136 (N_9136,N_8709,N_8230);
nand U9137 (N_9137,N_8824,N_8178);
xor U9138 (N_9138,N_8472,N_8605);
and U9139 (N_9139,N_8761,N_8233);
nand U9140 (N_9140,N_8990,N_8185);
or U9141 (N_9141,N_8384,N_8977);
or U9142 (N_9142,N_8087,N_8637);
nor U9143 (N_9143,N_8140,N_8499);
nor U9144 (N_9144,N_8764,N_8851);
xnor U9145 (N_9145,N_8985,N_8106);
xor U9146 (N_9146,N_8045,N_8033);
and U9147 (N_9147,N_8546,N_8341);
and U9148 (N_9148,N_8850,N_8165);
and U9149 (N_9149,N_8063,N_8523);
nor U9150 (N_9150,N_8912,N_8114);
nand U9151 (N_9151,N_8889,N_8247);
xnor U9152 (N_9152,N_8911,N_8723);
xnor U9153 (N_9153,N_8926,N_8330);
nand U9154 (N_9154,N_8658,N_8695);
and U9155 (N_9155,N_8123,N_8598);
nor U9156 (N_9156,N_8855,N_8947);
nand U9157 (N_9157,N_8796,N_8095);
nand U9158 (N_9158,N_8225,N_8685);
nor U9159 (N_9159,N_8860,N_8386);
xnor U9160 (N_9160,N_8311,N_8084);
or U9161 (N_9161,N_8018,N_8279);
nand U9162 (N_9162,N_8915,N_8121);
nand U9163 (N_9163,N_8218,N_8442);
nand U9164 (N_9164,N_8034,N_8963);
nor U9165 (N_9165,N_8488,N_8085);
nand U9166 (N_9166,N_8236,N_8213);
xnor U9167 (N_9167,N_8231,N_8455);
nor U9168 (N_9168,N_8253,N_8576);
or U9169 (N_9169,N_8522,N_8169);
xnor U9170 (N_9170,N_8244,N_8164);
or U9171 (N_9171,N_8214,N_8131);
or U9172 (N_9172,N_8370,N_8182);
or U9173 (N_9173,N_8356,N_8208);
nand U9174 (N_9174,N_8890,N_8014);
xor U9175 (N_9175,N_8611,N_8204);
nor U9176 (N_9176,N_8839,N_8656);
and U9177 (N_9177,N_8921,N_8715);
nand U9178 (N_9178,N_8027,N_8980);
nand U9179 (N_9179,N_8780,N_8199);
and U9180 (N_9180,N_8143,N_8539);
nand U9181 (N_9181,N_8544,N_8224);
and U9182 (N_9182,N_8593,N_8960);
nand U9183 (N_9183,N_8756,N_8916);
nor U9184 (N_9184,N_8562,N_8649);
nor U9185 (N_9185,N_8538,N_8597);
xnor U9186 (N_9186,N_8672,N_8609);
nor U9187 (N_9187,N_8120,N_8403);
xnor U9188 (N_9188,N_8240,N_8417);
and U9189 (N_9189,N_8809,N_8282);
nor U9190 (N_9190,N_8931,N_8717);
xnor U9191 (N_9191,N_8440,N_8675);
nor U9192 (N_9192,N_8591,N_8235);
or U9193 (N_9193,N_8877,N_8778);
nand U9194 (N_9194,N_8969,N_8834);
xnor U9195 (N_9195,N_8509,N_8798);
and U9196 (N_9196,N_8659,N_8206);
and U9197 (N_9197,N_8363,N_8704);
or U9198 (N_9198,N_8859,N_8210);
and U9199 (N_9199,N_8487,N_8388);
nor U9200 (N_9200,N_8655,N_8743);
or U9201 (N_9201,N_8667,N_8803);
nor U9202 (N_9202,N_8891,N_8202);
xnor U9203 (N_9203,N_8467,N_8807);
and U9204 (N_9204,N_8037,N_8445);
nand U9205 (N_9205,N_8643,N_8567);
or U9206 (N_9206,N_8741,N_8456);
nor U9207 (N_9207,N_8619,N_8585);
xor U9208 (N_9208,N_8082,N_8207);
or U9209 (N_9209,N_8574,N_8216);
and U9210 (N_9210,N_8699,N_8307);
or U9211 (N_9211,N_8390,N_8139);
or U9212 (N_9212,N_8117,N_8586);
nand U9213 (N_9213,N_8376,N_8489);
nand U9214 (N_9214,N_8423,N_8622);
xor U9215 (N_9215,N_8122,N_8382);
xnor U9216 (N_9216,N_8166,N_8661);
and U9217 (N_9217,N_8393,N_8359);
and U9218 (N_9218,N_8554,N_8320);
xor U9219 (N_9219,N_8854,N_8902);
nor U9220 (N_9220,N_8887,N_8880);
and U9221 (N_9221,N_8353,N_8943);
and U9222 (N_9222,N_8799,N_8334);
and U9223 (N_9223,N_8817,N_8418);
or U9224 (N_9224,N_8414,N_8580);
and U9225 (N_9225,N_8535,N_8868);
nor U9226 (N_9226,N_8507,N_8005);
nor U9227 (N_9227,N_8481,N_8735);
and U9228 (N_9228,N_8971,N_8494);
nand U9229 (N_9229,N_8149,N_8757);
or U9230 (N_9230,N_8399,N_8342);
or U9231 (N_9231,N_8929,N_8992);
nand U9232 (N_9232,N_8917,N_8621);
and U9233 (N_9233,N_8441,N_8042);
nand U9234 (N_9234,N_8510,N_8283);
and U9235 (N_9235,N_8325,N_8172);
xnor U9236 (N_9236,N_8974,N_8708);
xor U9237 (N_9237,N_8768,N_8674);
xor U9238 (N_9238,N_8239,N_8570);
and U9239 (N_9239,N_8345,N_8367);
xor U9240 (N_9240,N_8942,N_8410);
nor U9241 (N_9241,N_8010,N_8572);
or U9242 (N_9242,N_8556,N_8686);
and U9243 (N_9243,N_8331,N_8788);
and U9244 (N_9244,N_8624,N_8226);
nand U9245 (N_9245,N_8531,N_8263);
nand U9246 (N_9246,N_8616,N_8478);
and U9247 (N_9247,N_8221,N_8595);
or U9248 (N_9248,N_8938,N_8273);
nand U9249 (N_9249,N_8617,N_8453);
nor U9250 (N_9250,N_8566,N_8110);
or U9251 (N_9251,N_8227,N_8517);
and U9252 (N_9252,N_8404,N_8291);
nand U9253 (N_9253,N_8975,N_8898);
nand U9254 (N_9254,N_8340,N_8846);
nand U9255 (N_9255,N_8096,N_8579);
and U9256 (N_9256,N_8983,N_8051);
nor U9257 (N_9257,N_8997,N_8357);
and U9258 (N_9258,N_8258,N_8729);
and U9259 (N_9259,N_8793,N_8603);
and U9260 (N_9260,N_8521,N_8124);
and U9261 (N_9261,N_8430,N_8664);
xor U9262 (N_9262,N_8710,N_8787);
nor U9263 (N_9263,N_8323,N_8451);
xor U9264 (N_9264,N_8344,N_8332);
xnor U9265 (N_9265,N_8052,N_8924);
nand U9266 (N_9266,N_8612,N_8170);
nor U9267 (N_9267,N_8615,N_8304);
xor U9268 (N_9268,N_8257,N_8933);
nand U9269 (N_9269,N_8200,N_8553);
and U9270 (N_9270,N_8285,N_8186);
or U9271 (N_9271,N_8697,N_8520);
and U9272 (N_9272,N_8784,N_8491);
nor U9273 (N_9273,N_8670,N_8515);
nor U9274 (N_9274,N_8413,N_8726);
or U9275 (N_9275,N_8660,N_8542);
and U9276 (N_9276,N_8333,N_8061);
and U9277 (N_9277,N_8246,N_8671);
or U9278 (N_9278,N_8188,N_8770);
nand U9279 (N_9279,N_8271,N_8618);
nand U9280 (N_9280,N_8759,N_8049);
xor U9281 (N_9281,N_8754,N_8818);
xnor U9282 (N_9282,N_8783,N_8392);
nor U9283 (N_9283,N_8804,N_8127);
or U9284 (N_9284,N_8551,N_8537);
nor U9285 (N_9285,N_8377,N_8454);
nand U9286 (N_9286,N_8775,N_8705);
or U9287 (N_9287,N_8711,N_8462);
and U9288 (N_9288,N_8772,N_8657);
or U9289 (N_9289,N_8486,N_8973);
and U9290 (N_9290,N_8706,N_8716);
xor U9291 (N_9291,N_8959,N_8474);
xor U9292 (N_9292,N_8112,N_8490);
and U9293 (N_9293,N_8730,N_8346);
or U9294 (N_9294,N_8777,N_8907);
nor U9295 (N_9295,N_8540,N_8811);
nand U9296 (N_9296,N_8111,N_8460);
and U9297 (N_9297,N_8526,N_8719);
and U9298 (N_9298,N_8138,N_8217);
nand U9299 (N_9299,N_8141,N_8343);
and U9300 (N_9300,N_8368,N_8054);
nand U9301 (N_9301,N_8810,N_8081);
xor U9302 (N_9302,N_8568,N_8569);
nand U9303 (N_9303,N_8348,N_8004);
xnor U9304 (N_9304,N_8372,N_8189);
or U9305 (N_9305,N_8826,N_8080);
nand U9306 (N_9306,N_8970,N_8731);
nand U9307 (N_9307,N_8940,N_8177);
and U9308 (N_9308,N_8396,N_8802);
nor U9309 (N_9309,N_8508,N_8744);
nor U9310 (N_9310,N_8645,N_8774);
and U9311 (N_9311,N_8707,N_8545);
xor U9312 (N_9312,N_8019,N_8482);
xor U9313 (N_9313,N_8673,N_8518);
nor U9314 (N_9314,N_8310,N_8739);
nor U9315 (N_9315,N_8284,N_8352);
and U9316 (N_9316,N_8886,N_8881);
nand U9317 (N_9317,N_8296,N_8322);
nor U9318 (N_9318,N_8766,N_8436);
and U9319 (N_9319,N_8786,N_8435);
nand U9320 (N_9320,N_8862,N_8721);
xnor U9321 (N_9321,N_8424,N_8156);
and U9322 (N_9322,N_8949,N_8600);
and U9323 (N_9323,N_8443,N_8843);
and U9324 (N_9324,N_8152,N_8524);
xor U9325 (N_9325,N_8108,N_8415);
nor U9326 (N_9326,N_8391,N_8383);
or U9327 (N_9327,N_8920,N_8030);
nor U9328 (N_9328,N_8779,N_8560);
xnor U9329 (N_9329,N_8007,N_8176);
and U9330 (N_9330,N_8473,N_8944);
nand U9331 (N_9331,N_8146,N_8529);
and U9332 (N_9332,N_8314,N_8700);
and U9333 (N_9333,N_8301,N_8100);
and U9334 (N_9334,N_8137,N_8712);
and U9335 (N_9335,N_8349,N_8255);
and U9336 (N_9336,N_8471,N_8130);
nand U9337 (N_9337,N_8722,N_8895);
or U9338 (N_9338,N_8951,N_8892);
nand U9339 (N_9339,N_8444,N_8374);
or U9340 (N_9340,N_8613,N_8988);
nand U9341 (N_9341,N_8991,N_8053);
nand U9342 (N_9342,N_8434,N_8060);
nor U9343 (N_9343,N_8198,N_8767);
nor U9344 (N_9344,N_8548,N_8313);
nand U9345 (N_9345,N_8738,N_8025);
nand U9346 (N_9346,N_8590,N_8725);
or U9347 (N_9347,N_8387,N_8913);
nand U9348 (N_9348,N_8492,N_8290);
or U9349 (N_9349,N_8406,N_8930);
or U9350 (N_9350,N_8242,N_8126);
nand U9351 (N_9351,N_8946,N_8952);
or U9352 (N_9352,N_8914,N_8816);
nand U9353 (N_9353,N_8995,N_8858);
nor U9354 (N_9354,N_8259,N_8781);
nor U9355 (N_9355,N_8113,N_8996);
nand U9356 (N_9356,N_8328,N_8564);
or U9357 (N_9357,N_8024,N_8870);
or U9358 (N_9358,N_8447,N_8837);
and U9359 (N_9359,N_8651,N_8065);
nor U9360 (N_9360,N_8861,N_8058);
nor U9361 (N_9361,N_8820,N_8168);
nand U9362 (N_9362,N_8961,N_8268);
or U9363 (N_9363,N_8808,N_8646);
xnor U9364 (N_9364,N_8161,N_8505);
nor U9365 (N_9365,N_8962,N_8965);
nand U9366 (N_9366,N_8077,N_8409);
and U9367 (N_9367,N_8534,N_8662);
or U9368 (N_9368,N_8293,N_8116);
or U9369 (N_9369,N_8732,N_8461);
nand U9370 (N_9370,N_8822,N_8180);
xnor U9371 (N_9371,N_8677,N_8098);
or U9372 (N_9372,N_8469,N_8989);
xor U9373 (N_9373,N_8093,N_8557);
and U9374 (N_9374,N_8547,N_8450);
xnor U9375 (N_9375,N_8750,N_8280);
or U9376 (N_9376,N_8269,N_8982);
nor U9377 (N_9377,N_8753,N_8223);
or U9378 (N_9378,N_8679,N_8525);
xor U9379 (N_9379,N_8986,N_8703);
and U9380 (N_9380,N_8592,N_8792);
xor U9381 (N_9381,N_8957,N_8426);
nand U9382 (N_9382,N_8749,N_8599);
nor U9383 (N_9383,N_8583,N_8457);
nor U9384 (N_9384,N_8102,N_8602);
or U9385 (N_9385,N_8050,N_8589);
or U9386 (N_9386,N_8361,N_8201);
or U9387 (N_9387,N_8011,N_8885);
and U9388 (N_9388,N_8163,N_8394);
xnor U9389 (N_9389,N_8888,N_8541);
and U9390 (N_9390,N_8791,N_8800);
and U9391 (N_9391,N_8101,N_8256);
and U9392 (N_9392,N_8154,N_8252);
nor U9393 (N_9393,N_8683,N_8371);
nor U9394 (N_9394,N_8347,N_8153);
xor U9395 (N_9395,N_8932,N_8736);
nor U9396 (N_9396,N_8013,N_8628);
xor U9397 (N_9397,N_8873,N_8238);
nand U9398 (N_9398,N_8806,N_8790);
and U9399 (N_9399,N_8351,N_8727);
nand U9400 (N_9400,N_8823,N_8405);
xor U9401 (N_9401,N_8151,N_8561);
nand U9402 (N_9402,N_8976,N_8251);
or U9403 (N_9403,N_8243,N_8315);
nand U9404 (N_9404,N_8364,N_8513);
and U9405 (N_9405,N_8241,N_8896);
xnor U9406 (N_9406,N_8312,N_8771);
or U9407 (N_9407,N_8638,N_8663);
nor U9408 (N_9408,N_8044,N_8002);
xnor U9409 (N_9409,N_8691,N_8497);
and U9410 (N_9410,N_8857,N_8298);
nor U9411 (N_9411,N_8967,N_8501);
and U9412 (N_9412,N_8115,N_8633);
xor U9413 (N_9413,N_8302,N_8964);
xor U9414 (N_9414,N_8035,N_8484);
or U9415 (N_9415,N_8287,N_8578);
and U9416 (N_9416,N_8421,N_8563);
xor U9417 (N_9417,N_8836,N_8950);
and U9418 (N_9418,N_8316,N_8937);
xor U9419 (N_9419,N_8875,N_8555);
xor U9420 (N_9420,N_8292,N_8425);
nor U9421 (N_9421,N_8833,N_8380);
and U9422 (N_9422,N_8173,N_8919);
nand U9423 (N_9423,N_8966,N_8845);
and U9424 (N_9424,N_8159,N_8088);
or U9425 (N_9425,N_8366,N_8181);
xor U9426 (N_9426,N_8362,N_8894);
and U9427 (N_9427,N_8407,N_8993);
or U9428 (N_9428,N_8339,N_8694);
nand U9429 (N_9429,N_8134,N_8048);
xor U9430 (N_9430,N_8853,N_8872);
or U9431 (N_9431,N_8636,N_8905);
nor U9432 (N_9432,N_8630,N_8103);
xnor U9433 (N_9433,N_8549,N_8075);
or U9434 (N_9434,N_8678,N_8017);
nor U9435 (N_9435,N_8577,N_8125);
nand U9436 (N_9436,N_8953,N_8337);
nand U9437 (N_9437,N_8008,N_8797);
xor U9438 (N_9438,N_8245,N_8503);
nor U9439 (N_9439,N_8047,N_8688);
or U9440 (N_9440,N_8475,N_8431);
and U9441 (N_9441,N_8249,N_8500);
nand U9442 (N_9442,N_8530,N_8324);
xor U9443 (N_9443,N_8429,N_8635);
nand U9444 (N_9444,N_8698,N_8782);
xnor U9445 (N_9445,N_8194,N_8229);
nand U9446 (N_9446,N_8438,N_8682);
and U9447 (N_9447,N_8209,N_8237);
and U9448 (N_9448,N_8327,N_8175);
or U9449 (N_9449,N_8632,N_8516);
xnor U9450 (N_9450,N_8028,N_8594);
and U9451 (N_9451,N_8899,N_8900);
nor U9452 (N_9452,N_8922,N_8625);
or U9453 (N_9453,N_8411,N_8297);
nand U9454 (N_9454,N_8419,N_8665);
xor U9455 (N_9455,N_8884,N_8724);
or U9456 (N_9456,N_8648,N_8055);
nand U9457 (N_9457,N_8379,N_8696);
nor U9458 (N_9458,N_8511,N_8119);
nand U9459 (N_9459,N_8650,N_8128);
nor U9460 (N_9460,N_8155,N_8041);
xor U9461 (N_9461,N_8464,N_8653);
nand U9462 (N_9462,N_8016,N_8289);
xnor U9463 (N_9463,N_8821,N_8981);
nand U9464 (N_9464,N_8015,N_8690);
or U9465 (N_9465,N_8144,N_8876);
nand U9466 (N_9466,N_8897,N_8354);
nand U9467 (N_9467,N_8070,N_8059);
nand U9468 (N_9468,N_8107,N_8071);
nand U9469 (N_9469,N_8091,N_8588);
nor U9470 (N_9470,N_8179,N_8397);
xor U9471 (N_9471,N_8533,N_8785);
nand U9472 (N_9472,N_8335,N_8148);
or U9473 (N_9473,N_8449,N_8587);
or U9474 (N_9474,N_8994,N_8528);
or U9475 (N_9475,N_8681,N_8867);
or U9476 (N_9476,N_8498,N_8022);
xnor U9477 (N_9477,N_8856,N_8073);
nand U9478 (N_9478,N_8459,N_8067);
or U9479 (N_9479,N_8373,N_8439);
or U9480 (N_9480,N_8118,N_8831);
and U9481 (N_9481,N_8317,N_8145);
or U9482 (N_9482,N_8306,N_8760);
nor U9483 (N_9483,N_8196,N_8452);
and U9484 (N_9484,N_8776,N_8812);
and U9485 (N_9485,N_8300,N_8956);
nor U9486 (N_9486,N_8514,N_8476);
nor U9487 (N_9487,N_8260,N_8827);
or U9488 (N_9488,N_8437,N_8692);
xnor U9489 (N_9489,N_8078,N_8031);
and U9490 (N_9490,N_8211,N_8094);
nand U9491 (N_9491,N_8954,N_8848);
or U9492 (N_9492,N_8519,N_8718);
nor U9493 (N_9493,N_8072,N_8338);
and U9494 (N_9494,N_8582,N_8458);
nand U9495 (N_9495,N_8676,N_8832);
nor U9496 (N_9496,N_8190,N_8734);
or U9497 (N_9497,N_8046,N_8495);
xnor U9498 (N_9498,N_8968,N_8281);
or U9499 (N_9499,N_8036,N_8248);
nand U9500 (N_9500,N_8853,N_8432);
nand U9501 (N_9501,N_8890,N_8350);
and U9502 (N_9502,N_8839,N_8734);
and U9503 (N_9503,N_8122,N_8395);
xnor U9504 (N_9504,N_8424,N_8595);
nor U9505 (N_9505,N_8327,N_8325);
nor U9506 (N_9506,N_8520,N_8522);
xnor U9507 (N_9507,N_8406,N_8349);
nand U9508 (N_9508,N_8809,N_8636);
xor U9509 (N_9509,N_8413,N_8838);
xor U9510 (N_9510,N_8729,N_8458);
xor U9511 (N_9511,N_8972,N_8252);
or U9512 (N_9512,N_8468,N_8016);
nand U9513 (N_9513,N_8329,N_8493);
or U9514 (N_9514,N_8864,N_8293);
xnor U9515 (N_9515,N_8482,N_8683);
nor U9516 (N_9516,N_8487,N_8975);
or U9517 (N_9517,N_8696,N_8188);
and U9518 (N_9518,N_8745,N_8129);
nor U9519 (N_9519,N_8420,N_8387);
xor U9520 (N_9520,N_8330,N_8313);
nor U9521 (N_9521,N_8120,N_8421);
or U9522 (N_9522,N_8832,N_8085);
nor U9523 (N_9523,N_8616,N_8613);
and U9524 (N_9524,N_8571,N_8702);
nor U9525 (N_9525,N_8565,N_8316);
nand U9526 (N_9526,N_8505,N_8214);
xnor U9527 (N_9527,N_8742,N_8048);
or U9528 (N_9528,N_8612,N_8367);
nand U9529 (N_9529,N_8593,N_8258);
or U9530 (N_9530,N_8109,N_8138);
nand U9531 (N_9531,N_8168,N_8729);
nor U9532 (N_9532,N_8068,N_8846);
or U9533 (N_9533,N_8847,N_8859);
or U9534 (N_9534,N_8439,N_8877);
xor U9535 (N_9535,N_8322,N_8918);
nand U9536 (N_9536,N_8239,N_8643);
nand U9537 (N_9537,N_8153,N_8309);
and U9538 (N_9538,N_8721,N_8922);
xnor U9539 (N_9539,N_8158,N_8551);
nand U9540 (N_9540,N_8252,N_8992);
nand U9541 (N_9541,N_8240,N_8709);
nor U9542 (N_9542,N_8022,N_8137);
nor U9543 (N_9543,N_8635,N_8789);
nand U9544 (N_9544,N_8612,N_8932);
or U9545 (N_9545,N_8336,N_8685);
nand U9546 (N_9546,N_8189,N_8238);
and U9547 (N_9547,N_8810,N_8566);
xnor U9548 (N_9548,N_8307,N_8194);
nand U9549 (N_9549,N_8449,N_8817);
or U9550 (N_9550,N_8985,N_8214);
nor U9551 (N_9551,N_8167,N_8819);
or U9552 (N_9552,N_8972,N_8091);
nand U9553 (N_9553,N_8485,N_8884);
xor U9554 (N_9554,N_8285,N_8546);
nand U9555 (N_9555,N_8619,N_8720);
xor U9556 (N_9556,N_8075,N_8089);
xor U9557 (N_9557,N_8088,N_8781);
nor U9558 (N_9558,N_8014,N_8737);
nand U9559 (N_9559,N_8667,N_8317);
nand U9560 (N_9560,N_8724,N_8092);
and U9561 (N_9561,N_8473,N_8073);
nor U9562 (N_9562,N_8915,N_8608);
and U9563 (N_9563,N_8325,N_8270);
or U9564 (N_9564,N_8092,N_8233);
nor U9565 (N_9565,N_8206,N_8634);
nand U9566 (N_9566,N_8131,N_8887);
xor U9567 (N_9567,N_8046,N_8832);
nand U9568 (N_9568,N_8069,N_8032);
nand U9569 (N_9569,N_8849,N_8177);
xnor U9570 (N_9570,N_8114,N_8969);
and U9571 (N_9571,N_8430,N_8120);
xor U9572 (N_9572,N_8493,N_8649);
and U9573 (N_9573,N_8878,N_8827);
or U9574 (N_9574,N_8404,N_8285);
nand U9575 (N_9575,N_8778,N_8459);
or U9576 (N_9576,N_8081,N_8456);
xor U9577 (N_9577,N_8717,N_8355);
and U9578 (N_9578,N_8940,N_8220);
or U9579 (N_9579,N_8154,N_8845);
and U9580 (N_9580,N_8437,N_8803);
or U9581 (N_9581,N_8122,N_8984);
nor U9582 (N_9582,N_8473,N_8556);
xnor U9583 (N_9583,N_8826,N_8144);
xnor U9584 (N_9584,N_8174,N_8430);
and U9585 (N_9585,N_8973,N_8317);
xor U9586 (N_9586,N_8300,N_8057);
and U9587 (N_9587,N_8621,N_8169);
xor U9588 (N_9588,N_8777,N_8868);
nand U9589 (N_9589,N_8104,N_8307);
xor U9590 (N_9590,N_8689,N_8726);
xnor U9591 (N_9591,N_8141,N_8633);
or U9592 (N_9592,N_8382,N_8343);
xnor U9593 (N_9593,N_8583,N_8779);
or U9594 (N_9594,N_8100,N_8458);
nand U9595 (N_9595,N_8161,N_8433);
or U9596 (N_9596,N_8900,N_8759);
xor U9597 (N_9597,N_8692,N_8197);
and U9598 (N_9598,N_8779,N_8228);
and U9599 (N_9599,N_8055,N_8749);
or U9600 (N_9600,N_8667,N_8717);
nand U9601 (N_9601,N_8661,N_8957);
nor U9602 (N_9602,N_8876,N_8104);
nand U9603 (N_9603,N_8048,N_8204);
xor U9604 (N_9604,N_8144,N_8917);
or U9605 (N_9605,N_8179,N_8931);
and U9606 (N_9606,N_8772,N_8842);
nand U9607 (N_9607,N_8750,N_8214);
nand U9608 (N_9608,N_8984,N_8239);
xnor U9609 (N_9609,N_8510,N_8720);
and U9610 (N_9610,N_8448,N_8990);
and U9611 (N_9611,N_8986,N_8401);
nand U9612 (N_9612,N_8867,N_8679);
xnor U9613 (N_9613,N_8249,N_8636);
and U9614 (N_9614,N_8454,N_8370);
nand U9615 (N_9615,N_8209,N_8234);
nand U9616 (N_9616,N_8707,N_8290);
and U9617 (N_9617,N_8122,N_8901);
and U9618 (N_9618,N_8765,N_8345);
nor U9619 (N_9619,N_8696,N_8220);
nor U9620 (N_9620,N_8569,N_8774);
nand U9621 (N_9621,N_8721,N_8529);
or U9622 (N_9622,N_8533,N_8666);
and U9623 (N_9623,N_8492,N_8482);
nand U9624 (N_9624,N_8817,N_8034);
or U9625 (N_9625,N_8554,N_8464);
or U9626 (N_9626,N_8450,N_8078);
or U9627 (N_9627,N_8832,N_8040);
or U9628 (N_9628,N_8456,N_8629);
or U9629 (N_9629,N_8580,N_8733);
nand U9630 (N_9630,N_8264,N_8042);
nor U9631 (N_9631,N_8074,N_8388);
xnor U9632 (N_9632,N_8885,N_8235);
and U9633 (N_9633,N_8001,N_8664);
or U9634 (N_9634,N_8541,N_8784);
xnor U9635 (N_9635,N_8978,N_8179);
nor U9636 (N_9636,N_8283,N_8583);
nand U9637 (N_9637,N_8458,N_8599);
nor U9638 (N_9638,N_8373,N_8171);
or U9639 (N_9639,N_8394,N_8395);
nor U9640 (N_9640,N_8304,N_8426);
nor U9641 (N_9641,N_8547,N_8989);
or U9642 (N_9642,N_8419,N_8100);
and U9643 (N_9643,N_8119,N_8768);
xnor U9644 (N_9644,N_8978,N_8721);
and U9645 (N_9645,N_8985,N_8038);
xor U9646 (N_9646,N_8820,N_8753);
nor U9647 (N_9647,N_8869,N_8322);
or U9648 (N_9648,N_8856,N_8500);
nor U9649 (N_9649,N_8547,N_8940);
xor U9650 (N_9650,N_8627,N_8444);
xnor U9651 (N_9651,N_8206,N_8144);
nor U9652 (N_9652,N_8281,N_8137);
nand U9653 (N_9653,N_8403,N_8584);
or U9654 (N_9654,N_8278,N_8492);
xor U9655 (N_9655,N_8249,N_8259);
xor U9656 (N_9656,N_8762,N_8393);
or U9657 (N_9657,N_8907,N_8427);
nand U9658 (N_9658,N_8854,N_8726);
nor U9659 (N_9659,N_8691,N_8301);
or U9660 (N_9660,N_8411,N_8748);
and U9661 (N_9661,N_8329,N_8614);
nand U9662 (N_9662,N_8725,N_8214);
or U9663 (N_9663,N_8285,N_8540);
nor U9664 (N_9664,N_8453,N_8003);
nand U9665 (N_9665,N_8140,N_8711);
and U9666 (N_9666,N_8468,N_8819);
and U9667 (N_9667,N_8389,N_8381);
nand U9668 (N_9668,N_8154,N_8153);
or U9669 (N_9669,N_8192,N_8607);
and U9670 (N_9670,N_8773,N_8234);
nor U9671 (N_9671,N_8996,N_8130);
and U9672 (N_9672,N_8599,N_8890);
nor U9673 (N_9673,N_8620,N_8549);
nor U9674 (N_9674,N_8820,N_8407);
and U9675 (N_9675,N_8648,N_8970);
xnor U9676 (N_9676,N_8759,N_8396);
nor U9677 (N_9677,N_8125,N_8307);
xnor U9678 (N_9678,N_8751,N_8692);
or U9679 (N_9679,N_8146,N_8019);
or U9680 (N_9680,N_8990,N_8565);
and U9681 (N_9681,N_8529,N_8765);
nor U9682 (N_9682,N_8605,N_8904);
or U9683 (N_9683,N_8744,N_8369);
xnor U9684 (N_9684,N_8543,N_8486);
nand U9685 (N_9685,N_8082,N_8804);
xnor U9686 (N_9686,N_8504,N_8010);
or U9687 (N_9687,N_8558,N_8074);
nor U9688 (N_9688,N_8432,N_8475);
nand U9689 (N_9689,N_8595,N_8426);
or U9690 (N_9690,N_8276,N_8462);
nand U9691 (N_9691,N_8555,N_8202);
or U9692 (N_9692,N_8326,N_8177);
or U9693 (N_9693,N_8180,N_8224);
and U9694 (N_9694,N_8854,N_8989);
nor U9695 (N_9695,N_8310,N_8099);
and U9696 (N_9696,N_8632,N_8134);
nor U9697 (N_9697,N_8967,N_8948);
and U9698 (N_9698,N_8601,N_8005);
nor U9699 (N_9699,N_8373,N_8122);
nand U9700 (N_9700,N_8978,N_8375);
nand U9701 (N_9701,N_8823,N_8031);
xor U9702 (N_9702,N_8430,N_8589);
nand U9703 (N_9703,N_8131,N_8609);
nand U9704 (N_9704,N_8041,N_8671);
nor U9705 (N_9705,N_8532,N_8352);
nor U9706 (N_9706,N_8273,N_8322);
xor U9707 (N_9707,N_8003,N_8795);
nor U9708 (N_9708,N_8214,N_8247);
and U9709 (N_9709,N_8626,N_8091);
nand U9710 (N_9710,N_8124,N_8058);
and U9711 (N_9711,N_8729,N_8423);
nor U9712 (N_9712,N_8239,N_8927);
nand U9713 (N_9713,N_8829,N_8755);
or U9714 (N_9714,N_8568,N_8823);
or U9715 (N_9715,N_8156,N_8056);
nor U9716 (N_9716,N_8810,N_8179);
xor U9717 (N_9717,N_8681,N_8585);
nor U9718 (N_9718,N_8204,N_8608);
nand U9719 (N_9719,N_8766,N_8546);
nand U9720 (N_9720,N_8661,N_8518);
nand U9721 (N_9721,N_8448,N_8035);
xnor U9722 (N_9722,N_8891,N_8637);
or U9723 (N_9723,N_8019,N_8294);
xor U9724 (N_9724,N_8367,N_8170);
or U9725 (N_9725,N_8776,N_8272);
nor U9726 (N_9726,N_8287,N_8188);
or U9727 (N_9727,N_8164,N_8370);
nand U9728 (N_9728,N_8251,N_8061);
nand U9729 (N_9729,N_8832,N_8545);
xnor U9730 (N_9730,N_8997,N_8450);
or U9731 (N_9731,N_8722,N_8405);
or U9732 (N_9732,N_8415,N_8105);
xor U9733 (N_9733,N_8491,N_8876);
nand U9734 (N_9734,N_8373,N_8275);
and U9735 (N_9735,N_8495,N_8775);
or U9736 (N_9736,N_8153,N_8377);
or U9737 (N_9737,N_8803,N_8565);
or U9738 (N_9738,N_8211,N_8121);
and U9739 (N_9739,N_8604,N_8032);
xor U9740 (N_9740,N_8388,N_8379);
or U9741 (N_9741,N_8225,N_8126);
or U9742 (N_9742,N_8287,N_8581);
xor U9743 (N_9743,N_8335,N_8937);
or U9744 (N_9744,N_8767,N_8948);
or U9745 (N_9745,N_8755,N_8118);
and U9746 (N_9746,N_8003,N_8248);
or U9747 (N_9747,N_8965,N_8215);
xnor U9748 (N_9748,N_8994,N_8254);
xnor U9749 (N_9749,N_8300,N_8429);
nor U9750 (N_9750,N_8697,N_8488);
xor U9751 (N_9751,N_8599,N_8737);
nor U9752 (N_9752,N_8848,N_8183);
xor U9753 (N_9753,N_8971,N_8049);
xor U9754 (N_9754,N_8837,N_8794);
or U9755 (N_9755,N_8400,N_8692);
xor U9756 (N_9756,N_8389,N_8884);
and U9757 (N_9757,N_8417,N_8378);
or U9758 (N_9758,N_8662,N_8819);
or U9759 (N_9759,N_8909,N_8674);
or U9760 (N_9760,N_8539,N_8497);
and U9761 (N_9761,N_8540,N_8177);
or U9762 (N_9762,N_8210,N_8366);
nand U9763 (N_9763,N_8466,N_8993);
and U9764 (N_9764,N_8236,N_8542);
nand U9765 (N_9765,N_8119,N_8547);
xor U9766 (N_9766,N_8986,N_8531);
or U9767 (N_9767,N_8229,N_8496);
and U9768 (N_9768,N_8602,N_8941);
nand U9769 (N_9769,N_8755,N_8700);
or U9770 (N_9770,N_8343,N_8308);
nor U9771 (N_9771,N_8274,N_8108);
nand U9772 (N_9772,N_8911,N_8825);
or U9773 (N_9773,N_8243,N_8085);
nand U9774 (N_9774,N_8606,N_8891);
and U9775 (N_9775,N_8893,N_8895);
and U9776 (N_9776,N_8311,N_8324);
nand U9777 (N_9777,N_8506,N_8464);
or U9778 (N_9778,N_8981,N_8795);
and U9779 (N_9779,N_8147,N_8546);
xor U9780 (N_9780,N_8261,N_8620);
nand U9781 (N_9781,N_8282,N_8222);
or U9782 (N_9782,N_8793,N_8820);
and U9783 (N_9783,N_8761,N_8502);
or U9784 (N_9784,N_8605,N_8256);
and U9785 (N_9785,N_8941,N_8561);
or U9786 (N_9786,N_8395,N_8321);
or U9787 (N_9787,N_8190,N_8344);
and U9788 (N_9788,N_8059,N_8744);
nand U9789 (N_9789,N_8807,N_8591);
nand U9790 (N_9790,N_8539,N_8179);
nand U9791 (N_9791,N_8478,N_8284);
nand U9792 (N_9792,N_8579,N_8210);
xnor U9793 (N_9793,N_8589,N_8316);
xor U9794 (N_9794,N_8706,N_8492);
nand U9795 (N_9795,N_8460,N_8873);
nor U9796 (N_9796,N_8562,N_8407);
or U9797 (N_9797,N_8991,N_8501);
nand U9798 (N_9798,N_8040,N_8061);
nor U9799 (N_9799,N_8289,N_8778);
or U9800 (N_9800,N_8677,N_8700);
xor U9801 (N_9801,N_8593,N_8347);
or U9802 (N_9802,N_8850,N_8535);
nor U9803 (N_9803,N_8166,N_8373);
nand U9804 (N_9804,N_8335,N_8128);
nor U9805 (N_9805,N_8535,N_8469);
nor U9806 (N_9806,N_8269,N_8113);
or U9807 (N_9807,N_8065,N_8180);
and U9808 (N_9808,N_8656,N_8004);
or U9809 (N_9809,N_8143,N_8046);
nand U9810 (N_9810,N_8295,N_8810);
nand U9811 (N_9811,N_8753,N_8980);
nand U9812 (N_9812,N_8458,N_8736);
xor U9813 (N_9813,N_8976,N_8715);
nor U9814 (N_9814,N_8733,N_8951);
and U9815 (N_9815,N_8215,N_8685);
or U9816 (N_9816,N_8468,N_8337);
nand U9817 (N_9817,N_8087,N_8647);
or U9818 (N_9818,N_8307,N_8835);
nor U9819 (N_9819,N_8908,N_8774);
nand U9820 (N_9820,N_8470,N_8657);
or U9821 (N_9821,N_8647,N_8925);
xnor U9822 (N_9822,N_8369,N_8544);
xor U9823 (N_9823,N_8348,N_8262);
nand U9824 (N_9824,N_8929,N_8621);
nor U9825 (N_9825,N_8989,N_8324);
xnor U9826 (N_9826,N_8732,N_8419);
and U9827 (N_9827,N_8739,N_8172);
nand U9828 (N_9828,N_8932,N_8937);
xor U9829 (N_9829,N_8636,N_8492);
or U9830 (N_9830,N_8208,N_8813);
or U9831 (N_9831,N_8980,N_8711);
xnor U9832 (N_9832,N_8206,N_8006);
or U9833 (N_9833,N_8868,N_8042);
or U9834 (N_9834,N_8009,N_8877);
nand U9835 (N_9835,N_8442,N_8709);
nand U9836 (N_9836,N_8867,N_8336);
and U9837 (N_9837,N_8213,N_8057);
xor U9838 (N_9838,N_8260,N_8163);
nand U9839 (N_9839,N_8007,N_8240);
or U9840 (N_9840,N_8520,N_8921);
nor U9841 (N_9841,N_8617,N_8110);
nor U9842 (N_9842,N_8313,N_8915);
or U9843 (N_9843,N_8689,N_8161);
nor U9844 (N_9844,N_8403,N_8398);
nand U9845 (N_9845,N_8988,N_8737);
nand U9846 (N_9846,N_8852,N_8243);
nor U9847 (N_9847,N_8267,N_8576);
xnor U9848 (N_9848,N_8330,N_8245);
or U9849 (N_9849,N_8703,N_8902);
and U9850 (N_9850,N_8990,N_8554);
and U9851 (N_9851,N_8633,N_8061);
nor U9852 (N_9852,N_8059,N_8855);
xor U9853 (N_9853,N_8933,N_8497);
nand U9854 (N_9854,N_8072,N_8511);
and U9855 (N_9855,N_8059,N_8429);
nand U9856 (N_9856,N_8159,N_8150);
or U9857 (N_9857,N_8627,N_8517);
or U9858 (N_9858,N_8221,N_8441);
and U9859 (N_9859,N_8139,N_8096);
and U9860 (N_9860,N_8588,N_8836);
and U9861 (N_9861,N_8162,N_8151);
nor U9862 (N_9862,N_8283,N_8284);
nor U9863 (N_9863,N_8114,N_8010);
and U9864 (N_9864,N_8009,N_8961);
and U9865 (N_9865,N_8682,N_8566);
or U9866 (N_9866,N_8330,N_8018);
or U9867 (N_9867,N_8443,N_8889);
nor U9868 (N_9868,N_8451,N_8290);
xnor U9869 (N_9869,N_8930,N_8342);
and U9870 (N_9870,N_8146,N_8284);
xor U9871 (N_9871,N_8455,N_8218);
xnor U9872 (N_9872,N_8441,N_8092);
nand U9873 (N_9873,N_8061,N_8348);
xnor U9874 (N_9874,N_8359,N_8207);
nand U9875 (N_9875,N_8070,N_8164);
xnor U9876 (N_9876,N_8235,N_8576);
or U9877 (N_9877,N_8213,N_8619);
xor U9878 (N_9878,N_8662,N_8508);
nand U9879 (N_9879,N_8126,N_8310);
nand U9880 (N_9880,N_8285,N_8936);
nor U9881 (N_9881,N_8257,N_8464);
nor U9882 (N_9882,N_8500,N_8402);
xnor U9883 (N_9883,N_8602,N_8073);
and U9884 (N_9884,N_8002,N_8455);
or U9885 (N_9885,N_8112,N_8042);
nand U9886 (N_9886,N_8984,N_8745);
nor U9887 (N_9887,N_8299,N_8803);
or U9888 (N_9888,N_8976,N_8128);
xnor U9889 (N_9889,N_8102,N_8295);
xor U9890 (N_9890,N_8920,N_8454);
nand U9891 (N_9891,N_8589,N_8376);
xnor U9892 (N_9892,N_8734,N_8654);
xor U9893 (N_9893,N_8742,N_8177);
and U9894 (N_9894,N_8352,N_8540);
nand U9895 (N_9895,N_8711,N_8613);
and U9896 (N_9896,N_8326,N_8281);
nor U9897 (N_9897,N_8738,N_8113);
xor U9898 (N_9898,N_8542,N_8999);
or U9899 (N_9899,N_8721,N_8697);
or U9900 (N_9900,N_8002,N_8605);
nor U9901 (N_9901,N_8409,N_8546);
nand U9902 (N_9902,N_8472,N_8875);
xor U9903 (N_9903,N_8318,N_8747);
nor U9904 (N_9904,N_8167,N_8569);
nand U9905 (N_9905,N_8379,N_8132);
and U9906 (N_9906,N_8013,N_8798);
xor U9907 (N_9907,N_8094,N_8694);
xor U9908 (N_9908,N_8217,N_8210);
nor U9909 (N_9909,N_8852,N_8066);
nor U9910 (N_9910,N_8725,N_8275);
nand U9911 (N_9911,N_8078,N_8352);
xor U9912 (N_9912,N_8941,N_8884);
nand U9913 (N_9913,N_8654,N_8886);
nand U9914 (N_9914,N_8343,N_8100);
xnor U9915 (N_9915,N_8922,N_8143);
or U9916 (N_9916,N_8527,N_8623);
xnor U9917 (N_9917,N_8862,N_8989);
xor U9918 (N_9918,N_8789,N_8832);
nand U9919 (N_9919,N_8210,N_8361);
xor U9920 (N_9920,N_8193,N_8289);
nand U9921 (N_9921,N_8863,N_8248);
nor U9922 (N_9922,N_8798,N_8875);
xnor U9923 (N_9923,N_8490,N_8301);
and U9924 (N_9924,N_8412,N_8406);
or U9925 (N_9925,N_8641,N_8449);
and U9926 (N_9926,N_8501,N_8316);
or U9927 (N_9927,N_8333,N_8180);
nor U9928 (N_9928,N_8781,N_8572);
xnor U9929 (N_9929,N_8334,N_8958);
or U9930 (N_9930,N_8768,N_8323);
nand U9931 (N_9931,N_8902,N_8293);
or U9932 (N_9932,N_8970,N_8564);
xor U9933 (N_9933,N_8915,N_8436);
nor U9934 (N_9934,N_8534,N_8892);
nor U9935 (N_9935,N_8303,N_8561);
and U9936 (N_9936,N_8071,N_8789);
nor U9937 (N_9937,N_8864,N_8785);
and U9938 (N_9938,N_8484,N_8470);
or U9939 (N_9939,N_8221,N_8032);
xor U9940 (N_9940,N_8198,N_8927);
and U9941 (N_9941,N_8624,N_8473);
nand U9942 (N_9942,N_8412,N_8624);
nand U9943 (N_9943,N_8056,N_8458);
and U9944 (N_9944,N_8244,N_8206);
and U9945 (N_9945,N_8055,N_8392);
nor U9946 (N_9946,N_8198,N_8587);
nor U9947 (N_9947,N_8867,N_8776);
xor U9948 (N_9948,N_8519,N_8065);
xor U9949 (N_9949,N_8713,N_8491);
nand U9950 (N_9950,N_8218,N_8614);
and U9951 (N_9951,N_8610,N_8577);
and U9952 (N_9952,N_8501,N_8197);
xnor U9953 (N_9953,N_8479,N_8493);
xnor U9954 (N_9954,N_8485,N_8547);
xnor U9955 (N_9955,N_8670,N_8465);
nand U9956 (N_9956,N_8982,N_8683);
nor U9957 (N_9957,N_8804,N_8918);
xnor U9958 (N_9958,N_8315,N_8698);
nand U9959 (N_9959,N_8568,N_8049);
nor U9960 (N_9960,N_8316,N_8484);
nor U9961 (N_9961,N_8897,N_8724);
nand U9962 (N_9962,N_8359,N_8966);
xor U9963 (N_9963,N_8281,N_8841);
nor U9964 (N_9964,N_8893,N_8945);
nand U9965 (N_9965,N_8442,N_8724);
or U9966 (N_9966,N_8959,N_8619);
xor U9967 (N_9967,N_8816,N_8501);
xnor U9968 (N_9968,N_8588,N_8141);
or U9969 (N_9969,N_8618,N_8923);
nor U9970 (N_9970,N_8241,N_8783);
or U9971 (N_9971,N_8821,N_8947);
nand U9972 (N_9972,N_8200,N_8121);
or U9973 (N_9973,N_8609,N_8462);
nand U9974 (N_9974,N_8081,N_8362);
or U9975 (N_9975,N_8794,N_8579);
and U9976 (N_9976,N_8682,N_8106);
xnor U9977 (N_9977,N_8147,N_8176);
nand U9978 (N_9978,N_8399,N_8645);
or U9979 (N_9979,N_8287,N_8727);
nand U9980 (N_9980,N_8251,N_8659);
or U9981 (N_9981,N_8275,N_8037);
nor U9982 (N_9982,N_8621,N_8042);
and U9983 (N_9983,N_8518,N_8489);
xor U9984 (N_9984,N_8793,N_8235);
nand U9985 (N_9985,N_8358,N_8612);
or U9986 (N_9986,N_8842,N_8586);
and U9987 (N_9987,N_8089,N_8692);
xor U9988 (N_9988,N_8388,N_8915);
xor U9989 (N_9989,N_8541,N_8690);
xnor U9990 (N_9990,N_8324,N_8945);
xor U9991 (N_9991,N_8651,N_8400);
and U9992 (N_9992,N_8212,N_8069);
and U9993 (N_9993,N_8501,N_8080);
and U9994 (N_9994,N_8406,N_8897);
and U9995 (N_9995,N_8648,N_8290);
and U9996 (N_9996,N_8522,N_8555);
xnor U9997 (N_9997,N_8093,N_8078);
and U9998 (N_9998,N_8598,N_8327);
xor U9999 (N_9999,N_8726,N_8968);
or U10000 (N_10000,N_9330,N_9033);
or U10001 (N_10001,N_9374,N_9740);
nand U10002 (N_10002,N_9503,N_9287);
or U10003 (N_10003,N_9202,N_9825);
nor U10004 (N_10004,N_9274,N_9321);
nand U10005 (N_10005,N_9716,N_9613);
nor U10006 (N_10006,N_9098,N_9468);
and U10007 (N_10007,N_9393,N_9130);
and U10008 (N_10008,N_9451,N_9989);
nand U10009 (N_10009,N_9286,N_9601);
nor U10010 (N_10010,N_9345,N_9889);
nand U10011 (N_10011,N_9170,N_9789);
xnor U10012 (N_10012,N_9783,N_9419);
and U10013 (N_10013,N_9502,N_9172);
nand U10014 (N_10014,N_9077,N_9506);
nand U10015 (N_10015,N_9984,N_9223);
nand U10016 (N_10016,N_9311,N_9576);
or U10017 (N_10017,N_9416,N_9214);
and U10018 (N_10018,N_9895,N_9977);
nor U10019 (N_10019,N_9990,N_9869);
xor U10020 (N_10020,N_9937,N_9094);
nand U10021 (N_10021,N_9774,N_9204);
xnor U10022 (N_10022,N_9548,N_9616);
nor U10023 (N_10023,N_9779,N_9875);
or U10024 (N_10024,N_9743,N_9692);
nand U10025 (N_10025,N_9103,N_9925);
nor U10026 (N_10026,N_9087,N_9962);
and U10027 (N_10027,N_9864,N_9893);
and U10028 (N_10028,N_9426,N_9885);
nand U10029 (N_10029,N_9020,N_9310);
and U10030 (N_10030,N_9603,N_9195);
nor U10031 (N_10031,N_9487,N_9052);
xor U10032 (N_10032,N_9583,N_9014);
nand U10033 (N_10033,N_9557,N_9851);
or U10034 (N_10034,N_9032,N_9942);
nor U10035 (N_10035,N_9303,N_9436);
or U10036 (N_10036,N_9185,N_9654);
xor U10037 (N_10037,N_9134,N_9939);
nand U10038 (N_10038,N_9818,N_9376);
nand U10039 (N_10039,N_9600,N_9216);
or U10040 (N_10040,N_9674,N_9858);
nor U10041 (N_10041,N_9718,N_9882);
nand U10042 (N_10042,N_9703,N_9431);
and U10043 (N_10043,N_9000,N_9945);
nor U10044 (N_10044,N_9626,N_9715);
xnor U10045 (N_10045,N_9063,N_9235);
xor U10046 (N_10046,N_9517,N_9229);
and U10047 (N_10047,N_9272,N_9490);
or U10048 (N_10048,N_9566,N_9916);
and U10049 (N_10049,N_9335,N_9540);
and U10050 (N_10050,N_9403,N_9879);
nand U10051 (N_10051,N_9322,N_9242);
or U10052 (N_10052,N_9127,N_9960);
nand U10053 (N_10053,N_9846,N_9030);
and U10054 (N_10054,N_9791,N_9639);
and U10055 (N_10055,N_9293,N_9390);
and U10056 (N_10056,N_9731,N_9697);
xor U10057 (N_10057,N_9792,N_9051);
or U10058 (N_10058,N_9347,N_9594);
nand U10059 (N_10059,N_9057,N_9271);
nand U10060 (N_10060,N_9100,N_9702);
and U10061 (N_10061,N_9161,N_9258);
and U10062 (N_10062,N_9315,N_9480);
xor U10063 (N_10063,N_9435,N_9206);
or U10064 (N_10064,N_9773,N_9239);
xor U10065 (N_10065,N_9539,N_9927);
nand U10066 (N_10066,N_9580,N_9496);
or U10067 (N_10067,N_9084,N_9116);
and U10068 (N_10068,N_9061,N_9709);
nor U10069 (N_10069,N_9900,N_9831);
or U10070 (N_10070,N_9950,N_9920);
nand U10071 (N_10071,N_9289,N_9714);
nand U10072 (N_10072,N_9998,N_9447);
nor U10073 (N_10073,N_9081,N_9280);
xnor U10074 (N_10074,N_9821,N_9155);
and U10075 (N_10075,N_9649,N_9031);
xor U10076 (N_10076,N_9073,N_9633);
xor U10077 (N_10077,N_9296,N_9331);
or U10078 (N_10078,N_9406,N_9997);
nor U10079 (N_10079,N_9735,N_9001);
nand U10080 (N_10080,N_9290,N_9787);
and U10081 (N_10081,N_9295,N_9486);
or U10082 (N_10082,N_9737,N_9646);
nand U10083 (N_10083,N_9099,N_9949);
and U10084 (N_10084,N_9383,N_9838);
xnor U10085 (N_10085,N_9859,N_9364);
nor U10086 (N_10086,N_9154,N_9520);
nand U10087 (N_10087,N_9308,N_9993);
nor U10088 (N_10088,N_9189,N_9500);
nand U10089 (N_10089,N_9794,N_9260);
nand U10090 (N_10090,N_9277,N_9983);
xnor U10091 (N_10091,N_9568,N_9996);
or U10092 (N_10092,N_9698,N_9197);
or U10093 (N_10093,N_9750,N_9811);
and U10094 (N_10094,N_9733,N_9619);
xor U10095 (N_10095,N_9886,N_9809);
xnor U10096 (N_10096,N_9982,N_9294);
nand U10097 (N_10097,N_9726,N_9354);
nor U10098 (N_10098,N_9684,N_9163);
or U10099 (N_10099,N_9534,N_9346);
or U10100 (N_10100,N_9577,N_9527);
xor U10101 (N_10101,N_9333,N_9458);
nor U10102 (N_10102,N_9269,N_9704);
nand U10103 (N_10103,N_9824,N_9013);
and U10104 (N_10104,N_9002,N_9867);
nor U10105 (N_10105,N_9501,N_9117);
and U10106 (N_10106,N_9736,N_9054);
and U10107 (N_10107,N_9796,N_9834);
xnor U10108 (N_10108,N_9881,N_9037);
xnor U10109 (N_10109,N_9284,N_9123);
and U10110 (N_10110,N_9248,N_9378);
and U10111 (N_10111,N_9355,N_9379);
nand U10112 (N_10112,N_9399,N_9662);
or U10113 (N_10113,N_9911,N_9477);
or U10114 (N_10114,N_9976,N_9121);
xnor U10115 (N_10115,N_9327,N_9682);
xnor U10116 (N_10116,N_9251,N_9265);
xor U10117 (N_10117,N_9564,N_9083);
nand U10118 (N_10118,N_9917,N_9266);
or U10119 (N_10119,N_9660,N_9267);
or U10120 (N_10120,N_9168,N_9102);
nand U10121 (N_10121,N_9799,N_9012);
and U10122 (N_10122,N_9011,N_9781);
xor U10123 (N_10123,N_9659,N_9874);
or U10124 (N_10124,N_9391,N_9551);
nand U10125 (N_10125,N_9510,N_9689);
nand U10126 (N_10126,N_9201,N_9221);
nand U10127 (N_10127,N_9788,N_9860);
and U10128 (N_10128,N_9677,N_9456);
nor U10129 (N_10129,N_9086,N_9602);
and U10130 (N_10130,N_9699,N_9595);
xnor U10131 (N_10131,N_9428,N_9992);
nor U10132 (N_10132,N_9728,N_9048);
xor U10133 (N_10133,N_9617,N_9928);
nand U10134 (N_10134,N_9571,N_9805);
nand U10135 (N_10135,N_9592,N_9797);
and U10136 (N_10136,N_9299,N_9585);
nand U10137 (N_10137,N_9101,N_9957);
nor U10138 (N_10138,N_9301,N_9798);
or U10139 (N_10139,N_9375,N_9418);
and U10140 (N_10140,N_9777,N_9943);
and U10141 (N_10141,N_9400,N_9091);
nand U10142 (N_10142,N_9849,N_9681);
nor U10143 (N_10143,N_9902,N_9971);
nand U10144 (N_10144,N_9514,N_9146);
or U10145 (N_10145,N_9198,N_9363);
and U10146 (N_10146,N_9711,N_9505);
nand U10147 (N_10147,N_9870,N_9334);
nor U10148 (N_10148,N_9240,N_9298);
nand U10149 (N_10149,N_9723,N_9429);
and U10150 (N_10150,N_9285,N_9138);
or U10151 (N_10151,N_9524,N_9498);
or U10152 (N_10152,N_9856,N_9575);
or U10153 (N_10153,N_9464,N_9615);
nor U10154 (N_10154,N_9531,N_9782);
nand U10155 (N_10155,N_9912,N_9828);
nor U10156 (N_10156,N_9910,N_9466);
nand U10157 (N_10157,N_9222,N_9822);
xnor U10158 (N_10158,N_9397,N_9291);
nand U10159 (N_10159,N_9307,N_9224);
and U10160 (N_10160,N_9234,N_9455);
nand U10161 (N_10161,N_9956,N_9388);
xnor U10162 (N_10162,N_9452,N_9493);
xnor U10163 (N_10163,N_9437,N_9922);
nand U10164 (N_10164,N_9205,N_9663);
xor U10165 (N_10165,N_9629,N_9974);
or U10166 (N_10166,N_9096,N_9940);
nand U10167 (N_10167,N_9533,N_9283);
xnor U10168 (N_10168,N_9745,N_9358);
or U10169 (N_10169,N_9055,N_9572);
nor U10170 (N_10170,N_9817,N_9178);
nand U10171 (N_10171,N_9300,N_9761);
or U10172 (N_10172,N_9609,N_9730);
xnor U10173 (N_10173,N_9279,N_9395);
nor U10174 (N_10174,N_9582,N_9373);
xnor U10175 (N_10175,N_9385,N_9040);
or U10176 (N_10176,N_9316,N_9632);
nand U10177 (N_10177,N_9935,N_9407);
and U10178 (N_10178,N_9009,N_9541);
nor U10179 (N_10179,N_9739,N_9351);
nor U10180 (N_10180,N_9357,N_9752);
nor U10181 (N_10181,N_9836,N_9112);
xnor U10182 (N_10182,N_9144,N_9766);
xnor U10183 (N_10183,N_9412,N_9469);
nand U10184 (N_10184,N_9337,N_9156);
xor U10185 (N_10185,N_9901,N_9778);
nor U10186 (N_10186,N_9203,N_9166);
nand U10187 (N_10187,N_9471,N_9973);
and U10188 (N_10188,N_9732,N_9065);
nand U10189 (N_10189,N_9994,N_9010);
xor U10190 (N_10190,N_9965,N_9961);
and U10191 (N_10191,N_9196,N_9047);
or U10192 (N_10192,N_9705,N_9644);
and U10193 (N_10193,N_9710,N_9392);
nand U10194 (N_10194,N_9932,N_9213);
xor U10195 (N_10195,N_9350,N_9246);
nor U10196 (N_10196,N_9759,N_9394);
nand U10197 (N_10197,N_9765,N_9717);
nor U10198 (N_10198,N_9118,N_9210);
or U10199 (N_10199,N_9537,N_9133);
and U10200 (N_10200,N_9261,N_9685);
and U10201 (N_10201,N_9494,N_9148);
or U10202 (N_10202,N_9747,N_9670);
and U10203 (N_10203,N_9470,N_9948);
nand U10204 (N_10204,N_9866,N_9396);
xnor U10205 (N_10205,N_9512,N_9044);
and U10206 (N_10206,N_9323,N_9808);
or U10207 (N_10207,N_9402,N_9004);
and U10208 (N_10208,N_9946,N_9076);
xor U10209 (N_10209,N_9218,N_9529);
xor U10210 (N_10210,N_9446,N_9547);
nor U10211 (N_10211,N_9208,N_9245);
and U10212 (N_10212,N_9627,N_9693);
xnor U10213 (N_10213,N_9623,N_9596);
xnor U10214 (N_10214,N_9192,N_9230);
nor U10215 (N_10215,N_9405,N_9924);
or U10216 (N_10216,N_9905,N_9441);
nor U10217 (N_10217,N_9803,N_9748);
or U10218 (N_10218,N_9823,N_9495);
and U10219 (N_10219,N_9560,N_9854);
and U10220 (N_10220,N_9281,N_9970);
xor U10221 (N_10221,N_9309,N_9025);
nand U10222 (N_10222,N_9921,N_9381);
or U10223 (N_10223,N_9770,N_9833);
or U10224 (N_10224,N_9764,N_9482);
and U10225 (N_10225,N_9263,N_9814);
and U10226 (N_10226,N_9845,N_9069);
nor U10227 (N_10227,N_9071,N_9526);
or U10228 (N_10228,N_9590,N_9938);
or U10229 (N_10229,N_9741,N_9169);
nand U10230 (N_10230,N_9967,N_9078);
or U10231 (N_10231,N_9165,N_9827);
xor U10232 (N_10232,N_9656,N_9806);
nand U10233 (N_10233,N_9868,N_9411);
nand U10234 (N_10234,N_9636,N_9039);
xnor U10235 (N_10235,N_9558,N_9122);
and U10236 (N_10236,N_9349,N_9021);
nor U10237 (N_10237,N_9913,N_9164);
xnor U10238 (N_10238,N_9772,N_9143);
xor U10239 (N_10239,N_9963,N_9676);
nor U10240 (N_10240,N_9325,N_9367);
nand U10241 (N_10241,N_9304,N_9175);
or U10242 (N_10242,N_9080,N_9790);
or U10243 (N_10243,N_9622,N_9461);
xor U10244 (N_10244,N_9173,N_9604);
xnor U10245 (N_10245,N_9593,N_9135);
or U10246 (N_10246,N_9829,N_9929);
nand U10247 (N_10247,N_9588,N_9839);
or U10248 (N_10248,N_9516,N_9979);
and U10249 (N_10249,N_9729,N_9257);
nand U10250 (N_10250,N_9049,N_9694);
or U10251 (N_10251,N_9883,N_9926);
or U10252 (N_10252,N_9653,N_9137);
xor U10253 (N_10253,N_9085,N_9457);
nand U10254 (N_10254,N_9270,N_9092);
nor U10255 (N_10255,N_9687,N_9329);
or U10256 (N_10256,N_9158,N_9149);
and U10257 (N_10257,N_9578,N_9053);
or U10258 (N_10258,N_9819,N_9725);
nand U10259 (N_10259,N_9543,N_9319);
nor U10260 (N_10260,N_9093,N_9941);
xnor U10261 (N_10261,N_9262,N_9359);
nand U10262 (N_10262,N_9951,N_9584);
nor U10263 (N_10263,N_9986,N_9217);
nor U10264 (N_10264,N_9064,N_9273);
and U10265 (N_10265,N_9504,N_9415);
and U10266 (N_10266,N_9661,N_9022);
or U10267 (N_10267,N_9409,N_9306);
nor U10268 (N_10268,N_9150,N_9665);
or U10269 (N_10269,N_9988,N_9352);
and U10270 (N_10270,N_9252,N_9690);
nand U10271 (N_10271,N_9637,N_9519);
nand U10272 (N_10272,N_9876,N_9370);
or U10273 (N_10273,N_9862,N_9763);
or U10274 (N_10274,N_9795,N_9968);
nor U10275 (N_10275,N_9017,N_9389);
or U10276 (N_10276,N_9340,N_9066);
or U10277 (N_10277,N_9259,N_9691);
nor U10278 (N_10278,N_9947,N_9554);
nor U10279 (N_10279,N_9131,N_9522);
and U10280 (N_10280,N_9852,N_9671);
nand U10281 (N_10281,N_9847,N_9220);
or U10282 (N_10282,N_9414,N_9734);
or U10283 (N_10283,N_9755,N_9631);
or U10284 (N_10284,N_9784,N_9344);
or U10285 (N_10285,N_9673,N_9610);
or U10286 (N_10286,N_9362,N_9890);
nor U10287 (N_10287,N_9187,N_9499);
and U10288 (N_10288,N_9443,N_9128);
nor U10289 (N_10289,N_9918,N_9545);
and U10290 (N_10290,N_9145,N_9159);
and U10291 (N_10291,N_9966,N_9184);
nor U10292 (N_10292,N_9658,N_9621);
nor U10293 (N_10293,N_9802,N_9181);
nand U10294 (N_10294,N_9401,N_9445);
xor U10295 (N_10295,N_9591,N_9062);
nor U10296 (N_10296,N_9209,N_9785);
nor U10297 (N_10297,N_9059,N_9152);
and U10298 (N_10298,N_9721,N_9624);
nand U10299 (N_10299,N_9908,N_9183);
nand U10300 (N_10300,N_9141,N_9371);
nor U10301 (N_10301,N_9474,N_9872);
nand U10302 (N_10302,N_9276,N_9507);
or U10303 (N_10303,N_9018,N_9005);
or U10304 (N_10304,N_9919,N_9760);
or U10305 (N_10305,N_9147,N_9744);
nor U10306 (N_10306,N_9434,N_9573);
xnor U10307 (N_10307,N_9840,N_9342);
xor U10308 (N_10308,N_9598,N_9669);
or U10309 (N_10309,N_9645,N_9648);
or U10310 (N_10310,N_9372,N_9413);
or U10311 (N_10311,N_9638,N_9425);
nor U10312 (N_10312,N_9873,N_9140);
nand U10313 (N_10313,N_9706,N_9219);
and U10314 (N_10314,N_9453,N_9328);
or U10315 (N_10315,N_9029,N_9114);
and U10316 (N_10316,N_9933,N_9643);
nor U10317 (N_10317,N_9008,N_9683);
nor U10318 (N_10318,N_9800,N_9614);
and U10319 (N_10319,N_9769,N_9124);
nor U10320 (N_10320,N_9028,N_9511);
nand U10321 (N_10321,N_9440,N_9314);
xor U10322 (N_10322,N_9199,N_9625);
xor U10323 (N_10323,N_9892,N_9475);
and U10324 (N_10324,N_9556,N_9775);
or U10325 (N_10325,N_9459,N_9757);
and U10326 (N_10326,N_9820,N_9243);
nand U10327 (N_10327,N_9142,N_9043);
nand U10328 (N_10328,N_9404,N_9254);
xor U10329 (N_10329,N_9844,N_9410);
nand U10330 (N_10330,N_9871,N_9433);
nand U10331 (N_10331,N_9944,N_9587);
and U10332 (N_10332,N_9275,N_9233);
xnor U10333 (N_10333,N_9589,N_9225);
nand U10334 (N_10334,N_9980,N_9807);
nor U10335 (N_10335,N_9958,N_9953);
nor U10336 (N_10336,N_9125,N_9421);
or U10337 (N_10337,N_9481,N_9338);
xnor U10338 (N_10338,N_9640,N_9518);
nor U10339 (N_10339,N_9422,N_9136);
and U10340 (N_10340,N_9250,N_9525);
nor U10341 (N_10341,N_9036,N_9999);
xor U10342 (N_10342,N_9108,N_9975);
xor U10343 (N_10343,N_9454,N_9832);
xor U10344 (N_10344,N_9896,N_9768);
or U10345 (N_10345,N_9708,N_9720);
nor U10346 (N_10346,N_9353,N_9180);
nand U10347 (N_10347,N_9664,N_9110);
nand U10348 (N_10348,N_9082,N_9343);
and U10349 (N_10349,N_9462,N_9023);
or U10350 (N_10350,N_9176,N_9696);
nor U10351 (N_10351,N_9978,N_9835);
or U10352 (N_10352,N_9969,N_9200);
and U10353 (N_10353,N_9369,N_9536);
xor U10354 (N_10354,N_9278,N_9312);
nor U10355 (N_10355,N_9302,N_9105);
nor U10356 (N_10356,N_9894,N_9758);
xnor U10357 (N_10357,N_9226,N_9955);
nor U10358 (N_10358,N_9460,N_9567);
nand U10359 (N_10359,N_9542,N_9837);
or U10360 (N_10360,N_9597,N_9855);
and U10361 (N_10361,N_9088,N_9909);
nand U10362 (N_10362,N_9417,N_9478);
nand U10363 (N_10363,N_9003,N_9630);
and U10364 (N_10364,N_9007,N_9041);
nand U10365 (N_10365,N_9552,N_9045);
or U10366 (N_10366,N_9863,N_9570);
or U10367 (N_10367,N_9360,N_9247);
xnor U10368 (N_10368,N_9672,N_9467);
nor U10369 (N_10369,N_9700,N_9793);
nand U10370 (N_10370,N_9508,N_9813);
xnor U10371 (N_10371,N_9387,N_9581);
or U10372 (N_10372,N_9463,N_9380);
nand U10373 (N_10373,N_9857,N_9238);
xnor U10374 (N_10374,N_9804,N_9695);
nand U10375 (N_10375,N_9268,N_9565);
xor U10376 (N_10376,N_9104,N_9034);
nand U10377 (N_10377,N_9954,N_9878);
nor U10378 (N_10378,N_9897,N_9236);
nand U10379 (N_10379,N_9182,N_9132);
nand U10380 (N_10380,N_9751,N_9384);
or U10381 (N_10381,N_9153,N_9438);
xnor U10382 (N_10382,N_9848,N_9042);
xor U10383 (N_10383,N_9292,N_9550);
and U10384 (N_10384,N_9377,N_9074);
and U10385 (N_10385,N_9256,N_9923);
and U10386 (N_10386,N_9366,N_9607);
xnor U10387 (N_10387,N_9528,N_9212);
or U10388 (N_10388,N_9906,N_9079);
and U10389 (N_10389,N_9056,N_9476);
xor U10390 (N_10390,N_9424,N_9167);
and U10391 (N_10391,N_9015,N_9336);
and U10392 (N_10392,N_9249,N_9742);
or U10393 (N_10393,N_9877,N_9339);
nand U10394 (N_10394,N_9810,N_9126);
nand U10395 (N_10395,N_9050,N_9553);
nor U10396 (N_10396,N_9865,N_9521);
nor U10397 (N_10397,N_9194,N_9650);
nor U10398 (N_10398,N_9207,N_9667);
or U10399 (N_10399,N_9569,N_9151);
nand U10400 (N_10400,N_9341,N_9563);
nand U10401 (N_10401,N_9241,N_9738);
xnor U10402 (N_10402,N_9675,N_9850);
nand U10403 (N_10403,N_9599,N_9722);
or U10404 (N_10404,N_9106,N_9090);
xnor U10405 (N_10405,N_9068,N_9904);
and U10406 (N_10406,N_9801,N_9861);
nand U10407 (N_10407,N_9472,N_9324);
nor U10408 (N_10408,N_9513,N_9450);
nor U10409 (N_10409,N_9887,N_9915);
nor U10410 (N_10410,N_9964,N_9157);
xnor U10411 (N_10411,N_9561,N_9776);
nand U10412 (N_10412,N_9215,N_9952);
xor U10413 (N_10413,N_9492,N_9489);
or U10414 (N_10414,N_9688,N_9186);
xnor U10415 (N_10415,N_9538,N_9509);
xnor U10416 (N_10416,N_9841,N_9707);
or U10417 (N_10417,N_9326,N_9264);
or U10418 (N_10418,N_9420,N_9237);
or U10419 (N_10419,N_9686,N_9075);
xnor U10420 (N_10420,N_9934,N_9635);
or U10421 (N_10421,N_9060,N_9227);
nor U10422 (N_10422,N_9432,N_9067);
and U10423 (N_10423,N_9113,N_9724);
nor U10424 (N_10424,N_9408,N_9668);
and U10425 (N_10425,N_9016,N_9070);
nor U10426 (N_10426,N_9448,N_9898);
and U10427 (N_10427,N_9095,N_9812);
nand U10428 (N_10428,N_9006,N_9891);
xor U10429 (N_10429,N_9749,N_9657);
nor U10430 (N_10430,N_9771,N_9193);
or U10431 (N_10431,N_9853,N_9120);
nor U10432 (N_10432,N_9427,N_9930);
nand U10433 (N_10433,N_9985,N_9719);
or U10434 (N_10434,N_9318,N_9046);
and U10435 (N_10435,N_9666,N_9244);
nor U10436 (N_10436,N_9365,N_9097);
nor U10437 (N_10437,N_9972,N_9815);
or U10438 (N_10438,N_9439,N_9914);
nor U10439 (N_10439,N_9305,N_9109);
xor U10440 (N_10440,N_9713,N_9611);
nand U10441 (N_10441,N_9449,N_9931);
xnor U10442 (N_10442,N_9907,N_9652);
nor U10443 (N_10443,N_9382,N_9680);
or U10444 (N_10444,N_9058,N_9356);
nand U10445 (N_10445,N_9191,N_9701);
or U10446 (N_10446,N_9641,N_9995);
xnor U10447 (N_10447,N_9991,N_9562);
nor U10448 (N_10448,N_9473,N_9546);
nand U10449 (N_10449,N_9903,N_9727);
nand U10450 (N_10450,N_9488,N_9620);
nor U10451 (N_10451,N_9959,N_9177);
nor U10452 (N_10452,N_9026,N_9628);
nand U10453 (N_10453,N_9753,N_9139);
xnor U10454 (N_10454,N_9842,N_9317);
xor U10455 (N_10455,N_9574,N_9038);
nor U10456 (N_10456,N_9089,N_9348);
and U10457 (N_10457,N_9880,N_9712);
nor U10458 (N_10458,N_9549,N_9888);
xnor U10459 (N_10459,N_9444,N_9987);
nor U10460 (N_10460,N_9282,N_9612);
xor U10461 (N_10461,N_9232,N_9211);
or U10462 (N_10462,N_9497,N_9479);
nand U10463 (N_10463,N_9129,N_9190);
nor U10464 (N_10464,N_9756,N_9188);
and U10465 (N_10465,N_9936,N_9430);
nand U10466 (N_10466,N_9027,N_9555);
and U10467 (N_10467,N_9465,N_9608);
or U10468 (N_10468,N_9484,N_9160);
or U10469 (N_10469,N_9171,N_9762);
nor U10470 (N_10470,N_9162,N_9024);
nor U10471 (N_10471,N_9634,N_9754);
nor U10472 (N_10472,N_9830,N_9179);
nand U10473 (N_10473,N_9884,N_9386);
nor U10474 (N_10474,N_9780,N_9523);
or U10475 (N_10475,N_9231,N_9532);
nor U10476 (N_10476,N_9679,N_9361);
nand U10477 (N_10477,N_9255,N_9544);
and U10478 (N_10478,N_9228,N_9642);
nor U10479 (N_10479,N_9368,N_9606);
or U10480 (N_10480,N_9320,N_9119);
xor U10481 (N_10481,N_9288,N_9826);
nand U10482 (N_10482,N_9035,N_9332);
xnor U10483 (N_10483,N_9655,N_9786);
and U10484 (N_10484,N_9647,N_9746);
and U10485 (N_10485,N_9586,N_9174);
nor U10486 (N_10486,N_9530,N_9535);
xor U10487 (N_10487,N_9618,N_9559);
nand U10488 (N_10488,N_9485,N_9297);
and U10489 (N_10489,N_9491,N_9651);
xor U10490 (N_10490,N_9981,N_9816);
and U10491 (N_10491,N_9579,N_9423);
xor U10492 (N_10492,N_9253,N_9072);
and U10493 (N_10493,N_9605,N_9678);
and U10494 (N_10494,N_9019,N_9843);
nand U10495 (N_10495,N_9515,N_9115);
and U10496 (N_10496,N_9107,N_9442);
and U10497 (N_10497,N_9483,N_9899);
xor U10498 (N_10498,N_9111,N_9313);
and U10499 (N_10499,N_9767,N_9398);
xnor U10500 (N_10500,N_9762,N_9395);
nand U10501 (N_10501,N_9689,N_9174);
nor U10502 (N_10502,N_9115,N_9128);
xor U10503 (N_10503,N_9914,N_9453);
xnor U10504 (N_10504,N_9176,N_9591);
and U10505 (N_10505,N_9304,N_9408);
nand U10506 (N_10506,N_9578,N_9288);
xnor U10507 (N_10507,N_9551,N_9441);
nor U10508 (N_10508,N_9880,N_9647);
nor U10509 (N_10509,N_9665,N_9613);
nand U10510 (N_10510,N_9368,N_9854);
nand U10511 (N_10511,N_9752,N_9943);
nand U10512 (N_10512,N_9510,N_9112);
nor U10513 (N_10513,N_9988,N_9161);
or U10514 (N_10514,N_9065,N_9315);
and U10515 (N_10515,N_9166,N_9254);
xor U10516 (N_10516,N_9137,N_9777);
xnor U10517 (N_10517,N_9015,N_9840);
nor U10518 (N_10518,N_9930,N_9966);
and U10519 (N_10519,N_9581,N_9018);
xnor U10520 (N_10520,N_9433,N_9282);
nor U10521 (N_10521,N_9424,N_9292);
and U10522 (N_10522,N_9635,N_9776);
or U10523 (N_10523,N_9448,N_9334);
or U10524 (N_10524,N_9941,N_9108);
or U10525 (N_10525,N_9050,N_9700);
nand U10526 (N_10526,N_9938,N_9734);
nor U10527 (N_10527,N_9077,N_9364);
xnor U10528 (N_10528,N_9196,N_9838);
xnor U10529 (N_10529,N_9145,N_9820);
or U10530 (N_10530,N_9929,N_9978);
and U10531 (N_10531,N_9551,N_9679);
or U10532 (N_10532,N_9745,N_9923);
xor U10533 (N_10533,N_9228,N_9745);
nand U10534 (N_10534,N_9188,N_9750);
nor U10535 (N_10535,N_9845,N_9877);
or U10536 (N_10536,N_9119,N_9104);
xnor U10537 (N_10537,N_9109,N_9215);
and U10538 (N_10538,N_9588,N_9411);
nand U10539 (N_10539,N_9868,N_9634);
xnor U10540 (N_10540,N_9667,N_9709);
nor U10541 (N_10541,N_9964,N_9884);
nor U10542 (N_10542,N_9787,N_9436);
xnor U10543 (N_10543,N_9300,N_9924);
xnor U10544 (N_10544,N_9276,N_9014);
nor U10545 (N_10545,N_9302,N_9692);
nand U10546 (N_10546,N_9666,N_9073);
nand U10547 (N_10547,N_9064,N_9668);
and U10548 (N_10548,N_9624,N_9778);
and U10549 (N_10549,N_9023,N_9610);
nor U10550 (N_10550,N_9304,N_9212);
and U10551 (N_10551,N_9206,N_9070);
and U10552 (N_10552,N_9105,N_9166);
nor U10553 (N_10553,N_9378,N_9616);
nand U10554 (N_10554,N_9563,N_9022);
nor U10555 (N_10555,N_9782,N_9788);
nand U10556 (N_10556,N_9417,N_9725);
nor U10557 (N_10557,N_9086,N_9440);
nand U10558 (N_10558,N_9310,N_9012);
or U10559 (N_10559,N_9319,N_9976);
and U10560 (N_10560,N_9900,N_9913);
xnor U10561 (N_10561,N_9540,N_9791);
xor U10562 (N_10562,N_9551,N_9125);
or U10563 (N_10563,N_9460,N_9719);
xor U10564 (N_10564,N_9322,N_9712);
or U10565 (N_10565,N_9287,N_9190);
or U10566 (N_10566,N_9403,N_9616);
nand U10567 (N_10567,N_9168,N_9452);
and U10568 (N_10568,N_9990,N_9277);
xnor U10569 (N_10569,N_9361,N_9162);
or U10570 (N_10570,N_9459,N_9342);
or U10571 (N_10571,N_9186,N_9184);
and U10572 (N_10572,N_9272,N_9796);
nor U10573 (N_10573,N_9175,N_9171);
xnor U10574 (N_10574,N_9831,N_9470);
and U10575 (N_10575,N_9852,N_9876);
or U10576 (N_10576,N_9088,N_9578);
nor U10577 (N_10577,N_9883,N_9905);
or U10578 (N_10578,N_9926,N_9528);
nand U10579 (N_10579,N_9985,N_9898);
or U10580 (N_10580,N_9047,N_9058);
nand U10581 (N_10581,N_9222,N_9078);
or U10582 (N_10582,N_9727,N_9324);
and U10583 (N_10583,N_9526,N_9767);
and U10584 (N_10584,N_9051,N_9048);
nand U10585 (N_10585,N_9338,N_9907);
xor U10586 (N_10586,N_9336,N_9120);
and U10587 (N_10587,N_9103,N_9072);
xnor U10588 (N_10588,N_9530,N_9531);
nor U10589 (N_10589,N_9637,N_9063);
xnor U10590 (N_10590,N_9060,N_9787);
nor U10591 (N_10591,N_9716,N_9904);
nor U10592 (N_10592,N_9722,N_9032);
or U10593 (N_10593,N_9400,N_9336);
xnor U10594 (N_10594,N_9633,N_9369);
xnor U10595 (N_10595,N_9686,N_9019);
nor U10596 (N_10596,N_9098,N_9606);
and U10597 (N_10597,N_9791,N_9278);
or U10598 (N_10598,N_9816,N_9737);
nand U10599 (N_10599,N_9612,N_9954);
nand U10600 (N_10600,N_9285,N_9185);
xor U10601 (N_10601,N_9631,N_9453);
nand U10602 (N_10602,N_9935,N_9567);
xnor U10603 (N_10603,N_9753,N_9990);
nand U10604 (N_10604,N_9780,N_9917);
nor U10605 (N_10605,N_9857,N_9551);
nor U10606 (N_10606,N_9724,N_9042);
xnor U10607 (N_10607,N_9796,N_9006);
nor U10608 (N_10608,N_9212,N_9800);
nand U10609 (N_10609,N_9989,N_9188);
nor U10610 (N_10610,N_9091,N_9476);
and U10611 (N_10611,N_9451,N_9377);
xnor U10612 (N_10612,N_9689,N_9816);
nor U10613 (N_10613,N_9415,N_9051);
xnor U10614 (N_10614,N_9273,N_9458);
or U10615 (N_10615,N_9388,N_9818);
xnor U10616 (N_10616,N_9725,N_9557);
nand U10617 (N_10617,N_9651,N_9815);
nor U10618 (N_10618,N_9119,N_9508);
or U10619 (N_10619,N_9851,N_9099);
nor U10620 (N_10620,N_9033,N_9025);
nor U10621 (N_10621,N_9145,N_9974);
nand U10622 (N_10622,N_9478,N_9962);
nand U10623 (N_10623,N_9041,N_9426);
xor U10624 (N_10624,N_9857,N_9547);
or U10625 (N_10625,N_9314,N_9392);
xor U10626 (N_10626,N_9413,N_9074);
nand U10627 (N_10627,N_9825,N_9237);
or U10628 (N_10628,N_9917,N_9341);
xnor U10629 (N_10629,N_9063,N_9761);
nand U10630 (N_10630,N_9256,N_9445);
nor U10631 (N_10631,N_9222,N_9215);
nand U10632 (N_10632,N_9173,N_9191);
xnor U10633 (N_10633,N_9217,N_9706);
xnor U10634 (N_10634,N_9494,N_9588);
xnor U10635 (N_10635,N_9341,N_9863);
and U10636 (N_10636,N_9614,N_9887);
xor U10637 (N_10637,N_9959,N_9794);
nor U10638 (N_10638,N_9355,N_9086);
nand U10639 (N_10639,N_9844,N_9689);
or U10640 (N_10640,N_9953,N_9780);
nor U10641 (N_10641,N_9174,N_9714);
and U10642 (N_10642,N_9219,N_9138);
xnor U10643 (N_10643,N_9647,N_9734);
nand U10644 (N_10644,N_9289,N_9444);
or U10645 (N_10645,N_9285,N_9940);
and U10646 (N_10646,N_9339,N_9041);
nor U10647 (N_10647,N_9789,N_9592);
or U10648 (N_10648,N_9074,N_9627);
nand U10649 (N_10649,N_9285,N_9496);
xnor U10650 (N_10650,N_9149,N_9343);
nor U10651 (N_10651,N_9534,N_9880);
nor U10652 (N_10652,N_9551,N_9572);
xnor U10653 (N_10653,N_9249,N_9507);
or U10654 (N_10654,N_9334,N_9342);
xnor U10655 (N_10655,N_9019,N_9928);
xnor U10656 (N_10656,N_9288,N_9337);
nand U10657 (N_10657,N_9269,N_9215);
nor U10658 (N_10658,N_9202,N_9834);
and U10659 (N_10659,N_9295,N_9327);
and U10660 (N_10660,N_9544,N_9490);
nor U10661 (N_10661,N_9893,N_9668);
and U10662 (N_10662,N_9534,N_9046);
xnor U10663 (N_10663,N_9554,N_9534);
nand U10664 (N_10664,N_9653,N_9489);
xor U10665 (N_10665,N_9588,N_9340);
or U10666 (N_10666,N_9298,N_9345);
or U10667 (N_10667,N_9714,N_9871);
xor U10668 (N_10668,N_9035,N_9642);
xnor U10669 (N_10669,N_9533,N_9346);
and U10670 (N_10670,N_9446,N_9831);
nand U10671 (N_10671,N_9309,N_9753);
xor U10672 (N_10672,N_9597,N_9294);
nand U10673 (N_10673,N_9668,N_9935);
or U10674 (N_10674,N_9521,N_9860);
xor U10675 (N_10675,N_9542,N_9021);
nand U10676 (N_10676,N_9332,N_9935);
nor U10677 (N_10677,N_9512,N_9970);
nand U10678 (N_10678,N_9247,N_9073);
xor U10679 (N_10679,N_9663,N_9954);
and U10680 (N_10680,N_9238,N_9251);
and U10681 (N_10681,N_9395,N_9258);
nand U10682 (N_10682,N_9475,N_9220);
nand U10683 (N_10683,N_9572,N_9915);
xnor U10684 (N_10684,N_9206,N_9604);
or U10685 (N_10685,N_9320,N_9673);
nor U10686 (N_10686,N_9523,N_9677);
xnor U10687 (N_10687,N_9624,N_9452);
and U10688 (N_10688,N_9393,N_9114);
and U10689 (N_10689,N_9072,N_9165);
or U10690 (N_10690,N_9593,N_9889);
or U10691 (N_10691,N_9342,N_9035);
nor U10692 (N_10692,N_9669,N_9890);
xor U10693 (N_10693,N_9973,N_9358);
and U10694 (N_10694,N_9862,N_9896);
and U10695 (N_10695,N_9313,N_9633);
or U10696 (N_10696,N_9883,N_9107);
nand U10697 (N_10697,N_9272,N_9540);
or U10698 (N_10698,N_9629,N_9706);
nor U10699 (N_10699,N_9443,N_9985);
nand U10700 (N_10700,N_9329,N_9673);
xor U10701 (N_10701,N_9131,N_9833);
or U10702 (N_10702,N_9815,N_9365);
xnor U10703 (N_10703,N_9535,N_9203);
and U10704 (N_10704,N_9855,N_9652);
xor U10705 (N_10705,N_9406,N_9148);
nor U10706 (N_10706,N_9504,N_9279);
or U10707 (N_10707,N_9261,N_9208);
nor U10708 (N_10708,N_9188,N_9924);
and U10709 (N_10709,N_9543,N_9391);
nand U10710 (N_10710,N_9743,N_9601);
or U10711 (N_10711,N_9844,N_9206);
and U10712 (N_10712,N_9425,N_9742);
xor U10713 (N_10713,N_9766,N_9390);
nor U10714 (N_10714,N_9826,N_9778);
and U10715 (N_10715,N_9870,N_9526);
nor U10716 (N_10716,N_9611,N_9762);
nor U10717 (N_10717,N_9958,N_9853);
xnor U10718 (N_10718,N_9182,N_9288);
and U10719 (N_10719,N_9440,N_9753);
and U10720 (N_10720,N_9445,N_9366);
nor U10721 (N_10721,N_9805,N_9973);
xor U10722 (N_10722,N_9122,N_9795);
or U10723 (N_10723,N_9957,N_9802);
nor U10724 (N_10724,N_9501,N_9637);
nor U10725 (N_10725,N_9747,N_9136);
nand U10726 (N_10726,N_9259,N_9936);
nand U10727 (N_10727,N_9641,N_9273);
nand U10728 (N_10728,N_9017,N_9530);
and U10729 (N_10729,N_9594,N_9820);
nor U10730 (N_10730,N_9373,N_9794);
or U10731 (N_10731,N_9392,N_9957);
and U10732 (N_10732,N_9589,N_9442);
nand U10733 (N_10733,N_9185,N_9670);
nor U10734 (N_10734,N_9125,N_9567);
nand U10735 (N_10735,N_9110,N_9007);
or U10736 (N_10736,N_9493,N_9353);
nand U10737 (N_10737,N_9142,N_9439);
or U10738 (N_10738,N_9743,N_9848);
xnor U10739 (N_10739,N_9866,N_9780);
xor U10740 (N_10740,N_9047,N_9020);
nand U10741 (N_10741,N_9633,N_9154);
and U10742 (N_10742,N_9052,N_9870);
nand U10743 (N_10743,N_9098,N_9908);
or U10744 (N_10744,N_9913,N_9651);
and U10745 (N_10745,N_9004,N_9629);
and U10746 (N_10746,N_9213,N_9138);
and U10747 (N_10747,N_9187,N_9521);
xor U10748 (N_10748,N_9801,N_9356);
nand U10749 (N_10749,N_9160,N_9022);
and U10750 (N_10750,N_9517,N_9664);
and U10751 (N_10751,N_9164,N_9858);
or U10752 (N_10752,N_9628,N_9736);
or U10753 (N_10753,N_9133,N_9799);
xor U10754 (N_10754,N_9353,N_9460);
xnor U10755 (N_10755,N_9049,N_9586);
or U10756 (N_10756,N_9972,N_9491);
or U10757 (N_10757,N_9768,N_9462);
or U10758 (N_10758,N_9621,N_9189);
xor U10759 (N_10759,N_9563,N_9079);
and U10760 (N_10760,N_9265,N_9413);
xor U10761 (N_10761,N_9297,N_9798);
nor U10762 (N_10762,N_9239,N_9081);
or U10763 (N_10763,N_9845,N_9190);
xor U10764 (N_10764,N_9665,N_9396);
and U10765 (N_10765,N_9469,N_9076);
nand U10766 (N_10766,N_9308,N_9018);
or U10767 (N_10767,N_9750,N_9329);
nor U10768 (N_10768,N_9176,N_9785);
nand U10769 (N_10769,N_9776,N_9532);
xor U10770 (N_10770,N_9260,N_9201);
and U10771 (N_10771,N_9079,N_9914);
or U10772 (N_10772,N_9447,N_9747);
nand U10773 (N_10773,N_9966,N_9546);
or U10774 (N_10774,N_9142,N_9375);
and U10775 (N_10775,N_9057,N_9597);
nand U10776 (N_10776,N_9389,N_9089);
nor U10777 (N_10777,N_9542,N_9087);
and U10778 (N_10778,N_9049,N_9505);
xor U10779 (N_10779,N_9174,N_9353);
xor U10780 (N_10780,N_9886,N_9556);
nor U10781 (N_10781,N_9877,N_9886);
xor U10782 (N_10782,N_9432,N_9264);
nor U10783 (N_10783,N_9727,N_9724);
and U10784 (N_10784,N_9753,N_9046);
xnor U10785 (N_10785,N_9655,N_9177);
or U10786 (N_10786,N_9366,N_9746);
nand U10787 (N_10787,N_9967,N_9226);
nand U10788 (N_10788,N_9684,N_9460);
nor U10789 (N_10789,N_9832,N_9873);
nor U10790 (N_10790,N_9647,N_9840);
and U10791 (N_10791,N_9438,N_9878);
xor U10792 (N_10792,N_9904,N_9793);
xor U10793 (N_10793,N_9024,N_9479);
nor U10794 (N_10794,N_9829,N_9973);
or U10795 (N_10795,N_9436,N_9843);
or U10796 (N_10796,N_9657,N_9138);
nor U10797 (N_10797,N_9084,N_9615);
or U10798 (N_10798,N_9461,N_9762);
nor U10799 (N_10799,N_9433,N_9654);
nor U10800 (N_10800,N_9053,N_9627);
xnor U10801 (N_10801,N_9045,N_9217);
nor U10802 (N_10802,N_9330,N_9504);
xnor U10803 (N_10803,N_9670,N_9844);
nand U10804 (N_10804,N_9382,N_9274);
or U10805 (N_10805,N_9642,N_9617);
xnor U10806 (N_10806,N_9002,N_9986);
or U10807 (N_10807,N_9680,N_9466);
nor U10808 (N_10808,N_9966,N_9445);
or U10809 (N_10809,N_9784,N_9749);
and U10810 (N_10810,N_9215,N_9498);
or U10811 (N_10811,N_9649,N_9306);
or U10812 (N_10812,N_9811,N_9696);
xnor U10813 (N_10813,N_9921,N_9014);
nand U10814 (N_10814,N_9619,N_9706);
or U10815 (N_10815,N_9406,N_9649);
nor U10816 (N_10816,N_9520,N_9402);
nand U10817 (N_10817,N_9803,N_9285);
nor U10818 (N_10818,N_9938,N_9502);
nand U10819 (N_10819,N_9339,N_9022);
nor U10820 (N_10820,N_9509,N_9754);
xor U10821 (N_10821,N_9035,N_9223);
or U10822 (N_10822,N_9990,N_9709);
nor U10823 (N_10823,N_9764,N_9417);
nor U10824 (N_10824,N_9237,N_9002);
nor U10825 (N_10825,N_9051,N_9473);
xor U10826 (N_10826,N_9453,N_9697);
nor U10827 (N_10827,N_9029,N_9126);
nand U10828 (N_10828,N_9197,N_9881);
and U10829 (N_10829,N_9260,N_9404);
nor U10830 (N_10830,N_9503,N_9385);
or U10831 (N_10831,N_9982,N_9560);
xnor U10832 (N_10832,N_9645,N_9016);
nor U10833 (N_10833,N_9656,N_9371);
or U10834 (N_10834,N_9272,N_9170);
or U10835 (N_10835,N_9784,N_9093);
nand U10836 (N_10836,N_9479,N_9792);
nand U10837 (N_10837,N_9525,N_9339);
nor U10838 (N_10838,N_9331,N_9668);
xnor U10839 (N_10839,N_9068,N_9488);
or U10840 (N_10840,N_9943,N_9614);
xor U10841 (N_10841,N_9586,N_9519);
nand U10842 (N_10842,N_9516,N_9427);
nand U10843 (N_10843,N_9927,N_9511);
nand U10844 (N_10844,N_9790,N_9099);
nor U10845 (N_10845,N_9513,N_9104);
and U10846 (N_10846,N_9619,N_9501);
nand U10847 (N_10847,N_9116,N_9612);
xnor U10848 (N_10848,N_9741,N_9910);
or U10849 (N_10849,N_9631,N_9482);
or U10850 (N_10850,N_9667,N_9580);
nor U10851 (N_10851,N_9747,N_9406);
or U10852 (N_10852,N_9204,N_9823);
and U10853 (N_10853,N_9923,N_9910);
and U10854 (N_10854,N_9392,N_9679);
nand U10855 (N_10855,N_9475,N_9649);
or U10856 (N_10856,N_9089,N_9640);
xor U10857 (N_10857,N_9839,N_9508);
or U10858 (N_10858,N_9464,N_9687);
nand U10859 (N_10859,N_9767,N_9121);
or U10860 (N_10860,N_9677,N_9858);
or U10861 (N_10861,N_9636,N_9872);
nand U10862 (N_10862,N_9506,N_9158);
and U10863 (N_10863,N_9652,N_9773);
xor U10864 (N_10864,N_9953,N_9402);
and U10865 (N_10865,N_9034,N_9145);
and U10866 (N_10866,N_9140,N_9033);
nor U10867 (N_10867,N_9234,N_9831);
xnor U10868 (N_10868,N_9997,N_9500);
nor U10869 (N_10869,N_9578,N_9163);
nor U10870 (N_10870,N_9338,N_9771);
or U10871 (N_10871,N_9241,N_9159);
nand U10872 (N_10872,N_9117,N_9287);
nor U10873 (N_10873,N_9876,N_9247);
and U10874 (N_10874,N_9871,N_9133);
or U10875 (N_10875,N_9585,N_9815);
nand U10876 (N_10876,N_9689,N_9604);
nand U10877 (N_10877,N_9817,N_9013);
nor U10878 (N_10878,N_9906,N_9849);
nor U10879 (N_10879,N_9797,N_9286);
nand U10880 (N_10880,N_9300,N_9296);
nor U10881 (N_10881,N_9541,N_9243);
nor U10882 (N_10882,N_9682,N_9601);
xor U10883 (N_10883,N_9779,N_9820);
nand U10884 (N_10884,N_9610,N_9296);
nand U10885 (N_10885,N_9876,N_9277);
or U10886 (N_10886,N_9346,N_9315);
or U10887 (N_10887,N_9862,N_9011);
xor U10888 (N_10888,N_9919,N_9557);
xor U10889 (N_10889,N_9717,N_9086);
or U10890 (N_10890,N_9960,N_9538);
xnor U10891 (N_10891,N_9635,N_9233);
and U10892 (N_10892,N_9439,N_9089);
nor U10893 (N_10893,N_9363,N_9192);
or U10894 (N_10894,N_9152,N_9155);
xnor U10895 (N_10895,N_9613,N_9847);
nand U10896 (N_10896,N_9868,N_9327);
nand U10897 (N_10897,N_9795,N_9803);
or U10898 (N_10898,N_9640,N_9974);
xor U10899 (N_10899,N_9721,N_9145);
nand U10900 (N_10900,N_9570,N_9961);
xor U10901 (N_10901,N_9056,N_9395);
nand U10902 (N_10902,N_9678,N_9390);
and U10903 (N_10903,N_9823,N_9296);
nor U10904 (N_10904,N_9360,N_9175);
nor U10905 (N_10905,N_9611,N_9232);
or U10906 (N_10906,N_9065,N_9712);
xor U10907 (N_10907,N_9506,N_9163);
nor U10908 (N_10908,N_9787,N_9834);
xor U10909 (N_10909,N_9749,N_9453);
or U10910 (N_10910,N_9807,N_9591);
nand U10911 (N_10911,N_9706,N_9499);
xnor U10912 (N_10912,N_9477,N_9864);
nor U10913 (N_10913,N_9449,N_9736);
or U10914 (N_10914,N_9444,N_9749);
nor U10915 (N_10915,N_9488,N_9938);
and U10916 (N_10916,N_9337,N_9446);
xnor U10917 (N_10917,N_9061,N_9074);
nand U10918 (N_10918,N_9576,N_9920);
or U10919 (N_10919,N_9064,N_9699);
nor U10920 (N_10920,N_9042,N_9114);
nor U10921 (N_10921,N_9088,N_9648);
and U10922 (N_10922,N_9845,N_9724);
and U10923 (N_10923,N_9587,N_9296);
nand U10924 (N_10924,N_9278,N_9556);
and U10925 (N_10925,N_9697,N_9220);
nand U10926 (N_10926,N_9360,N_9967);
and U10927 (N_10927,N_9169,N_9116);
nand U10928 (N_10928,N_9611,N_9878);
and U10929 (N_10929,N_9502,N_9406);
and U10930 (N_10930,N_9594,N_9447);
nor U10931 (N_10931,N_9001,N_9374);
nand U10932 (N_10932,N_9000,N_9808);
or U10933 (N_10933,N_9213,N_9634);
xnor U10934 (N_10934,N_9290,N_9712);
and U10935 (N_10935,N_9836,N_9339);
xor U10936 (N_10936,N_9484,N_9454);
and U10937 (N_10937,N_9282,N_9160);
or U10938 (N_10938,N_9180,N_9430);
xor U10939 (N_10939,N_9494,N_9981);
or U10940 (N_10940,N_9108,N_9562);
nand U10941 (N_10941,N_9096,N_9385);
xnor U10942 (N_10942,N_9547,N_9426);
xor U10943 (N_10943,N_9562,N_9445);
or U10944 (N_10944,N_9447,N_9705);
nand U10945 (N_10945,N_9025,N_9578);
nand U10946 (N_10946,N_9331,N_9982);
and U10947 (N_10947,N_9818,N_9031);
and U10948 (N_10948,N_9172,N_9467);
and U10949 (N_10949,N_9580,N_9012);
nor U10950 (N_10950,N_9730,N_9219);
xnor U10951 (N_10951,N_9218,N_9724);
xnor U10952 (N_10952,N_9930,N_9322);
or U10953 (N_10953,N_9335,N_9929);
and U10954 (N_10954,N_9738,N_9189);
nand U10955 (N_10955,N_9624,N_9396);
nor U10956 (N_10956,N_9713,N_9159);
nand U10957 (N_10957,N_9531,N_9580);
xor U10958 (N_10958,N_9415,N_9812);
nand U10959 (N_10959,N_9101,N_9750);
or U10960 (N_10960,N_9136,N_9751);
nand U10961 (N_10961,N_9886,N_9577);
nor U10962 (N_10962,N_9792,N_9371);
nor U10963 (N_10963,N_9602,N_9933);
nor U10964 (N_10964,N_9431,N_9881);
nand U10965 (N_10965,N_9868,N_9163);
and U10966 (N_10966,N_9014,N_9285);
and U10967 (N_10967,N_9954,N_9034);
nand U10968 (N_10968,N_9753,N_9406);
nor U10969 (N_10969,N_9009,N_9946);
xor U10970 (N_10970,N_9610,N_9698);
nor U10971 (N_10971,N_9285,N_9757);
xnor U10972 (N_10972,N_9054,N_9849);
or U10973 (N_10973,N_9367,N_9987);
and U10974 (N_10974,N_9189,N_9113);
xnor U10975 (N_10975,N_9034,N_9708);
and U10976 (N_10976,N_9498,N_9357);
xnor U10977 (N_10977,N_9472,N_9575);
or U10978 (N_10978,N_9394,N_9309);
or U10979 (N_10979,N_9000,N_9982);
and U10980 (N_10980,N_9234,N_9586);
nor U10981 (N_10981,N_9839,N_9318);
nor U10982 (N_10982,N_9224,N_9129);
and U10983 (N_10983,N_9001,N_9857);
xnor U10984 (N_10984,N_9447,N_9627);
or U10985 (N_10985,N_9033,N_9787);
nor U10986 (N_10986,N_9228,N_9770);
nand U10987 (N_10987,N_9848,N_9155);
or U10988 (N_10988,N_9222,N_9345);
nor U10989 (N_10989,N_9182,N_9760);
xnor U10990 (N_10990,N_9019,N_9232);
and U10991 (N_10991,N_9071,N_9521);
xor U10992 (N_10992,N_9092,N_9293);
and U10993 (N_10993,N_9626,N_9764);
nand U10994 (N_10994,N_9532,N_9089);
nor U10995 (N_10995,N_9321,N_9090);
and U10996 (N_10996,N_9421,N_9780);
or U10997 (N_10997,N_9587,N_9655);
nand U10998 (N_10998,N_9817,N_9075);
nand U10999 (N_10999,N_9498,N_9154);
nor U11000 (N_11000,N_10613,N_10293);
and U11001 (N_11001,N_10443,N_10087);
or U11002 (N_11002,N_10980,N_10010);
xor U11003 (N_11003,N_10821,N_10681);
and U11004 (N_11004,N_10792,N_10409);
nand U11005 (N_11005,N_10202,N_10193);
and U11006 (N_11006,N_10045,N_10852);
and U11007 (N_11007,N_10510,N_10320);
nand U11008 (N_11008,N_10813,N_10748);
nor U11009 (N_11009,N_10548,N_10798);
xor U11010 (N_11010,N_10909,N_10873);
nor U11011 (N_11011,N_10250,N_10165);
or U11012 (N_11012,N_10492,N_10329);
nand U11013 (N_11013,N_10576,N_10172);
or U11014 (N_11014,N_10503,N_10338);
and U11015 (N_11015,N_10500,N_10220);
nand U11016 (N_11016,N_10358,N_10918);
xnor U11017 (N_11017,N_10116,N_10413);
and U11018 (N_11018,N_10461,N_10625);
and U11019 (N_11019,N_10023,N_10652);
and U11020 (N_11020,N_10296,N_10022);
xor U11021 (N_11021,N_10152,N_10251);
nand U11022 (N_11022,N_10407,N_10114);
and U11023 (N_11023,N_10458,N_10505);
and U11024 (N_11024,N_10267,N_10828);
nor U11025 (N_11025,N_10969,N_10680);
xnor U11026 (N_11026,N_10654,N_10089);
nor U11027 (N_11027,N_10121,N_10710);
or U11028 (N_11028,N_10683,N_10611);
or U11029 (N_11029,N_10014,N_10769);
and U11030 (N_11030,N_10782,N_10190);
nor U11031 (N_11031,N_10124,N_10770);
nor U11032 (N_11032,N_10965,N_10182);
and U11033 (N_11033,N_10192,N_10947);
and U11034 (N_11034,N_10000,N_10647);
and U11035 (N_11035,N_10478,N_10056);
and U11036 (N_11036,N_10118,N_10498);
and U11037 (N_11037,N_10765,N_10860);
nand U11038 (N_11038,N_10092,N_10411);
nor U11039 (N_11039,N_10968,N_10203);
nor U11040 (N_11040,N_10279,N_10558);
and U11041 (N_11041,N_10024,N_10051);
nor U11042 (N_11042,N_10110,N_10146);
nand U11043 (N_11043,N_10265,N_10093);
xor U11044 (N_11044,N_10357,N_10896);
xnor U11045 (N_11045,N_10583,N_10823);
or U11046 (N_11046,N_10878,N_10039);
and U11047 (N_11047,N_10672,N_10527);
nor U11048 (N_11048,N_10166,N_10509);
and U11049 (N_11049,N_10313,N_10630);
and U11050 (N_11050,N_10696,N_10222);
nor U11051 (N_11051,N_10434,N_10942);
nor U11052 (N_11052,N_10266,N_10585);
nand U11053 (N_11053,N_10833,N_10645);
nor U11054 (N_11054,N_10481,N_10164);
xnor U11055 (N_11055,N_10186,N_10106);
nor U11056 (N_11056,N_10890,N_10514);
or U11057 (N_11057,N_10030,N_10392);
or U11058 (N_11058,N_10479,N_10412);
and U11059 (N_11059,N_10759,N_10516);
or U11060 (N_11060,N_10950,N_10390);
and U11061 (N_11061,N_10290,N_10788);
nand U11062 (N_11062,N_10047,N_10758);
nor U11063 (N_11063,N_10996,N_10394);
nor U11064 (N_11064,N_10695,N_10634);
nand U11065 (N_11065,N_10231,N_10803);
nor U11066 (N_11066,N_10404,N_10662);
nand U11067 (N_11067,N_10818,N_10767);
and U11068 (N_11068,N_10998,N_10301);
nand U11069 (N_11069,N_10649,N_10447);
xnor U11070 (N_11070,N_10066,N_10774);
xnor U11071 (N_11071,N_10491,N_10825);
or U11072 (N_11072,N_10892,N_10620);
nor U11073 (N_11073,N_10819,N_10327);
nor U11074 (N_11074,N_10207,N_10610);
and U11075 (N_11075,N_10013,N_10960);
nand U11076 (N_11076,N_10371,N_10799);
and U11077 (N_11077,N_10167,N_10303);
xnor U11078 (N_11078,N_10168,N_10115);
and U11079 (N_11079,N_10869,N_10258);
xor U11080 (N_11080,N_10080,N_10525);
or U11081 (N_11081,N_10966,N_10851);
and U11082 (N_11082,N_10643,N_10460);
and U11083 (N_11083,N_10216,N_10981);
nand U11084 (N_11084,N_10016,N_10556);
nand U11085 (N_11085,N_10577,N_10276);
and U11086 (N_11086,N_10786,N_10011);
and U11087 (N_11087,N_10249,N_10101);
nor U11088 (N_11088,N_10686,N_10776);
nand U11089 (N_11089,N_10067,N_10651);
nand U11090 (N_11090,N_10017,N_10477);
xnor U11091 (N_11091,N_10836,N_10797);
xor U11092 (N_11092,N_10345,N_10719);
nor U11093 (N_11093,N_10440,N_10952);
nand U11094 (N_11094,N_10126,N_10424);
xor U11095 (N_11095,N_10480,N_10316);
and U11096 (N_11096,N_10377,N_10853);
xnor U11097 (N_11097,N_10230,N_10344);
nor U11098 (N_11098,N_10690,N_10554);
nor U11099 (N_11099,N_10910,N_10495);
nand U11100 (N_11100,N_10383,N_10507);
nor U11101 (N_11101,N_10711,N_10692);
nor U11102 (N_11102,N_10395,N_10897);
xnor U11103 (N_11103,N_10083,N_10032);
and U11104 (N_11104,N_10037,N_10761);
and U11105 (N_11105,N_10349,N_10336);
nand U11106 (N_11106,N_10579,N_10433);
xnor U11107 (N_11107,N_10086,N_10725);
or U11108 (N_11108,N_10923,N_10660);
nor U11109 (N_11109,N_10065,N_10730);
and U11110 (N_11110,N_10924,N_10564);
nand U11111 (N_11111,N_10841,N_10693);
and U11112 (N_11112,N_10062,N_10713);
or U11113 (N_11113,N_10551,N_10294);
nand U11114 (N_11114,N_10831,N_10973);
nand U11115 (N_11115,N_10224,N_10031);
nand U11116 (N_11116,N_10811,N_10367);
nand U11117 (N_11117,N_10309,N_10925);
xor U11118 (N_11118,N_10072,N_10351);
and U11119 (N_11119,N_10459,N_10578);
xnor U11120 (N_11120,N_10675,N_10627);
nand U11121 (N_11121,N_10096,N_10350);
and U11122 (N_11122,N_10600,N_10085);
or U11123 (N_11123,N_10260,N_10609);
or U11124 (N_11124,N_10866,N_10469);
nand U11125 (N_11125,N_10341,N_10663);
nand U11126 (N_11126,N_10314,N_10337);
or U11127 (N_11127,N_10317,N_10361);
or U11128 (N_11128,N_10637,N_10482);
and U11129 (N_11129,N_10687,N_10257);
nor U11130 (N_11130,N_10347,N_10252);
xor U11131 (N_11131,N_10355,N_10009);
nor U11132 (N_11132,N_10886,N_10330);
nor U11133 (N_11133,N_10817,N_10985);
or U11134 (N_11134,N_10468,N_10793);
or U11135 (N_11135,N_10536,N_10426);
or U11136 (N_11136,N_10927,N_10233);
nand U11137 (N_11137,N_10976,N_10606);
or U11138 (N_11138,N_10239,N_10034);
xnor U11139 (N_11139,N_10236,N_10905);
or U11140 (N_11140,N_10598,N_10493);
nand U11141 (N_11141,N_10242,N_10750);
and U11142 (N_11142,N_10162,N_10059);
and U11143 (N_11143,N_10670,N_10891);
or U11144 (N_11144,N_10561,N_10073);
or U11145 (N_11145,N_10908,N_10365);
xnor U11146 (N_11146,N_10139,N_10406);
nand U11147 (N_11147,N_10153,N_10999);
xor U11148 (N_11148,N_10832,N_10035);
nor U11149 (N_11149,N_10524,N_10553);
and U11150 (N_11150,N_10544,N_10179);
or U11151 (N_11151,N_10136,N_10074);
and U11152 (N_11152,N_10437,N_10213);
xor U11153 (N_11153,N_10715,N_10123);
or U11154 (N_11154,N_10784,N_10900);
or U11155 (N_11155,N_10006,N_10863);
nand U11156 (N_11156,N_10396,N_10682);
xor U11157 (N_11157,N_10570,N_10688);
or U11158 (N_11158,N_10785,N_10955);
or U11159 (N_11159,N_10655,N_10425);
or U11160 (N_11160,N_10839,N_10951);
nand U11161 (N_11161,N_10405,N_10895);
or U11162 (N_11162,N_10388,N_10027);
xnor U11163 (N_11163,N_10082,N_10874);
nor U11164 (N_11164,N_10993,N_10760);
nand U11165 (N_11165,N_10323,N_10824);
nand U11166 (N_11166,N_10604,N_10967);
or U11167 (N_11167,N_10929,N_10418);
and U11168 (N_11168,N_10467,N_10335);
and U11169 (N_11169,N_10804,N_10200);
xor U11170 (N_11170,N_10235,N_10472);
xor U11171 (N_11171,N_10608,N_10403);
nor U11172 (N_11172,N_10150,N_10444);
and U11173 (N_11173,N_10665,N_10992);
or U11174 (N_11174,N_10870,N_10812);
or U11175 (N_11175,N_10436,N_10633);
xor U11176 (N_11176,N_10378,N_10149);
nand U11177 (N_11177,N_10736,N_10724);
xnor U11178 (N_11178,N_10861,N_10684);
or U11179 (N_11179,N_10623,N_10452);
nand U11180 (N_11180,N_10272,N_10398);
and U11181 (N_11181,N_10125,N_10454);
nand U11182 (N_11182,N_10270,N_10937);
or U11183 (N_11183,N_10944,N_10593);
and U11184 (N_11184,N_10691,N_10312);
and U11185 (N_11185,N_10801,N_10989);
nand U11186 (N_11186,N_10120,N_10595);
xnor U11187 (N_11187,N_10094,N_10701);
nand U11188 (N_11188,N_10586,N_10281);
nor U11189 (N_11189,N_10169,N_10076);
xnor U11190 (N_11190,N_10020,N_10939);
xnor U11191 (N_11191,N_10129,N_10936);
or U11192 (N_11192,N_10802,N_10446);
nand U11193 (N_11193,N_10112,N_10780);
nor U11194 (N_11194,N_10240,N_10535);
or U11195 (N_11195,N_10151,N_10147);
or U11196 (N_11196,N_10285,N_10829);
or U11197 (N_11197,N_10614,N_10685);
xnor U11198 (N_11198,N_10990,N_10362);
nor U11199 (N_11199,N_10408,N_10397);
nand U11200 (N_11200,N_10143,N_10789);
xor U11201 (N_11201,N_10048,N_10835);
nor U11202 (N_11202,N_10745,N_10714);
xor U11203 (N_11203,N_10400,N_10209);
nor U11204 (N_11204,N_10912,N_10716);
xor U11205 (N_11205,N_10529,N_10640);
and U11206 (N_11206,N_10103,N_10588);
nor U11207 (N_11207,N_10226,N_10201);
nor U11208 (N_11208,N_10580,N_10133);
nor U11209 (N_11209,N_10310,N_10060);
xnor U11210 (N_11210,N_10015,N_10735);
nand U11211 (N_11211,N_10455,N_10858);
and U11212 (N_11212,N_10849,N_10539);
nand U11213 (N_11213,N_10679,N_10528);
nor U11214 (N_11214,N_10517,N_10484);
xor U11215 (N_11215,N_10420,N_10218);
xnor U11216 (N_11216,N_10068,N_10559);
xnor U11217 (N_11217,N_10644,N_10615);
nor U11218 (N_11218,N_10269,N_10738);
xnor U11219 (N_11219,N_10307,N_10783);
xor U11220 (N_11220,N_10806,N_10353);
nand U11221 (N_11221,N_10005,N_10555);
nor U11222 (N_11222,N_10273,N_10184);
and U11223 (N_11223,N_10487,N_10642);
nand U11224 (N_11224,N_10499,N_10287);
nor U11225 (N_11225,N_10042,N_10794);
nor U11226 (N_11226,N_10210,N_10844);
or U11227 (N_11227,N_10882,N_10913);
nor U11228 (N_11228,N_10840,N_10864);
nor U11229 (N_11229,N_10160,N_10919);
nand U11230 (N_11230,N_10698,N_10470);
or U11231 (N_11231,N_10826,N_10668);
or U11232 (N_11232,N_10331,N_10366);
and U11233 (N_11233,N_10275,N_10225);
or U11234 (N_11234,N_10175,N_10485);
nand U11235 (N_11235,N_10277,N_10628);
and U11236 (N_11236,N_10875,N_10261);
and U11237 (N_11237,N_10324,N_10100);
xnor U11238 (N_11238,N_10475,N_10621);
nand U11239 (N_11239,N_10865,N_10938);
and U11240 (N_11240,N_10019,N_10195);
nand U11241 (N_11241,N_10214,N_10626);
and U11242 (N_11242,N_10049,N_10234);
and U11243 (N_11243,N_10959,N_10515);
xnor U11244 (N_11244,N_10537,N_10755);
nand U11245 (N_11245,N_10709,N_10565);
and U11246 (N_11246,N_10862,N_10326);
nor U11247 (N_11247,N_10837,N_10208);
xnor U11248 (N_11248,N_10846,N_10943);
xor U11249 (N_11249,N_10787,N_10872);
nand U11250 (N_11250,N_10779,N_10174);
nor U11251 (N_11251,N_10917,N_10305);
nand U11252 (N_11252,N_10641,N_10549);
nor U11253 (N_11253,N_10752,N_10369);
xor U11254 (N_11254,N_10898,N_10757);
nor U11255 (N_11255,N_10489,N_10298);
and U11256 (N_11256,N_10359,N_10575);
nor U11257 (N_11257,N_10742,N_10328);
nand U11258 (N_11258,N_10971,N_10636);
or U11259 (N_11259,N_10734,N_10363);
and U11260 (N_11260,N_10368,N_10903);
xnor U11261 (N_11261,N_10930,N_10988);
and U11262 (N_11262,N_10007,N_10533);
and U11263 (N_11263,N_10243,N_10931);
nand U11264 (N_11264,N_10325,N_10531);
or U11265 (N_11265,N_10666,N_10340);
and U11266 (N_11266,N_10171,N_10494);
xor U11267 (N_11267,N_10227,N_10962);
or U11268 (N_11268,N_10843,N_10091);
or U11269 (N_11269,N_10954,N_10808);
or U11270 (N_11270,N_10712,N_10661);
or U11271 (N_11271,N_10753,N_10154);
and U11272 (N_11272,N_10248,N_10159);
xnor U11273 (N_11273,N_10135,N_10430);
and U11274 (N_11274,N_10380,N_10158);
and U11275 (N_11275,N_10963,N_10255);
nand U11276 (N_11276,N_10122,N_10763);
nand U11277 (N_11277,N_10722,N_10127);
or U11278 (N_11278,N_10809,N_10057);
and U11279 (N_11279,N_10071,N_10183);
xnor U11280 (N_11280,N_10970,N_10379);
and U11281 (N_11281,N_10283,N_10607);
or U11282 (N_11282,N_10194,N_10699);
nor U11283 (N_11283,N_10036,N_10393);
xor U11284 (N_11284,N_10972,N_10997);
nand U11285 (N_11285,N_10196,N_10311);
or U11286 (N_11286,N_10004,N_10185);
nand U11287 (N_11287,N_10948,N_10881);
nor U11288 (N_11288,N_10737,N_10102);
and U11289 (N_11289,N_10206,N_10348);
nand U11290 (N_11290,N_10814,N_10376);
nor U11291 (N_11291,N_10282,N_10263);
and U11292 (N_11292,N_10416,N_10958);
nor U11293 (N_11293,N_10717,N_10058);
nand U11294 (N_11294,N_10658,N_10271);
xor U11295 (N_11295,N_10117,N_10639);
nand U11296 (N_11296,N_10465,N_10098);
nand U11297 (N_11297,N_10474,N_10847);
or U11298 (N_11298,N_10935,N_10868);
and U11299 (N_11299,N_10212,N_10464);
or U11300 (N_11300,N_10689,N_10953);
nor U11301 (N_11301,N_10278,N_10956);
or U11302 (N_11302,N_10791,N_10704);
xor U11303 (N_11303,N_10423,N_10574);
xnor U11304 (N_11304,N_10887,N_10591);
nand U11305 (N_11305,N_10731,N_10673);
nor U11306 (N_11306,N_10046,N_10702);
xnor U11307 (N_11307,N_10664,N_10108);
and U11308 (N_11308,N_10563,N_10176);
nand U11309 (N_11309,N_10879,N_10486);
or U11310 (N_11310,N_10422,N_10572);
nand U11311 (N_11311,N_10384,N_10095);
xor U11312 (N_11312,N_10856,N_10070);
nand U11313 (N_11313,N_10697,N_10163);
and U11314 (N_11314,N_10211,N_10974);
or U11315 (N_11315,N_10375,N_10616);
nor U11316 (N_11316,N_10228,N_10262);
and U11317 (N_11317,N_10995,N_10820);
xnor U11318 (N_11318,N_10850,N_10546);
and U11319 (N_11319,N_10582,N_10932);
nor U11320 (N_11320,N_10914,N_10448);
nand U11321 (N_11321,N_10352,N_10771);
and U11322 (N_11322,N_10128,N_10822);
nor U11323 (N_11323,N_10427,N_10155);
nor U11324 (N_11324,N_10318,N_10300);
nor U11325 (N_11325,N_10617,N_10435);
nor U11326 (N_11326,N_10573,N_10188);
or U11327 (N_11327,N_10916,N_10597);
nand U11328 (N_11328,N_10677,N_10256);
nor U11329 (N_11329,N_10650,N_10041);
or U11330 (N_11330,N_10994,N_10244);
xor U11331 (N_11331,N_10867,N_10297);
or U11332 (N_11332,N_10883,N_10534);
and U11333 (N_11333,N_10830,N_10807);
xor U11334 (N_11334,N_10781,N_10854);
nor U11335 (N_11335,N_10321,N_10674);
or U11336 (N_11336,N_10456,N_10401);
and U11337 (N_11337,N_10569,N_10386);
and U11338 (N_11338,N_10274,N_10542);
xor U11339 (N_11339,N_10928,N_10922);
xnor U11340 (N_11340,N_10978,N_10532);
xnor U11341 (N_11341,N_10229,N_10957);
xnor U11342 (N_11342,N_10915,N_10333);
xnor U11343 (N_11343,N_10526,N_10302);
and U11344 (N_11344,N_10859,N_10247);
and U11345 (N_11345,N_10421,N_10343);
or U11346 (N_11346,N_10246,N_10523);
nand U11347 (N_11347,N_10088,N_10463);
and U11348 (N_11348,N_10221,N_10099);
or U11349 (N_11349,N_10084,N_10727);
nor U11350 (N_11350,N_10439,N_10933);
or U11351 (N_11351,N_10907,N_10571);
xor U11352 (N_11352,N_10871,N_10842);
nand U11353 (N_11353,N_10964,N_10519);
xor U11354 (N_11354,N_10198,N_10618);
or U11355 (N_11355,N_10827,N_10104);
nand U11356 (N_11356,N_10170,N_10596);
xor U11357 (N_11357,N_10148,N_10504);
xor U11358 (N_11358,N_10590,N_10718);
nor U11359 (N_11359,N_10857,N_10599);
or U11360 (N_11360,N_10483,N_10280);
nor U11361 (N_11361,N_10237,N_10217);
nor U11362 (N_11362,N_10946,N_10415);
nand U11363 (N_11363,N_10342,N_10410);
or U11364 (N_11364,N_10197,N_10291);
and U11365 (N_11365,N_10254,N_10669);
and U11366 (N_11366,N_10161,N_10920);
nand U11367 (N_11367,N_10417,N_10238);
and U11368 (N_11368,N_10215,N_10445);
and U11369 (N_11369,N_10138,N_10021);
nor U11370 (N_11370,N_10977,N_10471);
or U11371 (N_11371,N_10732,N_10205);
nand U11372 (N_11372,N_10877,N_10855);
or U11373 (N_11373,N_10466,N_10678);
and U11374 (N_11374,N_10315,N_10339);
nor U11375 (N_11375,N_10552,N_10502);
nand U11376 (N_11376,N_10543,N_10488);
nand U11377 (N_11377,N_10961,N_10079);
or U11378 (N_11378,N_10921,N_10044);
nand U11379 (N_11379,N_10845,N_10181);
and U11380 (N_11380,N_10097,N_10381);
nand U11381 (N_11381,N_10754,N_10657);
nand U11382 (N_11382,N_10442,N_10880);
or U11383 (N_11383,N_10901,N_10180);
or U11384 (N_11384,N_10986,N_10772);
nor U11385 (N_11385,N_10733,N_10295);
and U11386 (N_11386,N_10746,N_10008);
nand U11387 (N_11387,N_10834,N_10720);
xor U11388 (N_11388,N_10530,N_10449);
xor U11389 (N_11389,N_10512,N_10002);
nand U11390 (N_11390,N_10743,N_10253);
and U11391 (N_11391,N_10656,N_10612);
and U11392 (N_11392,N_10054,N_10584);
nand U11393 (N_11393,N_10040,N_10795);
nor U11394 (N_11394,N_10137,N_10764);
and U11395 (N_11395,N_10043,N_10659);
xor U11396 (N_11396,N_10132,N_10906);
nand U11397 (N_11397,N_10063,N_10299);
xnor U11398 (N_11398,N_10204,N_10025);
and U11399 (N_11399,N_10888,N_10268);
xnor U11400 (N_11400,N_10762,N_10773);
nor U11401 (N_11401,N_10382,N_10700);
and U11402 (N_11402,N_10726,N_10744);
and U11403 (N_11403,N_10721,N_10520);
and U11404 (N_11404,N_10457,N_10518);
or U11405 (N_11405,N_10003,N_10926);
nor U11406 (N_11406,N_10740,N_10131);
nor U11407 (N_11407,N_10145,N_10473);
nor U11408 (N_11408,N_10540,N_10245);
and U11409 (N_11409,N_10723,N_10428);
nand U11410 (N_11410,N_10144,N_10191);
nand U11411 (N_11411,N_10438,N_10741);
nand U11412 (N_11412,N_10728,N_10306);
or U11413 (N_11413,N_10777,N_10676);
nand U11414 (N_11414,N_10602,N_10756);
nor U11415 (N_11415,N_10241,N_10451);
xor U11416 (N_11416,N_10012,N_10157);
nand U11417 (N_11417,N_10360,N_10624);
xnor U11418 (N_11418,N_10441,N_10432);
nor U11419 (N_11419,N_10081,N_10538);
nor U11420 (N_11420,N_10052,N_10550);
or U11421 (N_11421,N_10508,N_10156);
and U11422 (N_11422,N_10134,N_10506);
nor U11423 (N_11423,N_10566,N_10810);
nand U11424 (N_11424,N_10055,N_10983);
and U11425 (N_11425,N_10838,N_10706);
and U11426 (N_11426,N_10934,N_10587);
or U11427 (N_11427,N_10346,N_10107);
or U11428 (N_11428,N_10501,N_10130);
and U11429 (N_11429,N_10815,N_10778);
xor U11430 (N_11430,N_10389,N_10631);
nor U11431 (N_11431,N_10982,N_10264);
xor U11432 (N_11432,N_10635,N_10075);
and U11433 (N_11433,N_10142,N_10026);
and U11434 (N_11434,N_10173,N_10638);
or U11435 (N_11435,N_10694,N_10402);
and U11436 (N_11436,N_10061,N_10547);
nand U11437 (N_11437,N_10703,N_10545);
nand U11438 (N_11438,N_10414,N_10141);
or U11439 (N_11439,N_10219,N_10028);
or U11440 (N_11440,N_10450,N_10001);
xor U11441 (N_11441,N_10889,N_10592);
nand U11442 (N_11442,N_10419,N_10018);
or U11443 (N_11443,N_10790,N_10667);
xnor U11444 (N_11444,N_10033,N_10705);
nor U11445 (N_11445,N_10385,N_10729);
xnor U11446 (N_11446,N_10111,N_10632);
and U11447 (N_11447,N_10601,N_10749);
nor U11448 (N_11448,N_10077,N_10334);
nand U11449 (N_11449,N_10286,N_10289);
nor U11450 (N_11450,N_10304,N_10991);
nor U11451 (N_11451,N_10177,N_10902);
nand U11452 (N_11452,N_10816,N_10453);
and U11453 (N_11453,N_10374,N_10622);
nand U11454 (N_11454,N_10568,N_10399);
and U11455 (N_11455,N_10805,N_10292);
nand U11456 (N_11456,N_10911,N_10322);
nand U11457 (N_11457,N_10557,N_10775);
xnor U11458 (N_11458,N_10391,N_10140);
or U11459 (N_11459,N_10053,N_10387);
nor U11460 (N_11460,N_10899,N_10050);
nor U11461 (N_11461,N_10490,N_10751);
xnor U11462 (N_11462,N_10603,N_10356);
nand U11463 (N_11463,N_10069,N_10708);
and U11464 (N_11464,N_10766,N_10370);
or U11465 (N_11465,N_10284,N_10187);
xnor U11466 (N_11466,N_10739,N_10288);
nand U11467 (N_11467,N_10768,N_10653);
or U11468 (N_11468,N_10945,N_10354);
nor U11469 (N_11469,N_10648,N_10521);
and U11470 (N_11470,N_10038,N_10984);
xor U11471 (N_11471,N_10090,N_10671);
and U11472 (N_11472,N_10884,N_10885);
or U11473 (N_11473,N_10646,N_10594);
and U11474 (N_11474,N_10605,N_10178);
nor U11475 (N_11475,N_10319,N_10522);
or U11476 (N_11476,N_10949,N_10078);
xor U11477 (N_11477,N_10496,N_10979);
or U11478 (N_11478,N_10747,N_10105);
nor U11479 (N_11479,N_10332,N_10796);
or U11480 (N_11480,N_10541,N_10029);
xnor U11481 (N_11481,N_10462,N_10876);
and U11482 (N_11482,N_10189,N_10431);
xnor U11483 (N_11483,N_10119,N_10560);
and U11484 (N_11484,N_10975,N_10941);
or U11485 (N_11485,N_10373,N_10199);
or U11486 (N_11486,N_10308,N_10707);
and U11487 (N_11487,N_10513,N_10562);
nor U11488 (N_11488,N_10476,N_10109);
and U11489 (N_11489,N_10987,N_10581);
or U11490 (N_11490,N_10589,N_10904);
or U11491 (N_11491,N_10893,N_10372);
and U11492 (N_11492,N_10567,N_10064);
xnor U11493 (N_11493,N_10232,N_10364);
or U11494 (N_11494,N_10511,N_10800);
and U11495 (N_11495,N_10223,N_10894);
and U11496 (N_11496,N_10259,N_10497);
xnor U11497 (N_11497,N_10940,N_10629);
nand U11498 (N_11498,N_10429,N_10848);
or U11499 (N_11499,N_10113,N_10619);
nand U11500 (N_11500,N_10349,N_10274);
nor U11501 (N_11501,N_10801,N_10824);
and U11502 (N_11502,N_10672,N_10483);
and U11503 (N_11503,N_10424,N_10393);
nand U11504 (N_11504,N_10679,N_10915);
nor U11505 (N_11505,N_10291,N_10269);
or U11506 (N_11506,N_10953,N_10998);
xnor U11507 (N_11507,N_10266,N_10877);
xor U11508 (N_11508,N_10471,N_10828);
nand U11509 (N_11509,N_10257,N_10394);
nor U11510 (N_11510,N_10019,N_10855);
nand U11511 (N_11511,N_10804,N_10012);
and U11512 (N_11512,N_10392,N_10348);
and U11513 (N_11513,N_10456,N_10332);
xnor U11514 (N_11514,N_10709,N_10010);
nand U11515 (N_11515,N_10075,N_10747);
nand U11516 (N_11516,N_10373,N_10614);
and U11517 (N_11517,N_10028,N_10327);
or U11518 (N_11518,N_10766,N_10034);
nor U11519 (N_11519,N_10383,N_10942);
xor U11520 (N_11520,N_10084,N_10535);
nor U11521 (N_11521,N_10076,N_10803);
xnor U11522 (N_11522,N_10555,N_10944);
and U11523 (N_11523,N_10880,N_10265);
nor U11524 (N_11524,N_10462,N_10656);
or U11525 (N_11525,N_10671,N_10254);
nor U11526 (N_11526,N_10269,N_10165);
nor U11527 (N_11527,N_10170,N_10075);
nor U11528 (N_11528,N_10756,N_10239);
and U11529 (N_11529,N_10039,N_10444);
xor U11530 (N_11530,N_10561,N_10890);
nand U11531 (N_11531,N_10745,N_10901);
nor U11532 (N_11532,N_10238,N_10109);
nor U11533 (N_11533,N_10460,N_10573);
xnor U11534 (N_11534,N_10914,N_10836);
nor U11535 (N_11535,N_10357,N_10630);
or U11536 (N_11536,N_10621,N_10798);
nand U11537 (N_11537,N_10563,N_10497);
and U11538 (N_11538,N_10116,N_10824);
nand U11539 (N_11539,N_10892,N_10621);
or U11540 (N_11540,N_10538,N_10835);
or U11541 (N_11541,N_10570,N_10150);
nand U11542 (N_11542,N_10628,N_10560);
nor U11543 (N_11543,N_10667,N_10779);
or U11544 (N_11544,N_10284,N_10578);
or U11545 (N_11545,N_10180,N_10760);
or U11546 (N_11546,N_10955,N_10394);
or U11547 (N_11547,N_10674,N_10947);
xor U11548 (N_11548,N_10458,N_10419);
or U11549 (N_11549,N_10738,N_10306);
nand U11550 (N_11550,N_10743,N_10727);
nor U11551 (N_11551,N_10006,N_10879);
or U11552 (N_11552,N_10832,N_10891);
xnor U11553 (N_11553,N_10535,N_10089);
or U11554 (N_11554,N_10480,N_10125);
xnor U11555 (N_11555,N_10470,N_10768);
nor U11556 (N_11556,N_10305,N_10293);
nand U11557 (N_11557,N_10608,N_10379);
and U11558 (N_11558,N_10148,N_10641);
nand U11559 (N_11559,N_10067,N_10782);
nor U11560 (N_11560,N_10248,N_10993);
and U11561 (N_11561,N_10746,N_10711);
or U11562 (N_11562,N_10430,N_10862);
and U11563 (N_11563,N_10987,N_10409);
nand U11564 (N_11564,N_10779,N_10715);
nor U11565 (N_11565,N_10950,N_10421);
nor U11566 (N_11566,N_10492,N_10654);
xor U11567 (N_11567,N_10831,N_10514);
nor U11568 (N_11568,N_10936,N_10993);
or U11569 (N_11569,N_10433,N_10127);
nor U11570 (N_11570,N_10007,N_10947);
or U11571 (N_11571,N_10837,N_10241);
and U11572 (N_11572,N_10847,N_10690);
and U11573 (N_11573,N_10027,N_10142);
xnor U11574 (N_11574,N_10217,N_10317);
nor U11575 (N_11575,N_10208,N_10476);
xor U11576 (N_11576,N_10179,N_10470);
nor U11577 (N_11577,N_10131,N_10060);
and U11578 (N_11578,N_10455,N_10749);
or U11579 (N_11579,N_10234,N_10271);
xnor U11580 (N_11580,N_10290,N_10388);
nand U11581 (N_11581,N_10718,N_10615);
nand U11582 (N_11582,N_10061,N_10738);
nand U11583 (N_11583,N_10844,N_10926);
nand U11584 (N_11584,N_10458,N_10797);
and U11585 (N_11585,N_10923,N_10817);
and U11586 (N_11586,N_10070,N_10435);
xor U11587 (N_11587,N_10765,N_10603);
xor U11588 (N_11588,N_10963,N_10648);
nor U11589 (N_11589,N_10362,N_10368);
nor U11590 (N_11590,N_10677,N_10414);
xnor U11591 (N_11591,N_10918,N_10319);
and U11592 (N_11592,N_10212,N_10993);
or U11593 (N_11593,N_10599,N_10866);
nor U11594 (N_11594,N_10640,N_10463);
and U11595 (N_11595,N_10135,N_10633);
and U11596 (N_11596,N_10009,N_10421);
or U11597 (N_11597,N_10068,N_10162);
xor U11598 (N_11598,N_10970,N_10884);
nor U11599 (N_11599,N_10102,N_10634);
xnor U11600 (N_11600,N_10652,N_10026);
xor U11601 (N_11601,N_10457,N_10593);
nand U11602 (N_11602,N_10771,N_10541);
or U11603 (N_11603,N_10241,N_10635);
and U11604 (N_11604,N_10181,N_10722);
or U11605 (N_11605,N_10934,N_10271);
nor U11606 (N_11606,N_10831,N_10274);
and U11607 (N_11607,N_10592,N_10847);
or U11608 (N_11608,N_10329,N_10904);
xnor U11609 (N_11609,N_10710,N_10991);
or U11610 (N_11610,N_10743,N_10860);
nor U11611 (N_11611,N_10774,N_10270);
and U11612 (N_11612,N_10090,N_10762);
and U11613 (N_11613,N_10404,N_10490);
nor U11614 (N_11614,N_10069,N_10040);
xnor U11615 (N_11615,N_10861,N_10271);
xnor U11616 (N_11616,N_10553,N_10053);
nand U11617 (N_11617,N_10646,N_10580);
or U11618 (N_11618,N_10730,N_10460);
xnor U11619 (N_11619,N_10999,N_10622);
xor U11620 (N_11620,N_10528,N_10676);
or U11621 (N_11621,N_10905,N_10408);
nand U11622 (N_11622,N_10900,N_10252);
nor U11623 (N_11623,N_10246,N_10836);
and U11624 (N_11624,N_10076,N_10565);
or U11625 (N_11625,N_10334,N_10818);
xor U11626 (N_11626,N_10154,N_10346);
xor U11627 (N_11627,N_10470,N_10716);
nor U11628 (N_11628,N_10609,N_10112);
nand U11629 (N_11629,N_10748,N_10219);
xnor U11630 (N_11630,N_10359,N_10473);
or U11631 (N_11631,N_10740,N_10153);
and U11632 (N_11632,N_10478,N_10824);
or U11633 (N_11633,N_10524,N_10242);
or U11634 (N_11634,N_10803,N_10999);
or U11635 (N_11635,N_10852,N_10946);
nor U11636 (N_11636,N_10605,N_10829);
and U11637 (N_11637,N_10176,N_10503);
or U11638 (N_11638,N_10600,N_10312);
and U11639 (N_11639,N_10849,N_10109);
nor U11640 (N_11640,N_10636,N_10447);
xor U11641 (N_11641,N_10228,N_10771);
nand U11642 (N_11642,N_10099,N_10232);
and U11643 (N_11643,N_10272,N_10510);
and U11644 (N_11644,N_10521,N_10091);
or U11645 (N_11645,N_10412,N_10038);
or U11646 (N_11646,N_10144,N_10180);
and U11647 (N_11647,N_10560,N_10043);
and U11648 (N_11648,N_10920,N_10424);
and U11649 (N_11649,N_10213,N_10697);
nor U11650 (N_11650,N_10246,N_10734);
nor U11651 (N_11651,N_10658,N_10441);
and U11652 (N_11652,N_10734,N_10618);
and U11653 (N_11653,N_10604,N_10366);
nor U11654 (N_11654,N_10900,N_10697);
and U11655 (N_11655,N_10010,N_10287);
xnor U11656 (N_11656,N_10373,N_10197);
xnor U11657 (N_11657,N_10676,N_10536);
xor U11658 (N_11658,N_10273,N_10683);
nor U11659 (N_11659,N_10733,N_10682);
xor U11660 (N_11660,N_10430,N_10605);
and U11661 (N_11661,N_10290,N_10117);
or U11662 (N_11662,N_10248,N_10444);
xnor U11663 (N_11663,N_10055,N_10001);
and U11664 (N_11664,N_10847,N_10575);
and U11665 (N_11665,N_10886,N_10967);
nor U11666 (N_11666,N_10570,N_10999);
or U11667 (N_11667,N_10025,N_10564);
nor U11668 (N_11668,N_10560,N_10212);
and U11669 (N_11669,N_10285,N_10263);
xor U11670 (N_11670,N_10084,N_10017);
nor U11671 (N_11671,N_10540,N_10375);
nand U11672 (N_11672,N_10713,N_10518);
nor U11673 (N_11673,N_10129,N_10058);
or U11674 (N_11674,N_10034,N_10118);
nor U11675 (N_11675,N_10152,N_10758);
and U11676 (N_11676,N_10728,N_10719);
nand U11677 (N_11677,N_10132,N_10703);
xnor U11678 (N_11678,N_10379,N_10572);
and U11679 (N_11679,N_10121,N_10157);
nand U11680 (N_11680,N_10739,N_10675);
nand U11681 (N_11681,N_10485,N_10710);
xor U11682 (N_11682,N_10756,N_10220);
nand U11683 (N_11683,N_10652,N_10161);
nor U11684 (N_11684,N_10740,N_10106);
nand U11685 (N_11685,N_10887,N_10716);
and U11686 (N_11686,N_10207,N_10173);
or U11687 (N_11687,N_10197,N_10060);
nand U11688 (N_11688,N_10857,N_10133);
nand U11689 (N_11689,N_10793,N_10224);
and U11690 (N_11690,N_10018,N_10113);
nor U11691 (N_11691,N_10038,N_10992);
or U11692 (N_11692,N_10659,N_10296);
nand U11693 (N_11693,N_10779,N_10095);
xor U11694 (N_11694,N_10612,N_10282);
xnor U11695 (N_11695,N_10125,N_10420);
or U11696 (N_11696,N_10952,N_10156);
or U11697 (N_11697,N_10815,N_10421);
nor U11698 (N_11698,N_10878,N_10943);
and U11699 (N_11699,N_10497,N_10119);
nand U11700 (N_11700,N_10612,N_10784);
nand U11701 (N_11701,N_10113,N_10725);
nor U11702 (N_11702,N_10005,N_10979);
and U11703 (N_11703,N_10887,N_10731);
xor U11704 (N_11704,N_10623,N_10153);
nand U11705 (N_11705,N_10868,N_10112);
xnor U11706 (N_11706,N_10189,N_10570);
and U11707 (N_11707,N_10617,N_10077);
nor U11708 (N_11708,N_10587,N_10037);
nand U11709 (N_11709,N_10584,N_10648);
or U11710 (N_11710,N_10060,N_10906);
nor U11711 (N_11711,N_10516,N_10211);
nand U11712 (N_11712,N_10474,N_10009);
or U11713 (N_11713,N_10698,N_10091);
and U11714 (N_11714,N_10627,N_10086);
or U11715 (N_11715,N_10455,N_10619);
or U11716 (N_11716,N_10468,N_10738);
xnor U11717 (N_11717,N_10047,N_10145);
nor U11718 (N_11718,N_10397,N_10069);
or U11719 (N_11719,N_10000,N_10688);
nand U11720 (N_11720,N_10168,N_10373);
or U11721 (N_11721,N_10777,N_10533);
nand U11722 (N_11722,N_10814,N_10136);
and U11723 (N_11723,N_10715,N_10051);
nand U11724 (N_11724,N_10840,N_10027);
xnor U11725 (N_11725,N_10143,N_10750);
and U11726 (N_11726,N_10232,N_10703);
and U11727 (N_11727,N_10556,N_10733);
nor U11728 (N_11728,N_10548,N_10956);
xor U11729 (N_11729,N_10203,N_10690);
and U11730 (N_11730,N_10683,N_10604);
and U11731 (N_11731,N_10842,N_10547);
nor U11732 (N_11732,N_10545,N_10980);
nand U11733 (N_11733,N_10693,N_10604);
xnor U11734 (N_11734,N_10349,N_10395);
and U11735 (N_11735,N_10005,N_10034);
or U11736 (N_11736,N_10696,N_10048);
and U11737 (N_11737,N_10527,N_10721);
and U11738 (N_11738,N_10511,N_10699);
nor U11739 (N_11739,N_10570,N_10677);
or U11740 (N_11740,N_10773,N_10789);
nand U11741 (N_11741,N_10825,N_10728);
and U11742 (N_11742,N_10465,N_10582);
and U11743 (N_11743,N_10888,N_10362);
and U11744 (N_11744,N_10849,N_10720);
nand U11745 (N_11745,N_10154,N_10903);
xnor U11746 (N_11746,N_10271,N_10577);
nor U11747 (N_11747,N_10194,N_10395);
and U11748 (N_11748,N_10391,N_10702);
and U11749 (N_11749,N_10332,N_10323);
xnor U11750 (N_11750,N_10854,N_10303);
nand U11751 (N_11751,N_10319,N_10992);
and U11752 (N_11752,N_10983,N_10608);
or U11753 (N_11753,N_10934,N_10898);
nand U11754 (N_11754,N_10746,N_10594);
and U11755 (N_11755,N_10402,N_10166);
nand U11756 (N_11756,N_10266,N_10613);
xor U11757 (N_11757,N_10050,N_10115);
xor U11758 (N_11758,N_10139,N_10411);
nand U11759 (N_11759,N_10767,N_10593);
or U11760 (N_11760,N_10917,N_10946);
and U11761 (N_11761,N_10535,N_10989);
xnor U11762 (N_11762,N_10328,N_10568);
and U11763 (N_11763,N_10991,N_10469);
and U11764 (N_11764,N_10895,N_10555);
xnor U11765 (N_11765,N_10561,N_10781);
or U11766 (N_11766,N_10652,N_10399);
nor U11767 (N_11767,N_10097,N_10728);
or U11768 (N_11768,N_10621,N_10151);
nor U11769 (N_11769,N_10853,N_10030);
or U11770 (N_11770,N_10025,N_10978);
xnor U11771 (N_11771,N_10269,N_10533);
nor U11772 (N_11772,N_10132,N_10608);
and U11773 (N_11773,N_10636,N_10944);
or U11774 (N_11774,N_10628,N_10414);
xnor U11775 (N_11775,N_10582,N_10462);
nor U11776 (N_11776,N_10077,N_10428);
or U11777 (N_11777,N_10951,N_10715);
and U11778 (N_11778,N_10255,N_10140);
nor U11779 (N_11779,N_10257,N_10839);
nand U11780 (N_11780,N_10063,N_10891);
and U11781 (N_11781,N_10052,N_10458);
and U11782 (N_11782,N_10405,N_10379);
and U11783 (N_11783,N_10617,N_10722);
xor U11784 (N_11784,N_10853,N_10492);
xnor U11785 (N_11785,N_10710,N_10423);
or U11786 (N_11786,N_10382,N_10426);
and U11787 (N_11787,N_10961,N_10861);
nand U11788 (N_11788,N_10163,N_10935);
or U11789 (N_11789,N_10584,N_10514);
nand U11790 (N_11790,N_10035,N_10093);
and U11791 (N_11791,N_10011,N_10325);
nor U11792 (N_11792,N_10664,N_10454);
and U11793 (N_11793,N_10897,N_10393);
nor U11794 (N_11794,N_10951,N_10164);
and U11795 (N_11795,N_10716,N_10896);
and U11796 (N_11796,N_10223,N_10338);
and U11797 (N_11797,N_10038,N_10457);
xor U11798 (N_11798,N_10094,N_10017);
nor U11799 (N_11799,N_10221,N_10539);
or U11800 (N_11800,N_10636,N_10858);
or U11801 (N_11801,N_10155,N_10437);
nor U11802 (N_11802,N_10786,N_10460);
xnor U11803 (N_11803,N_10197,N_10602);
nand U11804 (N_11804,N_10502,N_10601);
or U11805 (N_11805,N_10362,N_10864);
nand U11806 (N_11806,N_10573,N_10047);
or U11807 (N_11807,N_10180,N_10805);
xor U11808 (N_11808,N_10244,N_10986);
nor U11809 (N_11809,N_10412,N_10319);
nor U11810 (N_11810,N_10874,N_10847);
or U11811 (N_11811,N_10637,N_10570);
and U11812 (N_11812,N_10688,N_10300);
nor U11813 (N_11813,N_10351,N_10276);
and U11814 (N_11814,N_10510,N_10822);
xnor U11815 (N_11815,N_10921,N_10309);
or U11816 (N_11816,N_10820,N_10161);
nand U11817 (N_11817,N_10610,N_10142);
and U11818 (N_11818,N_10437,N_10610);
nor U11819 (N_11819,N_10609,N_10466);
nor U11820 (N_11820,N_10709,N_10493);
nor U11821 (N_11821,N_10147,N_10774);
nor U11822 (N_11822,N_10605,N_10055);
xnor U11823 (N_11823,N_10349,N_10293);
xor U11824 (N_11824,N_10633,N_10522);
or U11825 (N_11825,N_10421,N_10321);
nor U11826 (N_11826,N_10355,N_10488);
nor U11827 (N_11827,N_10375,N_10733);
or U11828 (N_11828,N_10985,N_10240);
nand U11829 (N_11829,N_10653,N_10261);
or U11830 (N_11830,N_10433,N_10246);
or U11831 (N_11831,N_10609,N_10304);
and U11832 (N_11832,N_10783,N_10859);
nor U11833 (N_11833,N_10774,N_10830);
nand U11834 (N_11834,N_10098,N_10787);
nor U11835 (N_11835,N_10813,N_10812);
nor U11836 (N_11836,N_10883,N_10462);
and U11837 (N_11837,N_10656,N_10945);
or U11838 (N_11838,N_10938,N_10374);
or U11839 (N_11839,N_10759,N_10924);
and U11840 (N_11840,N_10374,N_10934);
xnor U11841 (N_11841,N_10199,N_10293);
or U11842 (N_11842,N_10543,N_10294);
or U11843 (N_11843,N_10155,N_10432);
or U11844 (N_11844,N_10792,N_10523);
nand U11845 (N_11845,N_10903,N_10979);
nand U11846 (N_11846,N_10191,N_10294);
and U11847 (N_11847,N_10626,N_10591);
nor U11848 (N_11848,N_10331,N_10973);
nand U11849 (N_11849,N_10687,N_10906);
nor U11850 (N_11850,N_10270,N_10110);
or U11851 (N_11851,N_10909,N_10341);
xor U11852 (N_11852,N_10326,N_10504);
and U11853 (N_11853,N_10121,N_10259);
and U11854 (N_11854,N_10662,N_10316);
xor U11855 (N_11855,N_10601,N_10309);
and U11856 (N_11856,N_10689,N_10626);
xor U11857 (N_11857,N_10030,N_10785);
or U11858 (N_11858,N_10450,N_10215);
nor U11859 (N_11859,N_10660,N_10258);
nor U11860 (N_11860,N_10393,N_10180);
or U11861 (N_11861,N_10483,N_10065);
and U11862 (N_11862,N_10355,N_10589);
or U11863 (N_11863,N_10240,N_10026);
xnor U11864 (N_11864,N_10831,N_10390);
nand U11865 (N_11865,N_10414,N_10885);
nand U11866 (N_11866,N_10839,N_10522);
or U11867 (N_11867,N_10075,N_10288);
and U11868 (N_11868,N_10134,N_10056);
xnor U11869 (N_11869,N_10072,N_10850);
xnor U11870 (N_11870,N_10845,N_10485);
nand U11871 (N_11871,N_10942,N_10404);
or U11872 (N_11872,N_10630,N_10024);
nor U11873 (N_11873,N_10404,N_10153);
xor U11874 (N_11874,N_10379,N_10987);
nor U11875 (N_11875,N_10455,N_10356);
nor U11876 (N_11876,N_10689,N_10255);
and U11877 (N_11877,N_10395,N_10834);
nand U11878 (N_11878,N_10906,N_10199);
nand U11879 (N_11879,N_10522,N_10279);
or U11880 (N_11880,N_10520,N_10623);
nor U11881 (N_11881,N_10397,N_10688);
nor U11882 (N_11882,N_10938,N_10886);
xnor U11883 (N_11883,N_10057,N_10890);
nor U11884 (N_11884,N_10154,N_10512);
or U11885 (N_11885,N_10530,N_10864);
xor U11886 (N_11886,N_10416,N_10404);
or U11887 (N_11887,N_10860,N_10221);
and U11888 (N_11888,N_10754,N_10992);
and U11889 (N_11889,N_10368,N_10736);
xor U11890 (N_11890,N_10167,N_10864);
xnor U11891 (N_11891,N_10162,N_10499);
or U11892 (N_11892,N_10542,N_10527);
nand U11893 (N_11893,N_10115,N_10768);
nor U11894 (N_11894,N_10617,N_10320);
nand U11895 (N_11895,N_10108,N_10525);
and U11896 (N_11896,N_10120,N_10333);
or U11897 (N_11897,N_10434,N_10810);
xnor U11898 (N_11898,N_10112,N_10098);
xor U11899 (N_11899,N_10236,N_10153);
xnor U11900 (N_11900,N_10176,N_10779);
or U11901 (N_11901,N_10375,N_10176);
nor U11902 (N_11902,N_10076,N_10248);
xor U11903 (N_11903,N_10337,N_10815);
nand U11904 (N_11904,N_10935,N_10803);
xor U11905 (N_11905,N_10854,N_10858);
nand U11906 (N_11906,N_10401,N_10141);
xor U11907 (N_11907,N_10949,N_10230);
xor U11908 (N_11908,N_10731,N_10575);
xnor U11909 (N_11909,N_10177,N_10372);
nand U11910 (N_11910,N_10889,N_10479);
xor U11911 (N_11911,N_10972,N_10381);
nand U11912 (N_11912,N_10703,N_10903);
xnor U11913 (N_11913,N_10643,N_10910);
nand U11914 (N_11914,N_10623,N_10311);
xor U11915 (N_11915,N_10169,N_10746);
xor U11916 (N_11916,N_10465,N_10269);
or U11917 (N_11917,N_10042,N_10661);
or U11918 (N_11918,N_10715,N_10036);
or U11919 (N_11919,N_10669,N_10222);
nor U11920 (N_11920,N_10407,N_10576);
nand U11921 (N_11921,N_10979,N_10439);
and U11922 (N_11922,N_10257,N_10488);
nand U11923 (N_11923,N_10408,N_10516);
xor U11924 (N_11924,N_10747,N_10241);
and U11925 (N_11925,N_10093,N_10268);
and U11926 (N_11926,N_10086,N_10429);
nand U11927 (N_11927,N_10967,N_10922);
or U11928 (N_11928,N_10592,N_10000);
xor U11929 (N_11929,N_10113,N_10965);
or U11930 (N_11930,N_10815,N_10559);
nand U11931 (N_11931,N_10653,N_10052);
nand U11932 (N_11932,N_10158,N_10376);
xnor U11933 (N_11933,N_10617,N_10224);
or U11934 (N_11934,N_10464,N_10824);
and U11935 (N_11935,N_10812,N_10336);
and U11936 (N_11936,N_10527,N_10671);
and U11937 (N_11937,N_10807,N_10800);
nor U11938 (N_11938,N_10161,N_10343);
nor U11939 (N_11939,N_10150,N_10851);
and U11940 (N_11940,N_10170,N_10935);
nor U11941 (N_11941,N_10182,N_10111);
and U11942 (N_11942,N_10605,N_10849);
nand U11943 (N_11943,N_10503,N_10777);
or U11944 (N_11944,N_10701,N_10892);
nand U11945 (N_11945,N_10525,N_10222);
or U11946 (N_11946,N_10231,N_10457);
xor U11947 (N_11947,N_10659,N_10448);
or U11948 (N_11948,N_10197,N_10959);
and U11949 (N_11949,N_10443,N_10000);
or U11950 (N_11950,N_10910,N_10548);
xor U11951 (N_11951,N_10465,N_10505);
or U11952 (N_11952,N_10568,N_10685);
and U11953 (N_11953,N_10117,N_10808);
or U11954 (N_11954,N_10761,N_10996);
or U11955 (N_11955,N_10956,N_10015);
nand U11956 (N_11956,N_10716,N_10355);
xor U11957 (N_11957,N_10683,N_10625);
nor U11958 (N_11958,N_10401,N_10333);
xor U11959 (N_11959,N_10432,N_10922);
nand U11960 (N_11960,N_10254,N_10994);
or U11961 (N_11961,N_10755,N_10187);
nor U11962 (N_11962,N_10994,N_10602);
or U11963 (N_11963,N_10749,N_10914);
nand U11964 (N_11964,N_10201,N_10465);
or U11965 (N_11965,N_10713,N_10488);
or U11966 (N_11966,N_10456,N_10834);
xnor U11967 (N_11967,N_10228,N_10270);
and U11968 (N_11968,N_10099,N_10143);
xnor U11969 (N_11969,N_10218,N_10402);
or U11970 (N_11970,N_10486,N_10562);
or U11971 (N_11971,N_10470,N_10968);
and U11972 (N_11972,N_10626,N_10261);
nor U11973 (N_11973,N_10336,N_10982);
nor U11974 (N_11974,N_10205,N_10845);
nor U11975 (N_11975,N_10077,N_10533);
nor U11976 (N_11976,N_10010,N_10624);
nor U11977 (N_11977,N_10350,N_10237);
or U11978 (N_11978,N_10029,N_10224);
xnor U11979 (N_11979,N_10694,N_10448);
nand U11980 (N_11980,N_10376,N_10100);
or U11981 (N_11981,N_10586,N_10550);
and U11982 (N_11982,N_10959,N_10600);
and U11983 (N_11983,N_10169,N_10219);
xnor U11984 (N_11984,N_10964,N_10766);
and U11985 (N_11985,N_10209,N_10455);
nand U11986 (N_11986,N_10184,N_10294);
or U11987 (N_11987,N_10748,N_10650);
nor U11988 (N_11988,N_10773,N_10397);
nor U11989 (N_11989,N_10357,N_10580);
xnor U11990 (N_11990,N_10793,N_10114);
xnor U11991 (N_11991,N_10571,N_10189);
or U11992 (N_11992,N_10094,N_10340);
nor U11993 (N_11993,N_10949,N_10381);
xor U11994 (N_11994,N_10895,N_10253);
and U11995 (N_11995,N_10220,N_10673);
or U11996 (N_11996,N_10312,N_10659);
xor U11997 (N_11997,N_10797,N_10637);
and U11998 (N_11998,N_10873,N_10134);
or U11999 (N_11999,N_10667,N_10638);
and U12000 (N_12000,N_11330,N_11897);
xor U12001 (N_12001,N_11121,N_11580);
or U12002 (N_12002,N_11781,N_11606);
nand U12003 (N_12003,N_11226,N_11807);
nand U12004 (N_12004,N_11672,N_11675);
and U12005 (N_12005,N_11084,N_11274);
xor U12006 (N_12006,N_11837,N_11645);
nand U12007 (N_12007,N_11385,N_11736);
or U12008 (N_12008,N_11586,N_11549);
and U12009 (N_12009,N_11521,N_11783);
nand U12010 (N_12010,N_11924,N_11141);
nor U12011 (N_12011,N_11550,N_11304);
or U12012 (N_12012,N_11903,N_11231);
and U12013 (N_12013,N_11546,N_11523);
or U12014 (N_12014,N_11875,N_11701);
xor U12015 (N_12015,N_11557,N_11269);
nor U12016 (N_12016,N_11006,N_11631);
xnor U12017 (N_12017,N_11025,N_11734);
nand U12018 (N_12018,N_11848,N_11628);
xor U12019 (N_12019,N_11189,N_11356);
and U12020 (N_12020,N_11772,N_11241);
nor U12021 (N_12021,N_11756,N_11745);
nor U12022 (N_12022,N_11174,N_11265);
nand U12023 (N_12023,N_11284,N_11237);
xnor U12024 (N_12024,N_11207,N_11618);
and U12025 (N_12025,N_11162,N_11596);
or U12026 (N_12026,N_11011,N_11097);
or U12027 (N_12027,N_11238,N_11257);
or U12028 (N_12028,N_11967,N_11040);
and U12029 (N_12029,N_11020,N_11595);
or U12030 (N_12030,N_11272,N_11678);
and U12031 (N_12031,N_11735,N_11761);
and U12032 (N_12032,N_11451,N_11352);
and U12033 (N_12033,N_11372,N_11590);
nor U12034 (N_12034,N_11388,N_11473);
nand U12035 (N_12035,N_11988,N_11273);
nand U12036 (N_12036,N_11544,N_11540);
and U12037 (N_12037,N_11572,N_11996);
nor U12038 (N_12038,N_11424,N_11986);
nor U12039 (N_12039,N_11318,N_11125);
or U12040 (N_12040,N_11947,N_11299);
nor U12041 (N_12041,N_11686,N_11737);
nor U12042 (N_12042,N_11093,N_11294);
or U12043 (N_12043,N_11882,N_11629);
and U12044 (N_12044,N_11072,N_11743);
nor U12045 (N_12045,N_11437,N_11157);
or U12046 (N_12046,N_11357,N_11759);
nor U12047 (N_12047,N_11133,N_11476);
xnor U12048 (N_12048,N_11945,N_11514);
nand U12049 (N_12049,N_11055,N_11096);
nor U12050 (N_12050,N_11484,N_11012);
xor U12051 (N_12051,N_11977,N_11377);
and U12052 (N_12052,N_11927,N_11206);
or U12053 (N_12053,N_11828,N_11479);
and U12054 (N_12054,N_11496,N_11060);
nand U12055 (N_12055,N_11399,N_11229);
or U12056 (N_12056,N_11443,N_11113);
xor U12057 (N_12057,N_11918,N_11029);
xnor U12058 (N_12058,N_11128,N_11191);
xor U12059 (N_12059,N_11248,N_11487);
xnor U12060 (N_12060,N_11673,N_11884);
or U12061 (N_12061,N_11095,N_11916);
nand U12062 (N_12062,N_11511,N_11288);
nor U12063 (N_12063,N_11285,N_11449);
or U12064 (N_12064,N_11537,N_11512);
xnor U12065 (N_12065,N_11638,N_11341);
and U12066 (N_12066,N_11909,N_11723);
or U12067 (N_12067,N_11379,N_11270);
nand U12068 (N_12068,N_11682,N_11863);
and U12069 (N_12069,N_11069,N_11480);
xor U12070 (N_12070,N_11622,N_11957);
nand U12071 (N_12071,N_11731,N_11861);
or U12072 (N_12072,N_11180,N_11632);
xnor U12073 (N_12073,N_11371,N_11738);
and U12074 (N_12074,N_11887,N_11670);
and U12075 (N_12075,N_11669,N_11401);
nor U12076 (N_12076,N_11519,N_11109);
and U12077 (N_12077,N_11690,N_11732);
nand U12078 (N_12078,N_11555,N_11981);
nor U12079 (N_12079,N_11502,N_11446);
nor U12080 (N_12080,N_11130,N_11915);
nor U12081 (N_12081,N_11079,N_11845);
xnor U12082 (N_12082,N_11439,N_11931);
nor U12083 (N_12083,N_11951,N_11963);
or U12084 (N_12084,N_11472,N_11825);
and U12085 (N_12085,N_11431,N_11419);
xnor U12086 (N_12086,N_11777,N_11253);
xnor U12087 (N_12087,N_11317,N_11345);
or U12088 (N_12088,N_11001,N_11785);
nand U12089 (N_12089,N_11425,N_11007);
or U12090 (N_12090,N_11637,N_11906);
xor U12091 (N_12091,N_11538,N_11799);
or U12092 (N_12092,N_11244,N_11869);
nor U12093 (N_12093,N_11528,N_11470);
nor U12094 (N_12094,N_11225,N_11192);
and U12095 (N_12095,N_11074,N_11382);
nor U12096 (N_12096,N_11878,N_11374);
nand U12097 (N_12097,N_11111,N_11862);
and U12098 (N_12098,N_11491,N_11810);
nor U12099 (N_12099,N_11378,N_11668);
or U12100 (N_12100,N_11088,N_11859);
and U12101 (N_12101,N_11031,N_11393);
nand U12102 (N_12102,N_11752,N_11305);
and U12103 (N_12103,N_11936,N_11683);
and U12104 (N_12104,N_11126,N_11033);
nor U12105 (N_12105,N_11264,N_11455);
nor U12106 (N_12106,N_11856,N_11324);
xnor U12107 (N_12107,N_11803,N_11018);
nand U12108 (N_12108,N_11381,N_11214);
xnor U12109 (N_12109,N_11008,N_11010);
xnor U12110 (N_12110,N_11651,N_11529);
nor U12111 (N_12111,N_11623,N_11197);
nor U12112 (N_12112,N_11826,N_11598);
xnor U12113 (N_12113,N_11384,N_11250);
nand U12114 (N_12114,N_11004,N_11921);
xor U12115 (N_12115,N_11879,N_11985);
or U12116 (N_12116,N_11445,N_11753);
or U12117 (N_12117,N_11594,N_11085);
or U12118 (N_12118,N_11051,N_11534);
nand U12119 (N_12119,N_11423,N_11775);
and U12120 (N_12120,N_11043,N_11708);
xnor U12121 (N_12121,N_11187,N_11657);
or U12122 (N_12122,N_11014,N_11760);
and U12123 (N_12123,N_11448,N_11246);
and U12124 (N_12124,N_11642,N_11015);
xnor U12125 (N_12125,N_11561,N_11896);
or U12126 (N_12126,N_11486,N_11411);
nor U12127 (N_12127,N_11210,N_11108);
nor U12128 (N_12128,N_11478,N_11418);
or U12129 (N_12129,N_11205,N_11173);
or U12130 (N_12130,N_11677,N_11076);
nor U12131 (N_12131,N_11275,N_11368);
nand U12132 (N_12132,N_11913,N_11216);
nand U12133 (N_12133,N_11721,N_11497);
xor U12134 (N_12134,N_11578,N_11019);
nand U12135 (N_12135,N_11426,N_11765);
xor U12136 (N_12136,N_11755,N_11901);
xnor U12137 (N_12137,N_11297,N_11888);
nand U12138 (N_12138,N_11520,N_11220);
and U12139 (N_12139,N_11119,N_11083);
or U12140 (N_12140,N_11366,N_11005);
and U12141 (N_12141,N_11407,N_11616);
nand U12142 (N_12142,N_11905,N_11842);
nor U12143 (N_12143,N_11027,N_11868);
xor U12144 (N_12144,N_11349,N_11493);
xnor U12145 (N_12145,N_11791,N_11181);
nor U12146 (N_12146,N_11978,N_11792);
xnor U12147 (N_12147,N_11639,N_11347);
xor U12148 (N_12148,N_11458,N_11958);
and U12149 (N_12149,N_11087,N_11965);
nor U12150 (N_12150,N_11337,N_11498);
nor U12151 (N_12151,N_11416,N_11873);
or U12152 (N_12152,N_11808,N_11148);
and U12153 (N_12153,N_11917,N_11287);
xor U12154 (N_12154,N_11415,N_11459);
or U12155 (N_12155,N_11138,N_11147);
or U12156 (N_12156,N_11300,N_11260);
xnor U12157 (N_12157,N_11160,N_11864);
or U12158 (N_12158,N_11902,N_11698);
and U12159 (N_12159,N_11073,N_11070);
nand U12160 (N_12160,N_11744,N_11621);
nand U12161 (N_12161,N_11364,N_11268);
nand U12162 (N_12162,N_11570,N_11145);
nand U12163 (N_12163,N_11465,N_11505);
xor U12164 (N_12164,N_11463,N_11894);
and U12165 (N_12165,N_11794,N_11970);
xor U12166 (N_12166,N_11363,N_11102);
xnor U12167 (N_12167,N_11346,N_11234);
nor U12168 (N_12168,N_11199,N_11146);
and U12169 (N_12169,N_11195,N_11955);
nor U12170 (N_12170,N_11942,N_11624);
or U12171 (N_12171,N_11186,N_11649);
nor U12172 (N_12172,N_11310,N_11222);
and U12173 (N_12173,N_11203,N_11485);
nand U12174 (N_12174,N_11860,N_11560);
xor U12175 (N_12175,N_11768,N_11276);
xnor U12176 (N_12176,N_11249,N_11874);
nand U12177 (N_12177,N_11541,N_11440);
or U12178 (N_12178,N_11697,N_11802);
nor U12179 (N_12179,N_11608,N_11912);
nor U12180 (N_12180,N_11353,N_11311);
or U12181 (N_12181,N_11793,N_11442);
or U12182 (N_12182,N_11904,N_11836);
or U12183 (N_12183,N_11840,N_11571);
nand U12184 (N_12184,N_11948,N_11436);
xor U12185 (N_12185,N_11713,N_11240);
nand U12186 (N_12186,N_11575,N_11565);
nand U12187 (N_12187,N_11277,N_11468);
nor U12188 (N_12188,N_11714,N_11507);
nor U12189 (N_12189,N_11361,N_11987);
xnor U12190 (N_12190,N_11979,N_11919);
or U12191 (N_12191,N_11644,N_11002);
nor U12192 (N_12192,N_11815,N_11428);
or U12193 (N_12193,N_11030,N_11259);
nor U12194 (N_12194,N_11042,N_11930);
xnor U12195 (N_12195,N_11376,N_11597);
and U12196 (N_12196,N_11348,N_11143);
and U12197 (N_12197,N_11167,N_11123);
nand U12198 (N_12198,N_11438,N_11267);
nor U12199 (N_12199,N_11427,N_11078);
nor U12200 (N_12200,N_11188,N_11818);
nor U12201 (N_12201,N_11742,N_11747);
nand U12202 (N_12202,N_11266,N_11552);
and U12203 (N_12203,N_11821,N_11716);
xnor U12204 (N_12204,N_11643,N_11215);
or U12205 (N_12205,N_11086,N_11581);
xor U12206 (N_12206,N_11466,N_11634);
and U12207 (N_12207,N_11059,N_11679);
and U12208 (N_12208,N_11464,N_11920);
nor U12209 (N_12209,N_11066,N_11196);
xor U12210 (N_12210,N_11281,N_11057);
nand U12211 (N_12211,N_11016,N_11976);
and U12212 (N_12212,N_11530,N_11140);
nor U12213 (N_12213,N_11757,N_11671);
or U12214 (N_12214,N_11101,N_11218);
xor U12215 (N_12215,N_11230,N_11235);
nand U12216 (N_12216,N_11525,N_11023);
xor U12217 (N_12217,N_11889,N_11787);
nor U12218 (N_12218,N_11691,N_11129);
xor U12219 (N_12219,N_11080,N_11727);
and U12220 (N_12220,N_11647,N_11939);
xor U12221 (N_12221,N_11991,N_11726);
xnor U12222 (N_12222,N_11204,N_11386);
or U12223 (N_12223,N_11308,N_11252);
nor U12224 (N_12224,N_11243,N_11392);
xor U12225 (N_12225,N_11302,N_11327);
nand U12226 (N_12226,N_11653,N_11200);
xor U12227 (N_12227,N_11612,N_11805);
nand U12228 (N_12228,N_11636,N_11441);
and U12229 (N_12229,N_11796,N_11454);
nor U12230 (N_12230,N_11704,N_11801);
nand U12231 (N_12231,N_11433,N_11763);
and U12232 (N_12232,N_11773,N_11403);
nand U12233 (N_12233,N_11599,N_11469);
or U12234 (N_12234,N_11829,N_11137);
nor U12235 (N_12235,N_11247,N_11539);
xor U12236 (N_12236,N_11488,N_11058);
nor U12237 (N_12237,N_11293,N_11870);
nor U12238 (N_12238,N_11556,N_11283);
nor U12239 (N_12239,N_11256,N_11000);
nand U12240 (N_12240,N_11573,N_11165);
xor U12241 (N_12241,N_11475,N_11702);
nand U12242 (N_12242,N_11971,N_11279);
or U12243 (N_12243,N_11190,N_11664);
xor U12244 (N_12244,N_11232,N_11547);
or U12245 (N_12245,N_11417,N_11254);
nand U12246 (N_12246,N_11506,N_11494);
xor U12247 (N_12247,N_11367,N_11696);
nor U12248 (N_12248,N_11895,N_11532);
nand U12249 (N_12249,N_11591,N_11035);
nand U12250 (N_12250,N_11926,N_11886);
or U12251 (N_12251,N_11658,N_11340);
xnor U12252 (N_12252,N_11315,N_11408);
and U12253 (N_12253,N_11003,N_11115);
and U12254 (N_12254,N_11322,N_11554);
nor U12255 (N_12255,N_11858,N_11666);
or U12256 (N_12256,N_11922,N_11885);
nand U12257 (N_12257,N_11767,N_11960);
and U12258 (N_12258,N_11307,N_11798);
xor U12259 (N_12259,N_11333,N_11700);
xnor U12260 (N_12260,N_11460,N_11389);
nand U12261 (N_12261,N_11261,N_11396);
and U12262 (N_12262,N_11620,N_11749);
or U12263 (N_12263,N_11820,N_11390);
and U12264 (N_12264,N_11046,N_11219);
and U12265 (N_12265,N_11258,N_11208);
and U12266 (N_12266,N_11048,N_11457);
xor U12267 (N_12267,N_11579,N_11797);
xor U12268 (N_12268,N_11950,N_11944);
and U12269 (N_12269,N_11626,N_11871);
nor U12270 (N_12270,N_11569,N_11663);
and U12271 (N_12271,N_11091,N_11562);
nand U12272 (N_12272,N_11712,N_11962);
and U12273 (N_12273,N_11790,N_11321);
xnor U12274 (N_12274,N_11335,N_11127);
nand U12275 (N_12275,N_11037,N_11405);
nand U12276 (N_12276,N_11120,N_11660);
nand U12277 (N_12277,N_11420,N_11412);
and U12278 (N_12278,N_11617,N_11398);
nor U12279 (N_12279,N_11524,N_11312);
xor U12280 (N_12280,N_11509,N_11159);
xor U12281 (N_12281,N_11400,N_11911);
xnor U12282 (N_12282,N_11526,N_11343);
nor U12283 (N_12283,N_11176,N_11722);
nor U12284 (N_12284,N_11536,N_11516);
nor U12285 (N_12285,N_11375,N_11172);
nand U12286 (N_12286,N_11194,N_11394);
and U12287 (N_12287,N_11688,N_11584);
nor U12288 (N_12288,N_11313,N_11762);
nand U12289 (N_12289,N_11515,N_11202);
nand U12290 (N_12290,N_11314,N_11134);
nor U12291 (N_12291,N_11699,N_11245);
or U12292 (N_12292,N_11964,N_11329);
nand U12293 (N_12293,N_11680,N_11482);
and U12294 (N_12294,N_11703,N_11142);
nand U12295 (N_12295,N_11421,N_11332);
nand U12296 (N_12296,N_11136,N_11309);
nand U12297 (N_12297,N_11844,N_11490);
or U12298 (N_12298,N_11568,N_11492);
xor U12299 (N_12299,N_11891,N_11992);
nor U12300 (N_12300,N_11456,N_11228);
and U12301 (N_12301,N_11689,N_11508);
xor U12302 (N_12302,N_11839,N_11583);
or U12303 (N_12303,N_11429,N_11344);
xor U12304 (N_12304,N_11720,N_11851);
or U12305 (N_12305,N_11161,N_11943);
nand U12306 (N_12306,N_11154,N_11641);
and U12307 (N_12307,N_11907,N_11306);
and U12308 (N_12308,N_11531,N_11974);
and U12309 (N_12309,N_11748,N_11956);
or U12310 (N_12310,N_11914,N_11602);
nand U12311 (N_12311,N_11823,N_11667);
nor U12312 (N_12312,N_11064,N_11809);
and U12313 (N_12313,N_11153,N_11212);
or U12314 (N_12314,N_11843,N_11582);
or U12315 (N_12315,N_11477,N_11118);
and U12316 (N_12316,N_11510,N_11892);
xor U12317 (N_12317,N_11788,N_11328);
nor U12318 (N_12318,N_11106,N_11830);
and U12319 (N_12319,N_11567,N_11370);
xnor U12320 (N_12320,N_11937,N_11406);
and U12321 (N_12321,N_11946,N_11614);
or U12322 (N_12322,N_11593,N_11959);
xor U12323 (N_12323,N_11577,N_11184);
nor U12324 (N_12324,N_11741,N_11941);
or U12325 (N_12325,N_11576,N_11932);
nor U12326 (N_12326,N_11183,N_11961);
nand U12327 (N_12327,N_11404,N_11233);
nor U12328 (N_12328,N_11032,N_11350);
nor U12329 (N_12329,N_11925,N_11847);
and U12330 (N_12330,N_11075,N_11171);
xnor U12331 (N_12331,N_11211,N_11255);
or U12332 (N_12332,N_11185,N_11613);
xnor U12333 (N_12333,N_11359,N_11017);
nor U12334 (N_12334,N_11351,N_11301);
or U12335 (N_12335,N_11592,N_11893);
or U12336 (N_12336,N_11656,N_11898);
nand U12337 (N_12337,N_11718,N_11039);
xnor U12338 (N_12338,N_11298,N_11103);
nor U12339 (N_12339,N_11050,N_11542);
or U12340 (N_12340,N_11513,N_11295);
xnor U12341 (N_12341,N_11325,N_11601);
and U12342 (N_12342,N_11044,N_11813);
xor U12343 (N_12343,N_11380,N_11989);
nor U12344 (N_12344,N_11504,N_11650);
xor U12345 (N_12345,N_11227,N_11563);
or U12346 (N_12346,N_11966,N_11661);
nor U12347 (N_12347,N_11841,N_11414);
nand U12348 (N_12348,N_11342,N_11600);
and U12349 (N_12349,N_11646,N_11444);
nor U12350 (N_12350,N_11630,N_11131);
or U12351 (N_12351,N_11107,N_11164);
or U12352 (N_12352,N_11705,N_11814);
nor U12353 (N_12353,N_11263,N_11725);
nor U12354 (N_12354,N_11779,N_11290);
nor U12355 (N_12355,N_11495,N_11972);
or U12356 (N_12356,N_11435,N_11984);
nand U12357 (N_12357,N_11338,N_11709);
and U12358 (N_12358,N_11999,N_11063);
nor U12359 (N_12359,N_11013,N_11707);
nor U12360 (N_12360,N_11053,N_11135);
or U12361 (N_12361,N_11778,N_11271);
or U12362 (N_12362,N_11122,N_11627);
nand U12363 (N_12363,N_11089,N_11693);
xor U12364 (N_12364,N_11117,N_11223);
xor U12365 (N_12365,N_11280,N_11872);
xor U12366 (N_12366,N_11432,N_11834);
nand U12367 (N_12367,N_11890,N_11316);
nor U12368 (N_12368,N_11038,N_11804);
nor U12369 (N_12369,N_11640,N_11662);
xnor U12370 (N_12370,N_11832,N_11750);
or U12371 (N_12371,N_11110,N_11934);
xor U12372 (N_12372,N_11940,N_11036);
nand U12373 (N_12373,N_11949,N_11116);
nand U12374 (N_12374,N_11710,N_11262);
nor U12375 (N_12375,N_11564,N_11099);
or U12376 (N_12376,N_11846,N_11633);
and U12377 (N_12377,N_11533,N_11764);
or U12378 (N_12378,N_11052,N_11822);
nand U12379 (N_12379,N_11719,N_11499);
and U12380 (N_12380,N_11758,N_11471);
nand U12381 (N_12381,N_11067,N_11604);
and U12382 (N_12382,N_11610,N_11169);
nor U12383 (N_12383,N_11461,N_11151);
nand U12384 (N_12384,N_11094,N_11995);
nor U12385 (N_12385,N_11331,N_11838);
nand U12386 (N_12386,N_11553,N_11566);
and U12387 (N_12387,N_11409,N_11684);
nand U12388 (N_12388,N_11360,N_11251);
or U12389 (N_12389,N_11652,N_11865);
nand U12390 (N_12390,N_11855,N_11242);
nor U12391 (N_12391,N_11026,N_11733);
xor U12392 (N_12392,N_11817,N_11811);
or U12393 (N_12393,N_11397,N_11024);
nor U12394 (N_12394,N_11866,N_11453);
or U12395 (N_12395,N_11365,N_11062);
nor U12396 (N_12396,N_11434,N_11323);
and U12397 (N_12397,N_11224,N_11938);
nand U12398 (N_12398,N_11041,N_11201);
or U12399 (N_12399,N_11625,N_11383);
xor U12400 (N_12400,N_11447,N_11292);
nand U12401 (N_12401,N_11373,N_11462);
nand U12402 (N_12402,N_11588,N_11483);
xor U12403 (N_12403,N_11795,N_11835);
or U12404 (N_12404,N_11695,N_11800);
nand U12405 (N_12405,N_11022,N_11278);
and U12406 (N_12406,N_11980,N_11728);
and U12407 (N_12407,N_11993,N_11092);
nor U12408 (N_12408,N_11489,N_11994);
xnor U12409 (N_12409,N_11217,N_11786);
nand U12410 (N_12410,N_11150,N_11724);
and U12411 (N_12411,N_11090,N_11213);
xor U12412 (N_12412,N_11935,N_11694);
nand U12413 (N_12413,N_11236,N_11923);
xnor U12414 (N_12414,N_11422,N_11706);
xnor U12415 (N_12415,N_11819,N_11968);
or U12416 (N_12416,N_11973,N_11816);
and U12417 (N_12417,N_11149,N_11997);
nand U12418 (N_12418,N_11045,N_11193);
nor U12419 (N_12419,N_11009,N_11175);
or U12420 (N_12420,N_11827,N_11619);
nand U12421 (N_12421,N_11806,N_11876);
xnor U12422 (N_12422,N_11369,N_11170);
and U12423 (N_12423,N_11611,N_11158);
or U12424 (N_12424,N_11854,N_11481);
nor U12425 (N_12425,N_11098,N_11166);
or U12426 (N_12426,N_11715,N_11605);
nor U12427 (N_12427,N_11774,N_11177);
or U12428 (N_12428,N_11603,N_11607);
or U12429 (N_12429,N_11574,N_11585);
and U12430 (N_12430,N_11900,N_11056);
nor U12431 (N_12431,N_11168,N_11336);
nor U12432 (N_12432,N_11648,N_11517);
nand U12433 (N_12433,N_11751,N_11518);
nor U12434 (N_12434,N_11112,N_11077);
or U12435 (N_12435,N_11152,N_11155);
xor U12436 (N_12436,N_11609,N_11771);
nor U12437 (N_12437,N_11929,N_11975);
and U12438 (N_12438,N_11877,N_11387);
nor U12439 (N_12439,N_11319,N_11355);
and U12440 (N_12440,N_11402,N_11139);
or U12441 (N_12441,N_11061,N_11548);
or U12442 (N_12442,N_11105,N_11784);
nor U12443 (N_12443,N_11543,N_11474);
nand U12444 (N_12444,N_11717,N_11687);
and U12445 (N_12445,N_11692,N_11410);
xnor U12446 (N_12446,N_11789,N_11021);
nand U12447 (N_12447,N_11391,N_11239);
nor U12448 (N_12448,N_11559,N_11221);
and U12449 (N_12449,N_11065,N_11339);
nand U12450 (N_12450,N_11730,N_11665);
or U12451 (N_12451,N_11047,N_11358);
nor U12452 (N_12452,N_11867,N_11908);
nor U12453 (N_12453,N_11114,N_11163);
xnor U12454 (N_12454,N_11769,N_11635);
nor U12455 (N_12455,N_11081,N_11654);
xnor U12456 (N_12456,N_11899,N_11551);
and U12457 (N_12457,N_11144,N_11776);
nor U12458 (N_12458,N_11982,N_11812);
nor U12459 (N_12459,N_11334,N_11739);
nand U12460 (N_12460,N_11969,N_11054);
nand U12461 (N_12461,N_11766,N_11729);
or U12462 (N_12462,N_11291,N_11853);
nor U12463 (N_12463,N_11034,N_11100);
nor U12464 (N_12464,N_11881,N_11082);
or U12465 (N_12465,N_11711,N_11326);
nand U12466 (N_12466,N_11587,N_11209);
xor U12467 (N_12467,N_11156,N_11452);
xor U12468 (N_12468,N_11296,N_11450);
and U12469 (N_12469,N_11354,N_11685);
nor U12470 (N_12470,N_11503,N_11849);
and U12471 (N_12471,N_11527,N_11754);
xnor U12472 (N_12472,N_11198,N_11413);
nand U12473 (N_12473,N_11467,N_11952);
and U12474 (N_12474,N_11362,N_11303);
and U12475 (N_12475,N_11833,N_11740);
xor U12476 (N_12476,N_11852,N_11071);
xor U12477 (N_12477,N_11179,N_11395);
or U12478 (N_12478,N_11857,N_11953);
and U12479 (N_12479,N_11558,N_11983);
xor U12480 (N_12480,N_11655,N_11928);
nor U12481 (N_12481,N_11178,N_11831);
nor U12482 (N_12482,N_11681,N_11883);
or U12483 (N_12483,N_11770,N_11132);
nor U12484 (N_12484,N_11954,N_11068);
nand U12485 (N_12485,N_11501,N_11289);
xor U12486 (N_12486,N_11676,N_11282);
or U12487 (N_12487,N_11500,N_11782);
or U12488 (N_12488,N_11780,N_11286);
xnor U12489 (N_12489,N_11049,N_11746);
nor U12490 (N_12490,N_11545,N_11430);
nor U12491 (N_12491,N_11910,N_11998);
and U12492 (N_12492,N_11104,N_11589);
xor U12493 (N_12493,N_11028,N_11824);
or U12494 (N_12494,N_11182,N_11933);
xor U12495 (N_12495,N_11615,N_11522);
nor U12496 (N_12496,N_11850,N_11124);
and U12497 (N_12497,N_11535,N_11659);
nor U12498 (N_12498,N_11674,N_11880);
or U12499 (N_12499,N_11320,N_11990);
xor U12500 (N_12500,N_11246,N_11523);
xnor U12501 (N_12501,N_11082,N_11227);
and U12502 (N_12502,N_11925,N_11186);
or U12503 (N_12503,N_11262,N_11828);
and U12504 (N_12504,N_11256,N_11941);
and U12505 (N_12505,N_11723,N_11077);
nor U12506 (N_12506,N_11207,N_11442);
and U12507 (N_12507,N_11503,N_11876);
or U12508 (N_12508,N_11044,N_11613);
and U12509 (N_12509,N_11192,N_11375);
nand U12510 (N_12510,N_11438,N_11339);
nand U12511 (N_12511,N_11974,N_11253);
or U12512 (N_12512,N_11946,N_11671);
and U12513 (N_12513,N_11669,N_11043);
nor U12514 (N_12514,N_11889,N_11610);
xor U12515 (N_12515,N_11032,N_11366);
or U12516 (N_12516,N_11229,N_11973);
xor U12517 (N_12517,N_11214,N_11948);
nor U12518 (N_12518,N_11924,N_11544);
or U12519 (N_12519,N_11702,N_11557);
nand U12520 (N_12520,N_11761,N_11386);
nand U12521 (N_12521,N_11391,N_11133);
nor U12522 (N_12522,N_11745,N_11070);
and U12523 (N_12523,N_11267,N_11881);
nor U12524 (N_12524,N_11074,N_11152);
nand U12525 (N_12525,N_11659,N_11340);
nor U12526 (N_12526,N_11866,N_11342);
xnor U12527 (N_12527,N_11309,N_11399);
and U12528 (N_12528,N_11574,N_11631);
and U12529 (N_12529,N_11614,N_11874);
and U12530 (N_12530,N_11051,N_11992);
nor U12531 (N_12531,N_11532,N_11298);
and U12532 (N_12532,N_11181,N_11664);
nor U12533 (N_12533,N_11651,N_11742);
xnor U12534 (N_12534,N_11254,N_11725);
and U12535 (N_12535,N_11572,N_11177);
and U12536 (N_12536,N_11603,N_11723);
and U12537 (N_12537,N_11200,N_11132);
nand U12538 (N_12538,N_11733,N_11646);
nand U12539 (N_12539,N_11386,N_11669);
xor U12540 (N_12540,N_11778,N_11400);
nand U12541 (N_12541,N_11752,N_11217);
nand U12542 (N_12542,N_11664,N_11329);
or U12543 (N_12543,N_11426,N_11610);
nor U12544 (N_12544,N_11895,N_11761);
or U12545 (N_12545,N_11096,N_11879);
or U12546 (N_12546,N_11114,N_11778);
nor U12547 (N_12547,N_11361,N_11696);
nor U12548 (N_12548,N_11079,N_11570);
nand U12549 (N_12549,N_11275,N_11567);
and U12550 (N_12550,N_11507,N_11338);
nand U12551 (N_12551,N_11888,N_11492);
or U12552 (N_12552,N_11125,N_11148);
or U12553 (N_12553,N_11005,N_11068);
nor U12554 (N_12554,N_11175,N_11074);
and U12555 (N_12555,N_11150,N_11957);
or U12556 (N_12556,N_11886,N_11278);
or U12557 (N_12557,N_11548,N_11782);
or U12558 (N_12558,N_11921,N_11243);
nand U12559 (N_12559,N_11003,N_11389);
and U12560 (N_12560,N_11268,N_11659);
nor U12561 (N_12561,N_11192,N_11908);
or U12562 (N_12562,N_11379,N_11988);
nand U12563 (N_12563,N_11597,N_11764);
or U12564 (N_12564,N_11287,N_11498);
nor U12565 (N_12565,N_11877,N_11909);
or U12566 (N_12566,N_11381,N_11060);
or U12567 (N_12567,N_11277,N_11961);
xor U12568 (N_12568,N_11155,N_11275);
nand U12569 (N_12569,N_11561,N_11936);
or U12570 (N_12570,N_11453,N_11767);
xnor U12571 (N_12571,N_11090,N_11916);
and U12572 (N_12572,N_11700,N_11299);
and U12573 (N_12573,N_11151,N_11958);
or U12574 (N_12574,N_11059,N_11264);
or U12575 (N_12575,N_11258,N_11236);
xor U12576 (N_12576,N_11417,N_11659);
and U12577 (N_12577,N_11524,N_11825);
nor U12578 (N_12578,N_11636,N_11086);
and U12579 (N_12579,N_11256,N_11282);
or U12580 (N_12580,N_11037,N_11406);
and U12581 (N_12581,N_11776,N_11268);
xor U12582 (N_12582,N_11538,N_11524);
xnor U12583 (N_12583,N_11623,N_11826);
and U12584 (N_12584,N_11747,N_11036);
nor U12585 (N_12585,N_11919,N_11595);
nand U12586 (N_12586,N_11452,N_11445);
nor U12587 (N_12587,N_11296,N_11180);
or U12588 (N_12588,N_11597,N_11095);
nor U12589 (N_12589,N_11942,N_11471);
xor U12590 (N_12590,N_11125,N_11572);
xor U12591 (N_12591,N_11056,N_11217);
nor U12592 (N_12592,N_11609,N_11199);
nor U12593 (N_12593,N_11446,N_11330);
xnor U12594 (N_12594,N_11971,N_11656);
nand U12595 (N_12595,N_11766,N_11217);
nor U12596 (N_12596,N_11602,N_11893);
and U12597 (N_12597,N_11528,N_11234);
xnor U12598 (N_12598,N_11784,N_11537);
and U12599 (N_12599,N_11410,N_11358);
nand U12600 (N_12600,N_11499,N_11373);
or U12601 (N_12601,N_11177,N_11757);
nor U12602 (N_12602,N_11877,N_11679);
nand U12603 (N_12603,N_11563,N_11976);
and U12604 (N_12604,N_11967,N_11194);
nand U12605 (N_12605,N_11433,N_11528);
xor U12606 (N_12606,N_11544,N_11322);
xnor U12607 (N_12607,N_11510,N_11583);
and U12608 (N_12608,N_11266,N_11186);
and U12609 (N_12609,N_11014,N_11821);
xor U12610 (N_12610,N_11764,N_11384);
or U12611 (N_12611,N_11048,N_11884);
nand U12612 (N_12612,N_11812,N_11450);
nor U12613 (N_12613,N_11148,N_11135);
xor U12614 (N_12614,N_11490,N_11312);
nand U12615 (N_12615,N_11214,N_11785);
nor U12616 (N_12616,N_11709,N_11695);
and U12617 (N_12617,N_11922,N_11040);
nand U12618 (N_12618,N_11980,N_11641);
xnor U12619 (N_12619,N_11284,N_11655);
xnor U12620 (N_12620,N_11812,N_11178);
nor U12621 (N_12621,N_11103,N_11260);
nor U12622 (N_12622,N_11165,N_11239);
nor U12623 (N_12623,N_11442,N_11759);
nand U12624 (N_12624,N_11764,N_11019);
xor U12625 (N_12625,N_11357,N_11170);
nor U12626 (N_12626,N_11273,N_11752);
nand U12627 (N_12627,N_11786,N_11544);
xor U12628 (N_12628,N_11535,N_11587);
xnor U12629 (N_12629,N_11234,N_11077);
nand U12630 (N_12630,N_11312,N_11522);
or U12631 (N_12631,N_11499,N_11466);
xnor U12632 (N_12632,N_11784,N_11558);
or U12633 (N_12633,N_11116,N_11473);
xnor U12634 (N_12634,N_11688,N_11404);
nand U12635 (N_12635,N_11725,N_11137);
or U12636 (N_12636,N_11632,N_11076);
or U12637 (N_12637,N_11509,N_11867);
or U12638 (N_12638,N_11363,N_11625);
nand U12639 (N_12639,N_11578,N_11064);
nand U12640 (N_12640,N_11540,N_11233);
xnor U12641 (N_12641,N_11754,N_11014);
and U12642 (N_12642,N_11010,N_11864);
nand U12643 (N_12643,N_11031,N_11483);
nand U12644 (N_12644,N_11740,N_11963);
or U12645 (N_12645,N_11294,N_11241);
nand U12646 (N_12646,N_11866,N_11594);
nand U12647 (N_12647,N_11738,N_11440);
nand U12648 (N_12648,N_11228,N_11093);
and U12649 (N_12649,N_11280,N_11957);
xor U12650 (N_12650,N_11983,N_11387);
nand U12651 (N_12651,N_11607,N_11958);
xor U12652 (N_12652,N_11808,N_11608);
or U12653 (N_12653,N_11345,N_11651);
or U12654 (N_12654,N_11892,N_11219);
xnor U12655 (N_12655,N_11796,N_11093);
nand U12656 (N_12656,N_11882,N_11687);
and U12657 (N_12657,N_11774,N_11193);
and U12658 (N_12658,N_11296,N_11406);
nand U12659 (N_12659,N_11427,N_11751);
nor U12660 (N_12660,N_11213,N_11757);
nor U12661 (N_12661,N_11077,N_11459);
xor U12662 (N_12662,N_11883,N_11960);
nand U12663 (N_12663,N_11406,N_11984);
or U12664 (N_12664,N_11195,N_11762);
nand U12665 (N_12665,N_11437,N_11255);
nand U12666 (N_12666,N_11633,N_11185);
and U12667 (N_12667,N_11535,N_11951);
xnor U12668 (N_12668,N_11515,N_11986);
nor U12669 (N_12669,N_11753,N_11232);
xnor U12670 (N_12670,N_11214,N_11156);
xor U12671 (N_12671,N_11045,N_11937);
xnor U12672 (N_12672,N_11591,N_11721);
xor U12673 (N_12673,N_11295,N_11983);
and U12674 (N_12674,N_11935,N_11934);
xnor U12675 (N_12675,N_11739,N_11079);
or U12676 (N_12676,N_11997,N_11298);
or U12677 (N_12677,N_11297,N_11762);
or U12678 (N_12678,N_11187,N_11230);
or U12679 (N_12679,N_11917,N_11140);
nand U12680 (N_12680,N_11729,N_11749);
nand U12681 (N_12681,N_11443,N_11163);
nand U12682 (N_12682,N_11195,N_11947);
and U12683 (N_12683,N_11978,N_11092);
xor U12684 (N_12684,N_11924,N_11456);
or U12685 (N_12685,N_11095,N_11575);
xnor U12686 (N_12686,N_11256,N_11226);
and U12687 (N_12687,N_11698,N_11403);
and U12688 (N_12688,N_11946,N_11976);
and U12689 (N_12689,N_11743,N_11483);
nand U12690 (N_12690,N_11547,N_11715);
or U12691 (N_12691,N_11679,N_11603);
and U12692 (N_12692,N_11563,N_11622);
nor U12693 (N_12693,N_11194,N_11628);
nand U12694 (N_12694,N_11969,N_11351);
or U12695 (N_12695,N_11346,N_11182);
nand U12696 (N_12696,N_11836,N_11326);
nor U12697 (N_12697,N_11150,N_11662);
and U12698 (N_12698,N_11948,N_11726);
xnor U12699 (N_12699,N_11837,N_11466);
xor U12700 (N_12700,N_11585,N_11417);
nand U12701 (N_12701,N_11217,N_11977);
nor U12702 (N_12702,N_11809,N_11691);
and U12703 (N_12703,N_11788,N_11545);
or U12704 (N_12704,N_11266,N_11553);
nand U12705 (N_12705,N_11958,N_11807);
nand U12706 (N_12706,N_11772,N_11648);
xnor U12707 (N_12707,N_11680,N_11058);
nor U12708 (N_12708,N_11047,N_11642);
or U12709 (N_12709,N_11583,N_11651);
xor U12710 (N_12710,N_11640,N_11844);
nand U12711 (N_12711,N_11165,N_11415);
nor U12712 (N_12712,N_11825,N_11665);
xor U12713 (N_12713,N_11487,N_11759);
nor U12714 (N_12714,N_11351,N_11522);
or U12715 (N_12715,N_11121,N_11197);
xor U12716 (N_12716,N_11099,N_11296);
xnor U12717 (N_12717,N_11955,N_11426);
nor U12718 (N_12718,N_11402,N_11062);
nor U12719 (N_12719,N_11238,N_11744);
nand U12720 (N_12720,N_11756,N_11976);
nand U12721 (N_12721,N_11572,N_11162);
nor U12722 (N_12722,N_11522,N_11338);
xor U12723 (N_12723,N_11991,N_11039);
or U12724 (N_12724,N_11570,N_11936);
nor U12725 (N_12725,N_11841,N_11081);
xor U12726 (N_12726,N_11817,N_11887);
and U12727 (N_12727,N_11099,N_11817);
xor U12728 (N_12728,N_11353,N_11570);
nand U12729 (N_12729,N_11347,N_11327);
nor U12730 (N_12730,N_11481,N_11395);
xor U12731 (N_12731,N_11646,N_11021);
nor U12732 (N_12732,N_11059,N_11455);
nand U12733 (N_12733,N_11909,N_11638);
nor U12734 (N_12734,N_11718,N_11693);
nand U12735 (N_12735,N_11677,N_11020);
or U12736 (N_12736,N_11788,N_11004);
xnor U12737 (N_12737,N_11819,N_11879);
or U12738 (N_12738,N_11189,N_11969);
nor U12739 (N_12739,N_11469,N_11021);
and U12740 (N_12740,N_11910,N_11168);
nor U12741 (N_12741,N_11521,N_11405);
and U12742 (N_12742,N_11614,N_11540);
nor U12743 (N_12743,N_11669,N_11530);
and U12744 (N_12744,N_11938,N_11595);
xnor U12745 (N_12745,N_11317,N_11937);
nor U12746 (N_12746,N_11636,N_11635);
xnor U12747 (N_12747,N_11388,N_11568);
xnor U12748 (N_12748,N_11365,N_11342);
or U12749 (N_12749,N_11900,N_11677);
and U12750 (N_12750,N_11212,N_11375);
and U12751 (N_12751,N_11749,N_11048);
nand U12752 (N_12752,N_11140,N_11507);
nor U12753 (N_12753,N_11544,N_11132);
or U12754 (N_12754,N_11046,N_11678);
or U12755 (N_12755,N_11012,N_11267);
xor U12756 (N_12756,N_11722,N_11215);
nand U12757 (N_12757,N_11499,N_11425);
nor U12758 (N_12758,N_11608,N_11403);
nor U12759 (N_12759,N_11065,N_11716);
xor U12760 (N_12760,N_11856,N_11384);
and U12761 (N_12761,N_11006,N_11932);
and U12762 (N_12762,N_11988,N_11698);
xor U12763 (N_12763,N_11621,N_11947);
and U12764 (N_12764,N_11397,N_11912);
xor U12765 (N_12765,N_11317,N_11991);
or U12766 (N_12766,N_11898,N_11246);
or U12767 (N_12767,N_11705,N_11259);
and U12768 (N_12768,N_11335,N_11512);
and U12769 (N_12769,N_11558,N_11231);
nor U12770 (N_12770,N_11451,N_11852);
and U12771 (N_12771,N_11417,N_11952);
or U12772 (N_12772,N_11176,N_11233);
or U12773 (N_12773,N_11076,N_11913);
nand U12774 (N_12774,N_11733,N_11329);
or U12775 (N_12775,N_11958,N_11993);
xor U12776 (N_12776,N_11643,N_11836);
xor U12777 (N_12777,N_11950,N_11247);
and U12778 (N_12778,N_11817,N_11966);
or U12779 (N_12779,N_11296,N_11172);
nor U12780 (N_12780,N_11160,N_11840);
and U12781 (N_12781,N_11523,N_11185);
and U12782 (N_12782,N_11570,N_11824);
or U12783 (N_12783,N_11795,N_11980);
and U12784 (N_12784,N_11077,N_11842);
xnor U12785 (N_12785,N_11959,N_11010);
and U12786 (N_12786,N_11268,N_11661);
nand U12787 (N_12787,N_11908,N_11683);
xor U12788 (N_12788,N_11988,N_11272);
and U12789 (N_12789,N_11155,N_11296);
nand U12790 (N_12790,N_11141,N_11083);
xnor U12791 (N_12791,N_11260,N_11059);
xnor U12792 (N_12792,N_11452,N_11448);
nand U12793 (N_12793,N_11879,N_11549);
and U12794 (N_12794,N_11476,N_11502);
or U12795 (N_12795,N_11198,N_11935);
or U12796 (N_12796,N_11448,N_11979);
nor U12797 (N_12797,N_11100,N_11665);
or U12798 (N_12798,N_11995,N_11699);
xor U12799 (N_12799,N_11376,N_11441);
nor U12800 (N_12800,N_11836,N_11751);
or U12801 (N_12801,N_11252,N_11845);
or U12802 (N_12802,N_11749,N_11075);
and U12803 (N_12803,N_11754,N_11570);
nor U12804 (N_12804,N_11214,N_11178);
nor U12805 (N_12805,N_11415,N_11457);
nor U12806 (N_12806,N_11687,N_11908);
nor U12807 (N_12807,N_11610,N_11366);
nor U12808 (N_12808,N_11737,N_11590);
or U12809 (N_12809,N_11141,N_11872);
nor U12810 (N_12810,N_11922,N_11203);
and U12811 (N_12811,N_11879,N_11521);
and U12812 (N_12812,N_11693,N_11272);
and U12813 (N_12813,N_11755,N_11975);
or U12814 (N_12814,N_11978,N_11677);
xnor U12815 (N_12815,N_11017,N_11543);
or U12816 (N_12816,N_11580,N_11064);
and U12817 (N_12817,N_11049,N_11714);
nand U12818 (N_12818,N_11317,N_11891);
xnor U12819 (N_12819,N_11671,N_11588);
nor U12820 (N_12820,N_11998,N_11894);
and U12821 (N_12821,N_11325,N_11685);
or U12822 (N_12822,N_11070,N_11944);
or U12823 (N_12823,N_11884,N_11659);
xor U12824 (N_12824,N_11574,N_11385);
xnor U12825 (N_12825,N_11214,N_11442);
nand U12826 (N_12826,N_11024,N_11783);
or U12827 (N_12827,N_11286,N_11547);
and U12828 (N_12828,N_11371,N_11248);
or U12829 (N_12829,N_11435,N_11890);
and U12830 (N_12830,N_11862,N_11684);
or U12831 (N_12831,N_11853,N_11329);
or U12832 (N_12832,N_11519,N_11217);
nand U12833 (N_12833,N_11693,N_11764);
xor U12834 (N_12834,N_11190,N_11043);
xor U12835 (N_12835,N_11856,N_11526);
and U12836 (N_12836,N_11556,N_11655);
nor U12837 (N_12837,N_11796,N_11389);
nor U12838 (N_12838,N_11982,N_11120);
xor U12839 (N_12839,N_11122,N_11827);
nand U12840 (N_12840,N_11865,N_11471);
xnor U12841 (N_12841,N_11082,N_11116);
xor U12842 (N_12842,N_11766,N_11128);
xnor U12843 (N_12843,N_11744,N_11257);
nor U12844 (N_12844,N_11956,N_11764);
nor U12845 (N_12845,N_11634,N_11956);
xor U12846 (N_12846,N_11315,N_11814);
xor U12847 (N_12847,N_11628,N_11220);
or U12848 (N_12848,N_11287,N_11637);
nand U12849 (N_12849,N_11163,N_11772);
nor U12850 (N_12850,N_11411,N_11263);
and U12851 (N_12851,N_11672,N_11922);
nand U12852 (N_12852,N_11957,N_11005);
xnor U12853 (N_12853,N_11913,N_11537);
xnor U12854 (N_12854,N_11881,N_11182);
xnor U12855 (N_12855,N_11454,N_11983);
nand U12856 (N_12856,N_11062,N_11068);
nand U12857 (N_12857,N_11195,N_11233);
or U12858 (N_12858,N_11484,N_11441);
xor U12859 (N_12859,N_11218,N_11612);
or U12860 (N_12860,N_11520,N_11519);
and U12861 (N_12861,N_11941,N_11734);
or U12862 (N_12862,N_11576,N_11276);
or U12863 (N_12863,N_11818,N_11265);
or U12864 (N_12864,N_11913,N_11644);
or U12865 (N_12865,N_11040,N_11841);
nand U12866 (N_12866,N_11021,N_11004);
or U12867 (N_12867,N_11919,N_11754);
and U12868 (N_12868,N_11045,N_11531);
xor U12869 (N_12869,N_11814,N_11256);
and U12870 (N_12870,N_11296,N_11540);
or U12871 (N_12871,N_11501,N_11224);
and U12872 (N_12872,N_11369,N_11132);
xnor U12873 (N_12873,N_11758,N_11278);
and U12874 (N_12874,N_11034,N_11730);
nor U12875 (N_12875,N_11349,N_11967);
or U12876 (N_12876,N_11841,N_11606);
nand U12877 (N_12877,N_11697,N_11159);
nand U12878 (N_12878,N_11037,N_11894);
nand U12879 (N_12879,N_11032,N_11721);
nor U12880 (N_12880,N_11354,N_11988);
nand U12881 (N_12881,N_11204,N_11513);
or U12882 (N_12882,N_11805,N_11027);
nor U12883 (N_12883,N_11298,N_11614);
or U12884 (N_12884,N_11238,N_11320);
or U12885 (N_12885,N_11295,N_11029);
xor U12886 (N_12886,N_11329,N_11768);
and U12887 (N_12887,N_11589,N_11332);
or U12888 (N_12888,N_11029,N_11983);
nand U12889 (N_12889,N_11988,N_11154);
or U12890 (N_12890,N_11138,N_11590);
and U12891 (N_12891,N_11375,N_11672);
nand U12892 (N_12892,N_11290,N_11595);
xnor U12893 (N_12893,N_11007,N_11333);
nand U12894 (N_12894,N_11561,N_11405);
or U12895 (N_12895,N_11423,N_11744);
or U12896 (N_12896,N_11295,N_11478);
xnor U12897 (N_12897,N_11027,N_11894);
nor U12898 (N_12898,N_11129,N_11420);
and U12899 (N_12899,N_11735,N_11266);
nand U12900 (N_12900,N_11132,N_11221);
nor U12901 (N_12901,N_11740,N_11104);
and U12902 (N_12902,N_11940,N_11393);
nand U12903 (N_12903,N_11918,N_11319);
or U12904 (N_12904,N_11869,N_11513);
and U12905 (N_12905,N_11842,N_11416);
xor U12906 (N_12906,N_11740,N_11178);
or U12907 (N_12907,N_11937,N_11410);
nand U12908 (N_12908,N_11738,N_11324);
and U12909 (N_12909,N_11473,N_11970);
nand U12910 (N_12910,N_11069,N_11783);
nand U12911 (N_12911,N_11284,N_11475);
or U12912 (N_12912,N_11614,N_11268);
xnor U12913 (N_12913,N_11544,N_11662);
xnor U12914 (N_12914,N_11137,N_11252);
and U12915 (N_12915,N_11748,N_11437);
nand U12916 (N_12916,N_11741,N_11263);
or U12917 (N_12917,N_11929,N_11062);
nor U12918 (N_12918,N_11992,N_11960);
or U12919 (N_12919,N_11536,N_11496);
and U12920 (N_12920,N_11631,N_11148);
and U12921 (N_12921,N_11036,N_11056);
nand U12922 (N_12922,N_11632,N_11737);
and U12923 (N_12923,N_11116,N_11176);
or U12924 (N_12924,N_11864,N_11711);
nor U12925 (N_12925,N_11383,N_11256);
and U12926 (N_12926,N_11807,N_11603);
and U12927 (N_12927,N_11190,N_11540);
or U12928 (N_12928,N_11147,N_11947);
nor U12929 (N_12929,N_11532,N_11816);
xor U12930 (N_12930,N_11192,N_11919);
xnor U12931 (N_12931,N_11245,N_11887);
or U12932 (N_12932,N_11867,N_11705);
and U12933 (N_12933,N_11553,N_11405);
or U12934 (N_12934,N_11308,N_11111);
nand U12935 (N_12935,N_11487,N_11027);
nor U12936 (N_12936,N_11364,N_11114);
nand U12937 (N_12937,N_11126,N_11558);
nand U12938 (N_12938,N_11970,N_11492);
and U12939 (N_12939,N_11010,N_11360);
nand U12940 (N_12940,N_11711,N_11443);
and U12941 (N_12941,N_11950,N_11793);
nor U12942 (N_12942,N_11236,N_11992);
xnor U12943 (N_12943,N_11424,N_11624);
and U12944 (N_12944,N_11632,N_11681);
nor U12945 (N_12945,N_11148,N_11413);
or U12946 (N_12946,N_11550,N_11302);
or U12947 (N_12947,N_11945,N_11870);
nand U12948 (N_12948,N_11081,N_11044);
or U12949 (N_12949,N_11540,N_11588);
or U12950 (N_12950,N_11791,N_11299);
nand U12951 (N_12951,N_11972,N_11596);
nor U12952 (N_12952,N_11284,N_11519);
or U12953 (N_12953,N_11609,N_11916);
or U12954 (N_12954,N_11142,N_11434);
and U12955 (N_12955,N_11147,N_11326);
and U12956 (N_12956,N_11027,N_11039);
nor U12957 (N_12957,N_11060,N_11616);
nor U12958 (N_12958,N_11933,N_11594);
nor U12959 (N_12959,N_11829,N_11848);
and U12960 (N_12960,N_11309,N_11409);
or U12961 (N_12961,N_11686,N_11108);
nand U12962 (N_12962,N_11232,N_11923);
and U12963 (N_12963,N_11033,N_11683);
and U12964 (N_12964,N_11333,N_11485);
or U12965 (N_12965,N_11267,N_11166);
or U12966 (N_12966,N_11733,N_11571);
and U12967 (N_12967,N_11292,N_11223);
xnor U12968 (N_12968,N_11732,N_11550);
nand U12969 (N_12969,N_11077,N_11691);
and U12970 (N_12970,N_11061,N_11503);
xor U12971 (N_12971,N_11050,N_11918);
and U12972 (N_12972,N_11697,N_11114);
nor U12973 (N_12973,N_11198,N_11344);
and U12974 (N_12974,N_11240,N_11397);
nand U12975 (N_12975,N_11667,N_11747);
nor U12976 (N_12976,N_11596,N_11281);
or U12977 (N_12977,N_11823,N_11265);
or U12978 (N_12978,N_11691,N_11032);
xnor U12979 (N_12979,N_11950,N_11065);
nor U12980 (N_12980,N_11545,N_11140);
and U12981 (N_12981,N_11362,N_11701);
nor U12982 (N_12982,N_11699,N_11384);
or U12983 (N_12983,N_11145,N_11877);
or U12984 (N_12984,N_11672,N_11171);
or U12985 (N_12985,N_11642,N_11408);
nor U12986 (N_12986,N_11954,N_11916);
xor U12987 (N_12987,N_11647,N_11914);
nor U12988 (N_12988,N_11694,N_11231);
nand U12989 (N_12989,N_11792,N_11890);
or U12990 (N_12990,N_11617,N_11305);
and U12991 (N_12991,N_11742,N_11571);
and U12992 (N_12992,N_11560,N_11669);
and U12993 (N_12993,N_11689,N_11808);
nor U12994 (N_12994,N_11381,N_11858);
xor U12995 (N_12995,N_11156,N_11827);
and U12996 (N_12996,N_11489,N_11561);
and U12997 (N_12997,N_11749,N_11245);
nand U12998 (N_12998,N_11989,N_11691);
and U12999 (N_12999,N_11221,N_11379);
or U13000 (N_13000,N_12153,N_12084);
or U13001 (N_13001,N_12013,N_12208);
nor U13002 (N_13002,N_12272,N_12509);
and U13003 (N_13003,N_12814,N_12802);
nand U13004 (N_13004,N_12546,N_12493);
nor U13005 (N_13005,N_12124,N_12599);
or U13006 (N_13006,N_12350,N_12849);
and U13007 (N_13007,N_12897,N_12488);
nand U13008 (N_13008,N_12734,N_12742);
xnor U13009 (N_13009,N_12939,N_12641);
and U13010 (N_13010,N_12807,N_12579);
xor U13011 (N_13011,N_12673,N_12766);
nor U13012 (N_13012,N_12098,N_12291);
and U13013 (N_13013,N_12097,N_12868);
nand U13014 (N_13014,N_12068,N_12470);
nand U13015 (N_13015,N_12305,N_12838);
or U13016 (N_13016,N_12194,N_12709);
nand U13017 (N_13017,N_12569,N_12675);
nand U13018 (N_13018,N_12544,N_12558);
nand U13019 (N_13019,N_12358,N_12691);
xnor U13020 (N_13020,N_12292,N_12180);
and U13021 (N_13021,N_12765,N_12039);
or U13022 (N_13022,N_12732,N_12452);
nand U13023 (N_13023,N_12259,N_12988);
or U13024 (N_13024,N_12371,N_12937);
xnor U13025 (N_13025,N_12087,N_12037);
nand U13026 (N_13026,N_12888,N_12430);
nor U13027 (N_13027,N_12922,N_12933);
and U13028 (N_13028,N_12900,N_12007);
or U13029 (N_13029,N_12971,N_12143);
or U13030 (N_13030,N_12154,N_12150);
nor U13031 (N_13031,N_12095,N_12854);
nor U13032 (N_13032,N_12789,N_12425);
or U13033 (N_13033,N_12514,N_12030);
nand U13034 (N_13034,N_12716,N_12170);
nand U13035 (N_13035,N_12481,N_12820);
nand U13036 (N_13036,N_12835,N_12775);
xor U13037 (N_13037,N_12034,N_12252);
nand U13038 (N_13038,N_12307,N_12660);
and U13039 (N_13039,N_12472,N_12201);
nand U13040 (N_13040,N_12287,N_12202);
nor U13041 (N_13041,N_12676,N_12330);
or U13042 (N_13042,N_12998,N_12785);
nand U13043 (N_13043,N_12351,N_12538);
xnor U13044 (N_13044,N_12166,N_12889);
or U13045 (N_13045,N_12191,N_12815);
nor U13046 (N_13046,N_12256,N_12591);
nor U13047 (N_13047,N_12851,N_12562);
xor U13048 (N_13048,N_12772,N_12584);
nand U13049 (N_13049,N_12320,N_12184);
or U13050 (N_13050,N_12500,N_12271);
nand U13051 (N_13051,N_12042,N_12416);
xor U13052 (N_13052,N_12531,N_12883);
or U13053 (N_13053,N_12834,N_12739);
nor U13054 (N_13054,N_12915,N_12677);
xor U13055 (N_13055,N_12205,N_12419);
or U13056 (N_13056,N_12703,N_12961);
nor U13057 (N_13057,N_12678,N_12596);
nor U13058 (N_13058,N_12576,N_12125);
or U13059 (N_13059,N_12925,N_12974);
or U13060 (N_13060,N_12400,N_12795);
nand U13061 (N_13061,N_12265,N_12685);
nor U13062 (N_13062,N_12981,N_12704);
and U13063 (N_13063,N_12250,N_12701);
or U13064 (N_13064,N_12715,N_12659);
or U13065 (N_13065,N_12899,N_12951);
nor U13066 (N_13066,N_12636,N_12424);
or U13067 (N_13067,N_12592,N_12746);
or U13068 (N_13068,N_12484,N_12426);
nand U13069 (N_13069,N_12318,N_12188);
nand U13070 (N_13070,N_12916,N_12203);
nor U13071 (N_13071,N_12940,N_12080);
and U13072 (N_13072,N_12566,N_12295);
or U13073 (N_13073,N_12541,N_12075);
xnor U13074 (N_13074,N_12026,N_12163);
or U13075 (N_13075,N_12268,N_12130);
nor U13076 (N_13076,N_12520,N_12726);
nor U13077 (N_13077,N_12930,N_12829);
xor U13078 (N_13078,N_12453,N_12357);
xor U13079 (N_13079,N_12513,N_12662);
and U13080 (N_13080,N_12491,N_12728);
xor U13081 (N_13081,N_12323,N_12758);
and U13082 (N_13082,N_12244,N_12567);
xor U13083 (N_13083,N_12610,N_12864);
nor U13084 (N_13084,N_12078,N_12260);
nand U13085 (N_13085,N_12409,N_12114);
xnor U13086 (N_13086,N_12759,N_12539);
or U13087 (N_13087,N_12919,N_12668);
and U13088 (N_13088,N_12288,N_12324);
nor U13089 (N_13089,N_12984,N_12131);
nand U13090 (N_13090,N_12107,N_12861);
nor U13091 (N_13091,N_12833,N_12568);
or U13092 (N_13092,N_12683,N_12588);
or U13093 (N_13093,N_12870,N_12251);
or U13094 (N_13094,N_12370,N_12274);
or U13095 (N_13095,N_12178,N_12782);
nor U13096 (N_13096,N_12058,N_12386);
nor U13097 (N_13097,N_12947,N_12344);
and U13098 (N_13098,N_12471,N_12059);
nand U13099 (N_13099,N_12550,N_12101);
nor U13100 (N_13100,N_12924,N_12161);
and U13101 (N_13101,N_12905,N_12867);
xor U13102 (N_13102,N_12856,N_12245);
or U13103 (N_13103,N_12828,N_12760);
xnor U13104 (N_13104,N_12656,N_12317);
and U13105 (N_13105,N_12714,N_12985);
nor U13106 (N_13106,N_12233,N_12293);
and U13107 (N_13107,N_12296,N_12067);
xor U13108 (N_13108,N_12122,N_12139);
nand U13109 (N_13109,N_12556,N_12540);
nor U13110 (N_13110,N_12025,N_12956);
xnor U13111 (N_13111,N_12804,N_12010);
xor U13112 (N_13112,N_12247,N_12783);
and U13113 (N_13113,N_12816,N_12637);
or U13114 (N_13114,N_12149,N_12047);
xor U13115 (N_13115,N_12631,N_12118);
nand U13116 (N_13116,N_12222,N_12112);
nor U13117 (N_13117,N_12246,N_12780);
and U13118 (N_13118,N_12770,N_12092);
nor U13119 (N_13119,N_12031,N_12774);
or U13120 (N_13120,N_12137,N_12741);
nand U13121 (N_13121,N_12313,N_12962);
nand U13122 (N_13122,N_12411,N_12622);
xnor U13123 (N_13123,N_12696,N_12121);
or U13124 (N_13124,N_12088,N_12649);
nor U13125 (N_13125,N_12454,N_12601);
or U13126 (N_13126,N_12705,N_12434);
xnor U13127 (N_13127,N_12792,N_12938);
nor U13128 (N_13128,N_12492,N_12983);
nand U13129 (N_13129,N_12982,N_12955);
nor U13130 (N_13130,N_12748,N_12616);
or U13131 (N_13131,N_12308,N_12621);
nand U13132 (N_13132,N_12585,N_12410);
nand U13133 (N_13133,N_12496,N_12722);
xnor U13134 (N_13134,N_12439,N_12223);
or U13135 (N_13135,N_12022,N_12231);
and U13136 (N_13136,N_12160,N_12927);
and U13137 (N_13137,N_12482,N_12762);
xnor U13138 (N_13138,N_12960,N_12275);
or U13139 (N_13139,N_12263,N_12364);
or U13140 (N_13140,N_12526,N_12363);
xnor U13141 (N_13141,N_12487,N_12322);
xnor U13142 (N_13142,N_12229,N_12874);
nor U13143 (N_13143,N_12436,N_12427);
nor U13144 (N_13144,N_12447,N_12269);
and U13145 (N_13145,N_12549,N_12917);
nor U13146 (N_13146,N_12413,N_12301);
xnor U13147 (N_13147,N_12672,N_12489);
nand U13148 (N_13148,N_12336,N_12642);
nand U13149 (N_13149,N_12485,N_12060);
nand U13150 (N_13150,N_12328,N_12355);
and U13151 (N_13151,N_12294,N_12535);
nand U13152 (N_13152,N_12837,N_12950);
or U13153 (N_13153,N_12908,N_12614);
xnor U13154 (N_13154,N_12796,N_12926);
nand U13155 (N_13155,N_12183,N_12907);
or U13156 (N_13156,N_12803,N_12321);
and U13157 (N_13157,N_12629,N_12147);
nand U13158 (N_13158,N_12559,N_12063);
nor U13159 (N_13159,N_12083,N_12375);
xor U13160 (N_13160,N_12516,N_12634);
and U13161 (N_13161,N_12605,N_12199);
nand U13162 (N_13162,N_12749,N_12658);
and U13163 (N_13163,N_12994,N_12220);
nand U13164 (N_13164,N_12589,N_12182);
nand U13165 (N_13165,N_12109,N_12133);
nand U13166 (N_13166,N_12852,N_12906);
and U13167 (N_13167,N_12253,N_12127);
nor U13168 (N_13168,N_12467,N_12155);
nor U13169 (N_13169,N_12151,N_12727);
and U13170 (N_13170,N_12543,N_12992);
nand U13171 (N_13171,N_12209,N_12056);
nand U13172 (N_13172,N_12397,N_12946);
and U13173 (N_13173,N_12051,N_12811);
and U13174 (N_13174,N_12504,N_12967);
nand U13175 (N_13175,N_12561,N_12314);
nor U13176 (N_13176,N_12876,N_12192);
or U13177 (N_13177,N_12670,N_12942);
xnor U13178 (N_13178,N_12976,N_12718);
nor U13179 (N_13179,N_12573,N_12882);
xor U13180 (N_13180,N_12120,N_12412);
nor U13181 (N_13181,N_12128,N_12894);
nor U13182 (N_13182,N_12377,N_12359);
or U13183 (N_13183,N_12490,N_12141);
and U13184 (N_13184,N_12602,N_12327);
nand U13185 (N_13185,N_12999,N_12918);
nor U13186 (N_13186,N_12686,N_12764);
nand U13187 (N_13187,N_12473,N_12266);
xnor U13188 (N_13188,N_12590,N_12966);
or U13189 (N_13189,N_12819,N_12074);
and U13190 (N_13190,N_12360,N_12455);
nor U13191 (N_13191,N_12390,N_12054);
xor U13192 (N_13192,N_12587,N_12145);
and U13193 (N_13193,N_12529,N_12402);
or U13194 (N_13194,N_12171,N_12929);
or U13195 (N_13195,N_12625,N_12853);
xor U13196 (N_13196,N_12450,N_12329);
or U13197 (N_13197,N_12135,N_12699);
xnor U13198 (N_13198,N_12285,N_12255);
nor U13199 (N_13199,N_12639,N_12443);
xnor U13200 (N_13200,N_12763,N_12650);
and U13201 (N_13201,N_12624,N_12875);
or U13202 (N_13202,N_12018,N_12337);
or U13203 (N_13203,N_12957,N_12627);
or U13204 (N_13204,N_12666,N_12348);
nand U13205 (N_13205,N_12630,N_12494);
xnor U13206 (N_13206,N_12372,N_12415);
nor U13207 (N_13207,N_12707,N_12242);
and U13208 (N_13208,N_12527,N_12298);
nor U13209 (N_13209,N_12073,N_12560);
and U13210 (N_13210,N_12717,N_12657);
and U13211 (N_13211,N_12846,N_12302);
nand U13212 (N_13212,N_12794,N_12498);
and U13213 (N_13213,N_12196,N_12580);
and U13214 (N_13214,N_12928,N_12608);
and U13215 (N_13215,N_12089,N_12091);
nor U13216 (N_13216,N_12825,N_12033);
xnor U13217 (N_13217,N_12055,N_12679);
xor U13218 (N_13218,N_12214,N_12987);
or U13219 (N_13219,N_12847,N_12003);
nor U13220 (N_13220,N_12369,N_12381);
nor U13221 (N_13221,N_12700,N_12468);
xnor U13222 (N_13222,N_12647,N_12422);
nor U13223 (N_13223,N_12945,N_12440);
nand U13224 (N_13224,N_12028,N_12977);
nand U13225 (N_13225,N_12863,N_12609);
nand U13226 (N_13226,N_12167,N_12099);
and U13227 (N_13227,N_12206,N_12105);
nor U13228 (N_13228,N_12349,N_12552);
nand U13229 (N_13229,N_12423,N_12029);
and U13230 (N_13230,N_12019,N_12445);
or U13231 (N_13231,N_12248,N_12565);
nand U13232 (N_13232,N_12954,N_12653);
nand U13233 (N_13233,N_12532,N_12674);
nand U13234 (N_13234,N_12800,N_12667);
nand U13235 (N_13235,N_12048,N_12571);
nor U13236 (N_13236,N_12465,N_12462);
xnor U13237 (N_13237,N_12845,N_12923);
and U13238 (N_13238,N_12646,N_12618);
nand U13239 (N_13239,N_12404,N_12157);
or U13240 (N_13240,N_12784,N_12809);
and U13241 (N_13241,N_12973,N_12303);
nor U13242 (N_13242,N_12015,N_12689);
or U13243 (N_13243,N_12479,N_12389);
or U13244 (N_13244,N_12111,N_12175);
or U13245 (N_13245,N_12189,N_12378);
or U13246 (N_13246,N_12506,N_12551);
nor U13247 (N_13247,N_12510,N_12860);
xnor U13248 (N_13248,N_12881,N_12626);
nand U13249 (N_13249,N_12972,N_12172);
nand U13250 (N_13250,N_12093,N_12005);
nor U13251 (N_13251,N_12661,N_12286);
nor U13252 (N_13252,N_12790,N_12810);
xnor U13253 (N_13253,N_12264,N_12968);
or U13254 (N_13254,N_12574,N_12651);
nand U13255 (N_13255,N_12181,N_12451);
nand U13256 (N_13256,N_12177,N_12002);
xnor U13257 (N_13257,N_12200,N_12752);
nand U13258 (N_13258,N_12442,N_12799);
nor U13259 (N_13259,N_12258,N_12884);
xnor U13260 (N_13260,N_12776,N_12595);
and U13261 (N_13261,N_12781,N_12855);
xnor U13262 (N_13262,N_12949,N_12600);
nand U13263 (N_13263,N_12997,N_12499);
and U13264 (N_13264,N_12643,N_12195);
or U13265 (N_13265,N_12827,N_12038);
or U13266 (N_13266,N_12911,N_12553);
or U13267 (N_13267,N_12563,N_12207);
xor U13268 (N_13268,N_12542,N_12692);
xor U13269 (N_13269,N_12640,N_12212);
or U13270 (N_13270,N_12862,N_12697);
nand U13271 (N_13271,N_12335,N_12932);
nand U13272 (N_13272,N_12936,N_12433);
or U13273 (N_13273,N_12690,N_12289);
and U13274 (N_13274,N_12132,N_12986);
nor U13275 (N_13275,N_12980,N_12990);
nor U13276 (N_13276,N_12698,N_12332);
or U13277 (N_13277,N_12633,N_12645);
nor U13278 (N_13278,N_12354,N_12444);
nand U13279 (N_13279,N_12886,N_12197);
and U13280 (N_13280,N_12757,N_12831);
xor U13281 (N_13281,N_12594,N_12515);
nor U13282 (N_13282,N_12069,N_12094);
and U13283 (N_13283,N_12361,N_12964);
xnor U13284 (N_13284,N_12581,N_12779);
and U13285 (N_13285,N_12346,N_12943);
and U13286 (N_13286,N_12793,N_12952);
xnor U13287 (N_13287,N_12345,N_12036);
and U13288 (N_13288,N_12684,N_12116);
nor U13289 (N_13289,N_12437,N_12173);
nand U13290 (N_13290,N_12476,N_12613);
and U13291 (N_13291,N_12408,N_12877);
or U13292 (N_13292,N_12379,N_12747);
nand U13293 (N_13293,N_12041,N_12665);
nand U13294 (N_13294,N_12525,N_12719);
xnor U13295 (N_13295,N_12738,N_12431);
or U13296 (N_13296,N_12449,N_12428);
nand U13297 (N_13297,N_12777,N_12136);
and U13298 (N_13298,N_12575,N_12786);
nand U13299 (N_13299,N_12284,N_12388);
nand U13300 (N_13300,N_12458,N_12586);
nor U13301 (N_13301,N_12808,N_12989);
nor U13302 (N_13302,N_12912,N_12057);
xor U13303 (N_13303,N_12032,N_12866);
nand U13304 (N_13304,N_12934,N_12082);
nand U13305 (N_13305,N_12376,N_12680);
or U13306 (N_13306,N_12970,N_12230);
and U13307 (N_13307,N_12213,N_12469);
and U13308 (N_13308,N_12052,N_12228);
and U13309 (N_13309,N_12146,N_12953);
or U13310 (N_13310,N_12975,N_12459);
nand U13311 (N_13311,N_12909,N_12708);
and U13312 (N_13312,N_12832,N_12554);
nand U13313 (N_13313,N_12311,N_12024);
xnor U13314 (N_13314,N_12162,N_12090);
nor U13315 (N_13315,N_12713,N_12547);
nor U13316 (N_13316,N_12813,N_12570);
nor U13317 (N_13317,N_12309,N_12193);
xnor U13318 (N_13318,N_12306,N_12460);
or U13319 (N_13319,N_12237,N_12706);
xor U13320 (N_13320,N_12878,N_12046);
xor U13321 (N_13321,N_12014,N_12681);
nor U13322 (N_13322,N_12891,N_12035);
nand U13323 (N_13323,N_12577,N_12712);
nor U13324 (N_13324,N_12016,N_12027);
nand U13325 (N_13325,N_12695,N_12743);
and U13326 (N_13326,N_12343,N_12901);
and U13327 (N_13327,N_12339,N_12071);
nor U13328 (N_13328,N_12142,N_12021);
xnor U13329 (N_13329,N_12234,N_12395);
nand U13330 (N_13330,N_12316,N_12394);
and U13331 (N_13331,N_12232,N_12076);
nand U13332 (N_13332,N_12126,N_12227);
nand U13333 (N_13333,N_12903,N_12474);
xnor U13334 (N_13334,N_12420,N_12519);
and U13335 (N_13335,N_12996,N_12486);
nor U13336 (N_13336,N_12797,N_12902);
or U13337 (N_13337,N_12217,N_12300);
or U13338 (N_13338,N_12806,N_12805);
and U13339 (N_13339,N_12347,N_12597);
nor U13340 (N_13340,N_12582,N_12387);
xor U13341 (N_13341,N_12334,N_12898);
and U13342 (N_13342,N_12548,N_12963);
xor U13343 (N_13343,N_12865,N_12628);
or U13344 (N_13344,N_12115,N_12564);
nor U13345 (N_13345,N_12842,N_12545);
xor U13346 (N_13346,N_12935,N_12872);
and U13347 (N_13347,N_12096,N_12818);
or U13348 (N_13348,N_12262,N_12373);
nand U13349 (N_13349,N_12104,N_12297);
nor U13350 (N_13350,N_12312,N_12991);
nand U13351 (N_13351,N_12896,N_12761);
and U13352 (N_13352,N_12152,N_12839);
and U13353 (N_13353,N_12654,N_12755);
nor U13354 (N_13354,N_12848,N_12751);
nand U13355 (N_13355,N_12070,N_12771);
nor U13356 (N_13356,N_12687,N_12663);
xor U13357 (N_13357,N_12736,N_12393);
nand U13358 (N_13358,N_12403,N_12533);
and U13359 (N_13359,N_12857,N_12119);
xnor U13360 (N_13360,N_12017,N_12503);
and U13361 (N_13361,N_12249,N_12066);
and U13362 (N_13362,N_12277,N_12421);
or U13363 (N_13363,N_12081,N_12368);
nor U13364 (N_13364,N_12826,N_12744);
nor U13365 (N_13365,N_12100,N_12572);
nand U13366 (N_13366,N_12477,N_12843);
xnor U13367 (N_13367,N_12959,N_12521);
nor U13368 (N_13368,N_12969,N_12401);
xor U13369 (N_13369,N_12064,N_12108);
nor U13370 (N_13370,N_12004,N_12754);
or U13371 (N_13371,N_12085,N_12186);
xor U13372 (N_13372,N_12282,N_12768);
nor U13373 (N_13373,N_12235,N_12822);
xnor U13374 (N_13374,N_12356,N_12523);
nor U13375 (N_13375,N_12304,N_12148);
or U13376 (N_13376,N_12885,N_12528);
or U13377 (N_13377,N_12711,N_12921);
and U13378 (N_13378,N_12598,N_12362);
nor U13379 (N_13379,N_12483,N_12501);
and U13380 (N_13380,N_12261,N_12578);
nor U13381 (N_13381,N_12725,N_12914);
xnor U13382 (N_13382,N_12880,N_12710);
xnor U13383 (N_13383,N_12745,N_12257);
nand U13384 (N_13384,N_12391,N_12858);
xor U13385 (N_13385,N_12418,N_12380);
and U13386 (N_13386,N_12836,N_12607);
or U13387 (N_13387,N_12682,N_12049);
and U13388 (N_13388,N_12138,N_12756);
or U13389 (N_13389,N_12920,N_12464);
and U13390 (N_13390,N_12475,N_12910);
and U13391 (N_13391,N_12278,N_12224);
nor U13392 (N_13392,N_12507,N_12168);
and U13393 (N_13393,N_12044,N_12065);
nor U13394 (N_13394,N_12893,N_12216);
nor U13395 (N_13395,N_12478,N_12791);
xnor U13396 (N_13396,N_12185,N_12724);
nor U13397 (N_13397,N_12441,N_12179);
nor U13398 (N_13398,N_12432,N_12664);
nor U13399 (N_13399,N_12995,N_12435);
and U13400 (N_13400,N_12824,N_12617);
xnor U13401 (N_13401,N_12850,N_12011);
nand U13402 (N_13402,N_12965,N_12210);
and U13403 (N_13403,N_12366,N_12215);
nand U13404 (N_13404,N_12338,N_12398);
nor U13405 (N_13405,N_12254,N_12117);
xnor U13406 (N_13406,N_12406,N_12773);
and U13407 (N_13407,N_12737,N_12512);
nor U13408 (N_13408,N_12740,N_12315);
nand U13409 (N_13409,N_12517,N_12753);
or U13410 (N_13410,N_12632,N_12204);
and U13411 (N_13411,N_12446,N_12801);
or U13412 (N_13412,N_12012,N_12221);
and U13413 (N_13413,N_12009,N_12593);
xnor U13414 (N_13414,N_12729,N_12008);
or U13415 (N_13415,N_12669,N_12438);
xnor U13416 (N_13416,N_12352,N_12238);
or U13417 (N_13417,N_12638,N_12648);
xnor U13418 (N_13418,N_12890,N_12502);
nor U13419 (N_13419,N_12730,N_12045);
nand U13420 (N_13420,N_12382,N_12931);
or U13421 (N_13421,N_12944,N_12821);
nor U13422 (N_13422,N_12414,N_12341);
nor U13423 (N_13423,N_12399,N_12769);
nor U13424 (N_13424,N_12823,N_12405);
nand U13425 (N_13425,N_12140,N_12219);
or U13426 (N_13426,N_12767,N_12798);
nand U13427 (N_13427,N_12466,N_12383);
or U13428 (N_13428,N_12873,N_12169);
nor U13429 (N_13429,N_12536,N_12240);
and U13430 (N_13430,N_12655,N_12103);
nor U13431 (N_13431,N_12053,N_12325);
and U13432 (N_13432,N_12993,N_12077);
nor U13433 (N_13433,N_12392,N_12534);
and U13434 (N_13434,N_12006,N_12721);
nand U13435 (N_13435,N_12505,N_12623);
nand U13436 (N_13436,N_12270,N_12688);
nand U13437 (N_13437,N_12841,N_12895);
or U13438 (N_13438,N_12557,N_12106);
and U13439 (N_13439,N_12396,N_12720);
xnor U13440 (N_13440,N_12225,N_12461);
nor U13441 (N_13441,N_12694,N_12061);
or U13442 (N_13442,N_12830,N_12353);
xor U13443 (N_13443,N_12331,N_12652);
nand U13444 (N_13444,N_12457,N_12050);
nand U13445 (N_13445,N_12522,N_12273);
or U13446 (N_13446,N_12072,N_12040);
nor U13447 (N_13447,N_12279,N_12283);
and U13448 (N_13448,N_12787,N_12635);
xnor U13449 (N_13449,N_12524,N_12979);
xor U13450 (N_13450,N_12367,N_12913);
xor U13451 (N_13451,N_12310,N_12429);
or U13452 (N_13452,N_12384,N_12236);
and U13453 (N_13453,N_12508,N_12276);
or U13454 (N_13454,N_12859,N_12723);
and U13455 (N_13455,N_12144,N_12281);
nand U13456 (N_13456,N_12110,N_12495);
nor U13457 (N_13457,N_12644,N_12693);
nor U13458 (N_13458,N_12326,N_12537);
and U13459 (N_13459,N_12079,N_12280);
nand U13460 (N_13460,N_12319,N_12374);
xnor U13461 (N_13461,N_12174,N_12333);
xor U13462 (N_13462,N_12342,N_12243);
xnor U13463 (N_13463,N_12463,N_12407);
or U13464 (N_13464,N_12978,N_12892);
nor U13465 (N_13465,N_12456,N_12062);
xnor U13466 (N_13466,N_12176,N_12417);
and U13467 (N_13467,N_12165,N_12844);
xnor U13468 (N_13468,N_12129,N_12603);
and U13469 (N_13469,N_12904,N_12043);
and U13470 (N_13470,N_12001,N_12134);
nor U13471 (N_13471,N_12226,N_12123);
xnor U13472 (N_13472,N_12615,N_12000);
nor U13473 (N_13473,N_12948,N_12511);
nand U13474 (N_13474,N_12612,N_12788);
nand U13475 (N_13475,N_12340,N_12365);
xor U13476 (N_13476,N_12583,N_12158);
or U13477 (N_13477,N_12611,N_12480);
or U13478 (N_13478,N_12086,N_12750);
nor U13479 (N_13479,N_12731,N_12159);
and U13480 (N_13480,N_12555,N_12671);
and U13481 (N_13481,N_12156,N_12887);
and U13482 (N_13482,N_12211,N_12385);
and U13483 (N_13483,N_12198,N_12778);
and U13484 (N_13484,N_12871,N_12518);
xnor U13485 (N_13485,N_12620,N_12164);
xor U13486 (N_13486,N_12530,N_12020);
nand U13487 (N_13487,N_12812,N_12497);
xnor U13488 (N_13488,N_12941,N_12023);
nor U13489 (N_13489,N_12239,N_12113);
xor U13490 (N_13490,N_12817,N_12879);
nor U13491 (N_13491,N_12735,N_12619);
nor U13492 (N_13492,N_12606,N_12241);
nor U13493 (N_13493,N_12702,N_12604);
xnor U13494 (N_13494,N_12290,N_12187);
xnor U13495 (N_13495,N_12840,N_12733);
or U13496 (N_13496,N_12299,N_12448);
xor U13497 (N_13497,N_12958,N_12218);
or U13498 (N_13498,N_12267,N_12869);
nor U13499 (N_13499,N_12190,N_12102);
or U13500 (N_13500,N_12107,N_12707);
nand U13501 (N_13501,N_12403,N_12159);
xnor U13502 (N_13502,N_12439,N_12654);
or U13503 (N_13503,N_12408,N_12305);
nor U13504 (N_13504,N_12420,N_12752);
and U13505 (N_13505,N_12332,N_12980);
nor U13506 (N_13506,N_12124,N_12561);
xnor U13507 (N_13507,N_12460,N_12318);
nand U13508 (N_13508,N_12320,N_12847);
nor U13509 (N_13509,N_12821,N_12873);
xnor U13510 (N_13510,N_12626,N_12697);
nand U13511 (N_13511,N_12856,N_12697);
and U13512 (N_13512,N_12227,N_12100);
nand U13513 (N_13513,N_12989,N_12951);
and U13514 (N_13514,N_12010,N_12776);
or U13515 (N_13515,N_12280,N_12436);
xnor U13516 (N_13516,N_12891,N_12462);
and U13517 (N_13517,N_12932,N_12843);
and U13518 (N_13518,N_12195,N_12163);
nand U13519 (N_13519,N_12319,N_12066);
xor U13520 (N_13520,N_12996,N_12035);
nand U13521 (N_13521,N_12028,N_12793);
nand U13522 (N_13522,N_12551,N_12920);
and U13523 (N_13523,N_12211,N_12179);
nand U13524 (N_13524,N_12558,N_12830);
nor U13525 (N_13525,N_12601,N_12582);
nor U13526 (N_13526,N_12180,N_12289);
nor U13527 (N_13527,N_12506,N_12175);
nor U13528 (N_13528,N_12707,N_12920);
xor U13529 (N_13529,N_12286,N_12960);
or U13530 (N_13530,N_12657,N_12770);
nand U13531 (N_13531,N_12449,N_12024);
nand U13532 (N_13532,N_12158,N_12269);
nor U13533 (N_13533,N_12199,N_12744);
or U13534 (N_13534,N_12858,N_12572);
nand U13535 (N_13535,N_12945,N_12197);
or U13536 (N_13536,N_12527,N_12374);
or U13537 (N_13537,N_12712,N_12535);
nor U13538 (N_13538,N_12137,N_12516);
xor U13539 (N_13539,N_12537,N_12610);
nor U13540 (N_13540,N_12696,N_12134);
nor U13541 (N_13541,N_12022,N_12902);
nor U13542 (N_13542,N_12773,N_12181);
or U13543 (N_13543,N_12243,N_12624);
and U13544 (N_13544,N_12784,N_12213);
xnor U13545 (N_13545,N_12939,N_12532);
nor U13546 (N_13546,N_12911,N_12092);
xor U13547 (N_13547,N_12411,N_12471);
nand U13548 (N_13548,N_12936,N_12426);
or U13549 (N_13549,N_12129,N_12152);
and U13550 (N_13550,N_12550,N_12570);
nand U13551 (N_13551,N_12717,N_12053);
nand U13552 (N_13552,N_12656,N_12166);
nand U13553 (N_13553,N_12461,N_12891);
nor U13554 (N_13554,N_12199,N_12616);
or U13555 (N_13555,N_12092,N_12198);
and U13556 (N_13556,N_12648,N_12520);
and U13557 (N_13557,N_12812,N_12910);
and U13558 (N_13558,N_12113,N_12632);
or U13559 (N_13559,N_12536,N_12165);
and U13560 (N_13560,N_12762,N_12364);
nand U13561 (N_13561,N_12940,N_12814);
nand U13562 (N_13562,N_12648,N_12452);
or U13563 (N_13563,N_12024,N_12735);
xnor U13564 (N_13564,N_12329,N_12685);
or U13565 (N_13565,N_12602,N_12899);
and U13566 (N_13566,N_12225,N_12205);
and U13567 (N_13567,N_12439,N_12741);
and U13568 (N_13568,N_12829,N_12834);
and U13569 (N_13569,N_12869,N_12867);
nor U13570 (N_13570,N_12589,N_12993);
nor U13571 (N_13571,N_12880,N_12582);
xor U13572 (N_13572,N_12011,N_12660);
and U13573 (N_13573,N_12895,N_12437);
nor U13574 (N_13574,N_12165,N_12018);
nand U13575 (N_13575,N_12288,N_12220);
or U13576 (N_13576,N_12147,N_12619);
and U13577 (N_13577,N_12576,N_12717);
nor U13578 (N_13578,N_12265,N_12480);
or U13579 (N_13579,N_12961,N_12391);
or U13580 (N_13580,N_12964,N_12047);
xor U13581 (N_13581,N_12021,N_12998);
nor U13582 (N_13582,N_12726,N_12900);
and U13583 (N_13583,N_12170,N_12281);
and U13584 (N_13584,N_12356,N_12193);
and U13585 (N_13585,N_12216,N_12975);
or U13586 (N_13586,N_12602,N_12508);
nand U13587 (N_13587,N_12568,N_12918);
or U13588 (N_13588,N_12975,N_12031);
nand U13589 (N_13589,N_12415,N_12313);
or U13590 (N_13590,N_12872,N_12284);
nand U13591 (N_13591,N_12218,N_12397);
nand U13592 (N_13592,N_12872,N_12677);
and U13593 (N_13593,N_12109,N_12445);
nand U13594 (N_13594,N_12385,N_12836);
and U13595 (N_13595,N_12374,N_12534);
and U13596 (N_13596,N_12994,N_12672);
and U13597 (N_13597,N_12509,N_12712);
nand U13598 (N_13598,N_12850,N_12713);
and U13599 (N_13599,N_12209,N_12839);
nand U13600 (N_13600,N_12704,N_12793);
and U13601 (N_13601,N_12125,N_12292);
and U13602 (N_13602,N_12772,N_12699);
nor U13603 (N_13603,N_12618,N_12321);
nand U13604 (N_13604,N_12903,N_12730);
nor U13605 (N_13605,N_12463,N_12035);
nor U13606 (N_13606,N_12293,N_12976);
or U13607 (N_13607,N_12178,N_12758);
nor U13608 (N_13608,N_12309,N_12994);
or U13609 (N_13609,N_12067,N_12397);
nor U13610 (N_13610,N_12489,N_12915);
nand U13611 (N_13611,N_12556,N_12126);
nand U13612 (N_13612,N_12798,N_12006);
nand U13613 (N_13613,N_12355,N_12130);
nor U13614 (N_13614,N_12302,N_12431);
and U13615 (N_13615,N_12777,N_12990);
nor U13616 (N_13616,N_12623,N_12846);
and U13617 (N_13617,N_12685,N_12149);
or U13618 (N_13618,N_12198,N_12854);
xor U13619 (N_13619,N_12957,N_12001);
xnor U13620 (N_13620,N_12615,N_12176);
and U13621 (N_13621,N_12167,N_12535);
and U13622 (N_13622,N_12080,N_12768);
xnor U13623 (N_13623,N_12988,N_12929);
or U13624 (N_13624,N_12923,N_12184);
and U13625 (N_13625,N_12857,N_12218);
or U13626 (N_13626,N_12683,N_12080);
nand U13627 (N_13627,N_12349,N_12111);
and U13628 (N_13628,N_12514,N_12251);
or U13629 (N_13629,N_12649,N_12947);
xor U13630 (N_13630,N_12823,N_12933);
or U13631 (N_13631,N_12192,N_12151);
nand U13632 (N_13632,N_12146,N_12492);
and U13633 (N_13633,N_12210,N_12525);
nand U13634 (N_13634,N_12546,N_12812);
xor U13635 (N_13635,N_12380,N_12826);
nor U13636 (N_13636,N_12377,N_12954);
nand U13637 (N_13637,N_12243,N_12871);
nand U13638 (N_13638,N_12664,N_12167);
nand U13639 (N_13639,N_12153,N_12732);
and U13640 (N_13640,N_12074,N_12411);
nor U13641 (N_13641,N_12497,N_12818);
nor U13642 (N_13642,N_12376,N_12440);
and U13643 (N_13643,N_12078,N_12414);
or U13644 (N_13644,N_12809,N_12933);
nor U13645 (N_13645,N_12453,N_12293);
nor U13646 (N_13646,N_12035,N_12921);
nand U13647 (N_13647,N_12163,N_12843);
nor U13648 (N_13648,N_12943,N_12770);
xnor U13649 (N_13649,N_12683,N_12726);
or U13650 (N_13650,N_12056,N_12913);
nand U13651 (N_13651,N_12167,N_12397);
xor U13652 (N_13652,N_12901,N_12067);
or U13653 (N_13653,N_12929,N_12011);
xor U13654 (N_13654,N_12002,N_12150);
xnor U13655 (N_13655,N_12111,N_12234);
and U13656 (N_13656,N_12717,N_12981);
nor U13657 (N_13657,N_12299,N_12654);
or U13658 (N_13658,N_12612,N_12493);
and U13659 (N_13659,N_12821,N_12510);
or U13660 (N_13660,N_12860,N_12866);
nor U13661 (N_13661,N_12669,N_12915);
nand U13662 (N_13662,N_12973,N_12117);
nand U13663 (N_13663,N_12743,N_12852);
or U13664 (N_13664,N_12336,N_12652);
xnor U13665 (N_13665,N_12071,N_12002);
nor U13666 (N_13666,N_12570,N_12552);
or U13667 (N_13667,N_12689,N_12972);
xor U13668 (N_13668,N_12042,N_12162);
nor U13669 (N_13669,N_12023,N_12109);
and U13670 (N_13670,N_12614,N_12475);
and U13671 (N_13671,N_12584,N_12657);
nand U13672 (N_13672,N_12370,N_12595);
or U13673 (N_13673,N_12046,N_12709);
xor U13674 (N_13674,N_12126,N_12065);
or U13675 (N_13675,N_12767,N_12303);
xnor U13676 (N_13676,N_12593,N_12479);
and U13677 (N_13677,N_12487,N_12363);
and U13678 (N_13678,N_12337,N_12257);
nand U13679 (N_13679,N_12427,N_12581);
nor U13680 (N_13680,N_12927,N_12488);
and U13681 (N_13681,N_12134,N_12224);
nand U13682 (N_13682,N_12137,N_12257);
or U13683 (N_13683,N_12508,N_12563);
and U13684 (N_13684,N_12931,N_12742);
and U13685 (N_13685,N_12979,N_12743);
and U13686 (N_13686,N_12400,N_12083);
nand U13687 (N_13687,N_12995,N_12756);
nand U13688 (N_13688,N_12508,N_12323);
xnor U13689 (N_13689,N_12429,N_12464);
nand U13690 (N_13690,N_12878,N_12991);
xor U13691 (N_13691,N_12084,N_12867);
nor U13692 (N_13692,N_12482,N_12774);
xnor U13693 (N_13693,N_12332,N_12931);
nand U13694 (N_13694,N_12261,N_12416);
nand U13695 (N_13695,N_12153,N_12386);
and U13696 (N_13696,N_12094,N_12161);
nor U13697 (N_13697,N_12155,N_12725);
and U13698 (N_13698,N_12609,N_12253);
nor U13699 (N_13699,N_12164,N_12485);
xnor U13700 (N_13700,N_12978,N_12077);
nand U13701 (N_13701,N_12542,N_12862);
nand U13702 (N_13702,N_12916,N_12064);
or U13703 (N_13703,N_12905,N_12076);
nor U13704 (N_13704,N_12629,N_12784);
and U13705 (N_13705,N_12481,N_12108);
nand U13706 (N_13706,N_12382,N_12663);
and U13707 (N_13707,N_12814,N_12545);
xnor U13708 (N_13708,N_12110,N_12724);
nand U13709 (N_13709,N_12682,N_12222);
or U13710 (N_13710,N_12577,N_12587);
or U13711 (N_13711,N_12127,N_12358);
xnor U13712 (N_13712,N_12178,N_12797);
nor U13713 (N_13713,N_12608,N_12709);
and U13714 (N_13714,N_12654,N_12762);
xor U13715 (N_13715,N_12519,N_12716);
nand U13716 (N_13716,N_12852,N_12761);
xor U13717 (N_13717,N_12822,N_12724);
or U13718 (N_13718,N_12652,N_12028);
nor U13719 (N_13719,N_12967,N_12177);
xnor U13720 (N_13720,N_12846,N_12637);
xnor U13721 (N_13721,N_12354,N_12233);
xnor U13722 (N_13722,N_12005,N_12140);
nand U13723 (N_13723,N_12116,N_12904);
nand U13724 (N_13724,N_12681,N_12061);
and U13725 (N_13725,N_12436,N_12275);
or U13726 (N_13726,N_12487,N_12506);
xnor U13727 (N_13727,N_12034,N_12591);
xor U13728 (N_13728,N_12508,N_12346);
nor U13729 (N_13729,N_12634,N_12909);
nor U13730 (N_13730,N_12802,N_12139);
nand U13731 (N_13731,N_12756,N_12783);
xnor U13732 (N_13732,N_12022,N_12634);
nand U13733 (N_13733,N_12998,N_12959);
nand U13734 (N_13734,N_12517,N_12003);
xor U13735 (N_13735,N_12526,N_12893);
xor U13736 (N_13736,N_12088,N_12972);
nor U13737 (N_13737,N_12108,N_12671);
or U13738 (N_13738,N_12793,N_12950);
nor U13739 (N_13739,N_12807,N_12940);
nor U13740 (N_13740,N_12706,N_12529);
and U13741 (N_13741,N_12926,N_12130);
and U13742 (N_13742,N_12093,N_12498);
xnor U13743 (N_13743,N_12070,N_12986);
nor U13744 (N_13744,N_12052,N_12258);
or U13745 (N_13745,N_12317,N_12177);
and U13746 (N_13746,N_12283,N_12079);
xor U13747 (N_13747,N_12366,N_12805);
or U13748 (N_13748,N_12751,N_12562);
nor U13749 (N_13749,N_12368,N_12256);
xnor U13750 (N_13750,N_12756,N_12708);
or U13751 (N_13751,N_12718,N_12099);
xnor U13752 (N_13752,N_12433,N_12709);
nand U13753 (N_13753,N_12805,N_12989);
nand U13754 (N_13754,N_12857,N_12462);
nand U13755 (N_13755,N_12291,N_12666);
xor U13756 (N_13756,N_12135,N_12252);
nor U13757 (N_13757,N_12920,N_12445);
nor U13758 (N_13758,N_12396,N_12997);
or U13759 (N_13759,N_12369,N_12613);
or U13760 (N_13760,N_12086,N_12709);
nor U13761 (N_13761,N_12046,N_12731);
nor U13762 (N_13762,N_12266,N_12052);
and U13763 (N_13763,N_12067,N_12781);
xnor U13764 (N_13764,N_12272,N_12340);
nand U13765 (N_13765,N_12546,N_12908);
and U13766 (N_13766,N_12434,N_12155);
or U13767 (N_13767,N_12013,N_12983);
and U13768 (N_13768,N_12707,N_12651);
xor U13769 (N_13769,N_12564,N_12974);
and U13770 (N_13770,N_12069,N_12929);
xnor U13771 (N_13771,N_12343,N_12541);
and U13772 (N_13772,N_12377,N_12735);
nand U13773 (N_13773,N_12418,N_12193);
nand U13774 (N_13774,N_12562,N_12222);
nor U13775 (N_13775,N_12985,N_12317);
or U13776 (N_13776,N_12023,N_12090);
nand U13777 (N_13777,N_12510,N_12425);
nand U13778 (N_13778,N_12330,N_12427);
nor U13779 (N_13779,N_12157,N_12009);
xor U13780 (N_13780,N_12512,N_12736);
nand U13781 (N_13781,N_12927,N_12275);
nor U13782 (N_13782,N_12827,N_12555);
and U13783 (N_13783,N_12878,N_12497);
nor U13784 (N_13784,N_12486,N_12846);
nand U13785 (N_13785,N_12193,N_12242);
nor U13786 (N_13786,N_12408,N_12734);
and U13787 (N_13787,N_12928,N_12394);
and U13788 (N_13788,N_12296,N_12484);
nor U13789 (N_13789,N_12227,N_12437);
nand U13790 (N_13790,N_12032,N_12079);
xor U13791 (N_13791,N_12083,N_12950);
and U13792 (N_13792,N_12896,N_12422);
xor U13793 (N_13793,N_12069,N_12358);
nor U13794 (N_13794,N_12012,N_12672);
nand U13795 (N_13795,N_12168,N_12375);
nor U13796 (N_13796,N_12462,N_12585);
xor U13797 (N_13797,N_12617,N_12235);
or U13798 (N_13798,N_12294,N_12829);
or U13799 (N_13799,N_12469,N_12148);
nand U13800 (N_13800,N_12136,N_12650);
and U13801 (N_13801,N_12859,N_12377);
nor U13802 (N_13802,N_12607,N_12179);
and U13803 (N_13803,N_12347,N_12552);
or U13804 (N_13804,N_12669,N_12546);
and U13805 (N_13805,N_12817,N_12832);
or U13806 (N_13806,N_12647,N_12321);
and U13807 (N_13807,N_12746,N_12605);
xnor U13808 (N_13808,N_12324,N_12756);
xor U13809 (N_13809,N_12016,N_12853);
and U13810 (N_13810,N_12710,N_12385);
nor U13811 (N_13811,N_12731,N_12066);
or U13812 (N_13812,N_12833,N_12661);
or U13813 (N_13813,N_12429,N_12423);
nor U13814 (N_13814,N_12706,N_12843);
and U13815 (N_13815,N_12389,N_12266);
nand U13816 (N_13816,N_12129,N_12725);
and U13817 (N_13817,N_12097,N_12988);
nor U13818 (N_13818,N_12067,N_12850);
nand U13819 (N_13819,N_12754,N_12316);
or U13820 (N_13820,N_12280,N_12285);
nor U13821 (N_13821,N_12628,N_12224);
nand U13822 (N_13822,N_12007,N_12706);
or U13823 (N_13823,N_12787,N_12806);
nand U13824 (N_13824,N_12071,N_12192);
and U13825 (N_13825,N_12765,N_12471);
and U13826 (N_13826,N_12374,N_12245);
xnor U13827 (N_13827,N_12946,N_12728);
xnor U13828 (N_13828,N_12641,N_12809);
xor U13829 (N_13829,N_12181,N_12978);
or U13830 (N_13830,N_12047,N_12641);
and U13831 (N_13831,N_12376,N_12577);
and U13832 (N_13832,N_12113,N_12153);
xnor U13833 (N_13833,N_12389,N_12126);
and U13834 (N_13834,N_12127,N_12065);
or U13835 (N_13835,N_12532,N_12400);
or U13836 (N_13836,N_12623,N_12888);
nand U13837 (N_13837,N_12282,N_12176);
nor U13838 (N_13838,N_12964,N_12733);
nor U13839 (N_13839,N_12433,N_12047);
and U13840 (N_13840,N_12088,N_12014);
nand U13841 (N_13841,N_12592,N_12776);
nand U13842 (N_13842,N_12386,N_12711);
nand U13843 (N_13843,N_12722,N_12235);
and U13844 (N_13844,N_12766,N_12104);
nand U13845 (N_13845,N_12305,N_12124);
and U13846 (N_13846,N_12071,N_12518);
nand U13847 (N_13847,N_12910,N_12082);
xnor U13848 (N_13848,N_12154,N_12409);
nor U13849 (N_13849,N_12166,N_12657);
xor U13850 (N_13850,N_12514,N_12180);
nor U13851 (N_13851,N_12997,N_12294);
and U13852 (N_13852,N_12520,N_12293);
nor U13853 (N_13853,N_12642,N_12707);
xor U13854 (N_13854,N_12102,N_12281);
nand U13855 (N_13855,N_12461,N_12426);
and U13856 (N_13856,N_12907,N_12308);
nor U13857 (N_13857,N_12516,N_12020);
and U13858 (N_13858,N_12095,N_12806);
or U13859 (N_13859,N_12488,N_12671);
nor U13860 (N_13860,N_12166,N_12247);
and U13861 (N_13861,N_12785,N_12059);
nor U13862 (N_13862,N_12198,N_12649);
and U13863 (N_13863,N_12989,N_12866);
and U13864 (N_13864,N_12771,N_12001);
nor U13865 (N_13865,N_12988,N_12238);
xnor U13866 (N_13866,N_12871,N_12070);
nor U13867 (N_13867,N_12374,N_12986);
xnor U13868 (N_13868,N_12635,N_12903);
xnor U13869 (N_13869,N_12818,N_12907);
and U13870 (N_13870,N_12478,N_12099);
xor U13871 (N_13871,N_12648,N_12458);
xnor U13872 (N_13872,N_12282,N_12167);
or U13873 (N_13873,N_12103,N_12532);
and U13874 (N_13874,N_12420,N_12610);
and U13875 (N_13875,N_12657,N_12755);
nand U13876 (N_13876,N_12204,N_12996);
nand U13877 (N_13877,N_12288,N_12161);
or U13878 (N_13878,N_12354,N_12740);
nand U13879 (N_13879,N_12900,N_12983);
xor U13880 (N_13880,N_12365,N_12960);
or U13881 (N_13881,N_12078,N_12380);
nor U13882 (N_13882,N_12927,N_12108);
or U13883 (N_13883,N_12663,N_12568);
or U13884 (N_13884,N_12273,N_12209);
and U13885 (N_13885,N_12806,N_12524);
nor U13886 (N_13886,N_12595,N_12799);
or U13887 (N_13887,N_12296,N_12840);
and U13888 (N_13888,N_12821,N_12364);
nor U13889 (N_13889,N_12485,N_12967);
nor U13890 (N_13890,N_12060,N_12150);
xor U13891 (N_13891,N_12225,N_12485);
nor U13892 (N_13892,N_12729,N_12318);
or U13893 (N_13893,N_12043,N_12053);
nor U13894 (N_13894,N_12076,N_12957);
or U13895 (N_13895,N_12886,N_12643);
or U13896 (N_13896,N_12927,N_12594);
nor U13897 (N_13897,N_12289,N_12189);
or U13898 (N_13898,N_12399,N_12824);
nor U13899 (N_13899,N_12622,N_12612);
nand U13900 (N_13900,N_12929,N_12342);
nand U13901 (N_13901,N_12291,N_12457);
and U13902 (N_13902,N_12592,N_12828);
nand U13903 (N_13903,N_12628,N_12491);
and U13904 (N_13904,N_12651,N_12118);
nor U13905 (N_13905,N_12948,N_12482);
nor U13906 (N_13906,N_12083,N_12866);
and U13907 (N_13907,N_12375,N_12746);
nor U13908 (N_13908,N_12440,N_12026);
xor U13909 (N_13909,N_12179,N_12400);
nor U13910 (N_13910,N_12112,N_12703);
or U13911 (N_13911,N_12266,N_12873);
xor U13912 (N_13912,N_12882,N_12379);
xnor U13913 (N_13913,N_12622,N_12309);
nor U13914 (N_13914,N_12509,N_12692);
nor U13915 (N_13915,N_12566,N_12528);
nand U13916 (N_13916,N_12096,N_12341);
nor U13917 (N_13917,N_12359,N_12629);
nand U13918 (N_13918,N_12722,N_12200);
nand U13919 (N_13919,N_12192,N_12671);
nor U13920 (N_13920,N_12211,N_12842);
xor U13921 (N_13921,N_12395,N_12416);
nand U13922 (N_13922,N_12318,N_12517);
and U13923 (N_13923,N_12829,N_12788);
nor U13924 (N_13924,N_12754,N_12243);
nand U13925 (N_13925,N_12022,N_12339);
xnor U13926 (N_13926,N_12426,N_12205);
xnor U13927 (N_13927,N_12189,N_12886);
xnor U13928 (N_13928,N_12718,N_12863);
xnor U13929 (N_13929,N_12508,N_12080);
or U13930 (N_13930,N_12287,N_12487);
and U13931 (N_13931,N_12694,N_12322);
nor U13932 (N_13932,N_12622,N_12040);
or U13933 (N_13933,N_12106,N_12714);
xnor U13934 (N_13934,N_12425,N_12133);
or U13935 (N_13935,N_12864,N_12881);
nand U13936 (N_13936,N_12113,N_12229);
nand U13937 (N_13937,N_12229,N_12570);
and U13938 (N_13938,N_12508,N_12955);
or U13939 (N_13939,N_12859,N_12237);
and U13940 (N_13940,N_12228,N_12575);
and U13941 (N_13941,N_12904,N_12710);
xor U13942 (N_13942,N_12620,N_12909);
or U13943 (N_13943,N_12089,N_12173);
and U13944 (N_13944,N_12939,N_12844);
nor U13945 (N_13945,N_12801,N_12105);
xor U13946 (N_13946,N_12585,N_12773);
xor U13947 (N_13947,N_12931,N_12494);
and U13948 (N_13948,N_12057,N_12086);
and U13949 (N_13949,N_12705,N_12228);
and U13950 (N_13950,N_12088,N_12010);
and U13951 (N_13951,N_12707,N_12719);
nor U13952 (N_13952,N_12264,N_12412);
xor U13953 (N_13953,N_12508,N_12159);
xnor U13954 (N_13954,N_12709,N_12737);
nand U13955 (N_13955,N_12704,N_12075);
or U13956 (N_13956,N_12614,N_12959);
nor U13957 (N_13957,N_12219,N_12539);
nor U13958 (N_13958,N_12072,N_12071);
nor U13959 (N_13959,N_12936,N_12630);
or U13960 (N_13960,N_12021,N_12418);
and U13961 (N_13961,N_12513,N_12607);
xor U13962 (N_13962,N_12408,N_12321);
nor U13963 (N_13963,N_12694,N_12092);
or U13964 (N_13964,N_12694,N_12661);
xnor U13965 (N_13965,N_12698,N_12420);
xnor U13966 (N_13966,N_12480,N_12786);
and U13967 (N_13967,N_12673,N_12567);
nor U13968 (N_13968,N_12758,N_12546);
nor U13969 (N_13969,N_12384,N_12357);
nor U13970 (N_13970,N_12930,N_12090);
nor U13971 (N_13971,N_12697,N_12896);
or U13972 (N_13972,N_12715,N_12018);
nor U13973 (N_13973,N_12363,N_12386);
nor U13974 (N_13974,N_12973,N_12110);
nand U13975 (N_13975,N_12373,N_12941);
and U13976 (N_13976,N_12133,N_12792);
xnor U13977 (N_13977,N_12651,N_12687);
and U13978 (N_13978,N_12588,N_12475);
nor U13979 (N_13979,N_12364,N_12713);
xnor U13980 (N_13980,N_12985,N_12923);
and U13981 (N_13981,N_12096,N_12172);
nand U13982 (N_13982,N_12485,N_12318);
and U13983 (N_13983,N_12420,N_12441);
nand U13984 (N_13984,N_12106,N_12343);
or U13985 (N_13985,N_12047,N_12175);
xnor U13986 (N_13986,N_12604,N_12945);
xnor U13987 (N_13987,N_12189,N_12772);
xor U13988 (N_13988,N_12878,N_12782);
or U13989 (N_13989,N_12278,N_12543);
nand U13990 (N_13990,N_12294,N_12760);
or U13991 (N_13991,N_12709,N_12702);
nand U13992 (N_13992,N_12715,N_12708);
xnor U13993 (N_13993,N_12624,N_12779);
nor U13994 (N_13994,N_12295,N_12893);
xnor U13995 (N_13995,N_12877,N_12802);
or U13996 (N_13996,N_12874,N_12638);
nor U13997 (N_13997,N_12604,N_12562);
or U13998 (N_13998,N_12580,N_12269);
xnor U13999 (N_13999,N_12946,N_12240);
nor U14000 (N_14000,N_13861,N_13003);
nand U14001 (N_14001,N_13234,N_13675);
and U14002 (N_14002,N_13777,N_13493);
or U14003 (N_14003,N_13524,N_13960);
or U14004 (N_14004,N_13448,N_13324);
and U14005 (N_14005,N_13195,N_13866);
nor U14006 (N_14006,N_13564,N_13798);
xnor U14007 (N_14007,N_13659,N_13562);
nand U14008 (N_14008,N_13671,N_13552);
or U14009 (N_14009,N_13905,N_13949);
nand U14010 (N_14010,N_13953,N_13150);
and U14011 (N_14011,N_13964,N_13840);
nor U14012 (N_14012,N_13826,N_13471);
or U14013 (N_14013,N_13287,N_13405);
xnor U14014 (N_14014,N_13460,N_13321);
and U14015 (N_14015,N_13505,N_13213);
xnor U14016 (N_14016,N_13096,N_13909);
or U14017 (N_14017,N_13323,N_13898);
xnor U14018 (N_14018,N_13453,N_13247);
xor U14019 (N_14019,N_13259,N_13383);
nand U14020 (N_14020,N_13480,N_13972);
nor U14021 (N_14021,N_13119,N_13982);
nor U14022 (N_14022,N_13248,N_13832);
or U14023 (N_14023,N_13373,N_13482);
nor U14024 (N_14024,N_13961,N_13369);
or U14025 (N_14025,N_13151,N_13437);
xnor U14026 (N_14026,N_13956,N_13584);
xnor U14027 (N_14027,N_13566,N_13245);
nor U14028 (N_14028,N_13220,N_13520);
xor U14029 (N_14029,N_13468,N_13175);
and U14030 (N_14030,N_13320,N_13143);
and U14031 (N_14031,N_13906,N_13488);
or U14032 (N_14032,N_13241,N_13454);
and U14033 (N_14033,N_13262,N_13058);
and U14034 (N_14034,N_13492,N_13318);
or U14035 (N_14035,N_13180,N_13276);
or U14036 (N_14036,N_13108,N_13878);
nor U14037 (N_14037,N_13066,N_13963);
nand U14038 (N_14038,N_13715,N_13749);
and U14039 (N_14039,N_13186,N_13499);
xor U14040 (N_14040,N_13500,N_13424);
nand U14041 (N_14041,N_13966,N_13796);
nand U14042 (N_14042,N_13289,N_13126);
nand U14043 (N_14043,N_13490,N_13090);
xnor U14044 (N_14044,N_13112,N_13589);
or U14045 (N_14045,N_13804,N_13106);
and U14046 (N_14046,N_13604,N_13617);
nand U14047 (N_14047,N_13585,N_13809);
and U14048 (N_14048,N_13219,N_13797);
or U14049 (N_14049,N_13027,N_13434);
and U14050 (N_14050,N_13231,N_13355);
and U14051 (N_14051,N_13147,N_13372);
nand U14052 (N_14052,N_13496,N_13050);
nand U14053 (N_14053,N_13279,N_13770);
nand U14054 (N_14054,N_13733,N_13620);
nand U14055 (N_14055,N_13999,N_13013);
nor U14056 (N_14056,N_13548,N_13421);
nand U14057 (N_14057,N_13667,N_13033);
and U14058 (N_14058,N_13135,N_13529);
and U14059 (N_14059,N_13484,N_13943);
or U14060 (N_14060,N_13332,N_13427);
or U14061 (N_14061,N_13154,N_13461);
and U14062 (N_14062,N_13489,N_13860);
and U14063 (N_14063,N_13581,N_13225);
nand U14064 (N_14064,N_13140,N_13854);
or U14065 (N_14065,N_13300,N_13517);
xor U14066 (N_14066,N_13311,N_13212);
xor U14067 (N_14067,N_13766,N_13737);
xor U14068 (N_14068,N_13270,N_13178);
xnor U14069 (N_14069,N_13167,N_13590);
xnor U14070 (N_14070,N_13385,N_13346);
nor U14071 (N_14071,N_13726,N_13052);
nor U14072 (N_14072,N_13142,N_13165);
nand U14073 (N_14073,N_13221,N_13911);
nor U14074 (N_14074,N_13296,N_13538);
nor U14075 (N_14075,N_13012,N_13215);
nor U14076 (N_14076,N_13095,N_13417);
and U14077 (N_14077,N_13418,N_13670);
and U14078 (N_14078,N_13145,N_13301);
or U14079 (N_14079,N_13049,N_13759);
and U14080 (N_14080,N_13674,N_13720);
and U14081 (N_14081,N_13101,N_13694);
xnor U14082 (N_14082,N_13558,N_13088);
and U14083 (N_14083,N_13341,N_13556);
nand U14084 (N_14084,N_13495,N_13873);
and U14085 (N_14085,N_13696,N_13371);
and U14086 (N_14086,N_13985,N_13362);
nor U14087 (N_14087,N_13206,N_13312);
nand U14088 (N_14088,N_13356,N_13450);
nand U14089 (N_14089,N_13907,N_13638);
nor U14090 (N_14090,N_13286,N_13885);
xnor U14091 (N_14091,N_13244,N_13864);
and U14092 (N_14092,N_13543,N_13920);
nand U14093 (N_14093,N_13429,N_13926);
xnor U14094 (N_14094,N_13216,N_13077);
or U14095 (N_14095,N_13904,N_13394);
or U14096 (N_14096,N_13990,N_13193);
nand U14097 (N_14097,N_13516,N_13745);
xor U14098 (N_14098,N_13473,N_13577);
or U14099 (N_14099,N_13582,N_13007);
and U14100 (N_14100,N_13570,N_13204);
or U14101 (N_14101,N_13645,N_13340);
and U14102 (N_14102,N_13343,N_13021);
nor U14103 (N_14103,N_13650,N_13104);
and U14104 (N_14104,N_13326,N_13747);
nand U14105 (N_14105,N_13616,N_13807);
xnor U14106 (N_14106,N_13536,N_13941);
nor U14107 (N_14107,N_13974,N_13451);
nand U14108 (N_14108,N_13310,N_13704);
xor U14109 (N_14109,N_13821,N_13842);
nor U14110 (N_14110,N_13271,N_13462);
and U14111 (N_14111,N_13267,N_13419);
nor U14112 (N_14112,N_13976,N_13081);
and U14113 (N_14113,N_13389,N_13580);
nor U14114 (N_14114,N_13849,N_13883);
and U14115 (N_14115,N_13181,N_13565);
nor U14116 (N_14116,N_13728,N_13572);
and U14117 (N_14117,N_13541,N_13786);
or U14118 (N_14118,N_13975,N_13060);
or U14119 (N_14119,N_13933,N_13381);
nand U14120 (N_14120,N_13086,N_13993);
nand U14121 (N_14121,N_13386,N_13350);
xor U14122 (N_14122,N_13601,N_13593);
nand U14123 (N_14123,N_13712,N_13399);
or U14124 (N_14124,N_13535,N_13518);
nand U14125 (N_14125,N_13606,N_13138);
and U14126 (N_14126,N_13335,N_13962);
nand U14127 (N_14127,N_13455,N_13452);
xnor U14128 (N_14128,N_13504,N_13360);
and U14129 (N_14129,N_13398,N_13896);
nor U14130 (N_14130,N_13018,N_13487);
or U14131 (N_14131,N_13931,N_13872);
or U14132 (N_14132,N_13633,N_13478);
nand U14133 (N_14133,N_13641,N_13583);
or U14134 (N_14134,N_13020,N_13765);
nor U14135 (N_14135,N_13843,N_13830);
or U14136 (N_14136,N_13829,N_13844);
and U14137 (N_14137,N_13724,N_13578);
xnor U14138 (N_14138,N_13874,N_13875);
nand U14139 (N_14139,N_13137,N_13592);
and U14140 (N_14140,N_13711,N_13025);
and U14141 (N_14141,N_13261,N_13795);
or U14142 (N_14142,N_13443,N_13576);
or U14143 (N_14143,N_13550,N_13182);
and U14144 (N_14144,N_13121,N_13857);
nor U14145 (N_14145,N_13512,N_13788);
or U14146 (N_14146,N_13258,N_13059);
or U14147 (N_14147,N_13763,N_13422);
nor U14148 (N_14148,N_13100,N_13139);
and U14149 (N_14149,N_13651,N_13841);
or U14150 (N_14150,N_13599,N_13984);
or U14151 (N_14151,N_13436,N_13255);
xnor U14152 (N_14152,N_13103,N_13377);
and U14153 (N_14153,N_13664,N_13586);
nand U14154 (N_14154,N_13054,N_13122);
nand U14155 (N_14155,N_13407,N_13291);
xor U14156 (N_14156,N_13277,N_13769);
or U14157 (N_14157,N_13530,N_13363);
nor U14158 (N_14158,N_13000,N_13663);
or U14159 (N_14159,N_13727,N_13092);
nor U14160 (N_14160,N_13294,N_13380);
nand U14161 (N_14161,N_13004,N_13605);
and U14162 (N_14162,N_13329,N_13331);
or U14163 (N_14163,N_13858,N_13129);
nand U14164 (N_14164,N_13432,N_13622);
and U14165 (N_14165,N_13184,N_13131);
nand U14166 (N_14166,N_13867,N_13703);
or U14167 (N_14167,N_13315,N_13925);
nand U14168 (N_14168,N_13705,N_13992);
and U14169 (N_14169,N_13177,N_13947);
xor U14170 (N_14170,N_13944,N_13912);
nor U14171 (N_14171,N_13037,N_13814);
xnor U14172 (N_14172,N_13702,N_13024);
or U14173 (N_14173,N_13902,N_13116);
or U14174 (N_14174,N_13387,N_13044);
and U14175 (N_14175,N_13416,N_13236);
nor U14176 (N_14176,N_13476,N_13411);
nand U14177 (N_14177,N_13549,N_13806);
nand U14178 (N_14178,N_13540,N_13901);
or U14179 (N_14179,N_13313,N_13034);
or U14180 (N_14180,N_13611,N_13945);
xor U14181 (N_14181,N_13148,N_13657);
and U14182 (N_14182,N_13010,N_13032);
xnor U14183 (N_14183,N_13397,N_13899);
nor U14184 (N_14184,N_13268,N_13412);
nor U14185 (N_14185,N_13113,N_13850);
or U14186 (N_14186,N_13061,N_13205);
or U14187 (N_14187,N_13774,N_13345);
or U14188 (N_14188,N_13779,N_13439);
or U14189 (N_14189,N_13102,N_13075);
nand U14190 (N_14190,N_13557,N_13198);
nor U14191 (N_14191,N_13753,N_13097);
nand U14192 (N_14192,N_13751,N_13272);
and U14193 (N_14193,N_13924,N_13227);
xor U14194 (N_14194,N_13413,N_13870);
xor U14195 (N_14195,N_13787,N_13950);
nor U14196 (N_14196,N_13615,N_13008);
nor U14197 (N_14197,N_13598,N_13158);
and U14198 (N_14198,N_13414,N_13353);
nand U14199 (N_14199,N_13063,N_13574);
xor U14200 (N_14200,N_13402,N_13133);
or U14201 (N_14201,N_13977,N_13299);
xnor U14202 (N_14202,N_13477,N_13815);
xnor U14203 (N_14203,N_13430,N_13731);
nor U14204 (N_14204,N_13269,N_13141);
nor U14205 (N_14205,N_13783,N_13991);
nand U14206 (N_14206,N_13338,N_13845);
and U14207 (N_14207,N_13660,N_13082);
nand U14208 (N_14208,N_13036,N_13594);
and U14209 (N_14209,N_13794,N_13253);
nand U14210 (N_14210,N_13005,N_13201);
and U14211 (N_14211,N_13967,N_13202);
nor U14212 (N_14212,N_13958,N_13456);
and U14213 (N_14213,N_13676,N_13629);
and U14214 (N_14214,N_13936,N_13502);
and U14215 (N_14215,N_13995,N_13656);
or U14216 (N_14216,N_13742,N_13981);
or U14217 (N_14217,N_13072,N_13773);
and U14218 (N_14218,N_13908,N_13445);
nand U14219 (N_14219,N_13831,N_13740);
nand U14220 (N_14220,N_13406,N_13128);
and U14221 (N_14221,N_13374,N_13232);
and U14222 (N_14222,N_13681,N_13325);
nand U14223 (N_14223,N_13756,N_13628);
nand U14224 (N_14224,N_13643,N_13819);
nand U14225 (N_14225,N_13297,N_13144);
or U14226 (N_14226,N_13280,N_13725);
or U14227 (N_14227,N_13486,N_13458);
nand U14228 (N_14228,N_13852,N_13959);
nand U14229 (N_14229,N_13812,N_13636);
and U14230 (N_14230,N_13662,N_13706);
nand U14231 (N_14231,N_13686,N_13230);
and U14232 (N_14232,N_13192,N_13107);
nand U14233 (N_14233,N_13306,N_13683);
nor U14234 (N_14234,N_13479,N_13400);
and U14235 (N_14235,N_13501,N_13120);
xnor U14236 (N_14236,N_13188,N_13185);
nor U14237 (N_14237,N_13546,N_13624);
and U14238 (N_14238,N_13067,N_13149);
xor U14239 (N_14239,N_13778,N_13545);
nand U14240 (N_14240,N_13134,N_13687);
nor U14241 (N_14241,N_13275,N_13038);
nor U14242 (N_14242,N_13989,N_13612);
nor U14243 (N_14243,N_13894,N_13068);
or U14244 (N_14244,N_13080,N_13547);
nor U14245 (N_14245,N_13940,N_13314);
nand U14246 (N_14246,N_13093,N_13403);
or U14247 (N_14247,N_13738,N_13065);
nor U14248 (N_14248,N_13257,N_13876);
or U14249 (N_14249,N_13045,N_13240);
xnor U14250 (N_14250,N_13285,N_13146);
xor U14251 (N_14251,N_13483,N_13560);
and U14252 (N_14252,N_13089,N_13707);
nand U14253 (N_14253,N_13169,N_13877);
or U14254 (N_14254,N_13197,N_13746);
and U14255 (N_14255,N_13587,N_13893);
or U14256 (N_14256,N_13954,N_13238);
and U14257 (N_14257,N_13474,N_13309);
or U14258 (N_14258,N_13039,N_13689);
nand U14259 (N_14259,N_13695,N_13591);
xnor U14260 (N_14260,N_13189,N_13988);
nor U14261 (N_14261,N_13115,N_13457);
nand U14262 (N_14262,N_13079,N_13459);
nor U14263 (N_14263,N_13428,N_13750);
nor U14264 (N_14264,N_13827,N_13714);
nand U14265 (N_14265,N_13709,N_13948);
xor U14266 (N_14266,N_13031,N_13521);
nor U14267 (N_14267,N_13191,N_13523);
and U14268 (N_14268,N_13918,N_13528);
nand U14269 (N_14269,N_13994,N_13979);
and U14270 (N_14270,N_13359,N_13503);
nand U14271 (N_14271,N_13009,N_13304);
nor U14272 (N_14272,N_13697,N_13218);
xor U14273 (N_14273,N_13465,N_13250);
nand U14274 (N_14274,N_13915,N_13895);
and U14275 (N_14275,N_13357,N_13235);
and U14276 (N_14276,N_13161,N_13342);
and U14277 (N_14277,N_13514,N_13575);
nor U14278 (N_14278,N_13028,N_13987);
or U14279 (N_14279,N_13639,N_13118);
xnor U14280 (N_14280,N_13307,N_13035);
nor U14281 (N_14281,N_13123,N_13760);
and U14282 (N_14282,N_13464,N_13029);
or U14283 (N_14283,N_13608,N_13379);
or U14284 (N_14284,N_13431,N_13046);
and U14285 (N_14285,N_13016,N_13159);
xor U14286 (N_14286,N_13942,N_13824);
or U14287 (N_14287,N_13251,N_13467);
xnor U14288 (N_14288,N_13752,N_13846);
and U14289 (N_14289,N_13532,N_13784);
nor U14290 (N_14290,N_13207,N_13327);
or U14291 (N_14291,N_13472,N_13047);
nor U14292 (N_14292,N_13078,N_13919);
or U14293 (N_14293,N_13781,N_13098);
xnor U14294 (N_14294,N_13764,N_13983);
nand U14295 (N_14295,N_13498,N_13124);
nand U14296 (N_14296,N_13298,N_13408);
or U14297 (N_14297,N_13900,N_13721);
nand U14298 (N_14298,N_13654,N_13200);
and U14299 (N_14299,N_13132,N_13302);
and U14300 (N_14300,N_13162,N_13648);
and U14301 (N_14301,N_13157,N_13820);
nor U14302 (N_14302,N_13736,N_13761);
and U14303 (N_14303,N_13868,N_13692);
nand U14304 (N_14304,N_13070,N_13239);
or U14305 (N_14305,N_13927,N_13358);
nor U14306 (N_14306,N_13260,N_13719);
nand U14307 (N_14307,N_13996,N_13337);
or U14308 (N_14308,N_13333,N_13776);
or U14309 (N_14309,N_13396,N_13319);
nor U14310 (N_14310,N_13246,N_13263);
or U14311 (N_14311,N_13196,N_13409);
xnor U14312 (N_14312,N_13563,N_13537);
nor U14313 (N_14313,N_13222,N_13803);
nor U14314 (N_14314,N_13519,N_13595);
xor U14315 (N_14315,N_13017,N_13808);
nor U14316 (N_14316,N_13805,N_13839);
nor U14317 (N_14317,N_13305,N_13376);
xor U14318 (N_14318,N_13739,N_13168);
xor U14319 (N_14319,N_13627,N_13790);
and U14320 (N_14320,N_13237,N_13847);
or U14321 (N_14321,N_13644,N_13951);
and U14322 (N_14322,N_13506,N_13623);
xnor U14323 (N_14323,N_13952,N_13449);
nand U14324 (N_14324,N_13637,N_13567);
xnor U14325 (N_14325,N_13390,N_13816);
or U14326 (N_14326,N_13655,N_13923);
and U14327 (N_14327,N_13768,N_13515);
xor U14328 (N_14328,N_13684,N_13810);
nor U14329 (N_14329,N_13187,N_13882);
or U14330 (N_14330,N_13978,N_13690);
nor U14331 (N_14331,N_13554,N_13336);
nand U14332 (N_14332,N_13361,N_13190);
and U14333 (N_14333,N_13822,N_13672);
nand U14334 (N_14334,N_13210,N_13056);
or U14335 (N_14335,N_13266,N_13282);
and U14336 (N_14336,N_13833,N_13076);
or U14337 (N_14337,N_13109,N_13934);
xor U14338 (N_14338,N_13718,N_13791);
nor U14339 (N_14339,N_13242,N_13634);
nor U14340 (N_14340,N_13252,N_13055);
xnor U14341 (N_14341,N_13281,N_13762);
and U14342 (N_14342,N_13722,N_13264);
xnor U14343 (N_14343,N_13699,N_13074);
and U14344 (N_14344,N_13254,N_13729);
nand U14345 (N_14345,N_13176,N_13174);
nand U14346 (N_14346,N_13211,N_13283);
nor U14347 (N_14347,N_13836,N_13322);
nand U14348 (N_14348,N_13879,N_13354);
nand U14349 (N_14349,N_13630,N_13542);
or U14350 (N_14350,N_13828,N_13618);
or U14351 (N_14351,N_13965,N_13117);
nand U14352 (N_14352,N_13688,N_13388);
nand U14353 (N_14353,N_13051,N_13391);
nand U14354 (N_14354,N_13511,N_13732);
nor U14355 (N_14355,N_13913,N_13404);
xor U14356 (N_14356,N_13665,N_13401);
nor U14357 (N_14357,N_13223,N_13485);
or U14358 (N_14358,N_13344,N_13817);
and U14359 (N_14359,N_13642,N_13569);
and U14360 (N_14360,N_13316,N_13290);
or U14361 (N_14361,N_13596,N_13513);
xor U14362 (N_14362,N_13693,N_13288);
xnor U14363 (N_14363,N_13789,N_13447);
xnor U14364 (N_14364,N_13771,N_13023);
xnor U14365 (N_14365,N_13717,N_13160);
nor U14366 (N_14366,N_13892,N_13534);
or U14367 (N_14367,N_13811,N_13364);
nor U14368 (N_14368,N_13607,N_13441);
xor U14369 (N_14369,N_13544,N_13743);
xnor U14370 (N_14370,N_13292,N_13328);
nand U14371 (N_14371,N_13848,N_13932);
xnor U14372 (N_14372,N_13433,N_13835);
or U14373 (N_14373,N_13887,N_13799);
nor U14374 (N_14374,N_13347,N_13087);
nand U14375 (N_14375,N_13084,N_13710);
nor U14376 (N_14376,N_13597,N_13744);
xor U14377 (N_14377,N_13203,N_13652);
xor U14378 (N_14378,N_13802,N_13170);
nand U14379 (N_14379,N_13130,N_13265);
nor U14380 (N_14380,N_13910,N_13308);
nand U14381 (N_14381,N_13730,N_13573);
xor U14382 (N_14382,N_13040,N_13420);
nand U14383 (N_14383,N_13551,N_13348);
or U14384 (N_14384,N_13890,N_13057);
or U14385 (N_14385,N_13085,N_13754);
nor U14386 (N_14386,N_13825,N_13463);
nor U14387 (N_14387,N_13632,N_13669);
xnor U14388 (N_14388,N_13980,N_13646);
or U14389 (N_14389,N_13073,N_13571);
and U14390 (N_14390,N_13019,N_13946);
nand U14391 (N_14391,N_13613,N_13930);
xnor U14392 (N_14392,N_13243,N_13619);
nand U14393 (N_14393,N_13813,N_13680);
or U14394 (N_14394,N_13701,N_13475);
xor U14395 (N_14395,N_13658,N_13043);
nand U14396 (N_14396,N_13393,N_13767);
nor U14397 (N_14397,N_13625,N_13229);
nor U14398 (N_14398,N_13091,N_13561);
xnor U14399 (N_14399,N_13937,N_13600);
nand U14400 (N_14400,N_13273,N_13164);
or U14401 (N_14401,N_13837,N_13136);
nand U14402 (N_14402,N_13793,N_13368);
and U14403 (N_14403,N_13002,N_13973);
and U14404 (N_14404,N_13048,N_13929);
nand U14405 (N_14405,N_13071,N_13661);
nor U14406 (N_14406,N_13891,N_13792);
nand U14407 (N_14407,N_13713,N_13775);
and U14408 (N_14408,N_13317,N_13295);
nand U14409 (N_14409,N_13041,N_13856);
nor U14410 (N_14410,N_13865,N_13881);
nor U14411 (N_14411,N_13579,N_13152);
and U14412 (N_14412,N_13859,N_13179);
xor U14413 (N_14413,N_13446,N_13851);
or U14414 (N_14414,N_13351,N_13114);
xor U14415 (N_14415,N_13105,N_13610);
nand U14416 (N_14416,N_13274,N_13525);
nand U14417 (N_14417,N_13716,N_13838);
nor U14418 (N_14418,N_13171,N_13938);
nand U14419 (N_14419,N_13435,N_13349);
xor U14420 (N_14420,N_13531,N_13293);
xor U14421 (N_14421,N_13224,N_13970);
xnor U14422 (N_14422,N_13888,N_13862);
and U14423 (N_14423,N_13863,N_13968);
nand U14424 (N_14424,N_13603,N_13666);
nand U14425 (N_14425,N_13438,N_13208);
nor U14426 (N_14426,N_13957,N_13917);
xor U14427 (N_14427,N_13497,N_13510);
nor U14428 (N_14428,N_13395,N_13352);
and U14429 (N_14429,N_13935,N_13602);
and U14430 (N_14430,N_13442,N_13969);
nand U14431 (N_14431,N_13491,N_13916);
nand U14432 (N_14432,N_13673,N_13785);
nand U14433 (N_14433,N_13410,N_13568);
or U14434 (N_14434,N_13939,N_13470);
and U14435 (N_14435,N_13481,N_13640);
nor U14436 (N_14436,N_13780,N_13156);
xnor U14437 (N_14437,N_13698,N_13172);
xnor U14438 (N_14438,N_13588,N_13440);
nand U14439 (N_14439,N_13173,N_13209);
or U14440 (N_14440,N_13527,N_13559);
nand U14441 (N_14441,N_13233,N_13741);
xor U14442 (N_14442,N_13127,N_13800);
and U14443 (N_14443,N_13522,N_13685);
xnor U14444 (N_14444,N_13679,N_13922);
nor U14445 (N_14445,N_13782,N_13914);
and U14446 (N_14446,N_13886,N_13303);
nor U14447 (N_14447,N_13682,N_13370);
or U14448 (N_14448,N_13921,N_13426);
or U14449 (N_14449,N_13734,N_13677);
and U14450 (N_14450,N_13423,N_13631);
nand U14451 (N_14451,N_13365,N_13026);
and U14452 (N_14452,N_13022,N_13155);
or U14453 (N_14453,N_13415,N_13678);
nand U14454 (N_14454,N_13723,N_13194);
nor U14455 (N_14455,N_13494,N_13064);
nand U14456 (N_14456,N_13183,N_13855);
nand U14457 (N_14457,N_13163,N_13903);
xnor U14458 (N_14458,N_13834,N_13708);
and U14459 (N_14459,N_13507,N_13647);
xnor U14460 (N_14460,N_13199,N_13653);
and U14461 (N_14461,N_13339,N_13367);
or U14462 (N_14462,N_13649,N_13015);
or U14463 (N_14463,N_13509,N_13735);
xnor U14464 (N_14464,N_13014,N_13466);
or U14465 (N_14465,N_13955,N_13869);
or U14466 (N_14466,N_13284,N_13533);
and U14467 (N_14467,N_13700,N_13668);
nor U14468 (N_14468,N_13099,N_13626);
and U14469 (N_14469,N_13378,N_13384);
and U14470 (N_14470,N_13006,N_13226);
nor U14471 (N_14471,N_13986,N_13555);
nor U14472 (N_14472,N_13217,N_13772);
nand U14473 (N_14473,N_13880,N_13249);
or U14474 (N_14474,N_13539,N_13748);
and U14475 (N_14475,N_13928,N_13110);
xnor U14476 (N_14476,N_13801,N_13030);
and U14477 (N_14477,N_13757,N_13469);
or U14478 (N_14478,N_13971,N_13111);
or U14479 (N_14479,N_13011,N_13062);
xnor U14480 (N_14480,N_13001,N_13069);
nor U14481 (N_14481,N_13998,N_13166);
xnor U14482 (N_14482,N_13425,N_13614);
nand U14483 (N_14483,N_13621,N_13508);
xor U14484 (N_14484,N_13125,N_13823);
and U14485 (N_14485,N_13392,N_13897);
and U14486 (N_14486,N_13278,N_13758);
nand U14487 (N_14487,N_13755,N_13334);
and U14488 (N_14488,N_13444,N_13526);
xor U14489 (N_14489,N_13094,N_13691);
nor U14490 (N_14490,N_13818,N_13382);
nor U14491 (N_14491,N_13853,N_13375);
nand U14492 (N_14492,N_13153,N_13889);
nand U14493 (N_14493,N_13884,N_13997);
nand U14494 (N_14494,N_13083,N_13635);
xor U14495 (N_14495,N_13256,N_13053);
and U14496 (N_14496,N_13228,N_13871);
and U14497 (N_14497,N_13330,N_13042);
and U14498 (N_14498,N_13366,N_13553);
xnor U14499 (N_14499,N_13609,N_13214);
or U14500 (N_14500,N_13194,N_13837);
or U14501 (N_14501,N_13028,N_13809);
nand U14502 (N_14502,N_13070,N_13367);
and U14503 (N_14503,N_13796,N_13543);
xor U14504 (N_14504,N_13184,N_13967);
and U14505 (N_14505,N_13299,N_13829);
and U14506 (N_14506,N_13311,N_13746);
nand U14507 (N_14507,N_13751,N_13516);
xnor U14508 (N_14508,N_13599,N_13783);
nor U14509 (N_14509,N_13491,N_13267);
nor U14510 (N_14510,N_13986,N_13266);
or U14511 (N_14511,N_13167,N_13896);
or U14512 (N_14512,N_13704,N_13793);
nand U14513 (N_14513,N_13550,N_13091);
and U14514 (N_14514,N_13405,N_13320);
nor U14515 (N_14515,N_13079,N_13642);
and U14516 (N_14516,N_13449,N_13767);
nand U14517 (N_14517,N_13607,N_13644);
or U14518 (N_14518,N_13019,N_13067);
or U14519 (N_14519,N_13685,N_13678);
xor U14520 (N_14520,N_13027,N_13232);
xor U14521 (N_14521,N_13425,N_13991);
xor U14522 (N_14522,N_13319,N_13913);
and U14523 (N_14523,N_13066,N_13934);
xor U14524 (N_14524,N_13784,N_13796);
xnor U14525 (N_14525,N_13777,N_13099);
xor U14526 (N_14526,N_13738,N_13480);
xor U14527 (N_14527,N_13882,N_13855);
nor U14528 (N_14528,N_13013,N_13114);
or U14529 (N_14529,N_13121,N_13306);
or U14530 (N_14530,N_13373,N_13620);
xor U14531 (N_14531,N_13075,N_13570);
nor U14532 (N_14532,N_13747,N_13223);
xnor U14533 (N_14533,N_13333,N_13672);
or U14534 (N_14534,N_13524,N_13588);
and U14535 (N_14535,N_13663,N_13073);
or U14536 (N_14536,N_13819,N_13353);
and U14537 (N_14537,N_13863,N_13966);
xnor U14538 (N_14538,N_13391,N_13628);
or U14539 (N_14539,N_13348,N_13858);
or U14540 (N_14540,N_13439,N_13569);
nand U14541 (N_14541,N_13868,N_13152);
or U14542 (N_14542,N_13269,N_13607);
xor U14543 (N_14543,N_13734,N_13090);
or U14544 (N_14544,N_13348,N_13005);
nand U14545 (N_14545,N_13747,N_13027);
xor U14546 (N_14546,N_13450,N_13457);
xor U14547 (N_14547,N_13722,N_13429);
and U14548 (N_14548,N_13231,N_13310);
nand U14549 (N_14549,N_13772,N_13024);
xnor U14550 (N_14550,N_13273,N_13027);
nand U14551 (N_14551,N_13543,N_13482);
nand U14552 (N_14552,N_13445,N_13591);
or U14553 (N_14553,N_13688,N_13340);
nand U14554 (N_14554,N_13057,N_13672);
or U14555 (N_14555,N_13062,N_13079);
nor U14556 (N_14556,N_13395,N_13472);
or U14557 (N_14557,N_13550,N_13033);
or U14558 (N_14558,N_13602,N_13416);
and U14559 (N_14559,N_13959,N_13783);
or U14560 (N_14560,N_13893,N_13721);
and U14561 (N_14561,N_13411,N_13790);
nand U14562 (N_14562,N_13002,N_13602);
or U14563 (N_14563,N_13704,N_13326);
and U14564 (N_14564,N_13751,N_13216);
xnor U14565 (N_14565,N_13146,N_13315);
xnor U14566 (N_14566,N_13008,N_13980);
nand U14567 (N_14567,N_13635,N_13993);
and U14568 (N_14568,N_13999,N_13343);
or U14569 (N_14569,N_13325,N_13200);
or U14570 (N_14570,N_13420,N_13508);
nand U14571 (N_14571,N_13094,N_13533);
nor U14572 (N_14572,N_13139,N_13724);
nor U14573 (N_14573,N_13851,N_13813);
and U14574 (N_14574,N_13220,N_13538);
and U14575 (N_14575,N_13876,N_13061);
and U14576 (N_14576,N_13958,N_13652);
xnor U14577 (N_14577,N_13882,N_13950);
nand U14578 (N_14578,N_13297,N_13023);
or U14579 (N_14579,N_13975,N_13460);
nor U14580 (N_14580,N_13327,N_13124);
nand U14581 (N_14581,N_13821,N_13181);
and U14582 (N_14582,N_13335,N_13600);
nand U14583 (N_14583,N_13536,N_13790);
or U14584 (N_14584,N_13877,N_13367);
and U14585 (N_14585,N_13497,N_13320);
and U14586 (N_14586,N_13903,N_13720);
or U14587 (N_14587,N_13695,N_13456);
nor U14588 (N_14588,N_13101,N_13731);
xor U14589 (N_14589,N_13699,N_13823);
or U14590 (N_14590,N_13076,N_13144);
or U14591 (N_14591,N_13146,N_13982);
or U14592 (N_14592,N_13009,N_13409);
nand U14593 (N_14593,N_13966,N_13615);
and U14594 (N_14594,N_13693,N_13598);
nand U14595 (N_14595,N_13749,N_13675);
xnor U14596 (N_14596,N_13621,N_13149);
nor U14597 (N_14597,N_13517,N_13668);
or U14598 (N_14598,N_13466,N_13927);
nand U14599 (N_14599,N_13829,N_13151);
nor U14600 (N_14600,N_13386,N_13803);
xor U14601 (N_14601,N_13345,N_13222);
or U14602 (N_14602,N_13425,N_13716);
nand U14603 (N_14603,N_13025,N_13174);
nand U14604 (N_14604,N_13768,N_13217);
and U14605 (N_14605,N_13452,N_13053);
and U14606 (N_14606,N_13641,N_13222);
nand U14607 (N_14607,N_13358,N_13880);
nand U14608 (N_14608,N_13495,N_13950);
nand U14609 (N_14609,N_13012,N_13154);
nor U14610 (N_14610,N_13616,N_13942);
nand U14611 (N_14611,N_13043,N_13702);
nor U14612 (N_14612,N_13627,N_13296);
nor U14613 (N_14613,N_13330,N_13752);
nor U14614 (N_14614,N_13432,N_13653);
xor U14615 (N_14615,N_13677,N_13560);
nor U14616 (N_14616,N_13586,N_13726);
and U14617 (N_14617,N_13807,N_13788);
or U14618 (N_14618,N_13028,N_13575);
or U14619 (N_14619,N_13868,N_13415);
and U14620 (N_14620,N_13375,N_13065);
and U14621 (N_14621,N_13996,N_13484);
nand U14622 (N_14622,N_13268,N_13839);
or U14623 (N_14623,N_13742,N_13520);
xor U14624 (N_14624,N_13423,N_13982);
xor U14625 (N_14625,N_13385,N_13737);
nor U14626 (N_14626,N_13025,N_13524);
nand U14627 (N_14627,N_13842,N_13759);
nor U14628 (N_14628,N_13864,N_13612);
nand U14629 (N_14629,N_13665,N_13843);
xnor U14630 (N_14630,N_13660,N_13924);
nor U14631 (N_14631,N_13113,N_13435);
xor U14632 (N_14632,N_13852,N_13150);
nand U14633 (N_14633,N_13602,N_13706);
xnor U14634 (N_14634,N_13887,N_13145);
xor U14635 (N_14635,N_13009,N_13165);
xnor U14636 (N_14636,N_13572,N_13045);
and U14637 (N_14637,N_13733,N_13412);
nor U14638 (N_14638,N_13596,N_13469);
xor U14639 (N_14639,N_13788,N_13457);
nor U14640 (N_14640,N_13812,N_13161);
and U14641 (N_14641,N_13444,N_13904);
or U14642 (N_14642,N_13516,N_13203);
nor U14643 (N_14643,N_13813,N_13876);
and U14644 (N_14644,N_13094,N_13476);
xor U14645 (N_14645,N_13374,N_13849);
and U14646 (N_14646,N_13073,N_13898);
or U14647 (N_14647,N_13986,N_13885);
xnor U14648 (N_14648,N_13166,N_13521);
nand U14649 (N_14649,N_13979,N_13151);
nand U14650 (N_14650,N_13271,N_13239);
or U14651 (N_14651,N_13608,N_13529);
nand U14652 (N_14652,N_13952,N_13319);
nand U14653 (N_14653,N_13147,N_13783);
or U14654 (N_14654,N_13988,N_13810);
nand U14655 (N_14655,N_13515,N_13686);
xnor U14656 (N_14656,N_13392,N_13148);
or U14657 (N_14657,N_13336,N_13592);
xor U14658 (N_14658,N_13854,N_13545);
nand U14659 (N_14659,N_13672,N_13558);
nand U14660 (N_14660,N_13594,N_13782);
and U14661 (N_14661,N_13053,N_13760);
xnor U14662 (N_14662,N_13939,N_13078);
and U14663 (N_14663,N_13091,N_13677);
or U14664 (N_14664,N_13641,N_13327);
and U14665 (N_14665,N_13580,N_13549);
nand U14666 (N_14666,N_13161,N_13732);
or U14667 (N_14667,N_13648,N_13869);
xnor U14668 (N_14668,N_13804,N_13838);
xnor U14669 (N_14669,N_13979,N_13717);
xnor U14670 (N_14670,N_13942,N_13101);
or U14671 (N_14671,N_13414,N_13624);
or U14672 (N_14672,N_13161,N_13528);
and U14673 (N_14673,N_13132,N_13627);
nand U14674 (N_14674,N_13552,N_13159);
and U14675 (N_14675,N_13158,N_13392);
or U14676 (N_14676,N_13022,N_13042);
and U14677 (N_14677,N_13732,N_13321);
xnor U14678 (N_14678,N_13097,N_13360);
nor U14679 (N_14679,N_13514,N_13048);
xnor U14680 (N_14680,N_13367,N_13577);
and U14681 (N_14681,N_13504,N_13966);
xnor U14682 (N_14682,N_13219,N_13105);
or U14683 (N_14683,N_13431,N_13784);
and U14684 (N_14684,N_13656,N_13705);
nand U14685 (N_14685,N_13203,N_13279);
xnor U14686 (N_14686,N_13076,N_13976);
or U14687 (N_14687,N_13310,N_13031);
and U14688 (N_14688,N_13161,N_13310);
xnor U14689 (N_14689,N_13766,N_13518);
and U14690 (N_14690,N_13636,N_13642);
nand U14691 (N_14691,N_13295,N_13618);
nor U14692 (N_14692,N_13964,N_13193);
nand U14693 (N_14693,N_13040,N_13784);
nand U14694 (N_14694,N_13438,N_13166);
and U14695 (N_14695,N_13455,N_13918);
nor U14696 (N_14696,N_13745,N_13508);
nor U14697 (N_14697,N_13559,N_13073);
nand U14698 (N_14698,N_13484,N_13863);
xnor U14699 (N_14699,N_13165,N_13126);
xor U14700 (N_14700,N_13871,N_13112);
nor U14701 (N_14701,N_13703,N_13691);
nor U14702 (N_14702,N_13679,N_13122);
xor U14703 (N_14703,N_13038,N_13246);
or U14704 (N_14704,N_13985,N_13442);
nor U14705 (N_14705,N_13471,N_13178);
xnor U14706 (N_14706,N_13625,N_13940);
nor U14707 (N_14707,N_13985,N_13967);
nor U14708 (N_14708,N_13816,N_13238);
nand U14709 (N_14709,N_13935,N_13841);
nand U14710 (N_14710,N_13216,N_13081);
nand U14711 (N_14711,N_13856,N_13490);
xor U14712 (N_14712,N_13094,N_13713);
nand U14713 (N_14713,N_13991,N_13060);
xnor U14714 (N_14714,N_13660,N_13808);
nand U14715 (N_14715,N_13146,N_13299);
xor U14716 (N_14716,N_13825,N_13344);
nor U14717 (N_14717,N_13792,N_13548);
nor U14718 (N_14718,N_13874,N_13126);
and U14719 (N_14719,N_13361,N_13297);
and U14720 (N_14720,N_13548,N_13570);
nor U14721 (N_14721,N_13750,N_13791);
nor U14722 (N_14722,N_13336,N_13201);
and U14723 (N_14723,N_13001,N_13547);
xnor U14724 (N_14724,N_13826,N_13161);
nand U14725 (N_14725,N_13985,N_13793);
and U14726 (N_14726,N_13301,N_13673);
nor U14727 (N_14727,N_13080,N_13751);
or U14728 (N_14728,N_13382,N_13150);
nand U14729 (N_14729,N_13211,N_13073);
or U14730 (N_14730,N_13026,N_13232);
nor U14731 (N_14731,N_13881,N_13252);
nor U14732 (N_14732,N_13640,N_13449);
and U14733 (N_14733,N_13496,N_13507);
or U14734 (N_14734,N_13525,N_13332);
or U14735 (N_14735,N_13772,N_13505);
nor U14736 (N_14736,N_13259,N_13127);
and U14737 (N_14737,N_13617,N_13247);
xor U14738 (N_14738,N_13723,N_13243);
nand U14739 (N_14739,N_13396,N_13843);
and U14740 (N_14740,N_13047,N_13748);
nand U14741 (N_14741,N_13184,N_13482);
nor U14742 (N_14742,N_13082,N_13532);
or U14743 (N_14743,N_13775,N_13492);
xnor U14744 (N_14744,N_13167,N_13158);
nand U14745 (N_14745,N_13522,N_13770);
xnor U14746 (N_14746,N_13776,N_13657);
or U14747 (N_14747,N_13442,N_13528);
and U14748 (N_14748,N_13721,N_13798);
xor U14749 (N_14749,N_13910,N_13860);
or U14750 (N_14750,N_13668,N_13166);
or U14751 (N_14751,N_13020,N_13711);
and U14752 (N_14752,N_13442,N_13375);
or U14753 (N_14753,N_13543,N_13630);
and U14754 (N_14754,N_13521,N_13860);
and U14755 (N_14755,N_13776,N_13980);
xnor U14756 (N_14756,N_13207,N_13960);
nand U14757 (N_14757,N_13159,N_13347);
xor U14758 (N_14758,N_13864,N_13133);
xor U14759 (N_14759,N_13719,N_13197);
nand U14760 (N_14760,N_13654,N_13101);
xor U14761 (N_14761,N_13321,N_13817);
or U14762 (N_14762,N_13578,N_13195);
and U14763 (N_14763,N_13809,N_13728);
or U14764 (N_14764,N_13849,N_13222);
nand U14765 (N_14765,N_13339,N_13629);
nand U14766 (N_14766,N_13416,N_13432);
and U14767 (N_14767,N_13229,N_13007);
or U14768 (N_14768,N_13455,N_13028);
and U14769 (N_14769,N_13645,N_13984);
xor U14770 (N_14770,N_13247,N_13694);
xnor U14771 (N_14771,N_13834,N_13135);
or U14772 (N_14772,N_13986,N_13676);
or U14773 (N_14773,N_13763,N_13147);
nand U14774 (N_14774,N_13584,N_13235);
nand U14775 (N_14775,N_13946,N_13113);
xor U14776 (N_14776,N_13854,N_13112);
or U14777 (N_14777,N_13312,N_13641);
or U14778 (N_14778,N_13978,N_13201);
and U14779 (N_14779,N_13364,N_13494);
xnor U14780 (N_14780,N_13808,N_13331);
xor U14781 (N_14781,N_13828,N_13100);
or U14782 (N_14782,N_13576,N_13314);
xnor U14783 (N_14783,N_13098,N_13016);
xnor U14784 (N_14784,N_13212,N_13510);
or U14785 (N_14785,N_13902,N_13422);
or U14786 (N_14786,N_13539,N_13469);
xor U14787 (N_14787,N_13210,N_13085);
xnor U14788 (N_14788,N_13713,N_13157);
nand U14789 (N_14789,N_13374,N_13878);
and U14790 (N_14790,N_13185,N_13716);
or U14791 (N_14791,N_13933,N_13533);
xnor U14792 (N_14792,N_13683,N_13208);
or U14793 (N_14793,N_13728,N_13649);
xor U14794 (N_14794,N_13328,N_13555);
nand U14795 (N_14795,N_13919,N_13685);
xor U14796 (N_14796,N_13654,N_13580);
and U14797 (N_14797,N_13478,N_13036);
and U14798 (N_14798,N_13407,N_13522);
and U14799 (N_14799,N_13719,N_13156);
xnor U14800 (N_14800,N_13275,N_13642);
xnor U14801 (N_14801,N_13319,N_13930);
nor U14802 (N_14802,N_13838,N_13855);
nand U14803 (N_14803,N_13893,N_13232);
nor U14804 (N_14804,N_13334,N_13385);
xnor U14805 (N_14805,N_13133,N_13292);
nand U14806 (N_14806,N_13884,N_13966);
and U14807 (N_14807,N_13787,N_13557);
and U14808 (N_14808,N_13411,N_13187);
nand U14809 (N_14809,N_13898,N_13466);
nor U14810 (N_14810,N_13123,N_13580);
nor U14811 (N_14811,N_13232,N_13461);
xnor U14812 (N_14812,N_13690,N_13151);
nor U14813 (N_14813,N_13443,N_13165);
xnor U14814 (N_14814,N_13834,N_13430);
and U14815 (N_14815,N_13602,N_13555);
and U14816 (N_14816,N_13190,N_13000);
nand U14817 (N_14817,N_13893,N_13854);
nor U14818 (N_14818,N_13493,N_13679);
xor U14819 (N_14819,N_13553,N_13452);
nor U14820 (N_14820,N_13997,N_13663);
or U14821 (N_14821,N_13122,N_13460);
or U14822 (N_14822,N_13004,N_13884);
and U14823 (N_14823,N_13662,N_13892);
nand U14824 (N_14824,N_13162,N_13157);
and U14825 (N_14825,N_13790,N_13626);
nor U14826 (N_14826,N_13607,N_13417);
or U14827 (N_14827,N_13147,N_13983);
xor U14828 (N_14828,N_13831,N_13307);
and U14829 (N_14829,N_13418,N_13993);
and U14830 (N_14830,N_13022,N_13229);
xnor U14831 (N_14831,N_13243,N_13687);
xor U14832 (N_14832,N_13226,N_13409);
xnor U14833 (N_14833,N_13768,N_13497);
or U14834 (N_14834,N_13421,N_13886);
and U14835 (N_14835,N_13892,N_13380);
nand U14836 (N_14836,N_13213,N_13100);
and U14837 (N_14837,N_13249,N_13796);
xor U14838 (N_14838,N_13662,N_13997);
and U14839 (N_14839,N_13270,N_13462);
xor U14840 (N_14840,N_13099,N_13666);
or U14841 (N_14841,N_13582,N_13488);
or U14842 (N_14842,N_13919,N_13851);
or U14843 (N_14843,N_13819,N_13649);
nand U14844 (N_14844,N_13222,N_13575);
nand U14845 (N_14845,N_13618,N_13744);
xnor U14846 (N_14846,N_13971,N_13473);
nand U14847 (N_14847,N_13495,N_13580);
or U14848 (N_14848,N_13949,N_13203);
or U14849 (N_14849,N_13016,N_13125);
nand U14850 (N_14850,N_13044,N_13626);
or U14851 (N_14851,N_13787,N_13928);
and U14852 (N_14852,N_13778,N_13764);
nor U14853 (N_14853,N_13290,N_13352);
nand U14854 (N_14854,N_13105,N_13205);
or U14855 (N_14855,N_13201,N_13521);
or U14856 (N_14856,N_13024,N_13284);
nor U14857 (N_14857,N_13345,N_13680);
and U14858 (N_14858,N_13647,N_13625);
or U14859 (N_14859,N_13824,N_13701);
or U14860 (N_14860,N_13032,N_13708);
or U14861 (N_14861,N_13504,N_13089);
or U14862 (N_14862,N_13907,N_13010);
and U14863 (N_14863,N_13283,N_13655);
nor U14864 (N_14864,N_13817,N_13592);
xnor U14865 (N_14865,N_13314,N_13791);
nand U14866 (N_14866,N_13392,N_13291);
nor U14867 (N_14867,N_13051,N_13268);
nor U14868 (N_14868,N_13564,N_13159);
nand U14869 (N_14869,N_13934,N_13337);
nor U14870 (N_14870,N_13105,N_13467);
or U14871 (N_14871,N_13426,N_13009);
nand U14872 (N_14872,N_13223,N_13074);
xnor U14873 (N_14873,N_13646,N_13056);
and U14874 (N_14874,N_13614,N_13436);
xnor U14875 (N_14875,N_13225,N_13082);
nand U14876 (N_14876,N_13127,N_13952);
nor U14877 (N_14877,N_13420,N_13780);
and U14878 (N_14878,N_13820,N_13210);
nand U14879 (N_14879,N_13035,N_13299);
nand U14880 (N_14880,N_13245,N_13798);
and U14881 (N_14881,N_13103,N_13004);
xnor U14882 (N_14882,N_13011,N_13020);
and U14883 (N_14883,N_13182,N_13291);
nor U14884 (N_14884,N_13248,N_13839);
and U14885 (N_14885,N_13530,N_13460);
nand U14886 (N_14886,N_13139,N_13184);
xor U14887 (N_14887,N_13967,N_13048);
or U14888 (N_14888,N_13503,N_13904);
nand U14889 (N_14889,N_13561,N_13355);
nand U14890 (N_14890,N_13737,N_13024);
xor U14891 (N_14891,N_13461,N_13680);
xor U14892 (N_14892,N_13633,N_13753);
or U14893 (N_14893,N_13391,N_13883);
and U14894 (N_14894,N_13272,N_13162);
or U14895 (N_14895,N_13057,N_13730);
nand U14896 (N_14896,N_13222,N_13755);
xnor U14897 (N_14897,N_13589,N_13679);
and U14898 (N_14898,N_13987,N_13381);
xor U14899 (N_14899,N_13530,N_13377);
and U14900 (N_14900,N_13499,N_13538);
and U14901 (N_14901,N_13229,N_13925);
xnor U14902 (N_14902,N_13814,N_13120);
and U14903 (N_14903,N_13279,N_13603);
or U14904 (N_14904,N_13297,N_13276);
nand U14905 (N_14905,N_13725,N_13258);
nor U14906 (N_14906,N_13598,N_13039);
xor U14907 (N_14907,N_13019,N_13384);
xor U14908 (N_14908,N_13445,N_13587);
nor U14909 (N_14909,N_13679,N_13543);
nor U14910 (N_14910,N_13996,N_13702);
nand U14911 (N_14911,N_13717,N_13172);
nand U14912 (N_14912,N_13585,N_13177);
nand U14913 (N_14913,N_13714,N_13789);
xnor U14914 (N_14914,N_13178,N_13971);
nor U14915 (N_14915,N_13905,N_13321);
and U14916 (N_14916,N_13483,N_13283);
nor U14917 (N_14917,N_13635,N_13852);
and U14918 (N_14918,N_13177,N_13608);
or U14919 (N_14919,N_13364,N_13025);
nand U14920 (N_14920,N_13384,N_13753);
or U14921 (N_14921,N_13871,N_13461);
xor U14922 (N_14922,N_13075,N_13948);
or U14923 (N_14923,N_13929,N_13513);
nand U14924 (N_14924,N_13815,N_13570);
or U14925 (N_14925,N_13298,N_13200);
nand U14926 (N_14926,N_13379,N_13745);
nand U14927 (N_14927,N_13854,N_13900);
and U14928 (N_14928,N_13595,N_13653);
nand U14929 (N_14929,N_13120,N_13332);
nor U14930 (N_14930,N_13570,N_13397);
and U14931 (N_14931,N_13313,N_13941);
and U14932 (N_14932,N_13564,N_13289);
nand U14933 (N_14933,N_13889,N_13651);
xnor U14934 (N_14934,N_13604,N_13018);
nand U14935 (N_14935,N_13079,N_13793);
or U14936 (N_14936,N_13617,N_13383);
nor U14937 (N_14937,N_13396,N_13229);
nor U14938 (N_14938,N_13437,N_13742);
or U14939 (N_14939,N_13885,N_13213);
nand U14940 (N_14940,N_13790,N_13373);
xor U14941 (N_14941,N_13316,N_13531);
or U14942 (N_14942,N_13282,N_13396);
and U14943 (N_14943,N_13582,N_13356);
and U14944 (N_14944,N_13832,N_13628);
and U14945 (N_14945,N_13111,N_13926);
or U14946 (N_14946,N_13757,N_13763);
xnor U14947 (N_14947,N_13524,N_13465);
and U14948 (N_14948,N_13241,N_13484);
nand U14949 (N_14949,N_13951,N_13928);
nand U14950 (N_14950,N_13944,N_13269);
nor U14951 (N_14951,N_13205,N_13054);
or U14952 (N_14952,N_13020,N_13051);
xnor U14953 (N_14953,N_13119,N_13307);
and U14954 (N_14954,N_13408,N_13135);
nor U14955 (N_14955,N_13175,N_13813);
or U14956 (N_14956,N_13598,N_13857);
or U14957 (N_14957,N_13871,N_13487);
nor U14958 (N_14958,N_13288,N_13376);
xor U14959 (N_14959,N_13756,N_13920);
nor U14960 (N_14960,N_13283,N_13543);
and U14961 (N_14961,N_13794,N_13272);
nand U14962 (N_14962,N_13971,N_13441);
and U14963 (N_14963,N_13805,N_13389);
xnor U14964 (N_14964,N_13914,N_13316);
or U14965 (N_14965,N_13514,N_13478);
and U14966 (N_14966,N_13876,N_13271);
nand U14967 (N_14967,N_13635,N_13131);
nand U14968 (N_14968,N_13781,N_13493);
or U14969 (N_14969,N_13292,N_13398);
nor U14970 (N_14970,N_13063,N_13581);
and U14971 (N_14971,N_13507,N_13206);
nor U14972 (N_14972,N_13800,N_13534);
nor U14973 (N_14973,N_13045,N_13779);
xnor U14974 (N_14974,N_13905,N_13347);
xnor U14975 (N_14975,N_13291,N_13831);
nand U14976 (N_14976,N_13481,N_13873);
nor U14977 (N_14977,N_13596,N_13166);
nand U14978 (N_14978,N_13826,N_13549);
nor U14979 (N_14979,N_13434,N_13724);
xor U14980 (N_14980,N_13954,N_13412);
and U14981 (N_14981,N_13435,N_13506);
nand U14982 (N_14982,N_13621,N_13589);
nand U14983 (N_14983,N_13732,N_13434);
or U14984 (N_14984,N_13162,N_13754);
and U14985 (N_14985,N_13030,N_13681);
and U14986 (N_14986,N_13826,N_13128);
or U14987 (N_14987,N_13653,N_13056);
and U14988 (N_14988,N_13177,N_13420);
nor U14989 (N_14989,N_13128,N_13717);
and U14990 (N_14990,N_13225,N_13927);
nor U14991 (N_14991,N_13344,N_13641);
and U14992 (N_14992,N_13583,N_13234);
xor U14993 (N_14993,N_13043,N_13295);
nand U14994 (N_14994,N_13131,N_13511);
or U14995 (N_14995,N_13983,N_13312);
xor U14996 (N_14996,N_13534,N_13922);
or U14997 (N_14997,N_13140,N_13242);
xnor U14998 (N_14998,N_13236,N_13825);
xnor U14999 (N_14999,N_13621,N_13339);
xor U15000 (N_15000,N_14724,N_14722);
nand U15001 (N_15001,N_14266,N_14534);
nor U15002 (N_15002,N_14682,N_14910);
xnor U15003 (N_15003,N_14054,N_14090);
nor U15004 (N_15004,N_14779,N_14951);
and U15005 (N_15005,N_14042,N_14457);
and U15006 (N_15006,N_14752,N_14880);
or U15007 (N_15007,N_14484,N_14077);
or U15008 (N_15008,N_14933,N_14628);
and U15009 (N_15009,N_14255,N_14479);
nand U15010 (N_15010,N_14009,N_14284);
and U15011 (N_15011,N_14186,N_14818);
xor U15012 (N_15012,N_14893,N_14150);
xor U15013 (N_15013,N_14873,N_14633);
or U15014 (N_15014,N_14603,N_14028);
nor U15015 (N_15015,N_14698,N_14810);
xnor U15016 (N_15016,N_14902,N_14218);
and U15017 (N_15017,N_14812,N_14262);
nor U15018 (N_15018,N_14969,N_14317);
nor U15019 (N_15019,N_14907,N_14640);
nand U15020 (N_15020,N_14393,N_14421);
or U15021 (N_15021,N_14420,N_14816);
nor U15022 (N_15022,N_14161,N_14290);
and U15023 (N_15023,N_14587,N_14851);
or U15024 (N_15024,N_14076,N_14331);
or U15025 (N_15025,N_14430,N_14684);
or U15026 (N_15026,N_14449,N_14757);
nand U15027 (N_15027,N_14874,N_14746);
or U15028 (N_15028,N_14822,N_14855);
or U15029 (N_15029,N_14518,N_14794);
or U15030 (N_15030,N_14037,N_14462);
nand U15031 (N_15031,N_14216,N_14679);
nor U15032 (N_15032,N_14930,N_14013);
nand U15033 (N_15033,N_14945,N_14313);
or U15034 (N_15034,N_14738,N_14989);
or U15035 (N_15035,N_14413,N_14113);
or U15036 (N_15036,N_14120,N_14397);
nand U15037 (N_15037,N_14439,N_14777);
or U15038 (N_15038,N_14315,N_14440);
or U15039 (N_15039,N_14069,N_14596);
xnor U15040 (N_15040,N_14594,N_14972);
xnor U15041 (N_15041,N_14458,N_14140);
xnor U15042 (N_15042,N_14175,N_14012);
nand U15043 (N_15043,N_14645,N_14565);
nor U15044 (N_15044,N_14642,N_14775);
nor U15045 (N_15045,N_14342,N_14911);
nand U15046 (N_15046,N_14678,N_14423);
and U15047 (N_15047,N_14776,N_14731);
or U15048 (N_15048,N_14044,N_14387);
and U15049 (N_15049,N_14103,N_14233);
or U15050 (N_15050,N_14715,N_14496);
and U15051 (N_15051,N_14549,N_14477);
xnor U15052 (N_15052,N_14613,N_14735);
or U15053 (N_15053,N_14039,N_14916);
and U15054 (N_15054,N_14732,N_14490);
or U15055 (N_15055,N_14374,N_14510);
and U15056 (N_15056,N_14909,N_14192);
or U15057 (N_15057,N_14522,N_14996);
nor U15058 (N_15058,N_14174,N_14153);
nand U15059 (N_15059,N_14610,N_14048);
or U15060 (N_15060,N_14034,N_14629);
and U15061 (N_15061,N_14127,N_14723);
nor U15062 (N_15062,N_14124,N_14097);
nor U15063 (N_15063,N_14271,N_14520);
nor U15064 (N_15064,N_14714,N_14145);
and U15065 (N_15065,N_14657,N_14737);
nand U15066 (N_15066,N_14692,N_14562);
nor U15067 (N_15067,N_14859,N_14636);
or U15068 (N_15068,N_14986,N_14895);
or U15069 (N_15069,N_14553,N_14744);
xnor U15070 (N_15070,N_14027,N_14363);
nand U15071 (N_15071,N_14503,N_14237);
nor U15072 (N_15072,N_14303,N_14461);
nor U15073 (N_15073,N_14424,N_14672);
xnor U15074 (N_15074,N_14003,N_14478);
nor U15075 (N_15075,N_14059,N_14375);
or U15076 (N_15076,N_14292,N_14550);
and U15077 (N_15077,N_14924,N_14004);
nand U15078 (N_15078,N_14883,N_14295);
or U15079 (N_15079,N_14222,N_14592);
nor U15080 (N_15080,N_14858,N_14215);
and U15081 (N_15081,N_14452,N_14019);
and U15082 (N_15082,N_14083,N_14760);
xor U15083 (N_15083,N_14799,N_14041);
nand U15084 (N_15084,N_14551,N_14495);
nor U15085 (N_15085,N_14758,N_14730);
nor U15086 (N_15086,N_14343,N_14954);
xor U15087 (N_15087,N_14666,N_14467);
nor U15088 (N_15088,N_14489,N_14105);
or U15089 (N_15089,N_14182,N_14071);
or U15090 (N_15090,N_14991,N_14143);
nor U15091 (N_15091,N_14709,N_14507);
or U15092 (N_15092,N_14448,N_14024);
nor U15093 (N_15093,N_14780,N_14109);
or U15094 (N_15094,N_14185,N_14021);
and U15095 (N_15095,N_14767,N_14425);
xor U15096 (N_15096,N_14159,N_14095);
or U15097 (N_15097,N_14786,N_14035);
nor U15098 (N_15098,N_14288,N_14843);
or U15099 (N_15099,N_14371,N_14525);
and U15100 (N_15100,N_14789,N_14863);
and U15101 (N_15101,N_14414,N_14281);
xor U15102 (N_15102,N_14839,N_14405);
xnor U15103 (N_15103,N_14211,N_14166);
nand U15104 (N_15104,N_14253,N_14205);
nor U15105 (N_15105,N_14728,N_14199);
nor U15106 (N_15106,N_14871,N_14084);
and U15107 (N_15107,N_14649,N_14508);
and U15108 (N_15108,N_14154,N_14500);
and U15109 (N_15109,N_14572,N_14096);
nand U15110 (N_15110,N_14547,N_14849);
or U15111 (N_15111,N_14305,N_14241);
nand U15112 (N_15112,N_14395,N_14232);
xnor U15113 (N_15113,N_14400,N_14968);
nand U15114 (N_15114,N_14167,N_14614);
nor U15115 (N_15115,N_14260,N_14705);
or U15116 (N_15116,N_14514,N_14231);
xnor U15117 (N_15117,N_14959,N_14202);
nand U15118 (N_15118,N_14505,N_14408);
and U15119 (N_15119,N_14178,N_14023);
nand U15120 (N_15120,N_14051,N_14929);
xor U15121 (N_15121,N_14831,N_14604);
or U15122 (N_15122,N_14319,N_14415);
nor U15123 (N_15123,N_14686,N_14125);
xnor U15124 (N_15124,N_14234,N_14667);
nand U15125 (N_15125,N_14527,N_14653);
nand U15126 (N_15126,N_14378,N_14861);
or U15127 (N_15127,N_14569,N_14574);
nor U15128 (N_15128,N_14985,N_14402);
or U15129 (N_15129,N_14294,N_14743);
nand U15130 (N_15130,N_14245,N_14264);
xor U15131 (N_15131,N_14053,N_14468);
xnor U15132 (N_15132,N_14014,N_14509);
and U15133 (N_15133,N_14471,N_14618);
xnor U15134 (N_15134,N_14131,N_14598);
and U15135 (N_15135,N_14225,N_14310);
nor U15136 (N_15136,N_14312,N_14575);
nand U15137 (N_15137,N_14566,N_14783);
xor U15138 (N_15138,N_14011,N_14586);
xor U15139 (N_15139,N_14546,N_14325);
or U15140 (N_15140,N_14061,N_14309);
nand U15141 (N_15141,N_14302,N_14370);
nor U15142 (N_15142,N_14322,N_14516);
or U15143 (N_15143,N_14681,N_14208);
and U15144 (N_15144,N_14912,N_14064);
xnor U15145 (N_15145,N_14261,N_14632);
and U15146 (N_15146,N_14832,N_14155);
nand U15147 (N_15147,N_14060,N_14212);
xnor U15148 (N_15148,N_14038,N_14318);
nand U15149 (N_15149,N_14941,N_14755);
xor U15150 (N_15150,N_14570,N_14625);
xnor U15151 (N_15151,N_14904,N_14914);
xor U15152 (N_15152,N_14138,N_14918);
nor U15153 (N_15153,N_14357,N_14778);
or U15154 (N_15154,N_14114,N_14854);
nor U15155 (N_15155,N_14062,N_14339);
nand U15156 (N_15156,N_14406,N_14931);
nor U15157 (N_15157,N_14391,N_14938);
nor U15158 (N_15158,N_14943,N_14669);
nor U15159 (N_15159,N_14892,N_14967);
and U15160 (N_15160,N_14811,N_14431);
xnor U15161 (N_15161,N_14676,N_14382);
xor U15162 (N_15162,N_14144,N_14589);
xnor U15163 (N_15163,N_14079,N_14040);
nor U15164 (N_15164,N_14602,N_14360);
and U15165 (N_15165,N_14162,N_14187);
nand U15166 (N_15166,N_14773,N_14373);
nand U15167 (N_15167,N_14052,N_14285);
or U15168 (N_15168,N_14639,N_14739);
xor U15169 (N_15169,N_14726,N_14107);
nor U15170 (N_15170,N_14050,N_14944);
or U15171 (N_15171,N_14949,N_14541);
xnor U15172 (N_15172,N_14611,N_14492);
nand U15173 (N_15173,N_14635,N_14544);
nand U15174 (N_15174,N_14242,N_14803);
and U15175 (N_15175,N_14821,N_14427);
and U15176 (N_15176,N_14766,N_14085);
xnor U15177 (N_15177,N_14984,N_14273);
and U15178 (N_15178,N_14765,N_14976);
or U15179 (N_15179,N_14258,N_14022);
nand U15180 (N_15180,N_14134,N_14605);
nor U15181 (N_15181,N_14655,N_14963);
or U15182 (N_15182,N_14795,N_14227);
or U15183 (N_15183,N_14081,N_14354);
nor U15184 (N_15184,N_14734,N_14235);
nand U15185 (N_15185,N_14833,N_14422);
nor U15186 (N_15186,N_14180,N_14946);
nor U15187 (N_15187,N_14287,N_14117);
nand U15188 (N_15188,N_14286,N_14057);
nor U15189 (N_15189,N_14151,N_14512);
nor U15190 (N_15190,N_14136,N_14445);
nor U15191 (N_15191,N_14966,N_14361);
and U15192 (N_15192,N_14531,N_14224);
and U15193 (N_15193,N_14753,N_14919);
or U15194 (N_15194,N_14341,N_14671);
xor U15195 (N_15195,N_14497,N_14141);
and U15196 (N_15196,N_14046,N_14068);
or U15197 (N_15197,N_14030,N_14588);
nor U15198 (N_15198,N_14889,N_14875);
xor U15199 (N_15199,N_14089,N_14214);
xnor U15200 (N_15200,N_14769,N_14326);
xor U15201 (N_15201,N_14121,N_14072);
nand U15202 (N_15202,N_14868,N_14937);
nand U15203 (N_15203,N_14920,N_14501);
or U15204 (N_15204,N_14158,N_14947);
nand U15205 (N_15205,N_14763,N_14729);
xnor U15206 (N_15206,N_14321,N_14545);
and U15207 (N_15207,N_14538,N_14418);
or U15208 (N_15208,N_14813,N_14466);
nor U15209 (N_15209,N_14366,N_14523);
nor U15210 (N_15210,N_14965,N_14992);
or U15211 (N_15211,N_14239,N_14619);
and U15212 (N_15212,N_14164,N_14785);
or U15213 (N_15213,N_14680,N_14612);
or U15214 (N_15214,N_14349,N_14844);
nand U15215 (N_15215,N_14648,N_14189);
xor U15216 (N_15216,N_14915,N_14088);
xnor U15217 (N_15217,N_14700,N_14793);
or U15218 (N_15218,N_14787,N_14282);
xor U15219 (N_15219,N_14289,N_14369);
nand U15220 (N_15220,N_14656,N_14845);
or U15221 (N_15221,N_14177,N_14256);
nand U15222 (N_15222,N_14200,N_14116);
nand U15223 (N_15223,N_14383,N_14593);
xor U15224 (N_15224,N_14554,N_14848);
and U15225 (N_15225,N_14257,N_14459);
xor U15226 (N_15226,N_14555,N_14917);
xnor U15227 (N_15227,N_14974,N_14206);
and U15228 (N_15228,N_14197,N_14494);
nand U15229 (N_15229,N_14950,N_14364);
nor U15230 (N_15230,N_14396,N_14311);
nor U15231 (N_15231,N_14561,N_14008);
and U15232 (N_15232,N_14796,N_14517);
nor U15233 (N_15233,N_14198,N_14841);
or U15234 (N_15234,N_14171,N_14804);
or U15235 (N_15235,N_14830,N_14870);
and U15236 (N_15236,N_14623,N_14073);
and U15237 (N_15237,N_14470,N_14246);
or U15238 (N_15238,N_14480,N_14784);
or U15239 (N_15239,N_14228,N_14699);
nor U15240 (N_15240,N_14169,N_14377);
xor U15241 (N_15241,N_14270,N_14638);
or U15242 (N_15242,N_14347,N_14454);
or U15243 (N_15243,N_14998,N_14519);
nor U15244 (N_15244,N_14958,N_14754);
xor U15245 (N_15245,N_14721,N_14469);
nor U15246 (N_15246,N_14601,N_14647);
xor U15247 (N_15247,N_14579,N_14890);
and U15248 (N_15248,N_14674,N_14130);
and U15249 (N_15249,N_14564,N_14543);
nand U15250 (N_15250,N_14379,N_14573);
or U15251 (N_15251,N_14817,N_14390);
or U15252 (N_15252,N_14450,N_14314);
nor U15253 (N_15253,N_14316,N_14894);
or U15254 (N_15254,N_14328,N_14913);
xor U15255 (N_15255,N_14971,N_14711);
xnor U15256 (N_15256,N_14280,N_14372);
and U15257 (N_15257,N_14537,N_14176);
and U15258 (N_15258,N_14925,N_14112);
or U15259 (N_15259,N_14988,N_14923);
nand U15260 (N_15260,N_14173,N_14668);
nor U15261 (N_15261,N_14032,N_14007);
nor U15262 (N_15262,N_14908,N_14864);
nor U15263 (N_15263,N_14170,N_14590);
nand U15264 (N_15264,N_14359,N_14304);
and U15265 (N_15265,N_14617,N_14188);
or U15266 (N_15266,N_14350,N_14622);
xnor U15267 (N_15267,N_14641,N_14438);
nand U15268 (N_15268,N_14386,N_14165);
and U15269 (N_15269,N_14585,N_14903);
xor U15270 (N_15270,N_14720,N_14226);
xnor U15271 (N_15271,N_14394,N_14100);
and U15272 (N_15272,N_14269,N_14696);
xnor U15273 (N_15273,N_14005,N_14591);
or U15274 (N_15274,N_14993,N_14838);
xor U15275 (N_15275,N_14001,N_14230);
and U15276 (N_15276,N_14432,N_14825);
nor U15277 (N_15277,N_14901,N_14194);
or U15278 (N_15278,N_14719,N_14249);
and U15279 (N_15279,N_14788,N_14982);
or U15280 (N_15280,N_14884,N_14099);
xnor U15281 (N_15281,N_14987,N_14133);
nand U15282 (N_15282,N_14663,N_14745);
and U15283 (N_15283,N_14080,N_14184);
nor U15284 (N_15284,N_14535,N_14247);
xnor U15285 (N_15285,N_14797,N_14948);
and U15286 (N_15286,N_14482,N_14869);
nor U15287 (N_15287,N_14552,N_14092);
or U15288 (N_15288,N_14244,N_14798);
nand U15289 (N_15289,N_14823,N_14118);
xnor U15290 (N_15290,N_14981,N_14352);
xnor U15291 (N_15291,N_14957,N_14762);
nand U15292 (N_15292,N_14878,N_14536);
or U15293 (N_15293,N_14842,N_14101);
and U15294 (N_15294,N_14563,N_14278);
nor U15295 (N_15295,N_14142,N_14691);
or U15296 (N_15296,N_14970,N_14772);
nor U15297 (N_15297,N_14560,N_14263);
xnor U15298 (N_15298,N_14451,N_14163);
nand U15299 (N_15299,N_14486,N_14990);
or U15300 (N_15300,N_14559,N_14031);
nand U15301 (N_15301,N_14504,N_14111);
and U15302 (N_15302,N_14624,N_14333);
nand U15303 (N_15303,N_14540,N_14000);
or U15304 (N_15304,N_14195,N_14433);
and U15305 (N_15305,N_14733,N_14447);
nand U15306 (N_15306,N_14411,N_14267);
nand U15307 (N_15307,N_14621,N_14358);
nand U15308 (N_15308,N_14654,N_14529);
nor U15309 (N_15309,N_14389,N_14217);
or U15310 (N_15310,N_14781,N_14058);
and U15311 (N_15311,N_14710,N_14708);
and U15312 (N_15312,N_14661,N_14074);
and U15313 (N_15313,N_14856,N_14251);
and U15314 (N_15314,N_14324,N_14712);
nor U15315 (N_15315,N_14181,N_14082);
or U15316 (N_15316,N_14677,N_14275);
xnor U15317 (N_15317,N_14017,N_14835);
or U15318 (N_15318,N_14942,N_14026);
or U15319 (N_15319,N_14345,N_14337);
nand U15320 (N_15320,N_14646,N_14857);
or U15321 (N_15321,N_14355,N_14277);
nand U15322 (N_15322,N_14716,N_14401);
or U15323 (N_15323,N_14087,N_14702);
and U15324 (N_15324,N_14132,N_14906);
nand U15325 (N_15325,N_14637,N_14043);
and U15326 (N_15326,N_14558,N_14306);
nor U15327 (N_15327,N_14236,N_14221);
nor U15328 (N_15328,N_14147,N_14717);
xor U15329 (N_15329,N_14515,N_14664);
nand U15330 (N_15330,N_14977,N_14521);
or U15331 (N_15331,N_14932,N_14066);
nand U15332 (N_15332,N_14660,N_14827);
xor U15333 (N_15333,N_14814,N_14403);
nor U15334 (N_15334,N_14761,N_14606);
or U15335 (N_15335,N_14852,N_14344);
nand U15336 (N_15336,N_14476,N_14029);
or U15337 (N_15337,N_14706,N_14240);
or U15338 (N_15338,N_14921,N_14532);
and U15339 (N_15339,N_14539,N_14353);
or U15340 (N_15340,N_14940,N_14568);
and U15341 (N_15341,N_14876,N_14094);
and U15342 (N_15342,N_14297,N_14464);
or U15343 (N_15343,N_14928,N_14453);
or U15344 (N_15344,N_14036,N_14759);
or U15345 (N_15345,N_14768,N_14481);
or U15346 (N_15346,N_14407,N_14697);
xnor U15347 (N_15347,N_14608,N_14300);
nor U15348 (N_15348,N_14307,N_14701);
and U15349 (N_15349,N_14748,N_14102);
or U15350 (N_15350,N_14557,N_14475);
nand U15351 (N_15351,N_14973,N_14524);
and U15352 (N_15352,N_14888,N_14179);
nand U15353 (N_15353,N_14047,N_14882);
nand U15354 (N_15354,N_14877,N_14806);
nor U15355 (N_15355,N_14196,N_14056);
and U15356 (N_15356,N_14223,N_14980);
nand U15357 (N_15357,N_14815,N_14820);
nor U15358 (N_15358,N_14126,N_14460);
nor U15359 (N_15359,N_14293,N_14578);
xnor U15360 (N_15360,N_14276,N_14006);
nand U15361 (N_15361,N_14010,N_14528);
nand U15362 (N_15362,N_14254,N_14771);
or U15363 (N_15363,N_14191,N_14687);
xnor U15364 (N_15364,N_14417,N_14485);
xor U15365 (N_15365,N_14997,N_14493);
xnor U15366 (N_15366,N_14428,N_14577);
and U15367 (N_15367,N_14351,N_14152);
nor U15368 (N_15368,N_14110,N_14160);
nand U15369 (N_15369,N_14203,N_14220);
or U15370 (N_15370,N_14862,N_14805);
and U15371 (N_15371,N_14866,N_14620);
xor U15372 (N_15372,N_14093,N_14879);
or U15373 (N_15373,N_14850,N_14782);
and U15374 (N_15374,N_14867,N_14597);
or U15375 (N_15375,N_14123,N_14384);
xor U15376 (N_15376,N_14802,N_14675);
or U15377 (N_15377,N_14463,N_14491);
or U15378 (N_15378,N_14695,N_14499);
xor U15379 (N_15379,N_14872,N_14104);
xor U15380 (N_15380,N_14488,N_14513);
nor U15381 (N_15381,N_14502,N_14652);
nor U15382 (N_15382,N_14193,N_14826);
and U15383 (N_15383,N_14346,N_14749);
xnor U15384 (N_15384,N_14498,N_14533);
or U15385 (N_15385,N_14659,N_14961);
or U15386 (N_15386,N_14388,N_14900);
or U15387 (N_15387,N_14434,N_14576);
or U15388 (N_15388,N_14800,N_14999);
and U15389 (N_15389,N_14740,N_14172);
and U15390 (N_15390,N_14670,N_14248);
xnor U15391 (N_15391,N_14122,N_14335);
xor U15392 (N_15392,N_14381,N_14694);
xor U15393 (N_15393,N_14157,N_14704);
nor U15394 (N_15394,N_14398,N_14885);
xor U15395 (N_15395,N_14207,N_14129);
nor U15396 (N_15396,N_14443,N_14229);
xor U15397 (N_15397,N_14853,N_14268);
nand U15398 (N_15398,N_14824,N_14905);
and U15399 (N_15399,N_14658,N_14365);
nand U15400 (N_15400,N_14409,N_14149);
and U15401 (N_15401,N_14265,N_14025);
nand U15402 (N_15402,N_14334,N_14616);
xnor U15403 (N_15403,N_14119,N_14718);
xnor U15404 (N_15404,N_14530,N_14108);
nand U15405 (N_15405,N_14571,N_14086);
or U15406 (N_15406,N_14320,N_14329);
and U15407 (N_15407,N_14819,N_14376);
and U15408 (N_15408,N_14790,N_14340);
and U15409 (N_15409,N_14774,N_14033);
xnor U15410 (N_15410,N_14016,N_14444);
nand U15411 (N_15411,N_14472,N_14070);
and U15412 (N_15412,N_14455,N_14887);
and U15413 (N_15413,N_14156,N_14442);
and U15414 (N_15414,N_14688,N_14308);
nand U15415 (N_15415,N_14404,N_14627);
nand U15416 (N_15416,N_14091,N_14922);
nor U15417 (N_15417,N_14327,N_14898);
and U15418 (N_15418,N_14219,N_14741);
and U15419 (N_15419,N_14865,N_14630);
or U15420 (N_15420,N_14807,N_14446);
and U15421 (N_15421,N_14581,N_14926);
and U15422 (N_15422,N_14049,N_14065);
xor U15423 (N_15423,N_14747,N_14018);
or U15424 (N_15424,N_14332,N_14296);
or U15425 (N_15425,N_14756,N_14330);
or U15426 (N_15426,N_14201,N_14983);
nor U15427 (N_15427,N_14298,N_14367);
nand U15428 (N_15428,N_14429,N_14846);
or U15429 (N_15429,N_14956,N_14437);
or U15430 (N_15430,N_14272,N_14939);
nand U15431 (N_15431,N_14673,N_14736);
and U15432 (N_15432,N_14441,N_14392);
nor U15433 (N_15433,N_14809,N_14356);
nor U15434 (N_15434,N_14742,N_14209);
or U15435 (N_15435,N_14662,N_14210);
nand U15436 (N_15436,N_14801,N_14435);
and U15437 (N_15437,N_14526,N_14665);
nand U15438 (N_15438,N_14055,N_14582);
and U15439 (N_15439,N_14643,N_14764);
and U15440 (N_15440,N_14994,N_14483);
nor U15441 (N_15441,N_14808,N_14964);
nor U15442 (N_15442,N_14323,N_14836);
nand U15443 (N_15443,N_14583,N_14506);
or U15444 (N_15444,N_14045,N_14934);
nor U15445 (N_15445,N_14098,N_14979);
and U15446 (N_15446,N_14474,N_14259);
and U15447 (N_15447,N_14683,N_14338);
and U15448 (N_15448,N_14703,N_14927);
and U15449 (N_15449,N_14891,N_14567);
xor U15450 (N_15450,N_14301,N_14693);
or U15451 (N_15451,N_14975,N_14380);
and U15452 (N_15452,N_14600,N_14727);
and U15453 (N_15453,N_14713,N_14487);
nand U15454 (N_15454,N_14137,N_14135);
and U15455 (N_15455,N_14829,N_14580);
xnor U15456 (N_15456,N_14078,N_14115);
or U15457 (N_15457,N_14283,N_14274);
xnor U15458 (N_15458,N_14348,N_14650);
or U15459 (N_15459,N_14252,N_14542);
and U15460 (N_15460,N_14139,N_14751);
and U15461 (N_15461,N_14607,N_14584);
or U15462 (N_15462,N_14238,N_14634);
or U15463 (N_15463,N_14644,N_14243);
and U15464 (N_15464,N_14168,N_14626);
nor U15465 (N_15465,N_14412,N_14609);
nand U15466 (N_15466,N_14190,N_14955);
nand U15467 (N_15467,N_14615,N_14465);
nor U15468 (N_15468,N_14279,N_14899);
or U15469 (N_15469,N_14960,N_14419);
nand U15470 (N_15470,N_14399,N_14128);
or U15471 (N_15471,N_14426,N_14897);
xnor U15472 (N_15472,N_14436,N_14410);
nand U15473 (N_15473,N_14953,N_14631);
and U15474 (N_15474,N_14291,N_14886);
nand U15475 (N_15475,N_14935,N_14791);
and U15476 (N_15476,N_14881,N_14978);
or U15477 (N_15477,N_14690,N_14368);
and U15478 (N_15478,N_14792,N_14847);
nor U15479 (N_15479,N_14952,N_14595);
xnor U15480 (N_15480,N_14651,N_14015);
nor U15481 (N_15481,N_14962,N_14860);
nor U15482 (N_15482,N_14385,N_14299);
and U15483 (N_15483,N_14213,N_14896);
nand U15484 (N_15484,N_14548,N_14183);
xnor U15485 (N_15485,N_14685,N_14416);
nor U15486 (N_15486,N_14770,N_14148);
nand U15487 (N_15487,N_14362,N_14995);
nand U15488 (N_15488,N_14002,N_14067);
nor U15489 (N_15489,N_14511,N_14828);
nor U15490 (N_15490,N_14689,N_14336);
and U15491 (N_15491,N_14075,N_14837);
nor U15492 (N_15492,N_14840,N_14725);
xnor U15493 (N_15493,N_14456,N_14106);
nor U15494 (N_15494,N_14204,N_14250);
nand U15495 (N_15495,N_14599,N_14020);
and U15496 (N_15496,N_14063,N_14473);
or U15497 (N_15497,N_14936,N_14146);
xnor U15498 (N_15498,N_14834,N_14750);
nor U15499 (N_15499,N_14556,N_14707);
or U15500 (N_15500,N_14857,N_14065);
xnor U15501 (N_15501,N_14144,N_14037);
nand U15502 (N_15502,N_14941,N_14731);
nand U15503 (N_15503,N_14668,N_14673);
and U15504 (N_15504,N_14159,N_14872);
nand U15505 (N_15505,N_14980,N_14347);
nor U15506 (N_15506,N_14925,N_14175);
nor U15507 (N_15507,N_14504,N_14985);
or U15508 (N_15508,N_14158,N_14754);
or U15509 (N_15509,N_14384,N_14233);
nor U15510 (N_15510,N_14182,N_14357);
and U15511 (N_15511,N_14314,N_14440);
and U15512 (N_15512,N_14735,N_14894);
nor U15513 (N_15513,N_14272,N_14307);
xor U15514 (N_15514,N_14505,N_14281);
and U15515 (N_15515,N_14399,N_14032);
nand U15516 (N_15516,N_14313,N_14554);
nor U15517 (N_15517,N_14284,N_14792);
and U15518 (N_15518,N_14908,N_14112);
nand U15519 (N_15519,N_14914,N_14109);
and U15520 (N_15520,N_14434,N_14231);
nor U15521 (N_15521,N_14104,N_14834);
xnor U15522 (N_15522,N_14670,N_14990);
nor U15523 (N_15523,N_14910,N_14855);
and U15524 (N_15524,N_14586,N_14258);
or U15525 (N_15525,N_14223,N_14860);
or U15526 (N_15526,N_14517,N_14659);
nor U15527 (N_15527,N_14525,N_14717);
or U15528 (N_15528,N_14927,N_14466);
or U15529 (N_15529,N_14281,N_14952);
nand U15530 (N_15530,N_14568,N_14591);
nor U15531 (N_15531,N_14047,N_14524);
nor U15532 (N_15532,N_14467,N_14790);
xor U15533 (N_15533,N_14580,N_14348);
xnor U15534 (N_15534,N_14648,N_14392);
or U15535 (N_15535,N_14873,N_14522);
or U15536 (N_15536,N_14916,N_14343);
nand U15537 (N_15537,N_14282,N_14243);
or U15538 (N_15538,N_14710,N_14054);
or U15539 (N_15539,N_14453,N_14289);
nand U15540 (N_15540,N_14752,N_14811);
nor U15541 (N_15541,N_14084,N_14594);
nor U15542 (N_15542,N_14987,N_14303);
nand U15543 (N_15543,N_14612,N_14186);
xnor U15544 (N_15544,N_14925,N_14578);
nand U15545 (N_15545,N_14464,N_14875);
nand U15546 (N_15546,N_14064,N_14012);
nand U15547 (N_15547,N_14533,N_14440);
nand U15548 (N_15548,N_14122,N_14524);
xor U15549 (N_15549,N_14520,N_14925);
nand U15550 (N_15550,N_14179,N_14118);
or U15551 (N_15551,N_14831,N_14063);
and U15552 (N_15552,N_14160,N_14621);
nor U15553 (N_15553,N_14986,N_14839);
nor U15554 (N_15554,N_14209,N_14579);
nand U15555 (N_15555,N_14923,N_14110);
or U15556 (N_15556,N_14506,N_14393);
and U15557 (N_15557,N_14718,N_14907);
xor U15558 (N_15558,N_14819,N_14031);
and U15559 (N_15559,N_14967,N_14342);
and U15560 (N_15560,N_14872,N_14736);
and U15561 (N_15561,N_14397,N_14467);
nor U15562 (N_15562,N_14390,N_14832);
or U15563 (N_15563,N_14915,N_14491);
nor U15564 (N_15564,N_14006,N_14250);
nand U15565 (N_15565,N_14898,N_14307);
nor U15566 (N_15566,N_14286,N_14633);
nor U15567 (N_15567,N_14344,N_14078);
and U15568 (N_15568,N_14878,N_14720);
nand U15569 (N_15569,N_14608,N_14727);
nor U15570 (N_15570,N_14454,N_14261);
xnor U15571 (N_15571,N_14652,N_14435);
xor U15572 (N_15572,N_14762,N_14410);
nand U15573 (N_15573,N_14189,N_14458);
nor U15574 (N_15574,N_14257,N_14470);
and U15575 (N_15575,N_14065,N_14333);
nor U15576 (N_15576,N_14423,N_14686);
nor U15577 (N_15577,N_14317,N_14378);
or U15578 (N_15578,N_14135,N_14644);
xnor U15579 (N_15579,N_14101,N_14492);
nand U15580 (N_15580,N_14581,N_14058);
nor U15581 (N_15581,N_14334,N_14844);
or U15582 (N_15582,N_14771,N_14670);
xnor U15583 (N_15583,N_14315,N_14832);
and U15584 (N_15584,N_14504,N_14293);
nand U15585 (N_15585,N_14504,N_14039);
and U15586 (N_15586,N_14711,N_14479);
nor U15587 (N_15587,N_14254,N_14429);
xnor U15588 (N_15588,N_14390,N_14530);
nand U15589 (N_15589,N_14423,N_14618);
xnor U15590 (N_15590,N_14187,N_14898);
or U15591 (N_15591,N_14362,N_14220);
or U15592 (N_15592,N_14051,N_14345);
nor U15593 (N_15593,N_14618,N_14414);
xor U15594 (N_15594,N_14472,N_14301);
nand U15595 (N_15595,N_14883,N_14083);
xnor U15596 (N_15596,N_14365,N_14912);
and U15597 (N_15597,N_14760,N_14618);
xor U15598 (N_15598,N_14712,N_14990);
nor U15599 (N_15599,N_14056,N_14993);
nand U15600 (N_15600,N_14085,N_14275);
nor U15601 (N_15601,N_14654,N_14485);
nand U15602 (N_15602,N_14376,N_14079);
nor U15603 (N_15603,N_14598,N_14014);
nor U15604 (N_15604,N_14344,N_14597);
and U15605 (N_15605,N_14063,N_14847);
and U15606 (N_15606,N_14585,N_14825);
or U15607 (N_15607,N_14339,N_14483);
xor U15608 (N_15608,N_14776,N_14513);
and U15609 (N_15609,N_14617,N_14609);
and U15610 (N_15610,N_14293,N_14508);
or U15611 (N_15611,N_14554,N_14139);
nand U15612 (N_15612,N_14405,N_14846);
and U15613 (N_15613,N_14705,N_14289);
nor U15614 (N_15614,N_14098,N_14392);
xnor U15615 (N_15615,N_14564,N_14974);
xnor U15616 (N_15616,N_14777,N_14295);
xor U15617 (N_15617,N_14658,N_14049);
or U15618 (N_15618,N_14134,N_14142);
xor U15619 (N_15619,N_14112,N_14721);
nor U15620 (N_15620,N_14562,N_14259);
and U15621 (N_15621,N_14696,N_14998);
or U15622 (N_15622,N_14299,N_14359);
or U15623 (N_15623,N_14340,N_14711);
and U15624 (N_15624,N_14373,N_14884);
or U15625 (N_15625,N_14094,N_14490);
xor U15626 (N_15626,N_14686,N_14953);
nor U15627 (N_15627,N_14408,N_14521);
xor U15628 (N_15628,N_14688,N_14672);
and U15629 (N_15629,N_14957,N_14310);
nand U15630 (N_15630,N_14180,N_14234);
xnor U15631 (N_15631,N_14591,N_14429);
nand U15632 (N_15632,N_14104,N_14647);
xnor U15633 (N_15633,N_14566,N_14521);
and U15634 (N_15634,N_14121,N_14069);
or U15635 (N_15635,N_14453,N_14672);
or U15636 (N_15636,N_14518,N_14284);
nand U15637 (N_15637,N_14270,N_14971);
nand U15638 (N_15638,N_14078,N_14357);
and U15639 (N_15639,N_14173,N_14764);
nor U15640 (N_15640,N_14765,N_14827);
or U15641 (N_15641,N_14313,N_14916);
nor U15642 (N_15642,N_14993,N_14088);
and U15643 (N_15643,N_14244,N_14958);
xnor U15644 (N_15644,N_14478,N_14699);
or U15645 (N_15645,N_14358,N_14475);
or U15646 (N_15646,N_14802,N_14125);
nor U15647 (N_15647,N_14891,N_14254);
and U15648 (N_15648,N_14007,N_14086);
nor U15649 (N_15649,N_14973,N_14561);
nor U15650 (N_15650,N_14625,N_14526);
and U15651 (N_15651,N_14733,N_14818);
xor U15652 (N_15652,N_14386,N_14077);
nor U15653 (N_15653,N_14910,N_14727);
nand U15654 (N_15654,N_14813,N_14826);
nor U15655 (N_15655,N_14285,N_14950);
xor U15656 (N_15656,N_14872,N_14943);
and U15657 (N_15657,N_14996,N_14021);
xnor U15658 (N_15658,N_14357,N_14845);
or U15659 (N_15659,N_14055,N_14586);
and U15660 (N_15660,N_14935,N_14108);
and U15661 (N_15661,N_14744,N_14342);
nor U15662 (N_15662,N_14268,N_14359);
and U15663 (N_15663,N_14557,N_14968);
nand U15664 (N_15664,N_14689,N_14721);
and U15665 (N_15665,N_14304,N_14349);
nand U15666 (N_15666,N_14589,N_14802);
or U15667 (N_15667,N_14750,N_14889);
nand U15668 (N_15668,N_14093,N_14478);
xor U15669 (N_15669,N_14791,N_14202);
and U15670 (N_15670,N_14926,N_14735);
nor U15671 (N_15671,N_14969,N_14817);
nor U15672 (N_15672,N_14769,N_14156);
xor U15673 (N_15673,N_14151,N_14620);
or U15674 (N_15674,N_14023,N_14123);
or U15675 (N_15675,N_14751,N_14618);
nor U15676 (N_15676,N_14940,N_14057);
xor U15677 (N_15677,N_14531,N_14925);
nand U15678 (N_15678,N_14393,N_14659);
or U15679 (N_15679,N_14703,N_14880);
and U15680 (N_15680,N_14998,N_14630);
nor U15681 (N_15681,N_14723,N_14565);
and U15682 (N_15682,N_14834,N_14396);
nor U15683 (N_15683,N_14305,N_14913);
and U15684 (N_15684,N_14682,N_14421);
nor U15685 (N_15685,N_14575,N_14206);
nor U15686 (N_15686,N_14561,N_14158);
or U15687 (N_15687,N_14000,N_14129);
nor U15688 (N_15688,N_14068,N_14344);
or U15689 (N_15689,N_14318,N_14926);
and U15690 (N_15690,N_14736,N_14847);
or U15691 (N_15691,N_14803,N_14539);
nor U15692 (N_15692,N_14418,N_14998);
or U15693 (N_15693,N_14155,N_14056);
xnor U15694 (N_15694,N_14879,N_14821);
xnor U15695 (N_15695,N_14798,N_14972);
nand U15696 (N_15696,N_14039,N_14654);
xor U15697 (N_15697,N_14354,N_14960);
and U15698 (N_15698,N_14677,N_14729);
or U15699 (N_15699,N_14915,N_14677);
xor U15700 (N_15700,N_14936,N_14558);
nand U15701 (N_15701,N_14305,N_14734);
nand U15702 (N_15702,N_14984,N_14282);
nand U15703 (N_15703,N_14496,N_14195);
nor U15704 (N_15704,N_14068,N_14132);
xnor U15705 (N_15705,N_14776,N_14518);
or U15706 (N_15706,N_14763,N_14801);
and U15707 (N_15707,N_14571,N_14968);
nand U15708 (N_15708,N_14987,N_14063);
and U15709 (N_15709,N_14141,N_14048);
nor U15710 (N_15710,N_14683,N_14407);
nor U15711 (N_15711,N_14673,N_14451);
nand U15712 (N_15712,N_14874,N_14284);
nor U15713 (N_15713,N_14169,N_14019);
nor U15714 (N_15714,N_14812,N_14676);
xnor U15715 (N_15715,N_14732,N_14515);
nor U15716 (N_15716,N_14061,N_14365);
nand U15717 (N_15717,N_14451,N_14715);
xnor U15718 (N_15718,N_14520,N_14102);
xnor U15719 (N_15719,N_14417,N_14716);
nand U15720 (N_15720,N_14584,N_14165);
nor U15721 (N_15721,N_14849,N_14786);
xor U15722 (N_15722,N_14133,N_14343);
xnor U15723 (N_15723,N_14444,N_14501);
or U15724 (N_15724,N_14977,N_14069);
nand U15725 (N_15725,N_14795,N_14150);
or U15726 (N_15726,N_14041,N_14101);
or U15727 (N_15727,N_14351,N_14965);
or U15728 (N_15728,N_14625,N_14814);
and U15729 (N_15729,N_14530,N_14666);
nand U15730 (N_15730,N_14196,N_14875);
xor U15731 (N_15731,N_14923,N_14557);
nand U15732 (N_15732,N_14266,N_14043);
and U15733 (N_15733,N_14125,N_14593);
nand U15734 (N_15734,N_14704,N_14200);
xnor U15735 (N_15735,N_14523,N_14738);
and U15736 (N_15736,N_14742,N_14891);
nor U15737 (N_15737,N_14755,N_14877);
xor U15738 (N_15738,N_14892,N_14814);
or U15739 (N_15739,N_14519,N_14666);
and U15740 (N_15740,N_14327,N_14745);
nand U15741 (N_15741,N_14902,N_14154);
or U15742 (N_15742,N_14735,N_14294);
nor U15743 (N_15743,N_14148,N_14835);
nor U15744 (N_15744,N_14486,N_14584);
nor U15745 (N_15745,N_14040,N_14134);
nor U15746 (N_15746,N_14681,N_14918);
xnor U15747 (N_15747,N_14038,N_14099);
nand U15748 (N_15748,N_14200,N_14676);
nand U15749 (N_15749,N_14248,N_14337);
nor U15750 (N_15750,N_14963,N_14972);
xnor U15751 (N_15751,N_14131,N_14639);
and U15752 (N_15752,N_14233,N_14651);
xor U15753 (N_15753,N_14082,N_14548);
xnor U15754 (N_15754,N_14556,N_14465);
and U15755 (N_15755,N_14673,N_14862);
xnor U15756 (N_15756,N_14420,N_14876);
and U15757 (N_15757,N_14231,N_14023);
and U15758 (N_15758,N_14369,N_14691);
nor U15759 (N_15759,N_14749,N_14038);
nor U15760 (N_15760,N_14090,N_14185);
or U15761 (N_15761,N_14006,N_14156);
and U15762 (N_15762,N_14145,N_14480);
xor U15763 (N_15763,N_14456,N_14657);
nand U15764 (N_15764,N_14829,N_14524);
xor U15765 (N_15765,N_14718,N_14016);
xnor U15766 (N_15766,N_14329,N_14512);
nor U15767 (N_15767,N_14995,N_14239);
and U15768 (N_15768,N_14073,N_14080);
nor U15769 (N_15769,N_14378,N_14617);
nor U15770 (N_15770,N_14775,N_14351);
or U15771 (N_15771,N_14690,N_14863);
and U15772 (N_15772,N_14340,N_14272);
nand U15773 (N_15773,N_14586,N_14784);
and U15774 (N_15774,N_14013,N_14582);
nor U15775 (N_15775,N_14808,N_14806);
or U15776 (N_15776,N_14164,N_14113);
xor U15777 (N_15777,N_14159,N_14162);
and U15778 (N_15778,N_14623,N_14386);
nand U15779 (N_15779,N_14427,N_14125);
nor U15780 (N_15780,N_14055,N_14783);
and U15781 (N_15781,N_14724,N_14664);
or U15782 (N_15782,N_14185,N_14313);
nor U15783 (N_15783,N_14383,N_14573);
nand U15784 (N_15784,N_14159,N_14561);
nor U15785 (N_15785,N_14947,N_14349);
xor U15786 (N_15786,N_14220,N_14012);
nand U15787 (N_15787,N_14070,N_14096);
nand U15788 (N_15788,N_14887,N_14242);
or U15789 (N_15789,N_14090,N_14083);
or U15790 (N_15790,N_14616,N_14990);
nand U15791 (N_15791,N_14474,N_14886);
nor U15792 (N_15792,N_14300,N_14947);
or U15793 (N_15793,N_14774,N_14130);
or U15794 (N_15794,N_14727,N_14271);
or U15795 (N_15795,N_14209,N_14009);
and U15796 (N_15796,N_14818,N_14511);
or U15797 (N_15797,N_14688,N_14231);
or U15798 (N_15798,N_14737,N_14574);
nand U15799 (N_15799,N_14195,N_14081);
or U15800 (N_15800,N_14439,N_14285);
or U15801 (N_15801,N_14136,N_14478);
nand U15802 (N_15802,N_14154,N_14290);
or U15803 (N_15803,N_14169,N_14185);
nand U15804 (N_15804,N_14990,N_14499);
xor U15805 (N_15805,N_14587,N_14862);
nand U15806 (N_15806,N_14284,N_14315);
nand U15807 (N_15807,N_14903,N_14444);
xor U15808 (N_15808,N_14200,N_14726);
or U15809 (N_15809,N_14640,N_14363);
and U15810 (N_15810,N_14506,N_14431);
xnor U15811 (N_15811,N_14603,N_14837);
nor U15812 (N_15812,N_14681,N_14895);
or U15813 (N_15813,N_14619,N_14852);
nand U15814 (N_15814,N_14168,N_14070);
and U15815 (N_15815,N_14935,N_14963);
nand U15816 (N_15816,N_14797,N_14238);
xor U15817 (N_15817,N_14633,N_14087);
and U15818 (N_15818,N_14540,N_14043);
nor U15819 (N_15819,N_14456,N_14231);
and U15820 (N_15820,N_14011,N_14394);
xor U15821 (N_15821,N_14632,N_14111);
xnor U15822 (N_15822,N_14130,N_14436);
or U15823 (N_15823,N_14973,N_14246);
and U15824 (N_15824,N_14777,N_14493);
nor U15825 (N_15825,N_14048,N_14993);
xor U15826 (N_15826,N_14942,N_14441);
or U15827 (N_15827,N_14955,N_14662);
or U15828 (N_15828,N_14348,N_14777);
and U15829 (N_15829,N_14814,N_14384);
nor U15830 (N_15830,N_14606,N_14605);
nand U15831 (N_15831,N_14225,N_14282);
and U15832 (N_15832,N_14628,N_14459);
nand U15833 (N_15833,N_14888,N_14283);
nand U15834 (N_15834,N_14126,N_14050);
xor U15835 (N_15835,N_14317,N_14938);
nand U15836 (N_15836,N_14018,N_14200);
nor U15837 (N_15837,N_14954,N_14093);
and U15838 (N_15838,N_14901,N_14706);
nand U15839 (N_15839,N_14757,N_14274);
xnor U15840 (N_15840,N_14812,N_14883);
or U15841 (N_15841,N_14833,N_14107);
xnor U15842 (N_15842,N_14883,N_14957);
nand U15843 (N_15843,N_14962,N_14043);
xor U15844 (N_15844,N_14381,N_14024);
xor U15845 (N_15845,N_14125,N_14108);
xor U15846 (N_15846,N_14571,N_14825);
and U15847 (N_15847,N_14137,N_14917);
and U15848 (N_15848,N_14608,N_14145);
xnor U15849 (N_15849,N_14061,N_14468);
or U15850 (N_15850,N_14597,N_14396);
nand U15851 (N_15851,N_14897,N_14987);
or U15852 (N_15852,N_14678,N_14133);
and U15853 (N_15853,N_14371,N_14011);
nor U15854 (N_15854,N_14357,N_14034);
nor U15855 (N_15855,N_14138,N_14614);
nor U15856 (N_15856,N_14504,N_14323);
nor U15857 (N_15857,N_14021,N_14850);
xnor U15858 (N_15858,N_14069,N_14101);
or U15859 (N_15859,N_14367,N_14493);
or U15860 (N_15860,N_14991,N_14720);
nand U15861 (N_15861,N_14175,N_14543);
and U15862 (N_15862,N_14801,N_14144);
and U15863 (N_15863,N_14168,N_14292);
xor U15864 (N_15864,N_14919,N_14414);
xnor U15865 (N_15865,N_14918,N_14860);
nor U15866 (N_15866,N_14888,N_14778);
or U15867 (N_15867,N_14189,N_14529);
nor U15868 (N_15868,N_14892,N_14111);
and U15869 (N_15869,N_14214,N_14946);
nor U15870 (N_15870,N_14335,N_14189);
and U15871 (N_15871,N_14985,N_14962);
xnor U15872 (N_15872,N_14613,N_14534);
and U15873 (N_15873,N_14716,N_14675);
nand U15874 (N_15874,N_14904,N_14090);
or U15875 (N_15875,N_14069,N_14103);
xnor U15876 (N_15876,N_14682,N_14055);
or U15877 (N_15877,N_14066,N_14926);
and U15878 (N_15878,N_14233,N_14330);
nor U15879 (N_15879,N_14359,N_14110);
xor U15880 (N_15880,N_14114,N_14082);
and U15881 (N_15881,N_14652,N_14968);
or U15882 (N_15882,N_14055,N_14544);
or U15883 (N_15883,N_14377,N_14916);
and U15884 (N_15884,N_14378,N_14133);
xnor U15885 (N_15885,N_14202,N_14012);
nor U15886 (N_15886,N_14729,N_14336);
xor U15887 (N_15887,N_14476,N_14464);
or U15888 (N_15888,N_14184,N_14295);
nor U15889 (N_15889,N_14046,N_14652);
or U15890 (N_15890,N_14691,N_14494);
nor U15891 (N_15891,N_14182,N_14151);
xor U15892 (N_15892,N_14954,N_14882);
nor U15893 (N_15893,N_14993,N_14816);
and U15894 (N_15894,N_14038,N_14900);
nor U15895 (N_15895,N_14560,N_14496);
xor U15896 (N_15896,N_14988,N_14956);
nand U15897 (N_15897,N_14928,N_14458);
nor U15898 (N_15898,N_14897,N_14265);
or U15899 (N_15899,N_14842,N_14516);
or U15900 (N_15900,N_14957,N_14202);
or U15901 (N_15901,N_14480,N_14964);
or U15902 (N_15902,N_14600,N_14668);
or U15903 (N_15903,N_14923,N_14143);
xor U15904 (N_15904,N_14870,N_14400);
and U15905 (N_15905,N_14444,N_14722);
or U15906 (N_15906,N_14273,N_14052);
and U15907 (N_15907,N_14368,N_14711);
nor U15908 (N_15908,N_14611,N_14710);
nand U15909 (N_15909,N_14407,N_14112);
xnor U15910 (N_15910,N_14697,N_14676);
nand U15911 (N_15911,N_14929,N_14966);
or U15912 (N_15912,N_14191,N_14254);
and U15913 (N_15913,N_14775,N_14992);
and U15914 (N_15914,N_14294,N_14865);
and U15915 (N_15915,N_14328,N_14937);
and U15916 (N_15916,N_14629,N_14033);
and U15917 (N_15917,N_14921,N_14204);
xor U15918 (N_15918,N_14669,N_14231);
nor U15919 (N_15919,N_14487,N_14084);
or U15920 (N_15920,N_14923,N_14762);
xor U15921 (N_15921,N_14195,N_14174);
nor U15922 (N_15922,N_14982,N_14482);
nand U15923 (N_15923,N_14271,N_14287);
nor U15924 (N_15924,N_14855,N_14920);
nand U15925 (N_15925,N_14963,N_14644);
nand U15926 (N_15926,N_14132,N_14765);
xnor U15927 (N_15927,N_14144,N_14626);
and U15928 (N_15928,N_14136,N_14878);
nand U15929 (N_15929,N_14717,N_14934);
xor U15930 (N_15930,N_14846,N_14509);
xnor U15931 (N_15931,N_14955,N_14303);
and U15932 (N_15932,N_14466,N_14955);
or U15933 (N_15933,N_14233,N_14365);
nor U15934 (N_15934,N_14318,N_14367);
xor U15935 (N_15935,N_14093,N_14646);
xor U15936 (N_15936,N_14324,N_14138);
xnor U15937 (N_15937,N_14793,N_14168);
xor U15938 (N_15938,N_14756,N_14733);
nor U15939 (N_15939,N_14996,N_14535);
and U15940 (N_15940,N_14397,N_14465);
or U15941 (N_15941,N_14923,N_14561);
xor U15942 (N_15942,N_14267,N_14106);
xor U15943 (N_15943,N_14910,N_14090);
nand U15944 (N_15944,N_14449,N_14923);
xnor U15945 (N_15945,N_14415,N_14426);
or U15946 (N_15946,N_14537,N_14021);
xnor U15947 (N_15947,N_14268,N_14492);
nand U15948 (N_15948,N_14144,N_14931);
nand U15949 (N_15949,N_14810,N_14656);
or U15950 (N_15950,N_14628,N_14981);
and U15951 (N_15951,N_14697,N_14329);
nand U15952 (N_15952,N_14444,N_14907);
nor U15953 (N_15953,N_14640,N_14827);
xnor U15954 (N_15954,N_14121,N_14647);
and U15955 (N_15955,N_14378,N_14595);
xnor U15956 (N_15956,N_14577,N_14790);
nand U15957 (N_15957,N_14891,N_14007);
and U15958 (N_15958,N_14441,N_14997);
or U15959 (N_15959,N_14563,N_14115);
nor U15960 (N_15960,N_14206,N_14034);
nand U15961 (N_15961,N_14840,N_14524);
nor U15962 (N_15962,N_14623,N_14831);
nand U15963 (N_15963,N_14480,N_14803);
or U15964 (N_15964,N_14086,N_14527);
xnor U15965 (N_15965,N_14262,N_14611);
nand U15966 (N_15966,N_14111,N_14761);
or U15967 (N_15967,N_14380,N_14010);
nand U15968 (N_15968,N_14200,N_14206);
and U15969 (N_15969,N_14778,N_14232);
xnor U15970 (N_15970,N_14566,N_14264);
nand U15971 (N_15971,N_14955,N_14029);
and U15972 (N_15972,N_14791,N_14037);
and U15973 (N_15973,N_14122,N_14430);
xnor U15974 (N_15974,N_14126,N_14958);
or U15975 (N_15975,N_14139,N_14359);
nand U15976 (N_15976,N_14482,N_14162);
nor U15977 (N_15977,N_14577,N_14898);
nand U15978 (N_15978,N_14688,N_14195);
and U15979 (N_15979,N_14733,N_14970);
and U15980 (N_15980,N_14972,N_14878);
xnor U15981 (N_15981,N_14730,N_14711);
nand U15982 (N_15982,N_14337,N_14456);
or U15983 (N_15983,N_14933,N_14122);
and U15984 (N_15984,N_14497,N_14596);
and U15985 (N_15985,N_14159,N_14179);
nand U15986 (N_15986,N_14772,N_14085);
xor U15987 (N_15987,N_14160,N_14699);
nand U15988 (N_15988,N_14316,N_14803);
xnor U15989 (N_15989,N_14906,N_14648);
xor U15990 (N_15990,N_14256,N_14226);
or U15991 (N_15991,N_14271,N_14543);
nor U15992 (N_15992,N_14457,N_14336);
nand U15993 (N_15993,N_14422,N_14608);
xor U15994 (N_15994,N_14731,N_14501);
and U15995 (N_15995,N_14649,N_14255);
or U15996 (N_15996,N_14486,N_14660);
xnor U15997 (N_15997,N_14419,N_14013);
xnor U15998 (N_15998,N_14406,N_14507);
or U15999 (N_15999,N_14284,N_14095);
nor U16000 (N_16000,N_15538,N_15613);
nor U16001 (N_16001,N_15649,N_15922);
and U16002 (N_16002,N_15435,N_15745);
nor U16003 (N_16003,N_15446,N_15384);
xor U16004 (N_16004,N_15291,N_15262);
or U16005 (N_16005,N_15149,N_15899);
and U16006 (N_16006,N_15413,N_15898);
or U16007 (N_16007,N_15912,N_15390);
xnor U16008 (N_16008,N_15981,N_15924);
or U16009 (N_16009,N_15307,N_15071);
and U16010 (N_16010,N_15428,N_15814);
and U16011 (N_16011,N_15510,N_15812);
and U16012 (N_16012,N_15531,N_15969);
xnor U16013 (N_16013,N_15701,N_15058);
xor U16014 (N_16014,N_15250,N_15742);
xor U16015 (N_16015,N_15603,N_15209);
or U16016 (N_16016,N_15457,N_15949);
and U16017 (N_16017,N_15754,N_15865);
nand U16018 (N_16018,N_15686,N_15641);
and U16019 (N_16019,N_15550,N_15677);
xor U16020 (N_16020,N_15025,N_15840);
and U16021 (N_16021,N_15525,N_15959);
xor U16022 (N_16022,N_15393,N_15786);
and U16023 (N_16023,N_15204,N_15893);
nor U16024 (N_16024,N_15206,N_15312);
nor U16025 (N_16025,N_15859,N_15911);
xor U16026 (N_16026,N_15935,N_15261);
or U16027 (N_16027,N_15489,N_15228);
nand U16028 (N_16028,N_15001,N_15777);
and U16029 (N_16029,N_15746,N_15704);
nor U16030 (N_16030,N_15583,N_15294);
nand U16031 (N_16031,N_15028,N_15430);
nand U16032 (N_16032,N_15309,N_15243);
nor U16033 (N_16033,N_15275,N_15903);
and U16034 (N_16034,N_15093,N_15726);
or U16035 (N_16035,N_15144,N_15685);
nand U16036 (N_16036,N_15875,N_15886);
nor U16037 (N_16037,N_15425,N_15776);
nand U16038 (N_16038,N_15481,N_15241);
nor U16039 (N_16039,N_15353,N_15156);
nor U16040 (N_16040,N_15983,N_15456);
nor U16041 (N_16041,N_15574,N_15497);
xnor U16042 (N_16042,N_15637,N_15599);
nor U16043 (N_16043,N_15401,N_15696);
nor U16044 (N_16044,N_15295,N_15699);
xnor U16045 (N_16045,N_15468,N_15168);
or U16046 (N_16046,N_15545,N_15988);
xor U16047 (N_16047,N_15549,N_15589);
or U16048 (N_16048,N_15517,N_15439);
nand U16049 (N_16049,N_15064,N_15091);
or U16050 (N_16050,N_15923,N_15361);
xnor U16051 (N_16051,N_15824,N_15711);
or U16052 (N_16052,N_15744,N_15427);
and U16053 (N_16053,N_15639,N_15579);
xnor U16054 (N_16054,N_15593,N_15221);
xnor U16055 (N_16055,N_15046,N_15667);
and U16056 (N_16056,N_15993,N_15421);
nor U16057 (N_16057,N_15249,N_15519);
nor U16058 (N_16058,N_15129,N_15717);
or U16059 (N_16059,N_15815,N_15853);
and U16060 (N_16060,N_15304,N_15825);
nand U16061 (N_16061,N_15738,N_15161);
and U16062 (N_16062,N_15944,N_15917);
nor U16063 (N_16063,N_15326,N_15688);
nand U16064 (N_16064,N_15347,N_15966);
xnor U16065 (N_16065,N_15942,N_15775);
xor U16066 (N_16066,N_15086,N_15397);
and U16067 (N_16067,N_15410,N_15448);
or U16068 (N_16068,N_15089,N_15655);
nand U16069 (N_16069,N_15300,N_15470);
nand U16070 (N_16070,N_15120,N_15343);
or U16071 (N_16071,N_15873,N_15980);
nor U16072 (N_16072,N_15540,N_15765);
and U16073 (N_16073,N_15037,N_15488);
nor U16074 (N_16074,N_15956,N_15773);
xor U16075 (N_16075,N_15341,N_15547);
xor U16076 (N_16076,N_15163,N_15567);
xor U16077 (N_16077,N_15848,N_15118);
nand U16078 (N_16078,N_15672,N_15442);
xor U16079 (N_16079,N_15443,N_15679);
and U16080 (N_16080,N_15336,N_15978);
and U16081 (N_16081,N_15359,N_15648);
nand U16082 (N_16082,N_15965,N_15791);
nand U16083 (N_16083,N_15002,N_15143);
nor U16084 (N_16084,N_15405,N_15653);
nand U16085 (N_16085,N_15226,N_15654);
or U16086 (N_16086,N_15707,N_15344);
nor U16087 (N_16087,N_15061,N_15684);
xor U16088 (N_16088,N_15676,N_15330);
xor U16089 (N_16089,N_15996,N_15438);
xnor U16090 (N_16090,N_15392,N_15229);
xnor U16091 (N_16091,N_15609,N_15868);
xor U16092 (N_16092,N_15709,N_15458);
and U16093 (N_16093,N_15018,N_15887);
or U16094 (N_16094,N_15884,N_15635);
xor U16095 (N_16095,N_15819,N_15278);
xor U16096 (N_16096,N_15244,N_15755);
and U16097 (N_16097,N_15647,N_15069);
and U16098 (N_16098,N_15498,N_15533);
or U16099 (N_16099,N_15238,N_15260);
and U16100 (N_16100,N_15927,N_15124);
xnor U16101 (N_16101,N_15003,N_15495);
nand U16102 (N_16102,N_15175,N_15535);
xnor U16103 (N_16103,N_15346,N_15387);
nand U16104 (N_16104,N_15436,N_15863);
nor U16105 (N_16105,N_15584,N_15743);
xor U16106 (N_16106,N_15440,N_15400);
nand U16107 (N_16107,N_15728,N_15925);
nor U16108 (N_16108,N_15716,N_15408);
and U16109 (N_16109,N_15108,N_15740);
nand U16110 (N_16110,N_15720,N_15159);
nand U16111 (N_16111,N_15329,N_15461);
and U16112 (N_16112,N_15612,N_15009);
nand U16113 (N_16113,N_15422,N_15424);
or U16114 (N_16114,N_15659,N_15573);
xnor U16115 (N_16115,N_15693,N_15670);
xor U16116 (N_16116,N_15463,N_15013);
and U16117 (N_16117,N_15121,N_15842);
or U16118 (N_16118,N_15431,N_15571);
nor U16119 (N_16119,N_15551,N_15714);
and U16120 (N_16120,N_15809,N_15952);
or U16121 (N_16121,N_15102,N_15725);
and U16122 (N_16122,N_15587,N_15869);
nor U16123 (N_16123,N_15940,N_15317);
or U16124 (N_16124,N_15943,N_15795);
xnor U16125 (N_16125,N_15119,N_15065);
nor U16126 (N_16126,N_15762,N_15111);
or U16127 (N_16127,N_15059,N_15844);
nand U16128 (N_16128,N_15876,N_15181);
and U16129 (N_16129,N_15818,N_15817);
xor U16130 (N_16130,N_15565,N_15788);
nor U16131 (N_16131,N_15682,N_15896);
or U16132 (N_16132,N_15207,N_15205);
or U16133 (N_16133,N_15423,N_15713);
nor U16134 (N_16134,N_15114,N_15402);
nor U16135 (N_16135,N_15836,N_15130);
nor U16136 (N_16136,N_15789,N_15586);
xor U16137 (N_16137,N_15890,N_15476);
nand U16138 (N_16138,N_15872,N_15808);
and U16139 (N_16139,N_15039,N_15044);
nor U16140 (N_16140,N_15629,N_15147);
xnor U16141 (N_16141,N_15564,N_15308);
xor U16142 (N_16142,N_15076,N_15338);
and U16143 (N_16143,N_15792,N_15546);
and U16144 (N_16144,N_15878,N_15251);
xnor U16145 (N_16145,N_15697,N_15656);
xnor U16146 (N_16146,N_15332,N_15381);
and U16147 (N_16147,N_15866,N_15377);
or U16148 (N_16148,N_15841,N_15215);
xnor U16149 (N_16149,N_15881,N_15999);
or U16150 (N_16150,N_15813,N_15617);
and U16151 (N_16151,N_15211,N_15504);
nor U16152 (N_16152,N_15706,N_15727);
or U16153 (N_16153,N_15953,N_15802);
xor U16154 (N_16154,N_15874,N_15214);
nor U16155 (N_16155,N_15561,N_15210);
or U16156 (N_16156,N_15657,N_15715);
and U16157 (N_16157,N_15945,N_15350);
and U16158 (N_16158,N_15099,N_15608);
or U16159 (N_16159,N_15318,N_15462);
xor U16160 (N_16160,N_15766,N_15015);
nand U16161 (N_16161,N_15459,N_15254);
xnor U16162 (N_16162,N_15266,N_15169);
or U16163 (N_16163,N_15370,N_15152);
and U16164 (N_16164,N_15736,N_15882);
or U16165 (N_16165,N_15581,N_15253);
or U16166 (N_16166,N_15471,N_15918);
nor U16167 (N_16167,N_15734,N_15995);
xnor U16168 (N_16168,N_15477,N_15908);
nor U16169 (N_16169,N_15880,N_15939);
or U16170 (N_16170,N_15501,N_15673);
or U16171 (N_16171,N_15406,N_15588);
or U16172 (N_16172,N_15005,N_15831);
xor U16173 (N_16173,N_15178,N_15311);
nand U16174 (N_16174,N_15395,N_15897);
or U16175 (N_16175,N_15257,N_15165);
xor U16176 (N_16176,N_15113,N_15179);
nand U16177 (N_16177,N_15137,N_15625);
xnor U16178 (N_16178,N_15074,N_15732);
nand U16179 (N_16179,N_15695,N_15947);
xnor U16180 (N_16180,N_15004,N_15164);
and U16181 (N_16181,N_15258,N_15731);
and U16182 (N_16182,N_15748,N_15472);
nand U16183 (N_16183,N_15404,N_15323);
nand U16184 (N_16184,N_15123,N_15473);
xnor U16185 (N_16185,N_15515,N_15548);
xor U16186 (N_16186,N_15757,N_15378);
xor U16187 (N_16187,N_15449,N_15465);
xor U16188 (N_16188,N_15466,N_15364);
nor U16189 (N_16189,N_15062,N_15277);
and U16190 (N_16190,N_15373,N_15138);
nor U16191 (N_16191,N_15200,N_15045);
nor U16192 (N_16192,N_15246,N_15722);
xnor U16193 (N_16193,N_15984,N_15033);
nand U16194 (N_16194,N_15595,N_15371);
and U16195 (N_16195,N_15883,N_15630);
or U16196 (N_16196,N_15919,N_15753);
and U16197 (N_16197,N_15823,N_15528);
nand U16198 (N_16198,N_15365,N_15409);
nor U16199 (N_16199,N_15621,N_15623);
nand U16200 (N_16200,N_15516,N_15894);
nand U16201 (N_16201,N_15860,N_15877);
xnor U16202 (N_16202,N_15139,N_15990);
nor U16203 (N_16203,N_15160,N_15521);
or U16204 (N_16204,N_15098,N_15441);
xnor U16205 (N_16205,N_15694,N_15447);
xnor U16206 (N_16206,N_15145,N_15958);
and U16207 (N_16207,N_15954,N_15718);
or U16208 (N_16208,N_15543,N_15097);
xor U16209 (N_16209,N_15047,N_15281);
xnor U16210 (N_16210,N_15867,N_15627);
and U16211 (N_16211,N_15104,N_15691);
xnor U16212 (N_16212,N_15038,N_15712);
or U16213 (N_16213,N_15216,N_15314);
and U16214 (N_16214,N_15513,N_15232);
xor U16215 (N_16215,N_15772,N_15591);
nand U16216 (N_16216,N_15974,N_15920);
and U16217 (N_16217,N_15474,N_15166);
nand U16218 (N_16218,N_15665,N_15987);
and U16219 (N_16219,N_15851,N_15030);
nor U16220 (N_16220,N_15803,N_15492);
xnor U16221 (N_16221,N_15095,N_15217);
and U16222 (N_16222,N_15761,N_15298);
nor U16223 (N_16223,N_15509,N_15590);
xor U16224 (N_16224,N_15950,N_15019);
or U16225 (N_16225,N_15453,N_15043);
or U16226 (N_16226,N_15563,N_15434);
or U16227 (N_16227,N_15126,N_15146);
or U16228 (N_16228,N_15522,N_15601);
xor U16229 (N_16229,N_15508,N_15027);
and U16230 (N_16230,N_15871,N_15000);
or U16231 (N_16231,N_15154,N_15642);
or U16232 (N_16232,N_15026,N_15451);
and U16233 (N_16233,N_15455,N_15683);
nand U16234 (N_16234,N_15255,N_15827);
or U16235 (N_16235,N_15839,N_15680);
or U16236 (N_16236,N_15354,N_15930);
nand U16237 (N_16237,N_15968,N_15049);
and U16238 (N_16238,N_15085,N_15188);
xor U16239 (N_16239,N_15426,N_15838);
and U16240 (N_16240,N_15997,N_15926);
xnor U16241 (N_16241,N_15356,N_15646);
nand U16242 (N_16242,N_15087,N_15220);
or U16243 (N_16243,N_15783,N_15989);
xnor U16244 (N_16244,N_15756,N_15372);
and U16245 (N_16245,N_15668,N_15398);
nor U16246 (N_16246,N_15475,N_15932);
and U16247 (N_16247,N_15190,N_15223);
or U16248 (N_16248,N_15035,N_15285);
nand U16249 (N_16249,N_15901,N_15558);
or U16250 (N_16250,N_15060,N_15857);
nor U16251 (N_16251,N_15763,N_15011);
and U16252 (N_16252,N_15846,N_15107);
and U16253 (N_16253,N_15572,N_15342);
or U16254 (N_16254,N_15382,N_15057);
nor U16255 (N_16255,N_15063,N_15328);
nor U16256 (N_16256,N_15575,N_15798);
xor U16257 (N_16257,N_15915,N_15394);
and U16258 (N_16258,N_15847,N_15263);
xor U16259 (N_16259,N_15267,N_15801);
and U16260 (N_16260,N_15610,N_15921);
and U16261 (N_16261,N_15596,N_15358);
nor U16262 (N_16262,N_15532,N_15403);
xnor U16263 (N_16263,N_15799,N_15080);
nand U16264 (N_16264,N_15991,N_15067);
or U16265 (N_16265,N_15539,N_15585);
and U16266 (N_16266,N_15389,N_15702);
and U16267 (N_16267,N_15512,N_15692);
nand U16268 (N_16268,N_15034,N_15418);
and U16269 (N_16269,N_15661,N_15502);
nor U16270 (N_16270,N_15022,N_15088);
nor U16271 (N_16271,N_15643,N_15979);
and U16272 (N_16272,N_15345,N_15416);
or U16273 (N_16273,N_15905,N_15396);
or U16274 (N_16274,N_15781,N_15117);
and U16275 (N_16275,N_15376,N_15202);
and U16276 (N_16276,N_15131,N_15829);
or U16277 (N_16277,N_15592,N_15437);
and U16278 (N_16278,N_15325,N_15518);
xor U16279 (N_16279,N_15889,N_15994);
nor U16280 (N_16280,N_15615,N_15171);
or U16281 (N_16281,N_15806,N_15557);
or U16282 (N_16282,N_15885,N_15073);
nand U16283 (N_16283,N_15339,N_15928);
or U16284 (N_16284,N_15078,N_15235);
nand U16285 (N_16285,N_15816,N_15264);
or U16286 (N_16286,N_15195,N_15388);
nor U16287 (N_16287,N_15770,N_15577);
nor U16288 (N_16288,N_15213,N_15805);
nor U16289 (N_16289,N_15909,N_15380);
xnor U16290 (N_16290,N_15469,N_15083);
nand U16291 (N_16291,N_15849,N_15822);
and U16292 (N_16292,N_15391,N_15008);
or U16293 (N_16293,N_15559,N_15826);
or U16294 (N_16294,N_15794,N_15407);
nor U16295 (N_16295,N_15155,N_15904);
xor U16296 (N_16296,N_15505,N_15284);
and U16297 (N_16297,N_15769,N_15363);
xnor U16298 (N_16298,N_15967,N_15182);
and U16299 (N_16299,N_15189,N_15730);
xor U16300 (N_16300,N_15023,N_15556);
nor U16301 (N_16301,N_15937,N_15933);
and U16302 (N_16302,N_15212,N_15951);
nand U16303 (N_16303,N_15322,N_15598);
xor U16304 (N_16304,N_15176,N_15934);
nor U16305 (N_16305,N_15487,N_15618);
xnor U16306 (N_16306,N_15698,N_15313);
nor U16307 (N_16307,N_15334,N_15055);
xor U16308 (N_16308,N_15386,N_15961);
nor U16309 (N_16309,N_15172,N_15286);
and U16310 (N_16310,N_15383,N_15310);
nand U16311 (N_16311,N_15056,N_15429);
nand U16312 (N_16312,N_15106,N_15297);
nand U16313 (N_16313,N_15316,N_15931);
nand U16314 (N_16314,N_15315,N_15580);
xor U16315 (N_16315,N_15306,N_15499);
xnor U16316 (N_16316,N_15681,N_15302);
nand U16317 (N_16317,N_15024,N_15977);
nand U16318 (N_16318,N_15780,N_15636);
nor U16319 (N_16319,N_15821,N_15136);
or U16320 (N_16320,N_15602,N_15201);
or U16321 (N_16321,N_15197,N_15054);
nand U16322 (N_16322,N_15148,N_15500);
nor U16323 (N_16323,N_15767,N_15485);
xnor U16324 (N_16324,N_15768,N_15778);
nor U16325 (N_16325,N_15050,N_15520);
xnor U16326 (N_16326,N_15986,N_15374);
or U16327 (N_16327,N_15012,N_15072);
nor U16328 (N_16328,N_15631,N_15224);
or U16329 (N_16329,N_15666,N_15941);
nor U16330 (N_16330,N_15524,N_15719);
xor U16331 (N_16331,N_15052,N_15675);
nor U16332 (N_16332,N_15369,N_15331);
nor U16333 (N_16333,N_15412,N_15553);
nor U16334 (N_16334,N_15600,N_15084);
xnor U16335 (N_16335,N_15975,N_15231);
nand U16336 (N_16336,N_15963,N_15237);
nor U16337 (N_16337,N_15194,N_15582);
or U16338 (N_16338,N_15861,N_15494);
or U16339 (N_16339,N_15611,N_15735);
nand U16340 (N_16340,N_15319,N_15724);
or U16341 (N_16341,N_15858,N_15751);
and U16342 (N_16342,N_15219,N_15970);
and U16343 (N_16343,N_15491,N_15790);
and U16344 (N_16344,N_15110,N_15460);
xnor U16345 (N_16345,N_15782,N_15153);
xnor U16346 (N_16346,N_15016,N_15357);
xor U16347 (N_16347,N_15337,N_15810);
or U16348 (N_16348,N_15562,N_15192);
or U16349 (N_16349,N_15142,N_15218);
and U16350 (N_16350,N_15662,N_15737);
or U16351 (N_16351,N_15787,N_15900);
nand U16352 (N_16352,N_15158,N_15273);
or U16353 (N_16353,N_15555,N_15614);
and U16354 (N_16354,N_15483,N_15180);
or U16355 (N_16355,N_15703,N_15191);
xor U16356 (N_16356,N_15134,N_15607);
nor U16357 (N_16357,N_15797,N_15292);
xor U16358 (N_16358,N_15537,N_15031);
and U16359 (N_16359,N_15415,N_15268);
xnor U16360 (N_16360,N_15196,N_15747);
xor U16361 (N_16361,N_15710,N_15252);
or U16362 (N_16362,N_15651,N_15444);
nor U16363 (N_16363,N_15879,N_15321);
nor U16364 (N_16364,N_15283,N_15452);
and U16365 (N_16365,N_15578,N_15916);
or U16366 (N_16366,N_15222,N_15807);
nor U16367 (N_16367,N_15150,N_15351);
or U16368 (N_16368,N_15837,N_15101);
xor U16369 (N_16369,N_15992,N_15090);
nand U16370 (N_16370,N_15663,N_15367);
xor U16371 (N_16371,N_15523,N_15355);
and U16372 (N_16372,N_15420,N_15620);
xor U16373 (N_16373,N_15360,N_15042);
or U16374 (N_16374,N_15432,N_15948);
xnor U16375 (N_16375,N_15973,N_15269);
or U16376 (N_16376,N_15068,N_15606);
nand U16377 (N_16377,N_15774,N_15554);
xnor U16378 (N_16378,N_15705,N_15066);
nand U16379 (N_16379,N_15964,N_15203);
or U16380 (N_16380,N_15568,N_15233);
nand U16381 (N_16381,N_15287,N_15184);
xor U16382 (N_16382,N_15094,N_15785);
xnor U16383 (N_16383,N_15096,N_15576);
nand U16384 (N_16384,N_15010,N_15811);
nand U16385 (N_16385,N_15552,N_15605);
xnor U16386 (N_16386,N_15299,N_15542);
nand U16387 (N_16387,N_15616,N_15624);
xor U16388 (N_16388,N_15619,N_15955);
or U16389 (N_16389,N_15280,N_15723);
and U16390 (N_16390,N_15036,N_15247);
nor U16391 (N_16391,N_15296,N_15982);
xor U16392 (N_16392,N_15832,N_15892);
nor U16393 (N_16393,N_15536,N_15239);
or U16394 (N_16394,N_15414,N_15236);
nand U16395 (N_16395,N_15506,N_15833);
xor U16396 (N_16396,N_15484,N_15385);
and U16397 (N_16397,N_15834,N_15112);
nand U16398 (N_16398,N_15265,N_15327);
or U16399 (N_16399,N_15870,N_15041);
nand U16400 (N_16400,N_15855,N_15272);
xor U16401 (N_16401,N_15962,N_15450);
or U16402 (N_16402,N_15279,N_15368);
nor U16403 (N_16403,N_15051,N_15141);
nor U16404 (N_16404,N_15467,N_15417);
nor U16405 (N_16405,N_15193,N_15749);
and U16406 (N_16406,N_15632,N_15658);
and U16407 (N_16407,N_15077,N_15910);
nor U16408 (N_16408,N_15464,N_15862);
nand U16409 (N_16409,N_15914,N_15186);
and U16410 (N_16410,N_15208,N_15907);
and U16411 (N_16411,N_15079,N_15852);
nand U16412 (N_16412,N_15198,N_15162);
and U16413 (N_16413,N_15594,N_15784);
nand U16414 (N_16414,N_15324,N_15708);
xnor U16415 (N_16415,N_15971,N_15496);
and U16416 (N_16416,N_15480,N_15242);
nor U16417 (N_16417,N_15721,N_15796);
nor U16418 (N_16418,N_15362,N_15125);
nand U16419 (N_16419,N_15633,N_15301);
or U16420 (N_16420,N_15105,N_15913);
or U16421 (N_16421,N_15800,N_15622);
nand U16422 (N_16422,N_15109,N_15856);
nor U16423 (N_16423,N_15854,N_15029);
xnor U16424 (N_16424,N_15891,N_15007);
or U16425 (N_16425,N_15478,N_15366);
or U16426 (N_16426,N_15230,N_15173);
nor U16427 (N_16427,N_15626,N_15183);
or U16428 (N_16428,N_15700,N_15733);
nor U16429 (N_16429,N_15628,N_15375);
xnor U16430 (N_16430,N_15664,N_15644);
or U16431 (N_16431,N_15167,N_15503);
xor U16432 (N_16432,N_15225,N_15570);
and U16433 (N_16433,N_15760,N_15739);
and U16434 (N_16434,N_15764,N_15170);
xnor U16435 (N_16435,N_15100,N_15526);
and U16436 (N_16436,N_15690,N_15669);
or U16437 (N_16437,N_15021,N_15843);
nand U16438 (N_16438,N_15185,N_15527);
nor U16439 (N_16439,N_15678,N_15936);
or U16440 (N_16440,N_15135,N_15411);
nand U16441 (N_16441,N_15116,N_15530);
or U16442 (N_16442,N_15032,N_15759);
and U16443 (N_16443,N_15604,N_15534);
and U16444 (N_16444,N_15174,N_15128);
xnor U16445 (N_16445,N_15828,N_15132);
nor U16446 (N_16446,N_15245,N_15006);
and U16447 (N_16447,N_15946,N_15850);
nand U16448 (N_16448,N_15804,N_15115);
xnor U16449 (N_16449,N_15151,N_15081);
xnor U16450 (N_16450,N_15419,N_15276);
xnor U16451 (N_16451,N_15741,N_15187);
and U16452 (N_16452,N_15289,N_15689);
nor U16453 (N_16453,N_15288,N_15433);
nand U16454 (N_16454,N_15729,N_15399);
xnor U16455 (N_16455,N_15507,N_15048);
nor U16456 (N_16456,N_15333,N_15972);
xnor U16457 (N_16457,N_15902,N_15199);
or U16458 (N_16458,N_15634,N_15957);
nand U16459 (N_16459,N_15541,N_15671);
and U16460 (N_16460,N_15282,N_15335);
nor U16461 (N_16461,N_15305,N_15240);
nor U16462 (N_16462,N_15779,N_15674);
xor U16463 (N_16463,N_15998,N_15140);
and U16464 (N_16464,N_15127,N_15020);
nor U16465 (N_16465,N_15985,N_15234);
and U16466 (N_16466,N_15569,N_15075);
or U16467 (N_16467,N_15133,N_15645);
xor U16468 (N_16468,N_15895,N_15845);
nor U16469 (N_16469,N_15040,N_15511);
nand U16470 (N_16470,N_15352,N_15864);
xnor U16471 (N_16471,N_15976,N_15017);
or U16472 (N_16472,N_15340,N_15771);
xor U16473 (N_16473,N_15293,N_15349);
or U16474 (N_16474,N_15227,N_15660);
or U16475 (N_16475,N_15014,N_15544);
xnor U16476 (N_16476,N_15640,N_15379);
nor U16477 (N_16477,N_15270,N_15687);
nand U16478 (N_16478,N_15758,N_15938);
nor U16479 (N_16479,N_15157,N_15274);
and U16480 (N_16480,N_15103,N_15597);
nand U16481 (N_16481,N_15750,N_15820);
nand U16482 (N_16482,N_15248,N_15320);
and U16483 (N_16483,N_15256,N_15092);
nor U16484 (N_16484,N_15529,N_15493);
nand U16485 (N_16485,N_15053,N_15348);
nor U16486 (N_16486,N_15835,N_15929);
and U16487 (N_16487,N_15479,N_15888);
nand U16488 (N_16488,N_15259,N_15560);
xor U16489 (N_16489,N_15566,N_15652);
or U16490 (N_16490,N_15177,N_15082);
and U16491 (N_16491,N_15482,N_15070);
or U16492 (N_16492,N_15490,N_15486);
xor U16493 (N_16493,N_15122,N_15445);
nor U16494 (N_16494,N_15960,N_15303);
nand U16495 (N_16495,N_15638,N_15271);
nand U16496 (N_16496,N_15906,N_15830);
nand U16497 (N_16497,N_15650,N_15793);
and U16498 (N_16498,N_15290,N_15752);
xnor U16499 (N_16499,N_15454,N_15514);
or U16500 (N_16500,N_15507,N_15727);
xor U16501 (N_16501,N_15884,N_15465);
nand U16502 (N_16502,N_15743,N_15392);
nand U16503 (N_16503,N_15898,N_15324);
nand U16504 (N_16504,N_15303,N_15504);
xor U16505 (N_16505,N_15158,N_15334);
nand U16506 (N_16506,N_15899,N_15043);
xor U16507 (N_16507,N_15986,N_15499);
and U16508 (N_16508,N_15495,N_15022);
or U16509 (N_16509,N_15614,N_15563);
xnor U16510 (N_16510,N_15893,N_15979);
nor U16511 (N_16511,N_15048,N_15615);
or U16512 (N_16512,N_15018,N_15705);
or U16513 (N_16513,N_15233,N_15094);
nand U16514 (N_16514,N_15084,N_15892);
nand U16515 (N_16515,N_15217,N_15672);
xor U16516 (N_16516,N_15696,N_15169);
nor U16517 (N_16517,N_15706,N_15488);
nor U16518 (N_16518,N_15823,N_15029);
nand U16519 (N_16519,N_15288,N_15693);
nand U16520 (N_16520,N_15057,N_15563);
and U16521 (N_16521,N_15127,N_15616);
nand U16522 (N_16522,N_15730,N_15497);
nor U16523 (N_16523,N_15363,N_15630);
nand U16524 (N_16524,N_15186,N_15599);
or U16525 (N_16525,N_15009,N_15101);
xnor U16526 (N_16526,N_15605,N_15267);
nor U16527 (N_16527,N_15424,N_15803);
xnor U16528 (N_16528,N_15872,N_15972);
xor U16529 (N_16529,N_15713,N_15472);
xnor U16530 (N_16530,N_15269,N_15768);
nor U16531 (N_16531,N_15163,N_15364);
xor U16532 (N_16532,N_15617,N_15181);
xor U16533 (N_16533,N_15387,N_15037);
nor U16534 (N_16534,N_15262,N_15098);
or U16535 (N_16535,N_15748,N_15833);
and U16536 (N_16536,N_15394,N_15885);
xnor U16537 (N_16537,N_15706,N_15937);
and U16538 (N_16538,N_15328,N_15403);
or U16539 (N_16539,N_15485,N_15589);
or U16540 (N_16540,N_15593,N_15165);
nor U16541 (N_16541,N_15314,N_15641);
xor U16542 (N_16542,N_15724,N_15381);
and U16543 (N_16543,N_15454,N_15127);
or U16544 (N_16544,N_15893,N_15389);
or U16545 (N_16545,N_15665,N_15772);
nor U16546 (N_16546,N_15014,N_15729);
and U16547 (N_16547,N_15472,N_15244);
nor U16548 (N_16548,N_15591,N_15111);
or U16549 (N_16549,N_15328,N_15672);
or U16550 (N_16550,N_15790,N_15058);
xnor U16551 (N_16551,N_15994,N_15283);
nor U16552 (N_16552,N_15531,N_15932);
xnor U16553 (N_16553,N_15537,N_15652);
or U16554 (N_16554,N_15080,N_15946);
xor U16555 (N_16555,N_15092,N_15894);
or U16556 (N_16556,N_15907,N_15540);
nand U16557 (N_16557,N_15277,N_15203);
and U16558 (N_16558,N_15610,N_15020);
xnor U16559 (N_16559,N_15950,N_15358);
and U16560 (N_16560,N_15432,N_15081);
xor U16561 (N_16561,N_15282,N_15285);
nand U16562 (N_16562,N_15526,N_15421);
nand U16563 (N_16563,N_15033,N_15142);
xnor U16564 (N_16564,N_15841,N_15424);
xor U16565 (N_16565,N_15383,N_15594);
xor U16566 (N_16566,N_15503,N_15339);
and U16567 (N_16567,N_15434,N_15528);
or U16568 (N_16568,N_15655,N_15788);
or U16569 (N_16569,N_15378,N_15081);
or U16570 (N_16570,N_15265,N_15733);
xnor U16571 (N_16571,N_15270,N_15596);
nor U16572 (N_16572,N_15997,N_15597);
xor U16573 (N_16573,N_15302,N_15127);
or U16574 (N_16574,N_15013,N_15307);
or U16575 (N_16575,N_15330,N_15006);
nor U16576 (N_16576,N_15049,N_15577);
and U16577 (N_16577,N_15693,N_15910);
and U16578 (N_16578,N_15736,N_15448);
or U16579 (N_16579,N_15234,N_15028);
nand U16580 (N_16580,N_15595,N_15039);
and U16581 (N_16581,N_15143,N_15979);
and U16582 (N_16582,N_15412,N_15001);
or U16583 (N_16583,N_15122,N_15960);
nand U16584 (N_16584,N_15938,N_15041);
and U16585 (N_16585,N_15120,N_15734);
nor U16586 (N_16586,N_15789,N_15886);
nand U16587 (N_16587,N_15383,N_15393);
nand U16588 (N_16588,N_15020,N_15264);
xnor U16589 (N_16589,N_15213,N_15151);
and U16590 (N_16590,N_15700,N_15549);
and U16591 (N_16591,N_15387,N_15952);
nor U16592 (N_16592,N_15154,N_15498);
nor U16593 (N_16593,N_15378,N_15124);
or U16594 (N_16594,N_15963,N_15970);
and U16595 (N_16595,N_15198,N_15343);
or U16596 (N_16596,N_15215,N_15310);
nand U16597 (N_16597,N_15409,N_15279);
nor U16598 (N_16598,N_15602,N_15060);
xor U16599 (N_16599,N_15861,N_15483);
or U16600 (N_16600,N_15197,N_15424);
nor U16601 (N_16601,N_15026,N_15081);
xor U16602 (N_16602,N_15260,N_15630);
and U16603 (N_16603,N_15931,N_15739);
xor U16604 (N_16604,N_15427,N_15544);
nand U16605 (N_16605,N_15358,N_15355);
xor U16606 (N_16606,N_15863,N_15998);
nand U16607 (N_16607,N_15793,N_15546);
nand U16608 (N_16608,N_15932,N_15632);
or U16609 (N_16609,N_15340,N_15767);
xnor U16610 (N_16610,N_15549,N_15206);
nand U16611 (N_16611,N_15593,N_15060);
xnor U16612 (N_16612,N_15263,N_15636);
or U16613 (N_16613,N_15502,N_15245);
nor U16614 (N_16614,N_15316,N_15086);
nand U16615 (N_16615,N_15418,N_15031);
xnor U16616 (N_16616,N_15055,N_15942);
or U16617 (N_16617,N_15661,N_15373);
xor U16618 (N_16618,N_15058,N_15022);
and U16619 (N_16619,N_15883,N_15301);
nand U16620 (N_16620,N_15333,N_15273);
and U16621 (N_16621,N_15252,N_15763);
or U16622 (N_16622,N_15054,N_15435);
nor U16623 (N_16623,N_15379,N_15207);
or U16624 (N_16624,N_15951,N_15199);
and U16625 (N_16625,N_15173,N_15858);
and U16626 (N_16626,N_15681,N_15987);
nor U16627 (N_16627,N_15905,N_15724);
and U16628 (N_16628,N_15456,N_15175);
nor U16629 (N_16629,N_15022,N_15193);
nor U16630 (N_16630,N_15137,N_15298);
nor U16631 (N_16631,N_15987,N_15701);
xnor U16632 (N_16632,N_15092,N_15703);
xor U16633 (N_16633,N_15387,N_15014);
and U16634 (N_16634,N_15921,N_15772);
xnor U16635 (N_16635,N_15112,N_15396);
nand U16636 (N_16636,N_15328,N_15773);
xnor U16637 (N_16637,N_15771,N_15063);
xor U16638 (N_16638,N_15041,N_15554);
or U16639 (N_16639,N_15102,N_15161);
nor U16640 (N_16640,N_15006,N_15358);
or U16641 (N_16641,N_15279,N_15215);
or U16642 (N_16642,N_15705,N_15072);
nor U16643 (N_16643,N_15522,N_15755);
nor U16644 (N_16644,N_15201,N_15645);
nand U16645 (N_16645,N_15770,N_15963);
or U16646 (N_16646,N_15198,N_15428);
nor U16647 (N_16647,N_15057,N_15496);
nand U16648 (N_16648,N_15168,N_15563);
xor U16649 (N_16649,N_15711,N_15855);
or U16650 (N_16650,N_15356,N_15961);
nand U16651 (N_16651,N_15431,N_15574);
and U16652 (N_16652,N_15833,N_15365);
and U16653 (N_16653,N_15900,N_15609);
nand U16654 (N_16654,N_15265,N_15986);
nor U16655 (N_16655,N_15021,N_15582);
nand U16656 (N_16656,N_15360,N_15731);
or U16657 (N_16657,N_15500,N_15933);
nor U16658 (N_16658,N_15000,N_15688);
or U16659 (N_16659,N_15292,N_15021);
or U16660 (N_16660,N_15570,N_15875);
and U16661 (N_16661,N_15378,N_15025);
and U16662 (N_16662,N_15049,N_15259);
xnor U16663 (N_16663,N_15746,N_15283);
xor U16664 (N_16664,N_15455,N_15370);
and U16665 (N_16665,N_15432,N_15530);
nand U16666 (N_16666,N_15787,N_15395);
or U16667 (N_16667,N_15782,N_15772);
xor U16668 (N_16668,N_15860,N_15047);
nand U16669 (N_16669,N_15664,N_15574);
or U16670 (N_16670,N_15332,N_15337);
or U16671 (N_16671,N_15222,N_15903);
or U16672 (N_16672,N_15858,N_15754);
nor U16673 (N_16673,N_15465,N_15876);
nand U16674 (N_16674,N_15027,N_15509);
nand U16675 (N_16675,N_15996,N_15923);
xnor U16676 (N_16676,N_15085,N_15436);
nand U16677 (N_16677,N_15858,N_15107);
xor U16678 (N_16678,N_15219,N_15680);
xnor U16679 (N_16679,N_15170,N_15206);
xnor U16680 (N_16680,N_15043,N_15449);
and U16681 (N_16681,N_15323,N_15616);
and U16682 (N_16682,N_15671,N_15399);
nor U16683 (N_16683,N_15243,N_15720);
xor U16684 (N_16684,N_15574,N_15285);
nand U16685 (N_16685,N_15370,N_15172);
xnor U16686 (N_16686,N_15752,N_15713);
or U16687 (N_16687,N_15707,N_15711);
nor U16688 (N_16688,N_15449,N_15558);
or U16689 (N_16689,N_15444,N_15322);
or U16690 (N_16690,N_15339,N_15867);
xnor U16691 (N_16691,N_15753,N_15003);
nor U16692 (N_16692,N_15870,N_15690);
nor U16693 (N_16693,N_15546,N_15701);
and U16694 (N_16694,N_15131,N_15901);
or U16695 (N_16695,N_15030,N_15403);
or U16696 (N_16696,N_15628,N_15107);
nand U16697 (N_16697,N_15630,N_15780);
nand U16698 (N_16698,N_15409,N_15959);
xor U16699 (N_16699,N_15852,N_15696);
nand U16700 (N_16700,N_15729,N_15914);
nor U16701 (N_16701,N_15158,N_15836);
nor U16702 (N_16702,N_15902,N_15618);
and U16703 (N_16703,N_15048,N_15025);
nand U16704 (N_16704,N_15961,N_15068);
or U16705 (N_16705,N_15389,N_15757);
or U16706 (N_16706,N_15747,N_15868);
xnor U16707 (N_16707,N_15933,N_15246);
or U16708 (N_16708,N_15575,N_15227);
xnor U16709 (N_16709,N_15222,N_15307);
nand U16710 (N_16710,N_15343,N_15148);
and U16711 (N_16711,N_15977,N_15621);
nor U16712 (N_16712,N_15639,N_15816);
nand U16713 (N_16713,N_15284,N_15795);
and U16714 (N_16714,N_15880,N_15643);
xnor U16715 (N_16715,N_15956,N_15910);
or U16716 (N_16716,N_15024,N_15213);
and U16717 (N_16717,N_15556,N_15326);
and U16718 (N_16718,N_15077,N_15506);
xnor U16719 (N_16719,N_15133,N_15308);
nand U16720 (N_16720,N_15422,N_15761);
xor U16721 (N_16721,N_15791,N_15630);
and U16722 (N_16722,N_15977,N_15631);
and U16723 (N_16723,N_15155,N_15874);
and U16724 (N_16724,N_15720,N_15189);
nand U16725 (N_16725,N_15000,N_15901);
nand U16726 (N_16726,N_15416,N_15355);
nor U16727 (N_16727,N_15579,N_15827);
or U16728 (N_16728,N_15182,N_15131);
and U16729 (N_16729,N_15063,N_15287);
xor U16730 (N_16730,N_15549,N_15182);
nand U16731 (N_16731,N_15669,N_15240);
nor U16732 (N_16732,N_15072,N_15508);
and U16733 (N_16733,N_15857,N_15743);
or U16734 (N_16734,N_15243,N_15269);
xnor U16735 (N_16735,N_15764,N_15829);
or U16736 (N_16736,N_15785,N_15330);
xor U16737 (N_16737,N_15337,N_15437);
nor U16738 (N_16738,N_15858,N_15144);
xor U16739 (N_16739,N_15051,N_15048);
xnor U16740 (N_16740,N_15320,N_15624);
nand U16741 (N_16741,N_15044,N_15952);
nand U16742 (N_16742,N_15415,N_15364);
nand U16743 (N_16743,N_15655,N_15460);
or U16744 (N_16744,N_15091,N_15556);
nor U16745 (N_16745,N_15528,N_15361);
and U16746 (N_16746,N_15955,N_15949);
nand U16747 (N_16747,N_15254,N_15281);
nand U16748 (N_16748,N_15395,N_15243);
and U16749 (N_16749,N_15748,N_15657);
or U16750 (N_16750,N_15013,N_15006);
nor U16751 (N_16751,N_15654,N_15010);
xnor U16752 (N_16752,N_15244,N_15160);
nand U16753 (N_16753,N_15344,N_15462);
nand U16754 (N_16754,N_15622,N_15325);
xnor U16755 (N_16755,N_15558,N_15399);
xnor U16756 (N_16756,N_15304,N_15686);
and U16757 (N_16757,N_15291,N_15631);
nand U16758 (N_16758,N_15258,N_15494);
nand U16759 (N_16759,N_15818,N_15594);
nand U16760 (N_16760,N_15109,N_15407);
nor U16761 (N_16761,N_15231,N_15618);
and U16762 (N_16762,N_15362,N_15248);
and U16763 (N_16763,N_15391,N_15784);
xor U16764 (N_16764,N_15393,N_15370);
nor U16765 (N_16765,N_15154,N_15056);
nor U16766 (N_16766,N_15945,N_15352);
xnor U16767 (N_16767,N_15739,N_15935);
nor U16768 (N_16768,N_15757,N_15038);
nand U16769 (N_16769,N_15284,N_15900);
and U16770 (N_16770,N_15386,N_15915);
xor U16771 (N_16771,N_15779,N_15861);
xnor U16772 (N_16772,N_15558,N_15977);
and U16773 (N_16773,N_15467,N_15190);
and U16774 (N_16774,N_15733,N_15691);
or U16775 (N_16775,N_15683,N_15560);
xnor U16776 (N_16776,N_15814,N_15737);
nor U16777 (N_16777,N_15676,N_15105);
nor U16778 (N_16778,N_15052,N_15747);
nor U16779 (N_16779,N_15348,N_15097);
or U16780 (N_16780,N_15903,N_15012);
and U16781 (N_16781,N_15871,N_15447);
and U16782 (N_16782,N_15298,N_15595);
or U16783 (N_16783,N_15051,N_15510);
or U16784 (N_16784,N_15133,N_15618);
nand U16785 (N_16785,N_15107,N_15485);
xnor U16786 (N_16786,N_15117,N_15676);
nor U16787 (N_16787,N_15460,N_15328);
and U16788 (N_16788,N_15498,N_15939);
nand U16789 (N_16789,N_15028,N_15588);
nand U16790 (N_16790,N_15719,N_15267);
nand U16791 (N_16791,N_15524,N_15335);
and U16792 (N_16792,N_15245,N_15022);
nor U16793 (N_16793,N_15816,N_15851);
nand U16794 (N_16794,N_15890,N_15503);
nor U16795 (N_16795,N_15270,N_15312);
nand U16796 (N_16796,N_15230,N_15107);
and U16797 (N_16797,N_15958,N_15880);
nand U16798 (N_16798,N_15265,N_15465);
nand U16799 (N_16799,N_15528,N_15858);
xor U16800 (N_16800,N_15559,N_15111);
xor U16801 (N_16801,N_15352,N_15306);
xor U16802 (N_16802,N_15050,N_15708);
xor U16803 (N_16803,N_15678,N_15159);
and U16804 (N_16804,N_15013,N_15887);
and U16805 (N_16805,N_15936,N_15625);
and U16806 (N_16806,N_15470,N_15766);
xor U16807 (N_16807,N_15321,N_15535);
and U16808 (N_16808,N_15157,N_15949);
or U16809 (N_16809,N_15323,N_15866);
and U16810 (N_16810,N_15636,N_15288);
nor U16811 (N_16811,N_15350,N_15340);
xor U16812 (N_16812,N_15316,N_15860);
xor U16813 (N_16813,N_15033,N_15900);
and U16814 (N_16814,N_15839,N_15270);
xor U16815 (N_16815,N_15815,N_15429);
nor U16816 (N_16816,N_15000,N_15864);
or U16817 (N_16817,N_15238,N_15786);
xnor U16818 (N_16818,N_15482,N_15327);
nor U16819 (N_16819,N_15803,N_15038);
nand U16820 (N_16820,N_15312,N_15483);
or U16821 (N_16821,N_15645,N_15376);
xnor U16822 (N_16822,N_15910,N_15741);
and U16823 (N_16823,N_15956,N_15678);
nand U16824 (N_16824,N_15900,N_15584);
or U16825 (N_16825,N_15492,N_15517);
xnor U16826 (N_16826,N_15882,N_15777);
nand U16827 (N_16827,N_15226,N_15159);
nor U16828 (N_16828,N_15065,N_15539);
nor U16829 (N_16829,N_15982,N_15447);
nor U16830 (N_16830,N_15961,N_15997);
nand U16831 (N_16831,N_15029,N_15778);
nor U16832 (N_16832,N_15668,N_15167);
and U16833 (N_16833,N_15927,N_15420);
or U16834 (N_16834,N_15090,N_15274);
nor U16835 (N_16835,N_15764,N_15615);
nor U16836 (N_16836,N_15532,N_15695);
nand U16837 (N_16837,N_15974,N_15677);
nand U16838 (N_16838,N_15228,N_15344);
and U16839 (N_16839,N_15352,N_15179);
nor U16840 (N_16840,N_15776,N_15220);
nand U16841 (N_16841,N_15054,N_15458);
nand U16842 (N_16842,N_15681,N_15840);
nand U16843 (N_16843,N_15064,N_15316);
nand U16844 (N_16844,N_15869,N_15917);
or U16845 (N_16845,N_15439,N_15699);
xnor U16846 (N_16846,N_15129,N_15642);
nor U16847 (N_16847,N_15521,N_15923);
nor U16848 (N_16848,N_15218,N_15099);
xnor U16849 (N_16849,N_15231,N_15440);
nor U16850 (N_16850,N_15175,N_15677);
nor U16851 (N_16851,N_15712,N_15045);
nand U16852 (N_16852,N_15602,N_15087);
nor U16853 (N_16853,N_15426,N_15086);
xor U16854 (N_16854,N_15005,N_15073);
or U16855 (N_16855,N_15373,N_15362);
xor U16856 (N_16856,N_15319,N_15692);
xor U16857 (N_16857,N_15909,N_15160);
and U16858 (N_16858,N_15282,N_15413);
nand U16859 (N_16859,N_15804,N_15479);
nand U16860 (N_16860,N_15969,N_15559);
nand U16861 (N_16861,N_15775,N_15066);
xnor U16862 (N_16862,N_15517,N_15652);
and U16863 (N_16863,N_15356,N_15877);
nand U16864 (N_16864,N_15549,N_15608);
xor U16865 (N_16865,N_15260,N_15795);
nand U16866 (N_16866,N_15962,N_15455);
xnor U16867 (N_16867,N_15507,N_15803);
or U16868 (N_16868,N_15025,N_15715);
or U16869 (N_16869,N_15938,N_15510);
or U16870 (N_16870,N_15269,N_15328);
xnor U16871 (N_16871,N_15028,N_15195);
or U16872 (N_16872,N_15815,N_15933);
nand U16873 (N_16873,N_15606,N_15150);
nor U16874 (N_16874,N_15065,N_15788);
nor U16875 (N_16875,N_15958,N_15807);
nor U16876 (N_16876,N_15355,N_15054);
xnor U16877 (N_16877,N_15616,N_15806);
and U16878 (N_16878,N_15150,N_15947);
nand U16879 (N_16879,N_15696,N_15017);
nand U16880 (N_16880,N_15576,N_15142);
or U16881 (N_16881,N_15437,N_15631);
or U16882 (N_16882,N_15513,N_15591);
xor U16883 (N_16883,N_15835,N_15976);
nand U16884 (N_16884,N_15832,N_15533);
or U16885 (N_16885,N_15426,N_15431);
nor U16886 (N_16886,N_15412,N_15164);
nand U16887 (N_16887,N_15321,N_15104);
or U16888 (N_16888,N_15306,N_15433);
nand U16889 (N_16889,N_15286,N_15546);
or U16890 (N_16890,N_15031,N_15806);
nand U16891 (N_16891,N_15778,N_15231);
nor U16892 (N_16892,N_15477,N_15390);
nor U16893 (N_16893,N_15602,N_15744);
xnor U16894 (N_16894,N_15071,N_15113);
and U16895 (N_16895,N_15660,N_15292);
or U16896 (N_16896,N_15243,N_15467);
and U16897 (N_16897,N_15451,N_15024);
xnor U16898 (N_16898,N_15922,N_15566);
and U16899 (N_16899,N_15127,N_15071);
xor U16900 (N_16900,N_15503,N_15091);
or U16901 (N_16901,N_15484,N_15697);
or U16902 (N_16902,N_15967,N_15053);
xnor U16903 (N_16903,N_15338,N_15141);
nor U16904 (N_16904,N_15423,N_15944);
and U16905 (N_16905,N_15916,N_15976);
nor U16906 (N_16906,N_15018,N_15661);
xor U16907 (N_16907,N_15007,N_15152);
nor U16908 (N_16908,N_15573,N_15731);
nand U16909 (N_16909,N_15649,N_15345);
nand U16910 (N_16910,N_15706,N_15180);
nand U16911 (N_16911,N_15365,N_15804);
xor U16912 (N_16912,N_15153,N_15030);
nor U16913 (N_16913,N_15979,N_15547);
nor U16914 (N_16914,N_15485,N_15154);
xnor U16915 (N_16915,N_15335,N_15780);
and U16916 (N_16916,N_15799,N_15241);
nand U16917 (N_16917,N_15235,N_15524);
or U16918 (N_16918,N_15625,N_15032);
and U16919 (N_16919,N_15370,N_15910);
nand U16920 (N_16920,N_15293,N_15587);
nand U16921 (N_16921,N_15941,N_15555);
and U16922 (N_16922,N_15110,N_15790);
xor U16923 (N_16923,N_15886,N_15485);
nor U16924 (N_16924,N_15905,N_15211);
or U16925 (N_16925,N_15223,N_15488);
xnor U16926 (N_16926,N_15320,N_15061);
and U16927 (N_16927,N_15090,N_15533);
xnor U16928 (N_16928,N_15628,N_15606);
and U16929 (N_16929,N_15721,N_15824);
or U16930 (N_16930,N_15726,N_15899);
nor U16931 (N_16931,N_15122,N_15330);
xnor U16932 (N_16932,N_15670,N_15336);
and U16933 (N_16933,N_15092,N_15841);
nor U16934 (N_16934,N_15843,N_15923);
nor U16935 (N_16935,N_15829,N_15246);
and U16936 (N_16936,N_15503,N_15291);
or U16937 (N_16937,N_15683,N_15483);
nand U16938 (N_16938,N_15924,N_15124);
nand U16939 (N_16939,N_15933,N_15292);
nor U16940 (N_16940,N_15911,N_15228);
or U16941 (N_16941,N_15503,N_15980);
and U16942 (N_16942,N_15983,N_15135);
xor U16943 (N_16943,N_15743,N_15711);
xnor U16944 (N_16944,N_15449,N_15902);
nor U16945 (N_16945,N_15182,N_15930);
or U16946 (N_16946,N_15473,N_15565);
nand U16947 (N_16947,N_15980,N_15473);
xor U16948 (N_16948,N_15753,N_15268);
and U16949 (N_16949,N_15078,N_15462);
or U16950 (N_16950,N_15277,N_15139);
nand U16951 (N_16951,N_15433,N_15127);
xnor U16952 (N_16952,N_15800,N_15212);
nand U16953 (N_16953,N_15128,N_15762);
or U16954 (N_16954,N_15989,N_15385);
nor U16955 (N_16955,N_15554,N_15074);
or U16956 (N_16956,N_15643,N_15392);
and U16957 (N_16957,N_15054,N_15665);
nor U16958 (N_16958,N_15426,N_15341);
and U16959 (N_16959,N_15744,N_15558);
xor U16960 (N_16960,N_15742,N_15436);
nor U16961 (N_16961,N_15014,N_15375);
xor U16962 (N_16962,N_15904,N_15362);
xnor U16963 (N_16963,N_15605,N_15491);
nor U16964 (N_16964,N_15753,N_15709);
nand U16965 (N_16965,N_15504,N_15280);
and U16966 (N_16966,N_15636,N_15403);
nor U16967 (N_16967,N_15486,N_15848);
nor U16968 (N_16968,N_15839,N_15050);
xnor U16969 (N_16969,N_15280,N_15875);
xor U16970 (N_16970,N_15092,N_15249);
and U16971 (N_16971,N_15064,N_15350);
and U16972 (N_16972,N_15831,N_15170);
nor U16973 (N_16973,N_15576,N_15530);
nor U16974 (N_16974,N_15561,N_15426);
and U16975 (N_16975,N_15672,N_15954);
and U16976 (N_16976,N_15052,N_15797);
and U16977 (N_16977,N_15268,N_15524);
or U16978 (N_16978,N_15611,N_15080);
or U16979 (N_16979,N_15057,N_15306);
xnor U16980 (N_16980,N_15538,N_15359);
nor U16981 (N_16981,N_15394,N_15347);
xor U16982 (N_16982,N_15316,N_15553);
nand U16983 (N_16983,N_15689,N_15850);
nor U16984 (N_16984,N_15356,N_15684);
nand U16985 (N_16985,N_15455,N_15099);
xnor U16986 (N_16986,N_15599,N_15176);
nor U16987 (N_16987,N_15700,N_15245);
or U16988 (N_16988,N_15575,N_15105);
xor U16989 (N_16989,N_15015,N_15011);
nand U16990 (N_16990,N_15017,N_15360);
or U16991 (N_16991,N_15037,N_15999);
nor U16992 (N_16992,N_15795,N_15534);
nor U16993 (N_16993,N_15483,N_15816);
xor U16994 (N_16994,N_15269,N_15163);
xor U16995 (N_16995,N_15959,N_15167);
xor U16996 (N_16996,N_15695,N_15548);
nor U16997 (N_16997,N_15997,N_15826);
xor U16998 (N_16998,N_15652,N_15749);
nand U16999 (N_16999,N_15398,N_15265);
nand U17000 (N_17000,N_16955,N_16912);
and U17001 (N_17001,N_16257,N_16684);
and U17002 (N_17002,N_16054,N_16458);
nand U17003 (N_17003,N_16068,N_16470);
nand U17004 (N_17004,N_16208,N_16891);
or U17005 (N_17005,N_16484,N_16393);
and U17006 (N_17006,N_16771,N_16143);
xnor U17007 (N_17007,N_16327,N_16827);
or U17008 (N_17008,N_16815,N_16959);
nand U17009 (N_17009,N_16564,N_16268);
nor U17010 (N_17010,N_16873,N_16700);
or U17011 (N_17011,N_16028,N_16274);
nand U17012 (N_17012,N_16292,N_16016);
xor U17013 (N_17013,N_16619,N_16301);
nor U17014 (N_17014,N_16222,N_16382);
xnor U17015 (N_17015,N_16371,N_16581);
xor U17016 (N_17016,N_16296,N_16090);
xor U17017 (N_17017,N_16536,N_16887);
or U17018 (N_17018,N_16389,N_16014);
xor U17019 (N_17019,N_16971,N_16018);
nor U17020 (N_17020,N_16084,N_16707);
nor U17021 (N_17021,N_16752,N_16788);
nand U17022 (N_17022,N_16246,N_16990);
xnor U17023 (N_17023,N_16892,N_16394);
nor U17024 (N_17024,N_16510,N_16778);
and U17025 (N_17025,N_16335,N_16854);
and U17026 (N_17026,N_16218,N_16286);
nand U17027 (N_17027,N_16639,N_16941);
or U17028 (N_17028,N_16341,N_16863);
nor U17029 (N_17029,N_16422,N_16079);
nand U17030 (N_17030,N_16099,N_16435);
nand U17031 (N_17031,N_16361,N_16997);
nor U17032 (N_17032,N_16660,N_16488);
nand U17033 (N_17033,N_16176,N_16939);
nor U17034 (N_17034,N_16649,N_16739);
xor U17035 (N_17035,N_16515,N_16708);
or U17036 (N_17036,N_16446,N_16272);
xnor U17037 (N_17037,N_16356,N_16240);
nand U17038 (N_17038,N_16231,N_16372);
or U17039 (N_17039,N_16126,N_16800);
nor U17040 (N_17040,N_16859,N_16075);
xnor U17041 (N_17041,N_16065,N_16751);
nand U17042 (N_17042,N_16091,N_16819);
nand U17043 (N_17043,N_16063,N_16532);
nand U17044 (N_17044,N_16541,N_16963);
xor U17045 (N_17045,N_16251,N_16576);
or U17046 (N_17046,N_16768,N_16669);
nand U17047 (N_17047,N_16683,N_16501);
nor U17048 (N_17048,N_16001,N_16159);
nand U17049 (N_17049,N_16685,N_16385);
nor U17050 (N_17050,N_16678,N_16588);
nor U17051 (N_17051,N_16643,N_16217);
xor U17052 (N_17052,N_16568,N_16799);
xnor U17053 (N_17053,N_16808,N_16517);
nand U17054 (N_17054,N_16293,N_16438);
and U17055 (N_17055,N_16627,N_16557);
and U17056 (N_17056,N_16009,N_16747);
nor U17057 (N_17057,N_16164,N_16424);
and U17058 (N_17058,N_16279,N_16182);
or U17059 (N_17059,N_16258,N_16718);
nor U17060 (N_17060,N_16158,N_16152);
nand U17061 (N_17061,N_16428,N_16480);
nand U17062 (N_17062,N_16053,N_16398);
or U17063 (N_17063,N_16093,N_16066);
xor U17064 (N_17064,N_16156,N_16642);
nor U17065 (N_17065,N_16374,N_16089);
nor U17066 (N_17066,N_16400,N_16304);
nand U17067 (N_17067,N_16448,N_16624);
nand U17068 (N_17068,N_16761,N_16161);
nor U17069 (N_17069,N_16326,N_16670);
nor U17070 (N_17070,N_16154,N_16601);
nor U17071 (N_17071,N_16559,N_16291);
or U17072 (N_17072,N_16205,N_16414);
nor U17073 (N_17073,N_16225,N_16665);
or U17074 (N_17074,N_16734,N_16062);
and U17075 (N_17075,N_16467,N_16828);
nand U17076 (N_17076,N_16937,N_16621);
or U17077 (N_17077,N_16620,N_16789);
nor U17078 (N_17078,N_16043,N_16691);
nand U17079 (N_17079,N_16946,N_16085);
xnor U17080 (N_17080,N_16648,N_16204);
nor U17081 (N_17081,N_16727,N_16267);
or U17082 (N_17082,N_16634,N_16364);
or U17083 (N_17083,N_16375,N_16726);
xnor U17084 (N_17084,N_16954,N_16917);
and U17085 (N_17085,N_16696,N_16106);
nor U17086 (N_17086,N_16216,N_16852);
xor U17087 (N_17087,N_16979,N_16798);
or U17088 (N_17088,N_16343,N_16901);
or U17089 (N_17089,N_16040,N_16922);
or U17090 (N_17090,N_16228,N_16010);
or U17091 (N_17091,N_16289,N_16472);
nand U17092 (N_17092,N_16022,N_16762);
nor U17093 (N_17093,N_16898,N_16452);
xnor U17094 (N_17094,N_16060,N_16931);
or U17095 (N_17095,N_16109,N_16038);
or U17096 (N_17096,N_16985,N_16369);
nand U17097 (N_17097,N_16548,N_16650);
and U17098 (N_17098,N_16655,N_16841);
xnor U17099 (N_17099,N_16129,N_16077);
and U17100 (N_17100,N_16482,N_16058);
or U17101 (N_17101,N_16810,N_16881);
and U17102 (N_17102,N_16411,N_16527);
xnor U17103 (N_17103,N_16008,N_16086);
nor U17104 (N_17104,N_16029,N_16554);
xnor U17105 (N_17105,N_16951,N_16600);
or U17106 (N_17106,N_16410,N_16584);
nand U17107 (N_17107,N_16239,N_16462);
nor U17108 (N_17108,N_16977,N_16212);
xnor U17109 (N_17109,N_16763,N_16637);
or U17110 (N_17110,N_16500,N_16992);
nand U17111 (N_17111,N_16057,N_16017);
xor U17112 (N_17112,N_16549,N_16174);
xor U17113 (N_17113,N_16839,N_16249);
or U17114 (N_17114,N_16888,N_16036);
and U17115 (N_17115,N_16704,N_16333);
xor U17116 (N_17116,N_16623,N_16594);
or U17117 (N_17117,N_16920,N_16150);
and U17118 (N_17118,N_16117,N_16321);
xor U17119 (N_17119,N_16965,N_16653);
nand U17120 (N_17120,N_16320,N_16439);
and U17121 (N_17121,N_16259,N_16538);
and U17122 (N_17122,N_16509,N_16000);
nand U17123 (N_17123,N_16816,N_16262);
nor U17124 (N_17124,N_16373,N_16983);
nor U17125 (N_17125,N_16599,N_16135);
nand U17126 (N_17126,N_16777,N_16365);
nand U17127 (N_17127,N_16319,N_16714);
or U17128 (N_17128,N_16459,N_16546);
nand U17129 (N_17129,N_16139,N_16247);
and U17130 (N_17130,N_16664,N_16284);
and U17131 (N_17131,N_16157,N_16197);
or U17132 (N_17132,N_16379,N_16406);
or U17133 (N_17133,N_16605,N_16189);
xor U17134 (N_17134,N_16641,N_16468);
or U17135 (N_17135,N_16672,N_16032);
nor U17136 (N_17136,N_16862,N_16717);
or U17137 (N_17137,N_16048,N_16840);
nor U17138 (N_17138,N_16449,N_16166);
nor U17139 (N_17139,N_16377,N_16072);
nor U17140 (N_17140,N_16146,N_16209);
xnor U17141 (N_17141,N_16957,N_16023);
xnor U17142 (N_17142,N_16388,N_16535);
and U17143 (N_17143,N_16116,N_16552);
xnor U17144 (N_17144,N_16577,N_16645);
nor U17145 (N_17145,N_16453,N_16812);
or U17146 (N_17146,N_16460,N_16354);
and U17147 (N_17147,N_16450,N_16211);
xor U17148 (N_17148,N_16323,N_16263);
nand U17149 (N_17149,N_16674,N_16041);
nor U17150 (N_17150,N_16442,N_16806);
or U17151 (N_17151,N_16591,N_16473);
xnor U17152 (N_17152,N_16408,N_16826);
or U17153 (N_17153,N_16945,N_16606);
nor U17154 (N_17154,N_16030,N_16094);
or U17155 (N_17155,N_16646,N_16252);
nand U17156 (N_17156,N_16631,N_16928);
nor U17157 (N_17157,N_16167,N_16451);
nand U17158 (N_17158,N_16050,N_16681);
nand U17159 (N_17159,N_16614,N_16870);
xor U17160 (N_17160,N_16926,N_16195);
nand U17161 (N_17161,N_16479,N_16082);
nand U17162 (N_17162,N_16316,N_16924);
nor U17163 (N_17163,N_16475,N_16556);
nand U17164 (N_17164,N_16677,N_16310);
nor U17165 (N_17165,N_16780,N_16656);
nor U17166 (N_17166,N_16224,N_16953);
nor U17167 (N_17167,N_16942,N_16322);
xor U17168 (N_17168,N_16144,N_16698);
xor U17169 (N_17169,N_16261,N_16513);
and U17170 (N_17170,N_16330,N_16851);
and U17171 (N_17171,N_16002,N_16366);
and U17172 (N_17172,N_16838,N_16313);
xnor U17173 (N_17173,N_16709,N_16431);
xnor U17174 (N_17174,N_16007,N_16555);
xor U17175 (N_17175,N_16046,N_16042);
nor U17176 (N_17176,N_16171,N_16429);
or U17177 (N_17177,N_16626,N_16914);
nand U17178 (N_17178,N_16884,N_16142);
nor U17179 (N_17179,N_16096,N_16689);
nand U17180 (N_17180,N_16635,N_16618);
nor U17181 (N_17181,N_16845,N_16630);
nor U17182 (N_17182,N_16237,N_16260);
nor U17183 (N_17183,N_16622,N_16421);
nand U17184 (N_17184,N_16413,N_16534);
nor U17185 (N_17185,N_16775,N_16295);
nor U17186 (N_17186,N_16537,N_16351);
nand U17187 (N_17187,N_16332,N_16723);
nand U17188 (N_17188,N_16178,N_16785);
or U17189 (N_17189,N_16699,N_16035);
and U17190 (N_17190,N_16742,N_16900);
nor U17191 (N_17191,N_16602,N_16520);
or U17192 (N_17192,N_16514,N_16111);
nor U17193 (N_17193,N_16550,N_16185);
or U17194 (N_17194,N_16199,N_16409);
or U17195 (N_17195,N_16339,N_16434);
and U17196 (N_17196,N_16999,N_16947);
xor U17197 (N_17197,N_16682,N_16856);
xor U17198 (N_17198,N_16474,N_16934);
nor U17199 (N_17199,N_16746,N_16949);
and U17200 (N_17200,N_16047,N_16790);
nand U17201 (N_17201,N_16817,N_16350);
nor U17202 (N_17202,N_16506,N_16232);
xnor U17203 (N_17203,N_16889,N_16328);
or U17204 (N_17204,N_16006,N_16033);
or U17205 (N_17205,N_16749,N_16919);
nor U17206 (N_17206,N_16801,N_16991);
nor U17207 (N_17207,N_16151,N_16196);
nand U17208 (N_17208,N_16759,N_16352);
nand U17209 (N_17209,N_16551,N_16776);
nor U17210 (N_17210,N_16929,N_16179);
or U17211 (N_17211,N_16347,N_16308);
and U17212 (N_17212,N_16303,N_16741);
nand U17213 (N_17213,N_16565,N_16779);
or U17214 (N_17214,N_16781,N_16277);
xnor U17215 (N_17215,N_16574,N_16625);
or U17216 (N_17216,N_16960,N_16524);
or U17217 (N_17217,N_16758,N_16750);
or U17218 (N_17218,N_16346,N_16661);
or U17219 (N_17219,N_16478,N_16270);
or U17220 (N_17220,N_16202,N_16886);
nand U17221 (N_17221,N_16529,N_16464);
nor U17222 (N_17222,N_16219,N_16387);
xor U17223 (N_17223,N_16896,N_16080);
or U17224 (N_17224,N_16136,N_16105);
and U17225 (N_17225,N_16454,N_16792);
xor U17226 (N_17226,N_16744,N_16745);
or U17227 (N_17227,N_16730,N_16390);
and U17228 (N_17228,N_16397,N_16944);
xor U17229 (N_17229,N_16722,N_16611);
and U17230 (N_17230,N_16127,N_16724);
nand U17231 (N_17231,N_16617,N_16853);
or U17232 (N_17232,N_16269,N_16194);
xor U17233 (N_17233,N_16981,N_16287);
nor U17234 (N_17234,N_16753,N_16797);
nand U17235 (N_17235,N_16314,N_16972);
or U17236 (N_17236,N_16412,N_16894);
and U17237 (N_17237,N_16081,N_16445);
xnor U17238 (N_17238,N_16596,N_16399);
nand U17239 (N_17239,N_16294,N_16245);
xnor U17240 (N_17240,N_16358,N_16243);
nand U17241 (N_17241,N_16692,N_16710);
xnor U17242 (N_17242,N_16978,N_16415);
nand U17243 (N_17243,N_16019,N_16285);
or U17244 (N_17244,N_16420,N_16638);
and U17245 (N_17245,N_16507,N_16837);
and U17246 (N_17246,N_16141,N_16490);
nand U17247 (N_17247,N_16027,N_16864);
nor U17248 (N_17248,N_16074,N_16324);
nand U17249 (N_17249,N_16440,N_16271);
xor U17250 (N_17250,N_16469,N_16766);
nor U17251 (N_17251,N_16673,N_16795);
nand U17252 (N_17252,N_16813,N_16226);
nor U17253 (N_17253,N_16847,N_16051);
and U17254 (N_17254,N_16966,N_16866);
nand U17255 (N_17255,N_16265,N_16238);
and U17256 (N_17256,N_16015,N_16175);
nand U17257 (N_17257,N_16654,N_16497);
xor U17258 (N_17258,N_16561,N_16769);
and U17259 (N_17259,N_16402,N_16822);
and U17260 (N_17260,N_16070,N_16824);
nor U17261 (N_17261,N_16688,N_16748);
and U17262 (N_17262,N_16647,N_16553);
or U17263 (N_17263,N_16765,N_16984);
or U17264 (N_17264,N_16995,N_16842);
nor U17265 (N_17265,N_16498,N_16755);
or U17266 (N_17266,N_16633,N_16133);
xor U17267 (N_17267,N_16706,N_16875);
xor U17268 (N_17268,N_16880,N_16740);
and U17269 (N_17269,N_16119,N_16562);
or U17270 (N_17270,N_16976,N_16137);
or U17271 (N_17271,N_16802,N_16013);
nor U17272 (N_17272,N_16882,N_16160);
nor U17273 (N_17273,N_16299,N_16811);
nand U17274 (N_17274,N_16820,N_16629);
or U17275 (N_17275,N_16248,N_16034);
and U17276 (N_17276,N_16861,N_16457);
or U17277 (N_17277,N_16140,N_16604);
xor U17278 (N_17278,N_16483,N_16970);
nand U17279 (N_17279,N_16998,N_16128);
and U17280 (N_17280,N_16223,N_16067);
nand U17281 (N_17281,N_16021,N_16200);
nand U17282 (N_17282,N_16705,N_16834);
nand U17283 (N_17283,N_16502,N_16544);
or U17284 (N_17284,N_16465,N_16201);
nor U17285 (N_17285,N_16163,N_16615);
nand U17286 (N_17286,N_16256,N_16131);
or U17287 (N_17287,N_16676,N_16325);
xor U17288 (N_17288,N_16213,N_16297);
or U17289 (N_17289,N_16573,N_16757);
and U17290 (N_17290,N_16362,N_16904);
and U17291 (N_17291,N_16250,N_16547);
xor U17292 (N_17292,N_16585,N_16980);
or U17293 (N_17293,N_16101,N_16933);
nand U17294 (N_17294,N_16121,N_16503);
and U17295 (N_17295,N_16814,N_16850);
xnor U17296 (N_17296,N_16895,N_16906);
nand U17297 (N_17297,N_16613,N_16572);
or U17298 (N_17298,N_16902,N_16952);
nand U17299 (N_17299,N_16180,N_16113);
or U17300 (N_17300,N_16037,N_16242);
nor U17301 (N_17301,N_16721,N_16403);
and U17302 (N_17302,N_16426,N_16298);
and U17303 (N_17303,N_16872,N_16025);
and U17304 (N_17304,N_16485,N_16566);
and U17305 (N_17305,N_16214,N_16307);
xor U17306 (N_17306,N_16162,N_16064);
nor U17307 (N_17307,N_16416,N_16586);
nand U17308 (N_17308,N_16153,N_16533);
and U17309 (N_17309,N_16334,N_16363);
and U17310 (N_17310,N_16593,N_16783);
and U17311 (N_17311,N_16846,N_16729);
nor U17312 (N_17312,N_16932,N_16309);
and U17313 (N_17313,N_16969,N_16044);
nand U17314 (N_17314,N_16407,N_16049);
xor U17315 (N_17315,N_16918,N_16401);
and U17316 (N_17316,N_16110,N_16907);
nor U17317 (N_17317,N_16311,N_16367);
nand U17318 (N_17318,N_16395,N_16558);
xor U17319 (N_17319,N_16716,N_16825);
nor U17320 (N_17320,N_16312,N_16317);
xnor U17321 (N_17321,N_16234,N_16974);
xor U17322 (N_17322,N_16282,N_16188);
nor U17323 (N_17323,N_16940,N_16948);
or U17324 (N_17324,N_16496,N_16236);
and U17325 (N_17325,N_16908,N_16860);
xor U17326 (N_17326,N_16809,N_16276);
xor U17327 (N_17327,N_16345,N_16560);
and U17328 (N_17328,N_16526,N_16874);
nor U17329 (N_17329,N_16418,N_16982);
and U17330 (N_17330,N_16233,N_16512);
nor U17331 (N_17331,N_16612,N_16481);
nand U17332 (N_17332,N_16782,N_16134);
and U17333 (N_17333,N_16580,N_16805);
xnor U17334 (N_17334,N_16290,N_16930);
and U17335 (N_17335,N_16711,N_16658);
or U17336 (N_17336,N_16447,N_16690);
nand U17337 (N_17337,N_16651,N_16357);
xor U17338 (N_17338,N_16587,N_16181);
and U17339 (N_17339,N_16122,N_16370);
xnor U17340 (N_17340,N_16905,N_16495);
or U17341 (N_17341,N_16720,N_16786);
xnor U17342 (N_17342,N_16031,N_16471);
and U17343 (N_17343,N_16432,N_16857);
nand U17344 (N_17344,N_16885,N_16598);
nand U17345 (N_17345,N_16511,N_16349);
and U17346 (N_17346,N_16104,N_16165);
nor U17347 (N_17347,N_16754,N_16493);
or U17348 (N_17348,N_16943,N_16123);
nor U17349 (N_17349,N_16848,N_16417);
xnor U17350 (N_17350,N_16264,N_16210);
and U17351 (N_17351,N_16925,N_16996);
xnor U17352 (N_17352,N_16173,N_16461);
nand U17353 (N_17353,N_16575,N_16207);
or U17354 (N_17354,N_16280,N_16725);
nor U17355 (N_17355,N_16616,N_16732);
xor U17356 (N_17356,N_16518,N_16610);
and U17357 (N_17357,N_16712,N_16404);
nand U17358 (N_17358,N_16667,N_16773);
and U17359 (N_17359,N_16595,N_16657);
and U17360 (N_17360,N_16897,N_16628);
nand U17361 (N_17361,N_16071,N_16069);
nor U17362 (N_17362,N_16344,N_16423);
and U17363 (N_17363,N_16315,N_16190);
and U17364 (N_17364,N_16306,N_16697);
or U17365 (N_17365,N_16052,N_16437);
nor U17366 (N_17366,N_16731,N_16545);
or U17367 (N_17367,N_16386,N_16220);
and U17368 (N_17368,N_16355,N_16391);
nand U17369 (N_17369,N_16686,N_16938);
nor U17370 (N_17370,N_16958,N_16275);
nor U17371 (N_17371,N_16383,N_16590);
xnor U17372 (N_17372,N_16443,N_16793);
and U17373 (N_17373,N_16956,N_16571);
nor U17374 (N_17374,N_16570,N_16283);
and U17375 (N_17375,N_16491,N_16186);
and U17376 (N_17376,N_16336,N_16871);
or U17377 (N_17377,N_16563,N_16876);
and U17378 (N_17378,N_16916,N_16005);
nor U17379 (N_17379,N_16103,N_16112);
or U17380 (N_17380,N_16883,N_16441);
nand U17381 (N_17381,N_16427,N_16756);
nor U17382 (N_17382,N_16281,N_16184);
nand U17383 (N_17383,N_16737,N_16092);
or U17384 (N_17384,N_16170,N_16770);
nor U17385 (N_17385,N_16582,N_16120);
xor U17386 (N_17386,N_16348,N_16987);
or U17387 (N_17387,N_16523,N_16607);
and U17388 (N_17388,N_16230,N_16921);
xor U17389 (N_17389,N_16487,N_16936);
nor U17390 (N_17390,N_16254,N_16378);
and U17391 (N_17391,N_16796,N_16522);
nand U17392 (N_17392,N_16835,N_16078);
nor U17393 (N_17393,N_16519,N_16149);
nor U17394 (N_17394,N_16804,N_16868);
nor U17395 (N_17395,N_16318,N_16843);
nand U17396 (N_17396,N_16100,N_16359);
or U17397 (N_17397,N_16878,N_16396);
nor U17398 (N_17398,N_16011,N_16893);
nor U17399 (N_17399,N_16192,N_16155);
nand U17400 (N_17400,N_16003,N_16266);
and U17401 (N_17401,N_16659,N_16056);
xor U17402 (N_17402,N_16024,N_16993);
or U17403 (N_17403,N_16102,N_16662);
and U17404 (N_17404,N_16466,N_16994);
and U17405 (N_17405,N_16791,N_16767);
nor U17406 (N_17406,N_16803,N_16578);
nor U17407 (N_17407,N_16927,N_16384);
and U17408 (N_17408,N_16603,N_16494);
and U17409 (N_17409,N_16425,N_16733);
nor U17410 (N_17410,N_16124,N_16823);
nor U17411 (N_17411,N_16589,N_16302);
xor U17412 (N_17412,N_16147,N_16844);
xnor U17413 (N_17413,N_16542,N_16903);
nor U17414 (N_17414,N_16784,N_16198);
xnor U17415 (N_17415,N_16342,N_16499);
nand U17416 (N_17416,N_16492,N_16012);
nand U17417 (N_17417,N_16235,N_16713);
nand U17418 (N_17418,N_16477,N_16915);
xor U17419 (N_17419,N_16087,N_16540);
or U17420 (N_17420,N_16609,N_16026);
nand U17421 (N_17421,N_16592,N_16877);
xor U17422 (N_17422,N_16760,N_16743);
nand U17423 (N_17423,N_16715,N_16680);
nor U17424 (N_17424,N_16836,N_16890);
nor U17425 (N_17425,N_16858,N_16419);
nor U17426 (N_17426,N_16675,N_16337);
xor U17427 (N_17427,N_16433,N_16899);
xor U17428 (N_17428,N_16125,N_16539);
nand U17429 (N_17429,N_16118,N_16353);
xor U17430 (N_17430,N_16039,N_16076);
nor U17431 (N_17431,N_16183,N_16666);
nand U17432 (N_17432,N_16455,N_16807);
or U17433 (N_17433,N_16244,N_16879);
nor U17434 (N_17434,N_16597,N_16273);
or U17435 (N_17435,N_16392,N_16695);
and U17436 (N_17436,N_16148,N_16168);
and U17437 (N_17437,N_16055,N_16986);
nor U17438 (N_17438,N_16913,N_16701);
xnor U17439 (N_17439,N_16073,N_16215);
and U17440 (N_17440,N_16489,N_16193);
nor U17441 (N_17441,N_16694,N_16108);
and U17442 (N_17442,N_16687,N_16187);
and U17443 (N_17443,N_16405,N_16221);
nor U17444 (N_17444,N_16973,N_16107);
or U17445 (N_17445,N_16569,N_16504);
or U17446 (N_17446,N_16702,N_16278);
xor U17447 (N_17447,N_16935,N_16567);
or U17448 (N_17448,N_16305,N_16376);
nor U17449 (N_17449,N_16288,N_16004);
and U17450 (N_17450,N_16229,N_16968);
and U17451 (N_17451,N_16059,N_16368);
and U17452 (N_17452,N_16869,N_16950);
or U17453 (N_17453,N_16476,N_16830);
nor U17454 (N_17454,N_16821,N_16644);
nand U17455 (N_17455,N_16579,N_16338);
or U17456 (N_17456,N_16988,N_16115);
nor U17457 (N_17457,N_16169,N_16832);
nand U17458 (N_17458,N_16521,N_16463);
xnor U17459 (N_17459,N_16764,N_16331);
xnor U17460 (N_17460,N_16663,N_16255);
nand U17461 (N_17461,N_16911,N_16849);
nor U17462 (N_17462,N_16961,N_16865);
and U17463 (N_17463,N_16098,N_16516);
and U17464 (N_17464,N_16772,N_16095);
or U17465 (N_17465,N_16787,N_16989);
and U17466 (N_17466,N_16525,N_16505);
xnor U17467 (N_17467,N_16203,N_16583);
and U17468 (N_17468,N_16668,N_16083);
or U17469 (N_17469,N_16436,N_16671);
nand U17470 (N_17470,N_16829,N_16962);
and U17471 (N_17471,N_16909,N_16703);
xor U17472 (N_17472,N_16300,N_16975);
nor U17473 (N_17473,N_16172,N_16508);
xor U17474 (N_17474,N_16145,N_16097);
and U17475 (N_17475,N_16486,N_16738);
and U17476 (N_17476,N_16138,N_16045);
or U17477 (N_17477,N_16381,N_16543);
or U17478 (N_17478,N_16774,N_16114);
xor U17479 (N_17479,N_16910,N_16632);
nand U17480 (N_17480,N_16636,N_16177);
nor U17481 (N_17481,N_16640,N_16964);
or U17482 (N_17482,N_16456,N_16528);
or U17483 (N_17483,N_16430,N_16679);
nand U17484 (N_17484,N_16735,N_16818);
and U17485 (N_17485,N_16206,N_16020);
nor U17486 (N_17486,N_16867,N_16833);
xnor U17487 (N_17487,N_16794,N_16608);
nand U17488 (N_17488,N_16531,N_16736);
and U17489 (N_17489,N_16227,N_16967);
and U17490 (N_17490,N_16831,N_16380);
and U17491 (N_17491,N_16191,N_16088);
nand U17492 (N_17492,N_16530,N_16130);
nand U17493 (N_17493,N_16728,N_16340);
nor U17494 (N_17494,N_16923,N_16253);
xor U17495 (N_17495,N_16329,N_16132);
and U17496 (N_17496,N_16444,N_16360);
or U17497 (N_17497,N_16241,N_16693);
nand U17498 (N_17498,N_16719,N_16061);
xor U17499 (N_17499,N_16652,N_16855);
nand U17500 (N_17500,N_16783,N_16110);
or U17501 (N_17501,N_16013,N_16619);
nor U17502 (N_17502,N_16112,N_16966);
nor U17503 (N_17503,N_16879,N_16670);
and U17504 (N_17504,N_16064,N_16277);
and U17505 (N_17505,N_16655,N_16586);
or U17506 (N_17506,N_16614,N_16905);
or U17507 (N_17507,N_16322,N_16315);
or U17508 (N_17508,N_16666,N_16320);
xnor U17509 (N_17509,N_16786,N_16742);
and U17510 (N_17510,N_16073,N_16800);
nand U17511 (N_17511,N_16275,N_16867);
nor U17512 (N_17512,N_16512,N_16781);
and U17513 (N_17513,N_16390,N_16844);
nor U17514 (N_17514,N_16364,N_16153);
nand U17515 (N_17515,N_16692,N_16866);
xnor U17516 (N_17516,N_16330,N_16894);
xor U17517 (N_17517,N_16659,N_16909);
nand U17518 (N_17518,N_16802,N_16490);
and U17519 (N_17519,N_16054,N_16642);
xor U17520 (N_17520,N_16467,N_16515);
nand U17521 (N_17521,N_16197,N_16697);
and U17522 (N_17522,N_16785,N_16356);
and U17523 (N_17523,N_16671,N_16863);
nor U17524 (N_17524,N_16219,N_16582);
xor U17525 (N_17525,N_16325,N_16760);
nand U17526 (N_17526,N_16968,N_16568);
xor U17527 (N_17527,N_16802,N_16993);
xor U17528 (N_17528,N_16547,N_16195);
and U17529 (N_17529,N_16047,N_16694);
nand U17530 (N_17530,N_16882,N_16255);
and U17531 (N_17531,N_16127,N_16384);
nor U17532 (N_17532,N_16548,N_16291);
and U17533 (N_17533,N_16577,N_16209);
or U17534 (N_17534,N_16449,N_16012);
or U17535 (N_17535,N_16843,N_16314);
nand U17536 (N_17536,N_16630,N_16763);
xor U17537 (N_17537,N_16480,N_16255);
and U17538 (N_17538,N_16389,N_16341);
xnor U17539 (N_17539,N_16487,N_16907);
nand U17540 (N_17540,N_16031,N_16066);
and U17541 (N_17541,N_16605,N_16483);
nand U17542 (N_17542,N_16776,N_16988);
nor U17543 (N_17543,N_16379,N_16645);
or U17544 (N_17544,N_16474,N_16952);
and U17545 (N_17545,N_16080,N_16842);
nor U17546 (N_17546,N_16987,N_16799);
nor U17547 (N_17547,N_16329,N_16987);
and U17548 (N_17548,N_16203,N_16844);
and U17549 (N_17549,N_16155,N_16345);
xnor U17550 (N_17550,N_16839,N_16108);
nor U17551 (N_17551,N_16437,N_16383);
nand U17552 (N_17552,N_16920,N_16865);
nand U17553 (N_17553,N_16508,N_16930);
xor U17554 (N_17554,N_16917,N_16389);
xor U17555 (N_17555,N_16437,N_16464);
nor U17556 (N_17556,N_16353,N_16373);
xnor U17557 (N_17557,N_16137,N_16839);
xnor U17558 (N_17558,N_16260,N_16835);
and U17559 (N_17559,N_16648,N_16472);
xor U17560 (N_17560,N_16095,N_16031);
xnor U17561 (N_17561,N_16337,N_16039);
nor U17562 (N_17562,N_16959,N_16784);
nor U17563 (N_17563,N_16235,N_16041);
nor U17564 (N_17564,N_16372,N_16141);
and U17565 (N_17565,N_16914,N_16397);
and U17566 (N_17566,N_16310,N_16966);
nand U17567 (N_17567,N_16565,N_16694);
and U17568 (N_17568,N_16284,N_16599);
xor U17569 (N_17569,N_16613,N_16547);
and U17570 (N_17570,N_16080,N_16326);
and U17571 (N_17571,N_16645,N_16462);
or U17572 (N_17572,N_16455,N_16626);
or U17573 (N_17573,N_16502,N_16576);
xnor U17574 (N_17574,N_16487,N_16370);
nor U17575 (N_17575,N_16109,N_16796);
nor U17576 (N_17576,N_16354,N_16307);
xnor U17577 (N_17577,N_16728,N_16905);
and U17578 (N_17578,N_16819,N_16749);
xor U17579 (N_17579,N_16411,N_16899);
or U17580 (N_17580,N_16303,N_16699);
or U17581 (N_17581,N_16934,N_16286);
and U17582 (N_17582,N_16830,N_16661);
and U17583 (N_17583,N_16563,N_16236);
xnor U17584 (N_17584,N_16028,N_16648);
nand U17585 (N_17585,N_16709,N_16583);
nor U17586 (N_17586,N_16612,N_16696);
xor U17587 (N_17587,N_16171,N_16416);
nor U17588 (N_17588,N_16671,N_16891);
xnor U17589 (N_17589,N_16273,N_16080);
or U17590 (N_17590,N_16102,N_16254);
nor U17591 (N_17591,N_16334,N_16810);
xor U17592 (N_17592,N_16937,N_16768);
nand U17593 (N_17593,N_16556,N_16922);
nor U17594 (N_17594,N_16174,N_16096);
and U17595 (N_17595,N_16426,N_16286);
xor U17596 (N_17596,N_16729,N_16581);
or U17597 (N_17597,N_16419,N_16513);
and U17598 (N_17598,N_16578,N_16758);
nor U17599 (N_17599,N_16057,N_16863);
and U17600 (N_17600,N_16817,N_16558);
or U17601 (N_17601,N_16181,N_16160);
and U17602 (N_17602,N_16877,N_16324);
or U17603 (N_17603,N_16577,N_16222);
or U17604 (N_17604,N_16028,N_16143);
xnor U17605 (N_17605,N_16908,N_16850);
xnor U17606 (N_17606,N_16870,N_16158);
and U17607 (N_17607,N_16492,N_16165);
nor U17608 (N_17608,N_16845,N_16607);
and U17609 (N_17609,N_16863,N_16917);
nor U17610 (N_17610,N_16973,N_16095);
nor U17611 (N_17611,N_16514,N_16418);
xor U17612 (N_17612,N_16160,N_16067);
xnor U17613 (N_17613,N_16476,N_16168);
nand U17614 (N_17614,N_16888,N_16746);
or U17615 (N_17615,N_16791,N_16551);
nand U17616 (N_17616,N_16453,N_16791);
or U17617 (N_17617,N_16170,N_16277);
nor U17618 (N_17618,N_16930,N_16749);
nor U17619 (N_17619,N_16079,N_16019);
or U17620 (N_17620,N_16805,N_16128);
xor U17621 (N_17621,N_16992,N_16074);
xnor U17622 (N_17622,N_16472,N_16281);
xor U17623 (N_17623,N_16990,N_16790);
and U17624 (N_17624,N_16572,N_16004);
or U17625 (N_17625,N_16398,N_16518);
nand U17626 (N_17626,N_16762,N_16979);
nor U17627 (N_17627,N_16988,N_16342);
nor U17628 (N_17628,N_16164,N_16041);
or U17629 (N_17629,N_16142,N_16967);
nand U17630 (N_17630,N_16180,N_16439);
nor U17631 (N_17631,N_16446,N_16333);
xor U17632 (N_17632,N_16404,N_16481);
xnor U17633 (N_17633,N_16058,N_16128);
and U17634 (N_17634,N_16216,N_16119);
or U17635 (N_17635,N_16751,N_16445);
nand U17636 (N_17636,N_16095,N_16442);
nand U17637 (N_17637,N_16844,N_16890);
nor U17638 (N_17638,N_16623,N_16079);
nor U17639 (N_17639,N_16700,N_16998);
or U17640 (N_17640,N_16721,N_16887);
nand U17641 (N_17641,N_16010,N_16257);
and U17642 (N_17642,N_16115,N_16724);
xor U17643 (N_17643,N_16574,N_16806);
xnor U17644 (N_17644,N_16708,N_16456);
nor U17645 (N_17645,N_16149,N_16721);
nand U17646 (N_17646,N_16458,N_16549);
nand U17647 (N_17647,N_16343,N_16963);
nand U17648 (N_17648,N_16570,N_16937);
and U17649 (N_17649,N_16255,N_16403);
and U17650 (N_17650,N_16362,N_16844);
nand U17651 (N_17651,N_16600,N_16405);
xor U17652 (N_17652,N_16354,N_16102);
nor U17653 (N_17653,N_16402,N_16571);
and U17654 (N_17654,N_16683,N_16228);
or U17655 (N_17655,N_16928,N_16397);
and U17656 (N_17656,N_16502,N_16265);
and U17657 (N_17657,N_16989,N_16346);
nor U17658 (N_17658,N_16158,N_16422);
xnor U17659 (N_17659,N_16065,N_16570);
xor U17660 (N_17660,N_16545,N_16499);
xnor U17661 (N_17661,N_16717,N_16381);
xor U17662 (N_17662,N_16458,N_16042);
xor U17663 (N_17663,N_16537,N_16295);
xnor U17664 (N_17664,N_16040,N_16321);
or U17665 (N_17665,N_16221,N_16257);
or U17666 (N_17666,N_16390,N_16077);
and U17667 (N_17667,N_16047,N_16783);
xor U17668 (N_17668,N_16977,N_16742);
nand U17669 (N_17669,N_16967,N_16218);
or U17670 (N_17670,N_16101,N_16216);
and U17671 (N_17671,N_16135,N_16838);
xor U17672 (N_17672,N_16426,N_16383);
xor U17673 (N_17673,N_16081,N_16104);
or U17674 (N_17674,N_16935,N_16548);
or U17675 (N_17675,N_16827,N_16818);
and U17676 (N_17676,N_16426,N_16902);
xnor U17677 (N_17677,N_16740,N_16843);
and U17678 (N_17678,N_16750,N_16367);
and U17679 (N_17679,N_16857,N_16169);
and U17680 (N_17680,N_16198,N_16907);
or U17681 (N_17681,N_16868,N_16001);
or U17682 (N_17682,N_16216,N_16292);
nand U17683 (N_17683,N_16056,N_16751);
or U17684 (N_17684,N_16511,N_16514);
or U17685 (N_17685,N_16702,N_16811);
nand U17686 (N_17686,N_16743,N_16402);
or U17687 (N_17687,N_16894,N_16987);
or U17688 (N_17688,N_16823,N_16198);
xnor U17689 (N_17689,N_16307,N_16543);
xor U17690 (N_17690,N_16323,N_16163);
or U17691 (N_17691,N_16664,N_16701);
nand U17692 (N_17692,N_16739,N_16861);
xnor U17693 (N_17693,N_16987,N_16147);
xor U17694 (N_17694,N_16967,N_16028);
nor U17695 (N_17695,N_16298,N_16537);
or U17696 (N_17696,N_16687,N_16820);
xnor U17697 (N_17697,N_16816,N_16600);
and U17698 (N_17698,N_16628,N_16408);
nor U17699 (N_17699,N_16228,N_16830);
and U17700 (N_17700,N_16396,N_16823);
and U17701 (N_17701,N_16734,N_16426);
nand U17702 (N_17702,N_16426,N_16805);
and U17703 (N_17703,N_16188,N_16924);
nand U17704 (N_17704,N_16860,N_16686);
and U17705 (N_17705,N_16817,N_16621);
nand U17706 (N_17706,N_16930,N_16138);
and U17707 (N_17707,N_16055,N_16692);
and U17708 (N_17708,N_16443,N_16365);
and U17709 (N_17709,N_16512,N_16732);
or U17710 (N_17710,N_16039,N_16327);
xor U17711 (N_17711,N_16803,N_16498);
xor U17712 (N_17712,N_16867,N_16777);
and U17713 (N_17713,N_16201,N_16367);
nand U17714 (N_17714,N_16168,N_16545);
nor U17715 (N_17715,N_16154,N_16299);
or U17716 (N_17716,N_16570,N_16453);
xnor U17717 (N_17717,N_16772,N_16123);
or U17718 (N_17718,N_16903,N_16482);
nand U17719 (N_17719,N_16000,N_16749);
nor U17720 (N_17720,N_16217,N_16651);
nor U17721 (N_17721,N_16519,N_16428);
and U17722 (N_17722,N_16958,N_16926);
xor U17723 (N_17723,N_16499,N_16053);
and U17724 (N_17724,N_16454,N_16196);
or U17725 (N_17725,N_16950,N_16674);
and U17726 (N_17726,N_16866,N_16474);
and U17727 (N_17727,N_16828,N_16597);
or U17728 (N_17728,N_16485,N_16028);
nand U17729 (N_17729,N_16132,N_16793);
nand U17730 (N_17730,N_16689,N_16238);
or U17731 (N_17731,N_16387,N_16040);
xor U17732 (N_17732,N_16995,N_16811);
xor U17733 (N_17733,N_16253,N_16829);
or U17734 (N_17734,N_16256,N_16648);
or U17735 (N_17735,N_16116,N_16633);
nand U17736 (N_17736,N_16143,N_16565);
xnor U17737 (N_17737,N_16432,N_16201);
nand U17738 (N_17738,N_16108,N_16207);
xnor U17739 (N_17739,N_16866,N_16445);
or U17740 (N_17740,N_16121,N_16323);
or U17741 (N_17741,N_16958,N_16293);
and U17742 (N_17742,N_16124,N_16024);
nor U17743 (N_17743,N_16721,N_16802);
and U17744 (N_17744,N_16916,N_16784);
nand U17745 (N_17745,N_16285,N_16834);
nand U17746 (N_17746,N_16492,N_16323);
or U17747 (N_17747,N_16192,N_16291);
xnor U17748 (N_17748,N_16409,N_16628);
and U17749 (N_17749,N_16353,N_16455);
xnor U17750 (N_17750,N_16838,N_16916);
xor U17751 (N_17751,N_16008,N_16897);
nand U17752 (N_17752,N_16277,N_16425);
nand U17753 (N_17753,N_16982,N_16532);
nand U17754 (N_17754,N_16220,N_16289);
and U17755 (N_17755,N_16634,N_16724);
or U17756 (N_17756,N_16049,N_16677);
and U17757 (N_17757,N_16285,N_16903);
nor U17758 (N_17758,N_16237,N_16315);
or U17759 (N_17759,N_16827,N_16964);
nor U17760 (N_17760,N_16697,N_16635);
xnor U17761 (N_17761,N_16979,N_16517);
or U17762 (N_17762,N_16052,N_16192);
nor U17763 (N_17763,N_16100,N_16881);
xnor U17764 (N_17764,N_16343,N_16159);
nand U17765 (N_17765,N_16541,N_16224);
nor U17766 (N_17766,N_16612,N_16757);
nor U17767 (N_17767,N_16464,N_16159);
and U17768 (N_17768,N_16375,N_16875);
nand U17769 (N_17769,N_16996,N_16126);
or U17770 (N_17770,N_16552,N_16472);
xnor U17771 (N_17771,N_16696,N_16317);
nor U17772 (N_17772,N_16708,N_16256);
nand U17773 (N_17773,N_16283,N_16689);
or U17774 (N_17774,N_16818,N_16502);
nand U17775 (N_17775,N_16130,N_16687);
nand U17776 (N_17776,N_16567,N_16912);
xor U17777 (N_17777,N_16249,N_16996);
or U17778 (N_17778,N_16833,N_16386);
and U17779 (N_17779,N_16809,N_16844);
nand U17780 (N_17780,N_16977,N_16844);
nand U17781 (N_17781,N_16726,N_16580);
and U17782 (N_17782,N_16694,N_16135);
nand U17783 (N_17783,N_16151,N_16846);
or U17784 (N_17784,N_16896,N_16672);
or U17785 (N_17785,N_16116,N_16544);
xnor U17786 (N_17786,N_16803,N_16374);
nor U17787 (N_17787,N_16782,N_16768);
and U17788 (N_17788,N_16144,N_16487);
and U17789 (N_17789,N_16054,N_16479);
or U17790 (N_17790,N_16934,N_16418);
and U17791 (N_17791,N_16296,N_16960);
nor U17792 (N_17792,N_16702,N_16382);
xor U17793 (N_17793,N_16460,N_16667);
xnor U17794 (N_17794,N_16981,N_16688);
nand U17795 (N_17795,N_16423,N_16774);
nand U17796 (N_17796,N_16905,N_16523);
or U17797 (N_17797,N_16182,N_16764);
nor U17798 (N_17798,N_16513,N_16298);
nand U17799 (N_17799,N_16058,N_16268);
xnor U17800 (N_17800,N_16929,N_16056);
nor U17801 (N_17801,N_16907,N_16289);
nor U17802 (N_17802,N_16956,N_16087);
nand U17803 (N_17803,N_16221,N_16781);
nand U17804 (N_17804,N_16596,N_16710);
or U17805 (N_17805,N_16770,N_16733);
or U17806 (N_17806,N_16333,N_16674);
xnor U17807 (N_17807,N_16825,N_16181);
or U17808 (N_17808,N_16053,N_16062);
and U17809 (N_17809,N_16085,N_16011);
nand U17810 (N_17810,N_16035,N_16010);
xor U17811 (N_17811,N_16465,N_16008);
xor U17812 (N_17812,N_16968,N_16700);
and U17813 (N_17813,N_16599,N_16061);
xnor U17814 (N_17814,N_16749,N_16110);
xnor U17815 (N_17815,N_16359,N_16364);
nand U17816 (N_17816,N_16253,N_16432);
xor U17817 (N_17817,N_16389,N_16911);
or U17818 (N_17818,N_16443,N_16691);
or U17819 (N_17819,N_16036,N_16961);
or U17820 (N_17820,N_16730,N_16200);
nor U17821 (N_17821,N_16283,N_16640);
and U17822 (N_17822,N_16035,N_16599);
or U17823 (N_17823,N_16225,N_16015);
or U17824 (N_17824,N_16919,N_16628);
nor U17825 (N_17825,N_16659,N_16161);
nor U17826 (N_17826,N_16275,N_16451);
xnor U17827 (N_17827,N_16033,N_16212);
nor U17828 (N_17828,N_16628,N_16187);
nor U17829 (N_17829,N_16109,N_16947);
xor U17830 (N_17830,N_16245,N_16192);
xor U17831 (N_17831,N_16372,N_16146);
and U17832 (N_17832,N_16463,N_16249);
and U17833 (N_17833,N_16536,N_16983);
and U17834 (N_17834,N_16559,N_16490);
xnor U17835 (N_17835,N_16546,N_16174);
xnor U17836 (N_17836,N_16230,N_16183);
and U17837 (N_17837,N_16687,N_16626);
and U17838 (N_17838,N_16820,N_16597);
and U17839 (N_17839,N_16441,N_16972);
and U17840 (N_17840,N_16124,N_16522);
xnor U17841 (N_17841,N_16237,N_16328);
nor U17842 (N_17842,N_16432,N_16262);
and U17843 (N_17843,N_16704,N_16641);
or U17844 (N_17844,N_16687,N_16399);
or U17845 (N_17845,N_16925,N_16802);
nor U17846 (N_17846,N_16247,N_16202);
xor U17847 (N_17847,N_16830,N_16613);
xnor U17848 (N_17848,N_16205,N_16734);
or U17849 (N_17849,N_16136,N_16445);
and U17850 (N_17850,N_16496,N_16254);
and U17851 (N_17851,N_16491,N_16298);
or U17852 (N_17852,N_16615,N_16027);
or U17853 (N_17853,N_16079,N_16603);
and U17854 (N_17854,N_16711,N_16030);
and U17855 (N_17855,N_16813,N_16926);
xnor U17856 (N_17856,N_16967,N_16514);
xor U17857 (N_17857,N_16649,N_16734);
xor U17858 (N_17858,N_16770,N_16102);
or U17859 (N_17859,N_16607,N_16992);
and U17860 (N_17860,N_16422,N_16329);
and U17861 (N_17861,N_16665,N_16831);
and U17862 (N_17862,N_16200,N_16880);
or U17863 (N_17863,N_16106,N_16631);
or U17864 (N_17864,N_16039,N_16630);
nand U17865 (N_17865,N_16197,N_16747);
or U17866 (N_17866,N_16897,N_16410);
xnor U17867 (N_17867,N_16546,N_16618);
and U17868 (N_17868,N_16373,N_16031);
nand U17869 (N_17869,N_16173,N_16650);
nor U17870 (N_17870,N_16306,N_16884);
and U17871 (N_17871,N_16889,N_16419);
or U17872 (N_17872,N_16525,N_16721);
and U17873 (N_17873,N_16594,N_16340);
nor U17874 (N_17874,N_16263,N_16167);
nor U17875 (N_17875,N_16897,N_16668);
or U17876 (N_17876,N_16661,N_16524);
xor U17877 (N_17877,N_16655,N_16325);
and U17878 (N_17878,N_16170,N_16983);
or U17879 (N_17879,N_16112,N_16879);
xor U17880 (N_17880,N_16121,N_16788);
and U17881 (N_17881,N_16883,N_16642);
or U17882 (N_17882,N_16687,N_16676);
and U17883 (N_17883,N_16008,N_16812);
nand U17884 (N_17884,N_16096,N_16962);
nand U17885 (N_17885,N_16797,N_16177);
and U17886 (N_17886,N_16624,N_16665);
xnor U17887 (N_17887,N_16733,N_16611);
nor U17888 (N_17888,N_16465,N_16326);
nor U17889 (N_17889,N_16233,N_16471);
nand U17890 (N_17890,N_16435,N_16507);
or U17891 (N_17891,N_16562,N_16325);
and U17892 (N_17892,N_16904,N_16522);
nand U17893 (N_17893,N_16184,N_16287);
xor U17894 (N_17894,N_16034,N_16835);
nor U17895 (N_17895,N_16954,N_16253);
nand U17896 (N_17896,N_16523,N_16472);
or U17897 (N_17897,N_16083,N_16296);
nand U17898 (N_17898,N_16492,N_16725);
xnor U17899 (N_17899,N_16591,N_16445);
nor U17900 (N_17900,N_16935,N_16154);
nand U17901 (N_17901,N_16921,N_16055);
xor U17902 (N_17902,N_16849,N_16445);
and U17903 (N_17903,N_16571,N_16135);
and U17904 (N_17904,N_16690,N_16753);
nand U17905 (N_17905,N_16291,N_16202);
nand U17906 (N_17906,N_16362,N_16372);
or U17907 (N_17907,N_16019,N_16099);
and U17908 (N_17908,N_16540,N_16272);
and U17909 (N_17909,N_16770,N_16480);
nor U17910 (N_17910,N_16551,N_16693);
nor U17911 (N_17911,N_16286,N_16837);
and U17912 (N_17912,N_16542,N_16728);
xor U17913 (N_17913,N_16329,N_16279);
and U17914 (N_17914,N_16897,N_16140);
nand U17915 (N_17915,N_16330,N_16885);
xor U17916 (N_17916,N_16735,N_16652);
nand U17917 (N_17917,N_16748,N_16772);
xnor U17918 (N_17918,N_16876,N_16305);
xnor U17919 (N_17919,N_16925,N_16828);
nor U17920 (N_17920,N_16986,N_16919);
xnor U17921 (N_17921,N_16090,N_16429);
and U17922 (N_17922,N_16180,N_16478);
or U17923 (N_17923,N_16064,N_16559);
xor U17924 (N_17924,N_16292,N_16002);
nand U17925 (N_17925,N_16222,N_16099);
or U17926 (N_17926,N_16360,N_16300);
xnor U17927 (N_17927,N_16239,N_16835);
or U17928 (N_17928,N_16313,N_16414);
and U17929 (N_17929,N_16288,N_16131);
nand U17930 (N_17930,N_16823,N_16153);
xnor U17931 (N_17931,N_16680,N_16515);
nor U17932 (N_17932,N_16788,N_16605);
or U17933 (N_17933,N_16824,N_16054);
nor U17934 (N_17934,N_16863,N_16191);
and U17935 (N_17935,N_16026,N_16642);
nor U17936 (N_17936,N_16418,N_16321);
nor U17937 (N_17937,N_16652,N_16509);
xor U17938 (N_17938,N_16870,N_16936);
xnor U17939 (N_17939,N_16681,N_16081);
nor U17940 (N_17940,N_16611,N_16105);
nand U17941 (N_17941,N_16387,N_16462);
and U17942 (N_17942,N_16731,N_16185);
nor U17943 (N_17943,N_16013,N_16417);
nor U17944 (N_17944,N_16321,N_16302);
or U17945 (N_17945,N_16413,N_16196);
and U17946 (N_17946,N_16579,N_16382);
xor U17947 (N_17947,N_16370,N_16088);
or U17948 (N_17948,N_16305,N_16476);
nand U17949 (N_17949,N_16244,N_16301);
nand U17950 (N_17950,N_16394,N_16062);
xor U17951 (N_17951,N_16015,N_16261);
xor U17952 (N_17952,N_16745,N_16792);
and U17953 (N_17953,N_16348,N_16758);
nor U17954 (N_17954,N_16179,N_16103);
or U17955 (N_17955,N_16274,N_16550);
xor U17956 (N_17956,N_16351,N_16453);
xnor U17957 (N_17957,N_16301,N_16489);
and U17958 (N_17958,N_16491,N_16082);
nor U17959 (N_17959,N_16107,N_16282);
xnor U17960 (N_17960,N_16805,N_16953);
or U17961 (N_17961,N_16966,N_16399);
xnor U17962 (N_17962,N_16681,N_16388);
xor U17963 (N_17963,N_16218,N_16409);
xnor U17964 (N_17964,N_16943,N_16496);
nand U17965 (N_17965,N_16805,N_16213);
nand U17966 (N_17966,N_16406,N_16394);
xor U17967 (N_17967,N_16831,N_16821);
nand U17968 (N_17968,N_16936,N_16440);
nor U17969 (N_17969,N_16171,N_16770);
nor U17970 (N_17970,N_16267,N_16910);
nor U17971 (N_17971,N_16026,N_16623);
xor U17972 (N_17972,N_16850,N_16197);
nand U17973 (N_17973,N_16029,N_16139);
nand U17974 (N_17974,N_16384,N_16202);
and U17975 (N_17975,N_16035,N_16327);
xnor U17976 (N_17976,N_16242,N_16135);
nand U17977 (N_17977,N_16680,N_16087);
xor U17978 (N_17978,N_16830,N_16755);
xnor U17979 (N_17979,N_16445,N_16942);
nand U17980 (N_17980,N_16795,N_16825);
xnor U17981 (N_17981,N_16816,N_16193);
nand U17982 (N_17982,N_16876,N_16982);
and U17983 (N_17983,N_16468,N_16841);
nand U17984 (N_17984,N_16414,N_16320);
or U17985 (N_17985,N_16688,N_16943);
nand U17986 (N_17986,N_16642,N_16636);
xnor U17987 (N_17987,N_16975,N_16783);
xnor U17988 (N_17988,N_16094,N_16872);
or U17989 (N_17989,N_16875,N_16431);
xnor U17990 (N_17990,N_16183,N_16315);
and U17991 (N_17991,N_16845,N_16592);
nor U17992 (N_17992,N_16270,N_16785);
xor U17993 (N_17993,N_16828,N_16433);
nand U17994 (N_17994,N_16655,N_16162);
xnor U17995 (N_17995,N_16152,N_16387);
and U17996 (N_17996,N_16449,N_16720);
and U17997 (N_17997,N_16008,N_16066);
or U17998 (N_17998,N_16790,N_16690);
nor U17999 (N_17999,N_16572,N_16429);
nand U18000 (N_18000,N_17448,N_17657);
nand U18001 (N_18001,N_17420,N_17330);
or U18002 (N_18002,N_17469,N_17628);
or U18003 (N_18003,N_17207,N_17570);
and U18004 (N_18004,N_17611,N_17390);
xor U18005 (N_18005,N_17164,N_17740);
xnor U18006 (N_18006,N_17173,N_17272);
and U18007 (N_18007,N_17528,N_17388);
xor U18008 (N_18008,N_17102,N_17025);
and U18009 (N_18009,N_17226,N_17526);
nor U18010 (N_18010,N_17683,N_17160);
nand U18011 (N_18011,N_17853,N_17678);
nand U18012 (N_18012,N_17136,N_17763);
xnor U18013 (N_18013,N_17240,N_17615);
and U18014 (N_18014,N_17162,N_17950);
or U18015 (N_18015,N_17022,N_17108);
nand U18016 (N_18016,N_17064,N_17491);
or U18017 (N_18017,N_17197,N_17281);
nor U18018 (N_18018,N_17474,N_17905);
nand U18019 (N_18019,N_17057,N_17632);
nor U18020 (N_18020,N_17573,N_17396);
nor U18021 (N_18021,N_17534,N_17169);
nand U18022 (N_18022,N_17540,N_17708);
nand U18023 (N_18023,N_17716,N_17581);
xnor U18024 (N_18024,N_17253,N_17044);
xnor U18025 (N_18025,N_17159,N_17873);
nand U18026 (N_18026,N_17870,N_17441);
and U18027 (N_18027,N_17743,N_17705);
or U18028 (N_18028,N_17052,N_17063);
and U18029 (N_18029,N_17435,N_17781);
and U18030 (N_18030,N_17869,N_17826);
or U18031 (N_18031,N_17881,N_17867);
nor U18032 (N_18032,N_17908,N_17132);
xor U18033 (N_18033,N_17470,N_17978);
xnor U18034 (N_18034,N_17018,N_17962);
or U18035 (N_18035,N_17624,N_17868);
or U18036 (N_18036,N_17412,N_17142);
xor U18037 (N_18037,N_17183,N_17442);
or U18038 (N_18038,N_17587,N_17985);
nor U18039 (N_18039,N_17560,N_17871);
nor U18040 (N_18040,N_17092,N_17097);
nand U18041 (N_18041,N_17859,N_17239);
and U18042 (N_18042,N_17769,N_17537);
nand U18043 (N_18043,N_17995,N_17167);
or U18044 (N_18044,N_17328,N_17075);
and U18045 (N_18045,N_17454,N_17400);
xnor U18046 (N_18046,N_17710,N_17764);
and U18047 (N_18047,N_17619,N_17360);
nand U18048 (N_18048,N_17082,N_17280);
and U18049 (N_18049,N_17277,N_17742);
or U18050 (N_18050,N_17847,N_17128);
or U18051 (N_18051,N_17292,N_17228);
nand U18052 (N_18052,N_17898,N_17450);
nor U18053 (N_18053,N_17449,N_17012);
or U18054 (N_18054,N_17610,N_17294);
nand U18055 (N_18055,N_17154,N_17359);
and U18056 (N_18056,N_17204,N_17163);
or U18057 (N_18057,N_17760,N_17773);
or U18058 (N_18058,N_17917,N_17275);
nor U18059 (N_18059,N_17739,N_17753);
or U18060 (N_18060,N_17844,N_17089);
or U18061 (N_18061,N_17525,N_17947);
or U18062 (N_18062,N_17045,N_17172);
xor U18063 (N_18063,N_17673,N_17270);
xor U18064 (N_18064,N_17602,N_17952);
or U18065 (N_18065,N_17567,N_17814);
nor U18066 (N_18066,N_17895,N_17717);
nand U18067 (N_18067,N_17839,N_17120);
or U18068 (N_18068,N_17616,N_17013);
xnor U18069 (N_18069,N_17955,N_17279);
nor U18070 (N_18070,N_17234,N_17588);
and U18071 (N_18071,N_17195,N_17715);
or U18072 (N_18072,N_17429,N_17417);
xnor U18073 (N_18073,N_17332,N_17033);
nand U18074 (N_18074,N_17000,N_17016);
or U18075 (N_18075,N_17464,N_17325);
nor U18076 (N_18076,N_17501,N_17953);
nor U18077 (N_18077,N_17011,N_17631);
and U18078 (N_18078,N_17451,N_17783);
and U18079 (N_18079,N_17662,N_17067);
and U18080 (N_18080,N_17660,N_17669);
and U18081 (N_18081,N_17973,N_17079);
or U18082 (N_18082,N_17608,N_17688);
or U18083 (N_18083,N_17819,N_17860);
xnor U18084 (N_18084,N_17583,N_17285);
nor U18085 (N_18085,N_17741,N_17636);
and U18086 (N_18086,N_17046,N_17943);
xnor U18087 (N_18087,N_17048,N_17490);
nor U18088 (N_18088,N_17841,N_17327);
nor U18089 (N_18089,N_17344,N_17070);
xor U18090 (N_18090,N_17352,N_17023);
nand U18091 (N_18091,N_17314,N_17145);
or U18092 (N_18092,N_17105,N_17768);
or U18093 (N_18093,N_17324,N_17809);
or U18094 (N_18094,N_17322,N_17405);
xor U18095 (N_18095,N_17559,N_17062);
or U18096 (N_18096,N_17093,N_17912);
nor U18097 (N_18097,N_17776,N_17732);
xor U18098 (N_18098,N_17911,N_17211);
xor U18099 (N_18099,N_17446,N_17989);
or U18100 (N_18100,N_17290,N_17557);
xnor U18101 (N_18101,N_17891,N_17134);
or U18102 (N_18102,N_17182,N_17810);
and U18103 (N_18103,N_17366,N_17730);
or U18104 (N_18104,N_17475,N_17457);
or U18105 (N_18105,N_17496,N_17794);
nor U18106 (N_18106,N_17889,N_17152);
or U18107 (N_18107,N_17627,N_17553);
and U18108 (N_18108,N_17830,N_17519);
xor U18109 (N_18109,N_17775,N_17124);
nand U18110 (N_18110,N_17568,N_17107);
or U18111 (N_18111,N_17357,N_17480);
and U18112 (N_18112,N_17695,N_17112);
nand U18113 (N_18113,N_17759,N_17960);
nor U18114 (N_18114,N_17121,N_17458);
nor U18115 (N_18115,N_17224,N_17196);
nor U18116 (N_18116,N_17828,N_17267);
nor U18117 (N_18117,N_17722,N_17591);
nand U18118 (N_18118,N_17148,N_17158);
nor U18119 (N_18119,N_17382,N_17300);
nand U18120 (N_18120,N_17903,N_17893);
or U18121 (N_18121,N_17203,N_17422);
and U18122 (N_18122,N_17969,N_17576);
nand U18123 (N_18123,N_17691,N_17482);
xnor U18124 (N_18124,N_17961,N_17178);
or U18125 (N_18125,N_17094,N_17367);
nor U18126 (N_18126,N_17268,N_17646);
nor U18127 (N_18127,N_17605,N_17055);
or U18128 (N_18128,N_17579,N_17265);
xnor U18129 (N_18129,N_17372,N_17304);
nor U18130 (N_18130,N_17424,N_17970);
nor U18131 (N_18131,N_17051,N_17817);
nor U18132 (N_18132,N_17342,N_17397);
or U18133 (N_18133,N_17109,N_17346);
or U18134 (N_18134,N_17416,N_17373);
nor U18135 (N_18135,N_17404,N_17735);
nand U18136 (N_18136,N_17982,N_17243);
nand U18137 (N_18137,N_17655,N_17700);
or U18138 (N_18138,N_17190,N_17029);
or U18139 (N_18139,N_17822,N_17551);
and U18140 (N_18140,N_17736,N_17877);
nor U18141 (N_18141,N_17718,N_17797);
xor U18142 (N_18142,N_17361,N_17244);
and U18143 (N_18143,N_17820,N_17073);
and U18144 (N_18144,N_17625,N_17785);
or U18145 (N_18145,N_17084,N_17326);
or U18146 (N_18146,N_17241,N_17927);
and U18147 (N_18147,N_17473,N_17758);
xor U18148 (N_18148,N_17791,N_17129);
nand U18149 (N_18149,N_17536,N_17374);
xnor U18150 (N_18150,N_17507,N_17362);
nand U18151 (N_18151,N_17825,N_17702);
and U18152 (N_18152,N_17495,N_17233);
xor U18153 (N_18153,N_17336,N_17799);
nand U18154 (N_18154,N_17042,N_17863);
nor U18155 (N_18155,N_17353,N_17020);
and U18156 (N_18156,N_17365,N_17981);
nor U18157 (N_18157,N_17640,N_17452);
or U18158 (N_18158,N_17530,N_17897);
xnor U18159 (N_18159,N_17558,N_17509);
and U18160 (N_18160,N_17017,N_17484);
nand U18161 (N_18161,N_17437,N_17461);
nor U18162 (N_18162,N_17147,N_17410);
and U18163 (N_18163,N_17283,N_17793);
or U18164 (N_18164,N_17790,N_17149);
and U18165 (N_18165,N_17512,N_17569);
and U18166 (N_18166,N_17652,N_17585);
nor U18167 (N_18167,N_17979,N_17816);
and U18168 (N_18168,N_17836,N_17561);
and U18169 (N_18169,N_17254,N_17493);
and U18170 (N_18170,N_17489,N_17286);
xor U18171 (N_18171,N_17726,N_17175);
nor U18172 (N_18172,N_17804,N_17199);
nand U18173 (N_18173,N_17038,N_17987);
and U18174 (N_18174,N_17078,N_17888);
nor U18175 (N_18175,N_17185,N_17407);
nand U18176 (N_18176,N_17010,N_17676);
and U18177 (N_18177,N_17053,N_17837);
xnor U18178 (N_18178,N_17131,N_17237);
nand U18179 (N_18179,N_17137,N_17754);
or U18180 (N_18180,N_17750,N_17174);
xor U18181 (N_18181,N_17906,N_17377);
or U18182 (N_18182,N_17261,N_17208);
and U18183 (N_18183,N_17633,N_17476);
nor U18184 (N_18184,N_17513,N_17021);
xnor U18185 (N_18185,N_17005,N_17313);
xnor U18186 (N_18186,N_17032,N_17414);
or U18187 (N_18187,N_17737,N_17647);
or U18188 (N_18188,N_17645,N_17186);
nor U18189 (N_18189,N_17266,N_17545);
xnor U18190 (N_18190,N_17941,N_17824);
xor U18191 (N_18191,N_17503,N_17031);
xnor U18192 (N_18192,N_17620,N_17614);
or U18193 (N_18193,N_17642,N_17245);
nand U18194 (N_18194,N_17713,N_17289);
nor U18195 (N_18195,N_17780,N_17077);
nor U18196 (N_18196,N_17936,N_17395);
or U18197 (N_18197,N_17250,N_17418);
and U18198 (N_18198,N_17546,N_17983);
xnor U18199 (N_18199,N_17938,N_17571);
or U18200 (N_18200,N_17747,N_17946);
xnor U18201 (N_18201,N_17466,N_17100);
xor U18202 (N_18202,N_17217,N_17968);
or U18203 (N_18203,N_17096,N_17385);
xnor U18204 (N_18204,N_17638,N_17765);
nor U18205 (N_18205,N_17522,N_17161);
nor U18206 (N_18206,N_17685,N_17965);
nor U18207 (N_18207,N_17320,N_17692);
xor U18208 (N_18208,N_17238,N_17727);
nand U18209 (N_18209,N_17179,N_17368);
nor U18210 (N_18210,N_17498,N_17572);
nor U18211 (N_18211,N_17942,N_17278);
nor U18212 (N_18212,N_17861,N_17574);
nand U18213 (N_18213,N_17838,N_17219);
or U18214 (N_18214,N_17216,N_17842);
nor U18215 (N_18215,N_17684,N_17225);
nor U18216 (N_18216,N_17532,N_17904);
and U18217 (N_18217,N_17671,N_17260);
and U18218 (N_18218,N_17866,N_17709);
nor U18219 (N_18219,N_17659,N_17047);
and U18220 (N_18220,N_17883,N_17439);
nor U18221 (N_18221,N_17515,N_17375);
and U18222 (N_18222,N_17188,N_17915);
or U18223 (N_18223,N_17363,N_17609);
xnor U18224 (N_18224,N_17510,N_17399);
nand U18225 (N_18225,N_17643,N_17200);
nand U18226 (N_18226,N_17919,N_17287);
or U18227 (N_18227,N_17805,N_17933);
nor U18228 (N_18228,N_17271,N_17777);
nor U18229 (N_18229,N_17056,N_17607);
nor U18230 (N_18230,N_17019,N_17027);
nor U18231 (N_18231,N_17831,N_17213);
nor U18232 (N_18232,N_17263,N_17555);
or U18233 (N_18233,N_17544,N_17594);
or U18234 (N_18234,N_17311,N_17511);
nor U18235 (N_18235,N_17117,N_17098);
nor U18236 (N_18236,N_17974,N_17542);
xnor U18237 (N_18237,N_17623,N_17920);
nor U18238 (N_18238,N_17516,N_17913);
xnor U18239 (N_18239,N_17222,N_17663);
xor U18240 (N_18240,N_17187,N_17975);
xnor U18241 (N_18241,N_17194,N_17562);
nand U18242 (N_18242,N_17833,N_17026);
or U18243 (N_18243,N_17438,N_17116);
xnor U18244 (N_18244,N_17629,N_17181);
xnor U18245 (N_18245,N_17002,N_17894);
nand U18246 (N_18246,N_17258,N_17832);
nand U18247 (N_18247,N_17189,N_17066);
xnor U18248 (N_18248,N_17508,N_17923);
nor U18249 (N_18249,N_17004,N_17592);
nor U18250 (N_18250,N_17293,N_17909);
nor U18251 (N_18251,N_17305,N_17319);
nor U18252 (N_18252,N_17786,N_17231);
nor U18253 (N_18253,N_17566,N_17598);
or U18254 (N_18254,N_17850,N_17980);
or U18255 (N_18255,N_17813,N_17714);
nand U18256 (N_18256,N_17426,N_17101);
xor U18257 (N_18257,N_17472,N_17945);
or U18258 (N_18258,N_17745,N_17329);
nand U18259 (N_18259,N_17886,N_17015);
or U18260 (N_18260,N_17934,N_17811);
nor U18261 (N_18261,N_17580,N_17334);
or U18262 (N_18262,N_17994,N_17806);
and U18263 (N_18263,N_17180,N_17111);
nand U18264 (N_18264,N_17230,N_17041);
nand U18265 (N_18265,N_17977,N_17593);
and U18266 (N_18266,N_17302,N_17672);
nor U18267 (N_18267,N_17539,N_17988);
and U18268 (N_18268,N_17409,N_17331);
and U18269 (N_18269,N_17282,N_17921);
and U18270 (N_18270,N_17141,N_17523);
and U18271 (N_18271,N_17756,N_17256);
nor U18272 (N_18272,N_17689,N_17486);
xor U18273 (N_18273,N_17209,N_17310);
and U18274 (N_18274,N_17706,N_17113);
or U18275 (N_18275,N_17900,N_17612);
xor U18276 (N_18276,N_17419,N_17088);
nor U18277 (N_18277,N_17453,N_17383);
xnor U18278 (N_18278,N_17462,N_17341);
nand U18279 (N_18279,N_17854,N_17455);
or U18280 (N_18280,N_17925,N_17746);
or U18281 (N_18281,N_17192,N_17351);
nor U18282 (N_18282,N_17648,N_17220);
nand U18283 (N_18283,N_17876,N_17389);
and U18284 (N_18284,N_17531,N_17413);
xor U18285 (N_18285,N_17445,N_17381);
nor U18286 (N_18286,N_17144,N_17885);
and U18287 (N_18287,N_17902,N_17644);
xnor U18288 (N_18288,N_17698,N_17630);
nor U18289 (N_18289,N_17227,N_17795);
or U18290 (N_18290,N_17533,N_17527);
nand U18291 (N_18291,N_17043,N_17924);
nor U18292 (N_18292,N_17864,N_17703);
nor U18293 (N_18293,N_17661,N_17401);
and U18294 (N_18294,N_17049,N_17236);
nand U18295 (N_18295,N_17007,N_17488);
and U18296 (N_18296,N_17514,N_17951);
xor U18297 (N_18297,N_17494,N_17862);
or U18298 (N_18298,N_17087,N_17725);
or U18299 (N_18299,N_17316,N_17882);
xor U18300 (N_18300,N_17738,N_17303);
xor U18301 (N_18301,N_17554,N_17080);
or U18302 (N_18302,N_17114,N_17931);
nor U18303 (N_18303,N_17541,N_17036);
and U18304 (N_18304,N_17914,N_17001);
nor U18305 (N_18305,N_17734,N_17723);
nand U18306 (N_18306,N_17719,N_17411);
nor U18307 (N_18307,N_17991,N_17667);
nor U18308 (N_18308,N_17617,N_17170);
and U18309 (N_18309,N_17502,N_17637);
or U18310 (N_18310,N_17586,N_17323);
and U18311 (N_18311,N_17668,N_17402);
nand U18312 (N_18312,N_17784,N_17613);
nor U18313 (N_18313,N_17966,N_17459);
or U18314 (N_18314,N_17932,N_17964);
or U18315 (N_18315,N_17517,N_17364);
xnor U18316 (N_18316,N_17796,N_17699);
nand U18317 (N_18317,N_17724,N_17653);
nand U18318 (N_18318,N_17529,N_17297);
nand U18319 (N_18319,N_17037,N_17815);
or U18320 (N_18320,N_17284,N_17857);
nand U18321 (N_18321,N_17246,N_17301);
nand U18322 (N_18322,N_17818,N_17986);
nor U18323 (N_18323,N_17014,N_17807);
or U18324 (N_18324,N_17050,N_17690);
nor U18325 (N_18325,N_17890,N_17421);
and U18326 (N_18326,N_17879,N_17262);
nand U18327 (N_18327,N_17059,N_17299);
xnor U18328 (N_18328,N_17218,N_17345);
xnor U18329 (N_18329,N_17247,N_17778);
and U18330 (N_18330,N_17855,N_17076);
or U18331 (N_18331,N_17376,N_17595);
nor U18332 (N_18332,N_17939,N_17681);
and U18333 (N_18333,N_17058,N_17214);
nor U18334 (N_18334,N_17696,N_17369);
or U18335 (N_18335,N_17394,N_17339);
nand U18336 (N_18336,N_17497,N_17343);
or U18337 (N_18337,N_17878,N_17845);
or U18338 (N_18338,N_17639,N_17427);
and U18339 (N_18339,N_17601,N_17433);
or U18340 (N_18340,N_17210,N_17748);
nand U18341 (N_18341,N_17153,N_17596);
nor U18342 (N_18342,N_17193,N_17835);
and U18343 (N_18343,N_17584,N_17992);
nand U18344 (N_18344,N_17321,N_17762);
or U18345 (N_18345,N_17370,N_17679);
and U18346 (N_18346,N_17654,N_17798);
xor U18347 (N_18347,N_17099,N_17171);
nand U18348 (N_18348,N_17779,N_17431);
nor U18349 (N_18349,N_17852,N_17808);
and U18350 (N_18350,N_17752,N_17801);
and U18351 (N_18351,N_17317,N_17378);
nand U18352 (N_18352,N_17848,N_17150);
and U18353 (N_18353,N_17884,N_17133);
xnor U18354 (N_18354,N_17693,N_17039);
xnor U18355 (N_18355,N_17535,N_17701);
or U18356 (N_18356,N_17770,N_17907);
nor U18357 (N_18357,N_17772,N_17274);
or U18358 (N_18358,N_17130,N_17665);
xor U18359 (N_18359,N_17697,N_17168);
xor U18360 (N_18360,N_17926,N_17634);
nor U18361 (N_18361,N_17358,N_17252);
xor U18362 (N_18362,N_17967,N_17095);
or U18363 (N_18363,N_17916,N_17589);
xnor U18364 (N_18364,N_17465,N_17728);
or U18365 (N_18365,N_17935,N_17151);
or U18366 (N_18366,N_17674,N_17205);
xor U18367 (N_18367,N_17434,N_17959);
and U18368 (N_18368,N_17354,N_17350);
nor U18369 (N_18369,N_17590,N_17664);
nand U18370 (N_18370,N_17972,N_17788);
xnor U18371 (N_18371,N_17447,N_17547);
xnor U18372 (N_18372,N_17408,N_17744);
xor U18373 (N_18373,N_17687,N_17846);
or U18374 (N_18374,N_17849,N_17006);
nand U18375 (N_18375,N_17680,N_17471);
and U18376 (N_18376,N_17198,N_17035);
xor U18377 (N_18377,N_17298,N_17757);
xnor U18378 (N_18378,N_17720,N_17157);
and U18379 (N_18379,N_17963,N_17123);
nor U18380 (N_18380,N_17065,N_17201);
xor U18381 (N_18381,N_17221,N_17191);
nand U18382 (N_18382,N_17309,N_17312);
or U18383 (N_18383,N_17307,N_17563);
nor U18384 (N_18384,N_17125,N_17071);
and U18385 (N_18385,N_17749,N_17468);
xor U18386 (N_18386,N_17443,N_17651);
nand U18387 (N_18387,N_17415,N_17949);
nand U18388 (N_18388,N_17393,N_17139);
xnor U18389 (N_18389,N_17009,N_17269);
or U18390 (N_18390,N_17984,N_17649);
xnor U18391 (N_18391,N_17229,N_17255);
nor U18392 (N_18392,N_17937,N_17249);
nand U18393 (N_18393,N_17500,N_17957);
nand U18394 (N_18394,N_17349,N_17792);
or U18395 (N_18395,N_17899,N_17524);
and U18396 (N_18396,N_17575,N_17721);
xor U18397 (N_18397,N_17034,N_17140);
nand U18398 (N_18398,N_17295,N_17333);
nand U18399 (N_18399,N_17086,N_17812);
xor U18400 (N_18400,N_17520,N_17751);
nand U18401 (N_18401,N_17618,N_17892);
nor U18402 (N_18402,N_17843,N_17481);
nand U18403 (N_18403,N_17003,N_17729);
nand U18404 (N_18404,N_17787,N_17521);
xnor U18405 (N_18405,N_17565,N_17731);
or U18406 (N_18406,N_17436,N_17040);
xor U18407 (N_18407,N_17971,N_17851);
nand U18408 (N_18408,N_17887,N_17800);
nor U18409 (N_18409,N_17487,N_17548);
and U18410 (N_18410,N_17288,N_17296);
nand U18411 (N_18411,N_17264,N_17155);
or U18412 (N_18412,N_17430,N_17103);
nor U18413 (N_18413,N_17767,N_17090);
or U18414 (N_18414,N_17956,N_17380);
or U18415 (N_18415,N_17143,N_17081);
nor U18416 (N_18416,N_17666,N_17990);
xor U18417 (N_18417,N_17564,N_17930);
or U18418 (N_18418,N_17872,N_17928);
xnor U18419 (N_18419,N_17896,N_17337);
nor U18420 (N_18420,N_17083,N_17996);
nand U18421 (N_18421,N_17184,N_17235);
nand U18422 (N_18422,N_17257,N_17444);
nand U18423 (N_18423,N_17707,N_17335);
and U18424 (N_18424,N_17135,N_17406);
and U18425 (N_18425,N_17068,N_17165);
and U18426 (N_18426,N_17504,N_17242);
or U18427 (N_18427,N_17126,N_17771);
nand U18428 (N_18428,N_17318,N_17552);
xor U18429 (N_18429,N_17483,N_17348);
nor U18430 (N_18430,N_17834,N_17206);
nand U18431 (N_18431,N_17384,N_17069);
and U18432 (N_18432,N_17918,N_17371);
or U18433 (N_18433,N_17479,N_17024);
xor U18434 (N_18434,N_17929,N_17550);
and U18435 (N_18435,N_17658,N_17432);
nand U18436 (N_18436,N_17641,N_17944);
xnor U18437 (N_18437,N_17428,N_17232);
or U18438 (N_18438,N_17463,N_17597);
xnor U18439 (N_18439,N_17338,N_17626);
xnor U18440 (N_18440,N_17085,N_17998);
or U18441 (N_18441,N_17347,N_17340);
nor U18442 (N_18442,N_17291,N_17823);
xor U18443 (N_18443,N_17061,N_17603);
or U18444 (N_18444,N_17711,N_17072);
xor U18445 (N_18445,N_17379,N_17761);
xor U18446 (N_18446,N_17766,N_17177);
nand U18447 (N_18447,N_17122,N_17622);
or U18448 (N_18448,N_17492,N_17621);
xor U18449 (N_18449,N_17600,N_17577);
nor U18450 (N_18450,N_17518,N_17485);
nand U18451 (N_18451,N_17677,N_17856);
and U18452 (N_18452,N_17146,N_17789);
xnor U18453 (N_18453,N_17874,N_17119);
xnor U18454 (N_18454,N_17940,N_17803);
xnor U18455 (N_18455,N_17276,N_17403);
and U18456 (N_18456,N_17138,N_17355);
and U18457 (N_18457,N_17456,N_17308);
nand U18458 (N_18458,N_17306,N_17901);
and U18459 (N_18459,N_17875,N_17506);
or U18460 (N_18460,N_17176,N_17997);
nand U18461 (N_18461,N_17993,N_17840);
and U18462 (N_18462,N_17212,N_17202);
and U18463 (N_18463,N_17556,N_17273);
or U18464 (N_18464,N_17391,N_17110);
xnor U18465 (N_18465,N_17423,N_17115);
nor U18466 (N_18466,N_17315,N_17712);
and U18467 (N_18467,N_17156,N_17578);
xnor U18468 (N_18468,N_17091,N_17682);
or U18469 (N_18469,N_17865,N_17802);
and U18470 (N_18470,N_17599,N_17106);
or U18471 (N_18471,N_17543,N_17606);
or U18472 (N_18472,N_17251,N_17398);
and U18473 (N_18473,N_17477,N_17074);
or U18474 (N_18474,N_17704,N_17008);
and U18475 (N_18475,N_17215,N_17440);
nand U18476 (N_18476,N_17774,N_17538);
nor U18477 (N_18477,N_17829,N_17582);
xor U18478 (N_18478,N_17166,N_17392);
nand U18479 (N_18479,N_17976,N_17030);
or U18480 (N_18480,N_17954,N_17733);
and U18481 (N_18481,N_17604,N_17910);
and U18482 (N_18482,N_17675,N_17880);
or U18483 (N_18483,N_17460,N_17118);
and U18484 (N_18484,N_17670,N_17922);
nand U18485 (N_18485,N_17060,N_17650);
or U18486 (N_18486,N_17425,N_17356);
xor U18487 (N_18487,N_17223,N_17686);
and U18488 (N_18488,N_17387,N_17948);
xnor U18489 (N_18489,N_17821,N_17858);
xor U18490 (N_18490,N_17999,N_17755);
or U18491 (N_18491,N_17505,N_17782);
nand U18492 (N_18492,N_17958,N_17054);
or U18493 (N_18493,N_17028,N_17248);
and U18494 (N_18494,N_17478,N_17635);
and U18495 (N_18495,N_17104,N_17499);
xor U18496 (N_18496,N_17259,N_17386);
and U18497 (N_18497,N_17467,N_17127);
and U18498 (N_18498,N_17549,N_17694);
xnor U18499 (N_18499,N_17827,N_17656);
xnor U18500 (N_18500,N_17235,N_17048);
nand U18501 (N_18501,N_17651,N_17642);
or U18502 (N_18502,N_17899,N_17877);
xnor U18503 (N_18503,N_17803,N_17032);
nor U18504 (N_18504,N_17025,N_17856);
nand U18505 (N_18505,N_17285,N_17272);
nand U18506 (N_18506,N_17715,N_17022);
and U18507 (N_18507,N_17235,N_17749);
xor U18508 (N_18508,N_17512,N_17637);
nor U18509 (N_18509,N_17146,N_17558);
nand U18510 (N_18510,N_17478,N_17772);
xor U18511 (N_18511,N_17995,N_17532);
nor U18512 (N_18512,N_17454,N_17956);
or U18513 (N_18513,N_17687,N_17291);
nand U18514 (N_18514,N_17772,N_17402);
xor U18515 (N_18515,N_17267,N_17236);
nor U18516 (N_18516,N_17630,N_17135);
nand U18517 (N_18517,N_17511,N_17936);
nand U18518 (N_18518,N_17186,N_17214);
and U18519 (N_18519,N_17608,N_17910);
nor U18520 (N_18520,N_17224,N_17348);
xnor U18521 (N_18521,N_17791,N_17992);
and U18522 (N_18522,N_17405,N_17757);
or U18523 (N_18523,N_17587,N_17585);
or U18524 (N_18524,N_17733,N_17382);
or U18525 (N_18525,N_17351,N_17662);
nor U18526 (N_18526,N_17837,N_17571);
xor U18527 (N_18527,N_17985,N_17439);
or U18528 (N_18528,N_17061,N_17987);
or U18529 (N_18529,N_17350,N_17484);
nor U18530 (N_18530,N_17138,N_17116);
nor U18531 (N_18531,N_17634,N_17321);
and U18532 (N_18532,N_17363,N_17492);
and U18533 (N_18533,N_17313,N_17547);
nand U18534 (N_18534,N_17503,N_17061);
nor U18535 (N_18535,N_17001,N_17235);
or U18536 (N_18536,N_17322,N_17355);
nor U18537 (N_18537,N_17843,N_17490);
xnor U18538 (N_18538,N_17915,N_17806);
nor U18539 (N_18539,N_17969,N_17304);
and U18540 (N_18540,N_17063,N_17640);
or U18541 (N_18541,N_17712,N_17199);
or U18542 (N_18542,N_17987,N_17049);
or U18543 (N_18543,N_17145,N_17893);
and U18544 (N_18544,N_17729,N_17903);
and U18545 (N_18545,N_17077,N_17448);
xor U18546 (N_18546,N_17268,N_17690);
and U18547 (N_18547,N_17001,N_17469);
nor U18548 (N_18548,N_17685,N_17859);
or U18549 (N_18549,N_17864,N_17854);
nand U18550 (N_18550,N_17551,N_17874);
nand U18551 (N_18551,N_17354,N_17160);
nand U18552 (N_18552,N_17658,N_17843);
or U18553 (N_18553,N_17522,N_17983);
xor U18554 (N_18554,N_17342,N_17555);
or U18555 (N_18555,N_17989,N_17627);
and U18556 (N_18556,N_17075,N_17495);
nor U18557 (N_18557,N_17443,N_17998);
and U18558 (N_18558,N_17621,N_17954);
nor U18559 (N_18559,N_17979,N_17296);
and U18560 (N_18560,N_17195,N_17828);
nand U18561 (N_18561,N_17904,N_17424);
nor U18562 (N_18562,N_17581,N_17010);
nand U18563 (N_18563,N_17748,N_17145);
xor U18564 (N_18564,N_17345,N_17134);
nor U18565 (N_18565,N_17590,N_17126);
nand U18566 (N_18566,N_17817,N_17989);
nor U18567 (N_18567,N_17216,N_17882);
nor U18568 (N_18568,N_17552,N_17751);
or U18569 (N_18569,N_17834,N_17546);
nand U18570 (N_18570,N_17162,N_17707);
and U18571 (N_18571,N_17099,N_17146);
nand U18572 (N_18572,N_17534,N_17598);
and U18573 (N_18573,N_17148,N_17959);
nor U18574 (N_18574,N_17654,N_17185);
nor U18575 (N_18575,N_17996,N_17343);
and U18576 (N_18576,N_17391,N_17742);
or U18577 (N_18577,N_17134,N_17696);
nand U18578 (N_18578,N_17380,N_17002);
nand U18579 (N_18579,N_17377,N_17930);
nand U18580 (N_18580,N_17640,N_17251);
xor U18581 (N_18581,N_17366,N_17087);
and U18582 (N_18582,N_17688,N_17291);
and U18583 (N_18583,N_17240,N_17090);
nor U18584 (N_18584,N_17678,N_17130);
xnor U18585 (N_18585,N_17663,N_17408);
xor U18586 (N_18586,N_17861,N_17959);
nand U18587 (N_18587,N_17176,N_17474);
nor U18588 (N_18588,N_17097,N_17293);
or U18589 (N_18589,N_17975,N_17700);
or U18590 (N_18590,N_17229,N_17359);
xnor U18591 (N_18591,N_17965,N_17219);
nand U18592 (N_18592,N_17798,N_17985);
nor U18593 (N_18593,N_17954,N_17481);
xnor U18594 (N_18594,N_17200,N_17460);
or U18595 (N_18595,N_17638,N_17251);
or U18596 (N_18596,N_17442,N_17232);
nor U18597 (N_18597,N_17608,N_17576);
nand U18598 (N_18598,N_17710,N_17310);
nor U18599 (N_18599,N_17349,N_17555);
nand U18600 (N_18600,N_17599,N_17515);
or U18601 (N_18601,N_17212,N_17405);
or U18602 (N_18602,N_17943,N_17224);
xor U18603 (N_18603,N_17250,N_17289);
xnor U18604 (N_18604,N_17138,N_17803);
or U18605 (N_18605,N_17123,N_17563);
nand U18606 (N_18606,N_17529,N_17907);
and U18607 (N_18607,N_17791,N_17716);
nor U18608 (N_18608,N_17693,N_17764);
and U18609 (N_18609,N_17376,N_17648);
nand U18610 (N_18610,N_17889,N_17426);
xnor U18611 (N_18611,N_17179,N_17280);
nand U18612 (N_18612,N_17122,N_17078);
or U18613 (N_18613,N_17827,N_17292);
nand U18614 (N_18614,N_17971,N_17867);
or U18615 (N_18615,N_17093,N_17016);
xor U18616 (N_18616,N_17190,N_17849);
nor U18617 (N_18617,N_17778,N_17183);
and U18618 (N_18618,N_17000,N_17650);
nand U18619 (N_18619,N_17657,N_17220);
nand U18620 (N_18620,N_17621,N_17985);
nor U18621 (N_18621,N_17840,N_17541);
nand U18622 (N_18622,N_17332,N_17802);
nor U18623 (N_18623,N_17879,N_17276);
nand U18624 (N_18624,N_17140,N_17677);
or U18625 (N_18625,N_17711,N_17788);
nor U18626 (N_18626,N_17478,N_17803);
or U18627 (N_18627,N_17036,N_17226);
xor U18628 (N_18628,N_17184,N_17154);
or U18629 (N_18629,N_17227,N_17301);
or U18630 (N_18630,N_17451,N_17823);
and U18631 (N_18631,N_17179,N_17602);
and U18632 (N_18632,N_17316,N_17124);
or U18633 (N_18633,N_17766,N_17676);
nor U18634 (N_18634,N_17874,N_17967);
nor U18635 (N_18635,N_17237,N_17060);
and U18636 (N_18636,N_17143,N_17366);
and U18637 (N_18637,N_17109,N_17253);
nand U18638 (N_18638,N_17844,N_17973);
nor U18639 (N_18639,N_17441,N_17723);
xnor U18640 (N_18640,N_17942,N_17600);
nand U18641 (N_18641,N_17769,N_17964);
nor U18642 (N_18642,N_17464,N_17927);
nor U18643 (N_18643,N_17633,N_17861);
nand U18644 (N_18644,N_17755,N_17352);
xnor U18645 (N_18645,N_17239,N_17664);
xnor U18646 (N_18646,N_17568,N_17704);
or U18647 (N_18647,N_17305,N_17708);
xnor U18648 (N_18648,N_17091,N_17737);
and U18649 (N_18649,N_17018,N_17344);
or U18650 (N_18650,N_17377,N_17876);
nor U18651 (N_18651,N_17494,N_17736);
nand U18652 (N_18652,N_17417,N_17584);
and U18653 (N_18653,N_17693,N_17476);
nand U18654 (N_18654,N_17316,N_17534);
xnor U18655 (N_18655,N_17856,N_17541);
nor U18656 (N_18656,N_17968,N_17026);
nor U18657 (N_18657,N_17450,N_17266);
xor U18658 (N_18658,N_17599,N_17472);
nand U18659 (N_18659,N_17915,N_17424);
nor U18660 (N_18660,N_17051,N_17003);
nand U18661 (N_18661,N_17243,N_17489);
or U18662 (N_18662,N_17619,N_17074);
nand U18663 (N_18663,N_17606,N_17505);
or U18664 (N_18664,N_17934,N_17421);
nand U18665 (N_18665,N_17418,N_17375);
and U18666 (N_18666,N_17954,N_17162);
and U18667 (N_18667,N_17207,N_17441);
or U18668 (N_18668,N_17198,N_17697);
and U18669 (N_18669,N_17209,N_17560);
nor U18670 (N_18670,N_17421,N_17508);
nand U18671 (N_18671,N_17535,N_17196);
nor U18672 (N_18672,N_17683,N_17975);
nor U18673 (N_18673,N_17846,N_17672);
nor U18674 (N_18674,N_17341,N_17206);
xor U18675 (N_18675,N_17899,N_17752);
xor U18676 (N_18676,N_17302,N_17491);
xnor U18677 (N_18677,N_17593,N_17582);
nand U18678 (N_18678,N_17905,N_17006);
nor U18679 (N_18679,N_17618,N_17895);
nand U18680 (N_18680,N_17160,N_17344);
or U18681 (N_18681,N_17156,N_17864);
or U18682 (N_18682,N_17636,N_17661);
and U18683 (N_18683,N_17628,N_17000);
nand U18684 (N_18684,N_17013,N_17828);
nand U18685 (N_18685,N_17098,N_17356);
xor U18686 (N_18686,N_17944,N_17409);
nand U18687 (N_18687,N_17619,N_17415);
nor U18688 (N_18688,N_17700,N_17009);
nand U18689 (N_18689,N_17394,N_17698);
nor U18690 (N_18690,N_17929,N_17726);
xnor U18691 (N_18691,N_17197,N_17223);
nor U18692 (N_18692,N_17032,N_17118);
and U18693 (N_18693,N_17658,N_17704);
and U18694 (N_18694,N_17151,N_17853);
or U18695 (N_18695,N_17784,N_17772);
nor U18696 (N_18696,N_17761,N_17233);
nor U18697 (N_18697,N_17174,N_17223);
or U18698 (N_18698,N_17698,N_17179);
or U18699 (N_18699,N_17358,N_17652);
nand U18700 (N_18700,N_17541,N_17455);
nor U18701 (N_18701,N_17575,N_17270);
and U18702 (N_18702,N_17512,N_17222);
xnor U18703 (N_18703,N_17175,N_17705);
xor U18704 (N_18704,N_17124,N_17944);
nand U18705 (N_18705,N_17946,N_17433);
xnor U18706 (N_18706,N_17186,N_17122);
nand U18707 (N_18707,N_17885,N_17442);
xor U18708 (N_18708,N_17300,N_17473);
xor U18709 (N_18709,N_17876,N_17969);
nor U18710 (N_18710,N_17947,N_17682);
and U18711 (N_18711,N_17739,N_17480);
xor U18712 (N_18712,N_17187,N_17675);
nor U18713 (N_18713,N_17116,N_17768);
or U18714 (N_18714,N_17760,N_17113);
nor U18715 (N_18715,N_17317,N_17259);
nor U18716 (N_18716,N_17133,N_17075);
xnor U18717 (N_18717,N_17350,N_17455);
or U18718 (N_18718,N_17070,N_17289);
or U18719 (N_18719,N_17977,N_17765);
nor U18720 (N_18720,N_17584,N_17954);
and U18721 (N_18721,N_17685,N_17015);
nand U18722 (N_18722,N_17674,N_17651);
or U18723 (N_18723,N_17764,N_17661);
and U18724 (N_18724,N_17735,N_17252);
nand U18725 (N_18725,N_17207,N_17616);
nand U18726 (N_18726,N_17787,N_17895);
or U18727 (N_18727,N_17806,N_17058);
or U18728 (N_18728,N_17382,N_17906);
nand U18729 (N_18729,N_17479,N_17912);
or U18730 (N_18730,N_17502,N_17244);
nor U18731 (N_18731,N_17909,N_17947);
and U18732 (N_18732,N_17721,N_17688);
nor U18733 (N_18733,N_17706,N_17638);
and U18734 (N_18734,N_17434,N_17476);
or U18735 (N_18735,N_17233,N_17805);
xor U18736 (N_18736,N_17419,N_17458);
and U18737 (N_18737,N_17870,N_17300);
nor U18738 (N_18738,N_17770,N_17706);
xor U18739 (N_18739,N_17608,N_17173);
and U18740 (N_18740,N_17523,N_17491);
nand U18741 (N_18741,N_17254,N_17224);
xor U18742 (N_18742,N_17016,N_17556);
xnor U18743 (N_18743,N_17259,N_17427);
xnor U18744 (N_18744,N_17441,N_17054);
xnor U18745 (N_18745,N_17924,N_17970);
and U18746 (N_18746,N_17694,N_17708);
and U18747 (N_18747,N_17909,N_17692);
nand U18748 (N_18748,N_17011,N_17404);
or U18749 (N_18749,N_17129,N_17627);
or U18750 (N_18750,N_17681,N_17310);
nand U18751 (N_18751,N_17625,N_17724);
or U18752 (N_18752,N_17348,N_17836);
xnor U18753 (N_18753,N_17574,N_17592);
nand U18754 (N_18754,N_17661,N_17064);
xor U18755 (N_18755,N_17015,N_17544);
xor U18756 (N_18756,N_17674,N_17806);
or U18757 (N_18757,N_17929,N_17723);
and U18758 (N_18758,N_17119,N_17209);
or U18759 (N_18759,N_17884,N_17293);
or U18760 (N_18760,N_17741,N_17733);
and U18761 (N_18761,N_17549,N_17660);
and U18762 (N_18762,N_17528,N_17625);
and U18763 (N_18763,N_17170,N_17303);
and U18764 (N_18764,N_17798,N_17146);
nor U18765 (N_18765,N_17440,N_17552);
nor U18766 (N_18766,N_17294,N_17366);
nor U18767 (N_18767,N_17312,N_17037);
nand U18768 (N_18768,N_17433,N_17608);
or U18769 (N_18769,N_17283,N_17230);
or U18770 (N_18770,N_17881,N_17344);
xnor U18771 (N_18771,N_17625,N_17574);
and U18772 (N_18772,N_17926,N_17474);
nor U18773 (N_18773,N_17169,N_17055);
nor U18774 (N_18774,N_17380,N_17614);
xnor U18775 (N_18775,N_17610,N_17408);
xor U18776 (N_18776,N_17705,N_17214);
nand U18777 (N_18777,N_17680,N_17476);
and U18778 (N_18778,N_17854,N_17981);
or U18779 (N_18779,N_17379,N_17527);
xnor U18780 (N_18780,N_17432,N_17960);
nor U18781 (N_18781,N_17769,N_17179);
or U18782 (N_18782,N_17976,N_17538);
nand U18783 (N_18783,N_17852,N_17577);
nor U18784 (N_18784,N_17381,N_17155);
or U18785 (N_18785,N_17740,N_17038);
nor U18786 (N_18786,N_17307,N_17293);
xor U18787 (N_18787,N_17348,N_17214);
or U18788 (N_18788,N_17917,N_17582);
xnor U18789 (N_18789,N_17204,N_17662);
nand U18790 (N_18790,N_17092,N_17330);
and U18791 (N_18791,N_17995,N_17459);
or U18792 (N_18792,N_17685,N_17358);
nand U18793 (N_18793,N_17615,N_17207);
nor U18794 (N_18794,N_17359,N_17399);
nor U18795 (N_18795,N_17673,N_17213);
nand U18796 (N_18796,N_17588,N_17662);
or U18797 (N_18797,N_17579,N_17969);
nor U18798 (N_18798,N_17302,N_17575);
xor U18799 (N_18799,N_17935,N_17398);
and U18800 (N_18800,N_17173,N_17891);
nor U18801 (N_18801,N_17267,N_17494);
and U18802 (N_18802,N_17072,N_17931);
or U18803 (N_18803,N_17796,N_17801);
and U18804 (N_18804,N_17627,N_17209);
nor U18805 (N_18805,N_17599,N_17134);
and U18806 (N_18806,N_17488,N_17796);
nand U18807 (N_18807,N_17711,N_17077);
and U18808 (N_18808,N_17336,N_17280);
xor U18809 (N_18809,N_17351,N_17847);
nand U18810 (N_18810,N_17347,N_17019);
or U18811 (N_18811,N_17097,N_17495);
xnor U18812 (N_18812,N_17609,N_17841);
xor U18813 (N_18813,N_17404,N_17733);
and U18814 (N_18814,N_17755,N_17976);
nor U18815 (N_18815,N_17956,N_17647);
xnor U18816 (N_18816,N_17427,N_17875);
or U18817 (N_18817,N_17551,N_17570);
nor U18818 (N_18818,N_17711,N_17985);
nor U18819 (N_18819,N_17741,N_17688);
or U18820 (N_18820,N_17030,N_17907);
xor U18821 (N_18821,N_17919,N_17997);
and U18822 (N_18822,N_17354,N_17244);
xor U18823 (N_18823,N_17682,N_17434);
xor U18824 (N_18824,N_17407,N_17638);
nor U18825 (N_18825,N_17044,N_17847);
nand U18826 (N_18826,N_17156,N_17590);
xnor U18827 (N_18827,N_17831,N_17758);
xnor U18828 (N_18828,N_17608,N_17328);
or U18829 (N_18829,N_17830,N_17337);
xor U18830 (N_18830,N_17976,N_17261);
nand U18831 (N_18831,N_17673,N_17287);
xnor U18832 (N_18832,N_17547,N_17194);
nand U18833 (N_18833,N_17254,N_17510);
nand U18834 (N_18834,N_17706,N_17170);
nand U18835 (N_18835,N_17778,N_17848);
nor U18836 (N_18836,N_17756,N_17236);
xor U18837 (N_18837,N_17345,N_17574);
nand U18838 (N_18838,N_17643,N_17167);
nand U18839 (N_18839,N_17047,N_17879);
xor U18840 (N_18840,N_17409,N_17150);
nand U18841 (N_18841,N_17427,N_17504);
and U18842 (N_18842,N_17363,N_17193);
nor U18843 (N_18843,N_17800,N_17006);
nor U18844 (N_18844,N_17755,N_17163);
nor U18845 (N_18845,N_17938,N_17840);
or U18846 (N_18846,N_17554,N_17896);
or U18847 (N_18847,N_17950,N_17671);
xnor U18848 (N_18848,N_17483,N_17678);
xnor U18849 (N_18849,N_17482,N_17525);
xor U18850 (N_18850,N_17441,N_17349);
nor U18851 (N_18851,N_17152,N_17953);
and U18852 (N_18852,N_17814,N_17265);
xnor U18853 (N_18853,N_17808,N_17003);
and U18854 (N_18854,N_17423,N_17020);
or U18855 (N_18855,N_17053,N_17034);
xor U18856 (N_18856,N_17911,N_17081);
nor U18857 (N_18857,N_17341,N_17218);
xor U18858 (N_18858,N_17183,N_17532);
xnor U18859 (N_18859,N_17448,N_17013);
nor U18860 (N_18860,N_17380,N_17872);
and U18861 (N_18861,N_17165,N_17222);
and U18862 (N_18862,N_17621,N_17861);
or U18863 (N_18863,N_17658,N_17539);
nand U18864 (N_18864,N_17417,N_17322);
nor U18865 (N_18865,N_17389,N_17294);
and U18866 (N_18866,N_17852,N_17585);
nor U18867 (N_18867,N_17391,N_17310);
and U18868 (N_18868,N_17433,N_17690);
nand U18869 (N_18869,N_17123,N_17483);
and U18870 (N_18870,N_17137,N_17331);
nand U18871 (N_18871,N_17268,N_17969);
nor U18872 (N_18872,N_17050,N_17439);
nand U18873 (N_18873,N_17389,N_17253);
and U18874 (N_18874,N_17592,N_17120);
nand U18875 (N_18875,N_17234,N_17323);
xnor U18876 (N_18876,N_17466,N_17727);
nor U18877 (N_18877,N_17453,N_17843);
nand U18878 (N_18878,N_17090,N_17845);
and U18879 (N_18879,N_17024,N_17062);
and U18880 (N_18880,N_17407,N_17621);
or U18881 (N_18881,N_17202,N_17765);
and U18882 (N_18882,N_17731,N_17010);
and U18883 (N_18883,N_17877,N_17119);
or U18884 (N_18884,N_17925,N_17862);
xnor U18885 (N_18885,N_17565,N_17634);
or U18886 (N_18886,N_17238,N_17781);
nand U18887 (N_18887,N_17996,N_17034);
or U18888 (N_18888,N_17290,N_17454);
or U18889 (N_18889,N_17460,N_17861);
nand U18890 (N_18890,N_17372,N_17484);
nand U18891 (N_18891,N_17906,N_17773);
nor U18892 (N_18892,N_17655,N_17560);
nand U18893 (N_18893,N_17173,N_17322);
or U18894 (N_18894,N_17509,N_17397);
or U18895 (N_18895,N_17177,N_17969);
nand U18896 (N_18896,N_17439,N_17408);
and U18897 (N_18897,N_17320,N_17973);
and U18898 (N_18898,N_17683,N_17331);
or U18899 (N_18899,N_17054,N_17261);
nor U18900 (N_18900,N_17861,N_17942);
and U18901 (N_18901,N_17059,N_17441);
or U18902 (N_18902,N_17130,N_17122);
xor U18903 (N_18903,N_17491,N_17067);
nand U18904 (N_18904,N_17965,N_17877);
or U18905 (N_18905,N_17067,N_17616);
xnor U18906 (N_18906,N_17861,N_17409);
nand U18907 (N_18907,N_17734,N_17268);
nand U18908 (N_18908,N_17406,N_17287);
xor U18909 (N_18909,N_17536,N_17300);
or U18910 (N_18910,N_17695,N_17867);
nand U18911 (N_18911,N_17363,N_17911);
nor U18912 (N_18912,N_17865,N_17843);
nor U18913 (N_18913,N_17060,N_17372);
nor U18914 (N_18914,N_17015,N_17695);
nand U18915 (N_18915,N_17135,N_17498);
nor U18916 (N_18916,N_17808,N_17175);
nand U18917 (N_18917,N_17340,N_17677);
or U18918 (N_18918,N_17665,N_17457);
and U18919 (N_18919,N_17624,N_17124);
or U18920 (N_18920,N_17109,N_17867);
or U18921 (N_18921,N_17926,N_17656);
xor U18922 (N_18922,N_17902,N_17525);
and U18923 (N_18923,N_17474,N_17641);
or U18924 (N_18924,N_17187,N_17846);
nand U18925 (N_18925,N_17752,N_17012);
or U18926 (N_18926,N_17907,N_17343);
nand U18927 (N_18927,N_17560,N_17214);
or U18928 (N_18928,N_17971,N_17935);
nand U18929 (N_18929,N_17039,N_17026);
nor U18930 (N_18930,N_17422,N_17117);
nor U18931 (N_18931,N_17121,N_17928);
nor U18932 (N_18932,N_17299,N_17662);
or U18933 (N_18933,N_17499,N_17544);
nand U18934 (N_18934,N_17265,N_17757);
or U18935 (N_18935,N_17259,N_17651);
nor U18936 (N_18936,N_17799,N_17737);
nor U18937 (N_18937,N_17903,N_17222);
nand U18938 (N_18938,N_17399,N_17033);
xnor U18939 (N_18939,N_17267,N_17343);
or U18940 (N_18940,N_17757,N_17980);
xor U18941 (N_18941,N_17994,N_17626);
or U18942 (N_18942,N_17342,N_17453);
nor U18943 (N_18943,N_17568,N_17844);
and U18944 (N_18944,N_17457,N_17989);
xnor U18945 (N_18945,N_17403,N_17758);
xor U18946 (N_18946,N_17506,N_17332);
and U18947 (N_18947,N_17244,N_17343);
xnor U18948 (N_18948,N_17839,N_17426);
xnor U18949 (N_18949,N_17990,N_17888);
and U18950 (N_18950,N_17734,N_17752);
xor U18951 (N_18951,N_17393,N_17130);
xor U18952 (N_18952,N_17631,N_17435);
nor U18953 (N_18953,N_17309,N_17728);
xnor U18954 (N_18954,N_17752,N_17170);
and U18955 (N_18955,N_17221,N_17732);
nand U18956 (N_18956,N_17976,N_17936);
or U18957 (N_18957,N_17947,N_17557);
nor U18958 (N_18958,N_17330,N_17827);
or U18959 (N_18959,N_17795,N_17477);
nand U18960 (N_18960,N_17570,N_17347);
or U18961 (N_18961,N_17890,N_17264);
nor U18962 (N_18962,N_17942,N_17986);
and U18963 (N_18963,N_17411,N_17739);
nand U18964 (N_18964,N_17027,N_17941);
xor U18965 (N_18965,N_17918,N_17417);
nand U18966 (N_18966,N_17852,N_17216);
nand U18967 (N_18967,N_17790,N_17702);
and U18968 (N_18968,N_17064,N_17269);
and U18969 (N_18969,N_17596,N_17530);
or U18970 (N_18970,N_17781,N_17428);
and U18971 (N_18971,N_17441,N_17134);
and U18972 (N_18972,N_17104,N_17079);
and U18973 (N_18973,N_17724,N_17934);
or U18974 (N_18974,N_17072,N_17923);
xnor U18975 (N_18975,N_17528,N_17248);
xnor U18976 (N_18976,N_17127,N_17172);
nand U18977 (N_18977,N_17958,N_17551);
and U18978 (N_18978,N_17189,N_17773);
and U18979 (N_18979,N_17277,N_17531);
nand U18980 (N_18980,N_17531,N_17998);
and U18981 (N_18981,N_17154,N_17302);
nand U18982 (N_18982,N_17326,N_17289);
or U18983 (N_18983,N_17394,N_17982);
nor U18984 (N_18984,N_17975,N_17428);
nand U18985 (N_18985,N_17009,N_17804);
nand U18986 (N_18986,N_17067,N_17382);
xnor U18987 (N_18987,N_17058,N_17629);
nand U18988 (N_18988,N_17911,N_17238);
xor U18989 (N_18989,N_17324,N_17562);
and U18990 (N_18990,N_17195,N_17988);
nor U18991 (N_18991,N_17638,N_17268);
nor U18992 (N_18992,N_17559,N_17705);
nand U18993 (N_18993,N_17285,N_17769);
or U18994 (N_18994,N_17974,N_17557);
or U18995 (N_18995,N_17108,N_17362);
nand U18996 (N_18996,N_17685,N_17723);
and U18997 (N_18997,N_17334,N_17102);
xnor U18998 (N_18998,N_17501,N_17571);
nand U18999 (N_18999,N_17738,N_17025);
and U19000 (N_19000,N_18467,N_18455);
xor U19001 (N_19001,N_18807,N_18628);
or U19002 (N_19002,N_18328,N_18035);
xor U19003 (N_19003,N_18161,N_18978);
or U19004 (N_19004,N_18793,N_18634);
nor U19005 (N_19005,N_18546,N_18712);
nor U19006 (N_19006,N_18139,N_18813);
nand U19007 (N_19007,N_18864,N_18305);
xnor U19008 (N_19008,N_18986,N_18195);
nand U19009 (N_19009,N_18934,N_18721);
and U19010 (N_19010,N_18181,N_18832);
nand U19011 (N_19011,N_18112,N_18523);
nand U19012 (N_19012,N_18771,N_18209);
nor U19013 (N_19013,N_18925,N_18326);
or U19014 (N_19014,N_18587,N_18974);
nor U19015 (N_19015,N_18069,N_18822);
xor U19016 (N_19016,N_18030,N_18155);
nor U19017 (N_19017,N_18208,N_18143);
and U19018 (N_19018,N_18798,N_18754);
xnor U19019 (N_19019,N_18599,N_18503);
and U19020 (N_19020,N_18735,N_18073);
or U19021 (N_19021,N_18037,N_18084);
xnor U19022 (N_19022,N_18741,N_18412);
or U19023 (N_19023,N_18931,N_18508);
or U19024 (N_19024,N_18258,N_18626);
or U19025 (N_19025,N_18423,N_18074);
nand U19026 (N_19026,N_18133,N_18980);
xnor U19027 (N_19027,N_18781,N_18576);
nand U19028 (N_19028,N_18678,N_18196);
and U19029 (N_19029,N_18891,N_18111);
and U19030 (N_19030,N_18645,N_18180);
nand U19031 (N_19031,N_18178,N_18880);
or U19032 (N_19032,N_18094,N_18827);
xnor U19033 (N_19033,N_18722,N_18640);
or U19034 (N_19034,N_18558,N_18225);
nor U19035 (N_19035,N_18128,N_18550);
and U19036 (N_19036,N_18581,N_18386);
and U19037 (N_19037,N_18522,N_18226);
nor U19038 (N_19038,N_18706,N_18145);
or U19039 (N_19039,N_18159,N_18200);
nor U19040 (N_19040,N_18856,N_18473);
xor U19041 (N_19041,N_18374,N_18618);
and U19042 (N_19042,N_18666,N_18376);
or U19043 (N_19043,N_18372,N_18766);
nor U19044 (N_19044,N_18013,N_18897);
or U19045 (N_19045,N_18760,N_18416);
nand U19046 (N_19046,N_18095,N_18500);
nor U19047 (N_19047,N_18932,N_18402);
or U19048 (N_19048,N_18987,N_18730);
or U19049 (N_19049,N_18044,N_18905);
nand U19050 (N_19050,N_18883,N_18898);
xnor U19051 (N_19051,N_18293,N_18674);
nor U19052 (N_19052,N_18965,N_18555);
nand U19053 (N_19053,N_18688,N_18795);
or U19054 (N_19054,N_18782,N_18750);
nor U19055 (N_19055,N_18260,N_18907);
nand U19056 (N_19056,N_18241,N_18440);
nand U19057 (N_19057,N_18027,N_18332);
xor U19058 (N_19058,N_18909,N_18227);
xor U19059 (N_19059,N_18794,N_18485);
nor U19060 (N_19060,N_18025,N_18203);
xnor U19061 (N_19061,N_18691,N_18290);
xnor U19062 (N_19062,N_18452,N_18163);
xnor U19063 (N_19063,N_18427,N_18769);
or U19064 (N_19064,N_18580,N_18739);
xor U19065 (N_19065,N_18863,N_18690);
xor U19066 (N_19066,N_18803,N_18786);
xnor U19067 (N_19067,N_18101,N_18784);
or U19068 (N_19068,N_18316,N_18421);
or U19069 (N_19069,N_18253,N_18825);
nand U19070 (N_19070,N_18379,N_18017);
nand U19071 (N_19071,N_18132,N_18933);
or U19072 (N_19072,N_18973,N_18943);
nor U19073 (N_19073,N_18623,N_18903);
nand U19074 (N_19074,N_18855,N_18515);
xor U19075 (N_19075,N_18240,N_18611);
nor U19076 (N_19076,N_18829,N_18056);
nor U19077 (N_19077,N_18296,N_18177);
nor U19078 (N_19078,N_18363,N_18921);
or U19079 (N_19079,N_18872,N_18759);
xnor U19080 (N_19080,N_18926,N_18425);
nor U19081 (N_19081,N_18709,N_18090);
or U19082 (N_19082,N_18248,N_18673);
nand U19083 (N_19083,N_18853,N_18341);
nor U19084 (N_19084,N_18560,N_18049);
xor U19085 (N_19085,N_18207,N_18594);
or U19086 (N_19086,N_18811,N_18968);
nor U19087 (N_19087,N_18499,N_18837);
nor U19088 (N_19088,N_18800,N_18588);
nand U19089 (N_19089,N_18950,N_18469);
nand U19090 (N_19090,N_18011,N_18420);
nor U19091 (N_19091,N_18551,N_18121);
and U19092 (N_19092,N_18359,N_18616);
nor U19093 (N_19093,N_18681,N_18610);
and U19094 (N_19094,N_18086,N_18243);
nand U19095 (N_19095,N_18938,N_18670);
xnor U19096 (N_19096,N_18762,N_18361);
nor U19097 (N_19097,N_18637,N_18512);
xor U19098 (N_19098,N_18405,N_18646);
xnor U19099 (N_19099,N_18816,N_18572);
nor U19100 (N_19100,N_18780,N_18530);
and U19101 (N_19101,N_18282,N_18257);
nor U19102 (N_19102,N_18998,N_18172);
nand U19103 (N_19103,N_18672,N_18411);
nor U19104 (N_19104,N_18235,N_18068);
xnor U19105 (N_19105,N_18930,N_18511);
xnor U19106 (N_19106,N_18350,N_18748);
xor U19107 (N_19107,N_18692,N_18841);
xor U19108 (N_19108,N_18561,N_18642);
xnor U19109 (N_19109,N_18527,N_18449);
or U19110 (N_19110,N_18726,N_18220);
nor U19111 (N_19111,N_18788,N_18668);
nand U19112 (N_19112,N_18040,N_18929);
and U19113 (N_19113,N_18614,N_18117);
or U19114 (N_19114,N_18582,N_18461);
nor U19115 (N_19115,N_18937,N_18124);
nor U19116 (N_19116,N_18357,N_18230);
nor U19117 (N_19117,N_18629,N_18325);
or U19118 (N_19118,N_18912,N_18462);
or U19119 (N_19119,N_18399,N_18349);
and U19120 (N_19120,N_18565,N_18767);
xnor U19121 (N_19121,N_18447,N_18949);
nor U19122 (N_19122,N_18322,N_18573);
nor U19123 (N_19123,N_18886,N_18358);
or U19124 (N_19124,N_18996,N_18222);
xor U19125 (N_19125,N_18571,N_18888);
and U19126 (N_19126,N_18955,N_18173);
or U19127 (N_19127,N_18605,N_18644);
nor U19128 (N_19128,N_18439,N_18197);
or U19129 (N_19129,N_18353,N_18205);
nand U19130 (N_19130,N_18776,N_18635);
xnor U19131 (N_19131,N_18983,N_18545);
and U19132 (N_19132,N_18924,N_18088);
xor U19133 (N_19133,N_18860,N_18979);
nand U19134 (N_19134,N_18517,N_18658);
nor U19135 (N_19135,N_18024,N_18403);
and U19136 (N_19136,N_18956,N_18892);
and U19137 (N_19137,N_18687,N_18204);
or U19138 (N_19138,N_18179,N_18714);
or U19139 (N_19139,N_18851,N_18971);
xor U19140 (N_19140,N_18650,N_18833);
nand U19141 (N_19141,N_18152,N_18792);
nor U19142 (N_19142,N_18061,N_18466);
nor U19143 (N_19143,N_18773,N_18737);
nor U19144 (N_19144,N_18859,N_18480);
nor U19145 (N_19145,N_18433,N_18337);
nand U19146 (N_19146,N_18871,N_18419);
nand U19147 (N_19147,N_18664,N_18339);
nor U19148 (N_19148,N_18779,N_18575);
xnor U19149 (N_19149,N_18064,N_18055);
and U19150 (N_19150,N_18394,N_18414);
nor U19151 (N_19151,N_18481,N_18382);
and U19152 (N_19152,N_18757,N_18228);
and U19153 (N_19153,N_18187,N_18752);
nand U19154 (N_19154,N_18964,N_18409);
xor U19155 (N_19155,N_18893,N_18510);
xnor U19156 (N_19156,N_18823,N_18778);
and U19157 (N_19157,N_18654,N_18150);
and U19158 (N_19158,N_18595,N_18244);
nor U19159 (N_19159,N_18118,N_18016);
or U19160 (N_19160,N_18742,N_18866);
xnor U19161 (N_19161,N_18834,N_18320);
nor U19162 (N_19162,N_18774,N_18237);
xor U19163 (N_19163,N_18321,N_18216);
or U19164 (N_19164,N_18703,N_18135);
and U19165 (N_19165,N_18516,N_18005);
and U19166 (N_19166,N_18506,N_18665);
nor U19167 (N_19167,N_18099,N_18952);
nor U19168 (N_19168,N_18895,N_18944);
xor U19169 (N_19169,N_18424,N_18190);
xnor U19170 (N_19170,N_18657,N_18395);
nor U19171 (N_19171,N_18518,N_18946);
nor U19172 (N_19172,N_18600,N_18570);
xor U19173 (N_19173,N_18749,N_18304);
xor U19174 (N_19174,N_18504,N_18319);
nor U19175 (N_19175,N_18854,N_18162);
xor U19176 (N_19176,N_18875,N_18023);
or U19177 (N_19177,N_18553,N_18578);
nand U19178 (N_19178,N_18492,N_18335);
and U19179 (N_19179,N_18694,N_18362);
nand U19180 (N_19180,N_18753,N_18972);
nor U19181 (N_19181,N_18347,N_18529);
nand U19182 (N_19182,N_18345,N_18431);
xor U19183 (N_19183,N_18874,N_18476);
xnor U19184 (N_19184,N_18062,N_18410);
and U19185 (N_19185,N_18001,N_18951);
nor U19186 (N_19186,N_18393,N_18331);
or U19187 (N_19187,N_18842,N_18879);
and U19188 (N_19188,N_18519,N_18259);
nand U19189 (N_19189,N_18606,N_18169);
and U19190 (N_19190,N_18942,N_18540);
and U19191 (N_19191,N_18102,N_18078);
or U19192 (N_19192,N_18836,N_18223);
and U19193 (N_19193,N_18632,N_18093);
nand U19194 (N_19194,N_18928,N_18217);
or U19195 (N_19195,N_18478,N_18494);
and U19196 (N_19196,N_18020,N_18444);
nor U19197 (N_19197,N_18450,N_18266);
xor U19198 (N_19198,N_18464,N_18218);
xor U19199 (N_19199,N_18718,N_18271);
xnor U19200 (N_19200,N_18238,N_18039);
nand U19201 (N_19201,N_18589,N_18520);
nand U19202 (N_19202,N_18434,N_18415);
and U19203 (N_19203,N_18627,N_18671);
nand U19204 (N_19204,N_18817,N_18488);
nor U19205 (N_19205,N_18848,N_18961);
and U19206 (N_19206,N_18913,N_18840);
nand U19207 (N_19207,N_18988,N_18513);
nand U19208 (N_19208,N_18563,N_18922);
nor U19209 (N_19209,N_18022,N_18075);
nand U19210 (N_19210,N_18630,N_18373);
nor U19211 (N_19211,N_18388,N_18564);
xor U19212 (N_19212,N_18438,N_18543);
nor U19213 (N_19213,N_18923,N_18999);
nor U19214 (N_19214,N_18806,N_18059);
and U19215 (N_19215,N_18535,N_18904);
xnor U19216 (N_19216,N_18125,N_18114);
xor U19217 (N_19217,N_18083,N_18761);
nand U19218 (N_19218,N_18812,N_18324);
nor U19219 (N_19219,N_18622,N_18170);
and U19220 (N_19220,N_18483,N_18655);
or U19221 (N_19221,N_18314,N_18046);
xnor U19222 (N_19222,N_18239,N_18604);
and U19223 (N_19223,N_18597,N_18050);
and U19224 (N_19224,N_18877,N_18232);
or U19225 (N_19225,N_18598,N_18249);
nor U19226 (N_19226,N_18824,N_18725);
xnor U19227 (N_19227,N_18698,N_18103);
and U19228 (N_19228,N_18734,N_18060);
nand U19229 (N_19229,N_18865,N_18995);
xor U19230 (N_19230,N_18847,N_18336);
nor U19231 (N_19231,N_18495,N_18389);
nor U19232 (N_19232,N_18213,N_18149);
nor U19233 (N_19233,N_18477,N_18524);
nor U19234 (N_19234,N_18183,N_18474);
xnor U19235 (N_19235,N_18219,N_18413);
nand U19236 (N_19236,N_18306,N_18648);
nor U19237 (N_19237,N_18280,N_18066);
nor U19238 (N_19238,N_18501,N_18269);
and U19239 (N_19239,N_18935,N_18384);
nand U19240 (N_19240,N_18625,N_18652);
and U19241 (N_19241,N_18174,N_18541);
and U19242 (N_19242,N_18579,N_18291);
nor U19243 (N_19243,N_18138,N_18406);
or U19244 (N_19244,N_18662,N_18590);
xnor U19245 (N_19245,N_18911,N_18082);
and U19246 (N_19246,N_18343,N_18437);
nand U19247 (N_19247,N_18435,N_18033);
and U19248 (N_19248,N_18583,N_18254);
and U19249 (N_19249,N_18298,N_18902);
nand U19250 (N_19250,N_18015,N_18008);
xor U19251 (N_19251,N_18954,N_18176);
xnor U19252 (N_19252,N_18707,N_18053);
and U19253 (N_19253,N_18299,N_18081);
or U19254 (N_19254,N_18356,N_18945);
and U19255 (N_19255,N_18593,N_18963);
nor U19256 (N_19256,N_18505,N_18596);
and U19257 (N_19257,N_18028,N_18366);
nand U19258 (N_19258,N_18380,N_18171);
or U19259 (N_19259,N_18818,N_18072);
and U19260 (N_19260,N_18791,N_18772);
nand U19261 (N_19261,N_18746,N_18882);
nand U19262 (N_19262,N_18327,N_18639);
nor U19263 (N_19263,N_18723,N_18071);
nor U19264 (N_19264,N_18043,N_18479);
nor U19265 (N_19265,N_18482,N_18839);
and U19266 (N_19266,N_18936,N_18309);
nor U19267 (N_19267,N_18901,N_18468);
nand U19268 (N_19268,N_18957,N_18586);
and U19269 (N_19269,N_18609,N_18591);
or U19270 (N_19270,N_18164,N_18262);
nand U19271 (N_19271,N_18815,N_18430);
nand U19272 (N_19272,N_18279,N_18636);
and U19273 (N_19273,N_18157,N_18287);
xor U19274 (N_19274,N_18387,N_18521);
or U19275 (N_19275,N_18313,N_18284);
nor U19276 (N_19276,N_18426,N_18976);
nand U19277 (N_19277,N_18041,N_18689);
nor U19278 (N_19278,N_18021,N_18148);
xnor U19279 (N_19279,N_18231,N_18264);
xor U19280 (N_19280,N_18770,N_18982);
xnor U19281 (N_19281,N_18808,N_18910);
and U19282 (N_19282,N_18908,N_18106);
xnor U19283 (N_19283,N_18250,N_18255);
nand U19284 (N_19284,N_18079,N_18984);
or U19285 (N_19285,N_18004,N_18026);
or U19286 (N_19286,N_18843,N_18899);
or U19287 (N_19287,N_18568,N_18693);
nor U19288 (N_19288,N_18211,N_18113);
nor U19289 (N_19289,N_18686,N_18036);
nand U19290 (N_19290,N_18397,N_18697);
nand U19291 (N_19291,N_18619,N_18768);
nand U19292 (N_19292,N_18184,N_18014);
and U19293 (N_19293,N_18775,N_18710);
xnor U19294 (N_19294,N_18493,N_18289);
nor U19295 (N_19295,N_18539,N_18799);
nor U19296 (N_19296,N_18070,N_18428);
or U19297 (N_19297,N_18105,N_18206);
xnor U19298 (N_19298,N_18089,N_18751);
xnor U19299 (N_19299,N_18323,N_18104);
and U19300 (N_19300,N_18276,N_18042);
nor U19301 (N_19301,N_18318,N_18058);
xnor U19302 (N_19302,N_18894,N_18338);
or U19303 (N_19303,N_18992,N_18756);
or U19304 (N_19304,N_18679,N_18229);
nor U19305 (N_19305,N_18265,N_18960);
nand U19306 (N_19306,N_18303,N_18065);
nor U19307 (N_19307,N_18740,N_18436);
or U19308 (N_19308,N_18547,N_18396);
or U19309 (N_19309,N_18900,N_18802);
nand U19310 (N_19310,N_18708,N_18116);
nor U19311 (N_19311,N_18989,N_18977);
and U19312 (N_19312,N_18920,N_18615);
nand U19313 (N_19313,N_18067,N_18985);
or U19314 (N_19314,N_18002,N_18683);
xor U19315 (N_19315,N_18919,N_18051);
xnor U19316 (N_19316,N_18562,N_18007);
nand U19317 (N_19317,N_18034,N_18057);
xor U19318 (N_19318,N_18914,N_18878);
xor U19319 (N_19319,N_18621,N_18077);
and U19320 (N_19320,N_18019,N_18263);
nor U19321 (N_19321,N_18185,N_18283);
and U19322 (N_19322,N_18317,N_18368);
xor U19323 (N_19323,N_18012,N_18472);
and U19324 (N_19324,N_18365,N_18454);
xor U19325 (N_19325,N_18141,N_18453);
xnor U19326 (N_19326,N_18542,N_18785);
or U19327 (N_19327,N_18463,N_18385);
xor U19328 (N_19328,N_18994,N_18234);
or U19329 (N_19329,N_18729,N_18755);
and U19330 (N_19330,N_18294,N_18548);
nand U19331 (N_19331,N_18010,N_18215);
nor U19332 (N_19332,N_18432,N_18881);
or U19333 (N_19333,N_18407,N_18641);
and U19334 (N_19334,N_18607,N_18857);
and U19335 (N_19335,N_18783,N_18491);
and U19336 (N_19336,N_18054,N_18814);
and U19337 (N_19337,N_18981,N_18507);
or U19338 (N_19338,N_18038,N_18165);
nor U19339 (N_19339,N_18873,N_18838);
or U19340 (N_19340,N_18702,N_18097);
or U19341 (N_19341,N_18156,N_18647);
and U19342 (N_19342,N_18018,N_18533);
nor U19343 (N_19343,N_18273,N_18191);
nand U19344 (N_19344,N_18804,N_18108);
or U19345 (N_19345,N_18009,N_18631);
nor U19346 (N_19346,N_18927,N_18889);
or U19347 (N_19347,N_18375,N_18032);
nand U19348 (N_19348,N_18828,N_18490);
nand U19349 (N_19349,N_18821,N_18601);
nand U19350 (N_19350,N_18868,N_18715);
or U19351 (N_19351,N_18918,N_18344);
or U19352 (N_19352,N_18758,N_18392);
nand U19353 (N_19353,N_18110,N_18682);
nand U19354 (N_19354,N_18603,N_18354);
and U19355 (N_19355,N_18651,N_18252);
xnor U19356 (N_19356,N_18997,N_18502);
or U19357 (N_19357,N_18123,N_18092);
and U19358 (N_19358,N_18370,N_18991);
xor U19359 (N_19359,N_18745,N_18704);
nor U19360 (N_19360,N_18278,N_18175);
nor U19361 (N_19361,N_18251,N_18790);
and U19362 (N_19362,N_18224,N_18958);
or U19363 (N_19363,N_18819,N_18085);
and U19364 (N_19364,N_18566,N_18429);
nor U19365 (N_19365,N_18966,N_18369);
or U19366 (N_19366,N_18471,N_18096);
nor U19367 (N_19367,N_18484,N_18858);
and U19368 (N_19368,N_18701,N_18787);
nor U19369 (N_19369,N_18267,N_18297);
nor U19370 (N_19370,N_18826,N_18401);
nor U19371 (N_19371,N_18574,N_18302);
and U19372 (N_19372,N_18584,N_18810);
and U19373 (N_19373,N_18360,N_18939);
and U19374 (N_19374,N_18448,N_18136);
nor U19375 (N_19375,N_18805,N_18340);
nor U19376 (N_19376,N_18569,N_18869);
nor U19377 (N_19377,N_18906,N_18835);
xor U19378 (N_19378,N_18941,N_18967);
nor U19379 (N_19379,N_18346,N_18592);
xnor U19380 (N_19380,N_18885,N_18459);
or U19381 (N_19381,N_18194,N_18048);
or U19382 (N_19382,N_18534,N_18137);
xnor U19383 (N_19383,N_18301,N_18556);
nand U19384 (N_19384,N_18975,N_18182);
xor U19385 (N_19385,N_18656,N_18765);
xnor U19386 (N_19386,N_18390,N_18383);
and U19387 (N_19387,N_18602,N_18724);
xor U19388 (N_19388,N_18210,N_18567);
xnor U19389 (N_19389,N_18391,N_18809);
or U19390 (N_19390,N_18355,N_18684);
and U19391 (N_19391,N_18441,N_18158);
and U19392 (N_19392,N_18916,N_18160);
nand U19393 (N_19393,N_18727,N_18091);
or U19394 (N_19394,N_18398,N_18418);
and U19395 (N_19395,N_18352,N_18214);
xnor U19396 (N_19396,N_18720,N_18514);
nand U19397 (N_19397,N_18199,N_18381);
nor U19398 (N_19398,N_18371,N_18245);
nand U19399 (N_19399,N_18470,N_18852);
and U19400 (N_19400,N_18212,N_18489);
or U19401 (N_19401,N_18310,N_18126);
nand U19402 (N_19402,N_18509,N_18270);
or U19403 (N_19403,N_18192,N_18029);
nand U19404 (N_19404,N_18763,N_18649);
xor U19405 (N_19405,N_18465,N_18342);
nand U19406 (N_19406,N_18457,N_18367);
or U19407 (N_19407,N_18451,N_18154);
xnor U19408 (N_19408,N_18890,N_18528);
nand U19409 (N_19409,N_18475,N_18617);
xor U19410 (N_19410,N_18680,N_18695);
xor U19411 (N_19411,N_18559,N_18732);
or U19412 (N_19412,N_18292,N_18861);
or U19413 (N_19413,N_18408,N_18236);
xnor U19414 (N_19414,N_18940,N_18286);
nor U19415 (N_19415,N_18764,N_18277);
or U19416 (N_19416,N_18953,N_18700);
nand U19417 (N_19417,N_18486,N_18127);
nand U19418 (N_19418,N_18536,N_18549);
and U19419 (N_19419,N_18031,N_18677);
and U19420 (N_19420,N_18711,N_18400);
xor U19421 (N_19421,N_18959,N_18884);
and U19422 (N_19422,N_18728,N_18846);
xor U19423 (N_19423,N_18738,N_18624);
xnor U19424 (N_19424,N_18844,N_18544);
nor U19425 (N_19425,N_18532,N_18312);
nand U19426 (N_19426,N_18947,N_18585);
and U19427 (N_19427,N_18676,N_18063);
xnor U19428 (N_19428,N_18643,N_18830);
xor U19429 (N_19429,N_18201,N_18256);
nand U19430 (N_19430,N_18076,N_18300);
nand U19431 (N_19431,N_18142,N_18458);
nor U19432 (N_19432,N_18189,N_18948);
nor U19433 (N_19433,N_18867,N_18969);
or U19434 (N_19434,N_18801,N_18261);
and U19435 (N_19435,N_18000,N_18743);
or U19436 (N_19436,N_18422,N_18417);
and U19437 (N_19437,N_18777,N_18717);
and U19438 (N_19438,N_18531,N_18120);
nor U19439 (N_19439,N_18736,N_18917);
xor U19440 (N_19440,N_18147,N_18198);
nor U19441 (N_19441,N_18744,N_18663);
nand U19442 (N_19442,N_18443,N_18202);
xnor U19443 (N_19443,N_18311,N_18896);
and U19444 (N_19444,N_18557,N_18456);
nor U19445 (N_19445,N_18006,N_18887);
nor U19446 (N_19446,N_18188,N_18122);
xnor U19447 (N_19447,N_18330,N_18329);
nor U19448 (N_19448,N_18705,N_18850);
xnor U19449 (N_19449,N_18608,N_18281);
nand U19450 (N_19450,N_18334,N_18993);
nor U19451 (N_19451,N_18307,N_18849);
nor U19452 (N_19452,N_18538,N_18633);
or U19453 (N_19453,N_18696,N_18990);
xor U19454 (N_19454,N_18915,N_18377);
nor U19455 (N_19455,N_18446,N_18612);
or U19456 (N_19456,N_18554,N_18699);
xnor U19457 (N_19457,N_18130,N_18268);
or U19458 (N_19458,N_18168,N_18525);
and U19459 (N_19459,N_18247,N_18667);
and U19460 (N_19460,N_18107,N_18552);
nor U19461 (N_19461,N_18080,N_18140);
xnor U19462 (N_19462,N_18747,N_18333);
nor U19463 (N_19463,N_18167,N_18719);
xnor U19464 (N_19464,N_18460,N_18134);
and U19465 (N_19465,N_18620,N_18193);
and U19466 (N_19466,N_18870,N_18144);
or U19467 (N_19467,N_18308,N_18100);
nor U19468 (N_19468,N_18675,N_18288);
and U19469 (N_19469,N_18404,N_18796);
and U19470 (N_19470,N_18045,N_18862);
and U19471 (N_19471,N_18831,N_18351);
nand U19472 (N_19472,N_18242,N_18713);
nand U19473 (N_19473,N_18497,N_18526);
xnor U19474 (N_19474,N_18146,N_18845);
or U19475 (N_19475,N_18716,N_18378);
nor U19476 (N_19476,N_18445,N_18274);
nand U19477 (N_19477,N_18315,N_18087);
xor U19478 (N_19478,N_18498,N_18186);
nand U19479 (N_19479,N_18537,N_18653);
and U19480 (N_19480,N_18577,N_18496);
or U19481 (N_19481,N_18275,N_18487);
or U19482 (N_19482,N_18295,N_18233);
nand U19483 (N_19483,N_18153,N_18659);
and U19484 (N_19484,N_18285,N_18109);
nand U19485 (N_19485,N_18131,N_18364);
or U19486 (N_19486,N_18272,N_18731);
nor U19487 (N_19487,N_18660,N_18166);
or U19488 (N_19488,N_18613,N_18003);
and U19489 (N_19489,N_18789,N_18119);
or U19490 (N_19490,N_18129,N_18876);
or U19491 (N_19491,N_18047,N_18246);
nand U19492 (N_19492,N_18685,N_18098);
and U19493 (N_19493,N_18115,N_18052);
xnor U19494 (N_19494,N_18348,N_18797);
and U19495 (N_19495,N_18962,N_18820);
nand U19496 (N_19496,N_18661,N_18733);
or U19497 (N_19497,N_18151,N_18970);
or U19498 (N_19498,N_18638,N_18669);
nor U19499 (N_19499,N_18221,N_18442);
nand U19500 (N_19500,N_18339,N_18310);
and U19501 (N_19501,N_18187,N_18858);
nand U19502 (N_19502,N_18770,N_18134);
nor U19503 (N_19503,N_18702,N_18238);
nor U19504 (N_19504,N_18689,N_18405);
nor U19505 (N_19505,N_18238,N_18235);
and U19506 (N_19506,N_18010,N_18180);
xor U19507 (N_19507,N_18674,N_18348);
xnor U19508 (N_19508,N_18300,N_18476);
nand U19509 (N_19509,N_18719,N_18873);
and U19510 (N_19510,N_18295,N_18183);
nand U19511 (N_19511,N_18075,N_18313);
xnor U19512 (N_19512,N_18607,N_18944);
xor U19513 (N_19513,N_18934,N_18601);
nor U19514 (N_19514,N_18993,N_18748);
nand U19515 (N_19515,N_18933,N_18789);
nand U19516 (N_19516,N_18119,N_18467);
nor U19517 (N_19517,N_18924,N_18496);
or U19518 (N_19518,N_18064,N_18635);
xnor U19519 (N_19519,N_18598,N_18403);
and U19520 (N_19520,N_18999,N_18378);
nor U19521 (N_19521,N_18006,N_18112);
nor U19522 (N_19522,N_18917,N_18210);
nor U19523 (N_19523,N_18672,N_18828);
nand U19524 (N_19524,N_18898,N_18648);
or U19525 (N_19525,N_18460,N_18275);
nand U19526 (N_19526,N_18151,N_18349);
or U19527 (N_19527,N_18372,N_18264);
nor U19528 (N_19528,N_18573,N_18977);
xnor U19529 (N_19529,N_18764,N_18159);
xnor U19530 (N_19530,N_18452,N_18982);
and U19531 (N_19531,N_18204,N_18092);
and U19532 (N_19532,N_18936,N_18254);
and U19533 (N_19533,N_18482,N_18585);
nor U19534 (N_19534,N_18114,N_18189);
nand U19535 (N_19535,N_18247,N_18343);
nand U19536 (N_19536,N_18673,N_18680);
nor U19537 (N_19537,N_18764,N_18443);
and U19538 (N_19538,N_18711,N_18046);
and U19539 (N_19539,N_18586,N_18671);
nor U19540 (N_19540,N_18300,N_18072);
nand U19541 (N_19541,N_18464,N_18767);
nand U19542 (N_19542,N_18544,N_18396);
xnor U19543 (N_19543,N_18151,N_18856);
and U19544 (N_19544,N_18810,N_18652);
or U19545 (N_19545,N_18219,N_18505);
and U19546 (N_19546,N_18542,N_18632);
nor U19547 (N_19547,N_18827,N_18584);
and U19548 (N_19548,N_18242,N_18460);
nand U19549 (N_19549,N_18659,N_18507);
nor U19550 (N_19550,N_18793,N_18486);
and U19551 (N_19551,N_18733,N_18326);
or U19552 (N_19552,N_18494,N_18991);
xnor U19553 (N_19553,N_18279,N_18658);
nor U19554 (N_19554,N_18521,N_18132);
xnor U19555 (N_19555,N_18499,N_18079);
xnor U19556 (N_19556,N_18961,N_18612);
nor U19557 (N_19557,N_18548,N_18789);
nor U19558 (N_19558,N_18495,N_18566);
nand U19559 (N_19559,N_18321,N_18607);
nand U19560 (N_19560,N_18514,N_18838);
xor U19561 (N_19561,N_18351,N_18095);
nor U19562 (N_19562,N_18986,N_18871);
nand U19563 (N_19563,N_18978,N_18038);
nand U19564 (N_19564,N_18749,N_18624);
nand U19565 (N_19565,N_18968,N_18200);
or U19566 (N_19566,N_18443,N_18393);
nor U19567 (N_19567,N_18191,N_18375);
and U19568 (N_19568,N_18825,N_18773);
or U19569 (N_19569,N_18509,N_18700);
nor U19570 (N_19570,N_18954,N_18320);
or U19571 (N_19571,N_18016,N_18379);
or U19572 (N_19572,N_18218,N_18849);
or U19573 (N_19573,N_18208,N_18674);
or U19574 (N_19574,N_18814,N_18113);
and U19575 (N_19575,N_18757,N_18644);
nand U19576 (N_19576,N_18816,N_18841);
nand U19577 (N_19577,N_18401,N_18269);
or U19578 (N_19578,N_18882,N_18363);
nor U19579 (N_19579,N_18806,N_18180);
nand U19580 (N_19580,N_18723,N_18356);
xnor U19581 (N_19581,N_18827,N_18154);
and U19582 (N_19582,N_18683,N_18985);
and U19583 (N_19583,N_18564,N_18164);
and U19584 (N_19584,N_18782,N_18158);
and U19585 (N_19585,N_18262,N_18105);
or U19586 (N_19586,N_18721,N_18123);
nor U19587 (N_19587,N_18484,N_18722);
xnor U19588 (N_19588,N_18972,N_18984);
or U19589 (N_19589,N_18477,N_18181);
xnor U19590 (N_19590,N_18862,N_18369);
and U19591 (N_19591,N_18167,N_18248);
nor U19592 (N_19592,N_18267,N_18048);
xnor U19593 (N_19593,N_18228,N_18372);
or U19594 (N_19594,N_18914,N_18223);
nor U19595 (N_19595,N_18513,N_18706);
or U19596 (N_19596,N_18402,N_18251);
nor U19597 (N_19597,N_18237,N_18633);
and U19598 (N_19598,N_18132,N_18420);
nor U19599 (N_19599,N_18323,N_18764);
nor U19600 (N_19600,N_18305,N_18018);
xor U19601 (N_19601,N_18016,N_18054);
nor U19602 (N_19602,N_18079,N_18974);
nor U19603 (N_19603,N_18219,N_18693);
nor U19604 (N_19604,N_18659,N_18329);
and U19605 (N_19605,N_18988,N_18844);
and U19606 (N_19606,N_18342,N_18374);
or U19607 (N_19607,N_18883,N_18529);
nor U19608 (N_19608,N_18080,N_18659);
or U19609 (N_19609,N_18723,N_18332);
nor U19610 (N_19610,N_18591,N_18640);
or U19611 (N_19611,N_18220,N_18115);
nor U19612 (N_19612,N_18046,N_18246);
nor U19613 (N_19613,N_18642,N_18428);
nand U19614 (N_19614,N_18027,N_18723);
nor U19615 (N_19615,N_18419,N_18396);
xor U19616 (N_19616,N_18339,N_18497);
or U19617 (N_19617,N_18241,N_18568);
and U19618 (N_19618,N_18814,N_18718);
nor U19619 (N_19619,N_18592,N_18591);
and U19620 (N_19620,N_18098,N_18142);
or U19621 (N_19621,N_18667,N_18016);
nand U19622 (N_19622,N_18527,N_18886);
and U19623 (N_19623,N_18406,N_18146);
and U19624 (N_19624,N_18289,N_18998);
xor U19625 (N_19625,N_18774,N_18674);
and U19626 (N_19626,N_18261,N_18028);
and U19627 (N_19627,N_18877,N_18681);
nand U19628 (N_19628,N_18230,N_18665);
or U19629 (N_19629,N_18106,N_18674);
and U19630 (N_19630,N_18065,N_18204);
and U19631 (N_19631,N_18312,N_18009);
and U19632 (N_19632,N_18837,N_18714);
xnor U19633 (N_19633,N_18753,N_18206);
xnor U19634 (N_19634,N_18088,N_18118);
nor U19635 (N_19635,N_18149,N_18155);
or U19636 (N_19636,N_18293,N_18138);
nor U19637 (N_19637,N_18432,N_18015);
and U19638 (N_19638,N_18874,N_18567);
and U19639 (N_19639,N_18147,N_18106);
nand U19640 (N_19640,N_18702,N_18376);
and U19641 (N_19641,N_18845,N_18998);
and U19642 (N_19642,N_18158,N_18678);
xor U19643 (N_19643,N_18124,N_18585);
nand U19644 (N_19644,N_18104,N_18953);
xor U19645 (N_19645,N_18261,N_18054);
xnor U19646 (N_19646,N_18757,N_18612);
nand U19647 (N_19647,N_18518,N_18532);
xor U19648 (N_19648,N_18801,N_18009);
xnor U19649 (N_19649,N_18914,N_18780);
and U19650 (N_19650,N_18183,N_18522);
nor U19651 (N_19651,N_18874,N_18123);
or U19652 (N_19652,N_18890,N_18801);
nor U19653 (N_19653,N_18137,N_18599);
and U19654 (N_19654,N_18492,N_18487);
nand U19655 (N_19655,N_18255,N_18736);
xor U19656 (N_19656,N_18276,N_18567);
or U19657 (N_19657,N_18136,N_18518);
or U19658 (N_19658,N_18518,N_18237);
xnor U19659 (N_19659,N_18051,N_18306);
nand U19660 (N_19660,N_18117,N_18845);
and U19661 (N_19661,N_18452,N_18200);
nand U19662 (N_19662,N_18578,N_18219);
and U19663 (N_19663,N_18034,N_18938);
xor U19664 (N_19664,N_18854,N_18465);
xnor U19665 (N_19665,N_18326,N_18972);
nor U19666 (N_19666,N_18297,N_18895);
or U19667 (N_19667,N_18706,N_18836);
nand U19668 (N_19668,N_18263,N_18648);
and U19669 (N_19669,N_18708,N_18267);
nor U19670 (N_19670,N_18247,N_18690);
xnor U19671 (N_19671,N_18387,N_18210);
or U19672 (N_19672,N_18515,N_18950);
nor U19673 (N_19673,N_18770,N_18550);
xnor U19674 (N_19674,N_18389,N_18816);
and U19675 (N_19675,N_18131,N_18219);
xnor U19676 (N_19676,N_18200,N_18989);
nor U19677 (N_19677,N_18635,N_18347);
xnor U19678 (N_19678,N_18207,N_18624);
and U19679 (N_19679,N_18625,N_18823);
or U19680 (N_19680,N_18700,N_18216);
and U19681 (N_19681,N_18516,N_18761);
nor U19682 (N_19682,N_18186,N_18366);
or U19683 (N_19683,N_18757,N_18171);
or U19684 (N_19684,N_18843,N_18583);
nand U19685 (N_19685,N_18856,N_18091);
xor U19686 (N_19686,N_18987,N_18927);
or U19687 (N_19687,N_18273,N_18964);
or U19688 (N_19688,N_18607,N_18874);
and U19689 (N_19689,N_18062,N_18523);
and U19690 (N_19690,N_18518,N_18369);
xor U19691 (N_19691,N_18068,N_18812);
or U19692 (N_19692,N_18838,N_18761);
nor U19693 (N_19693,N_18957,N_18734);
nor U19694 (N_19694,N_18915,N_18135);
and U19695 (N_19695,N_18947,N_18146);
or U19696 (N_19696,N_18531,N_18773);
or U19697 (N_19697,N_18717,N_18224);
and U19698 (N_19698,N_18276,N_18899);
nand U19699 (N_19699,N_18852,N_18539);
nor U19700 (N_19700,N_18279,N_18033);
and U19701 (N_19701,N_18382,N_18397);
nor U19702 (N_19702,N_18205,N_18343);
or U19703 (N_19703,N_18966,N_18128);
nand U19704 (N_19704,N_18512,N_18682);
and U19705 (N_19705,N_18128,N_18302);
nor U19706 (N_19706,N_18957,N_18689);
nor U19707 (N_19707,N_18757,N_18945);
nor U19708 (N_19708,N_18640,N_18843);
nand U19709 (N_19709,N_18760,N_18858);
nor U19710 (N_19710,N_18546,N_18894);
nand U19711 (N_19711,N_18942,N_18395);
and U19712 (N_19712,N_18814,N_18828);
and U19713 (N_19713,N_18260,N_18071);
and U19714 (N_19714,N_18486,N_18417);
and U19715 (N_19715,N_18012,N_18495);
nand U19716 (N_19716,N_18720,N_18692);
nor U19717 (N_19717,N_18381,N_18527);
and U19718 (N_19718,N_18118,N_18362);
xnor U19719 (N_19719,N_18459,N_18547);
xor U19720 (N_19720,N_18175,N_18846);
xnor U19721 (N_19721,N_18279,N_18854);
nand U19722 (N_19722,N_18238,N_18883);
nor U19723 (N_19723,N_18454,N_18533);
xnor U19724 (N_19724,N_18356,N_18242);
xnor U19725 (N_19725,N_18093,N_18248);
or U19726 (N_19726,N_18423,N_18958);
xor U19727 (N_19727,N_18093,N_18116);
nand U19728 (N_19728,N_18471,N_18807);
nand U19729 (N_19729,N_18627,N_18764);
or U19730 (N_19730,N_18529,N_18918);
nand U19731 (N_19731,N_18917,N_18134);
or U19732 (N_19732,N_18665,N_18996);
xor U19733 (N_19733,N_18893,N_18122);
or U19734 (N_19734,N_18606,N_18802);
or U19735 (N_19735,N_18759,N_18047);
xnor U19736 (N_19736,N_18167,N_18723);
and U19737 (N_19737,N_18124,N_18389);
and U19738 (N_19738,N_18627,N_18933);
nand U19739 (N_19739,N_18453,N_18160);
xnor U19740 (N_19740,N_18559,N_18811);
and U19741 (N_19741,N_18099,N_18678);
nor U19742 (N_19742,N_18561,N_18941);
nand U19743 (N_19743,N_18522,N_18716);
xnor U19744 (N_19744,N_18339,N_18164);
nor U19745 (N_19745,N_18997,N_18628);
and U19746 (N_19746,N_18474,N_18152);
nand U19747 (N_19747,N_18630,N_18641);
nand U19748 (N_19748,N_18723,N_18515);
or U19749 (N_19749,N_18822,N_18443);
xor U19750 (N_19750,N_18554,N_18388);
nand U19751 (N_19751,N_18312,N_18293);
nor U19752 (N_19752,N_18963,N_18867);
or U19753 (N_19753,N_18550,N_18522);
nand U19754 (N_19754,N_18285,N_18313);
nand U19755 (N_19755,N_18622,N_18467);
or U19756 (N_19756,N_18131,N_18193);
xor U19757 (N_19757,N_18527,N_18027);
nor U19758 (N_19758,N_18080,N_18451);
nand U19759 (N_19759,N_18927,N_18857);
and U19760 (N_19760,N_18753,N_18672);
and U19761 (N_19761,N_18030,N_18575);
nor U19762 (N_19762,N_18896,N_18603);
and U19763 (N_19763,N_18008,N_18606);
and U19764 (N_19764,N_18225,N_18890);
nand U19765 (N_19765,N_18321,N_18487);
nand U19766 (N_19766,N_18698,N_18638);
xnor U19767 (N_19767,N_18235,N_18687);
and U19768 (N_19768,N_18584,N_18747);
nand U19769 (N_19769,N_18669,N_18075);
nor U19770 (N_19770,N_18005,N_18693);
nand U19771 (N_19771,N_18333,N_18766);
nor U19772 (N_19772,N_18289,N_18360);
nor U19773 (N_19773,N_18471,N_18118);
nor U19774 (N_19774,N_18882,N_18817);
and U19775 (N_19775,N_18906,N_18238);
and U19776 (N_19776,N_18864,N_18640);
xor U19777 (N_19777,N_18576,N_18048);
or U19778 (N_19778,N_18548,N_18487);
nor U19779 (N_19779,N_18690,N_18908);
and U19780 (N_19780,N_18052,N_18522);
nand U19781 (N_19781,N_18172,N_18955);
nor U19782 (N_19782,N_18452,N_18135);
nor U19783 (N_19783,N_18625,N_18760);
nand U19784 (N_19784,N_18634,N_18465);
or U19785 (N_19785,N_18736,N_18654);
xnor U19786 (N_19786,N_18278,N_18500);
xnor U19787 (N_19787,N_18326,N_18047);
nand U19788 (N_19788,N_18719,N_18902);
nand U19789 (N_19789,N_18002,N_18676);
xnor U19790 (N_19790,N_18278,N_18787);
xor U19791 (N_19791,N_18068,N_18363);
nor U19792 (N_19792,N_18896,N_18030);
nor U19793 (N_19793,N_18129,N_18912);
and U19794 (N_19794,N_18778,N_18268);
and U19795 (N_19795,N_18668,N_18613);
or U19796 (N_19796,N_18916,N_18634);
or U19797 (N_19797,N_18048,N_18253);
nand U19798 (N_19798,N_18786,N_18027);
nor U19799 (N_19799,N_18112,N_18971);
or U19800 (N_19800,N_18676,N_18591);
or U19801 (N_19801,N_18239,N_18586);
nor U19802 (N_19802,N_18357,N_18429);
and U19803 (N_19803,N_18793,N_18352);
nand U19804 (N_19804,N_18245,N_18819);
xor U19805 (N_19805,N_18529,N_18055);
and U19806 (N_19806,N_18553,N_18233);
or U19807 (N_19807,N_18632,N_18575);
and U19808 (N_19808,N_18618,N_18961);
xnor U19809 (N_19809,N_18475,N_18271);
or U19810 (N_19810,N_18528,N_18355);
nand U19811 (N_19811,N_18506,N_18928);
or U19812 (N_19812,N_18088,N_18090);
nand U19813 (N_19813,N_18770,N_18603);
or U19814 (N_19814,N_18214,N_18726);
nand U19815 (N_19815,N_18533,N_18542);
nand U19816 (N_19816,N_18427,N_18100);
nand U19817 (N_19817,N_18776,N_18312);
nor U19818 (N_19818,N_18559,N_18387);
nand U19819 (N_19819,N_18790,N_18248);
or U19820 (N_19820,N_18171,N_18734);
or U19821 (N_19821,N_18961,N_18195);
and U19822 (N_19822,N_18949,N_18137);
or U19823 (N_19823,N_18389,N_18738);
and U19824 (N_19824,N_18202,N_18352);
nor U19825 (N_19825,N_18070,N_18781);
nand U19826 (N_19826,N_18148,N_18499);
or U19827 (N_19827,N_18415,N_18186);
nor U19828 (N_19828,N_18498,N_18373);
nor U19829 (N_19829,N_18076,N_18796);
nand U19830 (N_19830,N_18839,N_18606);
and U19831 (N_19831,N_18818,N_18367);
or U19832 (N_19832,N_18455,N_18613);
xor U19833 (N_19833,N_18204,N_18366);
nor U19834 (N_19834,N_18129,N_18383);
and U19835 (N_19835,N_18134,N_18625);
or U19836 (N_19836,N_18766,N_18167);
or U19837 (N_19837,N_18474,N_18494);
or U19838 (N_19838,N_18517,N_18091);
and U19839 (N_19839,N_18883,N_18097);
nor U19840 (N_19840,N_18670,N_18500);
and U19841 (N_19841,N_18500,N_18518);
and U19842 (N_19842,N_18916,N_18304);
nor U19843 (N_19843,N_18153,N_18732);
nand U19844 (N_19844,N_18223,N_18094);
nand U19845 (N_19845,N_18337,N_18462);
or U19846 (N_19846,N_18449,N_18932);
nand U19847 (N_19847,N_18762,N_18995);
or U19848 (N_19848,N_18823,N_18437);
or U19849 (N_19849,N_18779,N_18038);
nand U19850 (N_19850,N_18287,N_18298);
or U19851 (N_19851,N_18488,N_18881);
nor U19852 (N_19852,N_18265,N_18651);
nor U19853 (N_19853,N_18824,N_18865);
xnor U19854 (N_19854,N_18791,N_18870);
or U19855 (N_19855,N_18690,N_18583);
or U19856 (N_19856,N_18705,N_18718);
nand U19857 (N_19857,N_18219,N_18122);
xor U19858 (N_19858,N_18464,N_18143);
or U19859 (N_19859,N_18529,N_18631);
nand U19860 (N_19860,N_18414,N_18888);
and U19861 (N_19861,N_18888,N_18961);
and U19862 (N_19862,N_18952,N_18079);
nand U19863 (N_19863,N_18468,N_18425);
and U19864 (N_19864,N_18079,N_18764);
or U19865 (N_19865,N_18403,N_18894);
or U19866 (N_19866,N_18783,N_18716);
xor U19867 (N_19867,N_18238,N_18351);
and U19868 (N_19868,N_18163,N_18064);
nor U19869 (N_19869,N_18354,N_18090);
and U19870 (N_19870,N_18979,N_18390);
xor U19871 (N_19871,N_18986,N_18776);
and U19872 (N_19872,N_18212,N_18588);
and U19873 (N_19873,N_18078,N_18733);
and U19874 (N_19874,N_18186,N_18070);
and U19875 (N_19875,N_18703,N_18645);
xor U19876 (N_19876,N_18648,N_18161);
or U19877 (N_19877,N_18301,N_18774);
nand U19878 (N_19878,N_18165,N_18094);
xor U19879 (N_19879,N_18422,N_18183);
nor U19880 (N_19880,N_18937,N_18016);
nand U19881 (N_19881,N_18067,N_18744);
and U19882 (N_19882,N_18955,N_18671);
or U19883 (N_19883,N_18271,N_18688);
nand U19884 (N_19884,N_18819,N_18005);
or U19885 (N_19885,N_18467,N_18610);
nand U19886 (N_19886,N_18645,N_18186);
xor U19887 (N_19887,N_18503,N_18982);
and U19888 (N_19888,N_18270,N_18039);
or U19889 (N_19889,N_18298,N_18002);
and U19890 (N_19890,N_18692,N_18024);
nand U19891 (N_19891,N_18454,N_18190);
xor U19892 (N_19892,N_18915,N_18386);
nand U19893 (N_19893,N_18754,N_18338);
xnor U19894 (N_19894,N_18497,N_18615);
nor U19895 (N_19895,N_18911,N_18074);
xnor U19896 (N_19896,N_18359,N_18558);
or U19897 (N_19897,N_18419,N_18623);
or U19898 (N_19898,N_18360,N_18476);
and U19899 (N_19899,N_18984,N_18992);
nor U19900 (N_19900,N_18393,N_18732);
or U19901 (N_19901,N_18019,N_18226);
and U19902 (N_19902,N_18574,N_18710);
or U19903 (N_19903,N_18808,N_18691);
nand U19904 (N_19904,N_18418,N_18789);
or U19905 (N_19905,N_18215,N_18175);
nand U19906 (N_19906,N_18636,N_18500);
and U19907 (N_19907,N_18638,N_18075);
nand U19908 (N_19908,N_18425,N_18820);
nand U19909 (N_19909,N_18366,N_18107);
nand U19910 (N_19910,N_18118,N_18532);
and U19911 (N_19911,N_18765,N_18625);
nand U19912 (N_19912,N_18384,N_18057);
xor U19913 (N_19913,N_18638,N_18690);
or U19914 (N_19914,N_18140,N_18275);
nand U19915 (N_19915,N_18923,N_18090);
or U19916 (N_19916,N_18378,N_18145);
nand U19917 (N_19917,N_18412,N_18158);
and U19918 (N_19918,N_18685,N_18987);
nor U19919 (N_19919,N_18826,N_18818);
and U19920 (N_19920,N_18868,N_18961);
or U19921 (N_19921,N_18585,N_18032);
nand U19922 (N_19922,N_18133,N_18577);
nor U19923 (N_19923,N_18033,N_18762);
xor U19924 (N_19924,N_18721,N_18242);
nand U19925 (N_19925,N_18191,N_18097);
xor U19926 (N_19926,N_18153,N_18792);
nor U19927 (N_19927,N_18556,N_18133);
and U19928 (N_19928,N_18271,N_18539);
or U19929 (N_19929,N_18863,N_18124);
nand U19930 (N_19930,N_18887,N_18932);
nand U19931 (N_19931,N_18615,N_18438);
or U19932 (N_19932,N_18855,N_18703);
nor U19933 (N_19933,N_18248,N_18169);
nor U19934 (N_19934,N_18931,N_18616);
or U19935 (N_19935,N_18011,N_18190);
and U19936 (N_19936,N_18354,N_18514);
xor U19937 (N_19937,N_18737,N_18057);
nor U19938 (N_19938,N_18889,N_18654);
nand U19939 (N_19939,N_18292,N_18744);
or U19940 (N_19940,N_18803,N_18415);
and U19941 (N_19941,N_18963,N_18280);
nor U19942 (N_19942,N_18631,N_18287);
xor U19943 (N_19943,N_18635,N_18885);
nor U19944 (N_19944,N_18564,N_18600);
and U19945 (N_19945,N_18229,N_18294);
xnor U19946 (N_19946,N_18072,N_18883);
xnor U19947 (N_19947,N_18907,N_18039);
nor U19948 (N_19948,N_18749,N_18232);
and U19949 (N_19949,N_18495,N_18522);
and U19950 (N_19950,N_18281,N_18437);
nand U19951 (N_19951,N_18085,N_18265);
or U19952 (N_19952,N_18918,N_18053);
xor U19953 (N_19953,N_18339,N_18314);
nand U19954 (N_19954,N_18657,N_18134);
and U19955 (N_19955,N_18085,N_18558);
or U19956 (N_19956,N_18737,N_18287);
nor U19957 (N_19957,N_18377,N_18492);
or U19958 (N_19958,N_18305,N_18786);
nor U19959 (N_19959,N_18162,N_18323);
xor U19960 (N_19960,N_18243,N_18094);
nor U19961 (N_19961,N_18182,N_18524);
xor U19962 (N_19962,N_18863,N_18211);
and U19963 (N_19963,N_18057,N_18026);
and U19964 (N_19964,N_18061,N_18317);
and U19965 (N_19965,N_18895,N_18056);
xor U19966 (N_19966,N_18669,N_18540);
nor U19967 (N_19967,N_18250,N_18405);
or U19968 (N_19968,N_18258,N_18073);
or U19969 (N_19969,N_18318,N_18072);
nand U19970 (N_19970,N_18008,N_18061);
xnor U19971 (N_19971,N_18767,N_18519);
and U19972 (N_19972,N_18234,N_18265);
nand U19973 (N_19973,N_18162,N_18952);
or U19974 (N_19974,N_18511,N_18350);
and U19975 (N_19975,N_18677,N_18699);
and U19976 (N_19976,N_18842,N_18072);
xor U19977 (N_19977,N_18722,N_18418);
or U19978 (N_19978,N_18071,N_18125);
xor U19979 (N_19979,N_18077,N_18071);
nor U19980 (N_19980,N_18343,N_18312);
and U19981 (N_19981,N_18489,N_18304);
nand U19982 (N_19982,N_18485,N_18337);
xnor U19983 (N_19983,N_18552,N_18210);
nor U19984 (N_19984,N_18804,N_18584);
xor U19985 (N_19985,N_18320,N_18962);
nor U19986 (N_19986,N_18076,N_18371);
nor U19987 (N_19987,N_18028,N_18930);
nor U19988 (N_19988,N_18391,N_18703);
nand U19989 (N_19989,N_18744,N_18433);
nor U19990 (N_19990,N_18426,N_18034);
nor U19991 (N_19991,N_18760,N_18183);
nand U19992 (N_19992,N_18890,N_18305);
xnor U19993 (N_19993,N_18239,N_18824);
or U19994 (N_19994,N_18961,N_18925);
xnor U19995 (N_19995,N_18322,N_18581);
nand U19996 (N_19996,N_18123,N_18145);
and U19997 (N_19997,N_18771,N_18609);
nor U19998 (N_19998,N_18143,N_18530);
nor U19999 (N_19999,N_18457,N_18353);
or U20000 (N_20000,N_19996,N_19403);
or U20001 (N_20001,N_19451,N_19689);
nand U20002 (N_20002,N_19673,N_19933);
xor U20003 (N_20003,N_19106,N_19148);
or U20004 (N_20004,N_19310,N_19138);
and U20005 (N_20005,N_19616,N_19128);
xor U20006 (N_20006,N_19150,N_19027);
and U20007 (N_20007,N_19255,N_19232);
nand U20008 (N_20008,N_19376,N_19246);
nor U20009 (N_20009,N_19647,N_19769);
or U20010 (N_20010,N_19773,N_19591);
nand U20011 (N_20011,N_19974,N_19176);
nand U20012 (N_20012,N_19558,N_19428);
and U20013 (N_20013,N_19546,N_19781);
nor U20014 (N_20014,N_19320,N_19585);
xor U20015 (N_20015,N_19044,N_19434);
nand U20016 (N_20016,N_19874,N_19031);
nor U20017 (N_20017,N_19118,N_19992);
and U20018 (N_20018,N_19482,N_19500);
or U20019 (N_20019,N_19812,N_19542);
nand U20020 (N_20020,N_19249,N_19790);
xor U20021 (N_20021,N_19340,N_19761);
xnor U20022 (N_20022,N_19530,N_19317);
xor U20023 (N_20023,N_19184,N_19486);
nor U20024 (N_20024,N_19254,N_19532);
and U20025 (N_20025,N_19337,N_19909);
nand U20026 (N_20026,N_19960,N_19285);
and U20027 (N_20027,N_19348,N_19124);
nor U20028 (N_20028,N_19405,N_19086);
nand U20029 (N_20029,N_19439,N_19935);
xnor U20030 (N_20030,N_19401,N_19608);
nand U20031 (N_20031,N_19997,N_19971);
nor U20032 (N_20032,N_19149,N_19518);
or U20033 (N_20033,N_19798,N_19905);
nor U20034 (N_20034,N_19442,N_19090);
nor U20035 (N_20035,N_19868,N_19737);
xnor U20036 (N_20036,N_19575,N_19201);
nand U20037 (N_20037,N_19295,N_19490);
nor U20038 (N_20038,N_19160,N_19768);
or U20039 (N_20039,N_19314,N_19488);
and U20040 (N_20040,N_19228,N_19889);
nand U20041 (N_20041,N_19586,N_19869);
nor U20042 (N_20042,N_19634,N_19598);
and U20043 (N_20043,N_19480,N_19389);
nand U20044 (N_20044,N_19876,N_19822);
nor U20045 (N_20045,N_19948,N_19025);
xnor U20046 (N_20046,N_19928,N_19499);
and U20047 (N_20047,N_19601,N_19067);
nor U20048 (N_20048,N_19581,N_19239);
nand U20049 (N_20049,N_19029,N_19925);
nor U20050 (N_20050,N_19719,N_19803);
nor U20051 (N_20051,N_19549,N_19977);
nand U20052 (N_20052,N_19022,N_19702);
and U20053 (N_20053,N_19784,N_19704);
xor U20054 (N_20054,N_19955,N_19521);
xnor U20055 (N_20055,N_19949,N_19155);
nand U20056 (N_20056,N_19056,N_19919);
and U20057 (N_20057,N_19849,N_19355);
xor U20058 (N_20058,N_19195,N_19567);
and U20059 (N_20059,N_19672,N_19087);
xnor U20060 (N_20060,N_19547,N_19880);
xor U20061 (N_20061,N_19233,N_19237);
xnor U20062 (N_20062,N_19194,N_19535);
xor U20063 (N_20063,N_19093,N_19374);
xnor U20064 (N_20064,N_19271,N_19460);
xnor U20065 (N_20065,N_19989,N_19832);
or U20066 (N_20066,N_19637,N_19133);
or U20067 (N_20067,N_19158,N_19402);
nand U20068 (N_20068,N_19851,N_19709);
nand U20069 (N_20069,N_19918,N_19892);
xor U20070 (N_20070,N_19074,N_19648);
and U20071 (N_20071,N_19189,N_19288);
xnor U20072 (N_20072,N_19198,N_19857);
xnor U20073 (N_20073,N_19813,N_19409);
or U20074 (N_20074,N_19009,N_19041);
xnor U20075 (N_20075,N_19404,N_19908);
and U20076 (N_20076,N_19145,N_19595);
xor U20077 (N_20077,N_19384,N_19491);
and U20078 (N_20078,N_19913,N_19131);
nand U20079 (N_20079,N_19327,N_19760);
or U20080 (N_20080,N_19720,N_19881);
xor U20081 (N_20081,N_19536,N_19639);
xor U20082 (N_20082,N_19185,N_19339);
or U20083 (N_20083,N_19004,N_19628);
xor U20084 (N_20084,N_19723,N_19831);
and U20085 (N_20085,N_19520,N_19212);
xnor U20086 (N_20086,N_19659,N_19561);
and U20087 (N_20087,N_19724,N_19739);
and U20088 (N_20088,N_19306,N_19219);
xnor U20089 (N_20089,N_19510,N_19522);
nand U20090 (N_20090,N_19268,N_19619);
nand U20091 (N_20091,N_19296,N_19172);
nand U20092 (N_20092,N_19018,N_19292);
nand U20093 (N_20093,N_19042,N_19627);
nor U20094 (N_20094,N_19240,N_19431);
nor U20095 (N_20095,N_19414,N_19688);
or U20096 (N_20096,N_19101,N_19350);
xor U20097 (N_20097,N_19003,N_19772);
or U20098 (N_20098,N_19531,N_19111);
nand U20099 (N_20099,N_19280,N_19452);
or U20100 (N_20100,N_19386,N_19808);
or U20101 (N_20101,N_19721,N_19293);
xnor U20102 (N_20102,N_19728,N_19511);
nor U20103 (N_20103,N_19926,N_19583);
nor U20104 (N_20104,N_19795,N_19275);
nand U20105 (N_20105,N_19024,N_19085);
and U20106 (N_20106,N_19330,N_19000);
and U20107 (N_20107,N_19694,N_19940);
nand U20108 (N_20108,N_19433,N_19710);
nand U20109 (N_20109,N_19590,N_19048);
and U20110 (N_20110,N_19907,N_19517);
and U20111 (N_20111,N_19764,N_19824);
xnor U20112 (N_20112,N_19171,N_19814);
xnor U20113 (N_20113,N_19801,N_19424);
xor U20114 (N_20114,N_19380,N_19045);
xor U20115 (N_20115,N_19653,N_19816);
nand U20116 (N_20116,N_19842,N_19277);
and U20117 (N_20117,N_19221,N_19756);
nor U20118 (N_20118,N_19623,N_19612);
nor U20119 (N_20119,N_19200,N_19286);
xor U20120 (N_20120,N_19323,N_19478);
and U20121 (N_20121,N_19758,N_19708);
xor U20122 (N_20122,N_19463,N_19065);
nand U20123 (N_20123,N_19611,N_19958);
or U20124 (N_20124,N_19733,N_19844);
xor U20125 (N_20125,N_19743,N_19416);
or U20126 (N_20126,N_19750,N_19862);
and U20127 (N_20127,N_19931,N_19788);
nor U20128 (N_20128,N_19257,N_19712);
xnor U20129 (N_20129,N_19779,N_19622);
xor U20130 (N_20130,N_19533,N_19089);
and U20131 (N_20131,N_19305,N_19109);
or U20132 (N_20132,N_19968,N_19923);
and U20133 (N_20133,N_19006,N_19661);
and U20134 (N_20134,N_19979,N_19599);
nand U20135 (N_20135,N_19407,N_19910);
xnor U20136 (N_20136,N_19061,N_19765);
and U20137 (N_20137,N_19924,N_19013);
or U20138 (N_20138,N_19681,N_19358);
nand U20139 (N_20139,N_19047,N_19963);
xnor U20140 (N_20140,N_19256,N_19572);
nor U20141 (N_20141,N_19058,N_19283);
and U20142 (N_20142,N_19193,N_19556);
nor U20143 (N_20143,N_19092,N_19726);
or U20144 (N_20144,N_19438,N_19731);
or U20145 (N_20145,N_19231,N_19853);
xor U20146 (N_20146,N_19315,N_19130);
or U20147 (N_20147,N_19199,N_19566);
nor U20148 (N_20148,N_19263,N_19369);
or U20149 (N_20149,N_19357,N_19961);
or U20150 (N_20150,N_19422,N_19064);
nand U20151 (N_20151,N_19338,N_19105);
nand U20152 (N_20152,N_19662,N_19457);
nand U20153 (N_20153,N_19748,N_19021);
or U20154 (N_20154,N_19367,N_19359);
or U20155 (N_20155,N_19860,N_19259);
nor U20156 (N_20156,N_19046,N_19649);
xor U20157 (N_20157,N_19843,N_19353);
nand U20158 (N_20158,N_19643,N_19505);
or U20159 (N_20159,N_19495,N_19448);
or U20160 (N_20160,N_19493,N_19373);
or U20161 (N_20161,N_19346,N_19698);
and U20162 (N_20162,N_19445,N_19341);
nor U20163 (N_20163,N_19391,N_19734);
and U20164 (N_20164,N_19551,N_19845);
and U20165 (N_20165,N_19620,N_19605);
nand U20166 (N_20166,N_19941,N_19774);
xnor U20167 (N_20167,N_19534,N_19169);
nor U20168 (N_20168,N_19883,N_19069);
and U20169 (N_20169,N_19217,N_19936);
xnor U20170 (N_20170,N_19991,N_19426);
and U20171 (N_20171,N_19902,N_19137);
nand U20172 (N_20172,N_19134,N_19570);
and U20173 (N_20173,N_19797,N_19618);
nand U20174 (N_20174,N_19363,N_19251);
or U20175 (N_20175,N_19789,N_19475);
and U20176 (N_20176,N_19055,N_19771);
nor U20177 (N_20177,N_19864,N_19565);
nor U20178 (N_20178,N_19423,N_19002);
and U20179 (N_20179,N_19554,N_19421);
and U20180 (N_20180,N_19226,N_19371);
and U20181 (N_20181,N_19379,N_19569);
xor U20182 (N_20182,N_19509,N_19210);
nand U20183 (N_20183,N_19593,N_19957);
or U20184 (N_20184,N_19103,N_19287);
or U20185 (N_20185,N_19494,N_19446);
or U20186 (N_20186,N_19316,N_19332);
nor U20187 (N_20187,N_19334,N_19023);
nor U20188 (N_20188,N_19990,N_19609);
nand U20189 (N_20189,N_19512,N_19664);
nand U20190 (N_20190,N_19929,N_19372);
nand U20191 (N_20191,N_19506,N_19076);
or U20192 (N_20192,N_19098,N_19785);
or U20193 (N_20193,N_19245,N_19584);
xnor U20194 (N_20194,N_19691,N_19040);
and U20195 (N_20195,N_19717,N_19787);
nor U20196 (N_20196,N_19944,N_19415);
xor U20197 (N_20197,N_19081,N_19904);
nor U20198 (N_20198,N_19998,N_19050);
nor U20199 (N_20199,N_19806,N_19250);
and U20200 (N_20200,N_19385,N_19008);
xnor U20201 (N_20201,N_19825,N_19587);
and U20202 (N_20202,N_19906,N_19888);
xnor U20203 (N_20203,N_19410,N_19035);
and U20204 (N_20204,N_19633,N_19886);
nand U20205 (N_20205,N_19503,N_19163);
and U20206 (N_20206,N_19519,N_19294);
and U20207 (N_20207,N_19266,N_19577);
and U20208 (N_20208,N_19950,N_19981);
xor U20209 (N_20209,N_19984,N_19011);
or U20210 (N_20210,N_19846,N_19701);
xor U20211 (N_20211,N_19388,N_19303);
nand U20212 (N_20212,N_19793,N_19987);
and U20213 (N_20213,N_19747,N_19485);
and U20214 (N_20214,N_19670,N_19225);
xnor U20215 (N_20215,N_19810,N_19516);
and U20216 (N_20216,N_19252,N_19878);
xor U20217 (N_20217,N_19147,N_19791);
xor U20218 (N_20218,N_19555,N_19140);
and U20219 (N_20219,N_19032,N_19687);
or U20220 (N_20220,N_19262,N_19049);
and U20221 (N_20221,N_19063,N_19121);
and U20222 (N_20222,N_19364,N_19139);
or U20223 (N_20223,N_19260,N_19328);
xnor U20224 (N_20224,N_19443,N_19116);
nor U20225 (N_20225,N_19986,N_19600);
or U20226 (N_20226,N_19677,N_19311);
or U20227 (N_20227,N_19084,N_19711);
and U20228 (N_20228,N_19079,N_19776);
nand U20229 (N_20229,N_19153,N_19216);
or U20230 (N_20230,N_19453,N_19967);
xor U20231 (N_20231,N_19281,N_19783);
or U20232 (N_20232,N_19538,N_19994);
or U20233 (N_20233,N_19807,N_19412);
or U20234 (N_20234,N_19576,N_19613);
xor U20235 (N_20235,N_19663,N_19496);
nand U20236 (N_20236,N_19930,N_19545);
nor U20237 (N_20237,N_19178,N_19307);
nand U20238 (N_20238,N_19333,N_19143);
nor U20239 (N_20239,N_19875,N_19912);
nor U20240 (N_20240,N_19449,N_19560);
nor U20241 (N_20241,N_19274,N_19916);
nor U20242 (N_20242,N_19901,N_19191);
nand U20243 (N_20243,N_19658,N_19954);
xor U20244 (N_20244,N_19513,N_19073);
nor U20245 (N_20245,N_19757,N_19548);
xor U20246 (N_20246,N_19070,N_19222);
or U20247 (N_20247,N_19982,N_19181);
nor U20248 (N_20248,N_19528,N_19945);
nor U20249 (N_20249,N_19615,N_19834);
or U20250 (N_20250,N_19804,N_19033);
nand U20251 (N_20251,N_19999,N_19179);
and U20252 (N_20252,N_19345,N_19652);
nand U20253 (N_20253,N_19173,N_19123);
or U20254 (N_20254,N_19447,N_19094);
nor U20255 (N_20255,N_19368,N_19187);
xor U20256 (N_20256,N_19470,N_19165);
and U20257 (N_20257,N_19951,N_19174);
and U20258 (N_20258,N_19541,N_19156);
nor U20259 (N_20259,N_19436,N_19248);
or U20260 (N_20260,N_19362,N_19291);
and U20261 (N_20261,N_19976,N_19895);
or U20262 (N_20262,N_19015,N_19716);
nand U20263 (N_20263,N_19767,N_19937);
nor U20264 (N_20264,N_19408,N_19243);
and U20265 (N_20265,N_19324,N_19484);
nor U20266 (N_20266,N_19899,N_19749);
or U20267 (N_20267,N_19543,N_19224);
and U20268 (N_20268,N_19437,N_19683);
nor U20269 (N_20269,N_19614,N_19481);
and U20270 (N_20270,N_19943,N_19603);
and U20271 (N_20271,N_19039,N_19780);
and U20272 (N_20272,N_19430,N_19034);
xnor U20273 (N_20273,N_19863,N_19927);
nor U20274 (N_20274,N_19290,N_19188);
nand U20275 (N_20275,N_19953,N_19030);
or U20276 (N_20276,N_19152,N_19043);
xnor U20277 (N_20277,N_19016,N_19877);
xor U20278 (N_20278,N_19596,N_19539);
nand U20279 (N_20279,N_19196,N_19469);
and U20280 (N_20280,N_19299,N_19885);
xnor U20281 (N_20281,N_19269,N_19696);
nor U20282 (N_20282,N_19301,N_19066);
xnor U20283 (N_20283,N_19730,N_19829);
and U20284 (N_20284,N_19455,N_19329);
nor U20285 (N_20285,N_19411,N_19762);
and U20286 (N_20286,N_19037,N_19164);
or U20287 (N_20287,N_19568,N_19897);
or U20288 (N_20288,N_19308,N_19597);
xor U20289 (N_20289,N_19208,N_19479);
or U20290 (N_20290,N_19223,N_19456);
nand U20291 (N_20291,N_19830,N_19477);
nand U20292 (N_20292,N_19592,N_19969);
nor U20293 (N_20293,N_19235,N_19242);
and U20294 (N_20294,N_19778,N_19141);
xor U20295 (N_20295,N_19057,N_19529);
and U20296 (N_20296,N_19203,N_19154);
nor U20297 (N_20297,N_19466,N_19001);
nand U20298 (N_20298,N_19993,N_19766);
nand U20299 (N_20299,N_19309,N_19903);
and U20300 (N_20300,N_19390,N_19417);
or U20301 (N_20301,N_19071,N_19082);
nand U20302 (N_20302,N_19896,N_19966);
nor U20303 (N_20303,N_19738,N_19640);
and U20304 (N_20304,N_19450,N_19604);
or U20305 (N_20305,N_19646,N_19523);
nand U20306 (N_20306,N_19080,N_19722);
and U20307 (N_20307,N_19365,N_19751);
xnor U20308 (N_20308,N_19489,N_19630);
nand U20309 (N_20309,N_19244,N_19097);
xor U20310 (N_20310,N_19238,N_19840);
and U20311 (N_20311,N_19939,N_19159);
nor U20312 (N_20312,N_19665,N_19632);
or U20313 (N_20313,N_19911,N_19852);
nor U20314 (N_20314,N_19441,N_19938);
nor U20315 (N_20315,N_19763,N_19192);
or U20316 (N_20316,N_19809,N_19799);
xor U20317 (N_20317,N_19859,N_19686);
xnor U20318 (N_20318,N_19186,N_19406);
nor U20319 (N_20319,N_19675,N_19054);
nor U20320 (N_20320,N_19395,N_19125);
and U20321 (N_20321,N_19959,N_19206);
nor U20322 (N_20322,N_19866,N_19841);
nor U20323 (N_20323,N_19072,N_19302);
or U20324 (N_20324,N_19474,N_19356);
or U20325 (N_20325,N_19427,N_19468);
nor U20326 (N_20326,N_19934,N_19377);
nand U20327 (N_20327,N_19017,N_19920);
nor U20328 (N_20328,N_19947,N_19540);
nor U20329 (N_20329,N_19654,N_19435);
or U20330 (N_20330,N_19537,N_19102);
nor U20331 (N_20331,N_19697,N_19626);
or U20332 (N_20332,N_19322,N_19679);
or U20333 (N_20333,N_19168,N_19343);
or U20334 (N_20334,N_19873,N_19279);
xnor U20335 (N_20335,N_19083,N_19588);
or U20336 (N_20336,N_19582,N_19100);
nand U20337 (N_20337,N_19745,N_19476);
xor U20338 (N_20338,N_19805,N_19775);
xnor U20339 (N_20339,N_19180,N_19400);
nor U20340 (N_20340,N_19879,N_19398);
nand U20341 (N_20341,N_19349,N_19800);
nor U20342 (N_20342,N_19113,N_19606);
or U20343 (N_20343,N_19336,N_19059);
nor U20344 (N_20344,N_19062,N_19504);
nand U20345 (N_20345,N_19574,N_19419);
or U20346 (N_20346,N_19051,N_19796);
or U20347 (N_20347,N_19454,N_19444);
or U20348 (N_20348,N_19550,N_19669);
xnor U20349 (N_20349,N_19366,N_19276);
nor U20350 (N_20350,N_19744,N_19264);
nand U20351 (N_20351,N_19360,N_19965);
nand U20352 (N_20352,N_19091,N_19674);
or U20353 (N_20353,N_19382,N_19387);
nand U20354 (N_20354,N_19273,N_19028);
nor U20355 (N_20355,N_19972,N_19706);
and U20356 (N_20356,N_19397,N_19502);
xnor U20357 (N_20357,N_19827,N_19699);
nor U20358 (N_20358,N_19732,N_19882);
or U20359 (N_20359,N_19132,N_19508);
and U20360 (N_20360,N_19942,N_19641);
nand U20361 (N_20361,N_19607,N_19298);
nor U20362 (N_20362,N_19352,N_19236);
and U20363 (N_20363,N_19891,N_19564);
xnor U20364 (N_20364,N_19563,N_19300);
or U20365 (N_20365,N_19399,N_19755);
or U20366 (N_20366,N_19684,N_19229);
nand U20367 (N_20367,N_19770,N_19112);
nand U20368 (N_20368,N_19552,N_19392);
or U20369 (N_20369,N_19854,N_19167);
nand U20370 (N_20370,N_19202,N_19837);
nand U20371 (N_20371,N_19425,N_19847);
or U20372 (N_20372,N_19660,N_19644);
nor U20373 (N_20373,N_19282,N_19802);
or U20374 (N_20374,N_19197,N_19289);
or U20375 (N_20375,N_19157,N_19492);
nor U20376 (N_20376,N_19828,N_19700);
xnor U20377 (N_20377,N_19507,N_19170);
nand U20378 (N_20378,N_19209,N_19635);
xnor U20379 (N_20379,N_19230,N_19331);
xor U20380 (N_20380,N_19676,N_19715);
or U20381 (N_20381,N_19515,N_19514);
xor U20382 (N_20382,N_19735,N_19284);
xnor U20383 (N_20383,N_19759,N_19861);
and U20384 (N_20384,N_19135,N_19685);
xnor U20385 (N_20385,N_19690,N_19151);
nand U20386 (N_20386,N_19978,N_19321);
or U20387 (N_20387,N_19884,N_19497);
xnor U20388 (N_20388,N_19077,N_19241);
and U20389 (N_20389,N_19746,N_19175);
and U20390 (N_20390,N_19740,N_19319);
and U20391 (N_20391,N_19544,N_19890);
nor U20392 (N_20392,N_19114,N_19579);
or U20393 (N_20393,N_19562,N_19394);
nor U20394 (N_20394,N_19819,N_19465);
xor U20395 (N_20395,N_19777,N_19095);
and U20396 (N_20396,N_19573,N_19893);
xor U20397 (N_20397,N_19161,N_19019);
xnor U20398 (N_20398,N_19326,N_19190);
nand U20399 (N_20399,N_19432,N_19858);
nand U20400 (N_20400,N_19347,N_19127);
and U20401 (N_20401,N_19975,N_19278);
and U20402 (N_20402,N_19820,N_19312);
nand U20403 (N_20403,N_19741,N_19848);
nand U20404 (N_20404,N_19638,N_19458);
nor U20405 (N_20405,N_19099,N_19162);
xor U20406 (N_20406,N_19970,N_19014);
or U20407 (N_20407,N_19693,N_19247);
nand U20408 (N_20408,N_19713,N_19578);
or U20409 (N_20409,N_19088,N_19526);
or U20410 (N_20410,N_19459,N_19297);
and U20411 (N_20411,N_19815,N_19678);
or U20412 (N_20412,N_19318,N_19917);
or U20413 (N_20413,N_19383,N_19115);
xnor U20414 (N_20414,N_19182,N_19351);
xnor U20415 (N_20415,N_19007,N_19211);
or U20416 (N_20416,N_19833,N_19922);
nand U20417 (N_20417,N_19214,N_19117);
nor U20418 (N_20418,N_19651,N_19396);
nor U20419 (N_20419,N_19786,N_19354);
and U20420 (N_20420,N_19501,N_19462);
nor U20421 (N_20421,N_19119,N_19393);
nand U20422 (N_20422,N_19122,N_19887);
or U20423 (N_20423,N_19218,N_19375);
and U20424 (N_20424,N_19036,N_19220);
xnor U20425 (N_20425,N_19205,N_19078);
nor U20426 (N_20426,N_19811,N_19068);
nand U20427 (N_20427,N_19335,N_19718);
xnor U20428 (N_20428,N_19108,N_19177);
xor U20429 (N_20429,N_19666,N_19253);
or U20430 (N_20430,N_19782,N_19729);
nor U20431 (N_20431,N_19855,N_19826);
or U20432 (N_20432,N_19580,N_19915);
nor U20433 (N_20433,N_19429,N_19342);
nand U20434 (N_20434,N_19136,N_19703);
nor U20435 (N_20435,N_19752,N_19836);
nor U20436 (N_20436,N_19483,N_19026);
or U20437 (N_20437,N_19707,N_19727);
nor U20438 (N_20438,N_19525,N_19589);
or U20439 (N_20439,N_19557,N_19107);
and U20440 (N_20440,N_19120,N_19461);
and U20441 (N_20441,N_19642,N_19617);
xor U20442 (N_20442,N_19129,N_19370);
xnor U20443 (N_20443,N_19872,N_19440);
and U20444 (N_20444,N_19420,N_19973);
nand U20445 (N_20445,N_19818,N_19553);
or U20446 (N_20446,N_19012,N_19344);
or U20447 (N_20447,N_19020,N_19667);
xnor U20448 (N_20448,N_19656,N_19418);
or U20449 (N_20449,N_19010,N_19571);
nand U20450 (N_20450,N_19900,N_19980);
and U20451 (N_20451,N_19473,N_19261);
or U20452 (N_20452,N_19625,N_19962);
or U20453 (N_20453,N_19668,N_19856);
nor U20454 (N_20454,N_19821,N_19624);
xnor U20455 (N_20455,N_19714,N_19464);
or U20456 (N_20456,N_19267,N_19995);
nor U20457 (N_20457,N_19524,N_19472);
or U20458 (N_20458,N_19142,N_19964);
nand U20459 (N_20459,N_19817,N_19682);
nand U20460 (N_20460,N_19655,N_19467);
or U20461 (N_20461,N_19629,N_19794);
nand U20462 (N_20462,N_19838,N_19610);
nand U20463 (N_20463,N_19498,N_19754);
or U20464 (N_20464,N_19823,N_19792);
and U20465 (N_20465,N_19126,N_19657);
and U20466 (N_20466,N_19146,N_19932);
or U20467 (N_20467,N_19870,N_19894);
or U20468 (N_20468,N_19038,N_19594);
or U20469 (N_20469,N_19207,N_19487);
nor U20470 (N_20470,N_19183,N_19645);
xnor U20471 (N_20471,N_19075,N_19096);
and U20472 (N_20472,N_19871,N_19680);
or U20473 (N_20473,N_19952,N_19914);
or U20474 (N_20474,N_19104,N_19985);
xnor U20475 (N_20475,N_19956,N_19234);
nand U20476 (N_20476,N_19378,N_19867);
and U20477 (N_20477,N_19060,N_19695);
or U20478 (N_20478,N_19053,N_19413);
and U20479 (N_20479,N_19272,N_19650);
nor U20480 (N_20480,N_19742,N_19636);
and U20481 (N_20481,N_19602,N_19144);
nand U20482 (N_20482,N_19381,N_19736);
xor U20483 (N_20483,N_19705,N_19946);
and U20484 (N_20484,N_19983,N_19270);
xnor U20485 (N_20485,N_19621,N_19527);
xnor U20486 (N_20486,N_19753,N_19361);
nor U20487 (N_20487,N_19839,N_19671);
nand U20488 (N_20488,N_19304,N_19631);
xnor U20489 (N_20489,N_19988,N_19835);
xor U20490 (N_20490,N_19265,N_19215);
nand U20491 (N_20491,N_19052,N_19559);
nand U20492 (N_20492,N_19213,N_19204);
nor U20493 (N_20493,N_19313,N_19725);
nor U20494 (N_20494,N_19325,N_19166);
nand U20495 (N_20495,N_19005,N_19850);
and U20496 (N_20496,N_19692,N_19258);
or U20497 (N_20497,N_19110,N_19471);
xor U20498 (N_20498,N_19921,N_19865);
xnor U20499 (N_20499,N_19898,N_19227);
xnor U20500 (N_20500,N_19400,N_19233);
nand U20501 (N_20501,N_19446,N_19295);
xnor U20502 (N_20502,N_19078,N_19083);
nand U20503 (N_20503,N_19199,N_19379);
or U20504 (N_20504,N_19781,N_19453);
and U20505 (N_20505,N_19166,N_19270);
and U20506 (N_20506,N_19359,N_19018);
or U20507 (N_20507,N_19370,N_19883);
or U20508 (N_20508,N_19809,N_19431);
or U20509 (N_20509,N_19244,N_19994);
xnor U20510 (N_20510,N_19821,N_19595);
or U20511 (N_20511,N_19398,N_19575);
xor U20512 (N_20512,N_19395,N_19249);
nand U20513 (N_20513,N_19480,N_19003);
nand U20514 (N_20514,N_19886,N_19231);
nand U20515 (N_20515,N_19685,N_19725);
or U20516 (N_20516,N_19131,N_19435);
xnor U20517 (N_20517,N_19116,N_19263);
nand U20518 (N_20518,N_19590,N_19483);
nor U20519 (N_20519,N_19771,N_19981);
nand U20520 (N_20520,N_19086,N_19554);
nand U20521 (N_20521,N_19051,N_19492);
or U20522 (N_20522,N_19438,N_19234);
xor U20523 (N_20523,N_19150,N_19546);
nor U20524 (N_20524,N_19691,N_19048);
nor U20525 (N_20525,N_19649,N_19481);
or U20526 (N_20526,N_19000,N_19495);
xor U20527 (N_20527,N_19228,N_19813);
nor U20528 (N_20528,N_19993,N_19055);
nand U20529 (N_20529,N_19528,N_19960);
nand U20530 (N_20530,N_19382,N_19222);
nand U20531 (N_20531,N_19735,N_19207);
xor U20532 (N_20532,N_19296,N_19893);
nor U20533 (N_20533,N_19836,N_19725);
nand U20534 (N_20534,N_19738,N_19035);
or U20535 (N_20535,N_19951,N_19847);
or U20536 (N_20536,N_19660,N_19236);
nor U20537 (N_20537,N_19561,N_19530);
or U20538 (N_20538,N_19836,N_19330);
nor U20539 (N_20539,N_19942,N_19820);
or U20540 (N_20540,N_19467,N_19882);
xor U20541 (N_20541,N_19917,N_19223);
and U20542 (N_20542,N_19111,N_19659);
and U20543 (N_20543,N_19291,N_19016);
xor U20544 (N_20544,N_19928,N_19759);
and U20545 (N_20545,N_19333,N_19282);
or U20546 (N_20546,N_19153,N_19929);
xnor U20547 (N_20547,N_19131,N_19030);
nand U20548 (N_20548,N_19326,N_19422);
xor U20549 (N_20549,N_19636,N_19998);
nor U20550 (N_20550,N_19688,N_19034);
nand U20551 (N_20551,N_19844,N_19113);
or U20552 (N_20552,N_19601,N_19000);
or U20553 (N_20553,N_19733,N_19668);
and U20554 (N_20554,N_19104,N_19378);
xnor U20555 (N_20555,N_19314,N_19240);
xnor U20556 (N_20556,N_19943,N_19606);
or U20557 (N_20557,N_19941,N_19683);
or U20558 (N_20558,N_19497,N_19138);
and U20559 (N_20559,N_19713,N_19210);
nand U20560 (N_20560,N_19572,N_19896);
and U20561 (N_20561,N_19350,N_19857);
or U20562 (N_20562,N_19822,N_19259);
or U20563 (N_20563,N_19533,N_19678);
nor U20564 (N_20564,N_19390,N_19746);
or U20565 (N_20565,N_19881,N_19157);
or U20566 (N_20566,N_19619,N_19214);
or U20567 (N_20567,N_19646,N_19390);
or U20568 (N_20568,N_19115,N_19682);
and U20569 (N_20569,N_19161,N_19386);
xnor U20570 (N_20570,N_19120,N_19144);
xnor U20571 (N_20571,N_19678,N_19577);
nor U20572 (N_20572,N_19527,N_19537);
nor U20573 (N_20573,N_19418,N_19521);
nor U20574 (N_20574,N_19343,N_19715);
and U20575 (N_20575,N_19499,N_19196);
or U20576 (N_20576,N_19800,N_19351);
nand U20577 (N_20577,N_19768,N_19159);
xor U20578 (N_20578,N_19132,N_19353);
nand U20579 (N_20579,N_19326,N_19510);
or U20580 (N_20580,N_19847,N_19066);
nor U20581 (N_20581,N_19755,N_19869);
xnor U20582 (N_20582,N_19167,N_19748);
and U20583 (N_20583,N_19635,N_19959);
nand U20584 (N_20584,N_19174,N_19034);
nand U20585 (N_20585,N_19343,N_19624);
nand U20586 (N_20586,N_19262,N_19296);
and U20587 (N_20587,N_19598,N_19849);
xor U20588 (N_20588,N_19856,N_19681);
xnor U20589 (N_20589,N_19057,N_19463);
and U20590 (N_20590,N_19818,N_19220);
and U20591 (N_20591,N_19243,N_19523);
nand U20592 (N_20592,N_19470,N_19925);
or U20593 (N_20593,N_19445,N_19822);
and U20594 (N_20594,N_19846,N_19952);
nor U20595 (N_20595,N_19875,N_19509);
nand U20596 (N_20596,N_19793,N_19583);
xor U20597 (N_20597,N_19326,N_19248);
nand U20598 (N_20598,N_19157,N_19590);
or U20599 (N_20599,N_19591,N_19394);
xor U20600 (N_20600,N_19549,N_19381);
or U20601 (N_20601,N_19936,N_19798);
xor U20602 (N_20602,N_19487,N_19440);
nor U20603 (N_20603,N_19137,N_19498);
or U20604 (N_20604,N_19477,N_19118);
and U20605 (N_20605,N_19919,N_19549);
xor U20606 (N_20606,N_19181,N_19577);
or U20607 (N_20607,N_19961,N_19585);
nand U20608 (N_20608,N_19325,N_19813);
and U20609 (N_20609,N_19644,N_19779);
nand U20610 (N_20610,N_19042,N_19965);
xor U20611 (N_20611,N_19359,N_19885);
nand U20612 (N_20612,N_19129,N_19532);
and U20613 (N_20613,N_19924,N_19206);
xor U20614 (N_20614,N_19385,N_19216);
and U20615 (N_20615,N_19624,N_19209);
nor U20616 (N_20616,N_19891,N_19103);
or U20617 (N_20617,N_19403,N_19881);
or U20618 (N_20618,N_19468,N_19579);
nand U20619 (N_20619,N_19552,N_19908);
xnor U20620 (N_20620,N_19741,N_19202);
and U20621 (N_20621,N_19094,N_19235);
nor U20622 (N_20622,N_19639,N_19492);
or U20623 (N_20623,N_19978,N_19989);
nand U20624 (N_20624,N_19118,N_19163);
and U20625 (N_20625,N_19843,N_19688);
and U20626 (N_20626,N_19213,N_19072);
xnor U20627 (N_20627,N_19881,N_19371);
or U20628 (N_20628,N_19737,N_19009);
xnor U20629 (N_20629,N_19654,N_19188);
nor U20630 (N_20630,N_19263,N_19830);
or U20631 (N_20631,N_19270,N_19163);
nor U20632 (N_20632,N_19960,N_19343);
xnor U20633 (N_20633,N_19554,N_19912);
or U20634 (N_20634,N_19655,N_19024);
nor U20635 (N_20635,N_19197,N_19738);
and U20636 (N_20636,N_19338,N_19681);
xor U20637 (N_20637,N_19385,N_19683);
xor U20638 (N_20638,N_19772,N_19179);
nor U20639 (N_20639,N_19156,N_19216);
and U20640 (N_20640,N_19393,N_19765);
xor U20641 (N_20641,N_19964,N_19237);
xor U20642 (N_20642,N_19932,N_19929);
or U20643 (N_20643,N_19472,N_19482);
or U20644 (N_20644,N_19862,N_19392);
and U20645 (N_20645,N_19740,N_19392);
nor U20646 (N_20646,N_19812,N_19087);
or U20647 (N_20647,N_19556,N_19806);
or U20648 (N_20648,N_19935,N_19164);
xnor U20649 (N_20649,N_19020,N_19670);
nor U20650 (N_20650,N_19729,N_19991);
and U20651 (N_20651,N_19606,N_19098);
nand U20652 (N_20652,N_19929,N_19057);
and U20653 (N_20653,N_19906,N_19345);
xor U20654 (N_20654,N_19822,N_19511);
nand U20655 (N_20655,N_19090,N_19137);
xnor U20656 (N_20656,N_19164,N_19231);
nand U20657 (N_20657,N_19028,N_19475);
nor U20658 (N_20658,N_19070,N_19118);
or U20659 (N_20659,N_19650,N_19561);
nand U20660 (N_20660,N_19785,N_19547);
nor U20661 (N_20661,N_19281,N_19921);
and U20662 (N_20662,N_19116,N_19259);
xor U20663 (N_20663,N_19720,N_19027);
xor U20664 (N_20664,N_19446,N_19492);
and U20665 (N_20665,N_19377,N_19002);
xor U20666 (N_20666,N_19310,N_19569);
xnor U20667 (N_20667,N_19033,N_19026);
and U20668 (N_20668,N_19421,N_19893);
nand U20669 (N_20669,N_19433,N_19634);
nand U20670 (N_20670,N_19510,N_19898);
xnor U20671 (N_20671,N_19171,N_19536);
xnor U20672 (N_20672,N_19841,N_19770);
nor U20673 (N_20673,N_19392,N_19873);
and U20674 (N_20674,N_19358,N_19496);
nand U20675 (N_20675,N_19747,N_19363);
nor U20676 (N_20676,N_19298,N_19300);
and U20677 (N_20677,N_19249,N_19918);
or U20678 (N_20678,N_19000,N_19261);
or U20679 (N_20679,N_19108,N_19270);
nand U20680 (N_20680,N_19280,N_19647);
nand U20681 (N_20681,N_19114,N_19899);
xnor U20682 (N_20682,N_19654,N_19534);
xnor U20683 (N_20683,N_19835,N_19563);
nor U20684 (N_20684,N_19587,N_19197);
and U20685 (N_20685,N_19503,N_19586);
nand U20686 (N_20686,N_19242,N_19594);
or U20687 (N_20687,N_19658,N_19880);
nor U20688 (N_20688,N_19486,N_19747);
nand U20689 (N_20689,N_19201,N_19044);
nor U20690 (N_20690,N_19139,N_19203);
nand U20691 (N_20691,N_19091,N_19217);
xor U20692 (N_20692,N_19452,N_19672);
nand U20693 (N_20693,N_19740,N_19274);
xnor U20694 (N_20694,N_19635,N_19965);
nor U20695 (N_20695,N_19749,N_19528);
and U20696 (N_20696,N_19546,N_19536);
nor U20697 (N_20697,N_19805,N_19283);
or U20698 (N_20698,N_19002,N_19540);
nor U20699 (N_20699,N_19520,N_19745);
xnor U20700 (N_20700,N_19957,N_19783);
nand U20701 (N_20701,N_19118,N_19698);
xor U20702 (N_20702,N_19644,N_19636);
nor U20703 (N_20703,N_19917,N_19911);
xnor U20704 (N_20704,N_19400,N_19570);
or U20705 (N_20705,N_19583,N_19695);
nor U20706 (N_20706,N_19196,N_19013);
or U20707 (N_20707,N_19450,N_19180);
or U20708 (N_20708,N_19998,N_19572);
nor U20709 (N_20709,N_19979,N_19932);
nand U20710 (N_20710,N_19503,N_19329);
nor U20711 (N_20711,N_19058,N_19810);
and U20712 (N_20712,N_19542,N_19610);
or U20713 (N_20713,N_19792,N_19421);
nor U20714 (N_20714,N_19181,N_19004);
and U20715 (N_20715,N_19474,N_19711);
or U20716 (N_20716,N_19747,N_19814);
or U20717 (N_20717,N_19724,N_19754);
and U20718 (N_20718,N_19509,N_19069);
and U20719 (N_20719,N_19224,N_19853);
nor U20720 (N_20720,N_19366,N_19111);
or U20721 (N_20721,N_19348,N_19199);
xor U20722 (N_20722,N_19298,N_19288);
nor U20723 (N_20723,N_19719,N_19465);
and U20724 (N_20724,N_19666,N_19843);
nand U20725 (N_20725,N_19956,N_19139);
or U20726 (N_20726,N_19557,N_19071);
and U20727 (N_20727,N_19669,N_19241);
nand U20728 (N_20728,N_19115,N_19878);
nand U20729 (N_20729,N_19484,N_19539);
or U20730 (N_20730,N_19033,N_19291);
or U20731 (N_20731,N_19356,N_19962);
nor U20732 (N_20732,N_19235,N_19351);
nor U20733 (N_20733,N_19761,N_19154);
or U20734 (N_20734,N_19610,N_19306);
nor U20735 (N_20735,N_19740,N_19134);
xor U20736 (N_20736,N_19911,N_19040);
xor U20737 (N_20737,N_19087,N_19899);
or U20738 (N_20738,N_19061,N_19205);
or U20739 (N_20739,N_19454,N_19799);
and U20740 (N_20740,N_19028,N_19290);
or U20741 (N_20741,N_19611,N_19515);
or U20742 (N_20742,N_19962,N_19074);
xor U20743 (N_20743,N_19041,N_19482);
or U20744 (N_20744,N_19422,N_19198);
xor U20745 (N_20745,N_19084,N_19772);
or U20746 (N_20746,N_19748,N_19258);
nand U20747 (N_20747,N_19370,N_19256);
xnor U20748 (N_20748,N_19387,N_19601);
nand U20749 (N_20749,N_19445,N_19864);
nor U20750 (N_20750,N_19697,N_19571);
and U20751 (N_20751,N_19843,N_19283);
xnor U20752 (N_20752,N_19538,N_19560);
nor U20753 (N_20753,N_19346,N_19261);
and U20754 (N_20754,N_19230,N_19574);
nand U20755 (N_20755,N_19650,N_19640);
nand U20756 (N_20756,N_19685,N_19684);
nor U20757 (N_20757,N_19678,N_19099);
nor U20758 (N_20758,N_19714,N_19691);
or U20759 (N_20759,N_19215,N_19351);
nand U20760 (N_20760,N_19987,N_19975);
nand U20761 (N_20761,N_19108,N_19368);
nand U20762 (N_20762,N_19242,N_19584);
or U20763 (N_20763,N_19135,N_19389);
nor U20764 (N_20764,N_19675,N_19353);
nor U20765 (N_20765,N_19719,N_19635);
nor U20766 (N_20766,N_19042,N_19006);
or U20767 (N_20767,N_19712,N_19515);
or U20768 (N_20768,N_19824,N_19237);
nor U20769 (N_20769,N_19541,N_19327);
xnor U20770 (N_20770,N_19930,N_19258);
and U20771 (N_20771,N_19911,N_19786);
nand U20772 (N_20772,N_19427,N_19982);
nand U20773 (N_20773,N_19071,N_19266);
nand U20774 (N_20774,N_19796,N_19068);
nor U20775 (N_20775,N_19484,N_19003);
nand U20776 (N_20776,N_19715,N_19276);
nor U20777 (N_20777,N_19796,N_19973);
nor U20778 (N_20778,N_19688,N_19348);
nor U20779 (N_20779,N_19260,N_19045);
or U20780 (N_20780,N_19096,N_19531);
nor U20781 (N_20781,N_19425,N_19208);
or U20782 (N_20782,N_19309,N_19741);
nand U20783 (N_20783,N_19417,N_19646);
xor U20784 (N_20784,N_19661,N_19202);
nand U20785 (N_20785,N_19543,N_19747);
or U20786 (N_20786,N_19113,N_19631);
or U20787 (N_20787,N_19014,N_19211);
or U20788 (N_20788,N_19706,N_19726);
nand U20789 (N_20789,N_19788,N_19678);
nand U20790 (N_20790,N_19586,N_19027);
and U20791 (N_20791,N_19614,N_19483);
xor U20792 (N_20792,N_19273,N_19609);
and U20793 (N_20793,N_19857,N_19334);
nor U20794 (N_20794,N_19405,N_19132);
nor U20795 (N_20795,N_19084,N_19809);
nor U20796 (N_20796,N_19473,N_19532);
and U20797 (N_20797,N_19848,N_19832);
and U20798 (N_20798,N_19555,N_19138);
nand U20799 (N_20799,N_19694,N_19968);
nand U20800 (N_20800,N_19952,N_19963);
nand U20801 (N_20801,N_19800,N_19627);
xor U20802 (N_20802,N_19361,N_19154);
nand U20803 (N_20803,N_19824,N_19367);
or U20804 (N_20804,N_19211,N_19486);
or U20805 (N_20805,N_19000,N_19648);
and U20806 (N_20806,N_19179,N_19581);
xor U20807 (N_20807,N_19548,N_19017);
nor U20808 (N_20808,N_19681,N_19446);
nand U20809 (N_20809,N_19189,N_19398);
nand U20810 (N_20810,N_19146,N_19594);
nand U20811 (N_20811,N_19860,N_19093);
nand U20812 (N_20812,N_19116,N_19529);
xnor U20813 (N_20813,N_19887,N_19625);
or U20814 (N_20814,N_19601,N_19508);
or U20815 (N_20815,N_19971,N_19987);
xnor U20816 (N_20816,N_19794,N_19411);
or U20817 (N_20817,N_19678,N_19497);
or U20818 (N_20818,N_19012,N_19900);
xnor U20819 (N_20819,N_19676,N_19374);
and U20820 (N_20820,N_19983,N_19288);
or U20821 (N_20821,N_19454,N_19009);
or U20822 (N_20822,N_19119,N_19285);
or U20823 (N_20823,N_19128,N_19255);
and U20824 (N_20824,N_19986,N_19512);
nor U20825 (N_20825,N_19666,N_19221);
nor U20826 (N_20826,N_19350,N_19957);
nor U20827 (N_20827,N_19448,N_19531);
nor U20828 (N_20828,N_19784,N_19774);
xnor U20829 (N_20829,N_19795,N_19441);
nand U20830 (N_20830,N_19797,N_19994);
nor U20831 (N_20831,N_19578,N_19515);
or U20832 (N_20832,N_19202,N_19168);
xnor U20833 (N_20833,N_19330,N_19011);
nand U20834 (N_20834,N_19290,N_19732);
nand U20835 (N_20835,N_19481,N_19973);
nor U20836 (N_20836,N_19216,N_19908);
nand U20837 (N_20837,N_19859,N_19363);
xor U20838 (N_20838,N_19056,N_19653);
xnor U20839 (N_20839,N_19675,N_19057);
or U20840 (N_20840,N_19659,N_19425);
nand U20841 (N_20841,N_19966,N_19120);
and U20842 (N_20842,N_19339,N_19632);
and U20843 (N_20843,N_19907,N_19809);
or U20844 (N_20844,N_19085,N_19865);
or U20845 (N_20845,N_19994,N_19409);
nor U20846 (N_20846,N_19267,N_19007);
nand U20847 (N_20847,N_19155,N_19483);
and U20848 (N_20848,N_19018,N_19491);
nor U20849 (N_20849,N_19949,N_19801);
nor U20850 (N_20850,N_19997,N_19295);
and U20851 (N_20851,N_19863,N_19193);
xor U20852 (N_20852,N_19068,N_19834);
xor U20853 (N_20853,N_19619,N_19543);
xnor U20854 (N_20854,N_19903,N_19917);
or U20855 (N_20855,N_19069,N_19500);
and U20856 (N_20856,N_19287,N_19108);
nor U20857 (N_20857,N_19027,N_19344);
and U20858 (N_20858,N_19166,N_19098);
nor U20859 (N_20859,N_19610,N_19994);
and U20860 (N_20860,N_19199,N_19030);
nor U20861 (N_20861,N_19384,N_19507);
xor U20862 (N_20862,N_19097,N_19182);
xor U20863 (N_20863,N_19049,N_19444);
and U20864 (N_20864,N_19136,N_19005);
and U20865 (N_20865,N_19457,N_19559);
and U20866 (N_20866,N_19121,N_19263);
xnor U20867 (N_20867,N_19408,N_19606);
nand U20868 (N_20868,N_19447,N_19219);
and U20869 (N_20869,N_19227,N_19442);
nor U20870 (N_20870,N_19297,N_19962);
nand U20871 (N_20871,N_19815,N_19862);
and U20872 (N_20872,N_19518,N_19200);
xnor U20873 (N_20873,N_19580,N_19228);
or U20874 (N_20874,N_19897,N_19892);
or U20875 (N_20875,N_19098,N_19544);
or U20876 (N_20876,N_19119,N_19998);
and U20877 (N_20877,N_19794,N_19084);
nor U20878 (N_20878,N_19731,N_19418);
nor U20879 (N_20879,N_19564,N_19849);
or U20880 (N_20880,N_19288,N_19680);
nand U20881 (N_20881,N_19153,N_19055);
nand U20882 (N_20882,N_19503,N_19736);
nor U20883 (N_20883,N_19448,N_19124);
nand U20884 (N_20884,N_19520,N_19159);
or U20885 (N_20885,N_19721,N_19604);
and U20886 (N_20886,N_19139,N_19856);
or U20887 (N_20887,N_19101,N_19899);
xor U20888 (N_20888,N_19235,N_19847);
and U20889 (N_20889,N_19346,N_19569);
nand U20890 (N_20890,N_19624,N_19109);
xor U20891 (N_20891,N_19845,N_19027);
and U20892 (N_20892,N_19491,N_19671);
and U20893 (N_20893,N_19785,N_19323);
or U20894 (N_20894,N_19466,N_19013);
xnor U20895 (N_20895,N_19152,N_19956);
and U20896 (N_20896,N_19242,N_19728);
or U20897 (N_20897,N_19816,N_19370);
nor U20898 (N_20898,N_19606,N_19963);
xnor U20899 (N_20899,N_19178,N_19157);
nand U20900 (N_20900,N_19575,N_19299);
and U20901 (N_20901,N_19591,N_19620);
nor U20902 (N_20902,N_19439,N_19828);
nor U20903 (N_20903,N_19666,N_19046);
xnor U20904 (N_20904,N_19704,N_19843);
xor U20905 (N_20905,N_19550,N_19154);
nor U20906 (N_20906,N_19340,N_19216);
nand U20907 (N_20907,N_19065,N_19086);
nor U20908 (N_20908,N_19325,N_19117);
nand U20909 (N_20909,N_19968,N_19321);
nor U20910 (N_20910,N_19531,N_19755);
xor U20911 (N_20911,N_19048,N_19470);
and U20912 (N_20912,N_19200,N_19081);
xnor U20913 (N_20913,N_19716,N_19675);
nand U20914 (N_20914,N_19895,N_19269);
nand U20915 (N_20915,N_19463,N_19566);
xnor U20916 (N_20916,N_19750,N_19533);
nor U20917 (N_20917,N_19441,N_19244);
xor U20918 (N_20918,N_19259,N_19153);
xor U20919 (N_20919,N_19726,N_19445);
or U20920 (N_20920,N_19728,N_19498);
and U20921 (N_20921,N_19528,N_19532);
nand U20922 (N_20922,N_19816,N_19717);
xnor U20923 (N_20923,N_19770,N_19385);
or U20924 (N_20924,N_19043,N_19467);
or U20925 (N_20925,N_19804,N_19963);
nor U20926 (N_20926,N_19910,N_19195);
and U20927 (N_20927,N_19905,N_19709);
or U20928 (N_20928,N_19614,N_19612);
nand U20929 (N_20929,N_19592,N_19403);
nor U20930 (N_20930,N_19492,N_19313);
or U20931 (N_20931,N_19328,N_19697);
xor U20932 (N_20932,N_19663,N_19490);
nand U20933 (N_20933,N_19440,N_19562);
nor U20934 (N_20934,N_19989,N_19807);
nor U20935 (N_20935,N_19397,N_19638);
nand U20936 (N_20936,N_19895,N_19537);
or U20937 (N_20937,N_19291,N_19528);
nor U20938 (N_20938,N_19916,N_19624);
or U20939 (N_20939,N_19778,N_19332);
or U20940 (N_20940,N_19731,N_19658);
or U20941 (N_20941,N_19191,N_19083);
nand U20942 (N_20942,N_19119,N_19669);
nor U20943 (N_20943,N_19469,N_19270);
nand U20944 (N_20944,N_19853,N_19453);
nor U20945 (N_20945,N_19281,N_19859);
or U20946 (N_20946,N_19440,N_19132);
nor U20947 (N_20947,N_19386,N_19705);
nor U20948 (N_20948,N_19599,N_19692);
nor U20949 (N_20949,N_19243,N_19736);
xor U20950 (N_20950,N_19736,N_19410);
or U20951 (N_20951,N_19572,N_19463);
nor U20952 (N_20952,N_19751,N_19412);
nand U20953 (N_20953,N_19536,N_19028);
or U20954 (N_20954,N_19279,N_19832);
nor U20955 (N_20955,N_19164,N_19768);
nor U20956 (N_20956,N_19374,N_19411);
nand U20957 (N_20957,N_19575,N_19320);
and U20958 (N_20958,N_19256,N_19464);
nand U20959 (N_20959,N_19557,N_19813);
nor U20960 (N_20960,N_19425,N_19188);
xor U20961 (N_20961,N_19505,N_19187);
xor U20962 (N_20962,N_19570,N_19150);
or U20963 (N_20963,N_19018,N_19537);
nor U20964 (N_20964,N_19373,N_19368);
nand U20965 (N_20965,N_19425,N_19331);
nor U20966 (N_20966,N_19777,N_19301);
and U20967 (N_20967,N_19021,N_19637);
nand U20968 (N_20968,N_19005,N_19525);
xnor U20969 (N_20969,N_19059,N_19204);
nand U20970 (N_20970,N_19969,N_19461);
nand U20971 (N_20971,N_19738,N_19372);
or U20972 (N_20972,N_19805,N_19711);
and U20973 (N_20973,N_19149,N_19402);
xor U20974 (N_20974,N_19967,N_19090);
or U20975 (N_20975,N_19086,N_19170);
xor U20976 (N_20976,N_19500,N_19269);
nor U20977 (N_20977,N_19280,N_19286);
xor U20978 (N_20978,N_19226,N_19815);
nand U20979 (N_20979,N_19809,N_19002);
and U20980 (N_20980,N_19571,N_19421);
or U20981 (N_20981,N_19308,N_19932);
xor U20982 (N_20982,N_19574,N_19279);
xor U20983 (N_20983,N_19734,N_19546);
or U20984 (N_20984,N_19024,N_19824);
or U20985 (N_20985,N_19694,N_19994);
and U20986 (N_20986,N_19717,N_19849);
nand U20987 (N_20987,N_19259,N_19296);
or U20988 (N_20988,N_19826,N_19013);
nand U20989 (N_20989,N_19057,N_19000);
nand U20990 (N_20990,N_19762,N_19410);
and U20991 (N_20991,N_19651,N_19405);
and U20992 (N_20992,N_19823,N_19671);
nor U20993 (N_20993,N_19102,N_19709);
nor U20994 (N_20994,N_19364,N_19093);
and U20995 (N_20995,N_19938,N_19029);
and U20996 (N_20996,N_19879,N_19342);
xnor U20997 (N_20997,N_19809,N_19330);
or U20998 (N_20998,N_19420,N_19765);
nor U20999 (N_20999,N_19431,N_19411);
and U21000 (N_21000,N_20293,N_20483);
and U21001 (N_21001,N_20491,N_20811);
nor U21002 (N_21002,N_20065,N_20095);
xor U21003 (N_21003,N_20568,N_20577);
or U21004 (N_21004,N_20130,N_20376);
xor U21005 (N_21005,N_20447,N_20575);
xnor U21006 (N_21006,N_20779,N_20285);
nor U21007 (N_21007,N_20528,N_20730);
or U21008 (N_21008,N_20451,N_20709);
and U21009 (N_21009,N_20386,N_20107);
nor U21010 (N_21010,N_20513,N_20727);
or U21011 (N_21011,N_20123,N_20714);
nand U21012 (N_21012,N_20196,N_20075);
nand U21013 (N_21013,N_20295,N_20452);
xnor U21014 (N_21014,N_20755,N_20847);
and U21015 (N_21015,N_20978,N_20237);
and U21016 (N_21016,N_20702,N_20383);
xnor U21017 (N_21017,N_20392,N_20300);
nor U21018 (N_21018,N_20445,N_20228);
nor U21019 (N_21019,N_20957,N_20203);
nand U21020 (N_21020,N_20630,N_20471);
and U21021 (N_21021,N_20002,N_20443);
nand U21022 (N_21022,N_20205,N_20360);
or U21023 (N_21023,N_20820,N_20052);
nor U21024 (N_21024,N_20043,N_20391);
or U21025 (N_21025,N_20686,N_20314);
nand U21026 (N_21026,N_20051,N_20519);
or U21027 (N_21027,N_20121,N_20348);
xor U21028 (N_21028,N_20692,N_20767);
or U21029 (N_21029,N_20098,N_20414);
nand U21030 (N_21030,N_20966,N_20637);
and U21031 (N_21031,N_20358,N_20380);
xor U21032 (N_21032,N_20803,N_20060);
nor U21033 (N_21033,N_20265,N_20101);
and U21034 (N_21034,N_20160,N_20061);
and U21035 (N_21035,N_20495,N_20674);
or U21036 (N_21036,N_20393,N_20835);
xnor U21037 (N_21037,N_20352,N_20961);
nor U21038 (N_21038,N_20777,N_20087);
nand U21039 (N_21039,N_20142,N_20673);
nor U21040 (N_21040,N_20343,N_20786);
xor U21041 (N_21041,N_20467,N_20959);
and U21042 (N_21042,N_20888,N_20639);
nor U21043 (N_21043,N_20849,N_20861);
nand U21044 (N_21044,N_20602,N_20970);
nor U21045 (N_21045,N_20603,N_20442);
or U21046 (N_21046,N_20643,N_20684);
and U21047 (N_21047,N_20672,N_20950);
and U21048 (N_21048,N_20748,N_20428);
or U21049 (N_21049,N_20449,N_20897);
or U21050 (N_21050,N_20817,N_20521);
and U21051 (N_21051,N_20553,N_20907);
nor U21052 (N_21052,N_20113,N_20222);
or U21053 (N_21053,N_20814,N_20944);
nor U21054 (N_21054,N_20766,N_20901);
nand U21055 (N_21055,N_20439,N_20598);
nor U21056 (N_21056,N_20865,N_20485);
and U21057 (N_21057,N_20517,N_20546);
nand U21058 (N_21058,N_20468,N_20063);
nor U21059 (N_21059,N_20460,N_20119);
and U21060 (N_21060,N_20241,N_20464);
nand U21061 (N_21061,N_20923,N_20840);
nand U21062 (N_21062,N_20206,N_20373);
xnor U21063 (N_21063,N_20789,N_20252);
and U21064 (N_21064,N_20932,N_20627);
nor U21065 (N_21065,N_20006,N_20289);
nand U21066 (N_21066,N_20470,N_20868);
xnor U21067 (N_21067,N_20039,N_20132);
and U21068 (N_21068,N_20220,N_20042);
or U21069 (N_21069,N_20848,N_20871);
xor U21070 (N_21070,N_20251,N_20448);
xor U21071 (N_21071,N_20930,N_20151);
nor U21072 (N_21072,N_20525,N_20836);
xnor U21073 (N_21073,N_20563,N_20677);
or U21074 (N_21074,N_20171,N_20009);
and U21075 (N_21075,N_20140,N_20549);
nand U21076 (N_21076,N_20083,N_20256);
nand U21077 (N_21077,N_20965,N_20004);
or U21078 (N_21078,N_20407,N_20413);
or U21079 (N_21079,N_20729,N_20921);
xor U21080 (N_21080,N_20790,N_20236);
or U21081 (N_21081,N_20510,N_20033);
nor U21082 (N_21082,N_20474,N_20813);
and U21083 (N_21083,N_20092,N_20557);
or U21084 (N_21084,N_20615,N_20906);
or U21085 (N_21085,N_20586,N_20411);
or U21086 (N_21086,N_20760,N_20512);
nand U21087 (N_21087,N_20867,N_20515);
and U21088 (N_21088,N_20096,N_20303);
nand U21089 (N_21089,N_20772,N_20860);
xnor U21090 (N_21090,N_20543,N_20926);
or U21091 (N_21091,N_20663,N_20556);
or U21092 (N_21092,N_20053,N_20079);
nor U21093 (N_21093,N_20209,N_20631);
xor U21094 (N_21094,N_20283,N_20642);
or U21095 (N_21095,N_20605,N_20272);
and U21096 (N_21096,N_20821,N_20987);
or U21097 (N_21097,N_20873,N_20403);
or U21098 (N_21098,N_20610,N_20902);
nor U21099 (N_21099,N_20010,N_20183);
xnor U21100 (N_21100,N_20837,N_20914);
or U21101 (N_21101,N_20698,N_20885);
xnor U21102 (N_21102,N_20658,N_20647);
xor U21103 (N_21103,N_20752,N_20405);
xor U21104 (N_21104,N_20437,N_20340);
or U21105 (N_21105,N_20750,N_20851);
nand U21106 (N_21106,N_20102,N_20170);
or U21107 (N_21107,N_20382,N_20090);
and U21108 (N_21108,N_20762,N_20511);
or U21109 (N_21109,N_20747,N_20131);
or U21110 (N_21110,N_20884,N_20030);
xor U21111 (N_21111,N_20336,N_20891);
or U21112 (N_21112,N_20980,N_20420);
xor U21113 (N_21113,N_20408,N_20216);
nand U21114 (N_21114,N_20450,N_20309);
nand U21115 (N_21115,N_20527,N_20943);
nand U21116 (N_21116,N_20623,N_20068);
xor U21117 (N_21117,N_20640,N_20255);
or U21118 (N_21118,N_20618,N_20812);
or U21119 (N_21119,N_20617,N_20355);
nor U21120 (N_21120,N_20955,N_20248);
xor U21121 (N_21121,N_20188,N_20286);
and U21122 (N_21122,N_20372,N_20981);
nor U21123 (N_21123,N_20863,N_20636);
and U21124 (N_21124,N_20224,N_20937);
xnor U21125 (N_21125,N_20167,N_20281);
and U21126 (N_21126,N_20818,N_20128);
nor U21127 (N_21127,N_20632,N_20192);
or U21128 (N_21128,N_20784,N_20889);
xnor U21129 (N_21129,N_20035,N_20280);
nor U21130 (N_21130,N_20975,N_20141);
nand U21131 (N_21131,N_20333,N_20268);
and U21132 (N_21132,N_20324,N_20184);
nand U21133 (N_21133,N_20362,N_20014);
and U21134 (N_21134,N_20387,N_20825);
xnor U21135 (N_21135,N_20080,N_20683);
nor U21136 (N_21136,N_20626,N_20735);
xor U21137 (N_21137,N_20609,N_20751);
and U21138 (N_21138,N_20562,N_20017);
nand U21139 (N_21139,N_20720,N_20866);
nand U21140 (N_21140,N_20354,N_20259);
nand U21141 (N_21141,N_20071,N_20593);
nand U21142 (N_21142,N_20328,N_20246);
and U21143 (N_21143,N_20941,N_20409);
nand U21144 (N_21144,N_20419,N_20581);
and U21145 (N_21145,N_20578,N_20505);
and U21146 (N_21146,N_20584,N_20041);
xnor U21147 (N_21147,N_20377,N_20179);
or U21148 (N_21148,N_20345,N_20230);
nor U21149 (N_21149,N_20958,N_20552);
nor U21150 (N_21150,N_20696,N_20652);
nand U21151 (N_21151,N_20815,N_20862);
xor U21152 (N_21152,N_20430,N_20768);
or U21153 (N_21153,N_20242,N_20590);
nor U21154 (N_21154,N_20124,N_20180);
and U21155 (N_21155,N_20369,N_20162);
and U21156 (N_21156,N_20995,N_20267);
or U21157 (N_21157,N_20507,N_20661);
nor U21158 (N_21158,N_20695,N_20298);
and U21159 (N_21159,N_20898,N_20534);
and U21160 (N_21160,N_20013,N_20899);
or U21161 (N_21161,N_20846,N_20879);
and U21162 (N_21162,N_20149,N_20843);
xor U21163 (N_21163,N_20560,N_20761);
or U21164 (N_21164,N_20582,N_20659);
and U21165 (N_21165,N_20500,N_20462);
xnor U21166 (N_21166,N_20839,N_20084);
nand U21167 (N_21167,N_20611,N_20669);
xor U21168 (N_21168,N_20478,N_20194);
xnor U21169 (N_21169,N_20480,N_20089);
nand U21170 (N_21170,N_20935,N_20435);
and U21171 (N_21171,N_20163,N_20019);
nor U21172 (N_21172,N_20415,N_20620);
and U21173 (N_21173,N_20774,N_20508);
nor U21174 (N_21174,N_20402,N_20667);
or U21175 (N_21175,N_20938,N_20799);
nand U21176 (N_21176,N_20954,N_20833);
nand U21177 (N_21177,N_20710,N_20368);
nor U21178 (N_21178,N_20134,N_20919);
nand U21179 (N_21179,N_20078,N_20091);
or U21180 (N_21180,N_20796,N_20262);
xnor U21181 (N_21181,N_20936,N_20335);
or U21182 (N_21182,N_20502,N_20423);
xor U21183 (N_21183,N_20506,N_20156);
nor U21184 (N_21184,N_20484,N_20493);
or U21185 (N_21185,N_20634,N_20133);
nand U21186 (N_21186,N_20308,N_20707);
and U21187 (N_21187,N_20600,N_20153);
nand U21188 (N_21188,N_20217,N_20759);
xor U21189 (N_21189,N_20214,N_20122);
nand U21190 (N_21190,N_20797,N_20622);
nand U21191 (N_21191,N_20773,N_20106);
nor U21192 (N_21192,N_20016,N_20597);
or U21193 (N_21193,N_20388,N_20972);
or U21194 (N_21194,N_20655,N_20794);
or U21195 (N_21195,N_20422,N_20145);
or U21196 (N_21196,N_20073,N_20573);
nor U21197 (N_21197,N_20296,N_20801);
or U21198 (N_21198,N_20390,N_20964);
or U21199 (N_21199,N_20226,N_20215);
or U21200 (N_21200,N_20099,N_20717);
nand U21201 (N_21201,N_20219,N_20742);
xnor U21202 (N_21202,N_20895,N_20644);
and U21203 (N_21203,N_20074,N_20317);
and U21204 (N_21204,N_20646,N_20271);
and U21205 (N_21205,N_20872,N_20116);
nor U21206 (N_21206,N_20713,N_20081);
nor U21207 (N_21207,N_20323,N_20304);
xor U21208 (N_21208,N_20931,N_20332);
and U21209 (N_21209,N_20998,N_20218);
xor U21210 (N_21210,N_20693,N_20595);
xnor U21211 (N_21211,N_20962,N_20136);
nand U21212 (N_21212,N_20208,N_20334);
xnor U21213 (N_21213,N_20278,N_20614);
and U21214 (N_21214,N_20723,N_20356);
and U21215 (N_21215,N_20800,N_20088);
nor U21216 (N_21216,N_20859,N_20886);
or U21217 (N_21217,N_20749,N_20746);
xor U21218 (N_21218,N_20986,N_20864);
and U21219 (N_21219,N_20533,N_20469);
xnor U21220 (N_21220,N_20910,N_20753);
xor U21221 (N_21221,N_20550,N_20370);
nand U21222 (N_21222,N_20441,N_20858);
nor U21223 (N_21223,N_20728,N_20971);
nor U21224 (N_21224,N_20745,N_20915);
nand U21225 (N_21225,N_20952,N_20911);
nand U21226 (N_21226,N_20706,N_20401);
nor U21227 (N_21227,N_20616,N_20488);
xor U21228 (N_21228,N_20651,N_20181);
nor U21229 (N_21229,N_20275,N_20664);
and U21230 (N_21230,N_20305,N_20904);
xor U21231 (N_21231,N_20487,N_20732);
or U21232 (N_21232,N_20680,N_20263);
or U21233 (N_21233,N_20307,N_20816);
and U21234 (N_21234,N_20887,N_20315);
nor U21235 (N_21235,N_20810,N_20780);
or U21236 (N_21236,N_20809,N_20892);
or U21237 (N_21237,N_20976,N_20571);
or U21238 (N_21238,N_20824,N_20031);
xnor U21239 (N_21239,N_20421,N_20077);
and U21240 (N_21240,N_20665,N_20754);
xnor U21241 (N_21241,N_20055,N_20537);
nor U21242 (N_21242,N_20249,N_20461);
nor U21243 (N_21243,N_20666,N_20114);
nand U21244 (N_21244,N_20704,N_20570);
or U21245 (N_21245,N_20700,N_20711);
nand U21246 (N_21246,N_20339,N_20979);
xor U21247 (N_21247,N_20601,N_20701);
xnor U21248 (N_21248,N_20826,N_20805);
or U21249 (N_21249,N_20604,N_20908);
or U21250 (N_21250,N_20266,N_20522);
xnor U21251 (N_21251,N_20118,N_20227);
nor U21252 (N_21252,N_20231,N_20139);
or U21253 (N_21253,N_20853,N_20044);
xnor U21254 (N_21254,N_20302,N_20086);
nand U21255 (N_21255,N_20486,N_20594);
and U21256 (N_21256,N_20771,N_20916);
nand U21257 (N_21257,N_20465,N_20148);
or U21258 (N_21258,N_20635,N_20558);
or U21259 (N_21259,N_20656,N_20318);
xor U21260 (N_21260,N_20679,N_20164);
nor U21261 (N_21261,N_20934,N_20791);
or U21262 (N_21262,N_20406,N_20621);
or U21263 (N_21263,N_20154,N_20040);
and U21264 (N_21264,N_20261,N_20829);
nor U21265 (N_21265,N_20662,N_20353);
nand U21266 (N_21266,N_20740,N_20798);
or U21267 (N_21267,N_20349,N_20518);
xor U21268 (N_21268,N_20769,N_20433);
xnor U21269 (N_21269,N_20776,N_20225);
nand U21270 (N_21270,N_20426,N_20011);
nor U21271 (N_21271,N_20947,N_20559);
xor U21272 (N_21272,N_20725,N_20320);
and U21273 (N_21273,N_20482,N_20808);
or U21274 (N_21274,N_20330,N_20765);
or U21275 (N_21275,N_20691,N_20221);
and U21276 (N_21276,N_20857,N_20120);
nand U21277 (N_21277,N_20306,N_20361);
and U21278 (N_21278,N_20182,N_20008);
nor U21279 (N_21279,N_20032,N_20440);
nand U21280 (N_21280,N_20366,N_20946);
nand U21281 (N_21281,N_20069,N_20492);
xnor U21282 (N_21282,N_20290,N_20681);
xor U21283 (N_21283,N_20240,N_20319);
xor U21284 (N_21284,N_20466,N_20172);
xor U21285 (N_21285,N_20007,N_20195);
and U21286 (N_21286,N_20424,N_20948);
nand U21287 (N_21287,N_20253,N_20175);
xnor U21288 (N_21288,N_20737,N_20516);
and U21289 (N_21289,N_20778,N_20158);
or U21290 (N_21290,N_20399,N_20325);
nand U21291 (N_21291,N_20731,N_20150);
nor U21292 (N_21292,N_20671,N_20375);
and U21293 (N_21293,N_20331,N_20456);
nand U21294 (N_21294,N_20363,N_20104);
or U21295 (N_21295,N_20381,N_20257);
nand U21296 (N_21296,N_20715,N_20574);
nor U21297 (N_21297,N_20223,N_20342);
nand U21298 (N_21298,N_20625,N_20876);
xnor U21299 (N_21299,N_20144,N_20384);
and U21300 (N_21300,N_20596,N_20347);
nand U21301 (N_21301,N_20279,N_20189);
nand U21302 (N_21302,N_20260,N_20210);
nor U21303 (N_21303,N_20024,N_20023);
or U21304 (N_21304,N_20992,N_20034);
nor U21305 (N_21305,N_20893,N_20193);
xnor U21306 (N_21306,N_20657,N_20988);
or U21307 (N_21307,N_20394,N_20481);
nand U21308 (N_21308,N_20057,N_20756);
nand U21309 (N_21309,N_20476,N_20579);
or U21310 (N_21310,N_20254,N_20722);
nand U21311 (N_21311,N_20135,N_20832);
or U21312 (N_21312,N_20870,N_20048);
and U21313 (N_21313,N_20496,N_20173);
nand U21314 (N_21314,N_20159,N_20933);
or U21315 (N_21315,N_20599,N_20770);
nand U21316 (N_21316,N_20125,N_20234);
nor U21317 (N_21317,N_20066,N_20690);
nor U21318 (N_21318,N_20344,N_20875);
xor U21319 (N_21319,N_20896,N_20292);
xor U21320 (N_21320,N_20564,N_20396);
and U21321 (N_21321,N_20269,N_20472);
nand U21322 (N_21322,N_20850,N_20997);
nand U21323 (N_21323,N_20067,N_20922);
or U21324 (N_21324,N_20878,N_20258);
nor U21325 (N_21325,N_20565,N_20416);
or U21326 (N_21326,N_20270,N_20346);
and U21327 (N_21327,N_20058,N_20412);
nor U21328 (N_21328,N_20022,N_20689);
xor U21329 (N_21329,N_20021,N_20912);
nor U21330 (N_21330,N_20338,N_20374);
or U21331 (N_21331,N_20903,N_20050);
or U21332 (N_21332,N_20494,N_20233);
xnor U21333 (N_21333,N_20956,N_20670);
xnor U21334 (N_21334,N_20977,N_20117);
nor U21335 (N_21335,N_20152,N_20991);
nor U21336 (N_21336,N_20070,N_20882);
or U21337 (N_21337,N_20458,N_20703);
or U21338 (N_21338,N_20350,N_20539);
and U21339 (N_21339,N_20327,N_20247);
and U21340 (N_21340,N_20112,N_20842);
or U21341 (N_21341,N_20554,N_20076);
nand U21342 (N_21342,N_20973,N_20201);
xor U21343 (N_21343,N_20400,N_20238);
and U21344 (N_21344,N_20498,N_20953);
xnor U21345 (N_21345,N_20688,N_20436);
nor U21346 (N_21346,N_20367,N_20479);
nand U21347 (N_21347,N_20186,N_20329);
and U21348 (N_21348,N_20744,N_20542);
and U21349 (N_21349,N_20446,N_20585);
and U21350 (N_21350,N_20326,N_20109);
and U21351 (N_21351,N_20029,N_20115);
xnor U21352 (N_21352,N_20294,N_20204);
and U21353 (N_21353,N_20037,N_20082);
and U21354 (N_21354,N_20675,N_20982);
or U21355 (N_21355,N_20273,N_20127);
xor U21356 (N_21356,N_20190,N_20503);
nor U21357 (N_21357,N_20883,N_20569);
and U21358 (N_21358,N_20477,N_20277);
nand U21359 (N_21359,N_20716,N_20687);
xor U21360 (N_21360,N_20100,N_20185);
and U21361 (N_21361,N_20489,N_20985);
xnor U21362 (N_21362,N_20245,N_20712);
or U21363 (N_21363,N_20807,N_20591);
or U21364 (N_21364,N_20705,N_20398);
and U21365 (N_21365,N_20459,N_20168);
nor U21366 (N_21366,N_20945,N_20660);
or U21367 (N_21367,N_20110,N_20138);
xor U21368 (N_21368,N_20782,N_20454);
xnor U21369 (N_21369,N_20589,N_20404);
nor U21370 (N_21370,N_20536,N_20645);
xor U21371 (N_21371,N_20845,N_20990);
and U21372 (N_21372,N_20576,N_20909);
or U21373 (N_21373,N_20619,N_20429);
nand U21374 (N_21374,N_20453,N_20996);
xor U21375 (N_21375,N_20566,N_20146);
nor U21376 (N_21376,N_20207,N_20551);
nand U21377 (N_21377,N_20178,N_20788);
or U21378 (N_21378,N_20359,N_20301);
or U21379 (N_21379,N_20905,N_20917);
nand U21380 (N_21380,N_20613,N_20097);
or U21381 (N_21381,N_20699,N_20795);
xnor U21382 (N_21382,N_20365,N_20020);
nand U21383 (N_21383,N_20624,N_20697);
and U21384 (N_21384,N_20852,N_20000);
nand U21385 (N_21385,N_20529,N_20969);
nor U21386 (N_21386,N_20137,N_20321);
nand U21387 (N_21387,N_20877,N_20607);
nor U21388 (N_21388,N_20927,N_20351);
or U21389 (N_21389,N_20567,N_20587);
nor U21390 (N_21390,N_20191,N_20025);
or U21391 (N_21391,N_20913,N_20758);
xnor U21392 (N_21392,N_20027,N_20900);
nor U21393 (N_21393,N_20918,N_20177);
nand U21394 (N_21394,N_20444,N_20721);
xor U21395 (N_21395,N_20741,N_20176);
or U21396 (N_21396,N_20583,N_20984);
or U21397 (N_21397,N_20804,N_20299);
nor U21398 (N_21398,N_20739,N_20555);
xor U21399 (N_21399,N_20960,N_20685);
nand U21400 (N_21400,N_20827,N_20874);
nor U21401 (N_21401,N_20499,N_20418);
nor U21402 (N_21402,N_20038,N_20062);
or U21403 (N_21403,N_20592,N_20337);
and U21404 (N_21404,N_20427,N_20763);
nand U21405 (N_21405,N_20783,N_20274);
or U21406 (N_21406,N_20432,N_20561);
nor U21407 (N_21407,N_20385,N_20650);
or U21408 (N_21408,N_20371,N_20920);
and U21409 (N_21409,N_20473,N_20417);
nor U21410 (N_21410,N_20654,N_20316);
xnor U21411 (N_21411,N_20802,N_20379);
or U21412 (N_21412,N_20572,N_20003);
xor U21413 (N_21413,N_20504,N_20046);
and U21414 (N_21414,N_20649,N_20924);
or U21415 (N_21415,N_20830,N_20054);
xor U21416 (N_21416,N_20856,N_20243);
nand U21417 (N_21417,N_20734,N_20284);
and U21418 (N_21418,N_20736,N_20668);
or U21419 (N_21419,N_20198,N_20520);
xnor U21420 (N_21420,N_20169,N_20297);
nor U21421 (N_21421,N_20588,N_20049);
nand U21422 (N_21422,N_20085,N_20881);
xnor U21423 (N_21423,N_20580,N_20854);
and U21424 (N_21424,N_20166,N_20841);
nand U21425 (N_21425,N_20831,N_20819);
nor U21426 (N_21426,N_20264,N_20925);
or U21427 (N_21427,N_20785,N_20457);
xnor U21428 (N_21428,N_20232,N_20229);
or U21429 (N_21429,N_20501,N_20928);
xor U21430 (N_21430,N_20056,N_20341);
nor U21431 (N_21431,N_20431,N_20047);
xnor U21432 (N_21432,N_20531,N_20781);
or U21433 (N_21433,N_20855,N_20397);
or U21434 (N_21434,N_20111,N_20822);
or U21435 (N_21435,N_20526,N_20165);
or U21436 (N_21436,N_20993,N_20103);
nor U21437 (N_21437,N_20202,N_20806);
or U21438 (N_21438,N_20288,N_20108);
and U21439 (N_21439,N_20028,N_20757);
and U21440 (N_21440,N_20678,N_20129);
nand U21441 (N_21441,N_20548,N_20235);
nor U21442 (N_21442,N_20395,N_20357);
or U21443 (N_21443,N_20793,N_20743);
nor U21444 (N_21444,N_20005,N_20844);
nor U21445 (N_21445,N_20282,N_20497);
nand U21446 (N_21446,N_20523,N_20276);
nand U21447 (N_21447,N_20015,N_20161);
xor U21448 (N_21448,N_20733,N_20514);
nand U21449 (N_21449,N_20641,N_20438);
nand U21450 (N_21450,N_20994,N_20434);
xnor U21451 (N_21451,N_20648,N_20838);
nand U21452 (N_21452,N_20983,N_20093);
xor U21453 (N_21453,N_20726,N_20147);
nand U21454 (N_21454,N_20547,N_20792);
nor U21455 (N_21455,N_20989,N_20239);
nor U21456 (N_21456,N_20187,N_20718);
and U21457 (N_21457,N_20869,N_20545);
nor U21458 (N_21458,N_20212,N_20764);
and U21459 (N_21459,N_20026,N_20942);
and U21460 (N_21460,N_20939,N_20828);
or U21461 (N_21461,N_20929,N_20463);
or U21462 (N_21462,N_20018,N_20197);
and U21463 (N_21463,N_20425,N_20951);
and U21464 (N_21464,N_20880,N_20532);
xor U21465 (N_21465,N_20682,N_20894);
or U21466 (N_21466,N_20312,N_20064);
xor U21467 (N_21467,N_20045,N_20940);
xnor U21468 (N_21468,N_20708,N_20105);
xor U21469 (N_21469,N_20157,N_20541);
or U21470 (N_21470,N_20738,N_20694);
or U21471 (N_21471,N_20638,N_20378);
or U21472 (N_21472,N_20834,N_20036);
and U21473 (N_21473,N_20968,N_20540);
nor U21474 (N_21474,N_20509,N_20143);
or U21475 (N_21475,N_20633,N_20126);
or U21476 (N_21476,N_20199,N_20389);
and U21477 (N_21477,N_20311,N_20544);
nor U21478 (N_21478,N_20538,N_20612);
xor U21479 (N_21479,N_20155,N_20012);
nor U21480 (N_21480,N_20999,N_20719);
xor U21481 (N_21481,N_20001,N_20535);
and U21482 (N_21482,N_20524,N_20291);
or U21483 (N_21483,N_20967,N_20364);
or U21484 (N_21484,N_20608,N_20322);
nand U21485 (N_21485,N_20211,N_20490);
nor U21486 (N_21486,N_20072,N_20310);
and U21487 (N_21487,N_20628,N_20724);
nor U21488 (N_21488,N_20250,N_20775);
or U21489 (N_21489,N_20455,N_20974);
nor U21490 (N_21490,N_20606,N_20213);
nand U21491 (N_21491,N_20629,N_20823);
nor U21492 (N_21492,N_20653,N_20787);
or U21493 (N_21493,N_20410,N_20963);
and U21494 (N_21494,N_20059,N_20949);
and U21495 (N_21495,N_20676,N_20244);
and U21496 (N_21496,N_20890,N_20174);
nor U21497 (N_21497,N_20530,N_20200);
or U21498 (N_21498,N_20094,N_20475);
nand U21499 (N_21499,N_20313,N_20287);
or U21500 (N_21500,N_20832,N_20826);
nand U21501 (N_21501,N_20058,N_20810);
and U21502 (N_21502,N_20688,N_20977);
xor U21503 (N_21503,N_20108,N_20639);
xnor U21504 (N_21504,N_20900,N_20430);
or U21505 (N_21505,N_20580,N_20296);
and U21506 (N_21506,N_20379,N_20528);
and U21507 (N_21507,N_20879,N_20936);
and U21508 (N_21508,N_20657,N_20619);
or U21509 (N_21509,N_20640,N_20346);
nor U21510 (N_21510,N_20227,N_20632);
or U21511 (N_21511,N_20329,N_20688);
nand U21512 (N_21512,N_20651,N_20655);
or U21513 (N_21513,N_20596,N_20888);
and U21514 (N_21514,N_20838,N_20452);
and U21515 (N_21515,N_20769,N_20087);
or U21516 (N_21516,N_20106,N_20090);
nor U21517 (N_21517,N_20437,N_20423);
nor U21518 (N_21518,N_20766,N_20546);
and U21519 (N_21519,N_20495,N_20456);
or U21520 (N_21520,N_20377,N_20979);
nor U21521 (N_21521,N_20096,N_20778);
or U21522 (N_21522,N_20548,N_20733);
or U21523 (N_21523,N_20379,N_20476);
or U21524 (N_21524,N_20212,N_20307);
nand U21525 (N_21525,N_20902,N_20978);
nand U21526 (N_21526,N_20267,N_20100);
xor U21527 (N_21527,N_20983,N_20143);
xor U21528 (N_21528,N_20581,N_20545);
nand U21529 (N_21529,N_20040,N_20509);
xor U21530 (N_21530,N_20941,N_20760);
nand U21531 (N_21531,N_20913,N_20949);
xnor U21532 (N_21532,N_20183,N_20425);
nand U21533 (N_21533,N_20688,N_20789);
and U21534 (N_21534,N_20153,N_20347);
and U21535 (N_21535,N_20119,N_20723);
nand U21536 (N_21536,N_20143,N_20040);
nand U21537 (N_21537,N_20606,N_20354);
nand U21538 (N_21538,N_20152,N_20505);
or U21539 (N_21539,N_20313,N_20354);
nand U21540 (N_21540,N_20835,N_20454);
and U21541 (N_21541,N_20842,N_20824);
and U21542 (N_21542,N_20634,N_20924);
nand U21543 (N_21543,N_20115,N_20444);
nor U21544 (N_21544,N_20531,N_20187);
or U21545 (N_21545,N_20750,N_20117);
xor U21546 (N_21546,N_20091,N_20445);
nor U21547 (N_21547,N_20648,N_20090);
and U21548 (N_21548,N_20600,N_20574);
nand U21549 (N_21549,N_20066,N_20301);
xnor U21550 (N_21550,N_20597,N_20188);
nor U21551 (N_21551,N_20420,N_20301);
and U21552 (N_21552,N_20709,N_20223);
nand U21553 (N_21553,N_20519,N_20096);
xor U21554 (N_21554,N_20769,N_20328);
and U21555 (N_21555,N_20756,N_20077);
nor U21556 (N_21556,N_20713,N_20213);
nor U21557 (N_21557,N_20889,N_20483);
or U21558 (N_21558,N_20277,N_20634);
and U21559 (N_21559,N_20384,N_20076);
nand U21560 (N_21560,N_20899,N_20704);
and U21561 (N_21561,N_20805,N_20986);
and U21562 (N_21562,N_20484,N_20681);
xor U21563 (N_21563,N_20169,N_20388);
or U21564 (N_21564,N_20301,N_20159);
xor U21565 (N_21565,N_20769,N_20015);
xor U21566 (N_21566,N_20039,N_20137);
xnor U21567 (N_21567,N_20707,N_20801);
nand U21568 (N_21568,N_20142,N_20770);
nand U21569 (N_21569,N_20874,N_20104);
nand U21570 (N_21570,N_20748,N_20908);
or U21571 (N_21571,N_20602,N_20373);
nand U21572 (N_21572,N_20774,N_20150);
or U21573 (N_21573,N_20756,N_20041);
nor U21574 (N_21574,N_20849,N_20993);
nand U21575 (N_21575,N_20708,N_20241);
and U21576 (N_21576,N_20187,N_20163);
nor U21577 (N_21577,N_20233,N_20105);
and U21578 (N_21578,N_20806,N_20909);
nor U21579 (N_21579,N_20975,N_20331);
or U21580 (N_21580,N_20861,N_20344);
nand U21581 (N_21581,N_20829,N_20043);
xnor U21582 (N_21582,N_20204,N_20187);
nor U21583 (N_21583,N_20296,N_20796);
nand U21584 (N_21584,N_20227,N_20214);
or U21585 (N_21585,N_20150,N_20732);
or U21586 (N_21586,N_20533,N_20968);
nor U21587 (N_21587,N_20290,N_20039);
and U21588 (N_21588,N_20580,N_20770);
xnor U21589 (N_21589,N_20268,N_20960);
xor U21590 (N_21590,N_20517,N_20362);
xnor U21591 (N_21591,N_20211,N_20077);
nor U21592 (N_21592,N_20947,N_20510);
or U21593 (N_21593,N_20630,N_20012);
and U21594 (N_21594,N_20959,N_20255);
and U21595 (N_21595,N_20894,N_20268);
nand U21596 (N_21596,N_20003,N_20378);
or U21597 (N_21597,N_20262,N_20456);
and U21598 (N_21598,N_20573,N_20455);
nor U21599 (N_21599,N_20076,N_20380);
and U21600 (N_21600,N_20351,N_20214);
nand U21601 (N_21601,N_20854,N_20622);
xor U21602 (N_21602,N_20400,N_20038);
xnor U21603 (N_21603,N_20684,N_20596);
or U21604 (N_21604,N_20705,N_20813);
nand U21605 (N_21605,N_20197,N_20627);
or U21606 (N_21606,N_20899,N_20588);
nand U21607 (N_21607,N_20304,N_20397);
nor U21608 (N_21608,N_20170,N_20183);
nor U21609 (N_21609,N_20537,N_20277);
nand U21610 (N_21610,N_20236,N_20485);
xor U21611 (N_21611,N_20246,N_20401);
xor U21612 (N_21612,N_20448,N_20052);
xnor U21613 (N_21613,N_20225,N_20919);
nor U21614 (N_21614,N_20124,N_20098);
nor U21615 (N_21615,N_20155,N_20358);
xnor U21616 (N_21616,N_20644,N_20702);
xor U21617 (N_21617,N_20741,N_20853);
and U21618 (N_21618,N_20417,N_20364);
or U21619 (N_21619,N_20395,N_20103);
or U21620 (N_21620,N_20374,N_20271);
xor U21621 (N_21621,N_20861,N_20193);
or U21622 (N_21622,N_20752,N_20860);
xor U21623 (N_21623,N_20581,N_20879);
nor U21624 (N_21624,N_20378,N_20698);
or U21625 (N_21625,N_20537,N_20670);
xor U21626 (N_21626,N_20112,N_20463);
or U21627 (N_21627,N_20077,N_20318);
xnor U21628 (N_21628,N_20048,N_20469);
nor U21629 (N_21629,N_20425,N_20607);
and U21630 (N_21630,N_20115,N_20907);
or U21631 (N_21631,N_20630,N_20058);
or U21632 (N_21632,N_20411,N_20087);
or U21633 (N_21633,N_20112,N_20941);
xnor U21634 (N_21634,N_20193,N_20154);
or U21635 (N_21635,N_20535,N_20117);
nand U21636 (N_21636,N_20785,N_20825);
nor U21637 (N_21637,N_20165,N_20329);
nand U21638 (N_21638,N_20416,N_20157);
and U21639 (N_21639,N_20737,N_20693);
nand U21640 (N_21640,N_20460,N_20952);
xnor U21641 (N_21641,N_20589,N_20367);
nor U21642 (N_21642,N_20158,N_20218);
or U21643 (N_21643,N_20388,N_20788);
and U21644 (N_21644,N_20926,N_20300);
or U21645 (N_21645,N_20969,N_20208);
xnor U21646 (N_21646,N_20030,N_20826);
or U21647 (N_21647,N_20664,N_20119);
xor U21648 (N_21648,N_20594,N_20231);
or U21649 (N_21649,N_20685,N_20938);
xnor U21650 (N_21650,N_20327,N_20777);
or U21651 (N_21651,N_20885,N_20288);
nand U21652 (N_21652,N_20573,N_20982);
nor U21653 (N_21653,N_20838,N_20933);
nor U21654 (N_21654,N_20229,N_20148);
and U21655 (N_21655,N_20346,N_20052);
or U21656 (N_21656,N_20741,N_20631);
nand U21657 (N_21657,N_20098,N_20892);
or U21658 (N_21658,N_20034,N_20046);
nor U21659 (N_21659,N_20215,N_20577);
nand U21660 (N_21660,N_20959,N_20134);
or U21661 (N_21661,N_20162,N_20418);
and U21662 (N_21662,N_20022,N_20430);
nor U21663 (N_21663,N_20526,N_20291);
xnor U21664 (N_21664,N_20075,N_20360);
or U21665 (N_21665,N_20753,N_20740);
nand U21666 (N_21666,N_20039,N_20206);
and U21667 (N_21667,N_20322,N_20224);
or U21668 (N_21668,N_20057,N_20450);
xor U21669 (N_21669,N_20692,N_20690);
nor U21670 (N_21670,N_20523,N_20480);
nand U21671 (N_21671,N_20639,N_20299);
and U21672 (N_21672,N_20677,N_20552);
or U21673 (N_21673,N_20545,N_20890);
or U21674 (N_21674,N_20779,N_20454);
or U21675 (N_21675,N_20697,N_20371);
or U21676 (N_21676,N_20578,N_20889);
nor U21677 (N_21677,N_20538,N_20968);
or U21678 (N_21678,N_20802,N_20550);
or U21679 (N_21679,N_20295,N_20088);
nor U21680 (N_21680,N_20587,N_20964);
and U21681 (N_21681,N_20464,N_20118);
nand U21682 (N_21682,N_20754,N_20730);
nand U21683 (N_21683,N_20167,N_20213);
nor U21684 (N_21684,N_20521,N_20868);
and U21685 (N_21685,N_20538,N_20287);
and U21686 (N_21686,N_20006,N_20849);
and U21687 (N_21687,N_20279,N_20733);
xor U21688 (N_21688,N_20153,N_20969);
nor U21689 (N_21689,N_20579,N_20234);
nand U21690 (N_21690,N_20509,N_20350);
nor U21691 (N_21691,N_20231,N_20311);
nand U21692 (N_21692,N_20673,N_20885);
xor U21693 (N_21693,N_20065,N_20805);
xnor U21694 (N_21694,N_20032,N_20097);
nor U21695 (N_21695,N_20217,N_20798);
and U21696 (N_21696,N_20613,N_20795);
nor U21697 (N_21697,N_20275,N_20626);
xnor U21698 (N_21698,N_20989,N_20197);
and U21699 (N_21699,N_20169,N_20050);
and U21700 (N_21700,N_20953,N_20748);
or U21701 (N_21701,N_20245,N_20246);
xor U21702 (N_21702,N_20678,N_20626);
and U21703 (N_21703,N_20500,N_20721);
nand U21704 (N_21704,N_20988,N_20205);
or U21705 (N_21705,N_20154,N_20533);
xor U21706 (N_21706,N_20041,N_20382);
and U21707 (N_21707,N_20820,N_20837);
xnor U21708 (N_21708,N_20996,N_20304);
or U21709 (N_21709,N_20965,N_20609);
nor U21710 (N_21710,N_20858,N_20606);
xnor U21711 (N_21711,N_20939,N_20845);
and U21712 (N_21712,N_20396,N_20887);
xnor U21713 (N_21713,N_20004,N_20126);
xor U21714 (N_21714,N_20432,N_20660);
nor U21715 (N_21715,N_20483,N_20999);
nor U21716 (N_21716,N_20176,N_20171);
nand U21717 (N_21717,N_20125,N_20039);
xnor U21718 (N_21718,N_20482,N_20320);
and U21719 (N_21719,N_20290,N_20322);
or U21720 (N_21720,N_20978,N_20480);
and U21721 (N_21721,N_20390,N_20212);
nand U21722 (N_21722,N_20034,N_20097);
xor U21723 (N_21723,N_20880,N_20711);
xnor U21724 (N_21724,N_20308,N_20068);
or U21725 (N_21725,N_20685,N_20256);
xnor U21726 (N_21726,N_20521,N_20744);
or U21727 (N_21727,N_20236,N_20421);
xor U21728 (N_21728,N_20013,N_20646);
nor U21729 (N_21729,N_20272,N_20262);
xnor U21730 (N_21730,N_20099,N_20410);
nor U21731 (N_21731,N_20311,N_20676);
nor U21732 (N_21732,N_20736,N_20872);
nor U21733 (N_21733,N_20570,N_20198);
nor U21734 (N_21734,N_20524,N_20314);
xor U21735 (N_21735,N_20494,N_20312);
or U21736 (N_21736,N_20817,N_20072);
xor U21737 (N_21737,N_20779,N_20122);
nand U21738 (N_21738,N_20539,N_20907);
or U21739 (N_21739,N_20538,N_20396);
and U21740 (N_21740,N_20920,N_20726);
or U21741 (N_21741,N_20755,N_20131);
or U21742 (N_21742,N_20188,N_20574);
or U21743 (N_21743,N_20540,N_20908);
or U21744 (N_21744,N_20954,N_20606);
nor U21745 (N_21745,N_20229,N_20765);
nand U21746 (N_21746,N_20962,N_20158);
xor U21747 (N_21747,N_20059,N_20051);
nand U21748 (N_21748,N_20720,N_20030);
or U21749 (N_21749,N_20240,N_20887);
nor U21750 (N_21750,N_20523,N_20105);
nand U21751 (N_21751,N_20983,N_20014);
nor U21752 (N_21752,N_20495,N_20755);
or U21753 (N_21753,N_20716,N_20659);
and U21754 (N_21754,N_20445,N_20117);
xor U21755 (N_21755,N_20757,N_20098);
nor U21756 (N_21756,N_20453,N_20183);
and U21757 (N_21757,N_20580,N_20392);
nand U21758 (N_21758,N_20354,N_20610);
xor U21759 (N_21759,N_20138,N_20484);
and U21760 (N_21760,N_20278,N_20764);
nand U21761 (N_21761,N_20870,N_20503);
and U21762 (N_21762,N_20907,N_20615);
nor U21763 (N_21763,N_20311,N_20886);
nor U21764 (N_21764,N_20305,N_20439);
nor U21765 (N_21765,N_20962,N_20792);
nor U21766 (N_21766,N_20417,N_20145);
nor U21767 (N_21767,N_20212,N_20284);
nor U21768 (N_21768,N_20337,N_20095);
or U21769 (N_21769,N_20746,N_20988);
nand U21770 (N_21770,N_20239,N_20262);
xor U21771 (N_21771,N_20262,N_20773);
xnor U21772 (N_21772,N_20194,N_20776);
or U21773 (N_21773,N_20073,N_20390);
or U21774 (N_21774,N_20611,N_20225);
and U21775 (N_21775,N_20730,N_20328);
nor U21776 (N_21776,N_20628,N_20076);
and U21777 (N_21777,N_20898,N_20714);
nand U21778 (N_21778,N_20608,N_20009);
nor U21779 (N_21779,N_20981,N_20967);
and U21780 (N_21780,N_20710,N_20903);
and U21781 (N_21781,N_20557,N_20089);
and U21782 (N_21782,N_20346,N_20259);
and U21783 (N_21783,N_20027,N_20324);
xnor U21784 (N_21784,N_20202,N_20027);
nor U21785 (N_21785,N_20663,N_20059);
nor U21786 (N_21786,N_20633,N_20374);
or U21787 (N_21787,N_20888,N_20208);
or U21788 (N_21788,N_20253,N_20003);
nand U21789 (N_21789,N_20887,N_20153);
nor U21790 (N_21790,N_20348,N_20483);
and U21791 (N_21791,N_20960,N_20568);
and U21792 (N_21792,N_20672,N_20139);
or U21793 (N_21793,N_20800,N_20572);
or U21794 (N_21794,N_20166,N_20840);
nand U21795 (N_21795,N_20133,N_20508);
or U21796 (N_21796,N_20885,N_20931);
and U21797 (N_21797,N_20393,N_20754);
xnor U21798 (N_21798,N_20415,N_20214);
nor U21799 (N_21799,N_20961,N_20596);
or U21800 (N_21800,N_20706,N_20064);
or U21801 (N_21801,N_20537,N_20340);
nand U21802 (N_21802,N_20363,N_20540);
nand U21803 (N_21803,N_20531,N_20418);
nand U21804 (N_21804,N_20715,N_20296);
or U21805 (N_21805,N_20342,N_20633);
xnor U21806 (N_21806,N_20119,N_20857);
or U21807 (N_21807,N_20512,N_20942);
nor U21808 (N_21808,N_20882,N_20829);
and U21809 (N_21809,N_20251,N_20252);
or U21810 (N_21810,N_20766,N_20326);
and U21811 (N_21811,N_20913,N_20473);
and U21812 (N_21812,N_20986,N_20353);
or U21813 (N_21813,N_20863,N_20795);
and U21814 (N_21814,N_20947,N_20908);
nand U21815 (N_21815,N_20157,N_20075);
or U21816 (N_21816,N_20186,N_20563);
xnor U21817 (N_21817,N_20220,N_20309);
nand U21818 (N_21818,N_20330,N_20531);
and U21819 (N_21819,N_20303,N_20149);
nand U21820 (N_21820,N_20704,N_20359);
xnor U21821 (N_21821,N_20651,N_20127);
nand U21822 (N_21822,N_20699,N_20271);
and U21823 (N_21823,N_20276,N_20635);
nand U21824 (N_21824,N_20198,N_20312);
or U21825 (N_21825,N_20584,N_20157);
xnor U21826 (N_21826,N_20855,N_20613);
or U21827 (N_21827,N_20477,N_20386);
and U21828 (N_21828,N_20864,N_20661);
xnor U21829 (N_21829,N_20038,N_20290);
nor U21830 (N_21830,N_20840,N_20150);
nand U21831 (N_21831,N_20029,N_20037);
nand U21832 (N_21832,N_20370,N_20392);
nand U21833 (N_21833,N_20796,N_20134);
and U21834 (N_21834,N_20896,N_20003);
or U21835 (N_21835,N_20672,N_20740);
xor U21836 (N_21836,N_20745,N_20963);
and U21837 (N_21837,N_20177,N_20804);
nor U21838 (N_21838,N_20462,N_20515);
and U21839 (N_21839,N_20471,N_20226);
xnor U21840 (N_21840,N_20666,N_20884);
xnor U21841 (N_21841,N_20623,N_20931);
nor U21842 (N_21842,N_20712,N_20170);
and U21843 (N_21843,N_20234,N_20189);
nor U21844 (N_21844,N_20307,N_20238);
nor U21845 (N_21845,N_20573,N_20468);
or U21846 (N_21846,N_20310,N_20874);
nor U21847 (N_21847,N_20531,N_20962);
or U21848 (N_21848,N_20752,N_20443);
and U21849 (N_21849,N_20781,N_20908);
or U21850 (N_21850,N_20817,N_20076);
xnor U21851 (N_21851,N_20805,N_20169);
nand U21852 (N_21852,N_20926,N_20587);
and U21853 (N_21853,N_20897,N_20199);
and U21854 (N_21854,N_20983,N_20933);
xor U21855 (N_21855,N_20685,N_20352);
or U21856 (N_21856,N_20517,N_20678);
xor U21857 (N_21857,N_20852,N_20396);
nor U21858 (N_21858,N_20041,N_20597);
and U21859 (N_21859,N_20653,N_20461);
nor U21860 (N_21860,N_20407,N_20735);
xnor U21861 (N_21861,N_20649,N_20713);
or U21862 (N_21862,N_20089,N_20425);
xnor U21863 (N_21863,N_20276,N_20284);
nor U21864 (N_21864,N_20711,N_20169);
nor U21865 (N_21865,N_20846,N_20837);
nand U21866 (N_21866,N_20809,N_20937);
nor U21867 (N_21867,N_20744,N_20895);
or U21868 (N_21868,N_20120,N_20482);
or U21869 (N_21869,N_20839,N_20952);
nand U21870 (N_21870,N_20330,N_20525);
xor U21871 (N_21871,N_20553,N_20478);
and U21872 (N_21872,N_20900,N_20916);
nand U21873 (N_21873,N_20113,N_20586);
nand U21874 (N_21874,N_20010,N_20616);
and U21875 (N_21875,N_20208,N_20050);
nand U21876 (N_21876,N_20044,N_20434);
or U21877 (N_21877,N_20186,N_20437);
and U21878 (N_21878,N_20069,N_20549);
or U21879 (N_21879,N_20239,N_20349);
xor U21880 (N_21880,N_20363,N_20258);
or U21881 (N_21881,N_20876,N_20937);
nor U21882 (N_21882,N_20364,N_20903);
nor U21883 (N_21883,N_20436,N_20229);
nand U21884 (N_21884,N_20635,N_20382);
nor U21885 (N_21885,N_20260,N_20217);
and U21886 (N_21886,N_20598,N_20895);
or U21887 (N_21887,N_20660,N_20068);
nor U21888 (N_21888,N_20888,N_20170);
and U21889 (N_21889,N_20844,N_20772);
nor U21890 (N_21890,N_20658,N_20429);
nor U21891 (N_21891,N_20422,N_20442);
and U21892 (N_21892,N_20603,N_20712);
and U21893 (N_21893,N_20657,N_20635);
and U21894 (N_21894,N_20416,N_20104);
or U21895 (N_21895,N_20064,N_20744);
xnor U21896 (N_21896,N_20863,N_20742);
xor U21897 (N_21897,N_20871,N_20125);
nor U21898 (N_21898,N_20574,N_20995);
xor U21899 (N_21899,N_20889,N_20363);
or U21900 (N_21900,N_20909,N_20915);
nand U21901 (N_21901,N_20861,N_20453);
nor U21902 (N_21902,N_20428,N_20391);
nor U21903 (N_21903,N_20190,N_20952);
or U21904 (N_21904,N_20217,N_20724);
or U21905 (N_21905,N_20619,N_20518);
and U21906 (N_21906,N_20686,N_20235);
nand U21907 (N_21907,N_20089,N_20272);
and U21908 (N_21908,N_20022,N_20876);
xnor U21909 (N_21909,N_20252,N_20702);
nand U21910 (N_21910,N_20767,N_20324);
nor U21911 (N_21911,N_20056,N_20657);
xnor U21912 (N_21912,N_20496,N_20289);
xor U21913 (N_21913,N_20342,N_20888);
nor U21914 (N_21914,N_20634,N_20462);
xnor U21915 (N_21915,N_20012,N_20158);
nand U21916 (N_21916,N_20067,N_20232);
or U21917 (N_21917,N_20643,N_20654);
nor U21918 (N_21918,N_20400,N_20332);
nand U21919 (N_21919,N_20008,N_20491);
nand U21920 (N_21920,N_20414,N_20363);
nand U21921 (N_21921,N_20901,N_20151);
nand U21922 (N_21922,N_20778,N_20525);
or U21923 (N_21923,N_20267,N_20253);
or U21924 (N_21924,N_20202,N_20812);
xor U21925 (N_21925,N_20390,N_20682);
or U21926 (N_21926,N_20824,N_20163);
xor U21927 (N_21927,N_20034,N_20991);
nor U21928 (N_21928,N_20569,N_20665);
nor U21929 (N_21929,N_20078,N_20001);
nor U21930 (N_21930,N_20748,N_20282);
and U21931 (N_21931,N_20984,N_20673);
or U21932 (N_21932,N_20691,N_20334);
xnor U21933 (N_21933,N_20800,N_20108);
xnor U21934 (N_21934,N_20504,N_20419);
or U21935 (N_21935,N_20991,N_20290);
nand U21936 (N_21936,N_20672,N_20805);
nand U21937 (N_21937,N_20311,N_20029);
nor U21938 (N_21938,N_20878,N_20583);
and U21939 (N_21939,N_20279,N_20606);
nor U21940 (N_21940,N_20949,N_20112);
nand U21941 (N_21941,N_20002,N_20049);
xor U21942 (N_21942,N_20081,N_20603);
nor U21943 (N_21943,N_20795,N_20720);
xor U21944 (N_21944,N_20233,N_20920);
and U21945 (N_21945,N_20801,N_20303);
xor U21946 (N_21946,N_20280,N_20453);
and U21947 (N_21947,N_20508,N_20328);
xnor U21948 (N_21948,N_20790,N_20981);
or U21949 (N_21949,N_20044,N_20073);
and U21950 (N_21950,N_20228,N_20408);
xnor U21951 (N_21951,N_20422,N_20513);
or U21952 (N_21952,N_20790,N_20352);
nor U21953 (N_21953,N_20596,N_20053);
nor U21954 (N_21954,N_20766,N_20728);
or U21955 (N_21955,N_20334,N_20256);
xor U21956 (N_21956,N_20882,N_20952);
xnor U21957 (N_21957,N_20426,N_20852);
and U21958 (N_21958,N_20521,N_20146);
nand U21959 (N_21959,N_20568,N_20418);
nor U21960 (N_21960,N_20851,N_20499);
xor U21961 (N_21961,N_20225,N_20122);
nor U21962 (N_21962,N_20083,N_20991);
or U21963 (N_21963,N_20466,N_20166);
nand U21964 (N_21964,N_20399,N_20356);
nor U21965 (N_21965,N_20275,N_20202);
nand U21966 (N_21966,N_20459,N_20192);
or U21967 (N_21967,N_20515,N_20099);
and U21968 (N_21968,N_20063,N_20511);
or U21969 (N_21969,N_20044,N_20009);
or U21970 (N_21970,N_20063,N_20962);
nand U21971 (N_21971,N_20103,N_20895);
xor U21972 (N_21972,N_20130,N_20156);
and U21973 (N_21973,N_20903,N_20091);
and U21974 (N_21974,N_20924,N_20988);
nand U21975 (N_21975,N_20322,N_20878);
nor U21976 (N_21976,N_20457,N_20972);
and U21977 (N_21977,N_20890,N_20869);
and U21978 (N_21978,N_20751,N_20485);
nor U21979 (N_21979,N_20523,N_20306);
and U21980 (N_21980,N_20712,N_20759);
nand U21981 (N_21981,N_20883,N_20810);
or U21982 (N_21982,N_20586,N_20119);
nand U21983 (N_21983,N_20685,N_20017);
and U21984 (N_21984,N_20128,N_20604);
nand U21985 (N_21985,N_20641,N_20121);
or U21986 (N_21986,N_20032,N_20424);
xor U21987 (N_21987,N_20003,N_20991);
or U21988 (N_21988,N_20036,N_20617);
xor U21989 (N_21989,N_20952,N_20377);
or U21990 (N_21990,N_20516,N_20070);
or U21991 (N_21991,N_20622,N_20376);
or U21992 (N_21992,N_20134,N_20463);
nand U21993 (N_21993,N_20462,N_20712);
or U21994 (N_21994,N_20827,N_20654);
or U21995 (N_21995,N_20830,N_20819);
nand U21996 (N_21996,N_20502,N_20757);
or U21997 (N_21997,N_20051,N_20794);
or U21998 (N_21998,N_20173,N_20346);
xor U21999 (N_21999,N_20520,N_20479);
and U22000 (N_22000,N_21292,N_21597);
nor U22001 (N_22001,N_21942,N_21699);
nor U22002 (N_22002,N_21009,N_21188);
and U22003 (N_22003,N_21420,N_21667);
xnor U22004 (N_22004,N_21720,N_21209);
nand U22005 (N_22005,N_21776,N_21178);
nor U22006 (N_22006,N_21523,N_21074);
nand U22007 (N_22007,N_21618,N_21885);
xnor U22008 (N_22008,N_21746,N_21498);
and U22009 (N_22009,N_21644,N_21829);
or U22010 (N_22010,N_21671,N_21494);
nor U22011 (N_22011,N_21750,N_21412);
nor U22012 (N_22012,N_21019,N_21106);
or U22013 (N_22013,N_21775,N_21172);
xor U22014 (N_22014,N_21300,N_21793);
xnor U22015 (N_22015,N_21993,N_21779);
nor U22016 (N_22016,N_21854,N_21262);
or U22017 (N_22017,N_21575,N_21410);
nand U22018 (N_22018,N_21033,N_21700);
or U22019 (N_22019,N_21390,N_21433);
xor U22020 (N_22020,N_21072,N_21913);
nor U22021 (N_22021,N_21249,N_21588);
xor U22022 (N_22022,N_21217,N_21109);
nand U22023 (N_22023,N_21992,N_21722);
or U22024 (N_22024,N_21623,N_21266);
nor U22025 (N_22025,N_21634,N_21711);
and U22026 (N_22026,N_21616,N_21935);
and U22027 (N_22027,N_21124,N_21245);
nor U22028 (N_22028,N_21731,N_21446);
xor U22029 (N_22029,N_21269,N_21396);
or U22030 (N_22030,N_21626,N_21367);
nand U22031 (N_22031,N_21451,N_21825);
nand U22032 (N_22032,N_21368,N_21151);
nand U22033 (N_22033,N_21280,N_21701);
or U22034 (N_22034,N_21631,N_21277);
nand U22035 (N_22035,N_21100,N_21838);
nand U22036 (N_22036,N_21159,N_21540);
or U22037 (N_22037,N_21984,N_21956);
or U22038 (N_22038,N_21195,N_21444);
nand U22039 (N_22039,N_21757,N_21022);
and U22040 (N_22040,N_21661,N_21924);
nand U22041 (N_22041,N_21107,N_21806);
or U22042 (N_22042,N_21371,N_21117);
nand U22043 (N_22043,N_21201,N_21818);
and U22044 (N_22044,N_21828,N_21902);
xnor U22045 (N_22045,N_21313,N_21718);
or U22046 (N_22046,N_21627,N_21353);
xnor U22047 (N_22047,N_21325,N_21813);
and U22048 (N_22048,N_21372,N_21286);
or U22049 (N_22049,N_21666,N_21729);
nor U22050 (N_22050,N_21120,N_21311);
and U22051 (N_22051,N_21535,N_21798);
xnor U22052 (N_22052,N_21977,N_21214);
nand U22053 (N_22053,N_21105,N_21415);
or U22054 (N_22054,N_21573,N_21783);
and U22055 (N_22055,N_21293,N_21321);
nor U22056 (N_22056,N_21594,N_21734);
xor U22057 (N_22057,N_21877,N_21872);
nor U22058 (N_22058,N_21721,N_21336);
xnor U22059 (N_22059,N_21108,N_21726);
xor U22060 (N_22060,N_21794,N_21570);
nand U22061 (N_22061,N_21708,N_21119);
xor U22062 (N_22062,N_21263,N_21436);
xor U22063 (N_22063,N_21492,N_21237);
nand U22064 (N_22064,N_21789,N_21118);
nor U22065 (N_22065,N_21154,N_21955);
nor U22066 (N_22066,N_21144,N_21974);
or U22067 (N_22067,N_21850,N_21847);
nor U22068 (N_22068,N_21760,N_21181);
or U22069 (N_22069,N_21128,N_21373);
nor U22070 (N_22070,N_21799,N_21474);
or U22071 (N_22071,N_21926,N_21542);
nand U22072 (N_22072,N_21682,N_21347);
and U22073 (N_22073,N_21018,N_21925);
and U22074 (N_22074,N_21255,N_21274);
xnor U22075 (N_22075,N_21233,N_21878);
xnor U22076 (N_22076,N_21511,N_21933);
or U22077 (N_22077,N_21267,N_21259);
and U22078 (N_22078,N_21569,N_21442);
or U22079 (N_22079,N_21213,N_21904);
nor U22080 (N_22080,N_21579,N_21907);
nor U22081 (N_22081,N_21330,N_21378);
and U22082 (N_22082,N_21075,N_21512);
nor U22083 (N_22083,N_21753,N_21026);
nand U22084 (N_22084,N_21554,N_21581);
or U22085 (N_22085,N_21969,N_21002);
nand U22086 (N_22086,N_21923,N_21463);
or U22087 (N_22087,N_21989,N_21884);
nand U22088 (N_22088,N_21205,N_21479);
nor U22089 (N_22089,N_21624,N_21745);
xnor U22090 (N_22090,N_21168,N_21417);
and U22091 (N_22091,N_21865,N_21583);
and U22092 (N_22092,N_21123,N_21524);
and U22093 (N_22093,N_21858,N_21224);
or U22094 (N_22094,N_21082,N_21180);
xnor U22095 (N_22095,N_21244,N_21797);
nor U22096 (N_22096,N_21846,N_21148);
xnor U22097 (N_22097,N_21495,N_21790);
xor U22098 (N_22098,N_21186,N_21355);
nand U22099 (N_22099,N_21756,N_21228);
nand U22100 (N_22100,N_21338,N_21025);
and U22101 (N_22101,N_21413,N_21045);
nand U22102 (N_22102,N_21149,N_21312);
and U22103 (N_22103,N_21778,N_21086);
nand U22104 (N_22104,N_21003,N_21152);
xor U22105 (N_22105,N_21946,N_21703);
xor U22106 (N_22106,N_21896,N_21239);
and U22107 (N_22107,N_21749,N_21342);
and U22108 (N_22108,N_21248,N_21717);
xnor U22109 (N_22109,N_21845,N_21559);
or U22110 (N_22110,N_21365,N_21894);
or U22111 (N_22111,N_21707,N_21005);
or U22112 (N_22112,N_21963,N_21219);
nor U22113 (N_22113,N_21546,N_21648);
or U22114 (N_22114,N_21678,N_21329);
or U22115 (N_22115,N_21875,N_21948);
xnor U22116 (N_22116,N_21081,N_21744);
and U22117 (N_22117,N_21695,N_21835);
or U22118 (N_22118,N_21027,N_21384);
and U22119 (N_22119,N_21339,N_21400);
or U22120 (N_22120,N_21472,N_21632);
or U22121 (N_22121,N_21654,N_21556);
nor U22122 (N_22122,N_21506,N_21918);
nand U22123 (N_22123,N_21997,N_21039);
nand U22124 (N_22124,N_21608,N_21537);
nor U22125 (N_22125,N_21803,N_21890);
and U22126 (N_22126,N_21099,N_21131);
nor U22127 (N_22127,N_21096,N_21246);
and U22128 (N_22128,N_21408,N_21965);
or U22129 (N_22129,N_21403,N_21053);
nor U22130 (N_22130,N_21958,N_21391);
nand U22131 (N_22131,N_21021,N_21879);
and U22132 (N_22132,N_21089,N_21059);
xor U22133 (N_22133,N_21723,N_21743);
or U22134 (N_22134,N_21903,N_21202);
or U22135 (N_22135,N_21370,N_21261);
and U22136 (N_22136,N_21522,N_21880);
nor U22137 (N_22137,N_21669,N_21136);
xor U22138 (N_22138,N_21194,N_21649);
nor U22139 (N_22139,N_21250,N_21369);
and U22140 (N_22140,N_21761,N_21138);
and U22141 (N_22141,N_21621,N_21358);
xnor U22142 (N_22142,N_21434,N_21668);
nor U22143 (N_22143,N_21464,N_21399);
xnor U22144 (N_22144,N_21834,N_21304);
and U22145 (N_22145,N_21327,N_21066);
nand U22146 (N_22146,N_21628,N_21121);
xor U22147 (N_22147,N_21314,N_21445);
nand U22148 (N_22148,N_21111,N_21203);
nor U22149 (N_22149,N_21625,N_21160);
and U22150 (N_22150,N_21802,N_21603);
nand U22151 (N_22151,N_21298,N_21919);
nor U22152 (N_22152,N_21502,N_21855);
nor U22153 (N_22153,N_21576,N_21754);
xnor U22154 (N_22154,N_21752,N_21476);
xor U22155 (N_22155,N_21218,N_21165);
nand U22156 (N_22156,N_21662,N_21816);
nor U22157 (N_22157,N_21742,N_21527);
nor U22158 (N_22158,N_21590,N_21437);
nand U22159 (N_22159,N_21031,N_21518);
or U22160 (N_22160,N_21422,N_21360);
nor U22161 (N_22161,N_21837,N_21363);
or U22162 (N_22162,N_21773,N_21866);
nor U22163 (N_22163,N_21538,N_21411);
nand U22164 (N_22164,N_21094,N_21792);
and U22165 (N_22165,N_21796,N_21548);
and U22166 (N_22166,N_21056,N_21823);
xor U22167 (N_22167,N_21800,N_21841);
or U22168 (N_22168,N_21097,N_21225);
or U22169 (N_22169,N_21780,N_21606);
or U22170 (N_22170,N_21937,N_21898);
and U22171 (N_22171,N_21819,N_21596);
or U22172 (N_22172,N_21281,N_21282);
nand U22173 (N_22173,N_21959,N_21764);
nand U22174 (N_22174,N_21859,N_21092);
nand U22175 (N_22175,N_21392,N_21715);
or U22176 (N_22176,N_21230,N_21012);
nand U22177 (N_22177,N_21612,N_21781);
xnor U22178 (N_22178,N_21448,N_21714);
or U22179 (N_22179,N_21060,N_21565);
nor U22180 (N_22180,N_21602,N_21449);
xnor U22181 (N_22181,N_21014,N_21968);
nand U22182 (N_22182,N_21470,N_21572);
nor U22183 (N_22183,N_21447,N_21348);
and U22184 (N_22184,N_21036,N_21155);
nand U22185 (N_22185,N_21197,N_21510);
and U22186 (N_22186,N_21461,N_21943);
and U22187 (N_22187,N_21740,N_21157);
nand U22188 (N_22188,N_21050,N_21784);
xnor U22189 (N_22189,N_21455,N_21536);
nand U22190 (N_22190,N_21112,N_21862);
nand U22191 (N_22191,N_21677,N_21385);
nand U22192 (N_22192,N_21211,N_21851);
nor U22193 (N_22193,N_21759,N_21465);
nor U22194 (N_22194,N_21234,N_21983);
and U22195 (N_22195,N_21947,N_21600);
or U22196 (N_22196,N_21636,N_21207);
nand U22197 (N_22197,N_21078,N_21037);
and U22198 (N_22198,N_21728,N_21807);
nor U22199 (N_22199,N_21619,N_21083);
and U22200 (N_22200,N_21297,N_21689);
xnor U22201 (N_22201,N_21639,N_21839);
nor U22202 (N_22202,N_21638,N_21549);
and U22203 (N_22203,N_21438,N_21712);
nand U22204 (N_22204,N_21652,N_21566);
or U22205 (N_22205,N_21737,N_21599);
nand U22206 (N_22206,N_21308,N_21589);
xor U22207 (N_22207,N_21024,N_21592);
nand U22208 (N_22208,N_21071,N_21344);
xor U22209 (N_22209,N_21539,N_21762);
xor U22210 (N_22210,N_21189,N_21307);
and U22211 (N_22211,N_21088,N_21204);
and U22212 (N_22212,N_21271,N_21115);
or U22213 (N_22213,N_21405,N_21317);
nor U22214 (N_22214,N_21440,N_21132);
or U22215 (N_22215,N_21299,N_21683);
nand U22216 (N_22216,N_21167,N_21232);
nand U22217 (N_22217,N_21273,N_21952);
xnor U22218 (N_22218,N_21966,N_21485);
and U22219 (N_22219,N_21134,N_21508);
and U22220 (N_22220,N_21268,N_21226);
nor U22221 (N_22221,N_21139,N_21331);
xnor U22222 (N_22222,N_21379,N_21670);
nand U22223 (N_22223,N_21135,N_21484);
or U22224 (N_22224,N_21931,N_21051);
xor U22225 (N_22225,N_21200,N_21285);
or U22226 (N_22226,N_21541,N_21503);
xnor U22227 (N_22227,N_21453,N_21376);
or U22228 (N_22228,N_21179,N_21477);
xor U22229 (N_22229,N_21725,N_21030);
and U22230 (N_22230,N_21543,N_21916);
xnor U22231 (N_22231,N_21288,N_21557);
nand U22232 (N_22232,N_21430,N_21719);
nand U22233 (N_22233,N_21156,N_21999);
and U22234 (N_22234,N_21316,N_21911);
nor U22235 (N_22235,N_21545,N_21694);
xnor U22236 (N_22236,N_21852,N_21673);
or U22237 (N_22237,N_21345,N_21637);
nand U22238 (N_22238,N_21227,N_21318);
or U22239 (N_22239,N_21733,N_21150);
nand U22240 (N_22240,N_21945,N_21551);
and U22241 (N_22241,N_21795,N_21251);
or U22242 (N_22242,N_21509,N_21801);
nand U22243 (N_22243,N_21844,N_21236);
nand U22244 (N_22244,N_21920,N_21362);
and U22245 (N_22245,N_21452,N_21961);
nand U22246 (N_22246,N_21651,N_21062);
or U22247 (N_22247,N_21295,N_21532);
nor U22248 (N_22248,N_21352,N_21486);
xor U22249 (N_22249,N_21777,N_21084);
xnor U22250 (N_22250,N_21291,N_21857);
nand U22251 (N_22251,N_21459,N_21450);
and U22252 (N_22252,N_21466,N_21040);
and U22253 (N_22253,N_21306,N_21874);
and U22254 (N_22254,N_21055,N_21769);
and U22255 (N_22255,N_21401,N_21986);
and U22256 (N_22256,N_21944,N_21264);
nor U22257 (N_22257,N_21864,N_21665);
and U22258 (N_22258,N_21351,N_21425);
and U22259 (N_22259,N_21791,N_21656);
xnor U22260 (N_22260,N_21553,N_21162);
nor U22261 (N_22261,N_21013,N_21895);
xor U22262 (N_22262,N_21967,N_21374);
nand U22263 (N_22263,N_21093,N_21125);
nor U22264 (N_22264,N_21070,N_21980);
nor U22265 (N_22265,N_21657,N_21229);
or U22266 (N_22266,N_21630,N_21861);
and U22267 (N_22267,N_21215,N_21531);
or U22268 (N_22268,N_21615,N_21960);
xor U22269 (N_22269,N_21870,N_21057);
nor U22270 (N_22270,N_21888,N_21614);
nand U22271 (N_22271,N_21685,N_21640);
xnor U22272 (N_22272,N_21921,N_21517);
xor U22273 (N_22273,N_21023,N_21755);
xnor U22274 (N_22274,N_21016,N_21418);
nand U22275 (N_22275,N_21361,N_21954);
and U22276 (N_22276,N_21130,N_21305);
or U22277 (N_22277,N_21617,N_21971);
nor U22278 (N_22278,N_21567,N_21810);
nor U22279 (N_22279,N_21595,N_21350);
xnor U22280 (N_22280,N_21017,N_21458);
or U22281 (N_22281,N_21198,N_21601);
or U22282 (N_22282,N_21586,N_21173);
and U22283 (N_22283,N_21951,N_21848);
nand U22284 (N_22284,N_21982,N_21141);
and U22285 (N_22285,N_21928,N_21061);
xor U22286 (N_22286,N_21253,N_21443);
nor U22287 (N_22287,N_21953,N_21521);
or U22288 (N_22288,N_21691,N_21513);
or U22289 (N_22289,N_21763,N_21891);
and U22290 (N_22290,N_21183,N_21635);
nor U22291 (N_22291,N_21876,N_21564);
nor U22292 (N_22292,N_21785,N_21140);
xor U22293 (N_22293,N_21552,N_21770);
or U22294 (N_22294,N_21525,N_21381);
or U22295 (N_22295,N_21515,N_21294);
xnor U22296 (N_22296,N_21990,N_21462);
nor U22297 (N_22297,N_21930,N_21704);
nor U22298 (N_22298,N_21278,N_21547);
and U22299 (N_22299,N_21126,N_21208);
and U22300 (N_22300,N_21964,N_21629);
or U22301 (N_22301,N_21998,N_21934);
nor U22302 (N_22302,N_21133,N_21067);
nor U22303 (N_22303,N_21110,N_21893);
nand U22304 (N_22304,N_21206,N_21320);
nand U22305 (N_22305,N_21221,N_21393);
nor U22306 (N_22306,N_21046,N_21697);
and U22307 (N_22307,N_21732,N_21315);
and U22308 (N_22308,N_21574,N_21398);
nor U22309 (N_22309,N_21970,N_21069);
nor U22310 (N_22310,N_21052,N_21301);
or U22311 (N_22311,N_21048,N_21011);
xor U22312 (N_22312,N_21558,N_21905);
xnor U22313 (N_22313,N_21840,N_21853);
nand U22314 (N_22314,N_21240,N_21912);
or U22315 (N_22315,N_21643,N_21812);
nand U22316 (N_22316,N_21426,N_21520);
nor U22317 (N_22317,N_21672,N_21469);
nand U22318 (N_22318,N_21129,N_21333);
and U22319 (N_22319,N_21058,N_21727);
and U22320 (N_22320,N_21471,N_21664);
and U22321 (N_22321,N_21786,N_21901);
xor U22322 (N_22322,N_21332,N_21222);
xor U22323 (N_22323,N_21482,N_21562);
or U22324 (N_22324,N_21402,N_21377);
or U22325 (N_22325,N_21193,N_21171);
xor U22326 (N_22326,N_21147,N_21758);
and U22327 (N_22327,N_21788,N_21272);
nand U22328 (N_22328,N_21578,N_21169);
xor U22329 (N_22329,N_21334,N_21686);
nor U22330 (N_22330,N_21354,N_21561);
nand U22331 (N_22331,N_21247,N_21483);
and U22332 (N_22332,N_21950,N_21421);
nand U22333 (N_22333,N_21199,N_21380);
and U22334 (N_22334,N_21153,N_21161);
nor U22335 (N_22335,N_21988,N_21473);
nor U22336 (N_22336,N_21191,N_21550);
nand U22337 (N_22337,N_21530,N_21319);
xor U22338 (N_22338,N_21979,N_21424);
or U22339 (N_22339,N_21241,N_21693);
nand U22340 (N_22340,N_21688,N_21283);
xor U22341 (N_22341,N_21808,N_21395);
or U22342 (N_22342,N_21481,N_21529);
and U22343 (N_22343,N_21177,N_21359);
nor U22344 (N_22344,N_21457,N_21035);
and U22345 (N_22345,N_21490,N_21647);
nand U22346 (N_22346,N_21220,N_21409);
nor U22347 (N_22347,N_21611,N_21653);
nand U22348 (N_22348,N_21768,N_21987);
or U22349 (N_22349,N_21054,N_21397);
or U22350 (N_22350,N_21419,N_21929);
and U22351 (N_22351,N_21642,N_21185);
nor U22352 (N_22352,N_21015,N_21079);
xor U22353 (N_22353,N_21416,N_21645);
nor U22354 (N_22354,N_21735,N_21235);
and U22355 (N_22355,N_21487,N_21975);
and U22356 (N_22356,N_21716,N_21713);
xnor U22357 (N_22357,N_21873,N_21568);
nor U22358 (N_22358,N_21910,N_21659);
and U22359 (N_22359,N_21076,N_21439);
and U22360 (N_22360,N_21322,N_21252);
nand U22361 (N_22361,N_21146,N_21504);
or U22362 (N_22362,N_21137,N_21279);
or U22363 (N_22363,N_21488,N_21063);
nand U22364 (N_22364,N_21533,N_21577);
nand U22365 (N_22365,N_21505,N_21815);
or U22366 (N_22366,N_21831,N_21309);
xor U22367 (N_22367,N_21692,N_21705);
and U22368 (N_22368,N_21406,N_21747);
nor U22369 (N_22369,N_21475,N_21932);
nor U22370 (N_22370,N_21607,N_21927);
nand U22371 (N_22371,N_21900,N_21323);
or U22372 (N_22372,N_21029,N_21454);
nand U22373 (N_22373,N_21674,N_21256);
or U22374 (N_22374,N_21526,N_21650);
or U22375 (N_22375,N_21748,N_21101);
nand U22376 (N_22376,N_21102,N_21499);
or U22377 (N_22377,N_21427,N_21480);
nor U22378 (N_22378,N_21867,N_21212);
and U22379 (N_22379,N_21343,N_21646);
xnor U22380 (N_22380,N_21043,N_21276);
nor U22381 (N_22381,N_21231,N_21922);
or U22382 (N_22382,N_21216,N_21468);
or U22383 (N_22383,N_21985,N_21836);
and U22384 (N_22384,N_21938,N_21897);
nand U22385 (N_22385,N_21571,N_21243);
nand U22386 (N_22386,N_21751,N_21658);
xor U22387 (N_22387,N_21114,N_21176);
nor U22388 (N_22388,N_21386,N_21698);
nand U22389 (N_22389,N_21098,N_21429);
xnor U22390 (N_22390,N_21145,N_21460);
xnor U22391 (N_22391,N_21337,N_21917);
nor U22392 (N_22392,N_21820,N_21899);
nor U22393 (N_22393,N_21028,N_21296);
and U22394 (N_22394,N_21184,N_21346);
nor U22395 (N_22395,N_21741,N_21767);
and U22396 (N_22396,N_21049,N_21387);
and U22397 (N_22397,N_21497,N_21765);
xnor U22398 (N_22398,N_21310,N_21257);
and U22399 (N_22399,N_21868,N_21001);
xor U22400 (N_22400,N_21340,N_21787);
or U22401 (N_22401,N_21441,N_21113);
and U22402 (N_22402,N_21882,N_21908);
nand U22403 (N_22403,N_21976,N_21388);
and U22404 (N_22404,N_21095,N_21881);
nand U22405 (N_22405,N_21302,N_21032);
and U22406 (N_22406,N_21906,N_21407);
or U22407 (N_22407,N_21706,N_21290);
nor U22408 (N_22408,N_21414,N_21004);
xor U22409 (N_22409,N_21771,N_21772);
and U22410 (N_22410,N_21260,N_21684);
nor U22411 (N_22411,N_21328,N_21843);
and U22412 (N_22412,N_21158,N_21604);
nand U22413 (N_22413,N_21182,N_21238);
xor U22414 (N_22414,N_21514,N_21814);
and U22415 (N_22415,N_21675,N_21432);
nand U22416 (N_22416,N_21860,N_21142);
and U22417 (N_22417,N_21357,N_21805);
or U22418 (N_22418,N_21680,N_21047);
nor U22419 (N_22419,N_21580,N_21341);
nand U22420 (N_22420,N_21914,N_21766);
and U22421 (N_22421,N_21507,N_21491);
and U22422 (N_22422,N_21613,N_21175);
and U22423 (N_22423,N_21994,N_21187);
nor U22424 (N_22424,N_21710,N_21609);
and U22425 (N_22425,N_21496,N_21270);
nor U22426 (N_22426,N_21830,N_21501);
nand U22427 (N_22427,N_21863,N_21622);
nand U22428 (N_22428,N_21641,N_21957);
nor U22429 (N_22429,N_21356,N_21389);
or U22430 (N_22430,N_21633,N_21655);
and U22431 (N_22431,N_21856,N_21824);
and U22432 (N_22432,N_21349,N_21822);
nor U22433 (N_22433,N_21324,N_21811);
or U22434 (N_22434,N_21516,N_21163);
and U22435 (N_22435,N_21493,N_21871);
or U22436 (N_22436,N_21949,N_21375);
nor U22437 (N_22437,N_21143,N_21679);
and U22438 (N_22438,N_21423,N_21724);
and U22439 (N_22439,N_21909,N_21832);
and U22440 (N_22440,N_21335,N_21326);
xnor U22441 (N_22441,N_21995,N_21041);
nand U22442 (N_22442,N_21582,N_21258);
nand U22443 (N_22443,N_21104,N_21289);
nand U22444 (N_22444,N_21842,N_21190);
or U22445 (N_22445,N_21736,N_21821);
xnor U22446 (N_22446,N_21489,N_21068);
xnor U22447 (N_22447,N_21660,N_21303);
and U22448 (N_22448,N_21170,N_21936);
nand U22449 (N_22449,N_21382,N_21103);
or U22450 (N_22450,N_21584,N_21038);
or U22451 (N_22451,N_21364,N_21940);
and U22452 (N_22452,N_21467,N_21404);
or U22453 (N_22453,N_21981,N_21431);
nand U22454 (N_22454,N_21738,N_21500);
nor U22455 (N_22455,N_21287,N_21702);
xnor U22456 (N_22456,N_21000,N_21833);
nor U22457 (N_22457,N_21774,N_21174);
nor U22458 (N_22458,N_21690,N_21883);
or U22459 (N_22459,N_21127,N_21192);
and U22460 (N_22460,N_21739,N_21696);
nor U22461 (N_22461,N_21366,N_21555);
xnor U22462 (N_22462,N_21428,N_21972);
or U22463 (N_22463,N_21978,N_21560);
nor U22464 (N_22464,N_21242,N_21534);
nor U22465 (N_22465,N_21122,N_21663);
nor U22466 (N_22466,N_21007,N_21605);
nand U22467 (N_22467,N_21887,N_21064);
and U22468 (N_22468,N_21210,N_21676);
and U22469 (N_22469,N_21010,N_21544);
and U22470 (N_22470,N_21610,N_21435);
xor U22471 (N_22471,N_21456,N_21585);
or U22472 (N_22472,N_21528,N_21709);
xor U22473 (N_22473,N_21827,N_21085);
and U22474 (N_22474,N_21962,N_21020);
xnor U22475 (N_22475,N_21782,N_21563);
or U22476 (N_22476,N_21196,N_21991);
nor U22477 (N_22477,N_21587,N_21090);
xor U22478 (N_22478,N_21265,N_21804);
xor U22479 (N_22479,N_21087,N_21166);
and U22480 (N_22480,N_21889,N_21091);
xor U22481 (N_22481,N_21006,N_21034);
and U22482 (N_22482,N_21080,N_21973);
nand U22483 (N_22483,N_21042,N_21116);
xnor U22484 (N_22484,N_21065,N_21008);
nor U22485 (N_22485,N_21164,N_21598);
and U22486 (N_22486,N_21478,N_21730);
and U22487 (N_22487,N_21223,N_21394);
xor U22488 (N_22488,N_21939,N_21254);
xor U22489 (N_22489,N_21275,N_21620);
nor U22490 (N_22490,N_21044,N_21809);
and U22491 (N_22491,N_21681,N_21996);
and U22492 (N_22492,N_21077,N_21826);
and U22493 (N_22493,N_21687,N_21915);
nor U22494 (N_22494,N_21886,N_21849);
nor U22495 (N_22495,N_21284,N_21892);
xnor U22496 (N_22496,N_21593,N_21869);
nand U22497 (N_22497,N_21383,N_21519);
xnor U22498 (N_22498,N_21817,N_21591);
or U22499 (N_22499,N_21073,N_21941);
nor U22500 (N_22500,N_21047,N_21787);
or U22501 (N_22501,N_21424,N_21697);
nand U22502 (N_22502,N_21441,N_21709);
or U22503 (N_22503,N_21767,N_21735);
xnor U22504 (N_22504,N_21086,N_21076);
xnor U22505 (N_22505,N_21338,N_21350);
or U22506 (N_22506,N_21709,N_21388);
and U22507 (N_22507,N_21239,N_21482);
or U22508 (N_22508,N_21882,N_21651);
nand U22509 (N_22509,N_21551,N_21350);
or U22510 (N_22510,N_21004,N_21392);
and U22511 (N_22511,N_21820,N_21996);
xnor U22512 (N_22512,N_21544,N_21049);
xor U22513 (N_22513,N_21453,N_21736);
or U22514 (N_22514,N_21548,N_21334);
nand U22515 (N_22515,N_21996,N_21028);
or U22516 (N_22516,N_21733,N_21818);
or U22517 (N_22517,N_21576,N_21364);
nor U22518 (N_22518,N_21010,N_21726);
and U22519 (N_22519,N_21103,N_21266);
or U22520 (N_22520,N_21750,N_21511);
nand U22521 (N_22521,N_21009,N_21549);
or U22522 (N_22522,N_21421,N_21711);
or U22523 (N_22523,N_21535,N_21627);
or U22524 (N_22524,N_21478,N_21925);
or U22525 (N_22525,N_21951,N_21455);
nand U22526 (N_22526,N_21881,N_21753);
or U22527 (N_22527,N_21626,N_21261);
xnor U22528 (N_22528,N_21248,N_21118);
xnor U22529 (N_22529,N_21052,N_21462);
nor U22530 (N_22530,N_21200,N_21219);
xor U22531 (N_22531,N_21323,N_21529);
and U22532 (N_22532,N_21243,N_21118);
nand U22533 (N_22533,N_21701,N_21264);
and U22534 (N_22534,N_21466,N_21250);
nand U22535 (N_22535,N_21080,N_21628);
nand U22536 (N_22536,N_21199,N_21334);
and U22537 (N_22537,N_21930,N_21898);
nand U22538 (N_22538,N_21476,N_21468);
and U22539 (N_22539,N_21834,N_21506);
xnor U22540 (N_22540,N_21152,N_21559);
and U22541 (N_22541,N_21394,N_21410);
nand U22542 (N_22542,N_21401,N_21600);
and U22543 (N_22543,N_21116,N_21053);
nand U22544 (N_22544,N_21829,N_21048);
or U22545 (N_22545,N_21432,N_21412);
and U22546 (N_22546,N_21603,N_21421);
nor U22547 (N_22547,N_21847,N_21160);
nor U22548 (N_22548,N_21212,N_21642);
nor U22549 (N_22549,N_21865,N_21558);
nor U22550 (N_22550,N_21894,N_21705);
nand U22551 (N_22551,N_21966,N_21594);
nand U22552 (N_22552,N_21686,N_21920);
or U22553 (N_22553,N_21489,N_21824);
xor U22554 (N_22554,N_21555,N_21371);
and U22555 (N_22555,N_21547,N_21468);
nor U22556 (N_22556,N_21804,N_21598);
xor U22557 (N_22557,N_21176,N_21333);
or U22558 (N_22558,N_21582,N_21553);
or U22559 (N_22559,N_21620,N_21132);
nand U22560 (N_22560,N_21286,N_21823);
nor U22561 (N_22561,N_21013,N_21315);
nor U22562 (N_22562,N_21757,N_21173);
nor U22563 (N_22563,N_21197,N_21905);
and U22564 (N_22564,N_21687,N_21794);
nand U22565 (N_22565,N_21752,N_21003);
nand U22566 (N_22566,N_21938,N_21799);
and U22567 (N_22567,N_21559,N_21127);
and U22568 (N_22568,N_21330,N_21906);
and U22569 (N_22569,N_21570,N_21359);
nor U22570 (N_22570,N_21647,N_21238);
nand U22571 (N_22571,N_21846,N_21742);
nor U22572 (N_22572,N_21091,N_21867);
or U22573 (N_22573,N_21697,N_21000);
xnor U22574 (N_22574,N_21519,N_21891);
xor U22575 (N_22575,N_21223,N_21035);
nand U22576 (N_22576,N_21756,N_21994);
or U22577 (N_22577,N_21342,N_21309);
or U22578 (N_22578,N_21307,N_21128);
xnor U22579 (N_22579,N_21183,N_21896);
nor U22580 (N_22580,N_21545,N_21910);
nand U22581 (N_22581,N_21594,N_21762);
and U22582 (N_22582,N_21890,N_21122);
nand U22583 (N_22583,N_21191,N_21289);
nand U22584 (N_22584,N_21491,N_21885);
xnor U22585 (N_22585,N_21082,N_21910);
xor U22586 (N_22586,N_21280,N_21174);
nand U22587 (N_22587,N_21931,N_21287);
or U22588 (N_22588,N_21734,N_21493);
and U22589 (N_22589,N_21124,N_21912);
nor U22590 (N_22590,N_21514,N_21886);
or U22591 (N_22591,N_21258,N_21755);
nor U22592 (N_22592,N_21718,N_21124);
or U22593 (N_22593,N_21924,N_21772);
or U22594 (N_22594,N_21067,N_21460);
and U22595 (N_22595,N_21624,N_21477);
xnor U22596 (N_22596,N_21974,N_21316);
xor U22597 (N_22597,N_21566,N_21011);
nor U22598 (N_22598,N_21643,N_21769);
xor U22599 (N_22599,N_21579,N_21860);
or U22600 (N_22600,N_21764,N_21874);
nor U22601 (N_22601,N_21882,N_21088);
nand U22602 (N_22602,N_21581,N_21992);
or U22603 (N_22603,N_21642,N_21856);
nand U22604 (N_22604,N_21096,N_21358);
or U22605 (N_22605,N_21537,N_21215);
or U22606 (N_22606,N_21808,N_21183);
or U22607 (N_22607,N_21872,N_21077);
nor U22608 (N_22608,N_21220,N_21793);
or U22609 (N_22609,N_21499,N_21797);
or U22610 (N_22610,N_21756,N_21676);
or U22611 (N_22611,N_21936,N_21184);
nor U22612 (N_22612,N_21587,N_21279);
xnor U22613 (N_22613,N_21182,N_21591);
or U22614 (N_22614,N_21323,N_21676);
nor U22615 (N_22615,N_21839,N_21168);
xnor U22616 (N_22616,N_21523,N_21930);
xor U22617 (N_22617,N_21989,N_21935);
nor U22618 (N_22618,N_21028,N_21062);
xnor U22619 (N_22619,N_21864,N_21356);
xor U22620 (N_22620,N_21445,N_21662);
nand U22621 (N_22621,N_21008,N_21487);
or U22622 (N_22622,N_21380,N_21681);
nor U22623 (N_22623,N_21206,N_21055);
xor U22624 (N_22624,N_21731,N_21418);
nor U22625 (N_22625,N_21721,N_21770);
xor U22626 (N_22626,N_21173,N_21942);
or U22627 (N_22627,N_21660,N_21823);
nand U22628 (N_22628,N_21486,N_21676);
xnor U22629 (N_22629,N_21088,N_21080);
nor U22630 (N_22630,N_21931,N_21923);
nand U22631 (N_22631,N_21265,N_21149);
nor U22632 (N_22632,N_21008,N_21863);
or U22633 (N_22633,N_21858,N_21509);
xor U22634 (N_22634,N_21400,N_21235);
nor U22635 (N_22635,N_21773,N_21027);
and U22636 (N_22636,N_21105,N_21281);
nand U22637 (N_22637,N_21928,N_21219);
or U22638 (N_22638,N_21907,N_21398);
nand U22639 (N_22639,N_21690,N_21566);
xor U22640 (N_22640,N_21753,N_21301);
xor U22641 (N_22641,N_21779,N_21248);
nand U22642 (N_22642,N_21573,N_21675);
nor U22643 (N_22643,N_21194,N_21208);
or U22644 (N_22644,N_21137,N_21412);
and U22645 (N_22645,N_21293,N_21960);
and U22646 (N_22646,N_21289,N_21140);
nor U22647 (N_22647,N_21134,N_21748);
xnor U22648 (N_22648,N_21627,N_21640);
and U22649 (N_22649,N_21035,N_21329);
or U22650 (N_22650,N_21037,N_21201);
nor U22651 (N_22651,N_21613,N_21391);
nand U22652 (N_22652,N_21920,N_21037);
xor U22653 (N_22653,N_21962,N_21052);
xnor U22654 (N_22654,N_21286,N_21307);
xnor U22655 (N_22655,N_21986,N_21830);
nor U22656 (N_22656,N_21274,N_21503);
xor U22657 (N_22657,N_21040,N_21967);
nand U22658 (N_22658,N_21686,N_21139);
nand U22659 (N_22659,N_21016,N_21326);
and U22660 (N_22660,N_21736,N_21680);
and U22661 (N_22661,N_21783,N_21899);
nand U22662 (N_22662,N_21267,N_21281);
nor U22663 (N_22663,N_21731,N_21379);
and U22664 (N_22664,N_21568,N_21944);
xnor U22665 (N_22665,N_21009,N_21132);
or U22666 (N_22666,N_21639,N_21801);
nand U22667 (N_22667,N_21439,N_21896);
and U22668 (N_22668,N_21953,N_21087);
xor U22669 (N_22669,N_21739,N_21543);
nor U22670 (N_22670,N_21941,N_21924);
and U22671 (N_22671,N_21740,N_21257);
and U22672 (N_22672,N_21125,N_21036);
or U22673 (N_22673,N_21160,N_21713);
nor U22674 (N_22674,N_21470,N_21009);
or U22675 (N_22675,N_21283,N_21857);
or U22676 (N_22676,N_21651,N_21673);
nor U22677 (N_22677,N_21885,N_21935);
nor U22678 (N_22678,N_21303,N_21908);
and U22679 (N_22679,N_21583,N_21601);
xor U22680 (N_22680,N_21608,N_21926);
nand U22681 (N_22681,N_21029,N_21524);
and U22682 (N_22682,N_21714,N_21207);
xor U22683 (N_22683,N_21089,N_21335);
nand U22684 (N_22684,N_21756,N_21782);
nor U22685 (N_22685,N_21058,N_21036);
xor U22686 (N_22686,N_21550,N_21237);
or U22687 (N_22687,N_21592,N_21407);
and U22688 (N_22688,N_21550,N_21667);
nand U22689 (N_22689,N_21352,N_21699);
nor U22690 (N_22690,N_21735,N_21815);
nor U22691 (N_22691,N_21998,N_21701);
nor U22692 (N_22692,N_21402,N_21876);
or U22693 (N_22693,N_21405,N_21823);
xor U22694 (N_22694,N_21911,N_21024);
nor U22695 (N_22695,N_21886,N_21636);
nand U22696 (N_22696,N_21797,N_21735);
nand U22697 (N_22697,N_21962,N_21690);
xor U22698 (N_22698,N_21383,N_21988);
nand U22699 (N_22699,N_21913,N_21974);
xnor U22700 (N_22700,N_21194,N_21461);
or U22701 (N_22701,N_21716,N_21360);
and U22702 (N_22702,N_21121,N_21170);
nand U22703 (N_22703,N_21329,N_21954);
nor U22704 (N_22704,N_21777,N_21725);
or U22705 (N_22705,N_21760,N_21756);
and U22706 (N_22706,N_21645,N_21490);
xnor U22707 (N_22707,N_21670,N_21292);
nor U22708 (N_22708,N_21734,N_21875);
or U22709 (N_22709,N_21126,N_21516);
and U22710 (N_22710,N_21473,N_21655);
and U22711 (N_22711,N_21855,N_21458);
nand U22712 (N_22712,N_21073,N_21701);
nor U22713 (N_22713,N_21141,N_21283);
xnor U22714 (N_22714,N_21716,N_21717);
nor U22715 (N_22715,N_21224,N_21274);
xnor U22716 (N_22716,N_21041,N_21220);
and U22717 (N_22717,N_21599,N_21432);
and U22718 (N_22718,N_21280,N_21981);
and U22719 (N_22719,N_21236,N_21212);
xor U22720 (N_22720,N_21702,N_21365);
nor U22721 (N_22721,N_21395,N_21563);
nand U22722 (N_22722,N_21444,N_21581);
or U22723 (N_22723,N_21130,N_21278);
and U22724 (N_22724,N_21159,N_21126);
or U22725 (N_22725,N_21720,N_21735);
nor U22726 (N_22726,N_21619,N_21384);
nand U22727 (N_22727,N_21948,N_21140);
nor U22728 (N_22728,N_21947,N_21617);
or U22729 (N_22729,N_21962,N_21923);
and U22730 (N_22730,N_21826,N_21027);
nand U22731 (N_22731,N_21890,N_21565);
or U22732 (N_22732,N_21386,N_21085);
nor U22733 (N_22733,N_21465,N_21823);
xor U22734 (N_22734,N_21222,N_21419);
and U22735 (N_22735,N_21158,N_21707);
xnor U22736 (N_22736,N_21252,N_21375);
or U22737 (N_22737,N_21229,N_21745);
or U22738 (N_22738,N_21533,N_21492);
or U22739 (N_22739,N_21511,N_21395);
xnor U22740 (N_22740,N_21541,N_21134);
or U22741 (N_22741,N_21889,N_21628);
nor U22742 (N_22742,N_21806,N_21808);
xnor U22743 (N_22743,N_21669,N_21092);
xor U22744 (N_22744,N_21469,N_21042);
xor U22745 (N_22745,N_21277,N_21065);
and U22746 (N_22746,N_21610,N_21524);
nor U22747 (N_22747,N_21495,N_21819);
or U22748 (N_22748,N_21615,N_21946);
nor U22749 (N_22749,N_21870,N_21506);
nand U22750 (N_22750,N_21062,N_21815);
and U22751 (N_22751,N_21151,N_21399);
nand U22752 (N_22752,N_21247,N_21090);
xnor U22753 (N_22753,N_21946,N_21694);
or U22754 (N_22754,N_21485,N_21916);
xor U22755 (N_22755,N_21177,N_21925);
xor U22756 (N_22756,N_21192,N_21666);
xor U22757 (N_22757,N_21442,N_21065);
and U22758 (N_22758,N_21987,N_21903);
and U22759 (N_22759,N_21193,N_21537);
or U22760 (N_22760,N_21328,N_21556);
and U22761 (N_22761,N_21508,N_21122);
nand U22762 (N_22762,N_21152,N_21937);
or U22763 (N_22763,N_21373,N_21024);
nand U22764 (N_22764,N_21513,N_21124);
nand U22765 (N_22765,N_21635,N_21431);
or U22766 (N_22766,N_21430,N_21479);
xnor U22767 (N_22767,N_21366,N_21224);
or U22768 (N_22768,N_21982,N_21366);
or U22769 (N_22769,N_21532,N_21789);
xnor U22770 (N_22770,N_21531,N_21120);
and U22771 (N_22771,N_21237,N_21093);
xnor U22772 (N_22772,N_21136,N_21641);
and U22773 (N_22773,N_21265,N_21411);
nor U22774 (N_22774,N_21910,N_21172);
nand U22775 (N_22775,N_21700,N_21971);
and U22776 (N_22776,N_21630,N_21096);
nand U22777 (N_22777,N_21733,N_21999);
xor U22778 (N_22778,N_21407,N_21627);
and U22779 (N_22779,N_21858,N_21047);
or U22780 (N_22780,N_21096,N_21470);
and U22781 (N_22781,N_21294,N_21449);
and U22782 (N_22782,N_21829,N_21374);
xnor U22783 (N_22783,N_21322,N_21427);
or U22784 (N_22784,N_21683,N_21254);
and U22785 (N_22785,N_21975,N_21141);
nor U22786 (N_22786,N_21302,N_21651);
xnor U22787 (N_22787,N_21528,N_21204);
nor U22788 (N_22788,N_21255,N_21467);
xor U22789 (N_22789,N_21690,N_21903);
and U22790 (N_22790,N_21155,N_21351);
nor U22791 (N_22791,N_21289,N_21188);
nor U22792 (N_22792,N_21050,N_21278);
nor U22793 (N_22793,N_21366,N_21146);
or U22794 (N_22794,N_21657,N_21907);
and U22795 (N_22795,N_21016,N_21274);
xnor U22796 (N_22796,N_21219,N_21435);
nand U22797 (N_22797,N_21226,N_21046);
nor U22798 (N_22798,N_21496,N_21482);
nor U22799 (N_22799,N_21730,N_21049);
nor U22800 (N_22800,N_21433,N_21224);
xnor U22801 (N_22801,N_21089,N_21564);
or U22802 (N_22802,N_21156,N_21197);
nor U22803 (N_22803,N_21208,N_21280);
and U22804 (N_22804,N_21386,N_21243);
nand U22805 (N_22805,N_21406,N_21613);
xnor U22806 (N_22806,N_21590,N_21088);
xnor U22807 (N_22807,N_21886,N_21726);
nor U22808 (N_22808,N_21097,N_21934);
or U22809 (N_22809,N_21923,N_21824);
and U22810 (N_22810,N_21553,N_21491);
and U22811 (N_22811,N_21643,N_21103);
nor U22812 (N_22812,N_21668,N_21244);
nand U22813 (N_22813,N_21391,N_21683);
nand U22814 (N_22814,N_21752,N_21470);
nor U22815 (N_22815,N_21752,N_21624);
or U22816 (N_22816,N_21505,N_21913);
and U22817 (N_22817,N_21716,N_21478);
and U22818 (N_22818,N_21893,N_21739);
and U22819 (N_22819,N_21359,N_21208);
and U22820 (N_22820,N_21892,N_21070);
nor U22821 (N_22821,N_21609,N_21945);
nor U22822 (N_22822,N_21442,N_21631);
xor U22823 (N_22823,N_21613,N_21096);
and U22824 (N_22824,N_21808,N_21360);
and U22825 (N_22825,N_21265,N_21317);
or U22826 (N_22826,N_21058,N_21865);
or U22827 (N_22827,N_21044,N_21790);
nand U22828 (N_22828,N_21612,N_21761);
nand U22829 (N_22829,N_21780,N_21072);
and U22830 (N_22830,N_21381,N_21355);
nor U22831 (N_22831,N_21953,N_21175);
or U22832 (N_22832,N_21742,N_21638);
and U22833 (N_22833,N_21291,N_21995);
nand U22834 (N_22834,N_21953,N_21427);
or U22835 (N_22835,N_21478,N_21350);
xnor U22836 (N_22836,N_21703,N_21450);
nand U22837 (N_22837,N_21363,N_21230);
nand U22838 (N_22838,N_21067,N_21282);
nor U22839 (N_22839,N_21191,N_21081);
nor U22840 (N_22840,N_21700,N_21958);
and U22841 (N_22841,N_21777,N_21234);
or U22842 (N_22842,N_21522,N_21237);
or U22843 (N_22843,N_21990,N_21077);
or U22844 (N_22844,N_21844,N_21417);
nor U22845 (N_22845,N_21223,N_21903);
nor U22846 (N_22846,N_21592,N_21737);
and U22847 (N_22847,N_21159,N_21759);
or U22848 (N_22848,N_21037,N_21176);
nor U22849 (N_22849,N_21670,N_21333);
and U22850 (N_22850,N_21928,N_21757);
nor U22851 (N_22851,N_21532,N_21546);
nand U22852 (N_22852,N_21740,N_21734);
nor U22853 (N_22853,N_21381,N_21965);
nand U22854 (N_22854,N_21937,N_21477);
and U22855 (N_22855,N_21342,N_21193);
nor U22856 (N_22856,N_21084,N_21187);
and U22857 (N_22857,N_21585,N_21392);
nand U22858 (N_22858,N_21678,N_21014);
xor U22859 (N_22859,N_21743,N_21678);
or U22860 (N_22860,N_21097,N_21807);
and U22861 (N_22861,N_21777,N_21983);
nand U22862 (N_22862,N_21499,N_21611);
nor U22863 (N_22863,N_21351,N_21478);
nand U22864 (N_22864,N_21144,N_21999);
xnor U22865 (N_22865,N_21384,N_21732);
and U22866 (N_22866,N_21600,N_21821);
and U22867 (N_22867,N_21835,N_21557);
xor U22868 (N_22868,N_21578,N_21310);
nand U22869 (N_22869,N_21702,N_21130);
xor U22870 (N_22870,N_21755,N_21130);
nor U22871 (N_22871,N_21554,N_21681);
xor U22872 (N_22872,N_21087,N_21091);
or U22873 (N_22873,N_21715,N_21840);
and U22874 (N_22874,N_21140,N_21045);
nand U22875 (N_22875,N_21288,N_21237);
or U22876 (N_22876,N_21047,N_21415);
nor U22877 (N_22877,N_21569,N_21616);
nand U22878 (N_22878,N_21003,N_21375);
nand U22879 (N_22879,N_21810,N_21100);
and U22880 (N_22880,N_21299,N_21024);
nand U22881 (N_22881,N_21317,N_21210);
or U22882 (N_22882,N_21696,N_21722);
or U22883 (N_22883,N_21525,N_21344);
nor U22884 (N_22884,N_21866,N_21293);
or U22885 (N_22885,N_21370,N_21026);
or U22886 (N_22886,N_21237,N_21352);
and U22887 (N_22887,N_21419,N_21425);
nand U22888 (N_22888,N_21388,N_21320);
nand U22889 (N_22889,N_21642,N_21521);
and U22890 (N_22890,N_21010,N_21115);
nand U22891 (N_22891,N_21112,N_21180);
and U22892 (N_22892,N_21267,N_21139);
nor U22893 (N_22893,N_21120,N_21359);
nand U22894 (N_22894,N_21799,N_21529);
nand U22895 (N_22895,N_21761,N_21530);
nand U22896 (N_22896,N_21279,N_21658);
nand U22897 (N_22897,N_21680,N_21017);
and U22898 (N_22898,N_21661,N_21284);
or U22899 (N_22899,N_21131,N_21013);
nor U22900 (N_22900,N_21763,N_21332);
nand U22901 (N_22901,N_21767,N_21410);
nand U22902 (N_22902,N_21242,N_21722);
xnor U22903 (N_22903,N_21963,N_21391);
nand U22904 (N_22904,N_21803,N_21096);
xor U22905 (N_22905,N_21157,N_21618);
or U22906 (N_22906,N_21167,N_21353);
nor U22907 (N_22907,N_21747,N_21414);
nor U22908 (N_22908,N_21639,N_21997);
nor U22909 (N_22909,N_21937,N_21016);
and U22910 (N_22910,N_21862,N_21393);
xor U22911 (N_22911,N_21121,N_21979);
nor U22912 (N_22912,N_21301,N_21531);
nor U22913 (N_22913,N_21661,N_21303);
or U22914 (N_22914,N_21118,N_21486);
nand U22915 (N_22915,N_21597,N_21315);
or U22916 (N_22916,N_21924,N_21521);
xnor U22917 (N_22917,N_21184,N_21842);
and U22918 (N_22918,N_21172,N_21083);
or U22919 (N_22919,N_21203,N_21124);
xnor U22920 (N_22920,N_21502,N_21578);
nor U22921 (N_22921,N_21319,N_21791);
and U22922 (N_22922,N_21273,N_21564);
nand U22923 (N_22923,N_21147,N_21455);
xor U22924 (N_22924,N_21587,N_21868);
xor U22925 (N_22925,N_21902,N_21487);
or U22926 (N_22926,N_21821,N_21073);
nor U22927 (N_22927,N_21729,N_21505);
nor U22928 (N_22928,N_21938,N_21722);
nand U22929 (N_22929,N_21658,N_21477);
nor U22930 (N_22930,N_21254,N_21703);
and U22931 (N_22931,N_21650,N_21068);
or U22932 (N_22932,N_21474,N_21238);
nand U22933 (N_22933,N_21804,N_21018);
and U22934 (N_22934,N_21123,N_21843);
or U22935 (N_22935,N_21229,N_21107);
xnor U22936 (N_22936,N_21430,N_21471);
nor U22937 (N_22937,N_21965,N_21113);
nand U22938 (N_22938,N_21519,N_21481);
nand U22939 (N_22939,N_21497,N_21789);
nand U22940 (N_22940,N_21416,N_21721);
or U22941 (N_22941,N_21879,N_21156);
nor U22942 (N_22942,N_21147,N_21846);
and U22943 (N_22943,N_21674,N_21685);
or U22944 (N_22944,N_21295,N_21359);
or U22945 (N_22945,N_21453,N_21424);
nor U22946 (N_22946,N_21856,N_21029);
and U22947 (N_22947,N_21020,N_21337);
nor U22948 (N_22948,N_21511,N_21425);
nor U22949 (N_22949,N_21666,N_21803);
nand U22950 (N_22950,N_21890,N_21290);
and U22951 (N_22951,N_21104,N_21167);
xnor U22952 (N_22952,N_21433,N_21324);
nor U22953 (N_22953,N_21965,N_21387);
xor U22954 (N_22954,N_21565,N_21909);
nor U22955 (N_22955,N_21782,N_21948);
or U22956 (N_22956,N_21029,N_21847);
or U22957 (N_22957,N_21069,N_21559);
or U22958 (N_22958,N_21819,N_21115);
xor U22959 (N_22959,N_21279,N_21905);
and U22960 (N_22960,N_21088,N_21730);
xnor U22961 (N_22961,N_21440,N_21645);
and U22962 (N_22962,N_21883,N_21342);
nor U22963 (N_22963,N_21561,N_21374);
nor U22964 (N_22964,N_21505,N_21562);
nand U22965 (N_22965,N_21074,N_21998);
nor U22966 (N_22966,N_21586,N_21612);
and U22967 (N_22967,N_21298,N_21809);
nand U22968 (N_22968,N_21396,N_21290);
nand U22969 (N_22969,N_21284,N_21922);
or U22970 (N_22970,N_21258,N_21420);
nor U22971 (N_22971,N_21672,N_21850);
xor U22972 (N_22972,N_21009,N_21700);
or U22973 (N_22973,N_21520,N_21873);
or U22974 (N_22974,N_21236,N_21755);
nand U22975 (N_22975,N_21804,N_21641);
and U22976 (N_22976,N_21282,N_21631);
xnor U22977 (N_22977,N_21064,N_21294);
nand U22978 (N_22978,N_21586,N_21542);
or U22979 (N_22979,N_21907,N_21320);
xnor U22980 (N_22980,N_21782,N_21408);
and U22981 (N_22981,N_21872,N_21341);
nor U22982 (N_22982,N_21641,N_21251);
xor U22983 (N_22983,N_21776,N_21658);
nor U22984 (N_22984,N_21730,N_21605);
nand U22985 (N_22985,N_21457,N_21095);
nand U22986 (N_22986,N_21899,N_21429);
and U22987 (N_22987,N_21134,N_21056);
nor U22988 (N_22988,N_21358,N_21948);
and U22989 (N_22989,N_21835,N_21345);
or U22990 (N_22990,N_21262,N_21696);
nand U22991 (N_22991,N_21166,N_21482);
or U22992 (N_22992,N_21901,N_21827);
or U22993 (N_22993,N_21219,N_21850);
nor U22994 (N_22994,N_21232,N_21181);
and U22995 (N_22995,N_21738,N_21640);
or U22996 (N_22996,N_21488,N_21523);
nand U22997 (N_22997,N_21284,N_21246);
or U22998 (N_22998,N_21280,N_21752);
or U22999 (N_22999,N_21887,N_21714);
or U23000 (N_23000,N_22070,N_22775);
nor U23001 (N_23001,N_22719,N_22909);
xor U23002 (N_23002,N_22529,N_22659);
nor U23003 (N_23003,N_22936,N_22415);
xor U23004 (N_23004,N_22481,N_22399);
or U23005 (N_23005,N_22258,N_22249);
nand U23006 (N_23006,N_22573,N_22537);
or U23007 (N_23007,N_22003,N_22710);
nor U23008 (N_23008,N_22228,N_22127);
nand U23009 (N_23009,N_22293,N_22066);
or U23010 (N_23010,N_22502,N_22947);
xnor U23011 (N_23011,N_22556,N_22044);
nand U23012 (N_23012,N_22711,N_22946);
and U23013 (N_23013,N_22793,N_22312);
or U23014 (N_23014,N_22584,N_22962);
nor U23015 (N_23015,N_22074,N_22208);
xor U23016 (N_23016,N_22037,N_22476);
nand U23017 (N_23017,N_22891,N_22534);
nand U23018 (N_23018,N_22542,N_22696);
and U23019 (N_23019,N_22553,N_22252);
or U23020 (N_23020,N_22482,N_22180);
and U23021 (N_23021,N_22002,N_22664);
xor U23022 (N_23022,N_22692,N_22177);
or U23023 (N_23023,N_22028,N_22164);
nand U23024 (N_23024,N_22192,N_22738);
and U23025 (N_23025,N_22301,N_22328);
xor U23026 (N_23026,N_22398,N_22352);
nor U23027 (N_23027,N_22675,N_22996);
or U23028 (N_23028,N_22004,N_22678);
or U23029 (N_23029,N_22205,N_22585);
or U23030 (N_23030,N_22467,N_22320);
and U23031 (N_23031,N_22688,N_22437);
or U23032 (N_23032,N_22876,N_22650);
and U23033 (N_23033,N_22651,N_22547);
nand U23034 (N_23034,N_22634,N_22552);
xnor U23035 (N_23035,N_22461,N_22948);
and U23036 (N_23036,N_22564,N_22364);
and U23037 (N_23037,N_22965,N_22158);
nand U23038 (N_23038,N_22985,N_22250);
and U23039 (N_23039,N_22818,N_22103);
or U23040 (N_23040,N_22338,N_22131);
or U23041 (N_23041,N_22102,N_22238);
nand U23042 (N_23042,N_22287,N_22087);
nand U23043 (N_23043,N_22539,N_22323);
xnor U23044 (N_23044,N_22754,N_22827);
and U23045 (N_23045,N_22939,N_22815);
or U23046 (N_23046,N_22434,N_22728);
and U23047 (N_23047,N_22196,N_22438);
or U23048 (N_23048,N_22605,N_22060);
nand U23049 (N_23049,N_22591,N_22737);
or U23050 (N_23050,N_22864,N_22852);
nand U23051 (N_23051,N_22630,N_22367);
nand U23052 (N_23052,N_22395,N_22752);
and U23053 (N_23053,N_22804,N_22247);
and U23054 (N_23054,N_22337,N_22075);
nor U23055 (N_23055,N_22823,N_22007);
nand U23056 (N_23056,N_22511,N_22483);
and U23057 (N_23057,N_22590,N_22078);
nor U23058 (N_23058,N_22642,N_22363);
nor U23059 (N_23059,N_22832,N_22197);
or U23060 (N_23060,N_22095,N_22978);
nand U23061 (N_23061,N_22824,N_22845);
xor U23062 (N_23062,N_22181,N_22175);
xor U23063 (N_23063,N_22491,N_22152);
nor U23064 (N_23064,N_22648,N_22612);
or U23065 (N_23065,N_22810,N_22418);
or U23066 (N_23066,N_22819,N_22530);
nor U23067 (N_23067,N_22681,N_22666);
nand U23068 (N_23068,N_22631,N_22785);
xor U23069 (N_23069,N_22967,N_22740);
nand U23070 (N_23070,N_22093,N_22052);
xor U23071 (N_23071,N_22492,N_22500);
xor U23072 (N_23072,N_22234,N_22883);
nor U23073 (N_23073,N_22774,N_22061);
nor U23074 (N_23074,N_22694,N_22910);
xnor U23075 (N_23075,N_22885,N_22527);
xnor U23076 (N_23076,N_22034,N_22430);
nand U23077 (N_23077,N_22772,N_22836);
xor U23078 (N_23078,N_22463,N_22148);
and U23079 (N_23079,N_22062,N_22551);
xnor U23080 (N_23080,N_22381,N_22041);
and U23081 (N_23081,N_22233,N_22941);
nor U23082 (N_23082,N_22391,N_22146);
nand U23083 (N_23083,N_22156,N_22118);
nor U23084 (N_23084,N_22643,N_22106);
xnor U23085 (N_23085,N_22445,N_22783);
or U23086 (N_23086,N_22270,N_22409);
and U23087 (N_23087,N_22667,N_22732);
and U23088 (N_23088,N_22767,N_22276);
xor U23089 (N_23089,N_22439,N_22566);
nand U23090 (N_23090,N_22045,N_22968);
nor U23091 (N_23091,N_22903,N_22105);
nor U23092 (N_23092,N_22092,N_22786);
and U23093 (N_23093,N_22682,N_22942);
nor U23094 (N_23094,N_22742,N_22302);
or U23095 (N_23095,N_22571,N_22730);
or U23096 (N_23096,N_22873,N_22023);
xnor U23097 (N_23097,N_22954,N_22030);
nor U23098 (N_23098,N_22884,N_22216);
xnor U23099 (N_23099,N_22218,N_22474);
and U23100 (N_23100,N_22330,N_22006);
nor U23101 (N_23101,N_22406,N_22424);
nor U23102 (N_23102,N_22859,N_22653);
or U23103 (N_23103,N_22230,N_22067);
nor U23104 (N_23104,N_22227,N_22874);
or U23105 (N_23105,N_22988,N_22402);
or U23106 (N_23106,N_22458,N_22318);
or U23107 (N_23107,N_22372,N_22248);
and U23108 (N_23108,N_22964,N_22531);
or U23109 (N_23109,N_22384,N_22160);
nand U23110 (N_23110,N_22897,N_22495);
xor U23111 (N_23111,N_22613,N_22351);
nand U23112 (N_23112,N_22206,N_22173);
and U23113 (N_23113,N_22262,N_22599);
nor U23114 (N_23114,N_22683,N_22453);
and U23115 (N_23115,N_22307,N_22188);
nor U23116 (N_23116,N_22280,N_22898);
or U23117 (N_23117,N_22207,N_22673);
xnor U23118 (N_23118,N_22532,N_22866);
xor U23119 (N_23119,N_22543,N_22271);
xor U23120 (N_23120,N_22149,N_22649);
nor U23121 (N_23121,N_22796,N_22782);
or U23122 (N_23122,N_22285,N_22360);
nand U23123 (N_23123,N_22282,N_22871);
xnor U23124 (N_23124,N_22494,N_22805);
nand U23125 (N_23125,N_22848,N_22171);
or U23126 (N_23126,N_22083,N_22563);
nand U23127 (N_23127,N_22935,N_22068);
xnor U23128 (N_23128,N_22038,N_22408);
xnor U23129 (N_23129,N_22615,N_22593);
and U23130 (N_23130,N_22830,N_22586);
nand U23131 (N_23131,N_22795,N_22436);
and U23132 (N_23132,N_22015,N_22776);
nor U23133 (N_23133,N_22700,N_22879);
nand U23134 (N_23134,N_22153,N_22569);
xnor U23135 (N_23135,N_22608,N_22908);
nand U23136 (N_23136,N_22905,N_22868);
nand U23137 (N_23137,N_22329,N_22315);
and U23138 (N_23138,N_22349,N_22524);
nand U23139 (N_23139,N_22843,N_22484);
and U23140 (N_23140,N_22291,N_22221);
and U23141 (N_23141,N_22707,N_22919);
xor U23142 (N_23142,N_22505,N_22178);
xor U23143 (N_23143,N_22575,N_22000);
or U23144 (N_23144,N_22844,N_22091);
and U23145 (N_23145,N_22231,N_22325);
nand U23146 (N_23146,N_22620,N_22841);
nor U23147 (N_23147,N_22369,N_22099);
xor U23148 (N_23148,N_22224,N_22410);
xnor U23149 (N_23149,N_22922,N_22598);
or U23150 (N_23150,N_22992,N_22993);
xnor U23151 (N_23151,N_22220,N_22375);
and U23152 (N_23152,N_22750,N_22400);
and U23153 (N_23153,N_22603,N_22284);
nor U23154 (N_23154,N_22472,N_22488);
nand U23155 (N_23155,N_22466,N_22264);
nand U23156 (N_23156,N_22656,N_22035);
and U23157 (N_23157,N_22899,N_22619);
nand U23158 (N_23158,N_22849,N_22385);
and U23159 (N_23159,N_22346,N_22961);
nor U23160 (N_23160,N_22272,N_22842);
xnor U23161 (N_23161,N_22089,N_22503);
nand U23162 (N_23162,N_22135,N_22036);
nor U23163 (N_23163,N_22456,N_22705);
nor U23164 (N_23164,N_22911,N_22746);
nand U23165 (N_23165,N_22404,N_22184);
nor U23166 (N_23166,N_22341,N_22888);
nand U23167 (N_23167,N_22016,N_22383);
or U23168 (N_23168,N_22469,N_22671);
xnor U23169 (N_23169,N_22441,N_22699);
or U23170 (N_23170,N_22257,N_22266);
and U23171 (N_23171,N_22283,N_22345);
nor U23172 (N_23172,N_22663,N_22155);
or U23173 (N_23173,N_22957,N_22595);
nand U23174 (N_23174,N_22588,N_22979);
or U23175 (N_23175,N_22535,N_22661);
nand U23176 (N_23176,N_22519,N_22626);
or U23177 (N_23177,N_22863,N_22689);
or U23178 (N_23178,N_22969,N_22596);
or U23179 (N_23179,N_22826,N_22421);
nand U23180 (N_23180,N_22557,N_22455);
or U23181 (N_23181,N_22142,N_22814);
or U23182 (N_23182,N_22803,N_22745);
and U23183 (N_23183,N_22520,N_22213);
nand U23184 (N_23184,N_22870,N_22869);
nand U23185 (N_23185,N_22239,N_22450);
nand U23186 (N_23186,N_22963,N_22063);
xor U23187 (N_23187,N_22020,N_22770);
or U23188 (N_23188,N_22447,N_22528);
and U23189 (N_23189,N_22057,N_22760);
or U23190 (N_23190,N_22674,N_22310);
xnor U23191 (N_23191,N_22636,N_22609);
or U23192 (N_23192,N_22151,N_22974);
nor U23193 (N_23193,N_22925,N_22555);
xor U23194 (N_23194,N_22422,N_22998);
or U23195 (N_23195,N_22693,N_22324);
nor U23196 (N_23196,N_22617,N_22332);
and U23197 (N_23197,N_22316,N_22607);
nand U23198 (N_23198,N_22644,N_22281);
xnor U23199 (N_23199,N_22702,N_22076);
xnor U23200 (N_23200,N_22995,N_22202);
xor U23201 (N_23201,N_22256,N_22669);
or U23202 (N_23202,N_22145,N_22778);
xnor U23203 (N_23203,N_22813,N_22183);
or U23204 (N_23204,N_22347,N_22241);
and U23205 (N_23205,N_22255,N_22670);
xnor U23206 (N_23206,N_22652,N_22983);
nand U23207 (N_23207,N_22713,N_22378);
nor U23208 (N_23208,N_22986,N_22881);
and U23209 (N_23209,N_22443,N_22377);
nand U23210 (N_23210,N_22460,N_22182);
xor U23211 (N_23211,N_22496,N_22420);
xor U23212 (N_23212,N_22565,N_22236);
nand U23213 (N_23213,N_22340,N_22017);
nor U23214 (N_23214,N_22254,N_22428);
nor U23215 (N_23215,N_22214,N_22751);
or U23216 (N_23216,N_22792,N_22574);
nand U23217 (N_23217,N_22762,N_22123);
nand U23218 (N_23218,N_22305,N_22896);
xor U23219 (N_23219,N_22677,N_22654);
nand U23220 (N_23220,N_22921,N_22319);
xor U23221 (N_23221,N_22514,N_22727);
nand U23222 (N_23222,N_22960,N_22261);
or U23223 (N_23223,N_22080,N_22309);
nor U23224 (N_23224,N_22433,N_22314);
and U23225 (N_23225,N_22163,N_22703);
and U23226 (N_23226,N_22971,N_22286);
nor U23227 (N_23227,N_22982,N_22121);
nand U23228 (N_23228,N_22718,N_22274);
xnor U23229 (N_23229,N_22950,N_22958);
or U23230 (N_23230,N_22684,N_22789);
and U23231 (N_23231,N_22244,N_22486);
or U23232 (N_23232,N_22934,N_22162);
and U23233 (N_23233,N_22594,N_22821);
and U23234 (N_23234,N_22457,N_22435);
nor U23235 (N_23235,N_22432,N_22051);
xor U23236 (N_23236,N_22984,N_22382);
or U23237 (N_23237,N_22582,N_22989);
xor U23238 (N_23238,N_22801,N_22886);
and U23239 (N_23239,N_22840,N_22096);
and U23240 (N_23240,N_22114,N_22655);
or U23241 (N_23241,N_22739,N_22024);
nor U23242 (N_23242,N_22943,N_22267);
or U23243 (N_23243,N_22311,N_22721);
and U23244 (N_23244,N_22056,N_22251);
xnor U23245 (N_23245,N_22465,N_22190);
nand U23246 (N_23246,N_22170,N_22082);
or U23247 (N_23247,N_22955,N_22508);
nand U23248 (N_23248,N_22298,N_22376);
nor U23249 (N_23249,N_22878,N_22839);
nand U23250 (N_23250,N_22211,N_22857);
xnor U23251 (N_23251,N_22209,N_22744);
and U23252 (N_23252,N_22907,N_22358);
nand U23253 (N_23253,N_22901,N_22734);
and U23254 (N_23254,N_22771,N_22956);
nand U23255 (N_23255,N_22129,N_22533);
nand U23256 (N_23256,N_22951,N_22366);
nor U23257 (N_23257,N_22449,N_22690);
and U23258 (N_23258,N_22223,N_22510);
nor U23259 (N_23259,N_22179,N_22829);
nand U23260 (N_23260,N_22454,N_22297);
and U23261 (N_23261,N_22212,N_22923);
nor U23262 (N_23262,N_22632,N_22225);
or U23263 (N_23263,N_22150,N_22614);
nand U23264 (N_23264,N_22572,N_22139);
xor U23265 (N_23265,N_22296,N_22865);
nand U23266 (N_23266,N_22781,N_22765);
or U23267 (N_23267,N_22959,N_22464);
or U23268 (N_23268,N_22906,N_22638);
xnor U23269 (N_23269,N_22541,N_22033);
nand U23270 (N_23270,N_22763,N_22949);
and U23271 (N_23271,N_22130,N_22368);
nor U23272 (N_23272,N_22576,N_22448);
xor U23273 (N_23273,N_22278,N_22854);
and U23274 (N_23274,N_22343,N_22440);
nor U23275 (N_23275,N_22379,N_22647);
xnor U23276 (N_23276,N_22549,N_22717);
nor U23277 (N_23277,N_22759,N_22773);
nor U23278 (N_23278,N_22097,N_22473);
xor U23279 (N_23279,N_22042,N_22867);
nor U23280 (N_23280,N_22085,N_22022);
nor U23281 (N_23281,N_22475,N_22788);
and U23282 (N_23282,N_22604,N_22507);
or U23283 (N_23283,N_22862,N_22232);
and U23284 (N_23284,N_22117,N_22065);
xor U23285 (N_23285,N_22359,N_22855);
xor U23286 (N_23286,N_22141,N_22902);
xor U23287 (N_23287,N_22545,N_22133);
and U23288 (N_23288,N_22090,N_22568);
and U23289 (N_23289,N_22111,N_22522);
nor U23290 (N_23290,N_22477,N_22392);
nand U23291 (N_23291,N_22720,N_22927);
nor U23292 (N_23292,N_22708,N_22412);
xnor U23293 (N_23293,N_22050,N_22685);
or U23294 (N_23294,N_22064,N_22622);
or U23295 (N_23295,N_22451,N_22640);
nand U23296 (N_23296,N_22446,N_22846);
xnor U23297 (N_23297,N_22790,N_22107);
or U23298 (N_23298,N_22665,N_22414);
xnor U23299 (N_23299,N_22386,N_22169);
xnor U23300 (N_23300,N_22975,N_22835);
nand U23301 (N_23301,N_22913,N_22723);
and U23302 (N_23302,N_22289,N_22210);
and U23303 (N_23303,N_22393,N_22147);
nor U23304 (N_23304,N_22729,N_22365);
or U23305 (N_23305,N_22561,N_22413);
and U23306 (N_23306,N_22926,N_22245);
and U23307 (N_23307,N_22932,N_22877);
and U23308 (N_23308,N_22116,N_22144);
or U23309 (N_23309,N_22388,N_22756);
nand U23310 (N_23310,N_22749,N_22515);
xnor U23311 (N_23311,N_22489,N_22242);
or U23312 (N_23312,N_22875,N_22073);
or U23313 (N_23313,N_22687,N_22990);
or U23314 (N_23314,N_22203,N_22081);
and U23315 (N_23315,N_22390,N_22672);
and U23316 (N_23316,N_22260,N_22478);
and U23317 (N_23317,N_22215,N_22108);
or U23318 (N_23318,N_22112,N_22602);
or U23319 (N_23319,N_22540,N_22820);
nor U23320 (N_23320,N_22904,N_22766);
or U23321 (N_23321,N_22370,N_22313);
xor U23322 (N_23322,N_22880,N_22322);
nor U23323 (N_23323,N_22980,N_22506);
nand U23324 (N_23324,N_22610,N_22554);
or U23325 (N_23325,N_22890,N_22295);
or U23326 (N_23326,N_22356,N_22748);
nand U23327 (N_23327,N_22342,N_22837);
nor U23328 (N_23328,N_22407,N_22861);
and U23329 (N_23329,N_22733,N_22847);
xnor U23330 (N_23330,N_22938,N_22025);
nor U23331 (N_23331,N_22353,N_22029);
and U23332 (N_23332,N_22047,N_22834);
and U23333 (N_23333,N_22431,N_22991);
xor U23334 (N_23334,N_22088,N_22526);
nor U23335 (N_23335,N_22726,N_22504);
and U23336 (N_23336,N_22094,N_22279);
and U23337 (N_23337,N_22010,N_22362);
and U23338 (N_23338,N_22999,N_22498);
nor U23339 (N_23339,N_22799,N_22558);
nand U23340 (N_23340,N_22137,N_22354);
and U23341 (N_23341,N_22419,N_22695);
nor U23342 (N_23342,N_22246,N_22119);
xnor U23343 (N_23343,N_22265,N_22485);
or U23344 (N_23344,N_22071,N_22597);
xnor U23345 (N_23345,N_22401,N_22816);
or U23346 (N_23346,N_22724,N_22668);
nor U23347 (N_23347,N_22791,N_22053);
nor U23348 (N_23348,N_22501,N_22931);
nor U23349 (N_23349,N_22509,N_22027);
nand U23350 (N_23350,N_22411,N_22929);
xor U23351 (N_23351,N_22187,N_22633);
or U23352 (N_23352,N_22189,N_22394);
xnor U23353 (N_23353,N_22058,N_22198);
nand U23354 (N_23354,N_22725,N_22973);
and U23355 (N_23355,N_22217,N_22933);
xnor U23356 (N_23356,N_22794,N_22120);
xnor U23357 (N_23357,N_22583,N_22976);
nand U23358 (N_23358,N_22981,N_22427);
nand U23359 (N_23359,N_22987,N_22624);
nor U23360 (N_23360,N_22755,N_22697);
or U23361 (N_23361,N_22335,N_22077);
or U23362 (N_23362,N_22397,N_22544);
nand U23363 (N_23363,N_22808,N_22525);
nand U23364 (N_23364,N_22807,N_22355);
nand U23365 (N_23365,N_22416,N_22780);
xnor U23366 (N_23366,N_22600,N_22014);
nor U23367 (N_23367,N_22658,N_22115);
nand U23368 (N_23368,N_22294,N_22109);
or U23369 (N_23369,N_22521,N_22019);
nand U23370 (N_23370,N_22470,N_22396);
xnor U23371 (N_23371,N_22743,N_22101);
nand U23372 (N_23372,N_22046,N_22299);
or U23373 (N_23373,N_22712,N_22166);
xnor U23374 (N_23374,N_22831,N_22100);
nor U23375 (N_23375,N_22021,N_22292);
or U23376 (N_23376,N_22680,N_22917);
nand U23377 (N_23377,N_22550,N_22657);
nor U23378 (N_23378,N_22308,N_22186);
xnor U23379 (N_23379,N_22200,N_22304);
and U23380 (N_23380,N_22578,N_22838);
nand U23381 (N_23381,N_22336,N_22833);
and U23382 (N_23382,N_22660,N_22581);
or U23383 (N_23383,N_22853,N_22997);
or U23384 (N_23384,N_22806,N_22893);
nor U23385 (N_23385,N_22193,N_22136);
and U23386 (N_23386,N_22303,N_22157);
xor U23387 (N_23387,N_22616,N_22442);
and U23388 (N_23388,N_22592,N_22185);
xnor U23389 (N_23389,N_22122,N_22167);
nor U23390 (N_23390,N_22784,N_22930);
or U23391 (N_23391,N_22779,N_22191);
xor U23392 (N_23392,N_22777,N_22425);
and U23393 (N_23393,N_22769,N_22499);
and U23394 (N_23394,N_22471,N_22048);
xnor U23395 (N_23395,N_22079,N_22199);
and U23396 (N_23396,N_22953,N_22900);
xnor U23397 (N_23397,N_22662,N_22005);
nand U23398 (N_23398,N_22012,N_22490);
nand U23399 (N_23399,N_22331,N_22032);
or U23400 (N_23400,N_22132,N_22300);
nand U23401 (N_23401,N_22161,N_22040);
nand U23402 (N_23402,N_22714,N_22676);
xor U23403 (N_23403,N_22741,N_22195);
nor U23404 (N_23404,N_22887,N_22290);
nor U23405 (N_23405,N_22001,N_22288);
and U23406 (N_23406,N_22374,N_22970);
nand U23407 (N_23407,N_22405,N_22452);
and U23408 (N_23408,N_22798,N_22444);
nor U23409 (N_23409,N_22237,N_22570);
and U23410 (N_23410,N_22009,N_22013);
xor U23411 (N_23411,N_22326,N_22479);
nor U23412 (N_23412,N_22516,N_22679);
nor U23413 (N_23413,N_22639,N_22621);
xor U23414 (N_23414,N_22043,N_22268);
xor U23415 (N_23415,N_22174,N_22086);
and U23416 (N_23416,N_22546,N_22159);
or U23417 (N_23417,N_22513,N_22124);
nor U23418 (N_23418,N_22275,N_22761);
xnor U23419 (N_23419,N_22892,N_22611);
or U23420 (N_23420,N_22426,N_22098);
xnor U23421 (N_23421,N_22850,N_22706);
and U23422 (N_23422,N_22731,N_22972);
nor U23423 (N_23423,N_22735,N_22937);
and U23424 (N_23424,N_22403,N_22856);
or U23425 (N_23425,N_22387,N_22882);
xnor U23426 (N_23426,N_22538,N_22860);
and U23427 (N_23427,N_22054,N_22625);
xor U23428 (N_23428,N_22125,N_22641);
xnor U23429 (N_23429,N_22559,N_22333);
nand U23430 (N_23430,N_22828,N_22113);
nand U23431 (N_23431,N_22327,N_22589);
xor U23432 (N_23432,N_22811,N_22273);
xor U23433 (N_23433,N_22587,N_22235);
or U23434 (N_23434,N_22172,N_22567);
xor U23435 (N_23435,N_22361,N_22914);
nand U23436 (N_23436,N_22577,N_22579);
nor U23437 (N_23437,N_22606,N_22176);
and U23438 (N_23438,N_22966,N_22277);
xor U23439 (N_23439,N_22459,N_22825);
or U23440 (N_23440,N_22915,N_22645);
nor U23441 (N_23441,N_22493,N_22138);
nor U23442 (N_23442,N_22259,N_22709);
or U23443 (N_23443,N_22548,N_22204);
nand U23444 (N_23444,N_22747,N_22417);
or U23445 (N_23445,N_22945,N_22134);
xnor U23446 (N_23446,N_22334,N_22357);
nand U23447 (N_23447,N_22110,N_22008);
xnor U23448 (N_23448,N_22306,N_22140);
xor U23449 (N_23449,N_22240,N_22698);
nand U23450 (N_23450,N_22618,N_22031);
or U23451 (N_23451,N_22629,N_22716);
and U23452 (N_23452,N_22764,N_22518);
and U23453 (N_23453,N_22928,N_22269);
xor U23454 (N_23454,N_22517,N_22201);
xnor U23455 (N_23455,N_22952,N_22072);
and U23456 (N_23456,N_22423,N_22536);
and U23457 (N_23457,N_22889,N_22894);
nor U23458 (N_23458,N_22222,N_22701);
nor U23459 (N_23459,N_22126,N_22462);
xor U23460 (N_23460,N_22851,N_22069);
and U23461 (N_23461,N_22084,N_22812);
nor U23462 (N_23462,N_22768,N_22920);
xor U23463 (N_23463,N_22194,N_22580);
nand U23464 (N_23464,N_22918,N_22736);
nand U23465 (N_23465,N_22317,N_22154);
nor U23466 (N_23466,N_22722,N_22623);
or U23467 (N_23467,N_22243,N_22371);
or U23468 (N_23468,N_22635,N_22601);
nand U23469 (N_23469,N_22344,N_22797);
or U23470 (N_23470,N_22940,N_22822);
and U23471 (N_23471,N_22055,N_22018);
and U23472 (N_23472,N_22226,N_22497);
or U23473 (N_23473,N_22039,N_22628);
xnor U23474 (N_23474,N_22916,N_22487);
nor U23475 (N_23475,N_22787,N_22523);
nor U23476 (N_23476,N_22373,N_22229);
or U23477 (N_23477,N_22165,N_22011);
xor U23478 (N_23478,N_22646,N_22704);
or U23479 (N_23479,N_22049,N_22389);
or U23480 (N_23480,N_22858,N_22380);
and U23481 (N_23481,N_22350,N_22253);
nand U23482 (N_23482,N_22429,N_22263);
nor U23483 (N_23483,N_22977,N_22994);
nor U23484 (N_23484,N_22562,N_22802);
or U23485 (N_23485,N_22560,N_22128);
or U23486 (N_23486,N_22757,N_22817);
nor U23487 (N_23487,N_22468,N_22753);
nand U23488 (N_23488,N_22480,N_22758);
nand U23489 (N_23489,N_22691,N_22026);
or U23490 (N_23490,N_22059,N_22912);
and U23491 (N_23491,N_22321,N_22219);
and U23492 (N_23492,N_22800,N_22627);
nor U23493 (N_23493,N_22348,N_22715);
or U23494 (N_23494,N_22895,N_22944);
or U23495 (N_23495,N_22512,N_22686);
or U23496 (N_23496,N_22104,N_22924);
nor U23497 (N_23497,N_22637,N_22143);
xor U23498 (N_23498,N_22339,N_22168);
or U23499 (N_23499,N_22809,N_22872);
nand U23500 (N_23500,N_22234,N_22541);
nor U23501 (N_23501,N_22704,N_22922);
or U23502 (N_23502,N_22221,N_22018);
nand U23503 (N_23503,N_22557,N_22894);
nor U23504 (N_23504,N_22444,N_22299);
and U23505 (N_23505,N_22996,N_22889);
nor U23506 (N_23506,N_22286,N_22808);
nor U23507 (N_23507,N_22308,N_22735);
xnor U23508 (N_23508,N_22847,N_22266);
nand U23509 (N_23509,N_22337,N_22344);
or U23510 (N_23510,N_22512,N_22415);
nand U23511 (N_23511,N_22420,N_22561);
nand U23512 (N_23512,N_22544,N_22234);
nor U23513 (N_23513,N_22163,N_22334);
nor U23514 (N_23514,N_22373,N_22702);
or U23515 (N_23515,N_22022,N_22408);
nand U23516 (N_23516,N_22602,N_22730);
and U23517 (N_23517,N_22143,N_22142);
or U23518 (N_23518,N_22287,N_22617);
nor U23519 (N_23519,N_22310,N_22226);
and U23520 (N_23520,N_22371,N_22166);
xnor U23521 (N_23521,N_22293,N_22320);
nor U23522 (N_23522,N_22925,N_22383);
xnor U23523 (N_23523,N_22378,N_22035);
or U23524 (N_23524,N_22689,N_22477);
xnor U23525 (N_23525,N_22375,N_22125);
or U23526 (N_23526,N_22435,N_22946);
xor U23527 (N_23527,N_22425,N_22491);
and U23528 (N_23528,N_22386,N_22019);
and U23529 (N_23529,N_22226,N_22516);
and U23530 (N_23530,N_22552,N_22883);
xnor U23531 (N_23531,N_22877,N_22321);
nand U23532 (N_23532,N_22491,N_22035);
nor U23533 (N_23533,N_22188,N_22103);
xnor U23534 (N_23534,N_22196,N_22044);
nand U23535 (N_23535,N_22801,N_22103);
or U23536 (N_23536,N_22691,N_22061);
or U23537 (N_23537,N_22590,N_22907);
xnor U23538 (N_23538,N_22032,N_22433);
and U23539 (N_23539,N_22645,N_22446);
or U23540 (N_23540,N_22616,N_22417);
or U23541 (N_23541,N_22776,N_22410);
xor U23542 (N_23542,N_22971,N_22868);
nor U23543 (N_23543,N_22348,N_22003);
nor U23544 (N_23544,N_22219,N_22197);
nor U23545 (N_23545,N_22111,N_22922);
nor U23546 (N_23546,N_22362,N_22125);
or U23547 (N_23547,N_22557,N_22196);
and U23548 (N_23548,N_22738,N_22947);
and U23549 (N_23549,N_22063,N_22834);
or U23550 (N_23550,N_22798,N_22991);
and U23551 (N_23551,N_22509,N_22966);
nand U23552 (N_23552,N_22986,N_22977);
and U23553 (N_23553,N_22632,N_22520);
xnor U23554 (N_23554,N_22106,N_22441);
and U23555 (N_23555,N_22783,N_22893);
and U23556 (N_23556,N_22557,N_22389);
xor U23557 (N_23557,N_22056,N_22857);
nand U23558 (N_23558,N_22039,N_22748);
or U23559 (N_23559,N_22693,N_22648);
or U23560 (N_23560,N_22955,N_22857);
and U23561 (N_23561,N_22860,N_22663);
and U23562 (N_23562,N_22643,N_22716);
nand U23563 (N_23563,N_22244,N_22032);
nand U23564 (N_23564,N_22855,N_22487);
and U23565 (N_23565,N_22399,N_22881);
xor U23566 (N_23566,N_22924,N_22345);
xnor U23567 (N_23567,N_22147,N_22246);
nor U23568 (N_23568,N_22011,N_22227);
nor U23569 (N_23569,N_22451,N_22540);
nand U23570 (N_23570,N_22066,N_22513);
xor U23571 (N_23571,N_22834,N_22869);
and U23572 (N_23572,N_22888,N_22355);
nor U23573 (N_23573,N_22479,N_22301);
and U23574 (N_23574,N_22936,N_22963);
or U23575 (N_23575,N_22872,N_22052);
nor U23576 (N_23576,N_22038,N_22538);
or U23577 (N_23577,N_22521,N_22225);
nand U23578 (N_23578,N_22536,N_22673);
or U23579 (N_23579,N_22946,N_22865);
nor U23580 (N_23580,N_22294,N_22886);
xor U23581 (N_23581,N_22995,N_22704);
nor U23582 (N_23582,N_22648,N_22844);
nand U23583 (N_23583,N_22280,N_22521);
xor U23584 (N_23584,N_22713,N_22152);
or U23585 (N_23585,N_22008,N_22565);
xnor U23586 (N_23586,N_22099,N_22230);
and U23587 (N_23587,N_22997,N_22385);
nor U23588 (N_23588,N_22739,N_22050);
nand U23589 (N_23589,N_22503,N_22947);
or U23590 (N_23590,N_22425,N_22901);
nand U23591 (N_23591,N_22626,N_22814);
nand U23592 (N_23592,N_22535,N_22587);
or U23593 (N_23593,N_22492,N_22815);
or U23594 (N_23594,N_22229,N_22004);
nor U23595 (N_23595,N_22885,N_22695);
xor U23596 (N_23596,N_22594,N_22816);
xor U23597 (N_23597,N_22567,N_22324);
nor U23598 (N_23598,N_22981,N_22995);
xnor U23599 (N_23599,N_22822,N_22561);
nor U23600 (N_23600,N_22557,N_22210);
nand U23601 (N_23601,N_22962,N_22430);
and U23602 (N_23602,N_22908,N_22390);
nor U23603 (N_23603,N_22067,N_22796);
xnor U23604 (N_23604,N_22946,N_22507);
nor U23605 (N_23605,N_22142,N_22315);
nand U23606 (N_23606,N_22919,N_22845);
xor U23607 (N_23607,N_22104,N_22679);
nor U23608 (N_23608,N_22527,N_22430);
nand U23609 (N_23609,N_22575,N_22943);
xor U23610 (N_23610,N_22384,N_22099);
nor U23611 (N_23611,N_22272,N_22049);
nor U23612 (N_23612,N_22037,N_22704);
nand U23613 (N_23613,N_22383,N_22969);
xnor U23614 (N_23614,N_22950,N_22263);
and U23615 (N_23615,N_22566,N_22181);
and U23616 (N_23616,N_22595,N_22434);
and U23617 (N_23617,N_22848,N_22041);
or U23618 (N_23618,N_22403,N_22391);
and U23619 (N_23619,N_22911,N_22939);
and U23620 (N_23620,N_22602,N_22358);
and U23621 (N_23621,N_22915,N_22749);
nand U23622 (N_23622,N_22766,N_22948);
and U23623 (N_23623,N_22063,N_22432);
and U23624 (N_23624,N_22644,N_22710);
nand U23625 (N_23625,N_22846,N_22532);
xor U23626 (N_23626,N_22492,N_22545);
nor U23627 (N_23627,N_22339,N_22927);
xor U23628 (N_23628,N_22998,N_22127);
or U23629 (N_23629,N_22348,N_22591);
and U23630 (N_23630,N_22560,N_22533);
or U23631 (N_23631,N_22878,N_22901);
xor U23632 (N_23632,N_22392,N_22708);
and U23633 (N_23633,N_22310,N_22986);
nor U23634 (N_23634,N_22768,N_22296);
and U23635 (N_23635,N_22348,N_22457);
xnor U23636 (N_23636,N_22893,N_22881);
nor U23637 (N_23637,N_22808,N_22450);
nand U23638 (N_23638,N_22577,N_22004);
nor U23639 (N_23639,N_22869,N_22903);
nor U23640 (N_23640,N_22812,N_22531);
and U23641 (N_23641,N_22445,N_22385);
xor U23642 (N_23642,N_22811,N_22805);
or U23643 (N_23643,N_22443,N_22496);
xnor U23644 (N_23644,N_22296,N_22970);
nand U23645 (N_23645,N_22396,N_22015);
nand U23646 (N_23646,N_22742,N_22212);
xor U23647 (N_23647,N_22749,N_22697);
xnor U23648 (N_23648,N_22131,N_22732);
or U23649 (N_23649,N_22410,N_22400);
nor U23650 (N_23650,N_22639,N_22263);
nand U23651 (N_23651,N_22360,N_22771);
and U23652 (N_23652,N_22077,N_22642);
nor U23653 (N_23653,N_22180,N_22684);
nand U23654 (N_23654,N_22468,N_22785);
or U23655 (N_23655,N_22481,N_22749);
and U23656 (N_23656,N_22996,N_22828);
and U23657 (N_23657,N_22768,N_22567);
nand U23658 (N_23658,N_22070,N_22515);
and U23659 (N_23659,N_22944,N_22248);
and U23660 (N_23660,N_22452,N_22928);
nor U23661 (N_23661,N_22832,N_22636);
nor U23662 (N_23662,N_22322,N_22406);
nand U23663 (N_23663,N_22633,N_22083);
and U23664 (N_23664,N_22152,N_22795);
nand U23665 (N_23665,N_22868,N_22796);
and U23666 (N_23666,N_22367,N_22760);
xnor U23667 (N_23667,N_22186,N_22138);
xnor U23668 (N_23668,N_22063,N_22629);
nand U23669 (N_23669,N_22128,N_22812);
nand U23670 (N_23670,N_22583,N_22155);
nand U23671 (N_23671,N_22660,N_22546);
nor U23672 (N_23672,N_22905,N_22844);
or U23673 (N_23673,N_22115,N_22854);
xnor U23674 (N_23674,N_22940,N_22625);
nand U23675 (N_23675,N_22712,N_22676);
nor U23676 (N_23676,N_22267,N_22060);
or U23677 (N_23677,N_22379,N_22943);
or U23678 (N_23678,N_22275,N_22421);
or U23679 (N_23679,N_22748,N_22058);
and U23680 (N_23680,N_22528,N_22985);
nand U23681 (N_23681,N_22082,N_22047);
or U23682 (N_23682,N_22452,N_22647);
nor U23683 (N_23683,N_22373,N_22554);
xnor U23684 (N_23684,N_22083,N_22919);
nor U23685 (N_23685,N_22737,N_22569);
or U23686 (N_23686,N_22213,N_22096);
nand U23687 (N_23687,N_22459,N_22960);
and U23688 (N_23688,N_22460,N_22624);
nor U23689 (N_23689,N_22994,N_22370);
nand U23690 (N_23690,N_22287,N_22772);
and U23691 (N_23691,N_22162,N_22059);
and U23692 (N_23692,N_22862,N_22084);
xnor U23693 (N_23693,N_22479,N_22632);
and U23694 (N_23694,N_22760,N_22691);
nand U23695 (N_23695,N_22406,N_22635);
nand U23696 (N_23696,N_22769,N_22569);
nand U23697 (N_23697,N_22863,N_22410);
xnor U23698 (N_23698,N_22273,N_22282);
or U23699 (N_23699,N_22647,N_22686);
xnor U23700 (N_23700,N_22206,N_22759);
nand U23701 (N_23701,N_22701,N_22839);
xnor U23702 (N_23702,N_22806,N_22971);
nand U23703 (N_23703,N_22371,N_22111);
and U23704 (N_23704,N_22923,N_22174);
xnor U23705 (N_23705,N_22315,N_22837);
and U23706 (N_23706,N_22921,N_22587);
and U23707 (N_23707,N_22104,N_22664);
or U23708 (N_23708,N_22424,N_22218);
nor U23709 (N_23709,N_22838,N_22833);
nor U23710 (N_23710,N_22259,N_22889);
nor U23711 (N_23711,N_22974,N_22582);
nor U23712 (N_23712,N_22945,N_22600);
nand U23713 (N_23713,N_22254,N_22186);
and U23714 (N_23714,N_22687,N_22922);
xor U23715 (N_23715,N_22285,N_22782);
nand U23716 (N_23716,N_22776,N_22412);
nand U23717 (N_23717,N_22291,N_22621);
nand U23718 (N_23718,N_22610,N_22803);
nand U23719 (N_23719,N_22028,N_22517);
nand U23720 (N_23720,N_22476,N_22879);
xnor U23721 (N_23721,N_22909,N_22586);
and U23722 (N_23722,N_22957,N_22268);
nand U23723 (N_23723,N_22642,N_22867);
and U23724 (N_23724,N_22017,N_22684);
nor U23725 (N_23725,N_22227,N_22922);
or U23726 (N_23726,N_22845,N_22961);
nand U23727 (N_23727,N_22048,N_22648);
xor U23728 (N_23728,N_22344,N_22696);
and U23729 (N_23729,N_22503,N_22938);
and U23730 (N_23730,N_22042,N_22706);
and U23731 (N_23731,N_22161,N_22581);
or U23732 (N_23732,N_22548,N_22080);
and U23733 (N_23733,N_22680,N_22664);
xnor U23734 (N_23734,N_22905,N_22170);
and U23735 (N_23735,N_22176,N_22719);
nand U23736 (N_23736,N_22059,N_22292);
nand U23737 (N_23737,N_22716,N_22420);
nor U23738 (N_23738,N_22425,N_22286);
or U23739 (N_23739,N_22663,N_22611);
nand U23740 (N_23740,N_22215,N_22698);
or U23741 (N_23741,N_22735,N_22902);
or U23742 (N_23742,N_22929,N_22807);
nand U23743 (N_23743,N_22297,N_22579);
or U23744 (N_23744,N_22642,N_22890);
nor U23745 (N_23745,N_22984,N_22589);
nor U23746 (N_23746,N_22308,N_22014);
or U23747 (N_23747,N_22004,N_22598);
xor U23748 (N_23748,N_22521,N_22109);
xor U23749 (N_23749,N_22234,N_22551);
or U23750 (N_23750,N_22071,N_22983);
nand U23751 (N_23751,N_22764,N_22521);
and U23752 (N_23752,N_22807,N_22040);
nand U23753 (N_23753,N_22115,N_22098);
nand U23754 (N_23754,N_22028,N_22174);
and U23755 (N_23755,N_22266,N_22572);
nand U23756 (N_23756,N_22427,N_22175);
or U23757 (N_23757,N_22326,N_22422);
xor U23758 (N_23758,N_22206,N_22295);
nand U23759 (N_23759,N_22405,N_22995);
xnor U23760 (N_23760,N_22972,N_22377);
nor U23761 (N_23761,N_22185,N_22164);
or U23762 (N_23762,N_22127,N_22884);
nand U23763 (N_23763,N_22875,N_22941);
or U23764 (N_23764,N_22518,N_22717);
and U23765 (N_23765,N_22804,N_22646);
nand U23766 (N_23766,N_22924,N_22809);
or U23767 (N_23767,N_22801,N_22258);
or U23768 (N_23768,N_22547,N_22450);
nor U23769 (N_23769,N_22830,N_22919);
xnor U23770 (N_23770,N_22705,N_22934);
and U23771 (N_23771,N_22439,N_22022);
xor U23772 (N_23772,N_22627,N_22821);
nand U23773 (N_23773,N_22906,N_22917);
and U23774 (N_23774,N_22283,N_22651);
nor U23775 (N_23775,N_22356,N_22033);
nand U23776 (N_23776,N_22008,N_22940);
xor U23777 (N_23777,N_22439,N_22374);
or U23778 (N_23778,N_22723,N_22481);
nor U23779 (N_23779,N_22215,N_22445);
and U23780 (N_23780,N_22020,N_22836);
and U23781 (N_23781,N_22974,N_22700);
nand U23782 (N_23782,N_22560,N_22894);
or U23783 (N_23783,N_22207,N_22834);
or U23784 (N_23784,N_22876,N_22306);
nor U23785 (N_23785,N_22476,N_22248);
nor U23786 (N_23786,N_22806,N_22626);
xnor U23787 (N_23787,N_22374,N_22242);
or U23788 (N_23788,N_22522,N_22134);
nor U23789 (N_23789,N_22025,N_22893);
and U23790 (N_23790,N_22495,N_22999);
xnor U23791 (N_23791,N_22737,N_22753);
and U23792 (N_23792,N_22171,N_22960);
nand U23793 (N_23793,N_22897,N_22923);
and U23794 (N_23794,N_22207,N_22975);
nor U23795 (N_23795,N_22426,N_22743);
nor U23796 (N_23796,N_22853,N_22670);
xor U23797 (N_23797,N_22305,N_22207);
and U23798 (N_23798,N_22724,N_22320);
nor U23799 (N_23799,N_22908,N_22949);
nor U23800 (N_23800,N_22016,N_22683);
nor U23801 (N_23801,N_22577,N_22771);
and U23802 (N_23802,N_22993,N_22258);
nor U23803 (N_23803,N_22950,N_22589);
and U23804 (N_23804,N_22537,N_22694);
nor U23805 (N_23805,N_22050,N_22171);
nand U23806 (N_23806,N_22831,N_22988);
or U23807 (N_23807,N_22896,N_22125);
xor U23808 (N_23808,N_22615,N_22099);
xor U23809 (N_23809,N_22576,N_22378);
or U23810 (N_23810,N_22175,N_22992);
nand U23811 (N_23811,N_22129,N_22652);
and U23812 (N_23812,N_22601,N_22021);
nor U23813 (N_23813,N_22964,N_22238);
nor U23814 (N_23814,N_22216,N_22581);
nor U23815 (N_23815,N_22593,N_22421);
nor U23816 (N_23816,N_22470,N_22324);
nor U23817 (N_23817,N_22418,N_22918);
and U23818 (N_23818,N_22877,N_22209);
or U23819 (N_23819,N_22693,N_22859);
nor U23820 (N_23820,N_22383,N_22708);
or U23821 (N_23821,N_22584,N_22895);
or U23822 (N_23822,N_22952,N_22006);
nand U23823 (N_23823,N_22286,N_22315);
xor U23824 (N_23824,N_22716,N_22530);
or U23825 (N_23825,N_22861,N_22566);
and U23826 (N_23826,N_22830,N_22393);
nor U23827 (N_23827,N_22827,N_22316);
xnor U23828 (N_23828,N_22167,N_22343);
xnor U23829 (N_23829,N_22921,N_22264);
nand U23830 (N_23830,N_22118,N_22552);
nand U23831 (N_23831,N_22842,N_22938);
and U23832 (N_23832,N_22590,N_22843);
nand U23833 (N_23833,N_22276,N_22740);
and U23834 (N_23834,N_22146,N_22737);
xor U23835 (N_23835,N_22311,N_22609);
and U23836 (N_23836,N_22611,N_22147);
xnor U23837 (N_23837,N_22602,N_22861);
nand U23838 (N_23838,N_22733,N_22586);
or U23839 (N_23839,N_22498,N_22181);
xnor U23840 (N_23840,N_22316,N_22175);
and U23841 (N_23841,N_22899,N_22350);
and U23842 (N_23842,N_22173,N_22352);
nand U23843 (N_23843,N_22271,N_22714);
xor U23844 (N_23844,N_22077,N_22367);
xor U23845 (N_23845,N_22352,N_22858);
and U23846 (N_23846,N_22254,N_22013);
or U23847 (N_23847,N_22374,N_22373);
and U23848 (N_23848,N_22531,N_22567);
or U23849 (N_23849,N_22332,N_22219);
and U23850 (N_23850,N_22200,N_22037);
or U23851 (N_23851,N_22856,N_22537);
or U23852 (N_23852,N_22524,N_22880);
or U23853 (N_23853,N_22130,N_22297);
nor U23854 (N_23854,N_22567,N_22680);
xnor U23855 (N_23855,N_22126,N_22323);
nand U23856 (N_23856,N_22658,N_22424);
or U23857 (N_23857,N_22104,N_22260);
or U23858 (N_23858,N_22249,N_22995);
and U23859 (N_23859,N_22543,N_22899);
or U23860 (N_23860,N_22728,N_22586);
xnor U23861 (N_23861,N_22126,N_22259);
xor U23862 (N_23862,N_22807,N_22015);
and U23863 (N_23863,N_22903,N_22779);
or U23864 (N_23864,N_22339,N_22891);
or U23865 (N_23865,N_22797,N_22763);
xnor U23866 (N_23866,N_22282,N_22474);
or U23867 (N_23867,N_22193,N_22859);
nand U23868 (N_23868,N_22202,N_22515);
xnor U23869 (N_23869,N_22069,N_22101);
or U23870 (N_23870,N_22304,N_22447);
and U23871 (N_23871,N_22476,N_22323);
nand U23872 (N_23872,N_22913,N_22595);
xor U23873 (N_23873,N_22021,N_22796);
or U23874 (N_23874,N_22613,N_22769);
and U23875 (N_23875,N_22526,N_22174);
xor U23876 (N_23876,N_22887,N_22666);
or U23877 (N_23877,N_22272,N_22325);
nor U23878 (N_23878,N_22934,N_22775);
xor U23879 (N_23879,N_22121,N_22128);
nand U23880 (N_23880,N_22589,N_22000);
or U23881 (N_23881,N_22054,N_22204);
xnor U23882 (N_23882,N_22586,N_22700);
xnor U23883 (N_23883,N_22946,N_22589);
and U23884 (N_23884,N_22767,N_22368);
or U23885 (N_23885,N_22131,N_22671);
nor U23886 (N_23886,N_22899,N_22032);
nor U23887 (N_23887,N_22348,N_22461);
nand U23888 (N_23888,N_22246,N_22752);
xor U23889 (N_23889,N_22654,N_22650);
or U23890 (N_23890,N_22022,N_22149);
or U23891 (N_23891,N_22625,N_22254);
xor U23892 (N_23892,N_22272,N_22518);
nand U23893 (N_23893,N_22555,N_22666);
nand U23894 (N_23894,N_22006,N_22731);
xor U23895 (N_23895,N_22328,N_22329);
nor U23896 (N_23896,N_22318,N_22395);
or U23897 (N_23897,N_22503,N_22550);
nand U23898 (N_23898,N_22878,N_22598);
or U23899 (N_23899,N_22656,N_22927);
nand U23900 (N_23900,N_22385,N_22552);
xnor U23901 (N_23901,N_22730,N_22546);
and U23902 (N_23902,N_22266,N_22015);
nor U23903 (N_23903,N_22781,N_22992);
and U23904 (N_23904,N_22287,N_22000);
nand U23905 (N_23905,N_22960,N_22993);
xor U23906 (N_23906,N_22416,N_22107);
xnor U23907 (N_23907,N_22988,N_22732);
nand U23908 (N_23908,N_22587,N_22922);
xnor U23909 (N_23909,N_22373,N_22886);
or U23910 (N_23910,N_22861,N_22649);
or U23911 (N_23911,N_22148,N_22486);
nor U23912 (N_23912,N_22772,N_22037);
nor U23913 (N_23913,N_22929,N_22120);
nor U23914 (N_23914,N_22937,N_22787);
and U23915 (N_23915,N_22215,N_22781);
and U23916 (N_23916,N_22762,N_22858);
or U23917 (N_23917,N_22481,N_22236);
or U23918 (N_23918,N_22395,N_22437);
and U23919 (N_23919,N_22665,N_22219);
nand U23920 (N_23920,N_22879,N_22795);
xnor U23921 (N_23921,N_22860,N_22294);
and U23922 (N_23922,N_22659,N_22482);
xor U23923 (N_23923,N_22390,N_22683);
nand U23924 (N_23924,N_22642,N_22101);
nor U23925 (N_23925,N_22575,N_22712);
and U23926 (N_23926,N_22631,N_22399);
and U23927 (N_23927,N_22873,N_22761);
and U23928 (N_23928,N_22468,N_22378);
xor U23929 (N_23929,N_22354,N_22519);
nand U23930 (N_23930,N_22764,N_22324);
nor U23931 (N_23931,N_22217,N_22392);
nand U23932 (N_23932,N_22638,N_22605);
xor U23933 (N_23933,N_22744,N_22092);
or U23934 (N_23934,N_22936,N_22650);
or U23935 (N_23935,N_22831,N_22052);
and U23936 (N_23936,N_22134,N_22847);
nand U23937 (N_23937,N_22655,N_22585);
or U23938 (N_23938,N_22389,N_22183);
xnor U23939 (N_23939,N_22617,N_22384);
or U23940 (N_23940,N_22302,N_22852);
xnor U23941 (N_23941,N_22557,N_22509);
nand U23942 (N_23942,N_22579,N_22063);
or U23943 (N_23943,N_22529,N_22900);
nor U23944 (N_23944,N_22957,N_22577);
nand U23945 (N_23945,N_22441,N_22770);
or U23946 (N_23946,N_22969,N_22929);
nand U23947 (N_23947,N_22426,N_22198);
nor U23948 (N_23948,N_22936,N_22428);
nand U23949 (N_23949,N_22320,N_22667);
nand U23950 (N_23950,N_22307,N_22395);
xnor U23951 (N_23951,N_22918,N_22308);
xnor U23952 (N_23952,N_22563,N_22590);
nand U23953 (N_23953,N_22754,N_22116);
or U23954 (N_23954,N_22206,N_22305);
nor U23955 (N_23955,N_22220,N_22216);
and U23956 (N_23956,N_22507,N_22567);
xnor U23957 (N_23957,N_22338,N_22871);
or U23958 (N_23958,N_22166,N_22172);
or U23959 (N_23959,N_22794,N_22044);
and U23960 (N_23960,N_22048,N_22567);
and U23961 (N_23961,N_22711,N_22845);
and U23962 (N_23962,N_22089,N_22907);
or U23963 (N_23963,N_22104,N_22149);
and U23964 (N_23964,N_22619,N_22782);
and U23965 (N_23965,N_22664,N_22774);
nand U23966 (N_23966,N_22963,N_22666);
and U23967 (N_23967,N_22144,N_22021);
or U23968 (N_23968,N_22117,N_22083);
nand U23969 (N_23969,N_22234,N_22568);
and U23970 (N_23970,N_22795,N_22083);
and U23971 (N_23971,N_22013,N_22932);
and U23972 (N_23972,N_22440,N_22441);
and U23973 (N_23973,N_22776,N_22496);
and U23974 (N_23974,N_22697,N_22644);
and U23975 (N_23975,N_22621,N_22466);
and U23976 (N_23976,N_22292,N_22031);
or U23977 (N_23977,N_22033,N_22353);
and U23978 (N_23978,N_22288,N_22941);
nor U23979 (N_23979,N_22701,N_22359);
nand U23980 (N_23980,N_22865,N_22185);
nand U23981 (N_23981,N_22355,N_22623);
nor U23982 (N_23982,N_22242,N_22529);
and U23983 (N_23983,N_22976,N_22953);
nor U23984 (N_23984,N_22055,N_22711);
or U23985 (N_23985,N_22040,N_22846);
nand U23986 (N_23986,N_22220,N_22588);
xnor U23987 (N_23987,N_22246,N_22839);
and U23988 (N_23988,N_22390,N_22426);
or U23989 (N_23989,N_22287,N_22624);
nor U23990 (N_23990,N_22649,N_22090);
nand U23991 (N_23991,N_22027,N_22630);
nor U23992 (N_23992,N_22277,N_22658);
nand U23993 (N_23993,N_22260,N_22234);
xnor U23994 (N_23994,N_22104,N_22881);
nand U23995 (N_23995,N_22939,N_22599);
or U23996 (N_23996,N_22780,N_22302);
xnor U23997 (N_23997,N_22790,N_22173);
and U23998 (N_23998,N_22660,N_22421);
and U23999 (N_23999,N_22591,N_22823);
nand U24000 (N_24000,N_23128,N_23442);
xnor U24001 (N_24001,N_23552,N_23394);
and U24002 (N_24002,N_23162,N_23400);
xor U24003 (N_24003,N_23401,N_23321);
or U24004 (N_24004,N_23123,N_23558);
nor U24005 (N_24005,N_23948,N_23513);
and U24006 (N_24006,N_23397,N_23872);
xor U24007 (N_24007,N_23979,N_23031);
or U24008 (N_24008,N_23177,N_23146);
nand U24009 (N_24009,N_23821,N_23911);
nand U24010 (N_24010,N_23882,N_23228);
nand U24011 (N_24011,N_23745,N_23692);
and U24012 (N_24012,N_23055,N_23797);
and U24013 (N_24013,N_23187,N_23635);
nor U24014 (N_24014,N_23761,N_23830);
xor U24015 (N_24015,N_23325,N_23013);
nand U24016 (N_24016,N_23993,N_23071);
and U24017 (N_24017,N_23267,N_23600);
or U24018 (N_24018,N_23689,N_23158);
nor U24019 (N_24019,N_23290,N_23305);
nor U24020 (N_24020,N_23721,N_23022);
or U24021 (N_24021,N_23493,N_23097);
nor U24022 (N_24022,N_23214,N_23512);
xnor U24023 (N_24023,N_23215,N_23796);
xor U24024 (N_24024,N_23679,N_23540);
or U24025 (N_24025,N_23915,N_23323);
or U24026 (N_24026,N_23186,N_23580);
nor U24027 (N_24027,N_23391,N_23634);
and U24028 (N_24028,N_23793,N_23842);
nor U24029 (N_24029,N_23962,N_23230);
or U24030 (N_24030,N_23567,N_23182);
nand U24031 (N_24031,N_23856,N_23181);
nor U24032 (N_24032,N_23585,N_23180);
nor U24033 (N_24033,N_23362,N_23795);
or U24034 (N_24034,N_23218,N_23366);
nor U24035 (N_24035,N_23563,N_23294);
nand U24036 (N_24036,N_23899,N_23212);
xnor U24037 (N_24037,N_23672,N_23981);
nor U24038 (N_24038,N_23084,N_23254);
nor U24039 (N_24039,N_23419,N_23386);
nor U24040 (N_24040,N_23010,N_23229);
nand U24041 (N_24041,N_23869,N_23346);
nor U24042 (N_24042,N_23538,N_23127);
and U24043 (N_24043,N_23355,N_23803);
or U24044 (N_24044,N_23311,N_23969);
or U24045 (N_24045,N_23933,N_23769);
xnor U24046 (N_24046,N_23877,N_23601);
or U24047 (N_24047,N_23562,N_23086);
and U24048 (N_24048,N_23518,N_23833);
nand U24049 (N_24049,N_23437,N_23360);
nand U24050 (N_24050,N_23713,N_23896);
xnor U24051 (N_24051,N_23317,N_23973);
nand U24052 (N_24052,N_23114,N_23787);
xor U24053 (N_24053,N_23396,N_23952);
nand U24054 (N_24054,N_23619,N_23859);
xnor U24055 (N_24055,N_23659,N_23488);
nor U24056 (N_24056,N_23646,N_23725);
or U24057 (N_24057,N_23372,N_23749);
nand U24058 (N_24058,N_23931,N_23698);
nand U24059 (N_24059,N_23261,N_23221);
and U24060 (N_24060,N_23040,N_23174);
nand U24061 (N_24061,N_23737,N_23522);
nand U24062 (N_24062,N_23154,N_23198);
xnor U24063 (N_24063,N_23743,N_23908);
or U24064 (N_24064,N_23754,N_23039);
xnor U24065 (N_24065,N_23895,N_23890);
and U24066 (N_24066,N_23062,N_23387);
nand U24067 (N_24067,N_23544,N_23253);
nand U24068 (N_24068,N_23104,N_23138);
nand U24069 (N_24069,N_23392,N_23612);
nor U24070 (N_24070,N_23695,N_23320);
nand U24071 (N_24071,N_23349,N_23383);
nand U24072 (N_24072,N_23555,N_23056);
xnor U24073 (N_24073,N_23237,N_23523);
nand U24074 (N_24074,N_23265,N_23696);
nand U24075 (N_24075,N_23959,N_23331);
and U24076 (N_24076,N_23773,N_23451);
and U24077 (N_24077,N_23395,N_23638);
and U24078 (N_24078,N_23077,N_23007);
or U24079 (N_24079,N_23117,N_23474);
nor U24080 (N_24080,N_23465,N_23731);
and U24081 (N_24081,N_23751,N_23529);
and U24082 (N_24082,N_23818,N_23102);
nand U24083 (N_24083,N_23134,N_23867);
or U24084 (N_24084,N_23834,N_23388);
xnor U24085 (N_24085,N_23614,N_23233);
and U24086 (N_24086,N_23945,N_23408);
nor U24087 (N_24087,N_23376,N_23716);
nor U24088 (N_24088,N_23135,N_23964);
xor U24089 (N_24089,N_23380,N_23333);
and U24090 (N_24090,N_23817,N_23815);
nor U24091 (N_24091,N_23242,N_23559);
nor U24092 (N_24092,N_23652,N_23357);
nor U24093 (N_24093,N_23501,N_23748);
nand U24094 (N_24094,N_23412,N_23129);
nor U24095 (N_24095,N_23155,N_23790);
nor U24096 (N_24096,N_23940,N_23209);
xor U24097 (N_24097,N_23938,N_23923);
nor U24098 (N_24098,N_23750,N_23204);
xnor U24099 (N_24099,N_23137,N_23484);
and U24100 (N_24100,N_23873,N_23482);
nand U24101 (N_24101,N_23537,N_23998);
or U24102 (N_24102,N_23416,N_23917);
or U24103 (N_24103,N_23628,N_23206);
nor U24104 (N_24104,N_23100,N_23650);
nand U24105 (N_24105,N_23132,N_23897);
nor U24106 (N_24106,N_23531,N_23076);
or U24107 (N_24107,N_23173,N_23118);
nand U24108 (N_24108,N_23201,N_23006);
nor U24109 (N_24109,N_23561,N_23343);
or U24110 (N_24110,N_23660,N_23857);
and U24111 (N_24111,N_23739,N_23615);
or U24112 (N_24112,N_23322,N_23900);
or U24113 (N_24113,N_23089,N_23985);
or U24114 (N_24114,N_23169,N_23812);
nor U24115 (N_24115,N_23093,N_23516);
or U24116 (N_24116,N_23337,N_23498);
xor U24117 (N_24117,N_23142,N_23080);
nand U24118 (N_24118,N_23909,N_23423);
and U24119 (N_24119,N_23051,N_23732);
nand U24120 (N_24120,N_23426,N_23236);
or U24121 (N_24121,N_23185,N_23618);
or U24122 (N_24122,N_23359,N_23608);
and U24123 (N_24123,N_23534,N_23175);
and U24124 (N_24124,N_23920,N_23956);
and U24125 (N_24125,N_23642,N_23048);
or U24126 (N_24126,N_23499,N_23332);
xnor U24127 (N_24127,N_23092,N_23999);
nor U24128 (N_24128,N_23313,N_23472);
or U24129 (N_24129,N_23109,N_23502);
or U24130 (N_24130,N_23219,N_23826);
or U24131 (N_24131,N_23008,N_23862);
nand U24132 (N_24132,N_23700,N_23982);
nor U24133 (N_24133,N_23947,N_23832);
and U24134 (N_24134,N_23514,N_23927);
or U24135 (N_24135,N_23837,N_23085);
nand U24136 (N_24136,N_23564,N_23028);
nor U24137 (N_24137,N_23464,N_23373);
and U24138 (N_24138,N_23605,N_23840);
or U24139 (N_24139,N_23458,N_23543);
nor U24140 (N_24140,N_23225,N_23786);
nand U24141 (N_24141,N_23038,N_23064);
nor U24142 (N_24142,N_23811,N_23413);
nand U24143 (N_24143,N_23798,N_23888);
nand U24144 (N_24144,N_23918,N_23824);
nand U24145 (N_24145,N_23620,N_23167);
nand U24146 (N_24146,N_23001,N_23189);
xnor U24147 (N_24147,N_23196,N_23418);
nand U24148 (N_24148,N_23264,N_23505);
and U24149 (N_24149,N_23588,N_23686);
or U24150 (N_24150,N_23298,N_23338);
xor U24151 (N_24151,N_23677,N_23368);
and U24152 (N_24152,N_23508,N_23115);
nor U24153 (N_24153,N_23524,N_23525);
and U24154 (N_24154,N_23980,N_23825);
nor U24155 (N_24155,N_23466,N_23053);
nand U24156 (N_24156,N_23170,N_23772);
or U24157 (N_24157,N_23542,N_23327);
and U24158 (N_24158,N_23319,N_23411);
xnor U24159 (N_24159,N_23611,N_23777);
xor U24160 (N_24160,N_23655,N_23549);
xnor U24161 (N_24161,N_23406,N_23178);
nand U24162 (N_24162,N_23766,N_23326);
or U24163 (N_24163,N_23708,N_23557);
and U24164 (N_24164,N_23823,N_23255);
nand U24165 (N_24165,N_23934,N_23044);
and U24166 (N_24166,N_23710,N_23768);
nand U24167 (N_24167,N_23607,N_23141);
xor U24168 (N_24168,N_23260,N_23393);
or U24169 (N_24169,N_23208,N_23030);
nand U24170 (N_24170,N_23992,N_23669);
and U24171 (N_24171,N_23262,N_23756);
nand U24172 (N_24172,N_23658,N_23238);
xnor U24173 (N_24173,N_23148,N_23143);
xor U24174 (N_24174,N_23520,N_23375);
and U24175 (N_24175,N_23415,N_23664);
nor U24176 (N_24176,N_23239,N_23626);
nor U24177 (N_24177,N_23893,N_23417);
and U24178 (N_24178,N_23921,N_23203);
or U24179 (N_24179,N_23342,N_23272);
xnor U24180 (N_24180,N_23582,N_23858);
nand U24181 (N_24181,N_23977,N_23340);
xor U24182 (N_24182,N_23407,N_23584);
nor U24183 (N_24183,N_23469,N_23259);
nand U24184 (N_24184,N_23547,N_23816);
xnor U24185 (N_24185,N_23976,N_23481);
nand U24186 (N_24186,N_23263,N_23479);
xor U24187 (N_24187,N_23081,N_23160);
and U24188 (N_24188,N_23110,N_23729);
and U24189 (N_24189,N_23112,N_23461);
nand U24190 (N_24190,N_23054,N_23536);
and U24191 (N_24191,N_23596,N_23864);
and U24192 (N_24192,N_23785,N_23309);
nor U24193 (N_24193,N_23901,N_23865);
nor U24194 (N_24194,N_23978,N_23234);
and U24195 (N_24195,N_23113,N_23667);
and U24196 (N_24196,N_23657,N_23995);
nor U24197 (N_24197,N_23356,N_23870);
nor U24198 (N_24198,N_23647,N_23566);
nor U24199 (N_24199,N_23345,N_23714);
nand U24200 (N_24200,N_23736,N_23783);
or U24201 (N_24201,N_23533,N_23497);
xnor U24202 (N_24202,N_23266,N_23404);
nand U24203 (N_24203,N_23009,N_23776);
and U24204 (N_24204,N_23223,N_23444);
xor U24205 (N_24205,N_23063,N_23315);
or U24206 (N_24206,N_23511,N_23382);
or U24207 (N_24207,N_23431,N_23220);
xnor U24208 (N_24208,N_23656,N_23595);
xor U24209 (N_24209,N_23485,N_23105);
or U24210 (N_24210,N_23662,N_23292);
nand U24211 (N_24211,N_23688,N_23427);
and U24212 (N_24212,N_23029,N_23649);
nor U24213 (N_24213,N_23843,N_23043);
or U24214 (N_24214,N_23280,N_23441);
and U24215 (N_24215,N_23344,N_23727);
and U24216 (N_24216,N_23300,N_23591);
or U24217 (N_24217,N_23072,N_23301);
xnor U24218 (N_24218,N_23248,N_23719);
or U24219 (N_24219,N_23951,N_23020);
xor U24220 (N_24220,N_23032,N_23389);
nand U24221 (N_24221,N_23963,N_23720);
and U24222 (N_24222,N_23057,N_23507);
and U24223 (N_24223,N_23633,N_23994);
nor U24224 (N_24224,N_23090,N_23930);
or U24225 (N_24225,N_23434,N_23252);
nor U24226 (N_24226,N_23027,N_23358);
nor U24227 (N_24227,N_23578,N_23207);
and U24228 (N_24228,N_23851,N_23712);
or U24229 (N_24229,N_23717,N_23576);
nor U24230 (N_24230,N_23569,N_23047);
or U24231 (N_24231,N_23473,N_23274);
nand U24232 (N_24232,N_23452,N_23735);
or U24233 (N_24233,N_23589,N_23004);
or U24234 (N_24234,N_23884,N_23486);
nor U24235 (N_24235,N_23402,N_23445);
or U24236 (N_24236,N_23804,N_23887);
xor U24237 (N_24237,N_23892,N_23651);
or U24238 (N_24238,N_23806,N_23829);
and U24239 (N_24239,N_23370,N_23810);
nor U24240 (N_24240,N_23405,N_23521);
nor U24241 (N_24241,N_23035,N_23779);
or U24242 (N_24242,N_23988,N_23450);
nand U24243 (N_24243,N_23183,N_23805);
xor U24244 (N_24244,N_23781,N_23184);
and U24245 (N_24245,N_23984,N_23987);
or U24246 (N_24246,N_23989,N_23583);
and U24247 (N_24247,N_23526,N_23673);
or U24248 (N_24248,N_23838,N_23025);
and U24249 (N_24249,N_23590,N_23453);
nor U24250 (N_24250,N_23866,N_23310);
or U24251 (N_24251,N_23049,N_23839);
xor U24252 (N_24252,N_23703,N_23966);
nor U24253 (N_24253,N_23621,N_23188);
or U24254 (N_24254,N_23088,N_23456);
xor U24255 (N_24255,N_23885,N_23683);
nor U24256 (N_24256,N_23844,N_23381);
or U24257 (N_24257,N_23771,N_23630);
xnor U24258 (N_24258,N_23161,N_23079);
xnor U24259 (N_24259,N_23075,N_23384);
or U24260 (N_24260,N_23070,N_23489);
nor U24261 (N_24261,N_23530,N_23699);
and U24262 (N_24262,N_23849,N_23707);
or U24263 (N_24263,N_23983,N_23907);
and U24264 (N_24264,N_23496,N_23133);
nand U24265 (N_24265,N_23641,N_23819);
xor U24266 (N_24266,N_23510,N_23961);
nand U24267 (N_24267,N_23680,N_23939);
nor U24268 (N_24268,N_23997,N_23879);
and U24269 (N_24269,N_23316,N_23448);
or U24270 (N_24270,N_23140,N_23875);
xnor U24271 (N_24271,N_23414,N_23506);
nor U24272 (N_24272,N_23269,N_23250);
or U24273 (N_24273,N_23808,N_23836);
and U24274 (N_24274,N_23653,N_23420);
nor U24275 (N_24275,N_23121,N_23046);
nand U24276 (N_24276,N_23024,N_23483);
nor U24277 (N_24277,N_23432,N_23539);
nand U24278 (N_24278,N_23016,N_23960);
nand U24279 (N_24279,N_23443,N_23568);
nand U24280 (N_24280,N_23706,N_23166);
and U24281 (N_24281,N_23058,N_23603);
or U24282 (N_24282,N_23718,N_23813);
or U24283 (N_24283,N_23033,N_23554);
xor U24284 (N_24284,N_23936,N_23285);
nor U24285 (N_24285,N_23059,N_23855);
and U24286 (N_24286,N_23066,N_23026);
nand U24287 (N_24287,N_23232,N_23436);
nand U24288 (N_24288,N_23809,N_23447);
nor U24289 (N_24289,N_23041,N_23957);
or U24290 (N_24290,N_23303,N_23289);
nor U24291 (N_24291,N_23517,N_23403);
and U24292 (N_24292,N_23487,N_23586);
nor U24293 (N_24293,N_23050,N_23631);
and U24294 (N_24294,N_23799,N_23975);
and U24295 (N_24295,N_23814,N_23663);
xnor U24296 (N_24296,N_23841,N_23205);
and U24297 (N_24297,N_23425,N_23774);
xor U24298 (N_24298,N_23922,N_23082);
xnor U24299 (N_24299,N_23150,N_23691);
nor U24300 (N_24300,N_23730,N_23347);
and U24301 (N_24301,N_23495,N_23752);
and U24302 (N_24302,N_23324,N_23307);
xor U24303 (N_24303,N_23579,N_23935);
or U24304 (N_24304,N_23304,N_23288);
xor U24305 (N_24305,N_23446,N_23409);
nand U24306 (N_24306,N_23968,N_23330);
and U24307 (N_24307,N_23928,N_23172);
xor U24308 (N_24308,N_23361,N_23565);
or U24309 (N_24309,N_23868,N_23932);
nand U24310 (N_24310,N_23728,N_23021);
and U24311 (N_24311,N_23942,N_23216);
nor U24312 (N_24312,N_23244,N_23599);
or U24313 (N_24313,N_23629,N_23850);
and U24314 (N_24314,N_23763,N_23535);
nand U24315 (N_24315,N_23871,N_23954);
or U24316 (N_24316,N_23256,N_23023);
nor U24317 (N_24317,N_23996,N_23211);
or U24318 (N_24318,N_23424,N_23293);
nand U24319 (N_24319,N_23891,N_23067);
nand U24320 (N_24320,N_23733,N_23297);
or U24321 (N_24321,N_23709,N_23011);
nand U24322 (N_24322,N_23492,N_23831);
nor U24323 (N_24323,N_23617,N_23224);
xnor U24324 (N_24324,N_23351,N_23697);
nand U24325 (N_24325,N_23005,N_23478);
nand U24326 (N_24326,N_23152,N_23622);
nand U24327 (N_24327,N_23801,N_23898);
xor U24328 (N_24328,N_23098,N_23246);
nand U24329 (N_24329,N_23273,N_23723);
nor U24330 (N_24330,N_23480,N_23278);
nand U24331 (N_24331,N_23581,N_23197);
xnor U24332 (N_24332,N_23339,N_23210);
nand U24333 (N_24333,N_23971,N_23822);
nand U24334 (N_24334,N_23861,N_23678);
xnor U24335 (N_24335,N_23247,N_23083);
and U24336 (N_24336,N_23528,N_23845);
and U24337 (N_24337,N_23126,N_23107);
nand U24338 (N_24338,N_23758,N_23640);
nor U24339 (N_24339,N_23550,N_23546);
nand U24340 (N_24340,N_23572,N_23190);
xnor U24341 (N_24341,N_23880,N_23609);
or U24342 (N_24342,N_23509,N_23958);
xor U24343 (N_24343,N_23592,N_23457);
nand U24344 (N_24344,N_23778,N_23095);
or U24345 (N_24345,N_23295,N_23715);
nand U24346 (N_24346,N_23746,N_23283);
or U24347 (N_24347,N_23570,N_23974);
xor U24348 (N_24348,N_23352,N_23950);
nand U24349 (N_24349,N_23052,N_23639);
nor U24350 (N_24350,N_23937,N_23671);
nand U24351 (N_24351,N_23296,N_23091);
nor U24352 (N_24352,N_23078,N_23666);
or U24353 (N_24353,N_23541,N_23257);
xor U24354 (N_24354,N_23335,N_23848);
nand U24355 (N_24355,N_23598,N_23643);
xor U24356 (N_24356,N_23243,N_23902);
and U24357 (N_24357,N_23328,N_23227);
nand U24358 (N_24358,N_23757,N_23788);
and U24359 (N_24359,N_23860,N_23287);
and U24360 (N_24360,N_23863,N_23759);
or U24361 (N_24361,N_23705,N_23199);
or U24362 (N_24362,N_23835,N_23604);
and U24363 (N_24363,N_23916,N_23103);
and U24364 (N_24364,N_23284,N_23551);
nor U24365 (N_24365,N_23770,N_23740);
or U24366 (N_24366,N_23645,N_23675);
or U24367 (N_24367,N_23925,N_23874);
xor U24368 (N_24368,N_23744,N_23202);
nand U24369 (N_24369,N_23245,N_23422);
nand U24370 (N_24370,N_23171,N_23363);
nor U24371 (N_24371,N_23654,N_23610);
and U24372 (N_24372,N_23676,N_23073);
and U24373 (N_24373,N_23440,N_23354);
xnor U24374 (N_24374,N_23704,N_23820);
nand U24375 (N_24375,N_23099,N_23632);
xnor U24376 (N_24376,N_23852,N_23130);
and U24377 (N_24377,N_23241,N_23784);
nand U24378 (N_24378,N_23792,N_23828);
and U24379 (N_24379,N_23306,N_23943);
and U24380 (N_24380,N_23045,N_23847);
or U24381 (N_24381,N_23762,N_23924);
and U24382 (N_24382,N_23379,N_23151);
xor U24383 (N_24383,N_23159,N_23136);
nor U24384 (N_24384,N_23460,N_23722);
nand U24385 (N_24385,N_23069,N_23760);
nor U24386 (N_24386,N_23794,N_23575);
nor U24387 (N_24387,N_23314,N_23015);
or U24388 (N_24388,N_23251,N_23019);
nor U24389 (N_24389,N_23494,N_23556);
nor U24390 (N_24390,N_23991,N_23854);
and U24391 (N_24391,N_23017,N_23800);
nand U24392 (N_24392,N_23527,N_23623);
xnor U24393 (N_24393,N_23276,N_23421);
or U24394 (N_24394,N_23467,N_23277);
nand U24395 (N_24395,N_23462,N_23912);
and U24396 (N_24396,N_23606,N_23702);
nand U24397 (N_24397,N_23226,N_23120);
or U24398 (N_24398,N_23299,N_23553);
nor U24399 (N_24399,N_23341,N_23385);
nand U24400 (N_24400,N_23500,N_23560);
or U24401 (N_24401,N_23275,N_23613);
and U24402 (N_24402,N_23986,N_23881);
nor U24403 (N_24403,N_23764,N_23122);
or U24404 (N_24404,N_23665,N_23889);
or U24405 (N_24405,N_23428,N_23944);
and U24406 (N_24406,N_23491,N_23222);
or U24407 (N_24407,N_23597,N_23116);
or U24408 (N_24408,N_23690,N_23377);
nor U24409 (N_24409,N_23399,N_23574);
nor U24410 (N_24410,N_23302,N_23477);
xnor U24411 (N_24411,N_23217,N_23687);
or U24412 (N_24412,N_23904,N_23374);
nand U24413 (N_24413,N_23545,N_23061);
nand U24414 (N_24414,N_23681,N_23648);
nand U24415 (N_24415,N_23433,N_23775);
or U24416 (N_24416,N_23972,N_23701);
and U24417 (N_24417,N_23350,N_23475);
or U24418 (N_24418,N_23685,N_23616);
or U24419 (N_24419,N_23571,N_23390);
nor U24420 (N_24420,N_23439,N_23176);
nor U24421 (N_24421,N_23191,N_23194);
and U24422 (N_24422,N_23213,N_23131);
and U24423 (N_24423,N_23883,N_23753);
nand U24424 (N_24424,N_23515,N_23037);
or U24425 (N_24425,N_23455,N_23532);
nor U24426 (N_24426,N_23694,N_23802);
or U24427 (N_24427,N_23036,N_23724);
xor U24428 (N_24428,N_23168,N_23476);
nand U24429 (N_24429,N_23014,N_23258);
xnor U24430 (N_24430,N_23065,N_23249);
xnor U24431 (N_24431,N_23336,N_23929);
nand U24432 (N_24432,N_23593,N_23153);
nand U24433 (N_24433,N_23192,N_23734);
nor U24434 (N_24434,N_23353,N_23449);
nand U24435 (N_24435,N_23435,N_23636);
xnor U24436 (N_24436,N_23738,N_23711);
nand U24437 (N_24437,N_23003,N_23573);
nor U24438 (N_24438,N_23119,N_23970);
and U24439 (N_24439,N_23068,N_23410);
nor U24440 (N_24440,N_23602,N_23459);
xnor U24441 (N_24441,N_23438,N_23644);
or U24442 (N_24442,N_23096,N_23125);
or U24443 (N_24443,N_23741,N_23108);
nor U24444 (N_24444,N_23018,N_23145);
and U24445 (N_24445,N_23780,N_23548);
nand U24446 (N_24446,N_23378,N_23329);
and U24447 (N_24447,N_23074,N_23164);
nand U24448 (N_24448,N_23594,N_23637);
xnor U24449 (N_24449,N_23002,N_23504);
nor U24450 (N_24450,N_23454,N_23334);
xnor U24451 (N_24451,N_23470,N_23919);
and U24452 (N_24452,N_23625,N_23106);
nand U24453 (N_24453,N_23430,N_23312);
or U24454 (N_24454,N_23367,N_23903);
and U24455 (N_24455,N_23807,N_23094);
nand U24456 (N_24456,N_23577,N_23042);
xor U24457 (N_24457,N_23364,N_23846);
nor U24458 (N_24458,N_23965,N_23291);
and U24459 (N_24459,N_23894,N_23124);
or U24460 (N_24460,N_23471,N_23627);
nor U24461 (N_24461,N_23286,N_23782);
nor U24462 (N_24462,N_23905,N_23318);
or U24463 (N_24463,N_23910,N_23726);
and U24464 (N_24464,N_23139,N_23941);
nand U24465 (N_24465,N_23149,N_23886);
nor U24466 (N_24466,N_23767,N_23468);
xor U24467 (N_24467,N_23490,N_23791);
or U24468 (N_24468,N_23670,N_23165);
or U24469 (N_24469,N_23913,N_23661);
or U24470 (N_24470,N_23953,N_23503);
or U24471 (N_24471,N_23365,N_23827);
nor U24472 (N_24472,N_23926,N_23398);
or U24473 (N_24473,N_23281,N_23684);
nand U24474 (N_24474,N_23878,N_23111);
nand U24475 (N_24475,N_23270,N_23101);
nor U24476 (N_24476,N_23587,N_23371);
or U24477 (N_24477,N_23279,N_23060);
and U24478 (N_24478,N_23348,N_23179);
nand U24479 (N_24479,N_23157,N_23853);
nor U24480 (N_24480,N_23949,N_23240);
or U24481 (N_24481,N_23682,N_23463);
xnor U24482 (N_24482,N_23193,N_23163);
xnor U24483 (N_24483,N_23268,N_23369);
and U24484 (N_24484,N_23955,N_23012);
and U24485 (N_24485,N_23308,N_23914);
nor U24486 (N_24486,N_23147,N_23034);
nor U24487 (N_24487,N_23624,N_23144);
xor U24488 (N_24488,N_23789,N_23668);
or U24489 (N_24489,N_23195,N_23087);
and U24490 (N_24490,N_23990,N_23156);
and U24491 (N_24491,N_23429,N_23946);
xor U24492 (N_24492,N_23765,N_23235);
or U24493 (N_24493,N_23519,N_23282);
or U24494 (N_24494,N_23906,N_23876);
xnor U24495 (N_24495,N_23271,N_23000);
and U24496 (N_24496,N_23674,N_23231);
or U24497 (N_24497,N_23200,N_23742);
nor U24498 (N_24498,N_23693,N_23747);
nand U24499 (N_24499,N_23967,N_23755);
nand U24500 (N_24500,N_23930,N_23495);
xor U24501 (N_24501,N_23767,N_23375);
or U24502 (N_24502,N_23445,N_23398);
nor U24503 (N_24503,N_23710,N_23245);
nand U24504 (N_24504,N_23258,N_23986);
and U24505 (N_24505,N_23822,N_23666);
or U24506 (N_24506,N_23775,N_23577);
xor U24507 (N_24507,N_23220,N_23298);
and U24508 (N_24508,N_23311,N_23306);
xnor U24509 (N_24509,N_23179,N_23710);
or U24510 (N_24510,N_23475,N_23526);
xnor U24511 (N_24511,N_23641,N_23874);
or U24512 (N_24512,N_23695,N_23222);
nand U24513 (N_24513,N_23368,N_23372);
and U24514 (N_24514,N_23168,N_23021);
nand U24515 (N_24515,N_23268,N_23158);
or U24516 (N_24516,N_23202,N_23190);
nor U24517 (N_24517,N_23269,N_23034);
and U24518 (N_24518,N_23543,N_23320);
and U24519 (N_24519,N_23558,N_23895);
and U24520 (N_24520,N_23498,N_23832);
nor U24521 (N_24521,N_23506,N_23279);
nor U24522 (N_24522,N_23559,N_23589);
xnor U24523 (N_24523,N_23546,N_23067);
xor U24524 (N_24524,N_23606,N_23766);
and U24525 (N_24525,N_23320,N_23628);
and U24526 (N_24526,N_23995,N_23882);
nor U24527 (N_24527,N_23602,N_23306);
nand U24528 (N_24528,N_23596,N_23815);
nand U24529 (N_24529,N_23894,N_23493);
nor U24530 (N_24530,N_23674,N_23597);
xnor U24531 (N_24531,N_23226,N_23113);
and U24532 (N_24532,N_23198,N_23197);
or U24533 (N_24533,N_23879,N_23781);
and U24534 (N_24534,N_23842,N_23972);
nand U24535 (N_24535,N_23688,N_23073);
nand U24536 (N_24536,N_23555,N_23565);
xnor U24537 (N_24537,N_23526,N_23973);
or U24538 (N_24538,N_23958,N_23471);
xnor U24539 (N_24539,N_23569,N_23570);
nand U24540 (N_24540,N_23320,N_23170);
nand U24541 (N_24541,N_23941,N_23581);
nand U24542 (N_24542,N_23304,N_23868);
nor U24543 (N_24543,N_23221,N_23056);
and U24544 (N_24544,N_23459,N_23719);
nand U24545 (N_24545,N_23615,N_23446);
nor U24546 (N_24546,N_23653,N_23382);
or U24547 (N_24547,N_23924,N_23174);
or U24548 (N_24548,N_23594,N_23598);
or U24549 (N_24549,N_23177,N_23800);
or U24550 (N_24550,N_23534,N_23108);
xnor U24551 (N_24551,N_23821,N_23682);
and U24552 (N_24552,N_23876,N_23775);
or U24553 (N_24553,N_23126,N_23740);
and U24554 (N_24554,N_23299,N_23454);
nand U24555 (N_24555,N_23468,N_23993);
and U24556 (N_24556,N_23112,N_23214);
or U24557 (N_24557,N_23097,N_23076);
nor U24558 (N_24558,N_23128,N_23542);
or U24559 (N_24559,N_23528,N_23517);
nand U24560 (N_24560,N_23319,N_23231);
xor U24561 (N_24561,N_23631,N_23320);
xnor U24562 (N_24562,N_23398,N_23645);
nand U24563 (N_24563,N_23556,N_23550);
nand U24564 (N_24564,N_23807,N_23425);
and U24565 (N_24565,N_23691,N_23856);
or U24566 (N_24566,N_23143,N_23767);
xnor U24567 (N_24567,N_23817,N_23684);
or U24568 (N_24568,N_23665,N_23339);
xnor U24569 (N_24569,N_23382,N_23530);
nor U24570 (N_24570,N_23975,N_23832);
or U24571 (N_24571,N_23996,N_23833);
or U24572 (N_24572,N_23333,N_23501);
or U24573 (N_24573,N_23802,N_23179);
or U24574 (N_24574,N_23455,N_23873);
xnor U24575 (N_24575,N_23398,N_23080);
and U24576 (N_24576,N_23192,N_23516);
xnor U24577 (N_24577,N_23015,N_23840);
or U24578 (N_24578,N_23228,N_23054);
xnor U24579 (N_24579,N_23952,N_23310);
nand U24580 (N_24580,N_23658,N_23051);
and U24581 (N_24581,N_23135,N_23875);
nand U24582 (N_24582,N_23866,N_23314);
xnor U24583 (N_24583,N_23665,N_23528);
nor U24584 (N_24584,N_23750,N_23257);
or U24585 (N_24585,N_23724,N_23232);
nor U24586 (N_24586,N_23544,N_23400);
and U24587 (N_24587,N_23625,N_23784);
xor U24588 (N_24588,N_23314,N_23355);
nand U24589 (N_24589,N_23392,N_23409);
or U24590 (N_24590,N_23243,N_23960);
nand U24591 (N_24591,N_23481,N_23455);
or U24592 (N_24592,N_23203,N_23326);
nand U24593 (N_24593,N_23022,N_23682);
nor U24594 (N_24594,N_23489,N_23033);
or U24595 (N_24595,N_23990,N_23185);
nand U24596 (N_24596,N_23941,N_23905);
nor U24597 (N_24597,N_23056,N_23833);
nand U24598 (N_24598,N_23428,N_23170);
and U24599 (N_24599,N_23517,N_23510);
and U24600 (N_24600,N_23245,N_23532);
xnor U24601 (N_24601,N_23560,N_23447);
xor U24602 (N_24602,N_23261,N_23498);
or U24603 (N_24603,N_23508,N_23414);
xnor U24604 (N_24604,N_23431,N_23358);
xnor U24605 (N_24605,N_23092,N_23822);
nor U24606 (N_24606,N_23801,N_23329);
nor U24607 (N_24607,N_23395,N_23950);
nand U24608 (N_24608,N_23864,N_23081);
xnor U24609 (N_24609,N_23663,N_23090);
nor U24610 (N_24610,N_23448,N_23107);
or U24611 (N_24611,N_23174,N_23336);
nor U24612 (N_24612,N_23802,N_23160);
xnor U24613 (N_24613,N_23404,N_23664);
nor U24614 (N_24614,N_23858,N_23983);
or U24615 (N_24615,N_23165,N_23756);
nand U24616 (N_24616,N_23171,N_23678);
xor U24617 (N_24617,N_23291,N_23935);
and U24618 (N_24618,N_23878,N_23754);
and U24619 (N_24619,N_23717,N_23310);
and U24620 (N_24620,N_23070,N_23635);
xor U24621 (N_24621,N_23408,N_23782);
xor U24622 (N_24622,N_23421,N_23449);
or U24623 (N_24623,N_23245,N_23143);
xor U24624 (N_24624,N_23894,N_23414);
and U24625 (N_24625,N_23999,N_23544);
xor U24626 (N_24626,N_23294,N_23938);
or U24627 (N_24627,N_23718,N_23569);
nor U24628 (N_24628,N_23944,N_23090);
nand U24629 (N_24629,N_23229,N_23966);
xnor U24630 (N_24630,N_23795,N_23191);
nor U24631 (N_24631,N_23405,N_23582);
or U24632 (N_24632,N_23973,N_23459);
nand U24633 (N_24633,N_23554,N_23301);
and U24634 (N_24634,N_23358,N_23298);
and U24635 (N_24635,N_23082,N_23340);
nand U24636 (N_24636,N_23817,N_23673);
nor U24637 (N_24637,N_23937,N_23356);
nor U24638 (N_24638,N_23989,N_23089);
or U24639 (N_24639,N_23696,N_23497);
nand U24640 (N_24640,N_23652,N_23867);
and U24641 (N_24641,N_23639,N_23757);
or U24642 (N_24642,N_23636,N_23432);
xnor U24643 (N_24643,N_23994,N_23098);
or U24644 (N_24644,N_23048,N_23013);
or U24645 (N_24645,N_23176,N_23796);
and U24646 (N_24646,N_23989,N_23424);
and U24647 (N_24647,N_23859,N_23504);
xor U24648 (N_24648,N_23157,N_23559);
or U24649 (N_24649,N_23897,N_23733);
nor U24650 (N_24650,N_23044,N_23191);
nand U24651 (N_24651,N_23232,N_23027);
xor U24652 (N_24652,N_23351,N_23700);
nor U24653 (N_24653,N_23490,N_23150);
nor U24654 (N_24654,N_23856,N_23585);
nor U24655 (N_24655,N_23878,N_23418);
and U24656 (N_24656,N_23716,N_23679);
xor U24657 (N_24657,N_23643,N_23198);
xnor U24658 (N_24658,N_23230,N_23011);
nor U24659 (N_24659,N_23421,N_23314);
nor U24660 (N_24660,N_23105,N_23607);
or U24661 (N_24661,N_23707,N_23942);
or U24662 (N_24662,N_23464,N_23026);
nand U24663 (N_24663,N_23414,N_23410);
nand U24664 (N_24664,N_23934,N_23542);
nor U24665 (N_24665,N_23728,N_23388);
and U24666 (N_24666,N_23610,N_23200);
xor U24667 (N_24667,N_23952,N_23315);
and U24668 (N_24668,N_23032,N_23833);
nand U24669 (N_24669,N_23680,N_23657);
and U24670 (N_24670,N_23609,N_23159);
and U24671 (N_24671,N_23173,N_23317);
or U24672 (N_24672,N_23842,N_23771);
nand U24673 (N_24673,N_23169,N_23657);
and U24674 (N_24674,N_23302,N_23009);
nor U24675 (N_24675,N_23528,N_23144);
and U24676 (N_24676,N_23849,N_23676);
nor U24677 (N_24677,N_23010,N_23123);
nor U24678 (N_24678,N_23766,N_23406);
or U24679 (N_24679,N_23486,N_23877);
and U24680 (N_24680,N_23705,N_23154);
or U24681 (N_24681,N_23545,N_23647);
nand U24682 (N_24682,N_23109,N_23952);
and U24683 (N_24683,N_23462,N_23409);
or U24684 (N_24684,N_23924,N_23245);
nand U24685 (N_24685,N_23509,N_23447);
or U24686 (N_24686,N_23727,N_23722);
nand U24687 (N_24687,N_23310,N_23936);
nor U24688 (N_24688,N_23233,N_23357);
and U24689 (N_24689,N_23771,N_23359);
nand U24690 (N_24690,N_23059,N_23369);
nand U24691 (N_24691,N_23372,N_23803);
or U24692 (N_24692,N_23472,N_23562);
nand U24693 (N_24693,N_23006,N_23707);
and U24694 (N_24694,N_23790,N_23457);
and U24695 (N_24695,N_23010,N_23109);
nor U24696 (N_24696,N_23380,N_23633);
nor U24697 (N_24697,N_23097,N_23723);
nor U24698 (N_24698,N_23848,N_23013);
nand U24699 (N_24699,N_23677,N_23465);
or U24700 (N_24700,N_23400,N_23573);
and U24701 (N_24701,N_23521,N_23801);
or U24702 (N_24702,N_23471,N_23829);
nand U24703 (N_24703,N_23004,N_23898);
nand U24704 (N_24704,N_23066,N_23274);
nand U24705 (N_24705,N_23481,N_23917);
xnor U24706 (N_24706,N_23415,N_23638);
or U24707 (N_24707,N_23772,N_23404);
or U24708 (N_24708,N_23764,N_23132);
or U24709 (N_24709,N_23443,N_23658);
xor U24710 (N_24710,N_23950,N_23452);
xnor U24711 (N_24711,N_23237,N_23932);
nand U24712 (N_24712,N_23396,N_23416);
nor U24713 (N_24713,N_23097,N_23857);
and U24714 (N_24714,N_23898,N_23548);
or U24715 (N_24715,N_23960,N_23785);
xnor U24716 (N_24716,N_23226,N_23349);
nand U24717 (N_24717,N_23353,N_23031);
nor U24718 (N_24718,N_23517,N_23956);
nand U24719 (N_24719,N_23425,N_23277);
nand U24720 (N_24720,N_23575,N_23758);
and U24721 (N_24721,N_23282,N_23322);
or U24722 (N_24722,N_23353,N_23003);
nor U24723 (N_24723,N_23932,N_23118);
and U24724 (N_24724,N_23308,N_23667);
xnor U24725 (N_24725,N_23986,N_23529);
nand U24726 (N_24726,N_23784,N_23718);
nor U24727 (N_24727,N_23638,N_23680);
or U24728 (N_24728,N_23307,N_23670);
or U24729 (N_24729,N_23719,N_23781);
xnor U24730 (N_24730,N_23679,N_23499);
and U24731 (N_24731,N_23050,N_23967);
nor U24732 (N_24732,N_23156,N_23021);
nand U24733 (N_24733,N_23993,N_23613);
nor U24734 (N_24734,N_23821,N_23736);
or U24735 (N_24735,N_23168,N_23689);
nand U24736 (N_24736,N_23315,N_23340);
and U24737 (N_24737,N_23127,N_23283);
nand U24738 (N_24738,N_23755,N_23118);
nand U24739 (N_24739,N_23568,N_23094);
and U24740 (N_24740,N_23808,N_23593);
and U24741 (N_24741,N_23807,N_23046);
and U24742 (N_24742,N_23147,N_23342);
nand U24743 (N_24743,N_23683,N_23256);
xor U24744 (N_24744,N_23410,N_23129);
or U24745 (N_24745,N_23761,N_23665);
nor U24746 (N_24746,N_23689,N_23328);
and U24747 (N_24747,N_23541,N_23488);
nor U24748 (N_24748,N_23582,N_23867);
and U24749 (N_24749,N_23061,N_23830);
xor U24750 (N_24750,N_23061,N_23626);
nor U24751 (N_24751,N_23357,N_23133);
and U24752 (N_24752,N_23848,N_23824);
nor U24753 (N_24753,N_23465,N_23736);
nand U24754 (N_24754,N_23628,N_23096);
xnor U24755 (N_24755,N_23729,N_23522);
and U24756 (N_24756,N_23825,N_23219);
and U24757 (N_24757,N_23430,N_23310);
nor U24758 (N_24758,N_23273,N_23600);
or U24759 (N_24759,N_23921,N_23585);
nor U24760 (N_24760,N_23218,N_23620);
nor U24761 (N_24761,N_23627,N_23140);
xor U24762 (N_24762,N_23407,N_23501);
nand U24763 (N_24763,N_23579,N_23700);
nand U24764 (N_24764,N_23928,N_23320);
or U24765 (N_24765,N_23451,N_23461);
and U24766 (N_24766,N_23417,N_23979);
xnor U24767 (N_24767,N_23476,N_23975);
nand U24768 (N_24768,N_23060,N_23910);
nand U24769 (N_24769,N_23899,N_23382);
nand U24770 (N_24770,N_23340,N_23759);
or U24771 (N_24771,N_23064,N_23491);
nor U24772 (N_24772,N_23023,N_23710);
nand U24773 (N_24773,N_23162,N_23513);
nand U24774 (N_24774,N_23089,N_23886);
nor U24775 (N_24775,N_23981,N_23433);
xor U24776 (N_24776,N_23701,N_23301);
nand U24777 (N_24777,N_23953,N_23307);
nor U24778 (N_24778,N_23414,N_23689);
nand U24779 (N_24779,N_23615,N_23629);
and U24780 (N_24780,N_23334,N_23758);
xor U24781 (N_24781,N_23455,N_23655);
or U24782 (N_24782,N_23564,N_23883);
nand U24783 (N_24783,N_23450,N_23290);
and U24784 (N_24784,N_23710,N_23592);
and U24785 (N_24785,N_23068,N_23980);
nand U24786 (N_24786,N_23027,N_23084);
nor U24787 (N_24787,N_23770,N_23088);
and U24788 (N_24788,N_23848,N_23094);
xnor U24789 (N_24789,N_23810,N_23954);
nand U24790 (N_24790,N_23616,N_23841);
nor U24791 (N_24791,N_23938,N_23418);
or U24792 (N_24792,N_23705,N_23326);
nand U24793 (N_24793,N_23805,N_23289);
and U24794 (N_24794,N_23637,N_23999);
and U24795 (N_24795,N_23500,N_23519);
xor U24796 (N_24796,N_23557,N_23467);
nor U24797 (N_24797,N_23551,N_23524);
or U24798 (N_24798,N_23987,N_23638);
or U24799 (N_24799,N_23828,N_23527);
and U24800 (N_24800,N_23077,N_23830);
nand U24801 (N_24801,N_23523,N_23952);
or U24802 (N_24802,N_23947,N_23767);
xnor U24803 (N_24803,N_23696,N_23119);
or U24804 (N_24804,N_23269,N_23876);
and U24805 (N_24805,N_23692,N_23663);
and U24806 (N_24806,N_23300,N_23196);
or U24807 (N_24807,N_23829,N_23349);
and U24808 (N_24808,N_23025,N_23151);
xnor U24809 (N_24809,N_23258,N_23089);
nor U24810 (N_24810,N_23074,N_23362);
nor U24811 (N_24811,N_23293,N_23118);
nor U24812 (N_24812,N_23182,N_23076);
and U24813 (N_24813,N_23141,N_23346);
nand U24814 (N_24814,N_23226,N_23229);
nor U24815 (N_24815,N_23430,N_23009);
and U24816 (N_24816,N_23634,N_23929);
xnor U24817 (N_24817,N_23510,N_23705);
nor U24818 (N_24818,N_23710,N_23063);
xnor U24819 (N_24819,N_23371,N_23867);
nor U24820 (N_24820,N_23788,N_23401);
and U24821 (N_24821,N_23299,N_23585);
nand U24822 (N_24822,N_23022,N_23549);
nand U24823 (N_24823,N_23744,N_23450);
xor U24824 (N_24824,N_23308,N_23706);
nand U24825 (N_24825,N_23276,N_23704);
nor U24826 (N_24826,N_23623,N_23747);
nor U24827 (N_24827,N_23511,N_23578);
xor U24828 (N_24828,N_23507,N_23145);
and U24829 (N_24829,N_23020,N_23833);
xnor U24830 (N_24830,N_23156,N_23385);
or U24831 (N_24831,N_23846,N_23242);
and U24832 (N_24832,N_23668,N_23803);
nand U24833 (N_24833,N_23657,N_23229);
nand U24834 (N_24834,N_23666,N_23915);
xnor U24835 (N_24835,N_23386,N_23823);
xnor U24836 (N_24836,N_23158,N_23130);
xor U24837 (N_24837,N_23355,N_23408);
xor U24838 (N_24838,N_23598,N_23188);
nand U24839 (N_24839,N_23657,N_23574);
or U24840 (N_24840,N_23915,N_23416);
and U24841 (N_24841,N_23795,N_23346);
xnor U24842 (N_24842,N_23447,N_23253);
and U24843 (N_24843,N_23664,N_23525);
xnor U24844 (N_24844,N_23378,N_23287);
nor U24845 (N_24845,N_23657,N_23347);
xor U24846 (N_24846,N_23097,N_23943);
xor U24847 (N_24847,N_23948,N_23366);
nand U24848 (N_24848,N_23528,N_23853);
and U24849 (N_24849,N_23317,N_23884);
and U24850 (N_24850,N_23504,N_23041);
and U24851 (N_24851,N_23997,N_23886);
nand U24852 (N_24852,N_23266,N_23575);
nand U24853 (N_24853,N_23583,N_23851);
xor U24854 (N_24854,N_23004,N_23046);
nor U24855 (N_24855,N_23270,N_23352);
xnor U24856 (N_24856,N_23303,N_23598);
and U24857 (N_24857,N_23340,N_23439);
and U24858 (N_24858,N_23812,N_23562);
and U24859 (N_24859,N_23654,N_23921);
and U24860 (N_24860,N_23281,N_23513);
or U24861 (N_24861,N_23917,N_23824);
nand U24862 (N_24862,N_23419,N_23273);
and U24863 (N_24863,N_23367,N_23744);
or U24864 (N_24864,N_23720,N_23643);
or U24865 (N_24865,N_23191,N_23723);
nor U24866 (N_24866,N_23439,N_23822);
xor U24867 (N_24867,N_23955,N_23628);
and U24868 (N_24868,N_23894,N_23347);
or U24869 (N_24869,N_23605,N_23557);
or U24870 (N_24870,N_23821,N_23913);
and U24871 (N_24871,N_23069,N_23398);
or U24872 (N_24872,N_23655,N_23123);
nor U24873 (N_24873,N_23468,N_23738);
nand U24874 (N_24874,N_23082,N_23553);
or U24875 (N_24875,N_23191,N_23157);
xor U24876 (N_24876,N_23192,N_23407);
nand U24877 (N_24877,N_23560,N_23701);
and U24878 (N_24878,N_23685,N_23099);
or U24879 (N_24879,N_23070,N_23905);
or U24880 (N_24880,N_23087,N_23091);
or U24881 (N_24881,N_23219,N_23637);
or U24882 (N_24882,N_23053,N_23921);
nand U24883 (N_24883,N_23906,N_23278);
xor U24884 (N_24884,N_23898,N_23957);
xnor U24885 (N_24885,N_23738,N_23772);
nand U24886 (N_24886,N_23519,N_23594);
and U24887 (N_24887,N_23380,N_23587);
nand U24888 (N_24888,N_23615,N_23955);
and U24889 (N_24889,N_23849,N_23284);
nor U24890 (N_24890,N_23006,N_23231);
xor U24891 (N_24891,N_23467,N_23857);
nor U24892 (N_24892,N_23519,N_23621);
or U24893 (N_24893,N_23226,N_23438);
or U24894 (N_24894,N_23555,N_23870);
nor U24895 (N_24895,N_23557,N_23098);
or U24896 (N_24896,N_23222,N_23307);
nand U24897 (N_24897,N_23500,N_23074);
nor U24898 (N_24898,N_23771,N_23068);
nor U24899 (N_24899,N_23017,N_23881);
xnor U24900 (N_24900,N_23933,N_23647);
or U24901 (N_24901,N_23344,N_23227);
nor U24902 (N_24902,N_23925,N_23034);
or U24903 (N_24903,N_23891,N_23508);
nand U24904 (N_24904,N_23359,N_23188);
and U24905 (N_24905,N_23330,N_23030);
and U24906 (N_24906,N_23699,N_23428);
xnor U24907 (N_24907,N_23067,N_23232);
xnor U24908 (N_24908,N_23006,N_23112);
xor U24909 (N_24909,N_23840,N_23049);
nand U24910 (N_24910,N_23175,N_23082);
and U24911 (N_24911,N_23994,N_23932);
nand U24912 (N_24912,N_23379,N_23127);
and U24913 (N_24913,N_23983,N_23593);
or U24914 (N_24914,N_23301,N_23456);
nor U24915 (N_24915,N_23724,N_23345);
or U24916 (N_24916,N_23837,N_23693);
nor U24917 (N_24917,N_23996,N_23662);
nand U24918 (N_24918,N_23932,N_23060);
nand U24919 (N_24919,N_23209,N_23392);
nand U24920 (N_24920,N_23436,N_23119);
or U24921 (N_24921,N_23535,N_23362);
nor U24922 (N_24922,N_23705,N_23981);
xor U24923 (N_24923,N_23812,N_23120);
nand U24924 (N_24924,N_23361,N_23665);
and U24925 (N_24925,N_23419,N_23930);
nand U24926 (N_24926,N_23230,N_23798);
and U24927 (N_24927,N_23757,N_23759);
and U24928 (N_24928,N_23727,N_23025);
nor U24929 (N_24929,N_23352,N_23117);
nor U24930 (N_24930,N_23921,N_23363);
xor U24931 (N_24931,N_23045,N_23499);
nand U24932 (N_24932,N_23679,N_23116);
or U24933 (N_24933,N_23256,N_23583);
and U24934 (N_24934,N_23507,N_23319);
nor U24935 (N_24935,N_23121,N_23484);
or U24936 (N_24936,N_23808,N_23728);
nand U24937 (N_24937,N_23260,N_23105);
or U24938 (N_24938,N_23367,N_23094);
or U24939 (N_24939,N_23840,N_23841);
or U24940 (N_24940,N_23603,N_23009);
xor U24941 (N_24941,N_23727,N_23541);
or U24942 (N_24942,N_23393,N_23798);
or U24943 (N_24943,N_23313,N_23922);
nor U24944 (N_24944,N_23410,N_23831);
nor U24945 (N_24945,N_23117,N_23995);
nand U24946 (N_24946,N_23933,N_23350);
nor U24947 (N_24947,N_23099,N_23052);
nor U24948 (N_24948,N_23291,N_23618);
nand U24949 (N_24949,N_23774,N_23004);
and U24950 (N_24950,N_23560,N_23787);
nand U24951 (N_24951,N_23347,N_23129);
nand U24952 (N_24952,N_23284,N_23759);
or U24953 (N_24953,N_23128,N_23741);
nor U24954 (N_24954,N_23974,N_23719);
nor U24955 (N_24955,N_23134,N_23640);
nor U24956 (N_24956,N_23614,N_23577);
nand U24957 (N_24957,N_23879,N_23597);
and U24958 (N_24958,N_23175,N_23034);
xnor U24959 (N_24959,N_23943,N_23893);
and U24960 (N_24960,N_23116,N_23468);
xnor U24961 (N_24961,N_23641,N_23265);
nor U24962 (N_24962,N_23508,N_23787);
nand U24963 (N_24963,N_23877,N_23093);
nor U24964 (N_24964,N_23822,N_23372);
nand U24965 (N_24965,N_23244,N_23035);
nand U24966 (N_24966,N_23361,N_23410);
xor U24967 (N_24967,N_23655,N_23889);
or U24968 (N_24968,N_23890,N_23571);
and U24969 (N_24969,N_23805,N_23927);
xnor U24970 (N_24970,N_23924,N_23459);
xnor U24971 (N_24971,N_23973,N_23431);
nand U24972 (N_24972,N_23780,N_23462);
and U24973 (N_24973,N_23365,N_23993);
nor U24974 (N_24974,N_23311,N_23046);
and U24975 (N_24975,N_23291,N_23341);
or U24976 (N_24976,N_23884,N_23695);
nor U24977 (N_24977,N_23813,N_23039);
xor U24978 (N_24978,N_23764,N_23202);
nand U24979 (N_24979,N_23628,N_23202);
xor U24980 (N_24980,N_23430,N_23733);
and U24981 (N_24981,N_23581,N_23572);
nand U24982 (N_24982,N_23630,N_23504);
and U24983 (N_24983,N_23276,N_23367);
xnor U24984 (N_24984,N_23663,N_23522);
or U24985 (N_24985,N_23907,N_23384);
and U24986 (N_24986,N_23780,N_23297);
or U24987 (N_24987,N_23507,N_23466);
nor U24988 (N_24988,N_23198,N_23750);
nand U24989 (N_24989,N_23076,N_23479);
and U24990 (N_24990,N_23932,N_23607);
and U24991 (N_24991,N_23098,N_23473);
nor U24992 (N_24992,N_23612,N_23802);
nand U24993 (N_24993,N_23027,N_23452);
nand U24994 (N_24994,N_23577,N_23097);
nor U24995 (N_24995,N_23942,N_23564);
and U24996 (N_24996,N_23901,N_23315);
xnor U24997 (N_24997,N_23057,N_23104);
and U24998 (N_24998,N_23228,N_23531);
nand U24999 (N_24999,N_23396,N_23907);
nand U25000 (N_25000,N_24658,N_24759);
xnor U25001 (N_25001,N_24833,N_24348);
and U25002 (N_25002,N_24425,N_24463);
and U25003 (N_25003,N_24068,N_24445);
nor U25004 (N_25004,N_24384,N_24170);
and U25005 (N_25005,N_24060,N_24590);
nor U25006 (N_25006,N_24048,N_24955);
nor U25007 (N_25007,N_24126,N_24930);
nor U25008 (N_25008,N_24529,N_24887);
nor U25009 (N_25009,N_24821,N_24981);
nor U25010 (N_25010,N_24488,N_24376);
or U25011 (N_25011,N_24765,N_24490);
nor U25012 (N_25012,N_24337,N_24233);
or U25013 (N_25013,N_24224,N_24883);
or U25014 (N_25014,N_24547,N_24796);
and U25015 (N_25015,N_24062,N_24303);
nand U25016 (N_25016,N_24896,N_24205);
nor U25017 (N_25017,N_24248,N_24357);
or U25018 (N_25018,N_24631,N_24564);
nor U25019 (N_25019,N_24092,N_24196);
nor U25020 (N_25020,N_24649,N_24360);
and U25021 (N_25021,N_24124,N_24526);
and U25022 (N_25022,N_24667,N_24251);
or U25023 (N_25023,N_24880,N_24652);
or U25024 (N_25024,N_24277,N_24733);
and U25025 (N_25025,N_24449,N_24640);
nand U25026 (N_25026,N_24828,N_24459);
and U25027 (N_25027,N_24975,N_24723);
nor U25028 (N_25028,N_24670,N_24568);
nand U25029 (N_25029,N_24996,N_24185);
nand U25030 (N_25030,N_24542,N_24687);
xor U25031 (N_25031,N_24097,N_24544);
or U25032 (N_25032,N_24415,N_24634);
nor U25033 (N_25033,N_24127,N_24099);
and U25034 (N_25034,N_24921,N_24025);
and U25035 (N_25035,N_24661,N_24301);
nand U25036 (N_25036,N_24339,N_24038);
or U25037 (N_25037,N_24150,N_24787);
or U25038 (N_25038,N_24232,N_24803);
or U25039 (N_25039,N_24627,N_24247);
or U25040 (N_25040,N_24279,N_24469);
nand U25041 (N_25041,N_24405,N_24399);
nand U25042 (N_25042,N_24487,N_24700);
nor U25043 (N_25043,N_24628,N_24822);
or U25044 (N_25044,N_24995,N_24203);
xor U25045 (N_25045,N_24788,N_24411);
nor U25046 (N_25046,N_24579,N_24178);
or U25047 (N_25047,N_24576,N_24418);
and U25048 (N_25048,N_24052,N_24964);
and U25049 (N_25049,N_24972,N_24409);
xor U25050 (N_25050,N_24329,N_24011);
or U25051 (N_25051,N_24750,N_24444);
xor U25052 (N_25052,N_24230,N_24088);
or U25053 (N_25053,N_24983,N_24245);
nand U25054 (N_25054,N_24431,N_24560);
or U25055 (N_25055,N_24748,N_24004);
or U25056 (N_25056,N_24446,N_24977);
nand U25057 (N_25057,N_24059,N_24924);
and U25058 (N_25058,N_24327,N_24452);
or U25059 (N_25059,N_24804,N_24282);
xnor U25060 (N_25060,N_24266,N_24585);
and U25061 (N_25061,N_24352,N_24300);
nand U25062 (N_25062,N_24932,N_24380);
xor U25063 (N_25063,N_24154,N_24437);
or U25064 (N_25064,N_24033,N_24274);
nor U25065 (N_25065,N_24501,N_24985);
and U25066 (N_25066,N_24507,N_24265);
nand U25067 (N_25067,N_24143,N_24486);
and U25068 (N_25068,N_24246,N_24864);
and U25069 (N_25069,N_24846,N_24443);
xnor U25070 (N_25070,N_24597,N_24118);
nand U25071 (N_25071,N_24306,N_24591);
or U25072 (N_25072,N_24604,N_24824);
or U25073 (N_25073,N_24729,N_24070);
xor U25074 (N_25074,N_24673,N_24939);
nand U25075 (N_25075,N_24622,N_24567);
and U25076 (N_25076,N_24696,N_24947);
nor U25077 (N_25077,N_24035,N_24087);
or U25078 (N_25078,N_24945,N_24807);
nor U25079 (N_25079,N_24863,N_24659);
nor U25080 (N_25080,N_24007,N_24779);
xor U25081 (N_25081,N_24367,N_24345);
nor U25082 (N_25082,N_24191,N_24332);
nor U25083 (N_25083,N_24288,N_24258);
or U25084 (N_25084,N_24356,N_24278);
nor U25085 (N_25085,N_24705,N_24517);
nand U25086 (N_25086,N_24394,N_24626);
nand U25087 (N_25087,N_24090,N_24297);
and U25088 (N_25088,N_24630,N_24682);
nor U25089 (N_25089,N_24882,N_24021);
and U25090 (N_25090,N_24386,N_24902);
or U25091 (N_25091,N_24112,N_24897);
or U25092 (N_25092,N_24582,N_24349);
nand U25093 (N_25093,N_24130,N_24000);
xor U25094 (N_25094,N_24322,N_24264);
nor U25095 (N_25095,N_24753,N_24014);
and U25096 (N_25096,N_24868,N_24812);
nor U25097 (N_25097,N_24173,N_24132);
xor U25098 (N_25098,N_24208,N_24987);
nor U25099 (N_25099,N_24869,N_24302);
xor U25100 (N_25100,N_24862,N_24694);
xor U25101 (N_25101,N_24504,N_24768);
nor U25102 (N_25102,N_24385,N_24806);
nor U25103 (N_25103,N_24785,N_24119);
or U25104 (N_25104,N_24034,N_24006);
xnor U25105 (N_25105,N_24872,N_24162);
xor U25106 (N_25106,N_24666,N_24049);
nand U25107 (N_25107,N_24984,N_24686);
xnor U25108 (N_25108,N_24428,N_24857);
nand U25109 (N_25109,N_24888,N_24054);
xnor U25110 (N_25110,N_24390,N_24678);
nand U25111 (N_25111,N_24892,N_24314);
or U25112 (N_25112,N_24260,N_24135);
nand U25113 (N_25113,N_24993,N_24636);
xnor U25114 (N_25114,N_24740,N_24164);
and U25115 (N_25115,N_24715,N_24480);
or U25116 (N_25116,N_24430,N_24878);
and U25117 (N_25117,N_24967,N_24216);
or U25118 (N_25118,N_24741,N_24586);
and U25119 (N_25119,N_24778,N_24657);
nand U25120 (N_25120,N_24476,N_24434);
or U25121 (N_25121,N_24506,N_24810);
nor U25122 (N_25122,N_24138,N_24063);
nor U25123 (N_25123,N_24198,N_24581);
nand U25124 (N_25124,N_24369,N_24294);
and U25125 (N_25125,N_24974,N_24919);
xnor U25126 (N_25126,N_24599,N_24843);
and U25127 (N_25127,N_24588,N_24295);
nand U25128 (N_25128,N_24761,N_24354);
nor U25129 (N_25129,N_24166,N_24147);
and U25130 (N_25130,N_24584,N_24262);
xnor U25131 (N_25131,N_24609,N_24091);
nand U25132 (N_25132,N_24650,N_24551);
nor U25133 (N_25133,N_24889,N_24226);
nor U25134 (N_25134,N_24844,N_24722);
xor U25135 (N_25135,N_24898,N_24886);
xor U25136 (N_25136,N_24387,N_24089);
nor U25137 (N_25137,N_24826,N_24858);
nor U25138 (N_25138,N_24766,N_24194);
nor U25139 (N_25139,N_24739,N_24937);
nand U25140 (N_25140,N_24479,N_24496);
xnor U25141 (N_25141,N_24607,N_24860);
and U25142 (N_25142,N_24031,N_24180);
and U25143 (N_25143,N_24891,N_24057);
xnor U25144 (N_25144,N_24681,N_24441);
or U25145 (N_25145,N_24414,N_24601);
or U25146 (N_25146,N_24471,N_24851);
or U25147 (N_25147,N_24848,N_24978);
and U25148 (N_25148,N_24953,N_24429);
or U25149 (N_25149,N_24085,N_24662);
and U25150 (N_25150,N_24637,N_24001);
nand U25151 (N_25151,N_24474,N_24566);
xnor U25152 (N_25152,N_24684,N_24982);
or U25153 (N_25153,N_24814,N_24461);
or U25154 (N_25154,N_24378,N_24527);
nand U25155 (N_25155,N_24256,N_24493);
nand U25156 (N_25156,N_24157,N_24508);
or U25157 (N_25157,N_24689,N_24123);
and U25158 (N_25158,N_24095,N_24020);
nand U25159 (N_25159,N_24885,N_24899);
nor U25160 (N_25160,N_24611,N_24076);
or U25161 (N_25161,N_24065,N_24677);
xnor U25162 (N_25162,N_24159,N_24370);
xnor U25163 (N_25163,N_24991,N_24933);
and U25164 (N_25164,N_24227,N_24513);
nand U25165 (N_25165,N_24381,N_24234);
nor U25166 (N_25166,N_24916,N_24613);
nor U25167 (N_25167,N_24713,N_24570);
nor U25168 (N_25168,N_24742,N_24388);
or U25169 (N_25169,N_24797,N_24697);
nand U25170 (N_25170,N_24594,N_24350);
xor U25171 (N_25171,N_24629,N_24758);
nor U25172 (N_25172,N_24557,N_24619);
nand U25173 (N_25173,N_24160,N_24942);
xor U25174 (N_25174,N_24745,N_24072);
nor U25175 (N_25175,N_24532,N_24552);
nand U25176 (N_25176,N_24683,N_24638);
nor U25177 (N_25177,N_24169,N_24511);
xor U25178 (N_25178,N_24894,N_24961);
nor U25179 (N_25179,N_24419,N_24269);
xnor U25180 (N_25180,N_24207,N_24075);
nand U25181 (N_25181,N_24510,N_24577);
or U25182 (N_25182,N_24962,N_24820);
and U25183 (N_25183,N_24424,N_24308);
xnor U25184 (N_25184,N_24877,N_24680);
and U25185 (N_25185,N_24144,N_24061);
or U25186 (N_25186,N_24478,N_24482);
or U25187 (N_25187,N_24403,N_24545);
xnor U25188 (N_25188,N_24201,N_24530);
nand U25189 (N_25189,N_24698,N_24602);
or U25190 (N_25190,N_24703,N_24976);
xnor U25191 (N_25191,N_24850,N_24859);
nor U25192 (N_25192,N_24375,N_24731);
xor U25193 (N_25193,N_24037,N_24559);
xnor U25194 (N_25194,N_24058,N_24215);
nor U25195 (N_25195,N_24284,N_24024);
and U25196 (N_25196,N_24676,N_24764);
nor U25197 (N_25197,N_24829,N_24500);
and U25198 (N_25198,N_24562,N_24465);
nor U25199 (N_25199,N_24136,N_24161);
xor U25200 (N_25200,N_24518,N_24793);
nor U25201 (N_25201,N_24798,N_24954);
nor U25202 (N_25202,N_24184,N_24324);
nor U25203 (N_25203,N_24728,N_24299);
or U25204 (N_25204,N_24298,N_24464);
or U25205 (N_25205,N_24556,N_24019);
and U25206 (N_25206,N_24719,N_24635);
nand U25207 (N_25207,N_24176,N_24240);
and U25208 (N_25208,N_24372,N_24692);
or U25209 (N_25209,N_24121,N_24710);
nor U25210 (N_25210,N_24875,N_24809);
or U25211 (N_25211,N_24755,N_24935);
nand U25212 (N_25212,N_24359,N_24081);
nor U25213 (N_25213,N_24218,N_24834);
or U25214 (N_25214,N_24669,N_24268);
nand U25215 (N_25215,N_24426,N_24811);
nor U25216 (N_25216,N_24286,N_24319);
nand U25217 (N_25217,N_24861,N_24771);
nor U25218 (N_25218,N_24813,N_24502);
nor U25219 (N_25219,N_24881,N_24690);
or U25220 (N_25220,N_24098,N_24223);
or U25221 (N_25221,N_24272,N_24468);
and U25222 (N_25222,N_24654,N_24943);
nor U25223 (N_25223,N_24546,N_24784);
nand U25224 (N_25224,N_24366,N_24537);
and U25225 (N_25225,N_24447,N_24603);
xor U25226 (N_25226,N_24010,N_24027);
xnor U25227 (N_25227,N_24046,N_24941);
and U25228 (N_25228,N_24318,N_24336);
nand U25229 (N_25229,N_24221,N_24204);
xor U25230 (N_25230,N_24895,N_24343);
or U25231 (N_25231,N_24412,N_24104);
nand U25232 (N_25232,N_24311,N_24340);
nor U25233 (N_25233,N_24101,N_24817);
and U25234 (N_25234,N_24315,N_24571);
xor U25235 (N_25235,N_24190,N_24515);
or U25236 (N_25236,N_24016,N_24131);
or U25237 (N_25237,N_24514,N_24053);
nand U25238 (N_25238,N_24794,N_24397);
xnor U25239 (N_25239,N_24435,N_24254);
nor U25240 (N_25240,N_24664,N_24077);
nor U25241 (N_25241,N_24492,N_24534);
or U25242 (N_25242,N_24029,N_24225);
nand U25243 (N_25243,N_24477,N_24906);
xnor U25244 (N_25244,N_24392,N_24032);
nor U25245 (N_25245,N_24093,N_24606);
or U25246 (N_25246,N_24956,N_24107);
and U25247 (N_25247,N_24321,N_24263);
xnor U25248 (N_25248,N_24725,N_24940);
and U25249 (N_25249,N_24317,N_24472);
nand U25250 (N_25250,N_24575,N_24767);
xnor U25251 (N_25251,N_24790,N_24328);
nand U25252 (N_25252,N_24106,N_24280);
nand U25253 (N_25253,N_24128,N_24992);
and U25254 (N_25254,N_24523,N_24938);
and U25255 (N_25255,N_24422,N_24134);
xor U25256 (N_25256,N_24931,N_24873);
and U25257 (N_25257,N_24365,N_24854);
xnor U25258 (N_25258,N_24856,N_24003);
and U25259 (N_25259,N_24838,N_24013);
nor U25260 (N_25260,N_24199,N_24361);
or U25261 (N_25261,N_24749,N_24738);
nand U25262 (N_25262,N_24776,N_24918);
nor U25263 (N_25263,N_24578,N_24165);
nor U25264 (N_25264,N_24287,N_24957);
nor U25265 (N_25265,N_24711,N_24427);
or U25266 (N_25266,N_24467,N_24457);
nor U25267 (N_25267,N_24313,N_24228);
nor U25268 (N_25268,N_24695,N_24172);
and U25269 (N_25269,N_24540,N_24358);
nor U25270 (N_25270,N_24837,N_24909);
xnor U25271 (N_25271,N_24125,N_24901);
or U25272 (N_25272,N_24639,N_24531);
or U25273 (N_25273,N_24774,N_24520);
nand U25274 (N_25274,N_24398,N_24675);
and U25275 (N_25275,N_24734,N_24999);
or U25276 (N_25276,N_24847,N_24616);
nor U25277 (N_25277,N_24979,N_24655);
nor U25278 (N_25278,N_24293,N_24718);
or U25279 (N_25279,N_24799,N_24117);
and U25280 (N_25280,N_24368,N_24792);
nor U25281 (N_25281,N_24831,N_24382);
xor U25282 (N_25282,N_24870,N_24113);
nor U25283 (N_25283,N_24805,N_24632);
and U25284 (N_25284,N_24716,N_24535);
nor U25285 (N_25285,N_24200,N_24835);
xor U25286 (N_25286,N_24653,N_24538);
and U25287 (N_25287,N_24926,N_24440);
nand U25288 (N_25288,N_24927,N_24780);
xnor U25289 (N_25289,N_24801,N_24707);
xnor U25290 (N_25290,N_24094,N_24549);
xnor U25291 (N_25291,N_24241,N_24389);
nand U25292 (N_25292,N_24083,N_24533);
or U25293 (N_25293,N_24338,N_24874);
xnor U25294 (N_25294,N_24815,N_24115);
nor U25295 (N_25295,N_24516,N_24786);
nor U25296 (N_25296,N_24044,N_24015);
and U25297 (N_25297,N_24563,N_24808);
nor U25298 (N_25298,N_24600,N_24079);
xor U25299 (N_25299,N_24420,N_24842);
and U25300 (N_25300,N_24122,N_24141);
nor U25301 (N_25301,N_24770,N_24222);
nor U25302 (N_25302,N_24968,N_24383);
nand U25303 (N_25303,N_24830,N_24146);
and U25304 (N_25304,N_24782,N_24679);
or U25305 (N_25305,N_24402,N_24840);
and U25306 (N_25306,N_24866,N_24644);
and U25307 (N_25307,N_24617,N_24290);
nand U25308 (N_25308,N_24206,N_24944);
or U25309 (N_25309,N_24853,N_24911);
and U25310 (N_25310,N_24724,N_24971);
nand U25311 (N_25311,N_24432,N_24952);
nor U25312 (N_25312,N_24273,N_24255);
or U25313 (N_25313,N_24296,N_24645);
and U25314 (N_25314,N_24149,N_24913);
nor U25315 (N_25315,N_24752,N_24111);
nor U25316 (N_25316,N_24271,N_24548);
and U25317 (N_25317,N_24353,N_24565);
or U25318 (N_25318,N_24867,N_24555);
and U25319 (N_25319,N_24691,N_24499);
or U25320 (N_25320,N_24819,N_24163);
or U25321 (N_25321,N_24168,N_24849);
xor U25322 (N_25322,N_24701,N_24494);
nand U25323 (N_25323,N_24410,N_24489);
xnor U25324 (N_25324,N_24220,N_24789);
nor U25325 (N_25325,N_24827,N_24051);
and U25326 (N_25326,N_24553,N_24460);
nor U25327 (N_25327,N_24922,N_24102);
nand U25328 (N_25328,N_24539,N_24067);
and U25329 (N_25329,N_24948,N_24876);
and U25330 (N_25330,N_24374,N_24291);
nor U25331 (N_25331,N_24005,N_24259);
nor U25332 (N_25332,N_24760,N_24481);
nand U25333 (N_25333,N_24592,N_24903);
xor U25334 (N_25334,N_24047,N_24746);
nand U25335 (N_25335,N_24304,N_24525);
and U25336 (N_25336,N_24528,N_24074);
nand U25337 (N_25337,N_24685,N_24002);
nand U25338 (N_25338,N_24043,N_24915);
xnor U25339 (N_25339,N_24416,N_24448);
nand U25340 (N_25340,N_24012,N_24949);
xor U25341 (N_25341,N_24073,N_24442);
or U25342 (N_25342,N_24145,N_24572);
nand U25343 (N_25343,N_24341,N_24022);
xnor U25344 (N_25344,N_24702,N_24139);
or U25345 (N_25345,N_24244,N_24276);
xnor U25346 (N_25346,N_24028,N_24116);
xor U25347 (N_25347,N_24156,N_24114);
nor U25348 (N_25348,N_24646,N_24777);
xor U25349 (N_25349,N_24721,N_24323);
and U25350 (N_25350,N_24800,N_24688);
nand U25351 (N_25351,N_24217,N_24036);
or U25352 (N_25352,N_24108,N_24351);
and U25353 (N_25353,N_24773,N_24129);
and U25354 (N_25354,N_24498,N_24699);
or U25355 (N_25355,N_24400,N_24998);
or U25356 (N_25356,N_24231,N_24148);
xor U25357 (N_25357,N_24708,N_24084);
xnor U25358 (N_25358,N_24404,N_24363);
and U25359 (N_25359,N_24064,N_24212);
xnor U25360 (N_25360,N_24307,N_24583);
and U25361 (N_25361,N_24717,N_24456);
nor U25362 (N_25362,N_24865,N_24393);
and U25363 (N_25363,N_24712,N_24473);
or U25364 (N_25364,N_24214,N_24633);
nor U25365 (N_25365,N_24377,N_24623);
xnor U25366 (N_25366,N_24153,N_24665);
or U25367 (N_25367,N_24485,N_24455);
and U25368 (N_25368,N_24598,N_24330);
or U25369 (N_25369,N_24973,N_24237);
and U25370 (N_25370,N_24171,N_24610);
and U25371 (N_25371,N_24934,N_24466);
nor U25372 (N_25372,N_24086,N_24648);
and U25373 (N_25373,N_24188,N_24615);
xor U25374 (N_25374,N_24709,N_24009);
and U25375 (N_25375,N_24396,N_24096);
and U25376 (N_25376,N_24069,N_24706);
or U25377 (N_25377,N_24197,N_24522);
nor U25378 (N_25378,N_24986,N_24026);
or U25379 (N_25379,N_24614,N_24519);
nand U25380 (N_25380,N_24334,N_24543);
and U25381 (N_25381,N_24417,N_24316);
and U25382 (N_25382,N_24100,N_24852);
and U25383 (N_25383,N_24320,N_24693);
nand U25384 (N_25384,N_24331,N_24371);
xnor U25385 (N_25385,N_24747,N_24018);
and U25386 (N_25386,N_24988,N_24726);
and U25387 (N_25387,N_24192,N_24561);
and U25388 (N_25388,N_24620,N_24174);
xor U25389 (N_25389,N_24347,N_24235);
nor U25390 (N_25390,N_24433,N_24050);
or U25391 (N_25391,N_24994,N_24621);
and U25392 (N_25392,N_24841,N_24960);
nor U25393 (N_25393,N_24651,N_24816);
or U25394 (N_25394,N_24855,N_24105);
and U25395 (N_25395,N_24066,N_24152);
nor U25396 (N_25396,N_24364,N_24503);
and U25397 (N_25397,N_24137,N_24912);
or U25398 (N_25398,N_24720,N_24080);
and U25399 (N_25399,N_24625,N_24714);
nor U25400 (N_25400,N_24509,N_24925);
nor U25401 (N_25401,N_24346,N_24550);
or U25402 (N_25402,N_24641,N_24140);
and U25403 (N_25403,N_24521,N_24242);
xnor U25404 (N_25404,N_24928,N_24495);
or U25405 (N_25405,N_24187,N_24605);
nor U25406 (N_25406,N_24177,N_24608);
nand U25407 (N_25407,N_24757,N_24936);
nor U25408 (N_25408,N_24959,N_24783);
nor U25409 (N_25409,N_24483,N_24071);
nor U25410 (N_25410,N_24905,N_24769);
nor U25411 (N_25411,N_24008,N_24167);
and U25412 (N_25412,N_24762,N_24823);
nor U25413 (N_25413,N_24155,N_24275);
and U25414 (N_25414,N_24175,N_24395);
and U25415 (N_25415,N_24186,N_24997);
or U25416 (N_25416,N_24946,N_24505);
and U25417 (N_25417,N_24039,N_24951);
and U25418 (N_25418,N_24672,N_24082);
nor U25419 (N_25419,N_24484,N_24253);
or U25420 (N_25420,N_24249,N_24989);
xor U25421 (N_25421,N_24871,N_24836);
nor U25422 (N_25422,N_24355,N_24023);
or U25423 (N_25423,N_24536,N_24454);
or U25424 (N_25424,N_24423,N_24379);
or U25425 (N_25425,N_24056,N_24236);
nand U25426 (N_25426,N_24907,N_24103);
and U25427 (N_25427,N_24373,N_24595);
xnor U25428 (N_25428,N_24289,N_24730);
nor U25429 (N_25429,N_24158,N_24183);
and U25430 (N_25430,N_24966,N_24775);
nand U25431 (N_25431,N_24257,N_24252);
nand U25432 (N_25432,N_24283,N_24671);
xnor U25433 (N_25433,N_24055,N_24238);
and U25434 (N_25434,N_24763,N_24391);
xnor U25435 (N_25435,N_24309,N_24333);
xnor U25436 (N_25436,N_24305,N_24893);
nor U25437 (N_25437,N_24587,N_24401);
nor U25438 (N_25438,N_24950,N_24884);
or U25439 (N_25439,N_24908,N_24407);
or U25440 (N_25440,N_24660,N_24890);
or U25441 (N_25441,N_24825,N_24754);
and U25442 (N_25442,N_24202,N_24596);
nor U25443 (N_25443,N_24413,N_24791);
xor U25444 (N_25444,N_24980,N_24270);
nand U25445 (N_25445,N_24142,N_24438);
or U25446 (N_25446,N_24406,N_24470);
or U25447 (N_25447,N_24737,N_24573);
and U25448 (N_25448,N_24110,N_24362);
nor U25449 (N_25449,N_24041,N_24042);
and U25450 (N_25450,N_24219,N_24541);
or U25451 (N_25451,N_24120,N_24569);
nor U25452 (N_25452,N_24990,N_24335);
nor U25453 (N_25453,N_24554,N_24450);
or U25454 (N_25454,N_24904,N_24642);
nor U25455 (N_25455,N_24781,N_24920);
nor U25456 (N_25456,N_24462,N_24929);
and U25457 (N_25457,N_24344,N_24408);
xor U25458 (N_25458,N_24732,N_24436);
nand U25459 (N_25459,N_24832,N_24795);
nor U25460 (N_25460,N_24109,N_24181);
xnor U25461 (N_25461,N_24580,N_24342);
or U25462 (N_25462,N_24751,N_24292);
nand U25463 (N_25463,N_24179,N_24453);
nor U25464 (N_25464,N_24193,N_24736);
nand U25465 (N_25465,N_24647,N_24845);
and U25466 (N_25466,N_24078,N_24243);
xor U25467 (N_25467,N_24189,N_24574);
nor U25468 (N_25468,N_24524,N_24656);
nor U25469 (N_25469,N_24151,N_24743);
nand U25470 (N_25470,N_24735,N_24910);
and U25471 (N_25471,N_24182,N_24618);
and U25472 (N_25472,N_24589,N_24211);
nor U25473 (N_25473,N_24312,N_24030);
or U25474 (N_25474,N_24704,N_24229);
nand U25475 (N_25475,N_24879,N_24727);
nor U25476 (N_25476,N_24970,N_24963);
nand U25477 (N_25477,N_24839,N_24674);
or U25478 (N_25478,N_24512,N_24475);
nor U25479 (N_25479,N_24209,N_24451);
nand U25480 (N_25480,N_24756,N_24497);
xnor U25481 (N_25481,N_24281,N_24239);
xnor U25482 (N_25482,N_24040,N_24917);
and U25483 (N_25483,N_24744,N_24958);
or U25484 (N_25484,N_24965,N_24668);
nand U25485 (N_25485,N_24772,N_24045);
xor U25486 (N_25486,N_24802,N_24900);
and U25487 (N_25487,N_24325,N_24612);
and U25488 (N_25488,N_24818,N_24017);
and U25489 (N_25489,N_24310,N_24285);
and U25490 (N_25490,N_24458,N_24624);
nand U25491 (N_25491,N_24213,N_24558);
and U25492 (N_25492,N_24210,N_24663);
and U25493 (N_25493,N_24643,N_24267);
nand U25494 (N_25494,N_24133,N_24261);
or U25495 (N_25495,N_24250,N_24969);
nor U25496 (N_25496,N_24195,N_24914);
or U25497 (N_25497,N_24593,N_24421);
or U25498 (N_25498,N_24439,N_24923);
xnor U25499 (N_25499,N_24491,N_24326);
and U25500 (N_25500,N_24725,N_24566);
nor U25501 (N_25501,N_24017,N_24507);
and U25502 (N_25502,N_24706,N_24123);
nor U25503 (N_25503,N_24759,N_24725);
xor U25504 (N_25504,N_24325,N_24624);
nor U25505 (N_25505,N_24273,N_24298);
and U25506 (N_25506,N_24576,N_24855);
nor U25507 (N_25507,N_24356,N_24434);
nor U25508 (N_25508,N_24961,N_24757);
or U25509 (N_25509,N_24466,N_24196);
nor U25510 (N_25510,N_24629,N_24387);
and U25511 (N_25511,N_24514,N_24087);
nor U25512 (N_25512,N_24146,N_24753);
nor U25513 (N_25513,N_24657,N_24224);
nand U25514 (N_25514,N_24385,N_24783);
nand U25515 (N_25515,N_24523,N_24007);
and U25516 (N_25516,N_24442,N_24789);
xor U25517 (N_25517,N_24723,N_24716);
nor U25518 (N_25518,N_24484,N_24810);
nand U25519 (N_25519,N_24421,N_24170);
xor U25520 (N_25520,N_24751,N_24518);
nand U25521 (N_25521,N_24284,N_24115);
or U25522 (N_25522,N_24432,N_24946);
nand U25523 (N_25523,N_24140,N_24735);
or U25524 (N_25524,N_24897,N_24750);
xor U25525 (N_25525,N_24166,N_24566);
nor U25526 (N_25526,N_24859,N_24037);
and U25527 (N_25527,N_24431,N_24706);
and U25528 (N_25528,N_24797,N_24492);
nor U25529 (N_25529,N_24260,N_24428);
xnor U25530 (N_25530,N_24660,N_24816);
nand U25531 (N_25531,N_24191,N_24892);
or U25532 (N_25532,N_24824,N_24246);
xor U25533 (N_25533,N_24908,N_24477);
or U25534 (N_25534,N_24350,N_24081);
xor U25535 (N_25535,N_24614,N_24997);
or U25536 (N_25536,N_24823,N_24736);
xnor U25537 (N_25537,N_24759,N_24410);
and U25538 (N_25538,N_24966,N_24926);
nor U25539 (N_25539,N_24917,N_24604);
xor U25540 (N_25540,N_24186,N_24276);
or U25541 (N_25541,N_24483,N_24145);
nor U25542 (N_25542,N_24026,N_24388);
xor U25543 (N_25543,N_24957,N_24779);
or U25544 (N_25544,N_24229,N_24749);
xor U25545 (N_25545,N_24252,N_24992);
nor U25546 (N_25546,N_24299,N_24328);
or U25547 (N_25547,N_24020,N_24272);
and U25548 (N_25548,N_24003,N_24929);
and U25549 (N_25549,N_24297,N_24859);
xnor U25550 (N_25550,N_24316,N_24155);
nor U25551 (N_25551,N_24176,N_24867);
or U25552 (N_25552,N_24753,N_24988);
nand U25553 (N_25553,N_24344,N_24359);
or U25554 (N_25554,N_24469,N_24972);
and U25555 (N_25555,N_24414,N_24599);
nor U25556 (N_25556,N_24583,N_24763);
nand U25557 (N_25557,N_24178,N_24080);
nor U25558 (N_25558,N_24706,N_24170);
xnor U25559 (N_25559,N_24408,N_24202);
or U25560 (N_25560,N_24243,N_24051);
xor U25561 (N_25561,N_24480,N_24193);
nand U25562 (N_25562,N_24046,N_24025);
or U25563 (N_25563,N_24533,N_24215);
or U25564 (N_25564,N_24895,N_24577);
and U25565 (N_25565,N_24651,N_24877);
and U25566 (N_25566,N_24790,N_24882);
and U25567 (N_25567,N_24198,N_24732);
and U25568 (N_25568,N_24577,N_24556);
xnor U25569 (N_25569,N_24121,N_24275);
and U25570 (N_25570,N_24255,N_24220);
nor U25571 (N_25571,N_24181,N_24871);
nor U25572 (N_25572,N_24383,N_24149);
or U25573 (N_25573,N_24831,N_24447);
or U25574 (N_25574,N_24218,N_24112);
and U25575 (N_25575,N_24789,N_24430);
nand U25576 (N_25576,N_24533,N_24980);
nand U25577 (N_25577,N_24812,N_24215);
nand U25578 (N_25578,N_24068,N_24314);
nand U25579 (N_25579,N_24374,N_24966);
or U25580 (N_25580,N_24069,N_24780);
nand U25581 (N_25581,N_24027,N_24389);
or U25582 (N_25582,N_24563,N_24959);
xor U25583 (N_25583,N_24906,N_24099);
nor U25584 (N_25584,N_24507,N_24988);
and U25585 (N_25585,N_24403,N_24247);
or U25586 (N_25586,N_24762,N_24447);
nor U25587 (N_25587,N_24031,N_24330);
nand U25588 (N_25588,N_24324,N_24977);
and U25589 (N_25589,N_24020,N_24321);
and U25590 (N_25590,N_24226,N_24117);
nand U25591 (N_25591,N_24495,N_24876);
or U25592 (N_25592,N_24606,N_24460);
xor U25593 (N_25593,N_24139,N_24418);
nor U25594 (N_25594,N_24463,N_24780);
nand U25595 (N_25595,N_24689,N_24910);
nand U25596 (N_25596,N_24273,N_24033);
nor U25597 (N_25597,N_24661,N_24171);
nand U25598 (N_25598,N_24536,N_24505);
xor U25599 (N_25599,N_24646,N_24897);
and U25600 (N_25600,N_24512,N_24853);
nor U25601 (N_25601,N_24651,N_24216);
xnor U25602 (N_25602,N_24004,N_24087);
nor U25603 (N_25603,N_24156,N_24621);
or U25604 (N_25604,N_24514,N_24828);
nand U25605 (N_25605,N_24091,N_24508);
nand U25606 (N_25606,N_24162,N_24964);
xor U25607 (N_25607,N_24599,N_24098);
and U25608 (N_25608,N_24044,N_24031);
nand U25609 (N_25609,N_24097,N_24055);
xor U25610 (N_25610,N_24143,N_24757);
and U25611 (N_25611,N_24954,N_24659);
or U25612 (N_25612,N_24761,N_24614);
nor U25613 (N_25613,N_24656,N_24438);
nor U25614 (N_25614,N_24535,N_24359);
and U25615 (N_25615,N_24950,N_24141);
nor U25616 (N_25616,N_24272,N_24119);
and U25617 (N_25617,N_24581,N_24995);
nor U25618 (N_25618,N_24864,N_24321);
and U25619 (N_25619,N_24099,N_24155);
nor U25620 (N_25620,N_24581,N_24659);
nand U25621 (N_25621,N_24054,N_24448);
xor U25622 (N_25622,N_24595,N_24344);
xor U25623 (N_25623,N_24528,N_24050);
nand U25624 (N_25624,N_24243,N_24368);
nand U25625 (N_25625,N_24061,N_24704);
nand U25626 (N_25626,N_24772,N_24228);
nor U25627 (N_25627,N_24954,N_24519);
nor U25628 (N_25628,N_24152,N_24249);
and U25629 (N_25629,N_24545,N_24184);
nor U25630 (N_25630,N_24941,N_24495);
and U25631 (N_25631,N_24163,N_24456);
nor U25632 (N_25632,N_24695,N_24959);
and U25633 (N_25633,N_24461,N_24584);
xor U25634 (N_25634,N_24895,N_24684);
nand U25635 (N_25635,N_24005,N_24777);
and U25636 (N_25636,N_24255,N_24452);
or U25637 (N_25637,N_24625,N_24388);
nor U25638 (N_25638,N_24988,N_24011);
nor U25639 (N_25639,N_24646,N_24756);
nor U25640 (N_25640,N_24018,N_24394);
nand U25641 (N_25641,N_24315,N_24738);
xor U25642 (N_25642,N_24457,N_24031);
and U25643 (N_25643,N_24260,N_24015);
nor U25644 (N_25644,N_24886,N_24601);
or U25645 (N_25645,N_24351,N_24243);
nand U25646 (N_25646,N_24707,N_24511);
or U25647 (N_25647,N_24955,N_24246);
nor U25648 (N_25648,N_24477,N_24423);
nand U25649 (N_25649,N_24309,N_24219);
xnor U25650 (N_25650,N_24398,N_24150);
or U25651 (N_25651,N_24820,N_24501);
xnor U25652 (N_25652,N_24081,N_24113);
nor U25653 (N_25653,N_24025,N_24677);
or U25654 (N_25654,N_24636,N_24771);
xnor U25655 (N_25655,N_24109,N_24549);
or U25656 (N_25656,N_24660,N_24447);
and U25657 (N_25657,N_24293,N_24602);
nand U25658 (N_25658,N_24952,N_24225);
nor U25659 (N_25659,N_24915,N_24189);
and U25660 (N_25660,N_24808,N_24656);
xor U25661 (N_25661,N_24630,N_24920);
and U25662 (N_25662,N_24506,N_24755);
nand U25663 (N_25663,N_24360,N_24838);
xor U25664 (N_25664,N_24003,N_24426);
or U25665 (N_25665,N_24649,N_24831);
or U25666 (N_25666,N_24249,N_24100);
and U25667 (N_25667,N_24823,N_24019);
nand U25668 (N_25668,N_24765,N_24951);
nand U25669 (N_25669,N_24264,N_24879);
or U25670 (N_25670,N_24291,N_24106);
xnor U25671 (N_25671,N_24789,N_24419);
xnor U25672 (N_25672,N_24834,N_24247);
xor U25673 (N_25673,N_24221,N_24972);
and U25674 (N_25674,N_24303,N_24329);
nor U25675 (N_25675,N_24963,N_24959);
or U25676 (N_25676,N_24747,N_24137);
nor U25677 (N_25677,N_24107,N_24590);
nor U25678 (N_25678,N_24388,N_24805);
xnor U25679 (N_25679,N_24941,N_24031);
nor U25680 (N_25680,N_24321,N_24572);
or U25681 (N_25681,N_24141,N_24217);
xnor U25682 (N_25682,N_24994,N_24990);
xnor U25683 (N_25683,N_24746,N_24647);
nor U25684 (N_25684,N_24751,N_24177);
or U25685 (N_25685,N_24111,N_24997);
or U25686 (N_25686,N_24396,N_24172);
nand U25687 (N_25687,N_24503,N_24387);
or U25688 (N_25688,N_24679,N_24577);
nor U25689 (N_25689,N_24104,N_24890);
nand U25690 (N_25690,N_24298,N_24857);
nand U25691 (N_25691,N_24809,N_24149);
nand U25692 (N_25692,N_24893,N_24656);
xnor U25693 (N_25693,N_24138,N_24110);
or U25694 (N_25694,N_24767,N_24990);
nor U25695 (N_25695,N_24355,N_24300);
nand U25696 (N_25696,N_24389,N_24227);
nor U25697 (N_25697,N_24832,N_24803);
nand U25698 (N_25698,N_24285,N_24494);
nand U25699 (N_25699,N_24012,N_24120);
and U25700 (N_25700,N_24086,N_24982);
and U25701 (N_25701,N_24419,N_24394);
and U25702 (N_25702,N_24343,N_24419);
or U25703 (N_25703,N_24779,N_24072);
and U25704 (N_25704,N_24805,N_24748);
nand U25705 (N_25705,N_24224,N_24982);
xor U25706 (N_25706,N_24625,N_24713);
and U25707 (N_25707,N_24737,N_24151);
or U25708 (N_25708,N_24921,N_24980);
xor U25709 (N_25709,N_24748,N_24857);
nor U25710 (N_25710,N_24244,N_24094);
nor U25711 (N_25711,N_24548,N_24183);
or U25712 (N_25712,N_24023,N_24225);
xor U25713 (N_25713,N_24625,N_24547);
nand U25714 (N_25714,N_24650,N_24754);
and U25715 (N_25715,N_24747,N_24314);
nand U25716 (N_25716,N_24608,N_24930);
xor U25717 (N_25717,N_24412,N_24001);
nor U25718 (N_25718,N_24397,N_24953);
xnor U25719 (N_25719,N_24664,N_24244);
and U25720 (N_25720,N_24599,N_24045);
and U25721 (N_25721,N_24665,N_24819);
nand U25722 (N_25722,N_24966,N_24948);
nor U25723 (N_25723,N_24649,N_24800);
or U25724 (N_25724,N_24646,N_24058);
or U25725 (N_25725,N_24143,N_24037);
nand U25726 (N_25726,N_24684,N_24957);
and U25727 (N_25727,N_24137,N_24088);
xnor U25728 (N_25728,N_24017,N_24143);
and U25729 (N_25729,N_24239,N_24426);
xor U25730 (N_25730,N_24019,N_24127);
xnor U25731 (N_25731,N_24546,N_24371);
or U25732 (N_25732,N_24394,N_24483);
and U25733 (N_25733,N_24412,N_24786);
nor U25734 (N_25734,N_24317,N_24715);
nor U25735 (N_25735,N_24466,N_24951);
or U25736 (N_25736,N_24055,N_24481);
and U25737 (N_25737,N_24796,N_24076);
or U25738 (N_25738,N_24635,N_24497);
nand U25739 (N_25739,N_24060,N_24902);
or U25740 (N_25740,N_24847,N_24208);
xnor U25741 (N_25741,N_24947,N_24779);
nor U25742 (N_25742,N_24259,N_24534);
xnor U25743 (N_25743,N_24263,N_24958);
nor U25744 (N_25744,N_24824,N_24170);
and U25745 (N_25745,N_24293,N_24305);
xor U25746 (N_25746,N_24062,N_24618);
nor U25747 (N_25747,N_24500,N_24325);
or U25748 (N_25748,N_24690,N_24971);
or U25749 (N_25749,N_24340,N_24072);
nor U25750 (N_25750,N_24768,N_24235);
nor U25751 (N_25751,N_24190,N_24167);
nor U25752 (N_25752,N_24701,N_24474);
xor U25753 (N_25753,N_24465,N_24077);
nand U25754 (N_25754,N_24952,N_24692);
nand U25755 (N_25755,N_24257,N_24185);
nor U25756 (N_25756,N_24512,N_24193);
xor U25757 (N_25757,N_24593,N_24460);
nand U25758 (N_25758,N_24356,N_24471);
nand U25759 (N_25759,N_24652,N_24675);
or U25760 (N_25760,N_24814,N_24382);
nand U25761 (N_25761,N_24451,N_24091);
xor U25762 (N_25762,N_24180,N_24958);
nand U25763 (N_25763,N_24171,N_24076);
nand U25764 (N_25764,N_24663,N_24274);
nand U25765 (N_25765,N_24407,N_24012);
nor U25766 (N_25766,N_24599,N_24219);
nand U25767 (N_25767,N_24577,N_24730);
or U25768 (N_25768,N_24940,N_24572);
nand U25769 (N_25769,N_24541,N_24809);
xor U25770 (N_25770,N_24655,N_24225);
xnor U25771 (N_25771,N_24410,N_24691);
xnor U25772 (N_25772,N_24081,N_24859);
xnor U25773 (N_25773,N_24673,N_24972);
xor U25774 (N_25774,N_24192,N_24515);
and U25775 (N_25775,N_24636,N_24793);
nand U25776 (N_25776,N_24566,N_24927);
and U25777 (N_25777,N_24000,N_24244);
nand U25778 (N_25778,N_24173,N_24588);
and U25779 (N_25779,N_24855,N_24528);
nor U25780 (N_25780,N_24193,N_24300);
xnor U25781 (N_25781,N_24703,N_24661);
nand U25782 (N_25782,N_24093,N_24652);
nand U25783 (N_25783,N_24916,N_24349);
nand U25784 (N_25784,N_24065,N_24093);
nor U25785 (N_25785,N_24917,N_24406);
or U25786 (N_25786,N_24159,N_24880);
nand U25787 (N_25787,N_24528,N_24220);
xnor U25788 (N_25788,N_24066,N_24021);
xor U25789 (N_25789,N_24388,N_24648);
and U25790 (N_25790,N_24758,N_24389);
or U25791 (N_25791,N_24691,N_24389);
or U25792 (N_25792,N_24161,N_24292);
or U25793 (N_25793,N_24972,N_24750);
and U25794 (N_25794,N_24029,N_24875);
xnor U25795 (N_25795,N_24627,N_24259);
and U25796 (N_25796,N_24805,N_24064);
and U25797 (N_25797,N_24665,N_24449);
nand U25798 (N_25798,N_24565,N_24823);
and U25799 (N_25799,N_24472,N_24587);
and U25800 (N_25800,N_24873,N_24704);
nand U25801 (N_25801,N_24395,N_24598);
or U25802 (N_25802,N_24615,N_24057);
nor U25803 (N_25803,N_24259,N_24545);
nor U25804 (N_25804,N_24785,N_24231);
xnor U25805 (N_25805,N_24778,N_24503);
or U25806 (N_25806,N_24662,N_24945);
xor U25807 (N_25807,N_24056,N_24123);
xnor U25808 (N_25808,N_24327,N_24583);
xor U25809 (N_25809,N_24979,N_24827);
and U25810 (N_25810,N_24285,N_24323);
nand U25811 (N_25811,N_24840,N_24943);
and U25812 (N_25812,N_24419,N_24778);
and U25813 (N_25813,N_24753,N_24339);
nand U25814 (N_25814,N_24740,N_24360);
or U25815 (N_25815,N_24472,N_24259);
and U25816 (N_25816,N_24102,N_24852);
nand U25817 (N_25817,N_24565,N_24526);
or U25818 (N_25818,N_24666,N_24827);
xor U25819 (N_25819,N_24301,N_24259);
xnor U25820 (N_25820,N_24626,N_24431);
nand U25821 (N_25821,N_24686,N_24764);
and U25822 (N_25822,N_24081,N_24051);
and U25823 (N_25823,N_24515,N_24550);
and U25824 (N_25824,N_24934,N_24567);
nor U25825 (N_25825,N_24703,N_24825);
nor U25826 (N_25826,N_24083,N_24684);
nor U25827 (N_25827,N_24210,N_24597);
xor U25828 (N_25828,N_24450,N_24137);
or U25829 (N_25829,N_24631,N_24164);
xor U25830 (N_25830,N_24217,N_24703);
nor U25831 (N_25831,N_24736,N_24684);
nor U25832 (N_25832,N_24233,N_24554);
nand U25833 (N_25833,N_24989,N_24326);
xnor U25834 (N_25834,N_24298,N_24995);
xnor U25835 (N_25835,N_24697,N_24101);
or U25836 (N_25836,N_24043,N_24538);
and U25837 (N_25837,N_24893,N_24215);
nand U25838 (N_25838,N_24113,N_24290);
and U25839 (N_25839,N_24005,N_24126);
nand U25840 (N_25840,N_24580,N_24532);
nand U25841 (N_25841,N_24513,N_24188);
nand U25842 (N_25842,N_24521,N_24027);
and U25843 (N_25843,N_24677,N_24774);
or U25844 (N_25844,N_24000,N_24271);
or U25845 (N_25845,N_24150,N_24292);
or U25846 (N_25846,N_24603,N_24442);
and U25847 (N_25847,N_24602,N_24132);
and U25848 (N_25848,N_24692,N_24991);
xor U25849 (N_25849,N_24421,N_24416);
or U25850 (N_25850,N_24681,N_24732);
and U25851 (N_25851,N_24778,N_24972);
xnor U25852 (N_25852,N_24111,N_24306);
or U25853 (N_25853,N_24814,N_24363);
and U25854 (N_25854,N_24382,N_24966);
xor U25855 (N_25855,N_24992,N_24490);
and U25856 (N_25856,N_24380,N_24307);
nor U25857 (N_25857,N_24730,N_24551);
and U25858 (N_25858,N_24657,N_24713);
xor U25859 (N_25859,N_24901,N_24086);
or U25860 (N_25860,N_24980,N_24053);
and U25861 (N_25861,N_24408,N_24347);
nand U25862 (N_25862,N_24671,N_24017);
and U25863 (N_25863,N_24415,N_24867);
or U25864 (N_25864,N_24265,N_24610);
or U25865 (N_25865,N_24946,N_24837);
or U25866 (N_25866,N_24584,N_24739);
nand U25867 (N_25867,N_24292,N_24993);
xor U25868 (N_25868,N_24038,N_24803);
nand U25869 (N_25869,N_24914,N_24915);
xor U25870 (N_25870,N_24483,N_24084);
xnor U25871 (N_25871,N_24427,N_24371);
or U25872 (N_25872,N_24066,N_24633);
xor U25873 (N_25873,N_24383,N_24123);
nor U25874 (N_25874,N_24264,N_24248);
and U25875 (N_25875,N_24179,N_24029);
and U25876 (N_25876,N_24271,N_24813);
or U25877 (N_25877,N_24563,N_24007);
or U25878 (N_25878,N_24459,N_24953);
or U25879 (N_25879,N_24725,N_24169);
xor U25880 (N_25880,N_24511,N_24850);
xnor U25881 (N_25881,N_24969,N_24216);
nand U25882 (N_25882,N_24017,N_24834);
nand U25883 (N_25883,N_24503,N_24684);
nand U25884 (N_25884,N_24274,N_24676);
xnor U25885 (N_25885,N_24680,N_24872);
nand U25886 (N_25886,N_24240,N_24308);
xor U25887 (N_25887,N_24148,N_24625);
nor U25888 (N_25888,N_24594,N_24266);
nor U25889 (N_25889,N_24119,N_24871);
or U25890 (N_25890,N_24470,N_24041);
and U25891 (N_25891,N_24481,N_24510);
nand U25892 (N_25892,N_24469,N_24621);
xnor U25893 (N_25893,N_24024,N_24421);
xnor U25894 (N_25894,N_24222,N_24055);
nor U25895 (N_25895,N_24892,N_24845);
and U25896 (N_25896,N_24352,N_24961);
nor U25897 (N_25897,N_24796,N_24144);
xnor U25898 (N_25898,N_24319,N_24497);
and U25899 (N_25899,N_24799,N_24951);
xnor U25900 (N_25900,N_24117,N_24399);
nand U25901 (N_25901,N_24678,N_24973);
or U25902 (N_25902,N_24193,N_24822);
xnor U25903 (N_25903,N_24068,N_24872);
xnor U25904 (N_25904,N_24633,N_24935);
nand U25905 (N_25905,N_24757,N_24959);
nand U25906 (N_25906,N_24186,N_24425);
or U25907 (N_25907,N_24674,N_24696);
and U25908 (N_25908,N_24488,N_24790);
or U25909 (N_25909,N_24498,N_24957);
nand U25910 (N_25910,N_24223,N_24018);
nor U25911 (N_25911,N_24113,N_24185);
nor U25912 (N_25912,N_24529,N_24289);
and U25913 (N_25913,N_24940,N_24319);
or U25914 (N_25914,N_24812,N_24940);
xor U25915 (N_25915,N_24724,N_24524);
nor U25916 (N_25916,N_24622,N_24372);
xor U25917 (N_25917,N_24431,N_24477);
xor U25918 (N_25918,N_24208,N_24016);
xor U25919 (N_25919,N_24268,N_24803);
nand U25920 (N_25920,N_24217,N_24888);
xor U25921 (N_25921,N_24346,N_24730);
xnor U25922 (N_25922,N_24117,N_24541);
xnor U25923 (N_25923,N_24132,N_24036);
nand U25924 (N_25924,N_24979,N_24245);
xnor U25925 (N_25925,N_24482,N_24963);
and U25926 (N_25926,N_24493,N_24804);
xor U25927 (N_25927,N_24454,N_24748);
nor U25928 (N_25928,N_24176,N_24616);
and U25929 (N_25929,N_24720,N_24002);
nand U25930 (N_25930,N_24506,N_24376);
xor U25931 (N_25931,N_24196,N_24356);
and U25932 (N_25932,N_24013,N_24657);
nand U25933 (N_25933,N_24039,N_24591);
nor U25934 (N_25934,N_24410,N_24278);
nand U25935 (N_25935,N_24580,N_24095);
xnor U25936 (N_25936,N_24883,N_24473);
or U25937 (N_25937,N_24827,N_24324);
xor U25938 (N_25938,N_24146,N_24515);
nor U25939 (N_25939,N_24411,N_24387);
or U25940 (N_25940,N_24833,N_24969);
xor U25941 (N_25941,N_24198,N_24937);
xnor U25942 (N_25942,N_24676,N_24235);
and U25943 (N_25943,N_24330,N_24194);
nor U25944 (N_25944,N_24071,N_24601);
and U25945 (N_25945,N_24277,N_24029);
or U25946 (N_25946,N_24798,N_24586);
or U25947 (N_25947,N_24102,N_24754);
nor U25948 (N_25948,N_24965,N_24189);
nand U25949 (N_25949,N_24176,N_24774);
xor U25950 (N_25950,N_24409,N_24526);
nand U25951 (N_25951,N_24731,N_24144);
nor U25952 (N_25952,N_24668,N_24048);
and U25953 (N_25953,N_24578,N_24026);
nor U25954 (N_25954,N_24968,N_24770);
and U25955 (N_25955,N_24822,N_24518);
xnor U25956 (N_25956,N_24266,N_24331);
nand U25957 (N_25957,N_24396,N_24071);
and U25958 (N_25958,N_24836,N_24965);
and U25959 (N_25959,N_24243,N_24485);
and U25960 (N_25960,N_24154,N_24342);
and U25961 (N_25961,N_24422,N_24636);
nand U25962 (N_25962,N_24301,N_24694);
nor U25963 (N_25963,N_24560,N_24222);
nor U25964 (N_25964,N_24806,N_24267);
xnor U25965 (N_25965,N_24185,N_24343);
and U25966 (N_25966,N_24815,N_24357);
xnor U25967 (N_25967,N_24210,N_24201);
and U25968 (N_25968,N_24729,N_24921);
nor U25969 (N_25969,N_24424,N_24879);
nand U25970 (N_25970,N_24337,N_24786);
nand U25971 (N_25971,N_24062,N_24824);
and U25972 (N_25972,N_24275,N_24587);
nor U25973 (N_25973,N_24151,N_24920);
and U25974 (N_25974,N_24746,N_24664);
xor U25975 (N_25975,N_24401,N_24005);
and U25976 (N_25976,N_24963,N_24768);
nor U25977 (N_25977,N_24869,N_24235);
or U25978 (N_25978,N_24568,N_24831);
and U25979 (N_25979,N_24236,N_24405);
nor U25980 (N_25980,N_24715,N_24488);
nand U25981 (N_25981,N_24902,N_24919);
or U25982 (N_25982,N_24613,N_24689);
nand U25983 (N_25983,N_24202,N_24577);
or U25984 (N_25984,N_24740,N_24174);
and U25985 (N_25985,N_24289,N_24162);
or U25986 (N_25986,N_24977,N_24460);
xnor U25987 (N_25987,N_24815,N_24342);
nor U25988 (N_25988,N_24664,N_24966);
or U25989 (N_25989,N_24326,N_24819);
xor U25990 (N_25990,N_24854,N_24763);
nor U25991 (N_25991,N_24173,N_24457);
xor U25992 (N_25992,N_24926,N_24942);
nor U25993 (N_25993,N_24040,N_24178);
and U25994 (N_25994,N_24665,N_24077);
or U25995 (N_25995,N_24927,N_24487);
and U25996 (N_25996,N_24553,N_24707);
xnor U25997 (N_25997,N_24955,N_24037);
xor U25998 (N_25998,N_24291,N_24629);
or U25999 (N_25999,N_24463,N_24829);
xnor U26000 (N_26000,N_25302,N_25168);
and U26001 (N_26001,N_25234,N_25856);
nand U26002 (N_26002,N_25265,N_25324);
and U26003 (N_26003,N_25182,N_25347);
xnor U26004 (N_26004,N_25707,N_25206);
xor U26005 (N_26005,N_25314,N_25608);
and U26006 (N_26006,N_25586,N_25441);
nor U26007 (N_26007,N_25431,N_25526);
nand U26008 (N_26008,N_25826,N_25846);
nor U26009 (N_26009,N_25120,N_25413);
xnor U26010 (N_26010,N_25782,N_25658);
and U26011 (N_26011,N_25590,N_25629);
nand U26012 (N_26012,N_25521,N_25337);
or U26013 (N_26013,N_25944,N_25779);
nor U26014 (N_26014,N_25794,N_25358);
and U26015 (N_26015,N_25949,N_25591);
and U26016 (N_26016,N_25085,N_25260);
xor U26017 (N_26017,N_25614,N_25972);
and U26018 (N_26018,N_25718,N_25200);
nand U26019 (N_26019,N_25800,N_25738);
nand U26020 (N_26020,N_25542,N_25346);
nor U26021 (N_26021,N_25508,N_25982);
xnor U26022 (N_26022,N_25634,N_25790);
nand U26023 (N_26023,N_25583,N_25550);
xnor U26024 (N_26024,N_25137,N_25049);
nand U26025 (N_26025,N_25559,N_25050);
nand U26026 (N_26026,N_25239,N_25088);
xnor U26027 (N_26027,N_25113,N_25369);
nor U26028 (N_26028,N_25666,N_25620);
and U26029 (N_26029,N_25451,N_25763);
xor U26030 (N_26030,N_25303,N_25000);
and U26031 (N_26031,N_25587,N_25636);
and U26032 (N_26032,N_25652,N_25639);
nand U26033 (N_26033,N_25321,N_25627);
nand U26034 (N_26034,N_25423,N_25169);
nor U26035 (N_26035,N_25453,N_25041);
and U26036 (N_26036,N_25199,N_25281);
and U26037 (N_26037,N_25389,N_25716);
or U26038 (N_26038,N_25975,N_25861);
nand U26039 (N_26039,N_25044,N_25893);
nand U26040 (N_26040,N_25961,N_25227);
xor U26041 (N_26041,N_25219,N_25020);
nor U26042 (N_26042,N_25802,N_25991);
and U26043 (N_26043,N_25998,N_25354);
xnor U26044 (N_26044,N_25053,N_25187);
and U26045 (N_26045,N_25214,N_25514);
or U26046 (N_26046,N_25886,N_25726);
or U26047 (N_26047,N_25921,N_25771);
nand U26048 (N_26048,N_25569,N_25135);
nand U26049 (N_26049,N_25563,N_25709);
nor U26050 (N_26050,N_25173,N_25640);
nor U26051 (N_26051,N_25390,N_25503);
xor U26052 (N_26052,N_25820,N_25458);
nor U26053 (N_26053,N_25136,N_25552);
nand U26054 (N_26054,N_25320,N_25683);
xor U26055 (N_26055,N_25250,N_25381);
nand U26056 (N_26056,N_25638,N_25637);
nor U26057 (N_26057,N_25145,N_25106);
nand U26058 (N_26058,N_25190,N_25114);
or U26059 (N_26059,N_25895,N_25979);
or U26060 (N_26060,N_25238,N_25124);
nand U26061 (N_26061,N_25697,N_25950);
nand U26062 (N_26062,N_25947,N_25421);
nor U26063 (N_26063,N_25330,N_25153);
nand U26064 (N_26064,N_25076,N_25964);
and U26065 (N_26065,N_25525,N_25329);
nor U26066 (N_26066,N_25537,N_25372);
xnor U26067 (N_26067,N_25099,N_25804);
nand U26068 (N_26068,N_25243,N_25967);
and U26069 (N_26069,N_25512,N_25613);
nor U26070 (N_26070,N_25147,N_25313);
nand U26071 (N_26071,N_25648,N_25345);
nor U26072 (N_26072,N_25725,N_25942);
nand U26073 (N_26073,N_25660,N_25777);
or U26074 (N_26074,N_25203,N_25612);
nor U26075 (N_26075,N_25315,N_25167);
or U26076 (N_26076,N_25499,N_25673);
nor U26077 (N_26077,N_25202,N_25622);
nor U26078 (N_26078,N_25244,N_25016);
or U26079 (N_26079,N_25891,N_25761);
and U26080 (N_26080,N_25655,N_25813);
and U26081 (N_26081,N_25576,N_25862);
or U26082 (N_26082,N_25141,N_25412);
nand U26083 (N_26083,N_25457,N_25693);
or U26084 (N_26084,N_25486,N_25284);
or U26085 (N_26085,N_25491,N_25215);
nor U26086 (N_26086,N_25519,N_25603);
and U26087 (N_26087,N_25805,N_25970);
or U26088 (N_26088,N_25459,N_25161);
nand U26089 (N_26089,N_25222,N_25128);
and U26090 (N_26090,N_25722,N_25523);
and U26091 (N_26091,N_25040,N_25405);
and U26092 (N_26092,N_25830,N_25792);
nand U26093 (N_26093,N_25326,N_25208);
nor U26094 (N_26094,N_25401,N_25767);
and U26095 (N_26095,N_25857,N_25855);
and U26096 (N_26096,N_25954,N_25799);
nand U26097 (N_26097,N_25122,N_25117);
nand U26098 (N_26098,N_25992,N_25840);
nand U26099 (N_26099,N_25286,N_25064);
nor U26100 (N_26100,N_25680,N_25750);
xnor U26101 (N_26101,N_25473,N_25185);
and U26102 (N_26102,N_25816,N_25466);
nor U26103 (N_26103,N_25256,N_25657);
and U26104 (N_26104,N_25823,N_25295);
nor U26105 (N_26105,N_25894,N_25362);
and U26106 (N_26106,N_25151,N_25531);
or U26107 (N_26107,N_25294,N_25887);
nor U26108 (N_26108,N_25352,N_25920);
nor U26109 (N_26109,N_25659,N_25513);
or U26110 (N_26110,N_25356,N_25116);
nor U26111 (N_26111,N_25807,N_25892);
xor U26112 (N_26112,N_25661,N_25695);
nand U26113 (N_26113,N_25868,N_25649);
or U26114 (N_26114,N_25084,N_25916);
and U26115 (N_26115,N_25605,N_25086);
xor U26116 (N_26116,N_25713,N_25101);
nor U26117 (N_26117,N_25630,N_25134);
or U26118 (N_26118,N_25102,N_25353);
and U26119 (N_26119,N_25841,N_25357);
or U26120 (N_26120,N_25270,N_25382);
or U26121 (N_26121,N_25984,N_25487);
or U26122 (N_26122,N_25558,N_25070);
or U26123 (N_26123,N_25753,N_25910);
nor U26124 (N_26124,N_25398,N_25299);
or U26125 (N_26125,N_25279,N_25584);
xnor U26126 (N_26126,N_25186,N_25934);
nor U26127 (N_26127,N_25618,N_25765);
and U26128 (N_26128,N_25388,N_25046);
and U26129 (N_26129,N_25383,N_25948);
xnor U26130 (N_26130,N_25287,N_25480);
nor U26131 (N_26131,N_25937,N_25283);
and U26132 (N_26132,N_25791,N_25069);
nand U26133 (N_26133,N_25484,N_25737);
and U26134 (N_26134,N_25119,N_25348);
and U26135 (N_26135,N_25676,N_25269);
xnor U26136 (N_26136,N_25367,N_25465);
xor U26137 (N_26137,N_25783,N_25034);
xnor U26138 (N_26138,N_25776,N_25340);
nand U26139 (N_26139,N_25560,N_25987);
or U26140 (N_26140,N_25030,N_25908);
nor U26141 (N_26141,N_25770,N_25429);
and U26142 (N_26142,N_25156,N_25745);
or U26143 (N_26143,N_25434,N_25705);
xor U26144 (N_26144,N_25838,N_25643);
xor U26145 (N_26145,N_25043,N_25848);
nor U26146 (N_26146,N_25175,N_25217);
and U26147 (N_26147,N_25607,N_25042);
and U26148 (N_26148,N_25306,N_25006);
nand U26149 (N_26149,N_25926,N_25481);
nand U26150 (N_26150,N_25598,N_25715);
nor U26151 (N_26151,N_25110,N_25739);
nand U26152 (N_26152,N_25571,N_25031);
nor U26153 (N_26153,N_25176,N_25140);
xnor U26154 (N_26154,N_25670,N_25812);
nand U26155 (N_26155,N_25827,N_25965);
nor U26156 (N_26156,N_25485,N_25562);
nor U26157 (N_26157,N_25157,N_25392);
and U26158 (N_26158,N_25593,N_25181);
or U26159 (N_26159,N_25829,N_25786);
and U26160 (N_26160,N_25759,N_25701);
or U26161 (N_26161,N_25541,N_25801);
and U26162 (N_26162,N_25544,N_25863);
or U26163 (N_26163,N_25564,N_25714);
nand U26164 (N_26164,N_25496,N_25758);
nand U26165 (N_26165,N_25619,N_25518);
nor U26166 (N_26166,N_25506,N_25532);
nor U26167 (N_26167,N_25834,N_25743);
xnor U26168 (N_26168,N_25323,N_25416);
xor U26169 (N_26169,N_25430,N_25796);
or U26170 (N_26170,N_25883,N_25308);
nand U26171 (N_26171,N_25195,N_25821);
xnor U26172 (N_26172,N_25242,N_25539);
nor U26173 (N_26173,N_25907,N_25818);
nand U26174 (N_26174,N_25798,N_25094);
nor U26175 (N_26175,N_25579,N_25305);
and U26176 (N_26176,N_25602,N_25817);
and U26177 (N_26177,N_25507,N_25689);
and U26178 (N_26178,N_25054,N_25568);
and U26179 (N_26179,N_25549,N_25078);
nor U26180 (N_26180,N_25927,N_25842);
and U26181 (N_26181,N_25939,N_25455);
xnor U26182 (N_26182,N_25177,N_25278);
or U26183 (N_26183,N_25425,N_25896);
and U26184 (N_26184,N_25824,N_25261);
nand U26185 (N_26185,N_25056,N_25148);
and U26186 (N_26186,N_25428,N_25255);
xnor U26187 (N_26187,N_25932,N_25860);
and U26188 (N_26188,N_25492,N_25529);
xnor U26189 (N_26189,N_25803,N_25712);
xor U26190 (N_26190,N_25873,N_25240);
nor U26191 (N_26191,N_25669,N_25062);
nand U26192 (N_26192,N_25500,N_25462);
nand U26193 (N_26193,N_25922,N_25454);
xor U26194 (N_26194,N_25610,N_25015);
xnor U26195 (N_26195,N_25617,N_25788);
nor U26196 (N_26196,N_25588,N_25501);
nand U26197 (N_26197,N_25280,N_25448);
xor U26198 (N_26198,N_25444,N_25865);
and U26199 (N_26199,N_25684,N_25387);
nand U26200 (N_26200,N_25159,N_25557);
nor U26201 (N_26201,N_25505,N_25418);
nor U26202 (N_26202,N_25223,N_25565);
and U26203 (N_26203,N_25325,N_25131);
and U26204 (N_26204,N_25164,N_25033);
or U26205 (N_26205,N_25074,N_25734);
nor U26206 (N_26206,N_25960,N_25300);
or U26207 (N_26207,N_25682,N_25079);
or U26208 (N_26208,N_25625,N_25780);
nor U26209 (N_26209,N_25566,N_25904);
or U26210 (N_26210,N_25983,N_25595);
nand U26211 (N_26211,N_25751,N_25476);
nand U26212 (N_26212,N_25914,N_25230);
and U26213 (N_26213,N_25273,N_25993);
or U26214 (N_26214,N_25377,N_25599);
and U26215 (N_26215,N_25004,N_25847);
nor U26216 (N_26216,N_25130,N_25058);
nand U26217 (N_26217,N_25338,N_25720);
and U26218 (N_26218,N_25365,N_25008);
xnor U26219 (N_26219,N_25364,N_25439);
or U26220 (N_26220,N_25845,N_25748);
or U26221 (N_26221,N_25014,N_25172);
nand U26222 (N_26222,N_25692,N_25010);
xor U26223 (N_26223,N_25297,N_25740);
nand U26224 (N_26224,N_25342,N_25098);
and U26225 (N_26225,N_25427,N_25933);
nor U26226 (N_26226,N_25374,N_25528);
or U26227 (N_26227,N_25730,N_25092);
and U26228 (N_26228,N_25201,N_25930);
xnor U26229 (N_26229,N_25142,N_25757);
nor U26230 (N_26230,N_25391,N_25424);
xor U26231 (N_26231,N_25951,N_25045);
nand U26232 (N_26232,N_25262,N_25246);
and U26233 (N_26233,N_25048,N_25112);
xor U26234 (N_26234,N_25941,N_25154);
xor U26235 (N_26235,N_25095,N_25482);
and U26236 (N_26236,N_25121,N_25881);
or U26237 (N_26237,N_25809,N_25166);
nand U26238 (N_26238,N_25005,N_25925);
nand U26239 (N_26239,N_25903,N_25498);
nor U26240 (N_26240,N_25837,N_25968);
xnor U26241 (N_26241,N_25450,N_25547);
and U26242 (N_26242,N_25118,N_25978);
nor U26243 (N_26243,N_25533,N_25994);
nor U26244 (N_26244,N_25996,N_25601);
xnor U26245 (N_26245,N_25665,N_25061);
nor U26246 (N_26246,N_25415,N_25055);
nor U26247 (N_26247,N_25986,N_25104);
xnor U26248 (N_26248,N_25854,N_25778);
or U26249 (N_26249,N_25577,N_25899);
xor U26250 (N_26250,N_25072,N_25490);
nor U26251 (N_26251,N_25277,N_25567);
nand U26252 (N_26252,N_25806,N_25879);
and U26253 (N_26253,N_25875,N_25997);
or U26254 (N_26254,N_25966,N_25057);
nand U26255 (N_26255,N_25700,N_25024);
nand U26256 (N_26256,N_25653,N_25858);
xor U26257 (N_26257,N_25775,N_25795);
or U26258 (N_26258,N_25911,N_25958);
xnor U26259 (N_26259,N_25561,N_25125);
nand U26260 (N_26260,N_25859,N_25535);
xnor U26261 (N_26261,N_25366,N_25133);
and U26262 (N_26262,N_25822,N_25023);
xor U26263 (N_26263,N_25403,N_25237);
nand U26264 (N_26264,N_25645,N_25013);
or U26265 (N_26265,N_25733,N_25882);
nand U26266 (N_26266,N_25343,N_25442);
xor U26267 (N_26267,N_25332,N_25475);
nand U26268 (N_26268,N_25411,N_25218);
and U26269 (N_26269,N_25426,N_25530);
nor U26270 (N_26270,N_25677,N_25980);
or U26271 (N_26271,N_25864,N_25832);
or U26272 (N_26272,N_25467,N_25241);
and U26273 (N_26273,N_25754,N_25408);
or U26274 (N_26274,N_25756,N_25463);
nand U26275 (N_26275,N_25721,N_25436);
nor U26276 (N_26276,N_25589,N_25472);
nor U26277 (N_26277,N_25376,N_25524);
nor U26278 (N_26278,N_25548,N_25204);
xor U26279 (N_26279,N_25679,N_25762);
or U26280 (N_26280,N_25065,N_25257);
nand U26281 (N_26281,N_25249,N_25139);
nand U26282 (N_26282,N_25385,N_25878);
nand U26283 (N_26283,N_25409,N_25616);
or U26284 (N_26284,N_25963,N_25546);
nor U26285 (N_26285,N_25582,N_25611);
or U26286 (N_26286,N_25728,N_25035);
xor U26287 (N_26287,N_25650,N_25704);
nand U26288 (N_26288,N_25163,N_25211);
or U26289 (N_26289,N_25336,N_25681);
and U26290 (N_26290,N_25394,N_25909);
nand U26291 (N_26291,N_25808,N_25724);
nor U26292 (N_26292,N_25307,N_25331);
or U26293 (N_26293,N_25959,N_25969);
nand U26294 (N_26294,N_25929,N_25289);
nor U26295 (N_26295,N_25690,N_25288);
nand U26296 (N_26296,N_25397,N_25461);
and U26297 (N_26297,N_25171,N_25772);
nor U26298 (N_26298,N_25370,N_25404);
xnor U26299 (N_26299,N_25063,N_25090);
xnor U26300 (N_26300,N_25871,N_25727);
xor U26301 (N_26301,N_25268,N_25236);
nand U26302 (N_26302,N_25368,N_25474);
nand U26303 (N_26303,N_25912,N_25296);
and U26304 (N_26304,N_25876,N_25621);
and U26305 (N_26305,N_25310,N_25609);
xnor U26306 (N_26306,N_25594,N_25210);
nor U26307 (N_26307,N_25974,N_25170);
and U26308 (N_26308,N_25688,N_25538);
nor U26309 (N_26309,N_25380,N_25600);
xnor U26310 (N_26310,N_25874,N_25363);
and U26311 (N_26311,N_25971,N_25489);
nand U26312 (N_26312,N_25460,N_25654);
nand U26313 (N_26313,N_25276,N_25096);
nor U26314 (N_26314,N_25025,N_25890);
or U26315 (N_26315,N_25853,N_25851);
and U26316 (N_26316,N_25127,N_25059);
nand U26317 (N_26317,N_25263,N_25604);
or U26318 (N_26318,N_25953,N_25833);
and U26319 (N_26319,N_25843,N_25386);
nand U26320 (N_26320,N_25111,N_25849);
and U26321 (N_26321,N_25752,N_25527);
nor U26322 (N_26322,N_25723,N_25438);
xor U26323 (N_26323,N_25885,N_25815);
and U26324 (N_26324,N_25869,N_25844);
or U26325 (N_26325,N_25596,N_25956);
xnor U26326 (N_26326,N_25360,N_25011);
or U26327 (N_26327,N_25298,N_25735);
xor U26328 (N_26328,N_25995,N_25433);
nand U26329 (N_26329,N_25350,N_25898);
and U26330 (N_26330,N_25852,N_25764);
or U26331 (N_26331,N_25447,N_25511);
nor U26332 (N_26332,N_25836,N_25067);
xnor U26333 (N_26333,N_25144,N_25935);
nor U26334 (N_26334,N_25977,N_25395);
or U26335 (N_26335,N_25384,N_25641);
nand U26336 (N_26336,N_25819,N_25691);
nand U26337 (N_26337,N_25973,N_25018);
xnor U26338 (N_26338,N_25355,N_25212);
or U26339 (N_26339,N_25319,N_25685);
xnor U26340 (N_26340,N_25766,N_25445);
nand U26341 (N_26341,N_25393,N_25793);
and U26342 (N_26342,N_25251,N_25699);
nor U26343 (N_26343,N_25115,N_25706);
or U26344 (N_26344,N_25510,N_25509);
nor U26345 (N_26345,N_25469,N_25985);
nor U26346 (N_26346,N_25301,N_25174);
and U26347 (N_26347,N_25624,N_25719);
xnor U26348 (N_26348,N_25087,N_25220);
nand U26349 (N_26349,N_25696,N_25290);
xor U26350 (N_26350,N_25943,N_25708);
xnor U26351 (N_26351,N_25742,N_25183);
or U26352 (N_26352,N_25488,N_25870);
nor U26353 (N_26353,N_25334,N_25226);
nand U26354 (N_26354,N_25009,N_25642);
or U26355 (N_26355,N_25225,N_25703);
or U26356 (N_26356,N_25036,N_25651);
nor U26357 (N_26357,N_25271,N_25435);
or U26358 (N_26358,N_25002,N_25686);
xor U26359 (N_26359,N_25440,N_25597);
nand U26360 (N_26360,N_25952,N_25188);
xnor U26361 (N_26361,N_25781,N_25919);
or U26362 (N_26362,N_25573,N_25452);
xnor U26363 (N_26363,N_25258,N_25228);
and U26364 (N_26364,N_25417,N_25205);
nand U26365 (N_26365,N_25626,N_25520);
nand U26366 (N_26366,N_25769,N_25497);
nor U26367 (N_26367,N_25717,N_25917);
xor U26368 (N_26368,N_25275,N_25109);
nor U26369 (N_26369,N_25522,N_25027);
nand U26370 (N_26370,N_25628,N_25311);
nor U26371 (N_26371,N_25410,N_25437);
nand U26372 (N_26372,N_25536,N_25252);
and U26373 (N_26373,N_25318,N_25312);
xnor U26374 (N_26374,N_25349,N_25344);
nand U26375 (N_26375,N_25493,N_25126);
nand U26376 (N_26376,N_25768,N_25931);
or U26377 (N_26377,N_25534,N_25266);
or U26378 (N_26378,N_25747,N_25180);
nor U26379 (N_26379,N_25155,N_25731);
xor U26380 (N_26380,N_25516,N_25003);
xnor U26381 (N_26381,N_25913,N_25021);
and U26382 (N_26382,N_25254,N_25160);
xor U26383 (N_26383,N_25632,N_25149);
nand U26384 (N_26384,N_25736,N_25235);
xnor U26385 (N_26385,N_25464,N_25456);
nand U26386 (N_26386,N_25468,N_25902);
xnor U26387 (N_26387,N_25667,N_25988);
nand U26388 (N_26388,N_25662,N_25132);
or U26389 (N_26389,N_25581,N_25414);
nand U26390 (N_26390,N_25184,N_25773);
and U26391 (N_26391,N_25554,N_25068);
nand U26392 (N_26392,N_25196,N_25787);
and U26393 (N_26393,N_25378,N_25198);
and U26394 (N_26394,N_25880,N_25292);
nor U26395 (N_26395,N_25744,N_25687);
nor U26396 (N_26396,N_25647,N_25828);
or U26397 (N_26397,N_25471,N_25406);
or U26398 (N_26398,N_25189,N_25073);
or U26399 (N_26399,N_25553,N_25052);
or U26400 (N_26400,N_25515,N_25399);
or U26401 (N_26401,N_25047,N_25990);
nand U26402 (N_26402,N_25158,N_25322);
nand U26403 (N_26403,N_25019,N_25540);
nor U26404 (N_26404,N_25711,N_25123);
and U26405 (N_26405,N_25197,N_25253);
xor U26406 (N_26406,N_25760,N_25585);
and U26407 (N_26407,N_25267,N_25233);
and U26408 (N_26408,N_25867,N_25037);
and U26409 (N_26409,N_25075,N_25888);
nand U26410 (N_26410,N_25946,N_25359);
nor U26411 (N_26411,N_25749,N_25032);
and U26412 (N_26412,N_25671,N_25209);
nor U26413 (N_26413,N_25884,N_25291);
and U26414 (N_26414,N_25213,N_25100);
xnor U26415 (N_26415,N_25103,N_25606);
and U26416 (N_26416,N_25333,N_25162);
or U26417 (N_26417,N_25957,N_25915);
and U26418 (N_26418,N_25193,N_25897);
nand U26419 (N_26419,N_25082,N_25432);
and U26420 (N_26420,N_25179,N_25746);
xor U26421 (N_26421,N_25839,N_25517);
or U26422 (N_26422,N_25668,N_25029);
or U26423 (N_26423,N_25811,N_25989);
nand U26424 (N_26424,N_25039,N_25077);
nor U26425 (N_26425,N_25129,N_25945);
or U26426 (N_26426,N_25774,N_25631);
or U26427 (N_26427,N_25420,N_25923);
nor U26428 (N_26428,N_25729,N_25784);
nand U26429 (N_26429,N_25678,N_25351);
and U26430 (N_26430,N_25570,N_25495);
nor U26431 (N_26431,N_25051,N_25814);
or U26432 (N_26432,N_25664,N_25091);
nand U26433 (N_26433,N_25371,N_25245);
nor U26434 (N_26434,N_25316,N_25232);
nand U26435 (N_26435,N_25906,N_25191);
or U26436 (N_26436,N_25905,N_25282);
nor U26437 (N_26437,N_25248,N_25976);
xnor U26438 (N_26438,N_25001,N_25741);
and U26439 (N_26439,N_25810,N_25107);
nand U26440 (N_26440,N_25060,N_25419);
nand U26441 (N_26441,N_25089,N_25216);
or U26442 (N_26442,N_25327,N_25443);
xor U26443 (N_26443,N_25574,N_25702);
nor U26444 (N_26444,N_25850,N_25592);
or U26445 (N_26445,N_25635,N_25402);
or U26446 (N_26446,N_25375,N_25710);
and U26447 (N_26447,N_25012,N_25789);
and U26448 (N_26448,N_25304,N_25835);
nor U26449 (N_26449,N_25293,N_25272);
or U26450 (N_26450,N_25672,N_25083);
or U26451 (N_26451,N_25007,N_25962);
nand U26452 (N_26452,N_25097,N_25143);
or U26453 (N_26453,N_25502,N_25877);
xnor U26454 (N_26454,N_25422,N_25494);
xnor U26455 (N_26455,N_25361,N_25999);
nand U26456 (N_26456,N_25981,N_25247);
and U26457 (N_26457,N_25825,N_25274);
nand U26458 (N_26458,N_25889,N_25938);
nand U26459 (N_26459,N_25900,N_25150);
nand U26460 (N_26460,N_25633,N_25165);
nor U26461 (N_26461,N_25555,N_25105);
or U26462 (N_26462,N_25285,N_25373);
or U26463 (N_26463,N_25901,N_25396);
or U26464 (N_26464,N_25698,N_25221);
nand U26465 (N_26465,N_25470,N_25446);
nand U26466 (N_26466,N_25646,N_25093);
xnor U26467 (N_26467,N_25572,N_25341);
or U26468 (N_26468,N_25674,N_25071);
nor U26469 (N_26469,N_25483,N_25477);
nand U26470 (N_26470,N_25259,N_25229);
or U26471 (N_26471,N_25955,N_25928);
or U26472 (N_26472,N_25224,N_25379);
nor U26473 (N_26473,N_25231,N_25339);
or U26474 (N_26474,N_25479,N_25407);
xnor U26475 (N_26475,N_25152,N_25138);
or U26476 (N_26476,N_25675,N_25580);
and U26477 (N_26477,N_25449,N_25400);
or U26478 (N_26478,N_25578,N_25694);
or U26479 (N_26479,N_25797,N_25028);
or U26480 (N_26480,N_25022,N_25026);
nor U26481 (N_26481,N_25785,N_25656);
nand U26482 (N_26482,N_25335,N_25066);
nand U26483 (N_26483,N_25575,N_25918);
and U26484 (N_26484,N_25872,N_25940);
and U26485 (N_26485,N_25478,N_25924);
nand U26486 (N_26486,N_25080,N_25545);
or U26487 (N_26487,N_25081,N_25623);
nand U26488 (N_26488,N_25831,N_25178);
and U26489 (N_26489,N_25551,N_25328);
xnor U26490 (N_26490,N_25866,N_25556);
and U26491 (N_26491,N_25017,N_25543);
or U26492 (N_26492,N_25644,N_25615);
xnor U26493 (N_26493,N_25317,N_25309);
and U26494 (N_26494,N_25108,N_25194);
or U26495 (N_26495,N_25755,N_25504);
nand U26496 (N_26496,N_25207,N_25146);
or U26497 (N_26497,N_25264,N_25936);
and U26498 (N_26498,N_25038,N_25663);
or U26499 (N_26499,N_25732,N_25192);
nor U26500 (N_26500,N_25637,N_25533);
and U26501 (N_26501,N_25739,N_25772);
nor U26502 (N_26502,N_25493,N_25598);
nor U26503 (N_26503,N_25879,N_25690);
nor U26504 (N_26504,N_25122,N_25584);
nand U26505 (N_26505,N_25614,N_25502);
nand U26506 (N_26506,N_25642,N_25062);
and U26507 (N_26507,N_25142,N_25982);
nand U26508 (N_26508,N_25716,N_25715);
and U26509 (N_26509,N_25203,N_25637);
xnor U26510 (N_26510,N_25709,N_25930);
xnor U26511 (N_26511,N_25626,N_25835);
or U26512 (N_26512,N_25049,N_25397);
xnor U26513 (N_26513,N_25226,N_25043);
xor U26514 (N_26514,N_25493,N_25819);
nand U26515 (N_26515,N_25586,N_25590);
nand U26516 (N_26516,N_25171,N_25815);
nand U26517 (N_26517,N_25957,N_25451);
nand U26518 (N_26518,N_25989,N_25264);
or U26519 (N_26519,N_25892,N_25071);
nor U26520 (N_26520,N_25575,N_25993);
nor U26521 (N_26521,N_25563,N_25095);
nor U26522 (N_26522,N_25879,N_25207);
xor U26523 (N_26523,N_25812,N_25429);
xor U26524 (N_26524,N_25541,N_25087);
nor U26525 (N_26525,N_25576,N_25620);
xor U26526 (N_26526,N_25928,N_25755);
and U26527 (N_26527,N_25094,N_25317);
xnor U26528 (N_26528,N_25445,N_25548);
or U26529 (N_26529,N_25820,N_25513);
and U26530 (N_26530,N_25497,N_25763);
and U26531 (N_26531,N_25095,N_25151);
and U26532 (N_26532,N_25617,N_25211);
and U26533 (N_26533,N_25098,N_25702);
xor U26534 (N_26534,N_25403,N_25418);
or U26535 (N_26535,N_25086,N_25495);
nor U26536 (N_26536,N_25691,N_25098);
nand U26537 (N_26537,N_25396,N_25264);
and U26538 (N_26538,N_25769,N_25140);
nand U26539 (N_26539,N_25567,N_25729);
or U26540 (N_26540,N_25024,N_25459);
xnor U26541 (N_26541,N_25509,N_25928);
or U26542 (N_26542,N_25636,N_25030);
and U26543 (N_26543,N_25728,N_25986);
and U26544 (N_26544,N_25108,N_25247);
xor U26545 (N_26545,N_25455,N_25070);
nor U26546 (N_26546,N_25034,N_25882);
nor U26547 (N_26547,N_25752,N_25266);
or U26548 (N_26548,N_25736,N_25666);
nor U26549 (N_26549,N_25756,N_25678);
xor U26550 (N_26550,N_25687,N_25633);
and U26551 (N_26551,N_25174,N_25954);
nand U26552 (N_26552,N_25611,N_25332);
and U26553 (N_26553,N_25175,N_25344);
and U26554 (N_26554,N_25817,N_25127);
or U26555 (N_26555,N_25203,N_25069);
or U26556 (N_26556,N_25175,N_25387);
nor U26557 (N_26557,N_25224,N_25347);
and U26558 (N_26558,N_25051,N_25596);
or U26559 (N_26559,N_25038,N_25727);
or U26560 (N_26560,N_25063,N_25338);
and U26561 (N_26561,N_25824,N_25870);
and U26562 (N_26562,N_25700,N_25494);
and U26563 (N_26563,N_25309,N_25905);
and U26564 (N_26564,N_25419,N_25507);
nand U26565 (N_26565,N_25818,N_25267);
xnor U26566 (N_26566,N_25573,N_25576);
nand U26567 (N_26567,N_25283,N_25312);
nor U26568 (N_26568,N_25099,N_25345);
or U26569 (N_26569,N_25057,N_25695);
nor U26570 (N_26570,N_25444,N_25597);
and U26571 (N_26571,N_25050,N_25961);
nor U26572 (N_26572,N_25001,N_25617);
or U26573 (N_26573,N_25000,N_25434);
xor U26574 (N_26574,N_25822,N_25315);
xnor U26575 (N_26575,N_25006,N_25803);
nor U26576 (N_26576,N_25503,N_25439);
or U26577 (N_26577,N_25286,N_25852);
xor U26578 (N_26578,N_25199,N_25932);
nand U26579 (N_26579,N_25696,N_25514);
or U26580 (N_26580,N_25682,N_25534);
or U26581 (N_26581,N_25483,N_25851);
xnor U26582 (N_26582,N_25074,N_25160);
or U26583 (N_26583,N_25100,N_25098);
xor U26584 (N_26584,N_25301,N_25161);
nor U26585 (N_26585,N_25293,N_25310);
or U26586 (N_26586,N_25790,N_25856);
nand U26587 (N_26587,N_25513,N_25844);
and U26588 (N_26588,N_25926,N_25410);
or U26589 (N_26589,N_25344,N_25195);
xor U26590 (N_26590,N_25864,N_25116);
or U26591 (N_26591,N_25871,N_25070);
nand U26592 (N_26592,N_25252,N_25977);
xnor U26593 (N_26593,N_25692,N_25211);
nand U26594 (N_26594,N_25958,N_25287);
xor U26595 (N_26595,N_25277,N_25204);
nand U26596 (N_26596,N_25230,N_25344);
or U26597 (N_26597,N_25169,N_25441);
or U26598 (N_26598,N_25272,N_25644);
or U26599 (N_26599,N_25033,N_25224);
nor U26600 (N_26600,N_25375,N_25120);
and U26601 (N_26601,N_25432,N_25470);
nor U26602 (N_26602,N_25878,N_25484);
or U26603 (N_26603,N_25954,N_25048);
nor U26604 (N_26604,N_25543,N_25218);
and U26605 (N_26605,N_25359,N_25317);
nor U26606 (N_26606,N_25389,N_25794);
nand U26607 (N_26607,N_25025,N_25745);
or U26608 (N_26608,N_25260,N_25129);
xor U26609 (N_26609,N_25187,N_25931);
nand U26610 (N_26610,N_25031,N_25925);
nand U26611 (N_26611,N_25909,N_25291);
nor U26612 (N_26612,N_25713,N_25570);
nor U26613 (N_26613,N_25995,N_25798);
nor U26614 (N_26614,N_25844,N_25736);
and U26615 (N_26615,N_25147,N_25595);
nor U26616 (N_26616,N_25626,N_25995);
or U26617 (N_26617,N_25108,N_25736);
xor U26618 (N_26618,N_25733,N_25397);
nor U26619 (N_26619,N_25957,N_25117);
and U26620 (N_26620,N_25793,N_25455);
nand U26621 (N_26621,N_25788,N_25089);
nand U26622 (N_26622,N_25603,N_25756);
nor U26623 (N_26623,N_25731,N_25321);
nand U26624 (N_26624,N_25232,N_25220);
nand U26625 (N_26625,N_25422,N_25562);
and U26626 (N_26626,N_25989,N_25710);
nor U26627 (N_26627,N_25514,N_25193);
or U26628 (N_26628,N_25224,N_25165);
xor U26629 (N_26629,N_25099,N_25802);
nand U26630 (N_26630,N_25582,N_25695);
nand U26631 (N_26631,N_25877,N_25554);
and U26632 (N_26632,N_25751,N_25006);
or U26633 (N_26633,N_25943,N_25789);
nor U26634 (N_26634,N_25854,N_25105);
or U26635 (N_26635,N_25053,N_25874);
and U26636 (N_26636,N_25402,N_25103);
nand U26637 (N_26637,N_25419,N_25552);
and U26638 (N_26638,N_25465,N_25318);
nand U26639 (N_26639,N_25582,N_25062);
nor U26640 (N_26640,N_25054,N_25875);
and U26641 (N_26641,N_25616,N_25436);
or U26642 (N_26642,N_25082,N_25393);
xnor U26643 (N_26643,N_25346,N_25132);
nand U26644 (N_26644,N_25299,N_25032);
xnor U26645 (N_26645,N_25006,N_25619);
and U26646 (N_26646,N_25039,N_25663);
and U26647 (N_26647,N_25936,N_25042);
or U26648 (N_26648,N_25663,N_25583);
or U26649 (N_26649,N_25155,N_25400);
or U26650 (N_26650,N_25038,N_25273);
nor U26651 (N_26651,N_25813,N_25773);
or U26652 (N_26652,N_25019,N_25157);
nor U26653 (N_26653,N_25638,N_25016);
and U26654 (N_26654,N_25294,N_25456);
xnor U26655 (N_26655,N_25490,N_25889);
and U26656 (N_26656,N_25517,N_25893);
nor U26657 (N_26657,N_25151,N_25862);
or U26658 (N_26658,N_25347,N_25392);
and U26659 (N_26659,N_25993,N_25186);
or U26660 (N_26660,N_25663,N_25661);
nand U26661 (N_26661,N_25434,N_25518);
nor U26662 (N_26662,N_25027,N_25300);
xor U26663 (N_26663,N_25857,N_25954);
or U26664 (N_26664,N_25568,N_25756);
or U26665 (N_26665,N_25944,N_25643);
nand U26666 (N_26666,N_25536,N_25770);
nor U26667 (N_26667,N_25143,N_25838);
xnor U26668 (N_26668,N_25564,N_25474);
nand U26669 (N_26669,N_25228,N_25850);
xor U26670 (N_26670,N_25014,N_25934);
nand U26671 (N_26671,N_25995,N_25184);
nor U26672 (N_26672,N_25104,N_25949);
xnor U26673 (N_26673,N_25460,N_25723);
or U26674 (N_26674,N_25830,N_25166);
nor U26675 (N_26675,N_25253,N_25679);
and U26676 (N_26676,N_25516,N_25732);
xor U26677 (N_26677,N_25161,N_25355);
or U26678 (N_26678,N_25345,N_25310);
xor U26679 (N_26679,N_25661,N_25244);
xor U26680 (N_26680,N_25341,N_25658);
nand U26681 (N_26681,N_25097,N_25086);
xnor U26682 (N_26682,N_25310,N_25666);
or U26683 (N_26683,N_25731,N_25508);
nand U26684 (N_26684,N_25744,N_25614);
or U26685 (N_26685,N_25175,N_25343);
xnor U26686 (N_26686,N_25717,N_25571);
nand U26687 (N_26687,N_25756,N_25607);
and U26688 (N_26688,N_25262,N_25346);
nor U26689 (N_26689,N_25142,N_25869);
nor U26690 (N_26690,N_25736,N_25424);
nor U26691 (N_26691,N_25141,N_25383);
nand U26692 (N_26692,N_25073,N_25799);
nor U26693 (N_26693,N_25742,N_25906);
nor U26694 (N_26694,N_25609,N_25307);
xnor U26695 (N_26695,N_25886,N_25044);
nor U26696 (N_26696,N_25371,N_25132);
xnor U26697 (N_26697,N_25391,N_25089);
nor U26698 (N_26698,N_25804,N_25823);
and U26699 (N_26699,N_25479,N_25783);
xor U26700 (N_26700,N_25316,N_25614);
xnor U26701 (N_26701,N_25537,N_25699);
xor U26702 (N_26702,N_25452,N_25894);
or U26703 (N_26703,N_25256,N_25492);
or U26704 (N_26704,N_25097,N_25560);
nand U26705 (N_26705,N_25952,N_25452);
or U26706 (N_26706,N_25186,N_25179);
and U26707 (N_26707,N_25797,N_25386);
xor U26708 (N_26708,N_25675,N_25513);
nand U26709 (N_26709,N_25019,N_25002);
or U26710 (N_26710,N_25974,N_25637);
xnor U26711 (N_26711,N_25751,N_25206);
nor U26712 (N_26712,N_25858,N_25760);
nor U26713 (N_26713,N_25319,N_25700);
xor U26714 (N_26714,N_25695,N_25991);
xor U26715 (N_26715,N_25896,N_25093);
and U26716 (N_26716,N_25240,N_25356);
or U26717 (N_26717,N_25232,N_25878);
xnor U26718 (N_26718,N_25376,N_25634);
or U26719 (N_26719,N_25633,N_25249);
xnor U26720 (N_26720,N_25342,N_25668);
nor U26721 (N_26721,N_25806,N_25805);
and U26722 (N_26722,N_25345,N_25272);
and U26723 (N_26723,N_25256,N_25073);
nor U26724 (N_26724,N_25339,N_25273);
nand U26725 (N_26725,N_25847,N_25647);
or U26726 (N_26726,N_25422,N_25062);
or U26727 (N_26727,N_25148,N_25641);
xor U26728 (N_26728,N_25207,N_25031);
nand U26729 (N_26729,N_25255,N_25199);
nor U26730 (N_26730,N_25933,N_25810);
nand U26731 (N_26731,N_25646,N_25835);
and U26732 (N_26732,N_25201,N_25006);
or U26733 (N_26733,N_25266,N_25781);
or U26734 (N_26734,N_25110,N_25892);
xnor U26735 (N_26735,N_25915,N_25793);
or U26736 (N_26736,N_25381,N_25409);
xor U26737 (N_26737,N_25063,N_25003);
or U26738 (N_26738,N_25476,N_25365);
nand U26739 (N_26739,N_25137,N_25850);
and U26740 (N_26740,N_25702,N_25840);
xor U26741 (N_26741,N_25352,N_25915);
and U26742 (N_26742,N_25721,N_25224);
xor U26743 (N_26743,N_25370,N_25926);
nand U26744 (N_26744,N_25036,N_25424);
nand U26745 (N_26745,N_25024,N_25238);
or U26746 (N_26746,N_25042,N_25024);
or U26747 (N_26747,N_25566,N_25141);
and U26748 (N_26748,N_25475,N_25922);
and U26749 (N_26749,N_25982,N_25626);
nor U26750 (N_26750,N_25566,N_25147);
nand U26751 (N_26751,N_25352,N_25922);
nor U26752 (N_26752,N_25961,N_25489);
nor U26753 (N_26753,N_25122,N_25942);
nand U26754 (N_26754,N_25995,N_25437);
or U26755 (N_26755,N_25985,N_25033);
nor U26756 (N_26756,N_25773,N_25073);
xnor U26757 (N_26757,N_25308,N_25055);
and U26758 (N_26758,N_25759,N_25903);
nand U26759 (N_26759,N_25278,N_25055);
nor U26760 (N_26760,N_25458,N_25064);
nor U26761 (N_26761,N_25627,N_25158);
nor U26762 (N_26762,N_25652,N_25469);
nor U26763 (N_26763,N_25929,N_25934);
or U26764 (N_26764,N_25566,N_25836);
nor U26765 (N_26765,N_25989,N_25656);
nand U26766 (N_26766,N_25401,N_25837);
nor U26767 (N_26767,N_25573,N_25606);
nand U26768 (N_26768,N_25085,N_25393);
nor U26769 (N_26769,N_25111,N_25534);
nand U26770 (N_26770,N_25297,N_25215);
and U26771 (N_26771,N_25943,N_25167);
xor U26772 (N_26772,N_25575,N_25883);
xor U26773 (N_26773,N_25375,N_25813);
nor U26774 (N_26774,N_25770,N_25698);
nor U26775 (N_26775,N_25756,N_25168);
or U26776 (N_26776,N_25799,N_25434);
xnor U26777 (N_26777,N_25097,N_25658);
and U26778 (N_26778,N_25437,N_25861);
nand U26779 (N_26779,N_25331,N_25962);
nor U26780 (N_26780,N_25339,N_25264);
xnor U26781 (N_26781,N_25600,N_25797);
xnor U26782 (N_26782,N_25322,N_25403);
nor U26783 (N_26783,N_25078,N_25041);
nor U26784 (N_26784,N_25292,N_25791);
and U26785 (N_26785,N_25202,N_25893);
nand U26786 (N_26786,N_25927,N_25943);
or U26787 (N_26787,N_25651,N_25842);
nor U26788 (N_26788,N_25064,N_25179);
or U26789 (N_26789,N_25062,N_25405);
xnor U26790 (N_26790,N_25354,N_25521);
and U26791 (N_26791,N_25244,N_25978);
nand U26792 (N_26792,N_25130,N_25439);
nor U26793 (N_26793,N_25069,N_25725);
or U26794 (N_26794,N_25613,N_25262);
and U26795 (N_26795,N_25879,N_25375);
and U26796 (N_26796,N_25478,N_25381);
xor U26797 (N_26797,N_25819,N_25564);
and U26798 (N_26798,N_25023,N_25524);
or U26799 (N_26799,N_25031,N_25968);
xor U26800 (N_26800,N_25575,N_25050);
xor U26801 (N_26801,N_25185,N_25505);
nor U26802 (N_26802,N_25217,N_25248);
xnor U26803 (N_26803,N_25380,N_25066);
or U26804 (N_26804,N_25112,N_25852);
and U26805 (N_26805,N_25145,N_25716);
xor U26806 (N_26806,N_25827,N_25141);
and U26807 (N_26807,N_25226,N_25239);
or U26808 (N_26808,N_25440,N_25372);
or U26809 (N_26809,N_25862,N_25695);
and U26810 (N_26810,N_25334,N_25949);
nor U26811 (N_26811,N_25735,N_25375);
nor U26812 (N_26812,N_25781,N_25966);
nand U26813 (N_26813,N_25770,N_25576);
xor U26814 (N_26814,N_25981,N_25194);
nand U26815 (N_26815,N_25014,N_25640);
xnor U26816 (N_26816,N_25199,N_25289);
and U26817 (N_26817,N_25335,N_25090);
xor U26818 (N_26818,N_25274,N_25128);
and U26819 (N_26819,N_25161,N_25342);
nand U26820 (N_26820,N_25404,N_25415);
nor U26821 (N_26821,N_25543,N_25353);
nand U26822 (N_26822,N_25341,N_25408);
or U26823 (N_26823,N_25572,N_25688);
and U26824 (N_26824,N_25843,N_25675);
or U26825 (N_26825,N_25563,N_25668);
nand U26826 (N_26826,N_25779,N_25694);
nor U26827 (N_26827,N_25194,N_25786);
nor U26828 (N_26828,N_25844,N_25262);
nand U26829 (N_26829,N_25566,N_25090);
nand U26830 (N_26830,N_25092,N_25639);
nor U26831 (N_26831,N_25535,N_25578);
xor U26832 (N_26832,N_25537,N_25058);
and U26833 (N_26833,N_25735,N_25292);
nor U26834 (N_26834,N_25622,N_25426);
nor U26835 (N_26835,N_25124,N_25081);
nand U26836 (N_26836,N_25723,N_25213);
nor U26837 (N_26837,N_25289,N_25539);
or U26838 (N_26838,N_25749,N_25914);
or U26839 (N_26839,N_25853,N_25059);
nand U26840 (N_26840,N_25235,N_25490);
xor U26841 (N_26841,N_25346,N_25389);
and U26842 (N_26842,N_25246,N_25895);
nor U26843 (N_26843,N_25884,N_25531);
xnor U26844 (N_26844,N_25369,N_25185);
nand U26845 (N_26845,N_25731,N_25507);
xnor U26846 (N_26846,N_25221,N_25022);
nor U26847 (N_26847,N_25474,N_25810);
and U26848 (N_26848,N_25410,N_25031);
xnor U26849 (N_26849,N_25764,N_25221);
nand U26850 (N_26850,N_25923,N_25581);
and U26851 (N_26851,N_25533,N_25593);
and U26852 (N_26852,N_25841,N_25522);
or U26853 (N_26853,N_25712,N_25777);
xor U26854 (N_26854,N_25308,N_25012);
and U26855 (N_26855,N_25485,N_25743);
and U26856 (N_26856,N_25772,N_25412);
nor U26857 (N_26857,N_25011,N_25574);
xor U26858 (N_26858,N_25843,N_25967);
nor U26859 (N_26859,N_25204,N_25618);
nand U26860 (N_26860,N_25736,N_25471);
or U26861 (N_26861,N_25024,N_25185);
nor U26862 (N_26862,N_25924,N_25023);
or U26863 (N_26863,N_25156,N_25909);
nand U26864 (N_26864,N_25821,N_25843);
and U26865 (N_26865,N_25958,N_25899);
or U26866 (N_26866,N_25072,N_25822);
xnor U26867 (N_26867,N_25370,N_25186);
nor U26868 (N_26868,N_25490,N_25162);
nor U26869 (N_26869,N_25594,N_25737);
and U26870 (N_26870,N_25140,N_25945);
xor U26871 (N_26871,N_25894,N_25074);
xor U26872 (N_26872,N_25595,N_25255);
xnor U26873 (N_26873,N_25962,N_25549);
nor U26874 (N_26874,N_25238,N_25872);
nor U26875 (N_26875,N_25079,N_25447);
xnor U26876 (N_26876,N_25913,N_25918);
or U26877 (N_26877,N_25867,N_25299);
xor U26878 (N_26878,N_25096,N_25123);
xor U26879 (N_26879,N_25294,N_25280);
nor U26880 (N_26880,N_25687,N_25494);
and U26881 (N_26881,N_25885,N_25827);
and U26882 (N_26882,N_25085,N_25040);
xnor U26883 (N_26883,N_25845,N_25875);
or U26884 (N_26884,N_25750,N_25288);
and U26885 (N_26885,N_25000,N_25277);
and U26886 (N_26886,N_25857,N_25938);
and U26887 (N_26887,N_25352,N_25579);
xnor U26888 (N_26888,N_25083,N_25845);
and U26889 (N_26889,N_25707,N_25663);
nand U26890 (N_26890,N_25248,N_25917);
nand U26891 (N_26891,N_25310,N_25772);
nor U26892 (N_26892,N_25379,N_25456);
xor U26893 (N_26893,N_25673,N_25484);
nor U26894 (N_26894,N_25875,N_25678);
or U26895 (N_26895,N_25636,N_25427);
or U26896 (N_26896,N_25507,N_25610);
nor U26897 (N_26897,N_25322,N_25895);
or U26898 (N_26898,N_25345,N_25654);
nand U26899 (N_26899,N_25453,N_25404);
and U26900 (N_26900,N_25316,N_25026);
nor U26901 (N_26901,N_25341,N_25440);
nor U26902 (N_26902,N_25077,N_25243);
and U26903 (N_26903,N_25246,N_25714);
or U26904 (N_26904,N_25620,N_25077);
and U26905 (N_26905,N_25625,N_25849);
nand U26906 (N_26906,N_25403,N_25027);
xor U26907 (N_26907,N_25503,N_25888);
xnor U26908 (N_26908,N_25580,N_25026);
or U26909 (N_26909,N_25938,N_25316);
xor U26910 (N_26910,N_25311,N_25833);
nand U26911 (N_26911,N_25897,N_25877);
nor U26912 (N_26912,N_25025,N_25824);
nor U26913 (N_26913,N_25667,N_25482);
and U26914 (N_26914,N_25021,N_25602);
xnor U26915 (N_26915,N_25759,N_25746);
and U26916 (N_26916,N_25407,N_25436);
nand U26917 (N_26917,N_25636,N_25782);
nor U26918 (N_26918,N_25479,N_25109);
or U26919 (N_26919,N_25399,N_25468);
and U26920 (N_26920,N_25090,N_25246);
or U26921 (N_26921,N_25803,N_25531);
or U26922 (N_26922,N_25449,N_25131);
nand U26923 (N_26923,N_25068,N_25623);
xor U26924 (N_26924,N_25436,N_25568);
and U26925 (N_26925,N_25781,N_25478);
and U26926 (N_26926,N_25093,N_25033);
nor U26927 (N_26927,N_25192,N_25379);
xnor U26928 (N_26928,N_25656,N_25291);
nand U26929 (N_26929,N_25575,N_25207);
and U26930 (N_26930,N_25962,N_25400);
nand U26931 (N_26931,N_25873,N_25596);
and U26932 (N_26932,N_25393,N_25773);
and U26933 (N_26933,N_25898,N_25711);
nor U26934 (N_26934,N_25376,N_25156);
nand U26935 (N_26935,N_25576,N_25025);
or U26936 (N_26936,N_25308,N_25171);
nand U26937 (N_26937,N_25341,N_25168);
xor U26938 (N_26938,N_25695,N_25898);
or U26939 (N_26939,N_25484,N_25816);
xor U26940 (N_26940,N_25986,N_25548);
and U26941 (N_26941,N_25475,N_25061);
nand U26942 (N_26942,N_25225,N_25336);
xor U26943 (N_26943,N_25632,N_25179);
and U26944 (N_26944,N_25907,N_25322);
nor U26945 (N_26945,N_25109,N_25127);
nor U26946 (N_26946,N_25562,N_25898);
nand U26947 (N_26947,N_25689,N_25171);
nand U26948 (N_26948,N_25877,N_25873);
xnor U26949 (N_26949,N_25657,N_25550);
nand U26950 (N_26950,N_25559,N_25660);
and U26951 (N_26951,N_25286,N_25148);
nor U26952 (N_26952,N_25911,N_25159);
nor U26953 (N_26953,N_25050,N_25736);
or U26954 (N_26954,N_25395,N_25147);
and U26955 (N_26955,N_25432,N_25323);
xnor U26956 (N_26956,N_25456,N_25749);
or U26957 (N_26957,N_25875,N_25325);
nand U26958 (N_26958,N_25942,N_25341);
nand U26959 (N_26959,N_25570,N_25824);
xor U26960 (N_26960,N_25831,N_25804);
and U26961 (N_26961,N_25288,N_25033);
and U26962 (N_26962,N_25638,N_25251);
nand U26963 (N_26963,N_25931,N_25686);
nand U26964 (N_26964,N_25415,N_25902);
or U26965 (N_26965,N_25103,N_25113);
and U26966 (N_26966,N_25267,N_25969);
and U26967 (N_26967,N_25889,N_25287);
and U26968 (N_26968,N_25641,N_25766);
nand U26969 (N_26969,N_25620,N_25869);
xor U26970 (N_26970,N_25078,N_25853);
xnor U26971 (N_26971,N_25757,N_25172);
nor U26972 (N_26972,N_25625,N_25550);
and U26973 (N_26973,N_25120,N_25758);
xor U26974 (N_26974,N_25326,N_25427);
and U26975 (N_26975,N_25059,N_25753);
nand U26976 (N_26976,N_25102,N_25407);
and U26977 (N_26977,N_25596,N_25699);
nand U26978 (N_26978,N_25547,N_25916);
or U26979 (N_26979,N_25061,N_25899);
nand U26980 (N_26980,N_25722,N_25367);
and U26981 (N_26981,N_25624,N_25265);
and U26982 (N_26982,N_25993,N_25621);
nand U26983 (N_26983,N_25426,N_25156);
or U26984 (N_26984,N_25836,N_25121);
and U26985 (N_26985,N_25980,N_25924);
nand U26986 (N_26986,N_25758,N_25560);
xor U26987 (N_26987,N_25655,N_25129);
or U26988 (N_26988,N_25940,N_25206);
nand U26989 (N_26989,N_25914,N_25574);
or U26990 (N_26990,N_25593,N_25948);
xnor U26991 (N_26991,N_25570,N_25705);
and U26992 (N_26992,N_25348,N_25484);
and U26993 (N_26993,N_25658,N_25181);
or U26994 (N_26994,N_25955,N_25599);
and U26995 (N_26995,N_25394,N_25419);
nor U26996 (N_26996,N_25174,N_25778);
or U26997 (N_26997,N_25412,N_25213);
nand U26998 (N_26998,N_25200,N_25899);
nor U26999 (N_26999,N_25107,N_25793);
xnor U27000 (N_27000,N_26649,N_26504);
or U27001 (N_27001,N_26363,N_26611);
nand U27002 (N_27002,N_26928,N_26344);
and U27003 (N_27003,N_26285,N_26130);
nor U27004 (N_27004,N_26280,N_26132);
and U27005 (N_27005,N_26311,N_26510);
xnor U27006 (N_27006,N_26924,N_26807);
nand U27007 (N_27007,N_26004,N_26824);
and U27008 (N_27008,N_26442,N_26937);
and U27009 (N_27009,N_26377,N_26333);
nand U27010 (N_27010,N_26567,N_26214);
nor U27011 (N_27011,N_26638,N_26658);
nand U27012 (N_27012,N_26262,N_26181);
nor U27013 (N_27013,N_26691,N_26418);
xnor U27014 (N_27014,N_26234,N_26952);
xnor U27015 (N_27015,N_26917,N_26195);
xnor U27016 (N_27016,N_26131,N_26610);
or U27017 (N_27017,N_26136,N_26783);
and U27018 (N_27018,N_26562,N_26506);
or U27019 (N_27019,N_26207,N_26967);
nor U27020 (N_27020,N_26478,N_26466);
xnor U27021 (N_27021,N_26727,N_26641);
or U27022 (N_27022,N_26468,N_26457);
xor U27023 (N_27023,N_26444,N_26317);
xnor U27024 (N_27024,N_26372,N_26695);
and U27025 (N_27025,N_26472,N_26339);
xnor U27026 (N_27026,N_26559,N_26375);
nor U27027 (N_27027,N_26310,N_26153);
nand U27028 (N_27028,N_26565,N_26165);
xor U27029 (N_27029,N_26979,N_26024);
nor U27030 (N_27030,N_26172,N_26349);
and U27031 (N_27031,N_26830,N_26011);
and U27032 (N_27032,N_26421,N_26841);
nand U27033 (N_27033,N_26705,N_26330);
and U27034 (N_27034,N_26495,N_26086);
xor U27035 (N_27035,N_26296,N_26536);
or U27036 (N_27036,N_26343,N_26001);
nor U27037 (N_27037,N_26817,N_26167);
nand U27038 (N_27038,N_26930,N_26081);
nand U27039 (N_27039,N_26028,N_26596);
or U27040 (N_27040,N_26885,N_26406);
xor U27041 (N_27041,N_26745,N_26038);
nand U27042 (N_27042,N_26821,N_26211);
nand U27043 (N_27043,N_26877,N_26387);
nor U27044 (N_27044,N_26835,N_26795);
and U27045 (N_27045,N_26867,N_26199);
and U27046 (N_27046,N_26757,N_26042);
or U27047 (N_27047,N_26045,N_26668);
and U27048 (N_27048,N_26057,N_26840);
or U27049 (N_27049,N_26603,N_26923);
or U27050 (N_27050,N_26200,N_26946);
or U27051 (N_27051,N_26424,N_26855);
nor U27052 (N_27052,N_26053,N_26522);
nand U27053 (N_27053,N_26751,N_26893);
xnor U27054 (N_27054,N_26755,N_26312);
and U27055 (N_27055,N_26742,N_26412);
and U27056 (N_27056,N_26104,N_26802);
nand U27057 (N_27057,N_26989,N_26164);
nor U27058 (N_27058,N_26530,N_26715);
xnor U27059 (N_27059,N_26579,N_26849);
nor U27060 (N_27060,N_26119,N_26222);
nand U27061 (N_27061,N_26679,N_26281);
or U27062 (N_27062,N_26798,N_26204);
xnor U27063 (N_27063,N_26607,N_26963);
and U27064 (N_27064,N_26079,N_26574);
nand U27065 (N_27065,N_26950,N_26772);
or U27066 (N_27066,N_26974,N_26360);
xnor U27067 (N_27067,N_26110,N_26461);
xor U27068 (N_27068,N_26689,N_26434);
or U27069 (N_27069,N_26275,N_26797);
xor U27070 (N_27070,N_26020,N_26077);
nor U27071 (N_27071,N_26487,N_26135);
and U27072 (N_27072,N_26650,N_26010);
and U27073 (N_27073,N_26429,N_26021);
nor U27074 (N_27074,N_26926,N_26463);
nand U27075 (N_27075,N_26098,N_26123);
and U27076 (N_27076,N_26118,N_26710);
nor U27077 (N_27077,N_26701,N_26949);
nor U27078 (N_27078,N_26904,N_26388);
nand U27079 (N_27079,N_26585,N_26456);
nor U27080 (N_27080,N_26051,N_26625);
nand U27081 (N_27081,N_26964,N_26364);
and U27082 (N_27082,N_26147,N_26269);
and U27083 (N_27083,N_26815,N_26270);
nand U27084 (N_27084,N_26188,N_26245);
xnor U27085 (N_27085,N_26183,N_26527);
xnor U27086 (N_27086,N_26752,N_26383);
and U27087 (N_27087,N_26314,N_26455);
nor U27088 (N_27088,N_26279,N_26956);
xnor U27089 (N_27089,N_26988,N_26758);
or U27090 (N_27090,N_26178,N_26055);
nand U27091 (N_27091,N_26620,N_26337);
nand U27092 (N_27092,N_26670,N_26366);
nor U27093 (N_27093,N_26212,N_26600);
nand U27094 (N_27094,N_26739,N_26336);
nand U27095 (N_27095,N_26552,N_26619);
xnor U27096 (N_27096,N_26012,N_26109);
or U27097 (N_27097,N_26392,N_26987);
or U27098 (N_27098,N_26627,N_26533);
xnor U27099 (N_27099,N_26728,N_26346);
and U27100 (N_27100,N_26939,N_26931);
xnor U27101 (N_27101,N_26002,N_26523);
and U27102 (N_27102,N_26577,N_26688);
and U27103 (N_27103,N_26850,N_26919);
and U27104 (N_27104,N_26432,N_26390);
or U27105 (N_27105,N_26676,N_26187);
and U27106 (N_27106,N_26244,N_26108);
nand U27107 (N_27107,N_26661,N_26420);
or U27108 (N_27108,N_26839,N_26379);
nand U27109 (N_27109,N_26368,N_26161);
or U27110 (N_27110,N_26238,N_26229);
or U27111 (N_27111,N_26725,N_26851);
nand U27112 (N_27112,N_26210,N_26060);
or U27113 (N_27113,N_26401,N_26194);
and U27114 (N_27114,N_26976,N_26790);
xnor U27115 (N_27115,N_26961,N_26291);
nor U27116 (N_27116,N_26588,N_26677);
nor U27117 (N_27117,N_26697,N_26206);
nor U27118 (N_27118,N_26908,N_26553);
nand U27119 (N_27119,N_26804,N_26288);
or U27120 (N_27120,N_26571,N_26277);
or U27121 (N_27121,N_26237,N_26407);
xor U27122 (N_27122,N_26485,N_26606);
and U27123 (N_27123,N_26373,N_26943);
or U27124 (N_27124,N_26174,N_26655);
or U27125 (N_27125,N_26062,N_26496);
nor U27126 (N_27126,N_26694,N_26580);
xor U27127 (N_27127,N_26729,N_26030);
xnor U27128 (N_27128,N_26292,N_26326);
and U27129 (N_27129,N_26575,N_26539);
xnor U27130 (N_27130,N_26814,N_26228);
nor U27131 (N_27131,N_26233,N_26891);
nand U27132 (N_27132,N_26756,N_26091);
and U27133 (N_27133,N_26308,N_26692);
and U27134 (N_27134,N_26747,N_26293);
xor U27135 (N_27135,N_26043,N_26769);
nor U27136 (N_27136,N_26716,N_26225);
and U27137 (N_27137,N_26965,N_26230);
xnor U27138 (N_27138,N_26584,N_26449);
xnor U27139 (N_27139,N_26791,N_26111);
and U27140 (N_27140,N_26185,N_26134);
nand U27141 (N_27141,N_26665,N_26662);
nor U27142 (N_27142,N_26543,N_26871);
xnor U27143 (N_27143,N_26730,N_26991);
and U27144 (N_27144,N_26675,N_26452);
or U27145 (N_27145,N_26529,N_26499);
and U27146 (N_27146,N_26342,N_26750);
or U27147 (N_27147,N_26591,N_26309);
xnor U27148 (N_27148,N_26122,N_26378);
and U27149 (N_27149,N_26525,N_26160);
nor U27150 (N_27150,N_26374,N_26301);
nor U27151 (N_27151,N_26217,N_26569);
nor U27152 (N_27152,N_26226,N_26166);
nor U27153 (N_27153,N_26707,N_26700);
xor U27154 (N_27154,N_26353,N_26634);
nand U27155 (N_27155,N_26307,N_26604);
and U27156 (N_27156,N_26106,N_26356);
and U27157 (N_27157,N_26984,N_26789);
or U27158 (N_27158,N_26905,N_26371);
or U27159 (N_27159,N_26345,N_26640);
or U27160 (N_27160,N_26394,N_26203);
xnor U27161 (N_27161,N_26819,N_26957);
or U27162 (N_27162,N_26545,N_26273);
and U27163 (N_27163,N_26663,N_26427);
nor U27164 (N_27164,N_26932,N_26143);
nand U27165 (N_27165,N_26329,N_26355);
xnor U27166 (N_27166,N_26083,N_26423);
and U27167 (N_27167,N_26486,N_26834);
nor U27168 (N_27168,N_26287,N_26706);
xor U27169 (N_27169,N_26327,N_26067);
or U27170 (N_27170,N_26760,N_26501);
and U27171 (N_27171,N_26537,N_26713);
or U27172 (N_27172,N_26737,N_26922);
nor U27173 (N_27173,N_26886,N_26405);
xor U27174 (N_27174,N_26402,N_26861);
nand U27175 (N_27175,N_26538,N_26248);
nor U27176 (N_27176,N_26911,N_26007);
and U27177 (N_27177,N_26828,N_26652);
or U27178 (N_27178,N_26561,N_26438);
or U27179 (N_27179,N_26682,N_26896);
xor U27180 (N_27180,N_26236,N_26792);
nor U27181 (N_27181,N_26027,N_26940);
or U27182 (N_27182,N_26786,N_26140);
nor U27183 (N_27183,N_26920,N_26605);
nand U27184 (N_27184,N_26986,N_26155);
nor U27185 (N_27185,N_26836,N_26115);
and U27186 (N_27186,N_26476,N_26031);
xor U27187 (N_27187,N_26482,N_26818);
nand U27188 (N_27188,N_26875,N_26032);
and U27189 (N_27189,N_26026,N_26628);
xnor U27190 (N_27190,N_26799,N_26286);
nand U27191 (N_27191,N_26256,N_26162);
xnor U27192 (N_27192,N_26094,N_26048);
nand U27193 (N_27193,N_26602,N_26838);
xor U27194 (N_27194,N_26735,N_26813);
or U27195 (N_27195,N_26549,N_26630);
xor U27196 (N_27196,N_26151,N_26622);
xor U27197 (N_27197,N_26177,N_26419);
or U27198 (N_27198,N_26544,N_26064);
nand U27199 (N_27199,N_26657,N_26820);
nand U27200 (N_27200,N_26144,N_26594);
and U27201 (N_27201,N_26744,N_26842);
or U27202 (N_27202,N_26914,N_26899);
or U27203 (N_27203,N_26411,N_26191);
or U27204 (N_27204,N_26089,N_26389);
xnor U27205 (N_27205,N_26776,N_26554);
or U27206 (N_27206,N_26127,N_26175);
xor U27207 (N_27207,N_26848,N_26491);
or U27208 (N_27208,N_26669,N_26599);
nand U27209 (N_27209,N_26105,N_26075);
nand U27210 (N_27210,N_26775,N_26071);
or U27211 (N_27211,N_26430,N_26832);
xnor U27212 (N_27212,N_26748,N_26260);
nor U27213 (N_27213,N_26464,N_26722);
nand U27214 (N_27214,N_26152,N_26399);
nor U27215 (N_27215,N_26039,N_26723);
and U27216 (N_27216,N_26994,N_26889);
or U27217 (N_27217,N_26741,N_26137);
and U27218 (N_27218,N_26445,N_26516);
xnor U27219 (N_27219,N_26141,N_26541);
or U27220 (N_27220,N_26431,N_26887);
nor U27221 (N_27221,N_26856,N_26008);
xor U27222 (N_27222,N_26489,N_26941);
nor U27223 (N_27223,N_26673,N_26146);
nor U27224 (N_27224,N_26381,N_26453);
nor U27225 (N_27225,N_26500,N_26816);
nor U27226 (N_27226,N_26947,N_26972);
and U27227 (N_27227,N_26568,N_26654);
nor U27228 (N_27228,N_26671,N_26044);
or U27229 (N_27229,N_26050,N_26202);
nand U27230 (N_27230,N_26171,N_26117);
nand U27231 (N_27231,N_26651,N_26873);
or U27232 (N_27232,N_26250,N_26023);
or U27233 (N_27233,N_26114,N_26515);
nor U27234 (N_27234,N_26825,N_26995);
or U27235 (N_27235,N_26408,N_26517);
and U27236 (N_27236,N_26653,N_26674);
and U27237 (N_27237,N_26274,N_26944);
and U27238 (N_27238,N_26921,N_26384);
nor U27239 (N_27239,N_26636,N_26428);
and U27240 (N_27240,N_26558,N_26014);
nand U27241 (N_27241,N_26782,N_26805);
nor U27242 (N_27242,N_26738,N_26107);
or U27243 (N_27243,N_26519,N_26054);
nor U27244 (N_27244,N_26416,N_26550);
nor U27245 (N_27245,N_26948,N_26929);
and U27246 (N_27246,N_26034,N_26266);
and U27247 (N_27247,N_26590,N_26702);
and U27248 (N_27248,N_26507,N_26255);
xnor U27249 (N_27249,N_26681,N_26810);
nor U27250 (N_27250,N_26708,N_26773);
nand U27251 (N_27251,N_26036,N_26469);
nor U27252 (N_27252,N_26582,N_26216);
nand U27253 (N_27253,N_26827,N_26357);
xor U27254 (N_27254,N_26268,N_26150);
and U27255 (N_27255,N_26564,N_26992);
xnor U27256 (N_27256,N_26168,N_26184);
or U27257 (N_27257,N_26765,N_26788);
and U27258 (N_27258,N_26912,N_26592);
nand U27259 (N_27259,N_26304,N_26078);
xor U27260 (N_27260,N_26321,N_26863);
and U27261 (N_27261,N_26724,N_26733);
nor U27262 (N_27262,N_26844,N_26714);
nand U27263 (N_27263,N_26736,N_26779);
nor U27264 (N_27264,N_26398,N_26335);
nand U27265 (N_27265,N_26693,N_26243);
or U27266 (N_27266,N_26121,N_26699);
and U27267 (N_27267,N_26521,N_26837);
xnor U27268 (N_27268,N_26595,N_26935);
nor U27269 (N_27269,N_26743,N_26581);
nand U27270 (N_27270,N_26099,N_26720);
nor U27271 (N_27271,N_26283,N_26126);
nor U27272 (N_27272,N_26158,N_26125);
nor U27273 (N_27273,N_26186,N_26148);
or U27274 (N_27274,N_26102,N_26511);
or U27275 (N_27275,N_26593,N_26843);
or U27276 (N_27276,N_26859,N_26660);
nand U27277 (N_27277,N_26801,N_26483);
and U27278 (N_27278,N_26953,N_26719);
nor U27279 (N_27279,N_26272,N_26305);
and U27280 (N_27280,N_26629,N_26382);
or U27281 (N_27281,N_26770,N_26112);
or U27282 (N_27282,N_26440,N_26936);
or U27283 (N_27283,N_26116,N_26883);
or U27284 (N_27284,N_26531,N_26473);
xnor U27285 (N_27285,N_26910,N_26085);
and U27286 (N_27286,N_26025,N_26197);
nand U27287 (N_27287,N_26916,N_26201);
nor U27288 (N_27288,N_26746,N_26997);
and U27289 (N_27289,N_26433,N_26477);
nor U27290 (N_27290,N_26598,N_26215);
and U27291 (N_27291,N_26909,N_26073);
nor U27292 (N_27292,N_26365,N_26493);
or U27293 (N_27293,N_26563,N_26734);
or U27294 (N_27294,N_26000,N_26915);
xor U27295 (N_27295,N_26954,N_26113);
xnor U27296 (N_27296,N_26481,N_26703);
nand U27297 (N_27297,N_26632,N_26809);
or U27298 (N_27298,N_26016,N_26639);
nand U27299 (N_27299,N_26978,N_26072);
nor U27300 (N_27300,N_26812,N_26803);
xor U27301 (N_27301,N_26220,N_26231);
and U27302 (N_27302,N_26767,N_26196);
nand U27303 (N_27303,N_26369,N_26348);
nor U27304 (N_27304,N_26898,N_26513);
xnor U27305 (N_27305,N_26858,N_26257);
xnor U27306 (N_27306,N_26492,N_26359);
or U27307 (N_27307,N_26823,N_26251);
and U27308 (N_27308,N_26993,N_26781);
xor U27309 (N_27309,N_26762,N_26509);
nand U27310 (N_27310,N_26560,N_26505);
xor U27311 (N_27311,N_26644,N_26557);
or U27312 (N_27312,N_26683,N_26124);
or U27313 (N_27313,N_26475,N_26497);
nand U27314 (N_27314,N_26686,N_26066);
and U27315 (N_27315,N_26621,N_26518);
and U27316 (N_27316,N_26555,N_26971);
nand U27317 (N_27317,N_26249,N_26768);
and U27318 (N_27318,N_26052,N_26065);
xor U27319 (N_27319,N_26721,N_26864);
or U27320 (N_27320,N_26731,N_26777);
or U27321 (N_27321,N_26895,N_26774);
nand U27322 (N_27322,N_26906,N_26862);
nor U27323 (N_27323,N_26945,N_26901);
and U27324 (N_27324,N_26415,N_26190);
nor U27325 (N_27325,N_26845,N_26460);
xnor U27326 (N_27326,N_26796,N_26213);
nand U27327 (N_27327,N_26446,N_26631);
and U27328 (N_27328,N_26800,N_26439);
and U27329 (N_27329,N_26242,N_26996);
nor U27330 (N_27330,N_26092,N_26865);
and U27331 (N_27331,N_26753,N_26316);
or U27332 (N_27332,N_26435,N_26880);
and U27333 (N_27333,N_26890,N_26391);
xor U27334 (N_27334,N_26436,N_26869);
nor U27335 (N_27335,N_26614,N_26951);
xor U27336 (N_27336,N_26985,N_26189);
nor U27337 (N_27337,N_26302,N_26656);
xnor U27338 (N_27338,N_26586,N_26955);
nor U27339 (N_27339,N_26219,N_26903);
xor U27340 (N_27340,N_26370,N_26637);
or U27341 (N_27341,N_26540,N_26981);
nor U27342 (N_27342,N_26074,N_26358);
or U27343 (N_27343,N_26087,N_26278);
xor U27344 (N_27344,N_26006,N_26354);
nand U27345 (N_27345,N_26037,N_26209);
nand U27346 (N_27346,N_26892,N_26218);
and U27347 (N_27347,N_26297,N_26049);
and U27348 (N_27348,N_26443,N_26331);
nor U27349 (N_27349,N_26626,N_26404);
or U27350 (N_27350,N_26300,N_26350);
nor U27351 (N_27351,N_26526,N_26528);
nand U27352 (N_27352,N_26340,N_26872);
xor U27353 (N_27353,N_26176,N_26860);
nand U27354 (N_27354,N_26341,N_26018);
xor U27355 (N_27355,N_26717,N_26019);
or U27356 (N_27356,N_26618,N_26409);
and U27357 (N_27357,N_26534,N_26712);
nor U27358 (N_27358,N_26942,N_26437);
xnor U27359 (N_27359,N_26458,N_26448);
and U27360 (N_27360,N_26041,N_26033);
and U27361 (N_27361,N_26982,N_26173);
nand U27362 (N_27362,N_26179,N_26462);
or U27363 (N_27363,N_26410,N_26902);
xnor U27364 (N_27364,N_26780,N_26646);
and U27365 (N_27365,N_26246,N_26267);
and U27366 (N_27366,N_26351,N_26857);
and U27367 (N_27367,N_26022,N_26088);
xnor U27368 (N_27368,N_26447,N_26938);
and U27369 (N_27369,N_26778,N_26400);
nor U27370 (N_27370,N_26573,N_26556);
or U27371 (N_27371,N_26223,N_26015);
nor U27372 (N_27372,N_26977,N_26422);
nor U27373 (N_27373,N_26395,N_26347);
and U27374 (N_27374,N_26385,N_26494);
and U27375 (N_27375,N_26253,N_26047);
nor U27376 (N_27376,N_26056,N_26264);
and U27377 (N_27377,N_26532,N_26298);
or U27378 (N_27378,N_26068,N_26450);
nand U27379 (N_27379,N_26154,N_26766);
or U27380 (N_27380,N_26484,N_26271);
xnor U27381 (N_27381,N_26069,N_26666);
nand U27382 (N_27382,N_26680,N_26009);
and U27383 (N_27383,N_26005,N_26076);
nand U27384 (N_27384,N_26058,N_26315);
nand U27385 (N_27385,N_26958,N_26925);
or U27386 (N_27386,N_26240,N_26361);
and U27387 (N_27387,N_26846,N_26740);
xnor U27388 (N_27388,N_26328,N_26470);
nand U27389 (N_27389,N_26542,N_26474);
nand U27390 (N_27390,N_26969,N_26601);
nand U27391 (N_27391,N_26624,N_26918);
nand U27392 (N_27392,N_26927,N_26403);
xnor U27393 (N_27393,N_26295,N_26794);
or U27394 (N_27394,N_26535,N_26138);
and U27395 (N_27395,N_26454,N_26589);
nand U27396 (N_27396,N_26096,N_26608);
nand U27397 (N_27397,N_26261,N_26913);
and U27398 (N_27398,N_26771,N_26870);
nor U27399 (N_27399,N_26247,N_26306);
or U27400 (N_27400,N_26672,N_26129);
and U27401 (N_27401,N_26142,N_26046);
or U27402 (N_27402,N_26612,N_26546);
and U27403 (N_27403,N_26718,N_26570);
nand U27404 (N_27404,N_26764,N_26061);
nor U27405 (N_27405,N_26959,N_26386);
nand U27406 (N_27406,N_26808,N_26498);
xor U27407 (N_27407,N_26459,N_26633);
and U27408 (N_27408,N_26894,N_26084);
xor U27409 (N_27409,N_26761,N_26696);
nand U27410 (N_27410,N_26063,N_26029);
xor U27411 (N_27411,N_26467,N_26367);
xnor U27412 (N_27412,N_26149,N_26684);
nor U27413 (N_27413,N_26881,N_26999);
xor U27414 (N_27414,N_26299,N_26876);
nand U27415 (N_27415,N_26678,N_26265);
nor U27416 (N_27416,N_26145,N_26749);
and U27417 (N_27417,N_26879,N_26193);
or U27418 (N_27418,N_26362,N_26471);
or U27419 (N_27419,N_26566,N_26451);
nor U27420 (N_27420,N_26097,N_26334);
or U27421 (N_27421,N_26396,N_26616);
and U27422 (N_27422,N_26617,N_26294);
nor U27423 (N_27423,N_26934,N_26352);
nor U27424 (N_27424,N_26100,N_26254);
nor U27425 (N_27425,N_26208,N_26259);
and U27426 (N_27426,N_26320,N_26139);
and U27427 (N_27427,N_26615,N_26664);
or U27428 (N_27428,N_26325,N_26829);
and U27429 (N_27429,N_26159,N_26290);
and U27430 (N_27430,N_26831,N_26040);
and U27431 (N_27431,N_26643,N_26082);
xor U27432 (N_27432,N_26303,N_26441);
nand U27433 (N_27433,N_26572,N_26785);
nand U27434 (N_27434,N_26017,N_26613);
and U27435 (N_27435,N_26503,N_26623);
xor U27436 (N_27436,N_26853,N_26170);
and U27437 (N_27437,N_26480,N_26983);
xor U27438 (N_27438,N_26276,N_26192);
or U27439 (N_27439,N_26465,N_26642);
and U27440 (N_27440,N_26547,N_26900);
xnor U27441 (N_27441,N_26426,N_26332);
or U27442 (N_27442,N_26488,N_26587);
nand U27443 (N_27443,N_26597,N_26239);
xnor U27444 (N_27444,N_26520,N_26414);
xor U27445 (N_27445,N_26157,N_26080);
xor U27446 (N_27446,N_26787,N_26338);
and U27447 (N_27447,N_26854,N_26508);
nor U27448 (N_27448,N_26711,N_26826);
or U27449 (N_27449,N_26578,N_26224);
and U27450 (N_27450,N_26980,N_26897);
and U27451 (N_27451,N_26282,N_26120);
nor U27452 (N_27452,N_26784,N_26322);
or U27453 (N_27453,N_26704,N_26013);
nand U27454 (N_27454,N_26490,N_26709);
or U27455 (N_27455,N_26754,N_26156);
nor U27456 (N_27456,N_26133,N_26998);
or U27457 (N_27457,N_26907,N_26397);
nor U27458 (N_27458,N_26198,N_26690);
nand U27459 (N_27459,N_26833,N_26884);
xnor U27460 (N_27460,N_26793,N_26070);
xor U27461 (N_27461,N_26659,N_26095);
or U27462 (N_27462,N_26323,N_26852);
xnor U27463 (N_27463,N_26221,N_26933);
xor U27464 (N_27464,N_26966,N_26968);
nor U27465 (N_27465,N_26090,N_26313);
or U27466 (N_27466,N_26847,N_26289);
or U27467 (N_27467,N_26235,N_26227);
nor U27468 (N_27468,N_26417,N_26003);
or U27469 (N_27469,N_26685,N_26479);
nand U27470 (N_27470,N_26576,N_26413);
xor U27471 (N_27471,N_26059,N_26882);
and U27472 (N_27472,N_26609,N_26973);
xor U27473 (N_27473,N_26376,N_26514);
or U27474 (N_27474,N_26868,N_26635);
and U27475 (N_27475,N_26888,N_26667);
xnor U27476 (N_27476,N_26687,N_26425);
nand U27477 (N_27477,N_26698,N_26975);
nor U27478 (N_27478,N_26284,N_26878);
and U27479 (N_27479,N_26732,N_26180);
xnor U27480 (N_27480,N_26252,N_26866);
nand U27481 (N_27481,N_26103,N_26182);
or U27482 (N_27482,N_26318,N_26319);
nand U27483 (N_27483,N_26232,N_26093);
nand U27484 (N_27484,N_26324,N_26035);
nand U27485 (N_27485,N_26524,N_26645);
nor U27486 (N_27486,N_26806,N_26241);
nand U27487 (N_27487,N_26960,N_26647);
or U27488 (N_27488,N_26380,N_26205);
nand U27489 (N_27489,N_26551,N_26726);
nand U27490 (N_27490,N_26990,N_26763);
xnor U27491 (N_27491,N_26169,N_26101);
nand U27492 (N_27492,N_26258,N_26811);
or U27493 (N_27493,N_26822,N_26583);
nor U27494 (N_27494,N_26263,N_26962);
and U27495 (N_27495,N_26548,N_26163);
nand U27496 (N_27496,N_26512,N_26128);
xnor U27497 (N_27497,N_26970,N_26759);
and U27498 (N_27498,N_26648,N_26874);
nand U27499 (N_27499,N_26393,N_26502);
and U27500 (N_27500,N_26601,N_26141);
xor U27501 (N_27501,N_26749,N_26365);
and U27502 (N_27502,N_26513,N_26952);
nor U27503 (N_27503,N_26216,N_26689);
or U27504 (N_27504,N_26170,N_26480);
or U27505 (N_27505,N_26222,N_26671);
xor U27506 (N_27506,N_26601,N_26098);
nor U27507 (N_27507,N_26147,N_26746);
nand U27508 (N_27508,N_26315,N_26647);
xnor U27509 (N_27509,N_26452,N_26409);
and U27510 (N_27510,N_26555,N_26002);
nor U27511 (N_27511,N_26886,N_26691);
xor U27512 (N_27512,N_26427,N_26065);
nand U27513 (N_27513,N_26307,N_26459);
and U27514 (N_27514,N_26981,N_26615);
nand U27515 (N_27515,N_26183,N_26426);
or U27516 (N_27516,N_26389,N_26308);
and U27517 (N_27517,N_26892,N_26148);
xnor U27518 (N_27518,N_26155,N_26013);
xnor U27519 (N_27519,N_26550,N_26675);
or U27520 (N_27520,N_26495,N_26214);
xor U27521 (N_27521,N_26704,N_26131);
nand U27522 (N_27522,N_26395,N_26895);
nor U27523 (N_27523,N_26095,N_26606);
xnor U27524 (N_27524,N_26491,N_26463);
nand U27525 (N_27525,N_26618,N_26082);
xor U27526 (N_27526,N_26569,N_26088);
nand U27527 (N_27527,N_26348,N_26911);
or U27528 (N_27528,N_26778,N_26248);
xnor U27529 (N_27529,N_26807,N_26597);
nor U27530 (N_27530,N_26988,N_26458);
nand U27531 (N_27531,N_26324,N_26140);
and U27532 (N_27532,N_26909,N_26866);
and U27533 (N_27533,N_26932,N_26437);
and U27534 (N_27534,N_26977,N_26702);
xor U27535 (N_27535,N_26941,N_26275);
and U27536 (N_27536,N_26276,N_26012);
nor U27537 (N_27537,N_26566,N_26531);
or U27538 (N_27538,N_26057,N_26648);
nor U27539 (N_27539,N_26520,N_26453);
nor U27540 (N_27540,N_26980,N_26732);
and U27541 (N_27541,N_26205,N_26362);
nor U27542 (N_27542,N_26108,N_26650);
and U27543 (N_27543,N_26795,N_26820);
nor U27544 (N_27544,N_26561,N_26463);
xnor U27545 (N_27545,N_26481,N_26155);
xnor U27546 (N_27546,N_26450,N_26282);
or U27547 (N_27547,N_26481,N_26850);
xor U27548 (N_27548,N_26014,N_26428);
and U27549 (N_27549,N_26965,N_26540);
nor U27550 (N_27550,N_26543,N_26345);
and U27551 (N_27551,N_26107,N_26591);
and U27552 (N_27552,N_26073,N_26538);
nand U27553 (N_27553,N_26042,N_26144);
xor U27554 (N_27554,N_26695,N_26131);
nand U27555 (N_27555,N_26271,N_26182);
xnor U27556 (N_27556,N_26857,N_26849);
or U27557 (N_27557,N_26099,N_26365);
and U27558 (N_27558,N_26525,N_26240);
xnor U27559 (N_27559,N_26563,N_26779);
nor U27560 (N_27560,N_26291,N_26754);
or U27561 (N_27561,N_26163,N_26295);
and U27562 (N_27562,N_26500,N_26434);
or U27563 (N_27563,N_26895,N_26829);
and U27564 (N_27564,N_26221,N_26110);
and U27565 (N_27565,N_26304,N_26185);
xor U27566 (N_27566,N_26279,N_26427);
and U27567 (N_27567,N_26548,N_26190);
nand U27568 (N_27568,N_26598,N_26928);
xnor U27569 (N_27569,N_26573,N_26569);
nor U27570 (N_27570,N_26499,N_26939);
or U27571 (N_27571,N_26108,N_26025);
nor U27572 (N_27572,N_26037,N_26623);
xnor U27573 (N_27573,N_26917,N_26827);
nand U27574 (N_27574,N_26691,N_26534);
and U27575 (N_27575,N_26796,N_26019);
xnor U27576 (N_27576,N_26854,N_26743);
nand U27577 (N_27577,N_26981,N_26834);
nand U27578 (N_27578,N_26428,N_26706);
nand U27579 (N_27579,N_26685,N_26404);
and U27580 (N_27580,N_26690,N_26598);
and U27581 (N_27581,N_26188,N_26541);
and U27582 (N_27582,N_26544,N_26900);
xor U27583 (N_27583,N_26492,N_26892);
xnor U27584 (N_27584,N_26771,N_26592);
nand U27585 (N_27585,N_26059,N_26335);
nor U27586 (N_27586,N_26929,N_26955);
and U27587 (N_27587,N_26145,N_26888);
nand U27588 (N_27588,N_26548,N_26301);
xor U27589 (N_27589,N_26720,N_26671);
nand U27590 (N_27590,N_26355,N_26334);
xnor U27591 (N_27591,N_26004,N_26837);
xor U27592 (N_27592,N_26093,N_26214);
nand U27593 (N_27593,N_26679,N_26953);
and U27594 (N_27594,N_26262,N_26285);
nand U27595 (N_27595,N_26610,N_26439);
or U27596 (N_27596,N_26509,N_26620);
or U27597 (N_27597,N_26686,N_26224);
nor U27598 (N_27598,N_26631,N_26346);
or U27599 (N_27599,N_26628,N_26060);
nor U27600 (N_27600,N_26281,N_26950);
nor U27601 (N_27601,N_26714,N_26201);
or U27602 (N_27602,N_26923,N_26029);
or U27603 (N_27603,N_26921,N_26161);
or U27604 (N_27604,N_26899,N_26070);
or U27605 (N_27605,N_26385,N_26188);
or U27606 (N_27606,N_26678,N_26396);
and U27607 (N_27607,N_26157,N_26842);
and U27608 (N_27608,N_26219,N_26041);
nand U27609 (N_27609,N_26500,N_26228);
or U27610 (N_27610,N_26024,N_26239);
and U27611 (N_27611,N_26820,N_26885);
nand U27612 (N_27612,N_26895,N_26442);
or U27613 (N_27613,N_26752,N_26198);
or U27614 (N_27614,N_26458,N_26310);
or U27615 (N_27615,N_26066,N_26919);
and U27616 (N_27616,N_26760,N_26473);
nand U27617 (N_27617,N_26100,N_26645);
nor U27618 (N_27618,N_26748,N_26419);
or U27619 (N_27619,N_26714,N_26150);
and U27620 (N_27620,N_26767,N_26283);
nor U27621 (N_27621,N_26275,N_26672);
and U27622 (N_27622,N_26625,N_26554);
xnor U27623 (N_27623,N_26235,N_26555);
nand U27624 (N_27624,N_26558,N_26229);
and U27625 (N_27625,N_26525,N_26898);
and U27626 (N_27626,N_26043,N_26771);
nand U27627 (N_27627,N_26391,N_26076);
and U27628 (N_27628,N_26209,N_26934);
nor U27629 (N_27629,N_26889,N_26724);
nor U27630 (N_27630,N_26874,N_26109);
and U27631 (N_27631,N_26650,N_26360);
or U27632 (N_27632,N_26381,N_26749);
xor U27633 (N_27633,N_26790,N_26355);
nor U27634 (N_27634,N_26234,N_26896);
xnor U27635 (N_27635,N_26268,N_26159);
xnor U27636 (N_27636,N_26059,N_26298);
or U27637 (N_27637,N_26233,N_26497);
and U27638 (N_27638,N_26463,N_26298);
xnor U27639 (N_27639,N_26732,N_26738);
xor U27640 (N_27640,N_26770,N_26283);
or U27641 (N_27641,N_26343,N_26678);
nor U27642 (N_27642,N_26312,N_26962);
and U27643 (N_27643,N_26859,N_26886);
and U27644 (N_27644,N_26722,N_26543);
or U27645 (N_27645,N_26018,N_26129);
xnor U27646 (N_27646,N_26998,N_26201);
or U27647 (N_27647,N_26698,N_26132);
xnor U27648 (N_27648,N_26898,N_26203);
or U27649 (N_27649,N_26530,N_26072);
or U27650 (N_27650,N_26800,N_26846);
xnor U27651 (N_27651,N_26356,N_26917);
and U27652 (N_27652,N_26447,N_26735);
or U27653 (N_27653,N_26217,N_26105);
xnor U27654 (N_27654,N_26321,N_26882);
nand U27655 (N_27655,N_26543,N_26542);
and U27656 (N_27656,N_26412,N_26891);
xnor U27657 (N_27657,N_26686,N_26431);
nor U27658 (N_27658,N_26614,N_26801);
xnor U27659 (N_27659,N_26279,N_26131);
nor U27660 (N_27660,N_26760,N_26111);
and U27661 (N_27661,N_26485,N_26058);
nand U27662 (N_27662,N_26376,N_26969);
and U27663 (N_27663,N_26462,N_26606);
or U27664 (N_27664,N_26252,N_26584);
nor U27665 (N_27665,N_26439,N_26783);
xor U27666 (N_27666,N_26378,N_26026);
xnor U27667 (N_27667,N_26609,N_26619);
xor U27668 (N_27668,N_26515,N_26320);
or U27669 (N_27669,N_26731,N_26099);
nand U27670 (N_27670,N_26449,N_26615);
nor U27671 (N_27671,N_26539,N_26728);
nor U27672 (N_27672,N_26078,N_26824);
nor U27673 (N_27673,N_26488,N_26455);
nand U27674 (N_27674,N_26962,N_26597);
and U27675 (N_27675,N_26886,N_26509);
or U27676 (N_27676,N_26751,N_26556);
and U27677 (N_27677,N_26941,N_26436);
nand U27678 (N_27678,N_26360,N_26313);
nor U27679 (N_27679,N_26867,N_26233);
or U27680 (N_27680,N_26565,N_26763);
nor U27681 (N_27681,N_26009,N_26132);
nor U27682 (N_27682,N_26724,N_26665);
xor U27683 (N_27683,N_26745,N_26957);
xnor U27684 (N_27684,N_26253,N_26068);
xor U27685 (N_27685,N_26366,N_26315);
xnor U27686 (N_27686,N_26705,N_26908);
and U27687 (N_27687,N_26019,N_26384);
nor U27688 (N_27688,N_26607,N_26465);
or U27689 (N_27689,N_26521,N_26734);
or U27690 (N_27690,N_26290,N_26785);
and U27691 (N_27691,N_26492,N_26805);
xor U27692 (N_27692,N_26835,N_26501);
nand U27693 (N_27693,N_26800,N_26228);
xor U27694 (N_27694,N_26543,N_26562);
nor U27695 (N_27695,N_26209,N_26199);
nand U27696 (N_27696,N_26428,N_26959);
or U27697 (N_27697,N_26068,N_26368);
xnor U27698 (N_27698,N_26104,N_26609);
xor U27699 (N_27699,N_26117,N_26542);
xor U27700 (N_27700,N_26995,N_26247);
nand U27701 (N_27701,N_26645,N_26356);
and U27702 (N_27702,N_26545,N_26234);
xnor U27703 (N_27703,N_26969,N_26442);
and U27704 (N_27704,N_26943,N_26977);
nor U27705 (N_27705,N_26478,N_26917);
nor U27706 (N_27706,N_26539,N_26386);
or U27707 (N_27707,N_26055,N_26002);
xnor U27708 (N_27708,N_26929,N_26386);
nand U27709 (N_27709,N_26551,N_26202);
and U27710 (N_27710,N_26107,N_26322);
and U27711 (N_27711,N_26385,N_26671);
nand U27712 (N_27712,N_26728,N_26104);
nand U27713 (N_27713,N_26910,N_26594);
nand U27714 (N_27714,N_26028,N_26254);
nand U27715 (N_27715,N_26136,N_26694);
and U27716 (N_27716,N_26587,N_26927);
or U27717 (N_27717,N_26828,N_26716);
or U27718 (N_27718,N_26727,N_26456);
nand U27719 (N_27719,N_26980,N_26918);
nor U27720 (N_27720,N_26941,N_26685);
nand U27721 (N_27721,N_26517,N_26655);
nand U27722 (N_27722,N_26086,N_26157);
xnor U27723 (N_27723,N_26591,N_26758);
and U27724 (N_27724,N_26039,N_26325);
and U27725 (N_27725,N_26137,N_26731);
or U27726 (N_27726,N_26721,N_26598);
nand U27727 (N_27727,N_26916,N_26310);
nor U27728 (N_27728,N_26988,N_26138);
or U27729 (N_27729,N_26724,N_26760);
nand U27730 (N_27730,N_26224,N_26006);
nand U27731 (N_27731,N_26064,N_26104);
xor U27732 (N_27732,N_26197,N_26179);
or U27733 (N_27733,N_26480,N_26771);
xor U27734 (N_27734,N_26513,N_26521);
xor U27735 (N_27735,N_26968,N_26278);
nor U27736 (N_27736,N_26952,N_26865);
xor U27737 (N_27737,N_26772,N_26996);
or U27738 (N_27738,N_26472,N_26314);
xor U27739 (N_27739,N_26562,N_26806);
xnor U27740 (N_27740,N_26755,N_26695);
nand U27741 (N_27741,N_26281,N_26268);
nand U27742 (N_27742,N_26507,N_26403);
nand U27743 (N_27743,N_26171,N_26256);
nand U27744 (N_27744,N_26396,N_26348);
and U27745 (N_27745,N_26628,N_26170);
xnor U27746 (N_27746,N_26121,N_26620);
nor U27747 (N_27747,N_26217,N_26219);
nor U27748 (N_27748,N_26197,N_26690);
xnor U27749 (N_27749,N_26064,N_26215);
and U27750 (N_27750,N_26848,N_26465);
nand U27751 (N_27751,N_26144,N_26980);
or U27752 (N_27752,N_26214,N_26722);
or U27753 (N_27753,N_26935,N_26498);
or U27754 (N_27754,N_26623,N_26529);
or U27755 (N_27755,N_26963,N_26380);
nand U27756 (N_27756,N_26550,N_26751);
nand U27757 (N_27757,N_26289,N_26962);
nand U27758 (N_27758,N_26014,N_26669);
nor U27759 (N_27759,N_26375,N_26468);
xor U27760 (N_27760,N_26216,N_26530);
and U27761 (N_27761,N_26035,N_26615);
nor U27762 (N_27762,N_26077,N_26797);
or U27763 (N_27763,N_26083,N_26987);
and U27764 (N_27764,N_26208,N_26886);
nand U27765 (N_27765,N_26935,N_26273);
nand U27766 (N_27766,N_26852,N_26648);
xnor U27767 (N_27767,N_26828,N_26359);
nand U27768 (N_27768,N_26916,N_26589);
and U27769 (N_27769,N_26947,N_26437);
nand U27770 (N_27770,N_26032,N_26754);
nor U27771 (N_27771,N_26225,N_26166);
nand U27772 (N_27772,N_26782,N_26262);
nand U27773 (N_27773,N_26387,N_26632);
nand U27774 (N_27774,N_26951,N_26727);
and U27775 (N_27775,N_26908,N_26352);
and U27776 (N_27776,N_26974,N_26471);
xor U27777 (N_27777,N_26686,N_26326);
nor U27778 (N_27778,N_26545,N_26094);
or U27779 (N_27779,N_26617,N_26229);
nand U27780 (N_27780,N_26426,N_26610);
and U27781 (N_27781,N_26402,N_26474);
nand U27782 (N_27782,N_26173,N_26193);
xnor U27783 (N_27783,N_26474,N_26665);
nand U27784 (N_27784,N_26746,N_26688);
xor U27785 (N_27785,N_26517,N_26977);
or U27786 (N_27786,N_26207,N_26179);
or U27787 (N_27787,N_26342,N_26593);
or U27788 (N_27788,N_26321,N_26503);
and U27789 (N_27789,N_26083,N_26550);
xor U27790 (N_27790,N_26270,N_26495);
or U27791 (N_27791,N_26133,N_26247);
nand U27792 (N_27792,N_26320,N_26469);
xnor U27793 (N_27793,N_26474,N_26395);
and U27794 (N_27794,N_26196,N_26707);
or U27795 (N_27795,N_26540,N_26782);
or U27796 (N_27796,N_26578,N_26767);
nor U27797 (N_27797,N_26907,N_26966);
nand U27798 (N_27798,N_26236,N_26213);
nand U27799 (N_27799,N_26129,N_26790);
or U27800 (N_27800,N_26285,N_26855);
and U27801 (N_27801,N_26563,N_26918);
or U27802 (N_27802,N_26523,N_26042);
nor U27803 (N_27803,N_26088,N_26535);
or U27804 (N_27804,N_26004,N_26211);
or U27805 (N_27805,N_26564,N_26630);
or U27806 (N_27806,N_26128,N_26131);
nor U27807 (N_27807,N_26336,N_26200);
nand U27808 (N_27808,N_26892,N_26769);
xor U27809 (N_27809,N_26683,N_26918);
and U27810 (N_27810,N_26919,N_26535);
nor U27811 (N_27811,N_26882,N_26856);
and U27812 (N_27812,N_26130,N_26722);
or U27813 (N_27813,N_26135,N_26089);
nor U27814 (N_27814,N_26892,N_26470);
or U27815 (N_27815,N_26309,N_26468);
nor U27816 (N_27816,N_26726,N_26362);
or U27817 (N_27817,N_26910,N_26927);
xor U27818 (N_27818,N_26819,N_26552);
xnor U27819 (N_27819,N_26833,N_26249);
or U27820 (N_27820,N_26099,N_26735);
xor U27821 (N_27821,N_26123,N_26685);
nand U27822 (N_27822,N_26117,N_26792);
xnor U27823 (N_27823,N_26732,N_26327);
and U27824 (N_27824,N_26952,N_26283);
nand U27825 (N_27825,N_26668,N_26958);
or U27826 (N_27826,N_26255,N_26974);
xor U27827 (N_27827,N_26866,N_26250);
nor U27828 (N_27828,N_26729,N_26828);
nand U27829 (N_27829,N_26122,N_26838);
nand U27830 (N_27830,N_26351,N_26807);
nor U27831 (N_27831,N_26878,N_26211);
and U27832 (N_27832,N_26912,N_26844);
nor U27833 (N_27833,N_26758,N_26301);
xor U27834 (N_27834,N_26784,N_26807);
and U27835 (N_27835,N_26476,N_26276);
or U27836 (N_27836,N_26319,N_26559);
nand U27837 (N_27837,N_26397,N_26172);
or U27838 (N_27838,N_26538,N_26242);
nor U27839 (N_27839,N_26346,N_26085);
or U27840 (N_27840,N_26332,N_26985);
or U27841 (N_27841,N_26039,N_26252);
nor U27842 (N_27842,N_26648,N_26685);
nor U27843 (N_27843,N_26539,N_26125);
nand U27844 (N_27844,N_26695,N_26430);
nor U27845 (N_27845,N_26205,N_26496);
nand U27846 (N_27846,N_26986,N_26203);
nor U27847 (N_27847,N_26240,N_26540);
xor U27848 (N_27848,N_26316,N_26728);
nand U27849 (N_27849,N_26025,N_26876);
and U27850 (N_27850,N_26726,N_26227);
or U27851 (N_27851,N_26595,N_26154);
and U27852 (N_27852,N_26531,N_26764);
nand U27853 (N_27853,N_26465,N_26347);
and U27854 (N_27854,N_26751,N_26540);
nor U27855 (N_27855,N_26080,N_26550);
nand U27856 (N_27856,N_26094,N_26020);
and U27857 (N_27857,N_26131,N_26224);
and U27858 (N_27858,N_26504,N_26439);
nand U27859 (N_27859,N_26981,N_26000);
or U27860 (N_27860,N_26011,N_26426);
xnor U27861 (N_27861,N_26688,N_26732);
or U27862 (N_27862,N_26026,N_26853);
nand U27863 (N_27863,N_26983,N_26526);
or U27864 (N_27864,N_26038,N_26823);
or U27865 (N_27865,N_26339,N_26182);
xnor U27866 (N_27866,N_26203,N_26913);
nand U27867 (N_27867,N_26318,N_26991);
xnor U27868 (N_27868,N_26654,N_26040);
nand U27869 (N_27869,N_26311,N_26475);
and U27870 (N_27870,N_26351,N_26593);
and U27871 (N_27871,N_26996,N_26802);
and U27872 (N_27872,N_26235,N_26718);
xnor U27873 (N_27873,N_26886,N_26658);
and U27874 (N_27874,N_26355,N_26077);
or U27875 (N_27875,N_26504,N_26559);
nand U27876 (N_27876,N_26070,N_26919);
or U27877 (N_27877,N_26369,N_26127);
nand U27878 (N_27878,N_26750,N_26752);
or U27879 (N_27879,N_26184,N_26079);
xor U27880 (N_27880,N_26380,N_26361);
and U27881 (N_27881,N_26142,N_26601);
nand U27882 (N_27882,N_26894,N_26852);
xnor U27883 (N_27883,N_26927,N_26647);
xor U27884 (N_27884,N_26686,N_26999);
nor U27885 (N_27885,N_26139,N_26292);
and U27886 (N_27886,N_26207,N_26782);
xnor U27887 (N_27887,N_26261,N_26329);
and U27888 (N_27888,N_26315,N_26551);
nor U27889 (N_27889,N_26914,N_26105);
xnor U27890 (N_27890,N_26343,N_26707);
and U27891 (N_27891,N_26593,N_26474);
nand U27892 (N_27892,N_26415,N_26004);
nor U27893 (N_27893,N_26679,N_26673);
xor U27894 (N_27894,N_26549,N_26206);
nor U27895 (N_27895,N_26423,N_26586);
or U27896 (N_27896,N_26632,N_26325);
and U27897 (N_27897,N_26916,N_26691);
xor U27898 (N_27898,N_26333,N_26300);
nand U27899 (N_27899,N_26081,N_26876);
or U27900 (N_27900,N_26433,N_26311);
xnor U27901 (N_27901,N_26614,N_26002);
and U27902 (N_27902,N_26401,N_26221);
nor U27903 (N_27903,N_26873,N_26054);
and U27904 (N_27904,N_26134,N_26123);
or U27905 (N_27905,N_26224,N_26259);
xor U27906 (N_27906,N_26515,N_26613);
xnor U27907 (N_27907,N_26939,N_26301);
or U27908 (N_27908,N_26235,N_26433);
and U27909 (N_27909,N_26293,N_26515);
and U27910 (N_27910,N_26248,N_26691);
xor U27911 (N_27911,N_26603,N_26967);
nand U27912 (N_27912,N_26973,N_26831);
nand U27913 (N_27913,N_26879,N_26000);
or U27914 (N_27914,N_26904,N_26649);
xnor U27915 (N_27915,N_26286,N_26301);
or U27916 (N_27916,N_26851,N_26377);
nand U27917 (N_27917,N_26401,N_26269);
and U27918 (N_27918,N_26801,N_26851);
nand U27919 (N_27919,N_26128,N_26264);
nand U27920 (N_27920,N_26050,N_26954);
and U27921 (N_27921,N_26333,N_26827);
and U27922 (N_27922,N_26208,N_26100);
or U27923 (N_27923,N_26333,N_26794);
xor U27924 (N_27924,N_26924,N_26647);
or U27925 (N_27925,N_26709,N_26248);
or U27926 (N_27926,N_26044,N_26577);
xor U27927 (N_27927,N_26060,N_26647);
xor U27928 (N_27928,N_26940,N_26204);
nor U27929 (N_27929,N_26580,N_26968);
and U27930 (N_27930,N_26413,N_26931);
and U27931 (N_27931,N_26434,N_26378);
or U27932 (N_27932,N_26573,N_26835);
nand U27933 (N_27933,N_26284,N_26795);
or U27934 (N_27934,N_26949,N_26171);
nor U27935 (N_27935,N_26643,N_26021);
and U27936 (N_27936,N_26161,N_26367);
xor U27937 (N_27937,N_26055,N_26220);
and U27938 (N_27938,N_26749,N_26689);
xor U27939 (N_27939,N_26332,N_26964);
nor U27940 (N_27940,N_26126,N_26206);
nor U27941 (N_27941,N_26893,N_26463);
nand U27942 (N_27942,N_26932,N_26993);
xnor U27943 (N_27943,N_26534,N_26943);
nand U27944 (N_27944,N_26099,N_26933);
xnor U27945 (N_27945,N_26831,N_26721);
and U27946 (N_27946,N_26134,N_26935);
and U27947 (N_27947,N_26129,N_26301);
nor U27948 (N_27948,N_26038,N_26530);
and U27949 (N_27949,N_26194,N_26043);
nor U27950 (N_27950,N_26255,N_26213);
nand U27951 (N_27951,N_26027,N_26387);
nor U27952 (N_27952,N_26227,N_26417);
nor U27953 (N_27953,N_26297,N_26706);
nand U27954 (N_27954,N_26416,N_26242);
xor U27955 (N_27955,N_26081,N_26241);
and U27956 (N_27956,N_26316,N_26568);
nor U27957 (N_27957,N_26869,N_26228);
or U27958 (N_27958,N_26763,N_26961);
xnor U27959 (N_27959,N_26994,N_26460);
or U27960 (N_27960,N_26649,N_26880);
and U27961 (N_27961,N_26794,N_26212);
nand U27962 (N_27962,N_26054,N_26742);
nor U27963 (N_27963,N_26822,N_26892);
nand U27964 (N_27964,N_26676,N_26213);
and U27965 (N_27965,N_26941,N_26452);
nand U27966 (N_27966,N_26179,N_26593);
nor U27967 (N_27967,N_26672,N_26428);
nand U27968 (N_27968,N_26631,N_26335);
or U27969 (N_27969,N_26408,N_26284);
and U27970 (N_27970,N_26847,N_26860);
and U27971 (N_27971,N_26379,N_26797);
nor U27972 (N_27972,N_26885,N_26779);
xor U27973 (N_27973,N_26080,N_26095);
and U27974 (N_27974,N_26968,N_26087);
xnor U27975 (N_27975,N_26311,N_26467);
or U27976 (N_27976,N_26418,N_26409);
nor U27977 (N_27977,N_26145,N_26366);
and U27978 (N_27978,N_26807,N_26438);
or U27979 (N_27979,N_26284,N_26827);
nand U27980 (N_27980,N_26951,N_26019);
or U27981 (N_27981,N_26438,N_26441);
and U27982 (N_27982,N_26989,N_26603);
xor U27983 (N_27983,N_26416,N_26278);
nor U27984 (N_27984,N_26832,N_26593);
xor U27985 (N_27985,N_26440,N_26433);
nor U27986 (N_27986,N_26424,N_26830);
nor U27987 (N_27987,N_26885,N_26312);
nand U27988 (N_27988,N_26901,N_26041);
nor U27989 (N_27989,N_26504,N_26625);
nand U27990 (N_27990,N_26825,N_26424);
and U27991 (N_27991,N_26998,N_26407);
and U27992 (N_27992,N_26113,N_26363);
nor U27993 (N_27993,N_26761,N_26411);
xor U27994 (N_27994,N_26116,N_26684);
nand U27995 (N_27995,N_26859,N_26970);
xnor U27996 (N_27996,N_26492,N_26971);
nand U27997 (N_27997,N_26680,N_26568);
nor U27998 (N_27998,N_26128,N_26482);
nand U27999 (N_27999,N_26540,N_26067);
or U28000 (N_28000,N_27928,N_27596);
xor U28001 (N_28001,N_27372,N_27697);
or U28002 (N_28002,N_27259,N_27598);
xnor U28003 (N_28003,N_27740,N_27823);
or U28004 (N_28004,N_27100,N_27907);
nor U28005 (N_28005,N_27338,N_27156);
nand U28006 (N_28006,N_27786,N_27929);
and U28007 (N_28007,N_27850,N_27896);
and U28008 (N_28008,N_27130,N_27451);
nand U28009 (N_28009,N_27638,N_27951);
nand U28010 (N_28010,N_27166,N_27087);
and U28011 (N_28011,N_27898,N_27049);
nand U28012 (N_28012,N_27600,N_27893);
and U28013 (N_28013,N_27542,N_27281);
xnor U28014 (N_28014,N_27273,N_27168);
xor U28015 (N_28015,N_27107,N_27840);
or U28016 (N_28016,N_27733,N_27766);
nor U28017 (N_28017,N_27413,N_27262);
and U28018 (N_28018,N_27198,N_27484);
or U28019 (N_28019,N_27367,N_27085);
and U28020 (N_28020,N_27362,N_27467);
nand U28021 (N_28021,N_27861,N_27426);
xor U28022 (N_28022,N_27543,N_27581);
or U28023 (N_28023,N_27872,N_27573);
xor U28024 (N_28024,N_27317,N_27300);
xor U28025 (N_28025,N_27780,N_27552);
nor U28026 (N_28026,N_27479,N_27836);
or U28027 (N_28027,N_27597,N_27221);
and U28028 (N_28028,N_27775,N_27180);
nand U28029 (N_28029,N_27278,N_27205);
nand U28030 (N_28030,N_27648,N_27003);
nor U28031 (N_28031,N_27718,N_27226);
nand U28032 (N_28032,N_27095,N_27975);
nor U28033 (N_28033,N_27422,N_27610);
xnor U28034 (N_28034,N_27029,N_27974);
xor U28035 (N_28035,N_27043,N_27093);
xor U28036 (N_28036,N_27193,N_27761);
xnor U28037 (N_28037,N_27556,N_27507);
or U28038 (N_28038,N_27480,N_27323);
nand U28039 (N_28039,N_27572,N_27591);
nor U28040 (N_28040,N_27537,N_27616);
nor U28041 (N_28041,N_27204,N_27751);
xnor U28042 (N_28042,N_27808,N_27113);
nand U28043 (N_28043,N_27634,N_27324);
nor U28044 (N_28044,N_27511,N_27941);
or U28045 (N_28045,N_27406,N_27510);
nand U28046 (N_28046,N_27777,N_27134);
nor U28047 (N_28047,N_27410,N_27835);
xor U28048 (N_28048,N_27343,N_27890);
or U28049 (N_28049,N_27456,N_27897);
nor U28050 (N_28050,N_27964,N_27949);
and U28051 (N_28051,N_27715,N_27576);
nor U28052 (N_28052,N_27187,N_27879);
nand U28053 (N_28053,N_27709,N_27584);
xor U28054 (N_28054,N_27499,N_27837);
nand U28055 (N_28055,N_27383,N_27473);
and U28056 (N_28056,N_27684,N_27371);
and U28057 (N_28057,N_27059,N_27826);
nor U28058 (N_28058,N_27517,N_27212);
xor U28059 (N_28059,N_27398,N_27141);
and U28060 (N_28060,N_27232,N_27934);
nor U28061 (N_28061,N_27647,N_27804);
or U28062 (N_28062,N_27178,N_27959);
and U28063 (N_28063,N_27120,N_27478);
nor U28064 (N_28064,N_27755,N_27233);
nand U28065 (N_28065,N_27989,N_27326);
or U28066 (N_28066,N_27864,N_27222);
xnor U28067 (N_28067,N_27830,N_27018);
nand U28068 (N_28068,N_27827,N_27615);
xor U28069 (N_28069,N_27284,N_27143);
nor U28070 (N_28070,N_27762,N_27287);
xnor U28071 (N_28071,N_27716,N_27844);
xnor U28072 (N_28072,N_27514,N_27612);
nand U28073 (N_28073,N_27158,N_27084);
or U28074 (N_28074,N_27917,N_27424);
nor U28075 (N_28075,N_27743,N_27668);
and U28076 (N_28076,N_27654,N_27435);
or U28077 (N_28077,N_27445,N_27485);
nand U28078 (N_28078,N_27902,N_27939);
nand U28079 (N_28079,N_27952,N_27161);
xnor U28080 (N_28080,N_27783,N_27117);
nor U28081 (N_28081,N_27956,N_27710);
xnor U28082 (N_28082,N_27194,N_27151);
xor U28083 (N_28083,N_27443,N_27729);
or U28084 (N_28084,N_27769,N_27725);
nand U28085 (N_28085,N_27595,N_27327);
nor U28086 (N_28086,N_27096,N_27454);
or U28087 (N_28087,N_27295,N_27901);
nand U28088 (N_28088,N_27381,N_27636);
nor U28089 (N_28089,N_27275,N_27046);
xor U28090 (N_28090,N_27070,N_27184);
and U28091 (N_28091,N_27782,N_27197);
or U28092 (N_28092,N_27258,N_27254);
nor U28093 (N_28093,N_27322,N_27308);
nand U28094 (N_28094,N_27720,N_27911);
or U28095 (N_28095,N_27968,N_27427);
nor U28096 (N_28096,N_27220,N_27544);
nand U28097 (N_28097,N_27759,N_27450);
and U28098 (N_28098,N_27539,N_27386);
nor U28099 (N_28099,N_27207,N_27345);
nand U28100 (N_28100,N_27878,N_27828);
or U28101 (N_28101,N_27051,N_27248);
or U28102 (N_28102,N_27298,N_27586);
nand U28103 (N_28103,N_27392,N_27779);
nand U28104 (N_28104,N_27501,N_27887);
nand U28105 (N_28105,N_27066,N_27493);
or U28106 (N_28106,N_27524,N_27138);
and U28107 (N_28107,N_27188,N_27519);
xnor U28108 (N_28108,N_27768,N_27081);
nand U28109 (N_28109,N_27671,N_27757);
nand U28110 (N_28110,N_27579,N_27854);
and U28111 (N_28111,N_27414,N_27148);
or U28112 (N_28112,N_27954,N_27267);
and U28113 (N_28113,N_27655,N_27102);
or U28114 (N_28114,N_27719,N_27019);
nand U28115 (N_28115,N_27303,N_27522);
xnor U28116 (N_28116,N_27179,N_27767);
or U28117 (N_28117,N_27881,N_27397);
nand U28118 (N_28118,N_27344,N_27428);
xor U28119 (N_28119,N_27223,N_27817);
or U28120 (N_28120,N_27006,N_27717);
nor U28121 (N_28121,N_27732,N_27238);
nor U28122 (N_28122,N_27466,N_27469);
nand U28123 (N_28123,N_27742,N_27170);
and U28124 (N_28124,N_27677,N_27870);
nand U28125 (N_28125,N_27602,N_27401);
xnor U28126 (N_28126,N_27293,N_27461);
xor U28127 (N_28127,N_27052,N_27492);
nor U28128 (N_28128,N_27944,N_27306);
nor U28129 (N_28129,N_27784,N_27476);
nor U28130 (N_28130,N_27809,N_27420);
nor U28131 (N_28131,N_27080,N_27181);
or U28132 (N_28132,N_27154,N_27673);
nor U28133 (N_28133,N_27877,N_27702);
nor U28134 (N_28134,N_27389,N_27394);
nand U28135 (N_28135,N_27583,N_27965);
and U28136 (N_28136,N_27566,N_27935);
nor U28137 (N_28137,N_27032,N_27366);
or U28138 (N_28138,N_27936,N_27693);
nor U28139 (N_28139,N_27853,N_27640);
nand U28140 (N_28140,N_27943,N_27905);
and U28141 (N_28141,N_27611,N_27588);
nand U28142 (N_28142,N_27892,N_27119);
nor U28143 (N_28143,N_27650,N_27497);
nand U28144 (N_28144,N_27924,N_27972);
nor U28145 (N_28145,N_27276,N_27665);
nor U28146 (N_28146,N_27438,N_27970);
nor U28147 (N_28147,N_27621,N_27149);
or U28148 (N_28148,N_27418,N_27244);
nand U28149 (N_28149,N_27508,N_27708);
and U28150 (N_28150,N_27055,N_27569);
and U28151 (N_28151,N_27155,N_27811);
or U28152 (N_28152,N_27498,N_27407);
nand U28153 (N_28153,N_27173,N_27302);
nor U28154 (N_28154,N_27988,N_27380);
xor U28155 (N_28155,N_27209,N_27721);
and U28156 (N_28156,N_27239,N_27447);
xnor U28157 (N_28157,N_27568,N_27503);
and U28158 (N_28158,N_27009,N_27171);
nor U28159 (N_28159,N_27625,N_27177);
nor U28160 (N_28160,N_27663,N_27599);
nor U28161 (N_28161,N_27578,N_27962);
or U28162 (N_28162,N_27067,N_27013);
and U28163 (N_28163,N_27747,N_27487);
xor U28164 (N_28164,N_27150,N_27040);
nand U28165 (N_28165,N_27139,N_27263);
and U28166 (N_28166,N_27641,N_27875);
nor U28167 (N_28167,N_27292,N_27201);
or U28168 (N_28168,N_27806,N_27976);
nand U28169 (N_28169,N_27182,N_27191);
and U28170 (N_28170,N_27162,N_27228);
xor U28171 (N_28171,N_27004,N_27871);
xnor U28172 (N_28172,N_27646,N_27411);
and U28173 (N_28173,N_27700,N_27520);
nor U28174 (N_28174,N_27235,N_27741);
xnor U28175 (N_28175,N_27352,N_27876);
nor U28176 (N_28176,N_27127,N_27409);
nor U28177 (N_28177,N_27031,N_27603);
xnor U28178 (N_28178,N_27685,N_27795);
and U28179 (N_28179,N_27913,N_27587);
nor U28180 (N_28180,N_27313,N_27210);
nand U28181 (N_28181,N_27342,N_27359);
nand U28182 (N_28182,N_27580,N_27269);
or U28183 (N_28183,N_27028,N_27057);
and U28184 (N_28184,N_27477,N_27666);
and U28185 (N_28185,N_27442,N_27231);
and U28186 (N_28186,N_27279,N_27042);
xor U28187 (N_28187,N_27983,N_27071);
or U28188 (N_28188,N_27252,N_27793);
xnor U28189 (N_28189,N_27405,N_27996);
nand U28190 (N_28190,N_27460,N_27379);
and U28191 (N_28191,N_27124,N_27068);
nor U28192 (N_28192,N_27883,N_27513);
nand U28193 (N_28193,N_27550,N_27370);
nor U28194 (N_28194,N_27947,N_27816);
or U28195 (N_28195,N_27475,N_27452);
nor U28196 (N_28196,N_27778,N_27946);
and U28197 (N_28197,N_27548,N_27789);
nor U28198 (N_28198,N_27538,N_27562);
xor U28199 (N_28199,N_27977,N_27803);
xnor U28200 (N_28200,N_27994,N_27855);
nand U28201 (N_28201,N_27140,N_27349);
xnor U28202 (N_28202,N_27076,N_27299);
and U28203 (N_28203,N_27489,N_27601);
nor U28204 (N_28204,N_27391,N_27528);
xor U28205 (N_28205,N_27812,N_27865);
or U28206 (N_28206,N_27667,N_27914);
and U28207 (N_28207,N_27416,N_27973);
nor U28208 (N_28208,N_27257,N_27289);
xnor U28209 (N_28209,N_27200,N_27926);
and U28210 (N_28210,N_27997,N_27121);
nand U28211 (N_28211,N_27754,N_27288);
nand U28212 (N_28212,N_27711,N_27726);
xor U28213 (N_28213,N_27859,N_27846);
or U28214 (N_28214,N_27190,N_27908);
nand U28215 (N_28215,N_27111,N_27157);
or U28216 (N_28216,N_27561,N_27737);
xnor U28217 (N_28217,N_27385,N_27689);
xor U28218 (N_28218,N_27565,N_27606);
and U28219 (N_28219,N_27110,N_27502);
nand U28220 (N_28220,N_27047,N_27833);
xnor U28221 (N_28221,N_27331,N_27570);
nor U28222 (N_28222,N_27294,N_27126);
nand U28223 (N_28223,N_27961,N_27982);
and U28224 (N_28224,N_27086,N_27094);
nor U28225 (N_28225,N_27108,N_27589);
or U28226 (N_28226,N_27133,N_27540);
xor U28227 (N_28227,N_27496,N_27571);
and U28228 (N_28228,N_27393,N_27867);
nand U28229 (N_28229,N_27314,N_27056);
or U28230 (N_28230,N_27745,N_27202);
or U28231 (N_28231,N_27750,N_27384);
and U28232 (N_28232,N_27651,N_27290);
nor U28233 (N_28233,N_27796,N_27264);
xor U28234 (N_28234,N_27064,N_27249);
nand U28235 (N_28235,N_27075,N_27787);
nand U28236 (N_28236,N_27353,N_27425);
xor U28237 (N_28237,N_27978,N_27132);
or U28238 (N_28238,N_27764,N_27347);
nand U28239 (N_28239,N_27674,N_27462);
and U28240 (N_28240,N_27658,N_27164);
and U28241 (N_28241,N_27167,N_27776);
nor U28242 (N_28242,N_27214,N_27404);
and U28243 (N_28243,N_27593,N_27304);
and U28244 (N_28244,N_27889,N_27703);
nor U28245 (N_28245,N_27984,N_27575);
nor U28246 (N_28246,N_27199,N_27695);
nand U28247 (N_28247,N_27705,N_27728);
nor U28248 (N_28248,N_27053,N_27436);
and U28249 (N_28249,N_27770,N_27839);
xnor U28250 (N_28250,N_27296,N_27521);
nor U28251 (N_28251,N_27585,N_27408);
nor U28252 (N_28252,N_27858,N_27660);
and U28253 (N_28253,N_27820,N_27727);
nor U28254 (N_28254,N_27131,N_27421);
xnor U28255 (N_28255,N_27559,N_27687);
nand U28256 (N_28256,N_27390,N_27465);
xnor U28257 (N_28257,N_27659,N_27361);
xnor U28258 (N_28258,N_27363,N_27169);
xnor U28259 (N_28259,N_27649,N_27862);
nand U28260 (N_28260,N_27628,N_27351);
nor U28261 (N_28261,N_27334,N_27567);
nand U28262 (N_28262,N_27860,N_27851);
nor U28263 (N_28263,N_27990,N_27050);
nor U28264 (N_28264,N_27642,N_27251);
xnor U28265 (N_28265,N_27712,N_27144);
nand U28266 (N_28266,N_27265,N_27781);
xnor U28267 (N_28267,N_27330,N_27841);
and U28268 (N_28268,N_27744,N_27886);
nand U28269 (N_28269,N_27546,N_27791);
or U28270 (N_28270,N_27724,N_27805);
or U28271 (N_28271,N_27335,N_27011);
and U28272 (N_28272,N_27657,N_27661);
nor U28273 (N_28273,N_27270,N_27172);
and U28274 (N_28274,N_27906,N_27063);
xnor U28275 (N_28275,N_27213,N_27843);
nand U28276 (N_28276,N_27535,N_27160);
xnor U28277 (N_28277,N_27802,N_27874);
nand U28278 (N_28278,N_27594,N_27310);
nand U28279 (N_28279,N_27564,N_27560);
xnor U28280 (N_28280,N_27021,N_27683);
nor U28281 (N_28281,N_27099,N_27518);
and U28282 (N_28282,N_27061,N_27038);
nand U28283 (N_28283,N_27396,N_27014);
xnor U28284 (N_28284,N_27950,N_27760);
or U28285 (N_28285,N_27992,N_27444);
or U28286 (N_28286,N_27165,N_27891);
nand U28287 (N_28287,N_27557,N_27533);
nor U28288 (N_28288,N_27079,N_27631);
nor U28289 (N_28289,N_27643,N_27266);
nand U28290 (N_28290,N_27626,N_27364);
and U28291 (N_28291,N_27922,N_27035);
nand U28292 (N_28292,N_27491,N_27319);
or U28293 (N_28293,N_27446,N_27919);
nand U28294 (N_28294,N_27756,N_27375);
nand U28295 (N_28295,N_27797,N_27955);
xor U28296 (N_28296,N_27790,N_27339);
or U28297 (N_28297,N_27822,N_27937);
and U28298 (N_28298,N_27838,N_27899);
and U28299 (N_28299,N_27000,N_27555);
xnor U28300 (N_28300,N_27995,N_27958);
nor U28301 (N_28301,N_27437,N_27065);
nor U28302 (N_28302,N_27921,N_27316);
xnor U28303 (N_28303,N_27532,N_27430);
nand U28304 (N_28304,N_27592,N_27525);
nand U28305 (N_28305,N_27174,N_27753);
nor U28306 (N_28306,N_27340,N_27692);
nor U28307 (N_28307,N_27483,N_27981);
nor U28308 (N_28308,N_27694,N_27176);
or U28309 (N_28309,N_27069,N_27993);
xor U28310 (N_28310,N_27240,N_27137);
or U28311 (N_28311,N_27849,N_27618);
nor U28312 (N_28312,N_27185,N_27285);
nand U28313 (N_28313,N_27073,N_27054);
and U28314 (N_28314,N_27880,N_27527);
or U28315 (N_28315,N_27309,N_27488);
xor U28316 (N_28316,N_27431,N_27365);
nor U28317 (N_28317,N_27966,N_27798);
nand U28318 (N_28318,N_27918,N_27940);
or U28319 (N_28319,N_27025,N_27909);
and U28320 (N_28320,N_27852,N_27163);
or U28321 (N_28321,N_27857,N_27842);
or U28322 (N_28322,N_27423,N_27688);
nor U28323 (N_28323,N_27082,N_27348);
nand U28324 (N_28324,N_27704,N_27474);
or U28325 (N_28325,N_27402,N_27261);
or U28326 (N_28326,N_27931,N_27399);
xor U28327 (N_28327,N_27536,N_27135);
nand U28328 (N_28328,N_27624,N_27077);
nor U28329 (N_28329,N_27623,N_27060);
nor U28330 (N_28330,N_27632,N_27274);
xor U28331 (N_28331,N_27114,N_27554);
nand U28332 (N_28332,N_27957,N_27558);
xnor U28333 (N_28333,N_27297,N_27792);
xor U28334 (N_28334,N_27748,N_27403);
and U28335 (N_28335,N_27229,N_27036);
nand U28336 (N_28336,N_27869,N_27932);
nand U28337 (N_28337,N_27246,N_27429);
xor U28338 (N_28338,N_27998,N_27884);
and U28339 (N_28339,N_27440,N_27175);
nand U28340 (N_28340,N_27346,N_27617);
or U28341 (N_28341,N_27136,N_27152);
xnor U28342 (N_28342,N_27925,N_27368);
and U28343 (N_28343,N_27387,N_27622);
or U28344 (N_28344,N_27738,N_27241);
and U28345 (N_28345,N_27664,N_27225);
xor U28346 (N_28346,N_27286,N_27788);
and U28347 (N_28347,N_27813,N_27186);
or U28348 (N_28348,N_27092,N_27101);
and U28349 (N_28349,N_27629,N_27044);
or U28350 (N_28350,N_27458,N_27814);
nand U28351 (N_28351,N_27807,N_27490);
and U28352 (N_28352,N_27930,N_27109);
nor U28353 (N_28353,N_27680,N_27236);
and U28354 (N_28354,N_27336,N_27801);
xnor U28355 (N_28355,N_27037,N_27283);
and U28356 (N_28356,N_27305,N_27312);
and U28357 (N_28357,N_27633,N_27432);
nand U28358 (N_28358,N_27328,N_27242);
and U28359 (N_28359,N_27923,N_27676);
xor U28360 (N_28360,N_27915,N_27464);
nor U28361 (N_28361,N_27329,N_27321);
or U28362 (N_28362,N_27644,N_27696);
nand U28363 (N_28363,N_27382,N_27341);
and U28364 (N_28364,N_27549,N_27834);
nand U28365 (N_28365,N_27072,N_27377);
and U28366 (N_28366,N_27986,N_27217);
or U28367 (N_28367,N_27682,N_27472);
or U28368 (N_28368,N_27500,N_27215);
or U28369 (N_28369,N_27417,N_27731);
xor U28370 (N_28370,N_27142,N_27608);
or U28371 (N_28371,N_27088,N_27690);
xor U28372 (N_28372,N_27504,N_27227);
nand U28373 (N_28373,N_27463,N_27669);
or U28374 (N_28374,N_27468,N_27991);
or U28375 (N_28375,N_27933,N_27530);
or U28376 (N_28376,N_27291,N_27459);
and U28377 (N_28377,N_27577,N_27627);
nor U28378 (N_28378,N_27613,N_27735);
and U28379 (N_28379,N_27574,N_27116);
or U28380 (N_28380,N_27698,N_27470);
nand U28381 (N_28381,N_27457,N_27218);
or U28382 (N_28382,N_27211,N_27619);
nor U28383 (N_28383,N_27016,N_27395);
xnor U28384 (N_28384,N_27448,N_27888);
nor U28385 (N_28385,N_27630,N_27523);
and U28386 (N_28386,N_27373,N_27900);
and U28387 (N_28387,N_27938,N_27045);
and U28388 (N_28388,N_27730,N_27010);
nand U28389 (N_28389,N_27635,N_27799);
xor U28390 (N_28390,N_27005,N_27681);
or U28391 (N_28391,N_27545,N_27062);
or U28392 (N_28392,N_27449,N_27903);
nand U28393 (N_28393,N_27505,N_27960);
nor U28394 (N_28394,N_27192,N_27333);
nand U28395 (N_28395,N_27216,N_27679);
xnor U28396 (N_28396,N_27752,N_27357);
xor U28397 (N_28397,N_27439,N_27774);
or U28398 (N_28398,N_27195,N_27129);
nand U28399 (N_28399,N_27125,N_27325);
and U28400 (N_28400,N_27369,N_27825);
nand U28401 (N_28401,N_27311,N_27714);
nor U28402 (N_28402,N_27495,N_27722);
or U28403 (N_28403,N_27916,N_27224);
nand U28404 (N_28404,N_27734,N_27253);
nor U28405 (N_28405,N_27271,N_27582);
xnor U28406 (N_28406,N_27971,N_27074);
nand U28407 (N_28407,N_27910,N_27848);
nand U28408 (N_28408,N_27486,N_27509);
xnor U28409 (N_28409,N_27206,N_27230);
nor U28410 (N_28410,N_27653,N_27453);
xnor U28411 (N_28411,N_27078,N_27039);
nor U28412 (N_28412,N_27237,N_27315);
nand U28413 (N_28413,N_27301,N_27058);
or U28414 (N_28414,N_27785,N_27856);
xor U28415 (N_28415,N_27307,N_27620);
nor U28416 (N_28416,N_27034,N_27953);
or U28417 (N_28417,N_27189,N_27017);
or U28418 (N_28418,N_27159,N_27219);
nand U28419 (N_28419,N_27810,N_27885);
and U28420 (N_28420,N_27128,N_27147);
nor U28421 (N_28421,N_27645,N_27736);
and U28422 (N_28422,N_27675,N_27882);
or U28423 (N_28423,N_27948,N_27048);
xnor U28424 (N_28424,N_27412,N_27607);
nor U28425 (N_28425,N_27701,N_27015);
xor U28426 (N_28426,N_27083,N_27847);
and U28427 (N_28427,N_27027,N_27243);
or U28428 (N_28428,N_27234,N_27614);
xnor U28429 (N_28429,N_27819,N_27097);
or U28430 (N_28430,N_27765,N_27374);
or U28431 (N_28431,N_27531,N_27277);
and U28432 (N_28432,N_27553,N_27208);
xnor U28433 (N_28433,N_27758,N_27105);
xor U28434 (N_28434,N_27547,N_27022);
xnor U28435 (N_28435,N_27146,N_27247);
nand U28436 (N_28436,N_27001,N_27773);
nand U28437 (N_28437,N_27007,N_27749);
and U28438 (N_28438,N_27033,N_27115);
nor U28439 (N_28439,N_27153,N_27318);
and U28440 (N_28440,N_27030,N_27866);
and U28441 (N_28441,N_27388,N_27104);
and U28442 (N_28442,N_27945,N_27455);
nand U28443 (N_28443,N_27699,N_27551);
and U28444 (N_28444,N_27203,N_27868);
nor U28445 (N_28445,N_27268,N_27320);
nor U28446 (N_28446,N_27829,N_27967);
nand U28447 (N_28447,N_27920,N_27845);
or U28448 (N_28448,N_27707,N_27441);
nor U28449 (N_28449,N_27821,N_27026);
nand U28450 (N_28450,N_27800,N_27656);
nor U28451 (N_28451,N_27350,N_27723);
nand U28452 (N_28452,N_27280,N_27089);
or U28453 (N_28453,N_27824,N_27512);
xor U28454 (N_28454,N_27118,N_27332);
nor U28455 (N_28455,N_27763,N_27098);
and U28456 (N_28456,N_27794,N_27979);
xor U28457 (N_28457,N_27378,N_27106);
and U28458 (N_28458,N_27250,N_27481);
xnor U28459 (N_28459,N_27541,N_27980);
xnor U28460 (N_28460,N_27494,N_27563);
or U28461 (N_28461,N_27832,N_27670);
nor U28462 (N_28462,N_27024,N_27023);
and U28463 (N_28463,N_27652,N_27008);
nor U28464 (N_28464,N_27196,N_27012);
xor U28465 (N_28465,N_27818,N_27894);
nor U28466 (N_28466,N_27863,N_27713);
xnor U28467 (N_28467,N_27260,N_27686);
nor U28468 (N_28468,N_27145,N_27482);
nor U28469 (N_28469,N_27434,N_27112);
nor U28470 (N_28470,N_27529,N_27590);
nand U28471 (N_28471,N_27002,N_27122);
nand U28472 (N_28472,N_27912,N_27256);
and U28473 (N_28473,N_27771,N_27534);
or U28474 (N_28474,N_27337,N_27604);
nand U28475 (N_28475,N_27609,N_27987);
nor U28476 (N_28476,N_27963,N_27739);
nor U28477 (N_28477,N_27183,N_27282);
and U28478 (N_28478,N_27400,N_27376);
nor U28479 (N_28479,N_27637,N_27506);
and U28480 (N_28480,N_27772,N_27691);
nand U28481 (N_28481,N_27515,N_27942);
nand U28482 (N_28482,N_27356,N_27662);
nor U28483 (N_28483,N_27706,N_27927);
nand U28484 (N_28484,N_27415,N_27020);
or U28485 (N_28485,N_27272,N_27091);
or U28486 (N_28486,N_27904,N_27672);
nand U28487 (N_28487,N_27526,N_27433);
or U28488 (N_28488,N_27103,N_27831);
or U28489 (N_28489,N_27354,N_27746);
nor U28490 (N_28490,N_27873,N_27360);
nand U28491 (N_28491,N_27245,N_27358);
xnor U28492 (N_28492,N_27255,N_27815);
or U28493 (N_28493,N_27090,N_27471);
and U28494 (N_28494,N_27605,N_27516);
nor U28495 (N_28495,N_27419,N_27355);
nor U28496 (N_28496,N_27969,N_27999);
nand U28497 (N_28497,N_27123,N_27639);
and U28498 (N_28498,N_27895,N_27678);
xor U28499 (N_28499,N_27041,N_27985);
xnor U28500 (N_28500,N_27964,N_27603);
and U28501 (N_28501,N_27605,N_27293);
nand U28502 (N_28502,N_27231,N_27210);
nor U28503 (N_28503,N_27762,N_27052);
and U28504 (N_28504,N_27124,N_27965);
nand U28505 (N_28505,N_27783,N_27459);
nand U28506 (N_28506,N_27267,N_27968);
and U28507 (N_28507,N_27828,N_27794);
xor U28508 (N_28508,N_27747,N_27781);
or U28509 (N_28509,N_27749,N_27329);
and U28510 (N_28510,N_27654,N_27824);
xnor U28511 (N_28511,N_27564,N_27773);
and U28512 (N_28512,N_27972,N_27102);
nand U28513 (N_28513,N_27110,N_27888);
nand U28514 (N_28514,N_27834,N_27886);
and U28515 (N_28515,N_27133,N_27682);
nand U28516 (N_28516,N_27675,N_27614);
nor U28517 (N_28517,N_27512,N_27267);
or U28518 (N_28518,N_27691,N_27256);
xor U28519 (N_28519,N_27392,N_27981);
xor U28520 (N_28520,N_27445,N_27215);
and U28521 (N_28521,N_27671,N_27557);
nand U28522 (N_28522,N_27230,N_27382);
nor U28523 (N_28523,N_27638,N_27856);
and U28524 (N_28524,N_27024,N_27783);
or U28525 (N_28525,N_27213,N_27470);
and U28526 (N_28526,N_27277,N_27648);
and U28527 (N_28527,N_27434,N_27082);
xnor U28528 (N_28528,N_27945,N_27391);
or U28529 (N_28529,N_27614,N_27601);
nor U28530 (N_28530,N_27175,N_27645);
and U28531 (N_28531,N_27947,N_27053);
and U28532 (N_28532,N_27895,N_27890);
nand U28533 (N_28533,N_27443,N_27368);
xnor U28534 (N_28534,N_27291,N_27806);
nor U28535 (N_28535,N_27555,N_27989);
or U28536 (N_28536,N_27402,N_27052);
or U28537 (N_28537,N_27911,N_27769);
or U28538 (N_28538,N_27435,N_27605);
or U28539 (N_28539,N_27882,N_27773);
nor U28540 (N_28540,N_27850,N_27825);
or U28541 (N_28541,N_27476,N_27980);
nand U28542 (N_28542,N_27897,N_27011);
nand U28543 (N_28543,N_27400,N_27395);
nor U28544 (N_28544,N_27340,N_27558);
and U28545 (N_28545,N_27800,N_27704);
or U28546 (N_28546,N_27113,N_27662);
xor U28547 (N_28547,N_27246,N_27321);
xor U28548 (N_28548,N_27633,N_27449);
and U28549 (N_28549,N_27401,N_27022);
nand U28550 (N_28550,N_27583,N_27100);
nor U28551 (N_28551,N_27209,N_27575);
xnor U28552 (N_28552,N_27453,N_27580);
nor U28553 (N_28553,N_27674,N_27066);
xnor U28554 (N_28554,N_27768,N_27436);
nand U28555 (N_28555,N_27100,N_27908);
xnor U28556 (N_28556,N_27375,N_27846);
nand U28557 (N_28557,N_27055,N_27197);
or U28558 (N_28558,N_27042,N_27315);
or U28559 (N_28559,N_27724,N_27124);
or U28560 (N_28560,N_27995,N_27504);
xor U28561 (N_28561,N_27254,N_27311);
and U28562 (N_28562,N_27453,N_27890);
nand U28563 (N_28563,N_27579,N_27515);
nand U28564 (N_28564,N_27781,N_27212);
and U28565 (N_28565,N_27190,N_27556);
nand U28566 (N_28566,N_27578,N_27580);
nor U28567 (N_28567,N_27558,N_27306);
nor U28568 (N_28568,N_27136,N_27833);
xnor U28569 (N_28569,N_27103,N_27482);
and U28570 (N_28570,N_27867,N_27151);
and U28571 (N_28571,N_27066,N_27644);
xnor U28572 (N_28572,N_27628,N_27877);
xor U28573 (N_28573,N_27056,N_27566);
or U28574 (N_28574,N_27840,N_27816);
nor U28575 (N_28575,N_27554,N_27484);
and U28576 (N_28576,N_27641,N_27346);
nor U28577 (N_28577,N_27144,N_27348);
or U28578 (N_28578,N_27506,N_27611);
nand U28579 (N_28579,N_27122,N_27915);
xor U28580 (N_28580,N_27320,N_27903);
and U28581 (N_28581,N_27080,N_27247);
nand U28582 (N_28582,N_27154,N_27603);
nor U28583 (N_28583,N_27629,N_27632);
xor U28584 (N_28584,N_27587,N_27957);
nor U28585 (N_28585,N_27176,N_27755);
nor U28586 (N_28586,N_27358,N_27429);
xnor U28587 (N_28587,N_27137,N_27870);
nand U28588 (N_28588,N_27894,N_27285);
or U28589 (N_28589,N_27524,N_27145);
nand U28590 (N_28590,N_27693,N_27565);
nor U28591 (N_28591,N_27437,N_27830);
or U28592 (N_28592,N_27589,N_27186);
nor U28593 (N_28593,N_27195,N_27663);
nor U28594 (N_28594,N_27700,N_27541);
or U28595 (N_28595,N_27846,N_27455);
nand U28596 (N_28596,N_27805,N_27368);
and U28597 (N_28597,N_27115,N_27098);
nor U28598 (N_28598,N_27403,N_27361);
or U28599 (N_28599,N_27689,N_27652);
nor U28600 (N_28600,N_27038,N_27353);
nand U28601 (N_28601,N_27465,N_27927);
xor U28602 (N_28602,N_27440,N_27137);
xor U28603 (N_28603,N_27934,N_27783);
nand U28604 (N_28604,N_27435,N_27249);
xor U28605 (N_28605,N_27814,N_27120);
or U28606 (N_28606,N_27761,N_27203);
or U28607 (N_28607,N_27179,N_27077);
or U28608 (N_28608,N_27353,N_27099);
or U28609 (N_28609,N_27363,N_27509);
and U28610 (N_28610,N_27132,N_27816);
xnor U28611 (N_28611,N_27031,N_27691);
or U28612 (N_28612,N_27441,N_27815);
nand U28613 (N_28613,N_27931,N_27594);
nor U28614 (N_28614,N_27029,N_27268);
nor U28615 (N_28615,N_27637,N_27910);
and U28616 (N_28616,N_27740,N_27423);
xor U28617 (N_28617,N_27812,N_27937);
nor U28618 (N_28618,N_27113,N_27990);
or U28619 (N_28619,N_27209,N_27785);
xnor U28620 (N_28620,N_27402,N_27149);
nand U28621 (N_28621,N_27213,N_27629);
or U28622 (N_28622,N_27448,N_27682);
or U28623 (N_28623,N_27545,N_27112);
xor U28624 (N_28624,N_27581,N_27140);
and U28625 (N_28625,N_27176,N_27065);
or U28626 (N_28626,N_27803,N_27656);
and U28627 (N_28627,N_27918,N_27119);
nor U28628 (N_28628,N_27435,N_27149);
xor U28629 (N_28629,N_27169,N_27514);
or U28630 (N_28630,N_27269,N_27665);
nor U28631 (N_28631,N_27411,N_27500);
nand U28632 (N_28632,N_27472,N_27713);
and U28633 (N_28633,N_27234,N_27871);
nor U28634 (N_28634,N_27560,N_27828);
xor U28635 (N_28635,N_27818,N_27988);
xor U28636 (N_28636,N_27435,N_27970);
nor U28637 (N_28637,N_27802,N_27862);
xnor U28638 (N_28638,N_27814,N_27613);
xnor U28639 (N_28639,N_27592,N_27687);
xor U28640 (N_28640,N_27037,N_27671);
or U28641 (N_28641,N_27004,N_27904);
nor U28642 (N_28642,N_27914,N_27266);
or U28643 (N_28643,N_27248,N_27564);
xnor U28644 (N_28644,N_27273,N_27431);
xnor U28645 (N_28645,N_27989,N_27210);
nand U28646 (N_28646,N_27133,N_27843);
nor U28647 (N_28647,N_27814,N_27019);
nand U28648 (N_28648,N_27148,N_27328);
nor U28649 (N_28649,N_27203,N_27529);
and U28650 (N_28650,N_27570,N_27481);
nand U28651 (N_28651,N_27536,N_27519);
and U28652 (N_28652,N_27922,N_27040);
or U28653 (N_28653,N_27251,N_27706);
nor U28654 (N_28654,N_27560,N_27837);
xnor U28655 (N_28655,N_27746,N_27822);
and U28656 (N_28656,N_27159,N_27807);
nand U28657 (N_28657,N_27142,N_27038);
nor U28658 (N_28658,N_27360,N_27472);
and U28659 (N_28659,N_27614,N_27011);
nor U28660 (N_28660,N_27383,N_27320);
and U28661 (N_28661,N_27386,N_27858);
and U28662 (N_28662,N_27092,N_27659);
or U28663 (N_28663,N_27274,N_27262);
and U28664 (N_28664,N_27353,N_27675);
xor U28665 (N_28665,N_27501,N_27951);
nand U28666 (N_28666,N_27254,N_27936);
and U28667 (N_28667,N_27642,N_27584);
nor U28668 (N_28668,N_27973,N_27002);
xnor U28669 (N_28669,N_27603,N_27433);
and U28670 (N_28670,N_27750,N_27581);
and U28671 (N_28671,N_27832,N_27546);
or U28672 (N_28672,N_27320,N_27805);
xor U28673 (N_28673,N_27941,N_27795);
or U28674 (N_28674,N_27070,N_27422);
nand U28675 (N_28675,N_27820,N_27462);
nor U28676 (N_28676,N_27959,N_27222);
nand U28677 (N_28677,N_27157,N_27401);
nand U28678 (N_28678,N_27402,N_27602);
or U28679 (N_28679,N_27163,N_27314);
nand U28680 (N_28680,N_27055,N_27785);
nor U28681 (N_28681,N_27098,N_27934);
xor U28682 (N_28682,N_27111,N_27016);
or U28683 (N_28683,N_27407,N_27758);
xor U28684 (N_28684,N_27614,N_27174);
nand U28685 (N_28685,N_27948,N_27105);
nor U28686 (N_28686,N_27764,N_27277);
and U28687 (N_28687,N_27255,N_27680);
and U28688 (N_28688,N_27739,N_27090);
nor U28689 (N_28689,N_27747,N_27832);
nor U28690 (N_28690,N_27828,N_27335);
and U28691 (N_28691,N_27911,N_27789);
nand U28692 (N_28692,N_27761,N_27273);
and U28693 (N_28693,N_27969,N_27317);
or U28694 (N_28694,N_27002,N_27112);
nor U28695 (N_28695,N_27120,N_27502);
or U28696 (N_28696,N_27281,N_27712);
and U28697 (N_28697,N_27702,N_27281);
or U28698 (N_28698,N_27879,N_27883);
xnor U28699 (N_28699,N_27949,N_27258);
nand U28700 (N_28700,N_27324,N_27099);
xor U28701 (N_28701,N_27407,N_27466);
or U28702 (N_28702,N_27291,N_27813);
xnor U28703 (N_28703,N_27436,N_27423);
xor U28704 (N_28704,N_27521,N_27412);
and U28705 (N_28705,N_27489,N_27311);
or U28706 (N_28706,N_27164,N_27412);
and U28707 (N_28707,N_27329,N_27653);
or U28708 (N_28708,N_27296,N_27205);
xor U28709 (N_28709,N_27065,N_27240);
nor U28710 (N_28710,N_27980,N_27878);
and U28711 (N_28711,N_27692,N_27491);
nor U28712 (N_28712,N_27126,N_27019);
and U28713 (N_28713,N_27325,N_27035);
nand U28714 (N_28714,N_27036,N_27441);
and U28715 (N_28715,N_27818,N_27955);
nand U28716 (N_28716,N_27604,N_27815);
or U28717 (N_28717,N_27410,N_27280);
and U28718 (N_28718,N_27476,N_27278);
xor U28719 (N_28719,N_27764,N_27815);
xnor U28720 (N_28720,N_27129,N_27615);
nand U28721 (N_28721,N_27166,N_27315);
xnor U28722 (N_28722,N_27264,N_27456);
nand U28723 (N_28723,N_27360,N_27435);
xor U28724 (N_28724,N_27295,N_27783);
and U28725 (N_28725,N_27286,N_27844);
nand U28726 (N_28726,N_27694,N_27728);
nor U28727 (N_28727,N_27255,N_27835);
nor U28728 (N_28728,N_27664,N_27434);
xnor U28729 (N_28729,N_27699,N_27956);
or U28730 (N_28730,N_27501,N_27737);
or U28731 (N_28731,N_27372,N_27317);
and U28732 (N_28732,N_27072,N_27566);
xor U28733 (N_28733,N_27904,N_27659);
nand U28734 (N_28734,N_27489,N_27935);
nand U28735 (N_28735,N_27244,N_27523);
nor U28736 (N_28736,N_27521,N_27865);
nor U28737 (N_28737,N_27560,N_27422);
or U28738 (N_28738,N_27939,N_27599);
xor U28739 (N_28739,N_27126,N_27622);
nor U28740 (N_28740,N_27674,N_27409);
nor U28741 (N_28741,N_27031,N_27899);
xor U28742 (N_28742,N_27133,N_27490);
xnor U28743 (N_28743,N_27499,N_27297);
nand U28744 (N_28744,N_27544,N_27674);
nand U28745 (N_28745,N_27867,N_27301);
and U28746 (N_28746,N_27838,N_27359);
and U28747 (N_28747,N_27540,N_27697);
nor U28748 (N_28748,N_27470,N_27279);
xnor U28749 (N_28749,N_27017,N_27963);
or U28750 (N_28750,N_27019,N_27576);
or U28751 (N_28751,N_27086,N_27548);
and U28752 (N_28752,N_27712,N_27049);
nor U28753 (N_28753,N_27344,N_27210);
xor U28754 (N_28754,N_27247,N_27253);
and U28755 (N_28755,N_27570,N_27571);
nand U28756 (N_28756,N_27159,N_27736);
and U28757 (N_28757,N_27436,N_27682);
nor U28758 (N_28758,N_27699,N_27279);
and U28759 (N_28759,N_27529,N_27547);
nand U28760 (N_28760,N_27231,N_27953);
or U28761 (N_28761,N_27117,N_27303);
or U28762 (N_28762,N_27939,N_27733);
and U28763 (N_28763,N_27470,N_27282);
or U28764 (N_28764,N_27287,N_27547);
nand U28765 (N_28765,N_27914,N_27220);
nand U28766 (N_28766,N_27098,N_27859);
nand U28767 (N_28767,N_27558,N_27154);
nor U28768 (N_28768,N_27020,N_27609);
or U28769 (N_28769,N_27591,N_27727);
xor U28770 (N_28770,N_27460,N_27790);
or U28771 (N_28771,N_27890,N_27488);
xnor U28772 (N_28772,N_27511,N_27253);
nand U28773 (N_28773,N_27711,N_27329);
and U28774 (N_28774,N_27304,N_27590);
nor U28775 (N_28775,N_27973,N_27408);
xor U28776 (N_28776,N_27343,N_27576);
or U28777 (N_28777,N_27824,N_27350);
nand U28778 (N_28778,N_27243,N_27214);
nand U28779 (N_28779,N_27943,N_27222);
or U28780 (N_28780,N_27060,N_27684);
nor U28781 (N_28781,N_27649,N_27571);
xor U28782 (N_28782,N_27964,N_27113);
xor U28783 (N_28783,N_27376,N_27312);
and U28784 (N_28784,N_27094,N_27031);
nor U28785 (N_28785,N_27312,N_27978);
and U28786 (N_28786,N_27554,N_27089);
xnor U28787 (N_28787,N_27815,N_27990);
or U28788 (N_28788,N_27928,N_27891);
xnor U28789 (N_28789,N_27124,N_27264);
nor U28790 (N_28790,N_27982,N_27668);
xnor U28791 (N_28791,N_27077,N_27741);
nand U28792 (N_28792,N_27460,N_27366);
xor U28793 (N_28793,N_27258,N_27858);
or U28794 (N_28794,N_27779,N_27490);
nor U28795 (N_28795,N_27309,N_27341);
xor U28796 (N_28796,N_27439,N_27234);
and U28797 (N_28797,N_27936,N_27340);
nor U28798 (N_28798,N_27171,N_27339);
nand U28799 (N_28799,N_27559,N_27547);
nand U28800 (N_28800,N_27671,N_27776);
xnor U28801 (N_28801,N_27225,N_27675);
nor U28802 (N_28802,N_27582,N_27224);
nand U28803 (N_28803,N_27168,N_27368);
nor U28804 (N_28804,N_27880,N_27336);
xor U28805 (N_28805,N_27638,N_27975);
xor U28806 (N_28806,N_27723,N_27525);
and U28807 (N_28807,N_27415,N_27593);
and U28808 (N_28808,N_27919,N_27623);
xnor U28809 (N_28809,N_27491,N_27437);
nand U28810 (N_28810,N_27920,N_27341);
nor U28811 (N_28811,N_27532,N_27745);
nor U28812 (N_28812,N_27600,N_27389);
nor U28813 (N_28813,N_27740,N_27777);
nor U28814 (N_28814,N_27153,N_27915);
or U28815 (N_28815,N_27873,N_27917);
and U28816 (N_28816,N_27189,N_27254);
nor U28817 (N_28817,N_27227,N_27119);
or U28818 (N_28818,N_27402,N_27396);
nor U28819 (N_28819,N_27245,N_27674);
nand U28820 (N_28820,N_27721,N_27160);
nor U28821 (N_28821,N_27777,N_27618);
or U28822 (N_28822,N_27209,N_27499);
nor U28823 (N_28823,N_27746,N_27929);
xor U28824 (N_28824,N_27803,N_27612);
nand U28825 (N_28825,N_27192,N_27431);
or U28826 (N_28826,N_27551,N_27358);
xor U28827 (N_28827,N_27450,N_27806);
and U28828 (N_28828,N_27281,N_27263);
and U28829 (N_28829,N_27373,N_27960);
nand U28830 (N_28830,N_27810,N_27503);
xnor U28831 (N_28831,N_27779,N_27522);
or U28832 (N_28832,N_27042,N_27746);
nand U28833 (N_28833,N_27806,N_27560);
nand U28834 (N_28834,N_27196,N_27729);
xnor U28835 (N_28835,N_27417,N_27255);
or U28836 (N_28836,N_27230,N_27058);
xor U28837 (N_28837,N_27298,N_27209);
or U28838 (N_28838,N_27614,N_27623);
xor U28839 (N_28839,N_27064,N_27059);
nor U28840 (N_28840,N_27419,N_27892);
and U28841 (N_28841,N_27273,N_27134);
nor U28842 (N_28842,N_27824,N_27234);
xor U28843 (N_28843,N_27681,N_27579);
xnor U28844 (N_28844,N_27292,N_27099);
nor U28845 (N_28845,N_27662,N_27326);
xnor U28846 (N_28846,N_27217,N_27185);
nor U28847 (N_28847,N_27467,N_27496);
xor U28848 (N_28848,N_27045,N_27813);
nand U28849 (N_28849,N_27123,N_27438);
and U28850 (N_28850,N_27604,N_27450);
nor U28851 (N_28851,N_27194,N_27913);
xnor U28852 (N_28852,N_27164,N_27746);
nor U28853 (N_28853,N_27597,N_27843);
nor U28854 (N_28854,N_27657,N_27481);
nor U28855 (N_28855,N_27920,N_27175);
nand U28856 (N_28856,N_27456,N_27609);
nand U28857 (N_28857,N_27203,N_27618);
or U28858 (N_28858,N_27063,N_27195);
and U28859 (N_28859,N_27329,N_27441);
nand U28860 (N_28860,N_27934,N_27509);
and U28861 (N_28861,N_27912,N_27269);
and U28862 (N_28862,N_27022,N_27828);
xnor U28863 (N_28863,N_27042,N_27806);
xor U28864 (N_28864,N_27985,N_27109);
or U28865 (N_28865,N_27221,N_27818);
nand U28866 (N_28866,N_27117,N_27987);
nor U28867 (N_28867,N_27280,N_27362);
xor U28868 (N_28868,N_27889,N_27575);
nor U28869 (N_28869,N_27915,N_27006);
and U28870 (N_28870,N_27478,N_27221);
or U28871 (N_28871,N_27337,N_27672);
nand U28872 (N_28872,N_27999,N_27661);
nand U28873 (N_28873,N_27488,N_27793);
or U28874 (N_28874,N_27817,N_27200);
nor U28875 (N_28875,N_27721,N_27620);
or U28876 (N_28876,N_27879,N_27147);
xnor U28877 (N_28877,N_27239,N_27225);
or U28878 (N_28878,N_27038,N_27496);
nand U28879 (N_28879,N_27365,N_27110);
or U28880 (N_28880,N_27753,N_27589);
nor U28881 (N_28881,N_27131,N_27124);
and U28882 (N_28882,N_27385,N_27344);
nand U28883 (N_28883,N_27138,N_27047);
nand U28884 (N_28884,N_27857,N_27206);
or U28885 (N_28885,N_27073,N_27234);
nor U28886 (N_28886,N_27824,N_27953);
or U28887 (N_28887,N_27639,N_27260);
or U28888 (N_28888,N_27180,N_27548);
nand U28889 (N_28889,N_27411,N_27164);
nand U28890 (N_28890,N_27378,N_27743);
nor U28891 (N_28891,N_27937,N_27413);
nand U28892 (N_28892,N_27755,N_27507);
or U28893 (N_28893,N_27629,N_27310);
or U28894 (N_28894,N_27221,N_27128);
and U28895 (N_28895,N_27947,N_27678);
nor U28896 (N_28896,N_27102,N_27641);
nor U28897 (N_28897,N_27389,N_27897);
and U28898 (N_28898,N_27581,N_27552);
xor U28899 (N_28899,N_27104,N_27428);
nor U28900 (N_28900,N_27819,N_27456);
nand U28901 (N_28901,N_27596,N_27033);
or U28902 (N_28902,N_27810,N_27055);
or U28903 (N_28903,N_27237,N_27045);
xnor U28904 (N_28904,N_27076,N_27612);
and U28905 (N_28905,N_27232,N_27079);
nor U28906 (N_28906,N_27752,N_27941);
xor U28907 (N_28907,N_27907,N_27156);
nand U28908 (N_28908,N_27052,N_27235);
nor U28909 (N_28909,N_27955,N_27928);
xor U28910 (N_28910,N_27013,N_27557);
nor U28911 (N_28911,N_27891,N_27204);
or U28912 (N_28912,N_27364,N_27695);
nor U28913 (N_28913,N_27924,N_27809);
xnor U28914 (N_28914,N_27165,N_27954);
xnor U28915 (N_28915,N_27694,N_27316);
and U28916 (N_28916,N_27219,N_27679);
xnor U28917 (N_28917,N_27973,N_27409);
and U28918 (N_28918,N_27863,N_27187);
or U28919 (N_28919,N_27965,N_27175);
nor U28920 (N_28920,N_27377,N_27058);
and U28921 (N_28921,N_27587,N_27686);
nand U28922 (N_28922,N_27056,N_27173);
or U28923 (N_28923,N_27024,N_27959);
nor U28924 (N_28924,N_27583,N_27192);
and U28925 (N_28925,N_27691,N_27306);
xor U28926 (N_28926,N_27590,N_27279);
or U28927 (N_28927,N_27262,N_27599);
xor U28928 (N_28928,N_27626,N_27747);
nand U28929 (N_28929,N_27954,N_27527);
nand U28930 (N_28930,N_27654,N_27536);
nand U28931 (N_28931,N_27855,N_27692);
nor U28932 (N_28932,N_27035,N_27067);
or U28933 (N_28933,N_27524,N_27557);
nand U28934 (N_28934,N_27678,N_27989);
or U28935 (N_28935,N_27083,N_27937);
xnor U28936 (N_28936,N_27879,N_27952);
nand U28937 (N_28937,N_27263,N_27404);
nor U28938 (N_28938,N_27262,N_27661);
xnor U28939 (N_28939,N_27795,N_27896);
xnor U28940 (N_28940,N_27453,N_27848);
nor U28941 (N_28941,N_27895,N_27956);
nand U28942 (N_28942,N_27055,N_27177);
or U28943 (N_28943,N_27829,N_27081);
xor U28944 (N_28944,N_27774,N_27031);
xnor U28945 (N_28945,N_27565,N_27842);
nand U28946 (N_28946,N_27541,N_27505);
nand U28947 (N_28947,N_27054,N_27756);
and U28948 (N_28948,N_27474,N_27141);
nor U28949 (N_28949,N_27543,N_27564);
nor U28950 (N_28950,N_27938,N_27095);
or U28951 (N_28951,N_27256,N_27808);
nand U28952 (N_28952,N_27147,N_27283);
nand U28953 (N_28953,N_27812,N_27163);
or U28954 (N_28954,N_27068,N_27092);
and U28955 (N_28955,N_27955,N_27926);
xnor U28956 (N_28956,N_27500,N_27910);
nand U28957 (N_28957,N_27894,N_27154);
or U28958 (N_28958,N_27626,N_27351);
and U28959 (N_28959,N_27888,N_27393);
nand U28960 (N_28960,N_27379,N_27633);
nand U28961 (N_28961,N_27872,N_27906);
nor U28962 (N_28962,N_27244,N_27387);
and U28963 (N_28963,N_27266,N_27238);
xnor U28964 (N_28964,N_27592,N_27524);
and U28965 (N_28965,N_27799,N_27113);
xor U28966 (N_28966,N_27450,N_27017);
and U28967 (N_28967,N_27489,N_27825);
and U28968 (N_28968,N_27196,N_27111);
or U28969 (N_28969,N_27394,N_27920);
nand U28970 (N_28970,N_27402,N_27010);
nand U28971 (N_28971,N_27369,N_27468);
nor U28972 (N_28972,N_27897,N_27819);
nor U28973 (N_28973,N_27807,N_27290);
nor U28974 (N_28974,N_27494,N_27013);
or U28975 (N_28975,N_27387,N_27482);
nor U28976 (N_28976,N_27753,N_27785);
nor U28977 (N_28977,N_27726,N_27725);
and U28978 (N_28978,N_27716,N_27240);
and U28979 (N_28979,N_27616,N_27804);
or U28980 (N_28980,N_27338,N_27413);
nor U28981 (N_28981,N_27520,N_27596);
and U28982 (N_28982,N_27295,N_27205);
xor U28983 (N_28983,N_27228,N_27444);
xnor U28984 (N_28984,N_27762,N_27207);
xor U28985 (N_28985,N_27442,N_27557);
and U28986 (N_28986,N_27508,N_27383);
and U28987 (N_28987,N_27716,N_27477);
nand U28988 (N_28988,N_27183,N_27609);
xor U28989 (N_28989,N_27418,N_27921);
and U28990 (N_28990,N_27744,N_27180);
or U28991 (N_28991,N_27433,N_27107);
xnor U28992 (N_28992,N_27729,N_27486);
nand U28993 (N_28993,N_27215,N_27412);
and U28994 (N_28994,N_27094,N_27588);
or U28995 (N_28995,N_27523,N_27094);
nand U28996 (N_28996,N_27175,N_27345);
nand U28997 (N_28997,N_27664,N_27567);
and U28998 (N_28998,N_27515,N_27057);
or U28999 (N_28999,N_27385,N_27790);
and U29000 (N_29000,N_28160,N_28835);
xnor U29001 (N_29001,N_28876,N_28270);
nor U29002 (N_29002,N_28786,N_28006);
nand U29003 (N_29003,N_28243,N_28384);
xor U29004 (N_29004,N_28434,N_28927);
nand U29005 (N_29005,N_28616,N_28059);
and U29006 (N_29006,N_28668,N_28954);
nor U29007 (N_29007,N_28889,N_28105);
and U29008 (N_29008,N_28859,N_28338);
and U29009 (N_29009,N_28665,N_28248);
nor U29010 (N_29010,N_28683,N_28689);
nand U29011 (N_29011,N_28694,N_28370);
and U29012 (N_29012,N_28381,N_28048);
nor U29013 (N_29013,N_28698,N_28556);
nor U29014 (N_29014,N_28332,N_28432);
nor U29015 (N_29015,N_28379,N_28378);
nand U29016 (N_29016,N_28608,N_28416);
nand U29017 (N_29017,N_28017,N_28162);
nor U29018 (N_29018,N_28041,N_28574);
and U29019 (N_29019,N_28977,N_28020);
nor U29020 (N_29020,N_28777,N_28083);
xnor U29021 (N_29021,N_28173,N_28039);
and U29022 (N_29022,N_28558,N_28337);
xor U29023 (N_29023,N_28074,N_28206);
or U29024 (N_29024,N_28620,N_28084);
or U29025 (N_29025,N_28455,N_28691);
nor U29026 (N_29026,N_28544,N_28203);
nor U29027 (N_29027,N_28983,N_28483);
xnor U29028 (N_29028,N_28759,N_28457);
nand U29029 (N_29029,N_28225,N_28877);
nand U29030 (N_29030,N_28198,N_28852);
or U29031 (N_29031,N_28797,N_28580);
nor U29032 (N_29032,N_28813,N_28976);
or U29033 (N_29033,N_28655,N_28134);
and U29034 (N_29034,N_28547,N_28176);
and U29035 (N_29035,N_28593,N_28179);
nand U29036 (N_29036,N_28314,N_28145);
nor U29037 (N_29037,N_28437,N_28000);
nor U29038 (N_29038,N_28785,N_28796);
and U29039 (N_29039,N_28949,N_28576);
xor U29040 (N_29040,N_28768,N_28043);
nor U29041 (N_29041,N_28501,N_28431);
nand U29042 (N_29042,N_28422,N_28201);
xor U29043 (N_29043,N_28891,N_28677);
xnor U29044 (N_29044,N_28819,N_28879);
nand U29045 (N_29045,N_28180,N_28319);
xnor U29046 (N_29046,N_28617,N_28426);
nor U29047 (N_29047,N_28118,N_28454);
xnor U29048 (N_29048,N_28867,N_28607);
nand U29049 (N_29049,N_28257,N_28327);
nor U29050 (N_29050,N_28227,N_28538);
nor U29051 (N_29051,N_28534,N_28478);
nor U29052 (N_29052,N_28304,N_28393);
nor U29053 (N_29053,N_28849,N_28202);
and U29054 (N_29054,N_28758,N_28102);
or U29055 (N_29055,N_28108,N_28512);
nor U29056 (N_29056,N_28472,N_28467);
xnor U29057 (N_29057,N_28602,N_28791);
and U29058 (N_29058,N_28448,N_28679);
nor U29059 (N_29059,N_28260,N_28656);
or U29060 (N_29060,N_28794,N_28709);
xnor U29061 (N_29061,N_28042,N_28387);
and U29062 (N_29062,N_28900,N_28050);
or U29063 (N_29063,N_28433,N_28971);
and U29064 (N_29064,N_28934,N_28924);
and U29065 (N_29065,N_28452,N_28740);
and U29066 (N_29066,N_28858,N_28653);
or U29067 (N_29067,N_28294,N_28840);
nand U29068 (N_29068,N_28832,N_28326);
nor U29069 (N_29069,N_28494,N_28894);
xor U29070 (N_29070,N_28579,N_28864);
xor U29071 (N_29071,N_28098,N_28936);
and U29072 (N_29072,N_28263,N_28559);
nand U29073 (N_29073,N_28303,N_28570);
nand U29074 (N_29074,N_28364,N_28253);
xor U29075 (N_29075,N_28897,N_28566);
or U29076 (N_29076,N_28860,N_28024);
xnor U29077 (N_29077,N_28333,N_28836);
nor U29078 (N_29078,N_28237,N_28443);
nor U29079 (N_29079,N_28533,N_28097);
xor U29080 (N_29080,N_28716,N_28030);
nor U29081 (N_29081,N_28763,N_28869);
xor U29082 (N_29082,N_28301,N_28634);
nand U29083 (N_29083,N_28101,N_28053);
xnor U29084 (N_29084,N_28619,N_28537);
nand U29085 (N_29085,N_28669,N_28535);
or U29086 (N_29086,N_28947,N_28204);
xor U29087 (N_29087,N_28769,N_28489);
xnor U29088 (N_29088,N_28506,N_28492);
xor U29089 (N_29089,N_28128,N_28584);
nand U29090 (N_29090,N_28838,N_28135);
xor U29091 (N_29091,N_28905,N_28708);
nor U29092 (N_29092,N_28845,N_28016);
nand U29093 (N_29093,N_28514,N_28543);
and U29094 (N_29094,N_28803,N_28414);
and U29095 (N_29095,N_28438,N_28407);
or U29096 (N_29096,N_28783,N_28571);
and U29097 (N_29097,N_28439,N_28088);
nand U29098 (N_29098,N_28502,N_28300);
xnor U29099 (N_29099,N_28562,N_28264);
nor U29100 (N_29100,N_28311,N_28831);
xor U29101 (N_29101,N_28729,N_28194);
or U29102 (N_29102,N_28563,N_28895);
nand U29103 (N_29103,N_28825,N_28545);
nand U29104 (N_29104,N_28136,N_28092);
or U29105 (N_29105,N_28621,N_28505);
nor U29106 (N_29106,N_28417,N_28681);
and U29107 (N_29107,N_28887,N_28355);
or U29108 (N_29108,N_28091,N_28047);
and U29109 (N_29109,N_28989,N_28241);
or U29110 (N_29110,N_28124,N_28415);
or U29111 (N_29111,N_28643,N_28126);
nand U29112 (N_29112,N_28396,N_28664);
and U29113 (N_29113,N_28274,N_28627);
nand U29114 (N_29114,N_28650,N_28187);
xnor U29115 (N_29115,N_28207,N_28651);
or U29116 (N_29116,N_28508,N_28703);
nor U29117 (N_29117,N_28344,N_28346);
xor U29118 (N_29118,N_28036,N_28246);
nor U29119 (N_29119,N_28335,N_28262);
or U29120 (N_29120,N_28406,N_28373);
nor U29121 (N_29121,N_28171,N_28799);
nor U29122 (N_29122,N_28518,N_28987);
xor U29123 (N_29123,N_28585,N_28710);
and U29124 (N_29124,N_28780,N_28998);
and U29125 (N_29125,N_28837,N_28955);
and U29126 (N_29126,N_28159,N_28220);
or U29127 (N_29127,N_28038,N_28610);
xnor U29128 (N_29128,N_28200,N_28318);
and U29129 (N_29129,N_28549,N_28660);
nor U29130 (N_29130,N_28857,N_28425);
nor U29131 (N_29131,N_28466,N_28696);
nand U29132 (N_29132,N_28833,N_28890);
nor U29133 (N_29133,N_28469,N_28312);
nor U29134 (N_29134,N_28412,N_28907);
or U29135 (N_29135,N_28586,N_28002);
or U29136 (N_29136,N_28941,N_28914);
and U29137 (N_29137,N_28992,N_28340);
or U29138 (N_29138,N_28163,N_28517);
and U29139 (N_29139,N_28328,N_28261);
nand U29140 (N_29140,N_28063,N_28626);
nand U29141 (N_29141,N_28361,N_28244);
nor U29142 (N_29142,N_28186,N_28181);
or U29143 (N_29143,N_28685,N_28368);
nand U29144 (N_29144,N_28427,N_28034);
or U29145 (N_29145,N_28408,N_28625);
or U29146 (N_29146,N_28009,N_28345);
nor U29147 (N_29147,N_28285,N_28666);
or U29148 (N_29148,N_28276,N_28037);
xor U29149 (N_29149,N_28464,N_28480);
nor U29150 (N_29150,N_28103,N_28398);
or U29151 (N_29151,N_28307,N_28223);
nand U29152 (N_29152,N_28875,N_28904);
or U29153 (N_29153,N_28386,N_28076);
xor U29154 (N_29154,N_28193,N_28968);
nand U29155 (N_29155,N_28140,N_28320);
or U29156 (N_29156,N_28131,N_28606);
and U29157 (N_29157,N_28429,N_28497);
and U29158 (N_29158,N_28411,N_28604);
nor U29159 (N_29159,N_28536,N_28741);
or U29160 (N_29160,N_28881,N_28357);
xnor U29161 (N_29161,N_28188,N_28463);
xnor U29162 (N_29162,N_28280,N_28143);
nor U29163 (N_29163,N_28067,N_28692);
xnor U29164 (N_29164,N_28259,N_28935);
nand U29165 (N_29165,N_28526,N_28903);
nand U29166 (N_29166,N_28116,N_28524);
xnor U29167 (N_29167,N_28779,N_28590);
xnor U29168 (N_29168,N_28766,N_28045);
nor U29169 (N_29169,N_28495,N_28376);
or U29170 (N_29170,N_28189,N_28049);
nand U29171 (N_29171,N_28657,N_28238);
or U29172 (N_29172,N_28155,N_28086);
nand U29173 (N_29173,N_28111,N_28459);
and U29174 (N_29174,N_28633,N_28525);
xnor U29175 (N_29175,N_28991,N_28937);
nand U29176 (N_29176,N_28075,N_28725);
and U29177 (N_29177,N_28476,N_28926);
nor U29178 (N_29178,N_28372,N_28212);
nand U29179 (N_29179,N_28749,N_28289);
nand U29180 (N_29180,N_28474,N_28295);
or U29181 (N_29181,N_28290,N_28151);
and U29182 (N_29182,N_28702,N_28343);
xnor U29183 (N_29183,N_28652,N_28814);
or U29184 (N_29184,N_28445,N_28224);
and U29185 (N_29185,N_28302,N_28070);
nor U29186 (N_29186,N_28945,N_28636);
nor U29187 (N_29187,N_28109,N_28156);
nor U29188 (N_29188,N_28771,N_28035);
or U29189 (N_29189,N_28458,N_28752);
and U29190 (N_29190,N_28292,N_28004);
and U29191 (N_29191,N_28470,N_28950);
nand U29192 (N_29192,N_28168,N_28614);
nor U29193 (N_29193,N_28435,N_28854);
nand U29194 (N_29194,N_28919,N_28921);
nand U29195 (N_29195,N_28583,N_28054);
nor U29196 (N_29196,N_28520,N_28883);
and U29197 (N_29197,N_28217,N_28028);
xor U29198 (N_29198,N_28296,N_28984);
nor U29199 (N_29199,N_28085,N_28704);
xor U29200 (N_29200,N_28231,N_28661);
nand U29201 (N_29201,N_28960,N_28021);
and U29202 (N_29202,N_28242,N_28965);
xor U29203 (N_29203,N_28866,N_28802);
or U29204 (N_29204,N_28137,N_28659);
and U29205 (N_29205,N_28675,N_28615);
and U29206 (N_29206,N_28603,N_28349);
and U29207 (N_29207,N_28951,N_28804);
and U29208 (N_29208,N_28213,N_28851);
and U29209 (N_29209,N_28450,N_28229);
nand U29210 (N_29210,N_28940,N_28946);
nor U29211 (N_29211,N_28449,N_28061);
nor U29212 (N_29212,N_28809,N_28258);
or U29213 (N_29213,N_28504,N_28719);
nand U29214 (N_29214,N_28527,N_28874);
xor U29215 (N_29215,N_28632,N_28532);
or U29216 (N_29216,N_28315,N_28888);
nand U29217 (N_29217,N_28649,N_28358);
or U29218 (N_29218,N_28667,N_28183);
or U29219 (N_29219,N_28226,N_28982);
or U29220 (N_29220,N_28060,N_28844);
or U29221 (N_29221,N_28447,N_28684);
nand U29222 (N_29222,N_28701,N_28909);
or U29223 (N_29223,N_28461,N_28993);
nand U29224 (N_29224,N_28715,N_28912);
or U29225 (N_29225,N_28008,N_28848);
xor U29226 (N_29226,N_28961,N_28601);
or U29227 (N_29227,N_28613,N_28847);
or U29228 (N_29228,N_28266,N_28671);
or U29229 (N_29229,N_28931,N_28596);
nand U29230 (N_29230,N_28161,N_28271);
nor U29231 (N_29231,N_28309,N_28823);
xnor U29232 (N_29232,N_28107,N_28529);
nor U29233 (N_29233,N_28753,N_28323);
xnor U29234 (N_29234,N_28239,N_28595);
nand U29235 (N_29235,N_28686,N_28997);
nand U29236 (N_29236,N_28025,N_28784);
or U29237 (N_29237,N_28399,N_28170);
and U29238 (N_29238,N_28404,N_28530);
nor U29239 (N_29239,N_28498,N_28722);
and U29240 (N_29240,N_28871,N_28388);
and U29241 (N_29241,N_28221,N_28436);
or U29242 (N_29242,N_28901,N_28569);
and U29243 (N_29243,N_28055,N_28023);
nor U29244 (N_29244,N_28999,N_28597);
nor U29245 (N_29245,N_28523,N_28915);
or U29246 (N_29246,N_28861,N_28598);
or U29247 (N_29247,N_28305,N_28058);
nor U29248 (N_29248,N_28029,N_28930);
nand U29249 (N_29249,N_28727,N_28308);
and U29250 (N_29250,N_28122,N_28939);
nand U29251 (N_29251,N_28690,N_28959);
xnor U29252 (N_29252,N_28870,N_28885);
xnor U29253 (N_29253,N_28932,N_28115);
xor U29254 (N_29254,N_28313,N_28591);
nand U29255 (N_29255,N_28743,N_28232);
xnor U29256 (N_29256,N_28078,N_28046);
nor U29257 (N_29257,N_28707,N_28933);
nand U29258 (N_29258,N_28277,N_28697);
or U29259 (N_29259,N_28139,N_28149);
xor U29260 (N_29260,N_28988,N_28430);
nor U29261 (N_29261,N_28868,N_28051);
and U29262 (N_29262,N_28268,N_28711);
xor U29263 (N_29263,N_28363,N_28321);
nor U29264 (N_29264,N_28995,N_28555);
or U29265 (N_29265,N_28963,N_28782);
xor U29266 (N_29266,N_28377,N_28878);
and U29267 (N_29267,N_28440,N_28418);
nor U29268 (N_29268,N_28351,N_28747);
nor U29269 (N_29269,N_28948,N_28575);
and U29270 (N_29270,N_28392,N_28141);
and U29271 (N_29271,N_28916,N_28734);
and U29272 (N_29272,N_28811,N_28104);
or U29273 (N_29273,N_28542,N_28521);
xor U29274 (N_29274,N_28682,N_28561);
xnor U29275 (N_29275,N_28428,N_28540);
nor U29276 (N_29276,N_28082,N_28631);
or U29277 (N_29277,N_28678,N_28382);
or U29278 (N_29278,N_28451,N_28639);
nand U29279 (N_29279,N_28979,N_28310);
xnor U29280 (N_29280,N_28423,N_28475);
or U29281 (N_29281,N_28830,N_28552);
nand U29282 (N_29282,N_28056,N_28772);
nand U29283 (N_29283,N_28245,N_28641);
nand U29284 (N_29284,N_28093,N_28695);
nand U29285 (N_29285,N_28487,N_28331);
nand U29286 (N_29286,N_28284,N_28442);
nor U29287 (N_29287,N_28917,N_28330);
xnor U29288 (N_29288,N_28190,N_28491);
and U29289 (N_29289,N_28594,N_28329);
xor U29290 (N_29290,N_28721,N_28884);
nand U29291 (N_29291,N_28353,N_28110);
or U29292 (N_29292,N_28040,N_28177);
nand U29293 (N_29293,N_28985,N_28745);
and U29294 (N_29294,N_28744,N_28397);
nor U29295 (N_29295,N_28577,N_28390);
or U29296 (N_29296,N_28027,N_28672);
or U29297 (N_29297,N_28252,N_28928);
or U29298 (N_29298,N_28676,N_28424);
nor U29299 (N_29299,N_28365,N_28962);
or U29300 (N_29300,N_28953,N_28567);
or U29301 (N_29301,N_28462,N_28756);
xor U29302 (N_29302,N_28609,N_28007);
xor U29303 (N_29303,N_28015,N_28150);
xor U29304 (N_29304,N_28693,N_28739);
nor U29305 (N_29305,N_28477,N_28587);
xnor U29306 (N_29306,N_28994,N_28119);
nor U29307 (N_29307,N_28647,N_28589);
nand U29308 (N_29308,N_28638,N_28283);
or U29309 (N_29309,N_28142,N_28215);
and U29310 (N_29310,N_28444,N_28389);
or U29311 (N_29311,N_28720,N_28925);
or U29312 (N_29312,N_28820,N_28850);
nand U29313 (N_29313,N_28205,N_28842);
and U29314 (N_29314,N_28922,N_28717);
or U29315 (N_29315,N_28637,N_28158);
and U29316 (N_29316,N_28642,N_28712);
xnor U29317 (N_29317,N_28500,N_28872);
nand U29318 (N_29318,N_28735,N_28485);
nand U29319 (N_29319,N_28964,N_28360);
nor U29320 (N_29320,N_28371,N_28724);
or U29321 (N_29321,N_28383,N_28781);
and U29322 (N_29322,N_28622,N_28421);
nand U29323 (N_29323,N_28882,N_28990);
nand U29324 (N_29324,N_28843,N_28908);
nor U29325 (N_29325,N_28279,N_28453);
or U29326 (N_29326,N_28099,N_28281);
nand U29327 (N_29327,N_28793,N_28635);
nand U29328 (N_29328,N_28297,N_28736);
nand U29329 (N_29329,N_28249,N_28564);
nor U29330 (N_29330,N_28503,N_28348);
nor U29331 (N_29331,N_28446,N_28172);
or U29332 (N_29332,N_28493,N_28582);
xnor U29333 (N_29333,N_28209,N_28862);
nor U29334 (N_29334,N_28460,N_28726);
nand U29335 (N_29335,N_28828,N_28420);
or U29336 (N_29336,N_28658,N_28072);
and U29337 (N_29337,N_28052,N_28810);
or U29338 (N_29338,N_28611,N_28488);
nand U29339 (N_29339,N_28853,N_28911);
nand U29340 (N_29340,N_28507,N_28751);
nor U29341 (N_29341,N_28550,N_28073);
or U29342 (N_29342,N_28568,N_28481);
xor U29343 (N_29343,N_28129,N_28762);
xnor U29344 (N_29344,N_28560,N_28479);
or U29345 (N_29345,N_28765,N_28293);
nand U29346 (N_29346,N_28509,N_28391);
and U29347 (N_29347,N_28247,N_28402);
xor U29348 (N_29348,N_28064,N_28623);
nor U29349 (N_29349,N_28286,N_28113);
nor U29350 (N_29350,N_28972,N_28792);
xnor U29351 (N_29351,N_28011,N_28282);
or U29352 (N_29352,N_28095,N_28673);
nand U29353 (N_29353,N_28841,N_28970);
or U29354 (N_29354,N_28920,N_28750);
xnor U29355 (N_29355,N_28026,N_28981);
or U29356 (N_29356,N_28554,N_28146);
or U29357 (N_29357,N_28322,N_28732);
xnor U29358 (N_29358,N_28663,N_28367);
and U29359 (N_29359,N_28898,N_28612);
nand U29360 (N_29360,N_28010,N_28336);
xor U29361 (N_29361,N_28013,N_28182);
nor U29362 (N_29362,N_28256,N_28062);
xnor U29363 (N_29363,N_28822,N_28800);
and U29364 (N_29364,N_28152,N_28272);
and U29365 (N_29365,N_28291,N_28090);
and U29366 (N_29366,N_28354,N_28978);
nor U29367 (N_29367,N_28531,N_28807);
xor U29368 (N_29368,N_28275,N_28148);
nor U29369 (N_29369,N_28513,N_28899);
nand U29370 (N_29370,N_28031,N_28005);
xor U29371 (N_29371,N_28401,N_28299);
and U29372 (N_29372,N_28746,N_28952);
nor U29373 (N_29373,N_28254,N_28199);
xnor U29374 (N_29374,N_28886,N_28410);
xnor U29375 (N_29375,N_28240,N_28032);
nor U29376 (N_29376,N_28821,N_28516);
xnor U29377 (N_29377,N_28185,N_28125);
or U29378 (N_29378,N_28700,N_28214);
and U29379 (N_29379,N_28730,N_28572);
nand U29380 (N_29380,N_28081,N_28748);
nor U29381 (N_29381,N_28385,N_28066);
nor U29382 (N_29382,N_28334,N_28094);
xor U29383 (N_29383,N_28640,N_28628);
nand U29384 (N_29384,N_28767,N_28255);
nor U29385 (N_29385,N_28068,N_28798);
and U29386 (N_29386,N_28528,N_28251);
xor U29387 (N_29387,N_28519,N_28133);
xnor U29388 (N_29388,N_28629,N_28374);
or U29389 (N_29389,N_28395,N_28588);
and U29390 (N_29390,N_28403,N_28468);
and U29391 (N_29391,N_28269,N_28644);
nor U29392 (N_29392,N_28630,N_28757);
or U29393 (N_29393,N_28077,N_28863);
nor U29394 (N_29394,N_28482,N_28773);
nor U29395 (N_29395,N_28069,N_28775);
nor U29396 (N_29396,N_28728,N_28958);
or U29397 (N_29397,N_28789,N_28778);
or U29398 (N_29398,N_28022,N_28117);
nor U29399 (N_29399,N_28236,N_28196);
or U29400 (N_29400,N_28742,N_28515);
or U29401 (N_29401,N_28918,N_28827);
nor U29402 (N_29402,N_28648,N_28906);
or U29403 (N_29403,N_28014,N_28705);
and U29404 (N_29404,N_28706,N_28581);
or U29405 (N_29405,N_28369,N_28646);
xor U29406 (N_29406,N_28120,N_28551);
xor U29407 (N_29407,N_28973,N_28896);
nor U29408 (N_29408,N_28755,N_28208);
nor U29409 (N_29409,N_28618,N_28166);
nor U29410 (N_29410,N_28754,N_28265);
and U29411 (N_29411,N_28347,N_28127);
nor U29412 (N_29412,N_28233,N_28165);
xor U29413 (N_29413,N_28071,N_28219);
nor U29414 (N_29414,N_28967,N_28057);
or U29415 (N_29415,N_28670,N_28174);
nand U29416 (N_29416,N_28923,N_28210);
nand U29417 (N_29417,N_28278,N_28624);
nor U29418 (N_29418,N_28818,N_28795);
nand U29419 (N_29419,N_28806,N_28147);
nand U29420 (N_29420,N_28287,N_28599);
nor U29421 (N_29421,N_28829,N_28824);
nand U29422 (N_29422,N_28132,N_28316);
nand U29423 (N_29423,N_28511,N_28801);
and U29424 (N_29424,N_28812,N_28153);
nand U29425 (N_29425,N_28892,N_28273);
and U29426 (N_29426,N_28565,N_28980);
xor U29427 (N_29427,N_28178,N_28130);
xor U29428 (N_29428,N_28169,N_28065);
or U29429 (N_29429,N_28966,N_28230);
nand U29430 (N_29430,N_28044,N_28938);
xnor U29431 (N_29431,N_28154,N_28816);
nor U29432 (N_29432,N_28902,N_28761);
xnor U29433 (N_29433,N_28731,N_28674);
or U29434 (N_29434,N_28087,N_28471);
nor U29435 (N_29435,N_28100,N_28893);
nor U29436 (N_29436,N_28834,N_28510);
nor U29437 (N_29437,N_28815,N_28197);
nand U29438 (N_29438,N_28600,N_28121);
nand U29439 (N_29439,N_28079,N_28456);
nand U29440 (N_29440,N_28164,N_28317);
nand U29441 (N_29441,N_28910,N_28218);
nor U29442 (N_29442,N_28211,N_28826);
nor U29443 (N_29443,N_28298,N_28548);
nor U29444 (N_29444,N_28366,N_28788);
xnor U29445 (N_29445,N_28342,N_28405);
nand U29446 (N_29446,N_28486,N_28112);
nor U29447 (N_29447,N_28913,N_28409);
and U29448 (N_29448,N_28856,N_28592);
nand U29449 (N_29449,N_28996,N_28688);
nor U29450 (N_29450,N_28359,N_28033);
or U29451 (N_29451,N_28645,N_28123);
xnor U29452 (N_29452,N_28541,N_28718);
xor U29453 (N_29453,N_28764,N_28228);
and U29454 (N_29454,N_28413,N_28394);
nand U29455 (N_29455,N_28774,N_28490);
nor U29456 (N_29456,N_28805,N_28484);
nand U29457 (N_29457,N_28654,N_28096);
nor U29458 (N_29458,N_28499,N_28114);
nand U29459 (N_29459,N_28019,N_28003);
or U29460 (N_29460,N_28080,N_28195);
or U29461 (N_29461,N_28738,N_28012);
nor U29462 (N_29462,N_28975,N_28400);
and U29463 (N_29463,N_28846,N_28986);
or U29464 (N_29464,N_28699,N_28714);
xnor U29465 (N_29465,N_28380,N_28865);
or U29466 (N_29466,N_28737,N_28341);
and U29467 (N_29467,N_28943,N_28350);
xor U29468 (N_29468,N_28873,N_28539);
xor U29469 (N_29469,N_28362,N_28557);
or U29470 (N_29470,N_28356,N_28306);
nor U29471 (N_29471,N_28713,N_28662);
and U29472 (N_29472,N_28855,N_28522);
or U29473 (N_29473,N_28944,N_28578);
or U29474 (N_29474,N_28733,N_28234);
xnor U29475 (N_29475,N_28419,N_28235);
and U29476 (N_29476,N_28473,N_28138);
nand U29477 (N_29477,N_28222,N_28089);
and U29478 (N_29478,N_28680,N_28605);
nand U29479 (N_29479,N_28496,N_28817);
nand U29480 (N_29480,N_28573,N_28776);
and U29481 (N_29481,N_28325,N_28546);
nand U29482 (N_29482,N_28839,N_28956);
or U29483 (N_29483,N_28106,N_28267);
nor U29484 (N_29484,N_28324,N_28465);
xnor U29485 (N_29485,N_28375,N_28352);
xor U29486 (N_29486,N_28790,N_28787);
and U29487 (N_29487,N_28167,N_28880);
and U29488 (N_29488,N_28929,N_28250);
xor U29489 (N_29489,N_28339,N_28942);
nand U29490 (N_29490,N_28216,N_28553);
and U29491 (N_29491,N_28191,N_28001);
or U29492 (N_29492,N_28723,N_28144);
xor U29493 (N_29493,N_28018,N_28441);
or U29494 (N_29494,N_28957,N_28157);
nand U29495 (N_29495,N_28770,N_28687);
nand U29496 (N_29496,N_28288,N_28974);
and U29497 (N_29497,N_28808,N_28184);
or U29498 (N_29498,N_28175,N_28969);
or U29499 (N_29499,N_28760,N_28192);
nor U29500 (N_29500,N_28206,N_28221);
or U29501 (N_29501,N_28606,N_28996);
or U29502 (N_29502,N_28892,N_28777);
nand U29503 (N_29503,N_28670,N_28019);
xnor U29504 (N_29504,N_28758,N_28142);
and U29505 (N_29505,N_28176,N_28967);
xnor U29506 (N_29506,N_28749,N_28330);
nand U29507 (N_29507,N_28922,N_28401);
or U29508 (N_29508,N_28325,N_28690);
nand U29509 (N_29509,N_28564,N_28445);
and U29510 (N_29510,N_28955,N_28647);
and U29511 (N_29511,N_28534,N_28340);
nor U29512 (N_29512,N_28235,N_28394);
nand U29513 (N_29513,N_28740,N_28373);
or U29514 (N_29514,N_28627,N_28985);
nand U29515 (N_29515,N_28527,N_28505);
or U29516 (N_29516,N_28699,N_28355);
xnor U29517 (N_29517,N_28481,N_28853);
and U29518 (N_29518,N_28143,N_28919);
xor U29519 (N_29519,N_28071,N_28711);
and U29520 (N_29520,N_28788,N_28010);
xor U29521 (N_29521,N_28675,N_28150);
xor U29522 (N_29522,N_28562,N_28813);
xnor U29523 (N_29523,N_28281,N_28593);
nand U29524 (N_29524,N_28482,N_28493);
nor U29525 (N_29525,N_28176,N_28169);
nand U29526 (N_29526,N_28690,N_28418);
or U29527 (N_29527,N_28361,N_28552);
or U29528 (N_29528,N_28971,N_28397);
nor U29529 (N_29529,N_28790,N_28175);
or U29530 (N_29530,N_28620,N_28326);
nor U29531 (N_29531,N_28222,N_28327);
and U29532 (N_29532,N_28936,N_28982);
xnor U29533 (N_29533,N_28459,N_28258);
xor U29534 (N_29534,N_28326,N_28854);
nand U29535 (N_29535,N_28211,N_28184);
nor U29536 (N_29536,N_28449,N_28949);
or U29537 (N_29537,N_28246,N_28184);
nor U29538 (N_29538,N_28295,N_28808);
nand U29539 (N_29539,N_28106,N_28355);
or U29540 (N_29540,N_28363,N_28231);
or U29541 (N_29541,N_28250,N_28624);
nand U29542 (N_29542,N_28228,N_28367);
and U29543 (N_29543,N_28609,N_28628);
and U29544 (N_29544,N_28025,N_28665);
nand U29545 (N_29545,N_28623,N_28813);
xor U29546 (N_29546,N_28685,N_28596);
nand U29547 (N_29547,N_28807,N_28864);
nor U29548 (N_29548,N_28136,N_28726);
xnor U29549 (N_29549,N_28581,N_28027);
nor U29550 (N_29550,N_28590,N_28037);
nor U29551 (N_29551,N_28173,N_28235);
or U29552 (N_29552,N_28503,N_28691);
and U29553 (N_29553,N_28137,N_28066);
and U29554 (N_29554,N_28255,N_28295);
xnor U29555 (N_29555,N_28935,N_28558);
and U29556 (N_29556,N_28692,N_28576);
or U29557 (N_29557,N_28365,N_28745);
and U29558 (N_29558,N_28350,N_28379);
or U29559 (N_29559,N_28022,N_28764);
xor U29560 (N_29560,N_28604,N_28201);
or U29561 (N_29561,N_28974,N_28449);
or U29562 (N_29562,N_28097,N_28478);
nor U29563 (N_29563,N_28106,N_28119);
nand U29564 (N_29564,N_28446,N_28955);
nand U29565 (N_29565,N_28045,N_28238);
or U29566 (N_29566,N_28005,N_28426);
or U29567 (N_29567,N_28509,N_28540);
and U29568 (N_29568,N_28134,N_28181);
nor U29569 (N_29569,N_28901,N_28344);
nor U29570 (N_29570,N_28065,N_28373);
nor U29571 (N_29571,N_28766,N_28609);
or U29572 (N_29572,N_28504,N_28481);
nand U29573 (N_29573,N_28701,N_28599);
and U29574 (N_29574,N_28190,N_28824);
nor U29575 (N_29575,N_28094,N_28844);
nor U29576 (N_29576,N_28450,N_28465);
xor U29577 (N_29577,N_28214,N_28183);
xnor U29578 (N_29578,N_28399,N_28565);
nor U29579 (N_29579,N_28914,N_28431);
and U29580 (N_29580,N_28039,N_28491);
nand U29581 (N_29581,N_28019,N_28773);
xor U29582 (N_29582,N_28311,N_28699);
nor U29583 (N_29583,N_28236,N_28692);
nor U29584 (N_29584,N_28273,N_28221);
and U29585 (N_29585,N_28171,N_28533);
nor U29586 (N_29586,N_28754,N_28075);
xnor U29587 (N_29587,N_28735,N_28392);
nor U29588 (N_29588,N_28666,N_28102);
nor U29589 (N_29589,N_28920,N_28118);
xnor U29590 (N_29590,N_28082,N_28218);
nand U29591 (N_29591,N_28609,N_28242);
xnor U29592 (N_29592,N_28293,N_28019);
or U29593 (N_29593,N_28432,N_28138);
nand U29594 (N_29594,N_28495,N_28308);
nor U29595 (N_29595,N_28691,N_28854);
or U29596 (N_29596,N_28909,N_28413);
nor U29597 (N_29597,N_28889,N_28538);
xor U29598 (N_29598,N_28173,N_28149);
nor U29599 (N_29599,N_28681,N_28147);
xnor U29600 (N_29600,N_28842,N_28379);
xor U29601 (N_29601,N_28042,N_28074);
nor U29602 (N_29602,N_28783,N_28772);
nand U29603 (N_29603,N_28317,N_28380);
nor U29604 (N_29604,N_28252,N_28309);
xor U29605 (N_29605,N_28107,N_28532);
or U29606 (N_29606,N_28559,N_28025);
nand U29607 (N_29607,N_28160,N_28481);
xnor U29608 (N_29608,N_28977,N_28285);
nand U29609 (N_29609,N_28934,N_28359);
xnor U29610 (N_29610,N_28452,N_28958);
nor U29611 (N_29611,N_28918,N_28442);
or U29612 (N_29612,N_28022,N_28122);
xnor U29613 (N_29613,N_28194,N_28781);
xnor U29614 (N_29614,N_28835,N_28884);
nor U29615 (N_29615,N_28938,N_28608);
xnor U29616 (N_29616,N_28472,N_28636);
nand U29617 (N_29617,N_28436,N_28566);
and U29618 (N_29618,N_28596,N_28415);
nand U29619 (N_29619,N_28381,N_28757);
or U29620 (N_29620,N_28140,N_28432);
xnor U29621 (N_29621,N_28449,N_28332);
xor U29622 (N_29622,N_28841,N_28718);
nand U29623 (N_29623,N_28752,N_28019);
or U29624 (N_29624,N_28904,N_28462);
xor U29625 (N_29625,N_28882,N_28931);
and U29626 (N_29626,N_28336,N_28045);
nand U29627 (N_29627,N_28674,N_28092);
nand U29628 (N_29628,N_28701,N_28940);
nor U29629 (N_29629,N_28374,N_28158);
xnor U29630 (N_29630,N_28788,N_28259);
and U29631 (N_29631,N_28935,N_28204);
or U29632 (N_29632,N_28644,N_28071);
xor U29633 (N_29633,N_28108,N_28295);
xor U29634 (N_29634,N_28806,N_28928);
nand U29635 (N_29635,N_28531,N_28055);
nand U29636 (N_29636,N_28710,N_28749);
or U29637 (N_29637,N_28849,N_28029);
xnor U29638 (N_29638,N_28042,N_28506);
or U29639 (N_29639,N_28285,N_28303);
or U29640 (N_29640,N_28293,N_28685);
nor U29641 (N_29641,N_28547,N_28763);
or U29642 (N_29642,N_28649,N_28712);
nand U29643 (N_29643,N_28060,N_28415);
and U29644 (N_29644,N_28214,N_28414);
nor U29645 (N_29645,N_28585,N_28808);
nor U29646 (N_29646,N_28367,N_28278);
or U29647 (N_29647,N_28837,N_28429);
nor U29648 (N_29648,N_28905,N_28761);
xnor U29649 (N_29649,N_28636,N_28004);
and U29650 (N_29650,N_28298,N_28873);
or U29651 (N_29651,N_28570,N_28973);
nand U29652 (N_29652,N_28214,N_28412);
nor U29653 (N_29653,N_28169,N_28355);
and U29654 (N_29654,N_28275,N_28743);
and U29655 (N_29655,N_28088,N_28290);
xor U29656 (N_29656,N_28824,N_28687);
nand U29657 (N_29657,N_28011,N_28618);
xor U29658 (N_29658,N_28790,N_28043);
and U29659 (N_29659,N_28004,N_28957);
and U29660 (N_29660,N_28081,N_28142);
xnor U29661 (N_29661,N_28717,N_28857);
xor U29662 (N_29662,N_28222,N_28139);
nor U29663 (N_29663,N_28595,N_28243);
nor U29664 (N_29664,N_28160,N_28138);
nand U29665 (N_29665,N_28050,N_28957);
nor U29666 (N_29666,N_28809,N_28459);
nor U29667 (N_29667,N_28033,N_28056);
and U29668 (N_29668,N_28706,N_28757);
and U29669 (N_29669,N_28048,N_28009);
nor U29670 (N_29670,N_28492,N_28305);
nand U29671 (N_29671,N_28627,N_28022);
nand U29672 (N_29672,N_28733,N_28599);
or U29673 (N_29673,N_28757,N_28766);
nor U29674 (N_29674,N_28880,N_28169);
or U29675 (N_29675,N_28662,N_28221);
nand U29676 (N_29676,N_28562,N_28482);
nor U29677 (N_29677,N_28380,N_28347);
or U29678 (N_29678,N_28678,N_28421);
and U29679 (N_29679,N_28031,N_28911);
nor U29680 (N_29680,N_28685,N_28563);
nand U29681 (N_29681,N_28536,N_28169);
nand U29682 (N_29682,N_28590,N_28728);
nand U29683 (N_29683,N_28658,N_28589);
xor U29684 (N_29684,N_28607,N_28672);
or U29685 (N_29685,N_28444,N_28273);
nor U29686 (N_29686,N_28348,N_28624);
nor U29687 (N_29687,N_28116,N_28205);
or U29688 (N_29688,N_28644,N_28730);
and U29689 (N_29689,N_28037,N_28340);
nand U29690 (N_29690,N_28011,N_28233);
and U29691 (N_29691,N_28582,N_28849);
nand U29692 (N_29692,N_28441,N_28471);
or U29693 (N_29693,N_28312,N_28005);
and U29694 (N_29694,N_28247,N_28803);
nor U29695 (N_29695,N_28451,N_28215);
nand U29696 (N_29696,N_28650,N_28302);
nand U29697 (N_29697,N_28579,N_28819);
and U29698 (N_29698,N_28025,N_28806);
xor U29699 (N_29699,N_28428,N_28099);
nor U29700 (N_29700,N_28819,N_28410);
and U29701 (N_29701,N_28229,N_28598);
nor U29702 (N_29702,N_28407,N_28872);
xor U29703 (N_29703,N_28910,N_28647);
or U29704 (N_29704,N_28296,N_28176);
and U29705 (N_29705,N_28123,N_28991);
xnor U29706 (N_29706,N_28422,N_28870);
xnor U29707 (N_29707,N_28956,N_28852);
nor U29708 (N_29708,N_28291,N_28766);
xnor U29709 (N_29709,N_28431,N_28527);
nand U29710 (N_29710,N_28650,N_28219);
or U29711 (N_29711,N_28693,N_28410);
xnor U29712 (N_29712,N_28977,N_28828);
nand U29713 (N_29713,N_28358,N_28263);
xor U29714 (N_29714,N_28714,N_28662);
and U29715 (N_29715,N_28335,N_28297);
or U29716 (N_29716,N_28919,N_28512);
nor U29717 (N_29717,N_28387,N_28480);
xnor U29718 (N_29718,N_28693,N_28567);
and U29719 (N_29719,N_28902,N_28727);
xor U29720 (N_29720,N_28627,N_28442);
or U29721 (N_29721,N_28921,N_28129);
and U29722 (N_29722,N_28412,N_28352);
nand U29723 (N_29723,N_28238,N_28686);
and U29724 (N_29724,N_28230,N_28956);
or U29725 (N_29725,N_28041,N_28423);
nor U29726 (N_29726,N_28634,N_28307);
nor U29727 (N_29727,N_28928,N_28697);
or U29728 (N_29728,N_28643,N_28447);
nor U29729 (N_29729,N_28420,N_28584);
xor U29730 (N_29730,N_28239,N_28059);
nand U29731 (N_29731,N_28342,N_28841);
nand U29732 (N_29732,N_28327,N_28592);
nor U29733 (N_29733,N_28331,N_28239);
nand U29734 (N_29734,N_28048,N_28281);
xnor U29735 (N_29735,N_28096,N_28918);
or U29736 (N_29736,N_28584,N_28498);
xnor U29737 (N_29737,N_28210,N_28891);
xor U29738 (N_29738,N_28493,N_28525);
or U29739 (N_29739,N_28502,N_28409);
or U29740 (N_29740,N_28780,N_28846);
nor U29741 (N_29741,N_28220,N_28690);
xnor U29742 (N_29742,N_28373,N_28551);
nor U29743 (N_29743,N_28858,N_28396);
nand U29744 (N_29744,N_28425,N_28658);
and U29745 (N_29745,N_28303,N_28210);
nor U29746 (N_29746,N_28665,N_28995);
nor U29747 (N_29747,N_28993,N_28716);
or U29748 (N_29748,N_28645,N_28809);
nor U29749 (N_29749,N_28695,N_28959);
nand U29750 (N_29750,N_28301,N_28322);
nor U29751 (N_29751,N_28155,N_28101);
and U29752 (N_29752,N_28930,N_28286);
and U29753 (N_29753,N_28854,N_28125);
nor U29754 (N_29754,N_28837,N_28308);
nor U29755 (N_29755,N_28861,N_28397);
nor U29756 (N_29756,N_28579,N_28979);
nand U29757 (N_29757,N_28843,N_28154);
xnor U29758 (N_29758,N_28024,N_28935);
xor U29759 (N_29759,N_28466,N_28137);
or U29760 (N_29760,N_28430,N_28167);
nor U29761 (N_29761,N_28330,N_28881);
nand U29762 (N_29762,N_28161,N_28694);
nand U29763 (N_29763,N_28571,N_28740);
xor U29764 (N_29764,N_28816,N_28218);
nand U29765 (N_29765,N_28254,N_28634);
or U29766 (N_29766,N_28868,N_28990);
or U29767 (N_29767,N_28421,N_28492);
and U29768 (N_29768,N_28704,N_28154);
nor U29769 (N_29769,N_28459,N_28607);
or U29770 (N_29770,N_28799,N_28490);
and U29771 (N_29771,N_28878,N_28010);
xor U29772 (N_29772,N_28627,N_28472);
or U29773 (N_29773,N_28901,N_28585);
xor U29774 (N_29774,N_28559,N_28725);
nand U29775 (N_29775,N_28181,N_28504);
xor U29776 (N_29776,N_28104,N_28719);
nand U29777 (N_29777,N_28278,N_28483);
or U29778 (N_29778,N_28417,N_28068);
nor U29779 (N_29779,N_28823,N_28834);
and U29780 (N_29780,N_28080,N_28400);
nand U29781 (N_29781,N_28799,N_28769);
or U29782 (N_29782,N_28672,N_28863);
xnor U29783 (N_29783,N_28128,N_28004);
or U29784 (N_29784,N_28540,N_28796);
xnor U29785 (N_29785,N_28668,N_28455);
and U29786 (N_29786,N_28407,N_28747);
or U29787 (N_29787,N_28278,N_28991);
nand U29788 (N_29788,N_28986,N_28315);
nor U29789 (N_29789,N_28656,N_28920);
or U29790 (N_29790,N_28411,N_28255);
xor U29791 (N_29791,N_28512,N_28963);
nand U29792 (N_29792,N_28417,N_28019);
nand U29793 (N_29793,N_28151,N_28875);
xnor U29794 (N_29794,N_28310,N_28931);
nor U29795 (N_29795,N_28975,N_28821);
nand U29796 (N_29796,N_28479,N_28100);
or U29797 (N_29797,N_28691,N_28187);
nor U29798 (N_29798,N_28981,N_28613);
xnor U29799 (N_29799,N_28634,N_28309);
xnor U29800 (N_29800,N_28655,N_28602);
or U29801 (N_29801,N_28296,N_28776);
nand U29802 (N_29802,N_28966,N_28335);
nand U29803 (N_29803,N_28254,N_28574);
xor U29804 (N_29804,N_28799,N_28714);
nand U29805 (N_29805,N_28543,N_28125);
or U29806 (N_29806,N_28915,N_28195);
nand U29807 (N_29807,N_28412,N_28312);
nor U29808 (N_29808,N_28004,N_28810);
nor U29809 (N_29809,N_28719,N_28335);
xnor U29810 (N_29810,N_28637,N_28638);
and U29811 (N_29811,N_28727,N_28909);
nand U29812 (N_29812,N_28415,N_28660);
nand U29813 (N_29813,N_28254,N_28290);
or U29814 (N_29814,N_28308,N_28302);
and U29815 (N_29815,N_28852,N_28170);
nor U29816 (N_29816,N_28067,N_28370);
xor U29817 (N_29817,N_28898,N_28889);
or U29818 (N_29818,N_28730,N_28946);
nand U29819 (N_29819,N_28201,N_28502);
nor U29820 (N_29820,N_28596,N_28158);
nand U29821 (N_29821,N_28173,N_28288);
nor U29822 (N_29822,N_28419,N_28292);
nand U29823 (N_29823,N_28171,N_28732);
nand U29824 (N_29824,N_28182,N_28884);
xor U29825 (N_29825,N_28865,N_28504);
and U29826 (N_29826,N_28548,N_28088);
nand U29827 (N_29827,N_28035,N_28220);
nor U29828 (N_29828,N_28105,N_28144);
and U29829 (N_29829,N_28984,N_28120);
or U29830 (N_29830,N_28590,N_28468);
and U29831 (N_29831,N_28453,N_28982);
or U29832 (N_29832,N_28031,N_28793);
and U29833 (N_29833,N_28394,N_28824);
and U29834 (N_29834,N_28821,N_28174);
xor U29835 (N_29835,N_28428,N_28017);
and U29836 (N_29836,N_28756,N_28072);
and U29837 (N_29837,N_28343,N_28558);
xor U29838 (N_29838,N_28748,N_28814);
xnor U29839 (N_29839,N_28272,N_28091);
nor U29840 (N_29840,N_28837,N_28450);
nor U29841 (N_29841,N_28685,N_28984);
nand U29842 (N_29842,N_28700,N_28817);
xnor U29843 (N_29843,N_28098,N_28983);
nand U29844 (N_29844,N_28428,N_28299);
or U29845 (N_29845,N_28749,N_28626);
xnor U29846 (N_29846,N_28318,N_28478);
nor U29847 (N_29847,N_28269,N_28803);
xor U29848 (N_29848,N_28985,N_28543);
and U29849 (N_29849,N_28695,N_28059);
nand U29850 (N_29850,N_28039,N_28185);
xor U29851 (N_29851,N_28142,N_28049);
nor U29852 (N_29852,N_28845,N_28850);
nor U29853 (N_29853,N_28849,N_28507);
and U29854 (N_29854,N_28491,N_28604);
or U29855 (N_29855,N_28311,N_28360);
xnor U29856 (N_29856,N_28223,N_28671);
or U29857 (N_29857,N_28886,N_28567);
or U29858 (N_29858,N_28397,N_28293);
nor U29859 (N_29859,N_28459,N_28373);
or U29860 (N_29860,N_28256,N_28348);
nand U29861 (N_29861,N_28525,N_28004);
nand U29862 (N_29862,N_28777,N_28004);
and U29863 (N_29863,N_28391,N_28086);
and U29864 (N_29864,N_28813,N_28552);
nand U29865 (N_29865,N_28996,N_28157);
xnor U29866 (N_29866,N_28198,N_28521);
and U29867 (N_29867,N_28648,N_28302);
xor U29868 (N_29868,N_28901,N_28845);
xor U29869 (N_29869,N_28111,N_28178);
nor U29870 (N_29870,N_28778,N_28210);
nand U29871 (N_29871,N_28481,N_28715);
nor U29872 (N_29872,N_28668,N_28778);
nand U29873 (N_29873,N_28785,N_28781);
nand U29874 (N_29874,N_28095,N_28296);
or U29875 (N_29875,N_28542,N_28306);
xnor U29876 (N_29876,N_28802,N_28709);
or U29877 (N_29877,N_28420,N_28345);
or U29878 (N_29878,N_28430,N_28420);
nor U29879 (N_29879,N_28542,N_28118);
or U29880 (N_29880,N_28037,N_28819);
or U29881 (N_29881,N_28106,N_28613);
or U29882 (N_29882,N_28891,N_28473);
nand U29883 (N_29883,N_28509,N_28485);
or U29884 (N_29884,N_28809,N_28800);
nand U29885 (N_29885,N_28164,N_28109);
xor U29886 (N_29886,N_28416,N_28724);
nor U29887 (N_29887,N_28804,N_28626);
and U29888 (N_29888,N_28783,N_28929);
nand U29889 (N_29889,N_28972,N_28838);
and U29890 (N_29890,N_28309,N_28277);
and U29891 (N_29891,N_28848,N_28618);
xnor U29892 (N_29892,N_28143,N_28964);
nor U29893 (N_29893,N_28063,N_28613);
xnor U29894 (N_29894,N_28503,N_28380);
and U29895 (N_29895,N_28968,N_28312);
nor U29896 (N_29896,N_28192,N_28518);
nand U29897 (N_29897,N_28847,N_28896);
nand U29898 (N_29898,N_28168,N_28321);
nor U29899 (N_29899,N_28180,N_28555);
or U29900 (N_29900,N_28410,N_28966);
nor U29901 (N_29901,N_28162,N_28137);
or U29902 (N_29902,N_28371,N_28808);
xnor U29903 (N_29903,N_28020,N_28195);
or U29904 (N_29904,N_28374,N_28380);
xnor U29905 (N_29905,N_28797,N_28519);
or U29906 (N_29906,N_28395,N_28870);
or U29907 (N_29907,N_28647,N_28532);
or U29908 (N_29908,N_28089,N_28050);
or U29909 (N_29909,N_28259,N_28710);
and U29910 (N_29910,N_28244,N_28697);
or U29911 (N_29911,N_28258,N_28524);
or U29912 (N_29912,N_28179,N_28662);
nand U29913 (N_29913,N_28184,N_28377);
nand U29914 (N_29914,N_28951,N_28198);
nor U29915 (N_29915,N_28256,N_28203);
nand U29916 (N_29916,N_28462,N_28420);
or U29917 (N_29917,N_28831,N_28675);
nor U29918 (N_29918,N_28369,N_28454);
nor U29919 (N_29919,N_28442,N_28786);
xor U29920 (N_29920,N_28189,N_28370);
xnor U29921 (N_29921,N_28637,N_28528);
nor U29922 (N_29922,N_28792,N_28014);
xnor U29923 (N_29923,N_28742,N_28955);
nor U29924 (N_29924,N_28673,N_28291);
and U29925 (N_29925,N_28790,N_28925);
and U29926 (N_29926,N_28972,N_28717);
nor U29927 (N_29927,N_28304,N_28186);
xor U29928 (N_29928,N_28668,N_28185);
nand U29929 (N_29929,N_28204,N_28611);
and U29930 (N_29930,N_28586,N_28749);
nor U29931 (N_29931,N_28325,N_28051);
or U29932 (N_29932,N_28489,N_28861);
and U29933 (N_29933,N_28847,N_28780);
xnor U29934 (N_29934,N_28209,N_28046);
nor U29935 (N_29935,N_28525,N_28872);
nor U29936 (N_29936,N_28217,N_28267);
and U29937 (N_29937,N_28400,N_28451);
nor U29938 (N_29938,N_28917,N_28616);
nor U29939 (N_29939,N_28646,N_28854);
nand U29940 (N_29940,N_28624,N_28015);
xor U29941 (N_29941,N_28156,N_28405);
or U29942 (N_29942,N_28481,N_28869);
and U29943 (N_29943,N_28071,N_28720);
nand U29944 (N_29944,N_28801,N_28368);
and U29945 (N_29945,N_28551,N_28184);
xor U29946 (N_29946,N_28745,N_28808);
nand U29947 (N_29947,N_28044,N_28934);
nand U29948 (N_29948,N_28045,N_28752);
nor U29949 (N_29949,N_28219,N_28513);
nor U29950 (N_29950,N_28560,N_28106);
or U29951 (N_29951,N_28981,N_28883);
nand U29952 (N_29952,N_28240,N_28116);
and U29953 (N_29953,N_28208,N_28561);
xnor U29954 (N_29954,N_28143,N_28092);
and U29955 (N_29955,N_28654,N_28535);
nor U29956 (N_29956,N_28185,N_28151);
xnor U29957 (N_29957,N_28757,N_28053);
or U29958 (N_29958,N_28049,N_28788);
and U29959 (N_29959,N_28363,N_28170);
nor U29960 (N_29960,N_28942,N_28686);
xnor U29961 (N_29961,N_28374,N_28686);
and U29962 (N_29962,N_28990,N_28636);
nor U29963 (N_29963,N_28419,N_28918);
nand U29964 (N_29964,N_28495,N_28012);
xnor U29965 (N_29965,N_28001,N_28254);
nor U29966 (N_29966,N_28056,N_28619);
or U29967 (N_29967,N_28127,N_28369);
xnor U29968 (N_29968,N_28198,N_28028);
xnor U29969 (N_29969,N_28646,N_28458);
or U29970 (N_29970,N_28548,N_28788);
and U29971 (N_29971,N_28699,N_28255);
nor U29972 (N_29972,N_28294,N_28982);
nand U29973 (N_29973,N_28605,N_28108);
and U29974 (N_29974,N_28033,N_28440);
xor U29975 (N_29975,N_28205,N_28769);
nor U29976 (N_29976,N_28070,N_28648);
nor U29977 (N_29977,N_28165,N_28208);
nor U29978 (N_29978,N_28295,N_28176);
or U29979 (N_29979,N_28018,N_28897);
nor U29980 (N_29980,N_28529,N_28044);
nor U29981 (N_29981,N_28816,N_28951);
and U29982 (N_29982,N_28467,N_28239);
nor U29983 (N_29983,N_28520,N_28680);
and U29984 (N_29984,N_28339,N_28688);
xor U29985 (N_29985,N_28735,N_28729);
xnor U29986 (N_29986,N_28773,N_28280);
nand U29987 (N_29987,N_28689,N_28642);
xnor U29988 (N_29988,N_28121,N_28969);
and U29989 (N_29989,N_28102,N_28936);
or U29990 (N_29990,N_28186,N_28468);
or U29991 (N_29991,N_28038,N_28933);
xnor U29992 (N_29992,N_28136,N_28986);
or U29993 (N_29993,N_28908,N_28076);
xnor U29994 (N_29994,N_28201,N_28536);
xor U29995 (N_29995,N_28378,N_28360);
nand U29996 (N_29996,N_28442,N_28173);
nand U29997 (N_29997,N_28253,N_28860);
xor U29998 (N_29998,N_28681,N_28254);
nand U29999 (N_29999,N_28112,N_28742);
and UO_0 (O_0,N_29394,N_29279);
and UO_1 (O_1,N_29542,N_29509);
or UO_2 (O_2,N_29699,N_29124);
nor UO_3 (O_3,N_29893,N_29309);
or UO_4 (O_4,N_29799,N_29220);
xnor UO_5 (O_5,N_29596,N_29785);
nor UO_6 (O_6,N_29564,N_29551);
or UO_7 (O_7,N_29110,N_29044);
or UO_8 (O_8,N_29190,N_29515);
or UO_9 (O_9,N_29683,N_29924);
nor UO_10 (O_10,N_29278,N_29718);
nor UO_11 (O_11,N_29069,N_29362);
xnor UO_12 (O_12,N_29797,N_29882);
and UO_13 (O_13,N_29817,N_29080);
nand UO_14 (O_14,N_29557,N_29415);
nand UO_15 (O_15,N_29584,N_29488);
xor UO_16 (O_16,N_29134,N_29098);
or UO_17 (O_17,N_29533,N_29318);
nand UO_18 (O_18,N_29296,N_29210);
nand UO_19 (O_19,N_29512,N_29518);
or UO_20 (O_20,N_29418,N_29894);
xor UO_21 (O_21,N_29475,N_29986);
nand UO_22 (O_22,N_29015,N_29087);
and UO_23 (O_23,N_29253,N_29746);
or UO_24 (O_24,N_29131,N_29376);
xor UO_25 (O_25,N_29631,N_29139);
nor UO_26 (O_26,N_29915,N_29874);
nand UO_27 (O_27,N_29822,N_29402);
and UO_28 (O_28,N_29917,N_29659);
and UO_29 (O_29,N_29627,N_29320);
and UO_30 (O_30,N_29965,N_29504);
nor UO_31 (O_31,N_29148,N_29848);
xnor UO_32 (O_32,N_29103,N_29492);
nor UO_33 (O_33,N_29706,N_29593);
xor UO_34 (O_34,N_29897,N_29623);
nand UO_35 (O_35,N_29328,N_29229);
and UO_36 (O_36,N_29899,N_29960);
nand UO_37 (O_37,N_29828,N_29469);
nor UO_38 (O_38,N_29448,N_29176);
xnor UO_39 (O_39,N_29733,N_29355);
xor UO_40 (O_40,N_29952,N_29454);
nand UO_41 (O_41,N_29634,N_29910);
and UO_42 (O_42,N_29081,N_29668);
nor UO_43 (O_43,N_29608,N_29294);
xnor UO_44 (O_44,N_29745,N_29552);
or UO_45 (O_45,N_29285,N_29249);
nor UO_46 (O_46,N_29671,N_29521);
or UO_47 (O_47,N_29796,N_29479);
nor UO_48 (O_48,N_29427,N_29128);
and UO_49 (O_49,N_29905,N_29648);
or UO_50 (O_50,N_29039,N_29616);
or UO_51 (O_51,N_29814,N_29034);
xnor UO_52 (O_52,N_29714,N_29510);
and UO_53 (O_53,N_29990,N_29638);
and UO_54 (O_54,N_29858,N_29072);
nor UO_55 (O_55,N_29674,N_29600);
xnor UO_56 (O_56,N_29381,N_29179);
nor UO_57 (O_57,N_29985,N_29261);
nand UO_58 (O_58,N_29613,N_29251);
nor UO_59 (O_59,N_29404,N_29686);
and UO_60 (O_60,N_29938,N_29624);
xnor UO_61 (O_61,N_29653,N_29763);
or UO_62 (O_62,N_29784,N_29168);
or UO_63 (O_63,N_29541,N_29277);
nand UO_64 (O_64,N_29793,N_29393);
nor UO_65 (O_65,N_29963,N_29703);
or UO_66 (O_66,N_29825,N_29004);
and UO_67 (O_67,N_29767,N_29651);
nor UO_68 (O_68,N_29480,N_29524);
nand UO_69 (O_69,N_29511,N_29574);
xor UO_70 (O_70,N_29269,N_29619);
nor UO_71 (O_71,N_29367,N_29676);
and UO_72 (O_72,N_29612,N_29478);
nand UO_73 (O_73,N_29871,N_29169);
nor UO_74 (O_74,N_29104,N_29038);
or UO_75 (O_75,N_29312,N_29156);
and UO_76 (O_76,N_29961,N_29931);
and UO_77 (O_77,N_29282,N_29097);
and UO_78 (O_78,N_29336,N_29006);
xnor UO_79 (O_79,N_29374,N_29430);
or UO_80 (O_80,N_29221,N_29747);
nand UO_81 (O_81,N_29424,N_29754);
or UO_82 (O_82,N_29735,N_29610);
nand UO_83 (O_83,N_29117,N_29423);
or UO_84 (O_84,N_29892,N_29888);
nor UO_85 (O_85,N_29774,N_29741);
nand UO_86 (O_86,N_29723,N_29209);
xor UO_87 (O_87,N_29725,N_29572);
or UO_88 (O_88,N_29060,N_29916);
nand UO_89 (O_89,N_29493,N_29839);
nor UO_90 (O_90,N_29020,N_29455);
nand UO_91 (O_91,N_29062,N_29982);
and UO_92 (O_92,N_29660,N_29935);
nand UO_93 (O_93,N_29936,N_29213);
and UO_94 (O_94,N_29476,N_29219);
nor UO_95 (O_95,N_29450,N_29245);
and UO_96 (O_96,N_29885,N_29452);
and UO_97 (O_97,N_29136,N_29732);
xor UO_98 (O_98,N_29724,N_29028);
and UO_99 (O_99,N_29335,N_29519);
nand UO_100 (O_100,N_29204,N_29116);
and UO_101 (O_101,N_29920,N_29482);
nand UO_102 (O_102,N_29993,N_29205);
or UO_103 (O_103,N_29140,N_29843);
and UO_104 (O_104,N_29491,N_29776);
xnor UO_105 (O_105,N_29144,N_29902);
nand UO_106 (O_106,N_29445,N_29456);
or UO_107 (O_107,N_29236,N_29658);
and UO_108 (O_108,N_29588,N_29705);
and UO_109 (O_109,N_29422,N_29912);
xnor UO_110 (O_110,N_29884,N_29389);
nor UO_111 (O_111,N_29319,N_29687);
nor UO_112 (O_112,N_29127,N_29760);
or UO_113 (O_113,N_29262,N_29365);
xnor UO_114 (O_114,N_29440,N_29762);
and UO_115 (O_115,N_29955,N_29397);
and UO_116 (O_116,N_29495,N_29721);
nand UO_117 (O_117,N_29949,N_29155);
or UO_118 (O_118,N_29435,N_29748);
xor UO_119 (O_119,N_29000,N_29925);
nand UO_120 (O_120,N_29013,N_29766);
nand UO_121 (O_121,N_29070,N_29941);
nor UO_122 (O_122,N_29537,N_29881);
nor UO_123 (O_123,N_29406,N_29715);
nand UO_124 (O_124,N_29323,N_29517);
nand UO_125 (O_125,N_29505,N_29343);
or UO_126 (O_126,N_29212,N_29869);
xnor UO_127 (O_127,N_29570,N_29577);
xor UO_128 (O_128,N_29956,N_29298);
xnor UO_129 (O_129,N_29759,N_29387);
nand UO_130 (O_130,N_29642,N_29820);
or UO_131 (O_131,N_29121,N_29535);
and UO_132 (O_132,N_29347,N_29696);
xor UO_133 (O_133,N_29022,N_29073);
nor UO_134 (O_134,N_29772,N_29942);
nand UO_135 (O_135,N_29466,N_29290);
or UO_136 (O_136,N_29161,N_29101);
and UO_137 (O_137,N_29033,N_29964);
nand UO_138 (O_138,N_29958,N_29314);
nand UO_139 (O_139,N_29354,N_29576);
or UO_140 (O_140,N_29149,N_29165);
and UO_141 (O_141,N_29031,N_29585);
or UO_142 (O_142,N_29603,N_29657);
and UO_143 (O_143,N_29755,N_29866);
nor UO_144 (O_144,N_29934,N_29348);
or UO_145 (O_145,N_29421,N_29840);
nor UO_146 (O_146,N_29904,N_29462);
and UO_147 (O_147,N_29673,N_29722);
xnor UO_148 (O_148,N_29199,N_29802);
xnor UO_149 (O_149,N_29607,N_29646);
or UO_150 (O_150,N_29991,N_29324);
xor UO_151 (O_151,N_29474,N_29891);
and UO_152 (O_152,N_29863,N_29114);
or UO_153 (O_153,N_29272,N_29556);
nand UO_154 (O_154,N_29182,N_29138);
and UO_155 (O_155,N_29630,N_29340);
xor UO_156 (O_156,N_29077,N_29494);
nor UO_157 (O_157,N_29447,N_29239);
xnor UO_158 (O_158,N_29325,N_29644);
or UO_159 (O_159,N_29043,N_29166);
and UO_160 (O_160,N_29856,N_29808);
and UO_161 (O_161,N_29566,N_29609);
or UO_162 (O_162,N_29014,N_29068);
or UO_163 (O_163,N_29194,N_29614);
xnor UO_164 (O_164,N_29377,N_29242);
nand UO_165 (O_165,N_29813,N_29943);
and UO_166 (O_166,N_29834,N_29266);
nand UO_167 (O_167,N_29226,N_29786);
xnor UO_168 (O_168,N_29313,N_29939);
nand UO_169 (O_169,N_29503,N_29366);
or UO_170 (O_170,N_29270,N_29907);
nand UO_171 (O_171,N_29661,N_29224);
nor UO_172 (O_172,N_29879,N_29851);
nand UO_173 (O_173,N_29057,N_29407);
and UO_174 (O_174,N_29976,N_29757);
nand UO_175 (O_175,N_29065,N_29024);
nor UO_176 (O_176,N_29717,N_29308);
nand UO_177 (O_177,N_29720,N_29559);
and UO_178 (O_178,N_29208,N_29716);
or UO_179 (O_179,N_29263,N_29781);
or UO_180 (O_180,N_29315,N_29231);
xnor UO_181 (O_181,N_29558,N_29586);
and UO_182 (O_182,N_29416,N_29102);
or UO_183 (O_183,N_29408,N_29790);
or UO_184 (O_184,N_29983,N_29940);
nand UO_185 (O_185,N_29522,N_29122);
nand UO_186 (O_186,N_29711,N_29052);
nand UO_187 (O_187,N_29777,N_29174);
or UO_188 (O_188,N_29458,N_29211);
or UO_189 (O_189,N_29453,N_29538);
xor UO_190 (O_190,N_29800,N_29185);
xnor UO_191 (O_191,N_29146,N_29092);
or UO_192 (O_192,N_29353,N_29841);
xor UO_193 (O_193,N_29049,N_29743);
xnor UO_194 (O_194,N_29944,N_29809);
nor UO_195 (O_195,N_29526,N_29280);
nand UO_196 (O_196,N_29041,N_29135);
xor UO_197 (O_197,N_29195,N_29369);
nor UO_198 (O_198,N_29051,N_29921);
nor UO_199 (O_199,N_29929,N_29967);
xnor UO_200 (O_200,N_29598,N_29734);
nor UO_201 (O_201,N_29898,N_29405);
or UO_202 (O_202,N_29361,N_29271);
nor UO_203 (O_203,N_29063,N_29597);
or UO_204 (O_204,N_29257,N_29801);
or UO_205 (O_205,N_29930,N_29787);
xor UO_206 (O_206,N_29216,N_29439);
xnor UO_207 (O_207,N_29988,N_29130);
or UO_208 (O_208,N_29048,N_29392);
xnor UO_209 (O_209,N_29580,N_29481);
and UO_210 (O_210,N_29305,N_29042);
xnor UO_211 (O_211,N_29547,N_29465);
or UO_212 (O_212,N_29019,N_29240);
nand UO_213 (O_213,N_29693,N_29622);
nor UO_214 (O_214,N_29287,N_29625);
nor UO_215 (O_215,N_29618,N_29247);
nand UO_216 (O_216,N_29339,N_29821);
nand UO_217 (O_217,N_29016,N_29700);
xor UO_218 (O_218,N_29370,N_29544);
and UO_219 (O_219,N_29922,N_29901);
nand UO_220 (O_220,N_29710,N_29691);
or UO_221 (O_221,N_29502,N_29667);
or UO_222 (O_222,N_29968,N_29021);
and UO_223 (O_223,N_29184,N_29291);
nor UO_224 (O_224,N_29845,N_29554);
and UO_225 (O_225,N_29143,N_29601);
xor UO_226 (O_226,N_29293,N_29730);
xor UO_227 (O_227,N_29030,N_29007);
and UO_228 (O_228,N_29548,N_29690);
xnor UO_229 (O_229,N_29911,N_29260);
or UO_230 (O_230,N_29876,N_29789);
or UO_231 (O_231,N_29560,N_29744);
xnor UO_232 (O_232,N_29273,N_29230);
nand UO_233 (O_233,N_29284,N_29937);
nand UO_234 (O_234,N_29275,N_29023);
or UO_235 (O_235,N_29563,N_29419);
nor UO_236 (O_236,N_29302,N_29680);
and UO_237 (O_237,N_29694,N_29579);
and UO_238 (O_238,N_29972,N_29933);
nand UO_239 (O_239,N_29948,N_29334);
and UO_240 (O_240,N_29133,N_29451);
or UO_241 (O_241,N_29443,N_29798);
nand UO_242 (O_242,N_29794,N_29286);
nand UO_243 (O_243,N_29599,N_29765);
xnor UO_244 (O_244,N_29909,N_29360);
xnor UO_245 (O_245,N_29297,N_29568);
nand UO_246 (O_246,N_29385,N_29573);
nand UO_247 (O_247,N_29643,N_29737);
nand UO_248 (O_248,N_29193,N_29567);
and UO_249 (O_249,N_29726,N_29977);
and UO_250 (O_250,N_29141,N_29463);
xnor UO_251 (O_251,N_29583,N_29636);
xor UO_252 (O_252,N_29886,N_29032);
or UO_253 (O_253,N_29974,N_29561);
nor UO_254 (O_254,N_29536,N_29791);
and UO_255 (O_255,N_29649,N_29788);
nor UO_256 (O_256,N_29803,N_29237);
and UO_257 (O_257,N_29107,N_29756);
nor UO_258 (O_258,N_29926,N_29973);
and UO_259 (O_259,N_29989,N_29578);
or UO_260 (O_260,N_29186,N_29356);
and UO_261 (O_261,N_29698,N_29352);
nand UO_262 (O_262,N_29047,N_29025);
and UO_263 (O_263,N_29132,N_29433);
xor UO_264 (O_264,N_29592,N_29233);
nand UO_265 (O_265,N_29464,N_29980);
nor UO_266 (O_266,N_29675,N_29395);
xnor UO_267 (O_267,N_29729,N_29299);
nand UO_268 (O_268,N_29662,N_29040);
nand UO_269 (O_269,N_29327,N_29095);
and UO_270 (O_270,N_29546,N_29532);
or UO_271 (O_271,N_29379,N_29241);
xnor UO_272 (O_272,N_29889,N_29029);
nor UO_273 (O_273,N_29903,N_29540);
nor UO_274 (O_274,N_29425,N_29962);
nand UO_275 (O_275,N_29358,N_29322);
and UO_276 (O_276,N_29046,N_29770);
xnor UO_277 (O_277,N_29966,N_29461);
xor UO_278 (O_278,N_29196,N_29078);
xor UO_279 (O_279,N_29534,N_29550);
nor UO_280 (O_280,N_29307,N_29664);
or UO_281 (O_281,N_29545,N_29112);
xnor UO_282 (O_282,N_29056,N_29970);
or UO_283 (O_283,N_29617,N_29105);
and UO_284 (O_284,N_29398,N_29652);
and UO_285 (O_285,N_29214,N_29151);
and UO_286 (O_286,N_29751,N_29238);
nand UO_287 (O_287,N_29164,N_29005);
or UO_288 (O_288,N_29349,N_29513);
nor UO_289 (O_289,N_29685,N_29002);
nand UO_290 (O_290,N_29345,N_29258);
nor UO_291 (O_291,N_29248,N_29152);
nor UO_292 (O_292,N_29525,N_29227);
xor UO_293 (O_293,N_29692,N_29203);
or UO_294 (O_294,N_29640,N_29444);
nand UO_295 (O_295,N_29371,N_29945);
xnor UO_296 (O_296,N_29816,N_29728);
xnor UO_297 (O_297,N_29838,N_29357);
nand UO_298 (O_298,N_29329,N_29264);
nor UO_299 (O_299,N_29677,N_29276);
nor UO_300 (O_300,N_29655,N_29633);
or UO_301 (O_301,N_29842,N_29108);
and UO_302 (O_302,N_29228,N_29341);
nand UO_303 (O_303,N_29632,N_29459);
nor UO_304 (O_304,N_29750,N_29120);
xnor UO_305 (O_305,N_29805,N_29332);
or UO_306 (O_306,N_29310,N_29987);
and UO_307 (O_307,N_29064,N_29234);
or UO_308 (O_308,N_29778,N_29665);
nand UO_309 (O_309,N_29859,N_29189);
and UO_310 (O_310,N_29806,N_29670);
nand UO_311 (O_311,N_29549,N_29429);
and UO_312 (O_312,N_29847,N_29947);
or UO_313 (O_313,N_29679,N_29927);
and UO_314 (O_314,N_29123,N_29626);
xnor UO_315 (O_315,N_29113,N_29217);
nor UO_316 (O_316,N_29951,N_29412);
nand UO_317 (O_317,N_29467,N_29094);
xor UO_318 (O_318,N_29890,N_29244);
or UO_319 (O_319,N_29388,N_29562);
nand UO_320 (O_320,N_29844,N_29089);
or UO_321 (O_321,N_29997,N_29071);
nand UO_322 (O_322,N_29850,N_29605);
nand UO_323 (O_323,N_29058,N_29984);
nand UO_324 (O_324,N_29218,N_29831);
xnor UO_325 (O_325,N_29391,N_29254);
nor UO_326 (O_326,N_29027,N_29037);
and UO_327 (O_327,N_29202,N_29295);
xnor UO_328 (O_328,N_29923,N_29913);
xor UO_329 (O_329,N_29639,N_29172);
or UO_330 (O_330,N_29872,N_29994);
xor UO_331 (O_331,N_29350,N_29153);
nand UO_332 (O_332,N_29701,N_29075);
and UO_333 (O_333,N_29830,N_29590);
or UO_334 (O_334,N_29682,N_29017);
or UO_335 (O_335,N_29157,N_29232);
and UO_336 (O_336,N_29292,N_29250);
and UO_337 (O_337,N_29018,N_29971);
and UO_338 (O_338,N_29088,N_29473);
nor UO_339 (O_339,N_29914,N_29485);
xnor UO_340 (O_340,N_29628,N_29697);
and UO_341 (O_341,N_29181,N_29399);
nor UO_342 (O_342,N_29066,N_29708);
and UO_343 (O_343,N_29835,N_29035);
xnor UO_344 (O_344,N_29528,N_29861);
xor UO_345 (O_345,N_29010,N_29900);
and UO_346 (O_346,N_29177,N_29629);
or UO_347 (O_347,N_29400,N_29647);
and UO_348 (O_348,N_29446,N_29301);
and UO_349 (O_349,N_29738,N_29222);
nand UO_350 (O_350,N_29595,N_29666);
or UO_351 (O_351,N_29832,N_29688);
and UO_352 (O_352,N_29581,N_29337);
xor UO_353 (O_353,N_29142,N_29530);
xnor UO_354 (O_354,N_29497,N_29752);
nand UO_355 (O_355,N_29235,N_29093);
or UO_356 (O_356,N_29198,N_29001);
and UO_357 (O_357,N_29853,N_29496);
nand UO_358 (O_358,N_29390,N_29602);
and UO_359 (O_359,N_29300,N_29867);
nand UO_360 (O_360,N_29160,N_29719);
and UO_361 (O_361,N_29565,N_29106);
nor UO_362 (O_362,N_29712,N_29126);
xnor UO_363 (O_363,N_29259,N_29115);
nand UO_364 (O_364,N_29200,N_29477);
nand UO_365 (O_365,N_29543,N_29672);
nor UO_366 (O_366,N_29995,N_29981);
nor UO_367 (O_367,N_29173,N_29096);
nor UO_368 (O_368,N_29836,N_29411);
or UO_369 (O_369,N_29099,N_29441);
xor UO_370 (O_370,N_29978,N_29436);
nor UO_371 (O_371,N_29074,N_29810);
or UO_372 (O_372,N_29084,N_29050);
xnor UO_373 (O_373,N_29873,N_29026);
nand UO_374 (O_374,N_29396,N_29317);
nand UO_375 (O_375,N_29527,N_29877);
and UO_376 (O_376,N_29768,N_29621);
or UO_377 (O_377,N_29191,N_29739);
nand UO_378 (O_378,N_29875,N_29188);
and UO_379 (O_379,N_29154,N_29896);
xor UO_380 (O_380,N_29243,N_29187);
nor UO_381 (O_381,N_29795,N_29306);
nand UO_382 (O_382,N_29773,N_29403);
and UO_383 (O_383,N_29742,N_29067);
or UO_384 (O_384,N_29118,N_29819);
nand UO_385 (O_385,N_29571,N_29351);
nor UO_386 (O_386,N_29162,N_29555);
nor UO_387 (O_387,N_29998,N_29959);
nor UO_388 (O_388,N_29431,N_29008);
xor UO_389 (O_389,N_29499,N_29256);
xor UO_390 (O_390,N_29109,N_29594);
nand UO_391 (O_391,N_29587,N_29484);
xnor UO_392 (O_392,N_29255,N_29589);
nand UO_393 (O_393,N_29650,N_29758);
nor UO_394 (O_394,N_29330,N_29582);
nor UO_395 (O_395,N_29782,N_29316);
and UO_396 (O_396,N_29531,N_29225);
or UO_397 (O_397,N_29125,N_29783);
and UO_398 (O_398,N_29486,N_29061);
nor UO_399 (O_399,N_29011,N_29727);
nor UO_400 (O_400,N_29620,N_29171);
xor UO_401 (O_401,N_29274,N_29695);
xnor UO_402 (O_402,N_29604,N_29992);
nand UO_403 (O_403,N_29950,N_29908);
or UO_404 (O_404,N_29333,N_29090);
nor UO_405 (O_405,N_29201,N_29383);
or UO_406 (O_406,N_29410,N_29457);
or UO_407 (O_407,N_29880,N_29471);
nor UO_408 (O_408,N_29183,N_29342);
or UO_409 (O_409,N_29771,N_29862);
nor UO_410 (O_410,N_29637,N_29434);
and UO_411 (O_411,N_29304,N_29740);
xnor UO_412 (O_412,N_29823,N_29003);
nand UO_413 (O_413,N_29331,N_29311);
nor UO_414 (O_414,N_29175,N_29368);
xor UO_415 (O_415,N_29999,N_29338);
and UO_416 (O_416,N_29569,N_29460);
and UO_417 (O_417,N_29147,N_29413);
nand UO_418 (O_418,N_29380,N_29846);
or UO_419 (O_419,N_29837,N_29807);
nand UO_420 (O_420,N_29707,N_29969);
xnor UO_421 (O_421,N_29827,N_29382);
or UO_422 (O_422,N_29178,N_29753);
and UO_423 (O_423,N_29975,N_29860);
nor UO_424 (O_424,N_29163,N_29812);
nor UO_425 (O_425,N_29870,N_29954);
and UO_426 (O_426,N_29854,N_29438);
nor UO_427 (O_427,N_29520,N_29326);
nor UO_428 (O_428,N_29615,N_29170);
or UO_429 (O_429,N_29575,N_29953);
nor UO_430 (O_430,N_29137,N_29414);
nor UO_431 (O_431,N_29887,N_29288);
xor UO_432 (O_432,N_29363,N_29386);
nor UO_433 (O_433,N_29684,N_29946);
nand UO_434 (O_434,N_29468,N_29826);
xor UO_435 (O_435,N_29129,N_29764);
xor UO_436 (O_436,N_29761,N_29483);
nand UO_437 (O_437,N_29516,N_29815);
nand UO_438 (O_438,N_29223,N_29996);
xor UO_439 (O_439,N_29702,N_29957);
nand UO_440 (O_440,N_29704,N_29437);
nand UO_441 (O_441,N_29145,N_29378);
nand UO_442 (O_442,N_29252,N_29100);
and UO_443 (O_443,N_29811,N_29818);
and UO_444 (O_444,N_29059,N_29076);
and UO_445 (O_445,N_29656,N_29792);
nand UO_446 (O_446,N_29045,N_29091);
nand UO_447 (O_447,N_29681,N_29498);
or UO_448 (O_448,N_29281,N_29489);
or UO_449 (O_449,N_29979,N_29833);
nor UO_450 (O_450,N_29553,N_29780);
xor UO_451 (O_451,N_29928,N_29036);
nand UO_452 (O_452,N_29267,N_29428);
and UO_453 (O_453,N_29663,N_29508);
nor UO_454 (O_454,N_29111,N_29906);
or UO_455 (O_455,N_29487,N_29506);
xnor UO_456 (O_456,N_29054,N_29359);
and UO_457 (O_457,N_29409,N_29215);
xor UO_458 (O_458,N_29180,N_29207);
and UO_459 (O_459,N_29932,N_29611);
and UO_460 (O_460,N_29514,N_29426);
and UO_461 (O_461,N_29401,N_29344);
nor UO_462 (O_462,N_29529,N_29736);
xnor UO_463 (O_463,N_29206,N_29829);
nor UO_464 (O_464,N_29775,N_29918);
and UO_465 (O_465,N_29082,N_29669);
or UO_466 (O_466,N_29432,N_29731);
nand UO_467 (O_467,N_29150,N_29364);
nand UO_468 (O_468,N_29878,N_29384);
or UO_469 (O_469,N_29265,N_29268);
nor UO_470 (O_470,N_29449,N_29009);
nor UO_471 (O_471,N_29470,N_29283);
nor UO_472 (O_472,N_29417,N_29192);
and UO_473 (O_473,N_29303,N_29159);
nor UO_474 (O_474,N_29375,N_29864);
nand UO_475 (O_475,N_29654,N_29855);
nor UO_476 (O_476,N_29420,N_29373);
nand UO_477 (O_477,N_29868,N_29919);
and UO_478 (O_478,N_29085,N_29769);
nand UO_479 (O_479,N_29895,N_29053);
nand UO_480 (O_480,N_29865,N_29804);
and UO_481 (O_481,N_29086,N_29606);
xnor UO_482 (O_482,N_29079,N_29500);
nor UO_483 (O_483,N_29883,N_29709);
or UO_484 (O_484,N_29197,N_29852);
xor UO_485 (O_485,N_29678,N_29713);
nor UO_486 (O_486,N_29158,N_29246);
xor UO_487 (O_487,N_29119,N_29167);
or UO_488 (O_488,N_29641,N_29055);
and UO_489 (O_489,N_29321,N_29749);
or UO_490 (O_490,N_29849,N_29779);
xnor UO_491 (O_491,N_29501,N_29857);
and UO_492 (O_492,N_29289,N_29490);
or UO_493 (O_493,N_29012,N_29372);
and UO_494 (O_494,N_29523,N_29824);
xor UO_495 (O_495,N_29507,N_29346);
xnor UO_496 (O_496,N_29083,N_29645);
and UO_497 (O_497,N_29689,N_29635);
nand UO_498 (O_498,N_29591,N_29472);
or UO_499 (O_499,N_29539,N_29442);
or UO_500 (O_500,N_29361,N_29507);
or UO_501 (O_501,N_29749,N_29095);
nand UO_502 (O_502,N_29523,N_29553);
nor UO_503 (O_503,N_29098,N_29827);
or UO_504 (O_504,N_29865,N_29623);
nand UO_505 (O_505,N_29504,N_29709);
xnor UO_506 (O_506,N_29816,N_29981);
or UO_507 (O_507,N_29865,N_29064);
or UO_508 (O_508,N_29008,N_29647);
nor UO_509 (O_509,N_29932,N_29518);
nor UO_510 (O_510,N_29187,N_29351);
nand UO_511 (O_511,N_29342,N_29144);
nand UO_512 (O_512,N_29635,N_29850);
xnor UO_513 (O_513,N_29190,N_29385);
and UO_514 (O_514,N_29929,N_29159);
nand UO_515 (O_515,N_29998,N_29280);
nand UO_516 (O_516,N_29371,N_29216);
xnor UO_517 (O_517,N_29441,N_29190);
and UO_518 (O_518,N_29248,N_29365);
and UO_519 (O_519,N_29725,N_29381);
nand UO_520 (O_520,N_29722,N_29469);
xor UO_521 (O_521,N_29335,N_29121);
and UO_522 (O_522,N_29065,N_29013);
xor UO_523 (O_523,N_29516,N_29819);
xnor UO_524 (O_524,N_29789,N_29589);
and UO_525 (O_525,N_29506,N_29490);
nand UO_526 (O_526,N_29970,N_29878);
nand UO_527 (O_527,N_29714,N_29873);
nor UO_528 (O_528,N_29728,N_29727);
and UO_529 (O_529,N_29045,N_29196);
or UO_530 (O_530,N_29239,N_29296);
nor UO_531 (O_531,N_29168,N_29033);
and UO_532 (O_532,N_29520,N_29555);
or UO_533 (O_533,N_29961,N_29855);
or UO_534 (O_534,N_29808,N_29116);
nor UO_535 (O_535,N_29722,N_29244);
xnor UO_536 (O_536,N_29015,N_29413);
nand UO_537 (O_537,N_29356,N_29605);
nand UO_538 (O_538,N_29678,N_29017);
nand UO_539 (O_539,N_29608,N_29382);
or UO_540 (O_540,N_29779,N_29001);
and UO_541 (O_541,N_29009,N_29313);
and UO_542 (O_542,N_29966,N_29873);
and UO_543 (O_543,N_29140,N_29058);
nand UO_544 (O_544,N_29965,N_29027);
nor UO_545 (O_545,N_29642,N_29157);
nor UO_546 (O_546,N_29314,N_29977);
nor UO_547 (O_547,N_29740,N_29907);
nand UO_548 (O_548,N_29067,N_29969);
nor UO_549 (O_549,N_29892,N_29623);
or UO_550 (O_550,N_29021,N_29535);
or UO_551 (O_551,N_29268,N_29825);
and UO_552 (O_552,N_29304,N_29454);
or UO_553 (O_553,N_29159,N_29249);
nand UO_554 (O_554,N_29231,N_29292);
nand UO_555 (O_555,N_29293,N_29485);
nand UO_556 (O_556,N_29451,N_29854);
and UO_557 (O_557,N_29428,N_29393);
nor UO_558 (O_558,N_29378,N_29186);
nand UO_559 (O_559,N_29192,N_29253);
xor UO_560 (O_560,N_29718,N_29085);
xor UO_561 (O_561,N_29024,N_29953);
nor UO_562 (O_562,N_29282,N_29226);
nor UO_563 (O_563,N_29543,N_29076);
nand UO_564 (O_564,N_29723,N_29453);
nand UO_565 (O_565,N_29291,N_29271);
nand UO_566 (O_566,N_29980,N_29705);
xnor UO_567 (O_567,N_29431,N_29107);
or UO_568 (O_568,N_29213,N_29343);
nor UO_569 (O_569,N_29098,N_29361);
xor UO_570 (O_570,N_29379,N_29947);
nor UO_571 (O_571,N_29501,N_29313);
nand UO_572 (O_572,N_29991,N_29065);
nor UO_573 (O_573,N_29193,N_29086);
nand UO_574 (O_574,N_29462,N_29460);
and UO_575 (O_575,N_29977,N_29518);
nand UO_576 (O_576,N_29701,N_29562);
nor UO_577 (O_577,N_29876,N_29930);
nor UO_578 (O_578,N_29013,N_29400);
and UO_579 (O_579,N_29838,N_29122);
nand UO_580 (O_580,N_29336,N_29400);
nor UO_581 (O_581,N_29668,N_29300);
nor UO_582 (O_582,N_29254,N_29363);
xnor UO_583 (O_583,N_29958,N_29553);
or UO_584 (O_584,N_29825,N_29450);
nor UO_585 (O_585,N_29211,N_29838);
nand UO_586 (O_586,N_29398,N_29473);
nand UO_587 (O_587,N_29309,N_29811);
or UO_588 (O_588,N_29676,N_29848);
and UO_589 (O_589,N_29151,N_29164);
nand UO_590 (O_590,N_29528,N_29877);
or UO_591 (O_591,N_29399,N_29210);
or UO_592 (O_592,N_29957,N_29576);
xnor UO_593 (O_593,N_29630,N_29672);
nand UO_594 (O_594,N_29444,N_29347);
xor UO_595 (O_595,N_29556,N_29523);
xnor UO_596 (O_596,N_29684,N_29204);
nand UO_597 (O_597,N_29385,N_29877);
xor UO_598 (O_598,N_29503,N_29058);
xor UO_599 (O_599,N_29956,N_29866);
or UO_600 (O_600,N_29941,N_29066);
nor UO_601 (O_601,N_29127,N_29479);
or UO_602 (O_602,N_29325,N_29995);
nand UO_603 (O_603,N_29183,N_29221);
or UO_604 (O_604,N_29291,N_29333);
xor UO_605 (O_605,N_29074,N_29171);
or UO_606 (O_606,N_29196,N_29106);
nand UO_607 (O_607,N_29960,N_29770);
nor UO_608 (O_608,N_29143,N_29040);
or UO_609 (O_609,N_29509,N_29364);
or UO_610 (O_610,N_29832,N_29356);
xnor UO_611 (O_611,N_29252,N_29526);
and UO_612 (O_612,N_29449,N_29331);
nand UO_613 (O_613,N_29403,N_29988);
or UO_614 (O_614,N_29988,N_29986);
nor UO_615 (O_615,N_29048,N_29931);
and UO_616 (O_616,N_29322,N_29561);
and UO_617 (O_617,N_29879,N_29952);
and UO_618 (O_618,N_29516,N_29373);
xor UO_619 (O_619,N_29553,N_29358);
and UO_620 (O_620,N_29605,N_29728);
nand UO_621 (O_621,N_29924,N_29208);
or UO_622 (O_622,N_29758,N_29015);
nand UO_623 (O_623,N_29778,N_29739);
or UO_624 (O_624,N_29312,N_29125);
and UO_625 (O_625,N_29908,N_29660);
and UO_626 (O_626,N_29411,N_29454);
xor UO_627 (O_627,N_29667,N_29259);
or UO_628 (O_628,N_29923,N_29520);
nand UO_629 (O_629,N_29396,N_29993);
and UO_630 (O_630,N_29740,N_29945);
and UO_631 (O_631,N_29385,N_29293);
nand UO_632 (O_632,N_29440,N_29736);
xor UO_633 (O_633,N_29730,N_29100);
xnor UO_634 (O_634,N_29969,N_29719);
nor UO_635 (O_635,N_29215,N_29940);
xor UO_636 (O_636,N_29172,N_29686);
nor UO_637 (O_637,N_29185,N_29595);
xnor UO_638 (O_638,N_29068,N_29268);
xnor UO_639 (O_639,N_29660,N_29363);
and UO_640 (O_640,N_29970,N_29322);
nand UO_641 (O_641,N_29880,N_29286);
nand UO_642 (O_642,N_29681,N_29570);
or UO_643 (O_643,N_29281,N_29332);
xor UO_644 (O_644,N_29234,N_29555);
nor UO_645 (O_645,N_29768,N_29180);
or UO_646 (O_646,N_29840,N_29764);
nand UO_647 (O_647,N_29722,N_29355);
and UO_648 (O_648,N_29238,N_29132);
or UO_649 (O_649,N_29193,N_29068);
or UO_650 (O_650,N_29271,N_29872);
nand UO_651 (O_651,N_29176,N_29709);
nand UO_652 (O_652,N_29099,N_29148);
nor UO_653 (O_653,N_29048,N_29131);
or UO_654 (O_654,N_29639,N_29251);
and UO_655 (O_655,N_29574,N_29577);
nor UO_656 (O_656,N_29432,N_29735);
nand UO_657 (O_657,N_29313,N_29770);
nor UO_658 (O_658,N_29591,N_29914);
nand UO_659 (O_659,N_29795,N_29096);
xnor UO_660 (O_660,N_29674,N_29631);
and UO_661 (O_661,N_29647,N_29325);
nor UO_662 (O_662,N_29298,N_29933);
and UO_663 (O_663,N_29899,N_29450);
nor UO_664 (O_664,N_29928,N_29152);
and UO_665 (O_665,N_29951,N_29067);
nand UO_666 (O_666,N_29181,N_29471);
or UO_667 (O_667,N_29338,N_29347);
nor UO_668 (O_668,N_29900,N_29165);
and UO_669 (O_669,N_29276,N_29247);
xor UO_670 (O_670,N_29594,N_29647);
or UO_671 (O_671,N_29170,N_29658);
nor UO_672 (O_672,N_29520,N_29573);
nor UO_673 (O_673,N_29274,N_29111);
xor UO_674 (O_674,N_29101,N_29995);
nor UO_675 (O_675,N_29769,N_29189);
nand UO_676 (O_676,N_29910,N_29930);
nor UO_677 (O_677,N_29874,N_29097);
xnor UO_678 (O_678,N_29307,N_29071);
xor UO_679 (O_679,N_29084,N_29562);
and UO_680 (O_680,N_29953,N_29019);
nor UO_681 (O_681,N_29705,N_29128);
xnor UO_682 (O_682,N_29035,N_29889);
nor UO_683 (O_683,N_29135,N_29585);
or UO_684 (O_684,N_29451,N_29142);
or UO_685 (O_685,N_29511,N_29116);
xor UO_686 (O_686,N_29732,N_29664);
nor UO_687 (O_687,N_29051,N_29588);
and UO_688 (O_688,N_29227,N_29152);
and UO_689 (O_689,N_29381,N_29513);
nor UO_690 (O_690,N_29626,N_29814);
and UO_691 (O_691,N_29028,N_29125);
or UO_692 (O_692,N_29104,N_29406);
nor UO_693 (O_693,N_29118,N_29562);
or UO_694 (O_694,N_29702,N_29887);
nand UO_695 (O_695,N_29001,N_29410);
or UO_696 (O_696,N_29455,N_29893);
xor UO_697 (O_697,N_29023,N_29999);
or UO_698 (O_698,N_29032,N_29129);
nor UO_699 (O_699,N_29096,N_29691);
and UO_700 (O_700,N_29851,N_29863);
xor UO_701 (O_701,N_29208,N_29571);
and UO_702 (O_702,N_29769,N_29063);
nor UO_703 (O_703,N_29189,N_29942);
xor UO_704 (O_704,N_29207,N_29974);
xor UO_705 (O_705,N_29579,N_29836);
nand UO_706 (O_706,N_29389,N_29501);
nor UO_707 (O_707,N_29699,N_29138);
or UO_708 (O_708,N_29062,N_29568);
nand UO_709 (O_709,N_29762,N_29656);
and UO_710 (O_710,N_29697,N_29763);
and UO_711 (O_711,N_29922,N_29230);
nand UO_712 (O_712,N_29206,N_29082);
xor UO_713 (O_713,N_29384,N_29844);
nand UO_714 (O_714,N_29321,N_29312);
xnor UO_715 (O_715,N_29227,N_29973);
nor UO_716 (O_716,N_29190,N_29884);
and UO_717 (O_717,N_29418,N_29943);
nor UO_718 (O_718,N_29917,N_29566);
xor UO_719 (O_719,N_29588,N_29241);
nor UO_720 (O_720,N_29432,N_29429);
or UO_721 (O_721,N_29351,N_29444);
or UO_722 (O_722,N_29198,N_29480);
and UO_723 (O_723,N_29701,N_29611);
or UO_724 (O_724,N_29558,N_29679);
nor UO_725 (O_725,N_29747,N_29219);
nand UO_726 (O_726,N_29534,N_29863);
nor UO_727 (O_727,N_29510,N_29158);
or UO_728 (O_728,N_29637,N_29799);
nor UO_729 (O_729,N_29267,N_29729);
nor UO_730 (O_730,N_29841,N_29883);
nor UO_731 (O_731,N_29966,N_29227);
xnor UO_732 (O_732,N_29300,N_29996);
xnor UO_733 (O_733,N_29757,N_29827);
xnor UO_734 (O_734,N_29923,N_29185);
nor UO_735 (O_735,N_29821,N_29366);
nand UO_736 (O_736,N_29027,N_29624);
xnor UO_737 (O_737,N_29593,N_29808);
or UO_738 (O_738,N_29046,N_29760);
and UO_739 (O_739,N_29619,N_29989);
nor UO_740 (O_740,N_29387,N_29488);
or UO_741 (O_741,N_29002,N_29454);
xor UO_742 (O_742,N_29381,N_29461);
and UO_743 (O_743,N_29387,N_29825);
nand UO_744 (O_744,N_29745,N_29351);
xor UO_745 (O_745,N_29764,N_29880);
nor UO_746 (O_746,N_29181,N_29414);
nor UO_747 (O_747,N_29856,N_29155);
and UO_748 (O_748,N_29105,N_29541);
xnor UO_749 (O_749,N_29066,N_29112);
nand UO_750 (O_750,N_29216,N_29838);
xnor UO_751 (O_751,N_29766,N_29970);
nor UO_752 (O_752,N_29594,N_29879);
nand UO_753 (O_753,N_29941,N_29026);
nor UO_754 (O_754,N_29803,N_29930);
nand UO_755 (O_755,N_29714,N_29871);
and UO_756 (O_756,N_29204,N_29224);
nor UO_757 (O_757,N_29829,N_29298);
nor UO_758 (O_758,N_29107,N_29618);
or UO_759 (O_759,N_29107,N_29078);
xnor UO_760 (O_760,N_29660,N_29661);
or UO_761 (O_761,N_29482,N_29857);
nand UO_762 (O_762,N_29934,N_29533);
and UO_763 (O_763,N_29101,N_29358);
nand UO_764 (O_764,N_29435,N_29057);
nand UO_765 (O_765,N_29706,N_29179);
or UO_766 (O_766,N_29414,N_29500);
and UO_767 (O_767,N_29362,N_29986);
nor UO_768 (O_768,N_29060,N_29653);
xnor UO_769 (O_769,N_29648,N_29481);
nor UO_770 (O_770,N_29635,N_29833);
xor UO_771 (O_771,N_29791,N_29098);
xnor UO_772 (O_772,N_29354,N_29235);
and UO_773 (O_773,N_29996,N_29605);
xor UO_774 (O_774,N_29504,N_29850);
xnor UO_775 (O_775,N_29812,N_29042);
nor UO_776 (O_776,N_29346,N_29936);
or UO_777 (O_777,N_29633,N_29254);
nor UO_778 (O_778,N_29092,N_29193);
nor UO_779 (O_779,N_29357,N_29289);
nand UO_780 (O_780,N_29326,N_29553);
or UO_781 (O_781,N_29646,N_29430);
or UO_782 (O_782,N_29386,N_29343);
nor UO_783 (O_783,N_29869,N_29885);
nor UO_784 (O_784,N_29922,N_29568);
xor UO_785 (O_785,N_29376,N_29270);
or UO_786 (O_786,N_29812,N_29616);
or UO_787 (O_787,N_29603,N_29822);
xnor UO_788 (O_788,N_29667,N_29121);
nand UO_789 (O_789,N_29085,N_29498);
and UO_790 (O_790,N_29639,N_29674);
nand UO_791 (O_791,N_29366,N_29953);
xnor UO_792 (O_792,N_29321,N_29950);
nand UO_793 (O_793,N_29589,N_29663);
nand UO_794 (O_794,N_29645,N_29959);
or UO_795 (O_795,N_29636,N_29577);
nor UO_796 (O_796,N_29411,N_29088);
xor UO_797 (O_797,N_29394,N_29126);
nand UO_798 (O_798,N_29422,N_29040);
nor UO_799 (O_799,N_29862,N_29759);
or UO_800 (O_800,N_29393,N_29854);
nand UO_801 (O_801,N_29903,N_29438);
and UO_802 (O_802,N_29487,N_29878);
or UO_803 (O_803,N_29313,N_29745);
or UO_804 (O_804,N_29865,N_29191);
nand UO_805 (O_805,N_29764,N_29517);
nand UO_806 (O_806,N_29987,N_29102);
nor UO_807 (O_807,N_29195,N_29223);
and UO_808 (O_808,N_29309,N_29913);
nand UO_809 (O_809,N_29258,N_29438);
or UO_810 (O_810,N_29783,N_29429);
and UO_811 (O_811,N_29340,N_29364);
or UO_812 (O_812,N_29847,N_29011);
and UO_813 (O_813,N_29394,N_29669);
xnor UO_814 (O_814,N_29336,N_29468);
xnor UO_815 (O_815,N_29057,N_29980);
and UO_816 (O_816,N_29455,N_29609);
xnor UO_817 (O_817,N_29617,N_29419);
or UO_818 (O_818,N_29023,N_29720);
xnor UO_819 (O_819,N_29697,N_29229);
and UO_820 (O_820,N_29499,N_29211);
or UO_821 (O_821,N_29987,N_29567);
and UO_822 (O_822,N_29418,N_29197);
nor UO_823 (O_823,N_29687,N_29218);
nor UO_824 (O_824,N_29504,N_29066);
nor UO_825 (O_825,N_29765,N_29238);
and UO_826 (O_826,N_29414,N_29580);
nor UO_827 (O_827,N_29474,N_29061);
or UO_828 (O_828,N_29296,N_29487);
nor UO_829 (O_829,N_29847,N_29309);
nand UO_830 (O_830,N_29157,N_29770);
or UO_831 (O_831,N_29600,N_29804);
nor UO_832 (O_832,N_29603,N_29998);
xnor UO_833 (O_833,N_29958,N_29063);
nor UO_834 (O_834,N_29395,N_29681);
nor UO_835 (O_835,N_29667,N_29358);
nor UO_836 (O_836,N_29499,N_29314);
nand UO_837 (O_837,N_29892,N_29609);
and UO_838 (O_838,N_29185,N_29661);
xor UO_839 (O_839,N_29341,N_29723);
nand UO_840 (O_840,N_29234,N_29340);
nor UO_841 (O_841,N_29024,N_29231);
nand UO_842 (O_842,N_29588,N_29623);
nor UO_843 (O_843,N_29827,N_29810);
nor UO_844 (O_844,N_29507,N_29172);
nand UO_845 (O_845,N_29115,N_29354);
nor UO_846 (O_846,N_29986,N_29457);
or UO_847 (O_847,N_29893,N_29418);
or UO_848 (O_848,N_29781,N_29472);
nand UO_849 (O_849,N_29872,N_29262);
or UO_850 (O_850,N_29790,N_29611);
or UO_851 (O_851,N_29454,N_29523);
nor UO_852 (O_852,N_29274,N_29027);
xnor UO_853 (O_853,N_29746,N_29827);
nand UO_854 (O_854,N_29322,N_29349);
nand UO_855 (O_855,N_29695,N_29441);
and UO_856 (O_856,N_29879,N_29443);
or UO_857 (O_857,N_29603,N_29458);
nand UO_858 (O_858,N_29701,N_29080);
xnor UO_859 (O_859,N_29694,N_29438);
nand UO_860 (O_860,N_29665,N_29122);
or UO_861 (O_861,N_29465,N_29266);
xor UO_862 (O_862,N_29077,N_29473);
nand UO_863 (O_863,N_29434,N_29574);
nand UO_864 (O_864,N_29212,N_29249);
nand UO_865 (O_865,N_29481,N_29486);
or UO_866 (O_866,N_29965,N_29306);
and UO_867 (O_867,N_29771,N_29375);
xnor UO_868 (O_868,N_29151,N_29144);
nand UO_869 (O_869,N_29842,N_29528);
nand UO_870 (O_870,N_29409,N_29367);
nor UO_871 (O_871,N_29569,N_29107);
and UO_872 (O_872,N_29709,N_29004);
and UO_873 (O_873,N_29910,N_29798);
xnor UO_874 (O_874,N_29798,N_29724);
or UO_875 (O_875,N_29916,N_29336);
nor UO_876 (O_876,N_29096,N_29653);
nor UO_877 (O_877,N_29473,N_29275);
xor UO_878 (O_878,N_29183,N_29797);
and UO_879 (O_879,N_29149,N_29188);
and UO_880 (O_880,N_29761,N_29152);
nor UO_881 (O_881,N_29429,N_29860);
or UO_882 (O_882,N_29952,N_29173);
and UO_883 (O_883,N_29729,N_29991);
nor UO_884 (O_884,N_29405,N_29595);
xor UO_885 (O_885,N_29552,N_29260);
xor UO_886 (O_886,N_29286,N_29468);
or UO_887 (O_887,N_29697,N_29533);
nand UO_888 (O_888,N_29356,N_29769);
or UO_889 (O_889,N_29767,N_29206);
and UO_890 (O_890,N_29486,N_29333);
and UO_891 (O_891,N_29882,N_29892);
xor UO_892 (O_892,N_29214,N_29790);
or UO_893 (O_893,N_29663,N_29434);
nor UO_894 (O_894,N_29283,N_29214);
nand UO_895 (O_895,N_29045,N_29771);
or UO_896 (O_896,N_29973,N_29615);
or UO_897 (O_897,N_29195,N_29733);
nor UO_898 (O_898,N_29061,N_29261);
nor UO_899 (O_899,N_29194,N_29438);
and UO_900 (O_900,N_29868,N_29419);
nand UO_901 (O_901,N_29684,N_29572);
nor UO_902 (O_902,N_29845,N_29815);
xnor UO_903 (O_903,N_29311,N_29742);
or UO_904 (O_904,N_29254,N_29059);
and UO_905 (O_905,N_29015,N_29688);
and UO_906 (O_906,N_29864,N_29652);
and UO_907 (O_907,N_29260,N_29631);
xnor UO_908 (O_908,N_29017,N_29337);
xnor UO_909 (O_909,N_29694,N_29341);
xor UO_910 (O_910,N_29661,N_29277);
or UO_911 (O_911,N_29112,N_29640);
nand UO_912 (O_912,N_29748,N_29419);
nand UO_913 (O_913,N_29469,N_29210);
or UO_914 (O_914,N_29368,N_29865);
and UO_915 (O_915,N_29174,N_29822);
nand UO_916 (O_916,N_29884,N_29268);
or UO_917 (O_917,N_29336,N_29112);
nand UO_918 (O_918,N_29850,N_29114);
nor UO_919 (O_919,N_29715,N_29812);
nand UO_920 (O_920,N_29908,N_29528);
or UO_921 (O_921,N_29378,N_29301);
xor UO_922 (O_922,N_29259,N_29776);
nor UO_923 (O_923,N_29740,N_29121);
nand UO_924 (O_924,N_29689,N_29920);
and UO_925 (O_925,N_29353,N_29495);
xnor UO_926 (O_926,N_29386,N_29480);
nand UO_927 (O_927,N_29110,N_29037);
nor UO_928 (O_928,N_29627,N_29551);
or UO_929 (O_929,N_29136,N_29765);
or UO_930 (O_930,N_29425,N_29451);
nand UO_931 (O_931,N_29806,N_29435);
or UO_932 (O_932,N_29169,N_29044);
nor UO_933 (O_933,N_29195,N_29886);
and UO_934 (O_934,N_29441,N_29890);
and UO_935 (O_935,N_29262,N_29287);
nand UO_936 (O_936,N_29532,N_29939);
or UO_937 (O_937,N_29734,N_29814);
nor UO_938 (O_938,N_29101,N_29428);
xnor UO_939 (O_939,N_29288,N_29515);
nand UO_940 (O_940,N_29116,N_29708);
and UO_941 (O_941,N_29501,N_29381);
or UO_942 (O_942,N_29573,N_29787);
xor UO_943 (O_943,N_29944,N_29203);
nor UO_944 (O_944,N_29019,N_29649);
nand UO_945 (O_945,N_29742,N_29284);
nand UO_946 (O_946,N_29498,N_29922);
nand UO_947 (O_947,N_29079,N_29255);
nand UO_948 (O_948,N_29464,N_29434);
or UO_949 (O_949,N_29068,N_29178);
xor UO_950 (O_950,N_29734,N_29880);
and UO_951 (O_951,N_29713,N_29547);
nor UO_952 (O_952,N_29651,N_29703);
nor UO_953 (O_953,N_29861,N_29649);
and UO_954 (O_954,N_29433,N_29067);
nor UO_955 (O_955,N_29126,N_29967);
or UO_956 (O_956,N_29695,N_29476);
and UO_957 (O_957,N_29934,N_29910);
or UO_958 (O_958,N_29477,N_29094);
and UO_959 (O_959,N_29255,N_29681);
xnor UO_960 (O_960,N_29602,N_29728);
or UO_961 (O_961,N_29359,N_29288);
nor UO_962 (O_962,N_29728,N_29422);
xnor UO_963 (O_963,N_29635,N_29501);
nor UO_964 (O_964,N_29447,N_29859);
and UO_965 (O_965,N_29282,N_29914);
nand UO_966 (O_966,N_29465,N_29719);
or UO_967 (O_967,N_29611,N_29763);
and UO_968 (O_968,N_29387,N_29744);
or UO_969 (O_969,N_29647,N_29709);
or UO_970 (O_970,N_29364,N_29252);
nor UO_971 (O_971,N_29474,N_29579);
and UO_972 (O_972,N_29399,N_29684);
nor UO_973 (O_973,N_29618,N_29660);
or UO_974 (O_974,N_29347,N_29048);
or UO_975 (O_975,N_29173,N_29688);
nand UO_976 (O_976,N_29318,N_29212);
xor UO_977 (O_977,N_29624,N_29403);
nor UO_978 (O_978,N_29840,N_29440);
nor UO_979 (O_979,N_29089,N_29661);
nor UO_980 (O_980,N_29464,N_29193);
and UO_981 (O_981,N_29869,N_29577);
and UO_982 (O_982,N_29328,N_29702);
or UO_983 (O_983,N_29001,N_29241);
nor UO_984 (O_984,N_29263,N_29368);
nand UO_985 (O_985,N_29758,N_29983);
nand UO_986 (O_986,N_29160,N_29638);
nor UO_987 (O_987,N_29664,N_29102);
and UO_988 (O_988,N_29670,N_29983);
and UO_989 (O_989,N_29941,N_29658);
or UO_990 (O_990,N_29384,N_29860);
nand UO_991 (O_991,N_29049,N_29890);
nor UO_992 (O_992,N_29957,N_29097);
or UO_993 (O_993,N_29854,N_29944);
xor UO_994 (O_994,N_29241,N_29599);
xnor UO_995 (O_995,N_29610,N_29155);
nand UO_996 (O_996,N_29713,N_29064);
xnor UO_997 (O_997,N_29398,N_29675);
or UO_998 (O_998,N_29844,N_29668);
xor UO_999 (O_999,N_29935,N_29340);
nor UO_1000 (O_1000,N_29440,N_29522);
and UO_1001 (O_1001,N_29896,N_29648);
nand UO_1002 (O_1002,N_29108,N_29201);
nand UO_1003 (O_1003,N_29384,N_29378);
and UO_1004 (O_1004,N_29494,N_29469);
nand UO_1005 (O_1005,N_29474,N_29260);
or UO_1006 (O_1006,N_29105,N_29886);
nand UO_1007 (O_1007,N_29785,N_29694);
xnor UO_1008 (O_1008,N_29438,N_29272);
or UO_1009 (O_1009,N_29676,N_29748);
nor UO_1010 (O_1010,N_29815,N_29826);
and UO_1011 (O_1011,N_29726,N_29840);
nor UO_1012 (O_1012,N_29065,N_29789);
xor UO_1013 (O_1013,N_29637,N_29894);
or UO_1014 (O_1014,N_29643,N_29298);
and UO_1015 (O_1015,N_29589,N_29917);
xnor UO_1016 (O_1016,N_29295,N_29791);
nand UO_1017 (O_1017,N_29860,N_29739);
or UO_1018 (O_1018,N_29975,N_29100);
or UO_1019 (O_1019,N_29031,N_29183);
and UO_1020 (O_1020,N_29915,N_29737);
nand UO_1021 (O_1021,N_29494,N_29746);
nor UO_1022 (O_1022,N_29357,N_29666);
nand UO_1023 (O_1023,N_29979,N_29730);
nor UO_1024 (O_1024,N_29431,N_29973);
nand UO_1025 (O_1025,N_29944,N_29751);
and UO_1026 (O_1026,N_29285,N_29092);
xor UO_1027 (O_1027,N_29535,N_29950);
nand UO_1028 (O_1028,N_29471,N_29412);
or UO_1029 (O_1029,N_29792,N_29737);
and UO_1030 (O_1030,N_29849,N_29431);
xnor UO_1031 (O_1031,N_29666,N_29785);
or UO_1032 (O_1032,N_29776,N_29815);
xnor UO_1033 (O_1033,N_29348,N_29197);
nand UO_1034 (O_1034,N_29751,N_29054);
nand UO_1035 (O_1035,N_29357,N_29496);
nor UO_1036 (O_1036,N_29792,N_29003);
or UO_1037 (O_1037,N_29914,N_29806);
and UO_1038 (O_1038,N_29313,N_29460);
or UO_1039 (O_1039,N_29499,N_29759);
and UO_1040 (O_1040,N_29498,N_29062);
or UO_1041 (O_1041,N_29539,N_29130);
nor UO_1042 (O_1042,N_29314,N_29377);
or UO_1043 (O_1043,N_29478,N_29408);
and UO_1044 (O_1044,N_29605,N_29408);
and UO_1045 (O_1045,N_29490,N_29368);
or UO_1046 (O_1046,N_29013,N_29823);
and UO_1047 (O_1047,N_29916,N_29994);
nand UO_1048 (O_1048,N_29938,N_29821);
or UO_1049 (O_1049,N_29589,N_29303);
nand UO_1050 (O_1050,N_29963,N_29536);
nor UO_1051 (O_1051,N_29880,N_29802);
xor UO_1052 (O_1052,N_29588,N_29404);
or UO_1053 (O_1053,N_29989,N_29326);
nor UO_1054 (O_1054,N_29663,N_29126);
or UO_1055 (O_1055,N_29502,N_29122);
and UO_1056 (O_1056,N_29043,N_29872);
nor UO_1057 (O_1057,N_29126,N_29926);
nand UO_1058 (O_1058,N_29338,N_29588);
and UO_1059 (O_1059,N_29036,N_29379);
and UO_1060 (O_1060,N_29056,N_29840);
xnor UO_1061 (O_1061,N_29175,N_29225);
nor UO_1062 (O_1062,N_29875,N_29007);
nand UO_1063 (O_1063,N_29612,N_29996);
and UO_1064 (O_1064,N_29940,N_29772);
nor UO_1065 (O_1065,N_29505,N_29144);
and UO_1066 (O_1066,N_29807,N_29072);
and UO_1067 (O_1067,N_29865,N_29032);
or UO_1068 (O_1068,N_29251,N_29659);
and UO_1069 (O_1069,N_29100,N_29171);
and UO_1070 (O_1070,N_29129,N_29696);
or UO_1071 (O_1071,N_29256,N_29056);
nor UO_1072 (O_1072,N_29146,N_29703);
or UO_1073 (O_1073,N_29732,N_29486);
or UO_1074 (O_1074,N_29124,N_29554);
nor UO_1075 (O_1075,N_29201,N_29479);
or UO_1076 (O_1076,N_29611,N_29715);
and UO_1077 (O_1077,N_29774,N_29802);
or UO_1078 (O_1078,N_29551,N_29755);
xor UO_1079 (O_1079,N_29999,N_29530);
or UO_1080 (O_1080,N_29141,N_29991);
nand UO_1081 (O_1081,N_29157,N_29539);
nand UO_1082 (O_1082,N_29772,N_29525);
nor UO_1083 (O_1083,N_29494,N_29832);
or UO_1084 (O_1084,N_29956,N_29160);
and UO_1085 (O_1085,N_29499,N_29699);
or UO_1086 (O_1086,N_29914,N_29369);
nor UO_1087 (O_1087,N_29155,N_29379);
and UO_1088 (O_1088,N_29652,N_29139);
or UO_1089 (O_1089,N_29515,N_29240);
or UO_1090 (O_1090,N_29832,N_29416);
or UO_1091 (O_1091,N_29804,N_29176);
or UO_1092 (O_1092,N_29759,N_29207);
and UO_1093 (O_1093,N_29993,N_29732);
nor UO_1094 (O_1094,N_29687,N_29420);
nand UO_1095 (O_1095,N_29408,N_29804);
or UO_1096 (O_1096,N_29345,N_29521);
or UO_1097 (O_1097,N_29745,N_29555);
xor UO_1098 (O_1098,N_29654,N_29611);
and UO_1099 (O_1099,N_29399,N_29774);
nand UO_1100 (O_1100,N_29875,N_29677);
nor UO_1101 (O_1101,N_29541,N_29902);
nand UO_1102 (O_1102,N_29722,N_29246);
nand UO_1103 (O_1103,N_29255,N_29755);
nand UO_1104 (O_1104,N_29852,N_29094);
or UO_1105 (O_1105,N_29483,N_29046);
xnor UO_1106 (O_1106,N_29329,N_29825);
or UO_1107 (O_1107,N_29172,N_29408);
nor UO_1108 (O_1108,N_29723,N_29434);
nor UO_1109 (O_1109,N_29328,N_29852);
and UO_1110 (O_1110,N_29949,N_29216);
nand UO_1111 (O_1111,N_29913,N_29596);
nand UO_1112 (O_1112,N_29054,N_29348);
nor UO_1113 (O_1113,N_29115,N_29616);
or UO_1114 (O_1114,N_29459,N_29511);
and UO_1115 (O_1115,N_29418,N_29535);
nor UO_1116 (O_1116,N_29293,N_29299);
and UO_1117 (O_1117,N_29113,N_29973);
or UO_1118 (O_1118,N_29854,N_29059);
nor UO_1119 (O_1119,N_29633,N_29152);
xor UO_1120 (O_1120,N_29994,N_29245);
nand UO_1121 (O_1121,N_29459,N_29864);
and UO_1122 (O_1122,N_29107,N_29575);
and UO_1123 (O_1123,N_29723,N_29134);
nor UO_1124 (O_1124,N_29141,N_29493);
nand UO_1125 (O_1125,N_29058,N_29410);
nand UO_1126 (O_1126,N_29050,N_29659);
and UO_1127 (O_1127,N_29102,N_29148);
or UO_1128 (O_1128,N_29535,N_29685);
nor UO_1129 (O_1129,N_29188,N_29832);
nor UO_1130 (O_1130,N_29341,N_29973);
and UO_1131 (O_1131,N_29031,N_29202);
or UO_1132 (O_1132,N_29419,N_29725);
nand UO_1133 (O_1133,N_29743,N_29331);
or UO_1134 (O_1134,N_29624,N_29539);
xor UO_1135 (O_1135,N_29594,N_29304);
xnor UO_1136 (O_1136,N_29840,N_29323);
nor UO_1137 (O_1137,N_29346,N_29579);
xor UO_1138 (O_1138,N_29070,N_29208);
and UO_1139 (O_1139,N_29955,N_29984);
xnor UO_1140 (O_1140,N_29803,N_29632);
nor UO_1141 (O_1141,N_29319,N_29128);
nor UO_1142 (O_1142,N_29771,N_29195);
and UO_1143 (O_1143,N_29086,N_29180);
xor UO_1144 (O_1144,N_29786,N_29245);
or UO_1145 (O_1145,N_29052,N_29927);
and UO_1146 (O_1146,N_29602,N_29573);
or UO_1147 (O_1147,N_29906,N_29129);
nand UO_1148 (O_1148,N_29717,N_29782);
or UO_1149 (O_1149,N_29490,N_29844);
and UO_1150 (O_1150,N_29035,N_29555);
and UO_1151 (O_1151,N_29981,N_29643);
or UO_1152 (O_1152,N_29245,N_29007);
nor UO_1153 (O_1153,N_29442,N_29319);
xor UO_1154 (O_1154,N_29016,N_29640);
or UO_1155 (O_1155,N_29625,N_29774);
and UO_1156 (O_1156,N_29911,N_29812);
nor UO_1157 (O_1157,N_29345,N_29503);
nand UO_1158 (O_1158,N_29762,N_29371);
or UO_1159 (O_1159,N_29634,N_29999);
or UO_1160 (O_1160,N_29644,N_29473);
or UO_1161 (O_1161,N_29222,N_29221);
xor UO_1162 (O_1162,N_29132,N_29030);
nor UO_1163 (O_1163,N_29513,N_29646);
nor UO_1164 (O_1164,N_29938,N_29494);
and UO_1165 (O_1165,N_29466,N_29805);
or UO_1166 (O_1166,N_29808,N_29459);
or UO_1167 (O_1167,N_29618,N_29063);
xor UO_1168 (O_1168,N_29450,N_29991);
or UO_1169 (O_1169,N_29547,N_29201);
xor UO_1170 (O_1170,N_29239,N_29507);
xor UO_1171 (O_1171,N_29241,N_29140);
nand UO_1172 (O_1172,N_29043,N_29409);
xnor UO_1173 (O_1173,N_29690,N_29464);
and UO_1174 (O_1174,N_29704,N_29428);
nor UO_1175 (O_1175,N_29350,N_29087);
nor UO_1176 (O_1176,N_29941,N_29184);
xnor UO_1177 (O_1177,N_29622,N_29730);
xor UO_1178 (O_1178,N_29189,N_29343);
xor UO_1179 (O_1179,N_29457,N_29373);
xnor UO_1180 (O_1180,N_29069,N_29682);
or UO_1181 (O_1181,N_29429,N_29353);
nand UO_1182 (O_1182,N_29175,N_29116);
and UO_1183 (O_1183,N_29197,N_29030);
xnor UO_1184 (O_1184,N_29579,N_29125);
nor UO_1185 (O_1185,N_29111,N_29148);
xor UO_1186 (O_1186,N_29458,N_29307);
nor UO_1187 (O_1187,N_29050,N_29150);
and UO_1188 (O_1188,N_29453,N_29874);
xor UO_1189 (O_1189,N_29884,N_29274);
xnor UO_1190 (O_1190,N_29149,N_29020);
nor UO_1191 (O_1191,N_29785,N_29349);
xor UO_1192 (O_1192,N_29115,N_29850);
nor UO_1193 (O_1193,N_29852,N_29678);
nor UO_1194 (O_1194,N_29992,N_29113);
and UO_1195 (O_1195,N_29861,N_29951);
xnor UO_1196 (O_1196,N_29303,N_29671);
or UO_1197 (O_1197,N_29428,N_29418);
xnor UO_1198 (O_1198,N_29720,N_29871);
nor UO_1199 (O_1199,N_29364,N_29830);
nand UO_1200 (O_1200,N_29451,N_29903);
or UO_1201 (O_1201,N_29029,N_29682);
nor UO_1202 (O_1202,N_29390,N_29461);
nand UO_1203 (O_1203,N_29569,N_29233);
nor UO_1204 (O_1204,N_29117,N_29083);
or UO_1205 (O_1205,N_29468,N_29727);
and UO_1206 (O_1206,N_29032,N_29144);
nor UO_1207 (O_1207,N_29008,N_29970);
or UO_1208 (O_1208,N_29720,N_29815);
nand UO_1209 (O_1209,N_29750,N_29242);
nand UO_1210 (O_1210,N_29467,N_29046);
and UO_1211 (O_1211,N_29222,N_29400);
and UO_1212 (O_1212,N_29864,N_29124);
nand UO_1213 (O_1213,N_29536,N_29677);
nand UO_1214 (O_1214,N_29076,N_29046);
nand UO_1215 (O_1215,N_29649,N_29486);
or UO_1216 (O_1216,N_29495,N_29666);
or UO_1217 (O_1217,N_29326,N_29196);
or UO_1218 (O_1218,N_29493,N_29487);
nor UO_1219 (O_1219,N_29034,N_29878);
nand UO_1220 (O_1220,N_29872,N_29630);
xnor UO_1221 (O_1221,N_29602,N_29996);
xnor UO_1222 (O_1222,N_29857,N_29346);
or UO_1223 (O_1223,N_29348,N_29552);
nand UO_1224 (O_1224,N_29564,N_29571);
and UO_1225 (O_1225,N_29554,N_29674);
nand UO_1226 (O_1226,N_29892,N_29439);
and UO_1227 (O_1227,N_29926,N_29487);
nand UO_1228 (O_1228,N_29747,N_29997);
nand UO_1229 (O_1229,N_29597,N_29913);
nand UO_1230 (O_1230,N_29114,N_29419);
nor UO_1231 (O_1231,N_29919,N_29702);
xor UO_1232 (O_1232,N_29324,N_29687);
nand UO_1233 (O_1233,N_29538,N_29836);
xnor UO_1234 (O_1234,N_29591,N_29058);
and UO_1235 (O_1235,N_29760,N_29320);
and UO_1236 (O_1236,N_29460,N_29843);
or UO_1237 (O_1237,N_29496,N_29130);
nor UO_1238 (O_1238,N_29678,N_29118);
xor UO_1239 (O_1239,N_29210,N_29283);
and UO_1240 (O_1240,N_29942,N_29213);
nand UO_1241 (O_1241,N_29929,N_29917);
or UO_1242 (O_1242,N_29127,N_29049);
nor UO_1243 (O_1243,N_29603,N_29719);
nor UO_1244 (O_1244,N_29582,N_29048);
nand UO_1245 (O_1245,N_29661,N_29097);
or UO_1246 (O_1246,N_29820,N_29871);
nand UO_1247 (O_1247,N_29511,N_29787);
nand UO_1248 (O_1248,N_29918,N_29791);
nor UO_1249 (O_1249,N_29391,N_29811);
nand UO_1250 (O_1250,N_29619,N_29171);
nor UO_1251 (O_1251,N_29363,N_29913);
nor UO_1252 (O_1252,N_29826,N_29382);
and UO_1253 (O_1253,N_29939,N_29166);
nand UO_1254 (O_1254,N_29798,N_29087);
nor UO_1255 (O_1255,N_29100,N_29731);
or UO_1256 (O_1256,N_29211,N_29086);
or UO_1257 (O_1257,N_29185,N_29588);
nand UO_1258 (O_1258,N_29794,N_29568);
xor UO_1259 (O_1259,N_29345,N_29459);
xor UO_1260 (O_1260,N_29216,N_29231);
and UO_1261 (O_1261,N_29034,N_29631);
nor UO_1262 (O_1262,N_29233,N_29392);
nor UO_1263 (O_1263,N_29451,N_29714);
xnor UO_1264 (O_1264,N_29341,N_29069);
nor UO_1265 (O_1265,N_29602,N_29900);
nand UO_1266 (O_1266,N_29247,N_29900);
or UO_1267 (O_1267,N_29716,N_29750);
xor UO_1268 (O_1268,N_29234,N_29660);
nor UO_1269 (O_1269,N_29277,N_29680);
nor UO_1270 (O_1270,N_29132,N_29396);
xor UO_1271 (O_1271,N_29405,N_29768);
or UO_1272 (O_1272,N_29577,N_29884);
nor UO_1273 (O_1273,N_29259,N_29287);
nand UO_1274 (O_1274,N_29404,N_29849);
nand UO_1275 (O_1275,N_29063,N_29447);
or UO_1276 (O_1276,N_29246,N_29149);
xnor UO_1277 (O_1277,N_29766,N_29865);
and UO_1278 (O_1278,N_29876,N_29511);
or UO_1279 (O_1279,N_29949,N_29645);
nand UO_1280 (O_1280,N_29993,N_29047);
or UO_1281 (O_1281,N_29180,N_29055);
xor UO_1282 (O_1282,N_29974,N_29206);
or UO_1283 (O_1283,N_29858,N_29735);
nor UO_1284 (O_1284,N_29643,N_29932);
nor UO_1285 (O_1285,N_29433,N_29241);
nor UO_1286 (O_1286,N_29385,N_29983);
or UO_1287 (O_1287,N_29029,N_29339);
and UO_1288 (O_1288,N_29984,N_29139);
or UO_1289 (O_1289,N_29249,N_29486);
nor UO_1290 (O_1290,N_29264,N_29431);
or UO_1291 (O_1291,N_29287,N_29279);
nand UO_1292 (O_1292,N_29639,N_29275);
nor UO_1293 (O_1293,N_29117,N_29594);
and UO_1294 (O_1294,N_29448,N_29535);
and UO_1295 (O_1295,N_29871,N_29984);
and UO_1296 (O_1296,N_29450,N_29805);
and UO_1297 (O_1297,N_29897,N_29145);
nor UO_1298 (O_1298,N_29409,N_29741);
and UO_1299 (O_1299,N_29135,N_29445);
or UO_1300 (O_1300,N_29205,N_29889);
nor UO_1301 (O_1301,N_29966,N_29651);
and UO_1302 (O_1302,N_29125,N_29491);
nor UO_1303 (O_1303,N_29278,N_29429);
nand UO_1304 (O_1304,N_29929,N_29579);
nand UO_1305 (O_1305,N_29976,N_29084);
and UO_1306 (O_1306,N_29098,N_29354);
nand UO_1307 (O_1307,N_29088,N_29085);
nand UO_1308 (O_1308,N_29278,N_29508);
nor UO_1309 (O_1309,N_29619,N_29461);
nand UO_1310 (O_1310,N_29131,N_29101);
nand UO_1311 (O_1311,N_29510,N_29958);
nor UO_1312 (O_1312,N_29576,N_29017);
and UO_1313 (O_1313,N_29557,N_29145);
or UO_1314 (O_1314,N_29364,N_29758);
xor UO_1315 (O_1315,N_29838,N_29117);
and UO_1316 (O_1316,N_29439,N_29630);
and UO_1317 (O_1317,N_29673,N_29792);
nor UO_1318 (O_1318,N_29229,N_29966);
and UO_1319 (O_1319,N_29551,N_29393);
nor UO_1320 (O_1320,N_29979,N_29128);
or UO_1321 (O_1321,N_29158,N_29225);
nand UO_1322 (O_1322,N_29720,N_29232);
and UO_1323 (O_1323,N_29286,N_29509);
nor UO_1324 (O_1324,N_29912,N_29744);
nand UO_1325 (O_1325,N_29936,N_29790);
nand UO_1326 (O_1326,N_29264,N_29850);
nand UO_1327 (O_1327,N_29364,N_29727);
or UO_1328 (O_1328,N_29275,N_29513);
or UO_1329 (O_1329,N_29451,N_29839);
nand UO_1330 (O_1330,N_29975,N_29780);
nor UO_1331 (O_1331,N_29163,N_29027);
xnor UO_1332 (O_1332,N_29162,N_29019);
or UO_1333 (O_1333,N_29147,N_29961);
and UO_1334 (O_1334,N_29321,N_29634);
nand UO_1335 (O_1335,N_29804,N_29429);
and UO_1336 (O_1336,N_29407,N_29718);
or UO_1337 (O_1337,N_29755,N_29259);
xor UO_1338 (O_1338,N_29393,N_29240);
nor UO_1339 (O_1339,N_29822,N_29440);
nor UO_1340 (O_1340,N_29490,N_29617);
or UO_1341 (O_1341,N_29731,N_29428);
and UO_1342 (O_1342,N_29288,N_29167);
nand UO_1343 (O_1343,N_29757,N_29943);
and UO_1344 (O_1344,N_29135,N_29272);
and UO_1345 (O_1345,N_29483,N_29194);
nor UO_1346 (O_1346,N_29159,N_29818);
and UO_1347 (O_1347,N_29407,N_29047);
nand UO_1348 (O_1348,N_29418,N_29050);
nand UO_1349 (O_1349,N_29263,N_29178);
nand UO_1350 (O_1350,N_29843,N_29695);
and UO_1351 (O_1351,N_29831,N_29196);
nand UO_1352 (O_1352,N_29123,N_29328);
and UO_1353 (O_1353,N_29223,N_29202);
or UO_1354 (O_1354,N_29547,N_29520);
xnor UO_1355 (O_1355,N_29876,N_29968);
nor UO_1356 (O_1356,N_29691,N_29847);
or UO_1357 (O_1357,N_29950,N_29539);
nand UO_1358 (O_1358,N_29228,N_29930);
xor UO_1359 (O_1359,N_29411,N_29689);
nand UO_1360 (O_1360,N_29512,N_29865);
and UO_1361 (O_1361,N_29587,N_29999);
xnor UO_1362 (O_1362,N_29095,N_29439);
nor UO_1363 (O_1363,N_29083,N_29523);
nor UO_1364 (O_1364,N_29869,N_29249);
nor UO_1365 (O_1365,N_29918,N_29470);
or UO_1366 (O_1366,N_29726,N_29709);
nor UO_1367 (O_1367,N_29202,N_29738);
xnor UO_1368 (O_1368,N_29329,N_29977);
xnor UO_1369 (O_1369,N_29804,N_29944);
nand UO_1370 (O_1370,N_29541,N_29015);
or UO_1371 (O_1371,N_29628,N_29582);
or UO_1372 (O_1372,N_29821,N_29357);
or UO_1373 (O_1373,N_29890,N_29297);
nor UO_1374 (O_1374,N_29009,N_29680);
xnor UO_1375 (O_1375,N_29010,N_29400);
xnor UO_1376 (O_1376,N_29455,N_29579);
nor UO_1377 (O_1377,N_29394,N_29755);
nand UO_1378 (O_1378,N_29557,N_29443);
xor UO_1379 (O_1379,N_29632,N_29174);
nand UO_1380 (O_1380,N_29591,N_29373);
or UO_1381 (O_1381,N_29268,N_29212);
nor UO_1382 (O_1382,N_29694,N_29861);
xor UO_1383 (O_1383,N_29783,N_29645);
and UO_1384 (O_1384,N_29868,N_29899);
xor UO_1385 (O_1385,N_29674,N_29742);
or UO_1386 (O_1386,N_29586,N_29107);
xnor UO_1387 (O_1387,N_29154,N_29039);
and UO_1388 (O_1388,N_29486,N_29378);
and UO_1389 (O_1389,N_29819,N_29203);
xnor UO_1390 (O_1390,N_29090,N_29660);
and UO_1391 (O_1391,N_29081,N_29566);
xor UO_1392 (O_1392,N_29625,N_29383);
nand UO_1393 (O_1393,N_29152,N_29662);
or UO_1394 (O_1394,N_29949,N_29036);
or UO_1395 (O_1395,N_29829,N_29196);
or UO_1396 (O_1396,N_29555,N_29235);
nand UO_1397 (O_1397,N_29072,N_29271);
or UO_1398 (O_1398,N_29268,N_29164);
or UO_1399 (O_1399,N_29888,N_29528);
and UO_1400 (O_1400,N_29210,N_29196);
nor UO_1401 (O_1401,N_29871,N_29452);
nand UO_1402 (O_1402,N_29692,N_29574);
nor UO_1403 (O_1403,N_29208,N_29569);
xnor UO_1404 (O_1404,N_29643,N_29286);
nor UO_1405 (O_1405,N_29805,N_29695);
nand UO_1406 (O_1406,N_29154,N_29779);
or UO_1407 (O_1407,N_29872,N_29635);
xor UO_1408 (O_1408,N_29925,N_29878);
nand UO_1409 (O_1409,N_29758,N_29397);
xor UO_1410 (O_1410,N_29882,N_29740);
nor UO_1411 (O_1411,N_29334,N_29685);
nor UO_1412 (O_1412,N_29984,N_29755);
or UO_1413 (O_1413,N_29305,N_29153);
and UO_1414 (O_1414,N_29843,N_29936);
xor UO_1415 (O_1415,N_29523,N_29591);
nand UO_1416 (O_1416,N_29591,N_29704);
xor UO_1417 (O_1417,N_29757,N_29736);
nand UO_1418 (O_1418,N_29562,N_29825);
nor UO_1419 (O_1419,N_29830,N_29420);
and UO_1420 (O_1420,N_29233,N_29847);
nor UO_1421 (O_1421,N_29709,N_29572);
nand UO_1422 (O_1422,N_29485,N_29801);
xor UO_1423 (O_1423,N_29737,N_29693);
nand UO_1424 (O_1424,N_29381,N_29010);
and UO_1425 (O_1425,N_29206,N_29383);
or UO_1426 (O_1426,N_29894,N_29688);
xnor UO_1427 (O_1427,N_29970,N_29605);
or UO_1428 (O_1428,N_29536,N_29518);
nor UO_1429 (O_1429,N_29720,N_29211);
xnor UO_1430 (O_1430,N_29705,N_29863);
and UO_1431 (O_1431,N_29470,N_29017);
and UO_1432 (O_1432,N_29740,N_29781);
nor UO_1433 (O_1433,N_29753,N_29632);
nand UO_1434 (O_1434,N_29245,N_29850);
nand UO_1435 (O_1435,N_29256,N_29000);
nand UO_1436 (O_1436,N_29209,N_29948);
and UO_1437 (O_1437,N_29159,N_29541);
nand UO_1438 (O_1438,N_29740,N_29869);
xnor UO_1439 (O_1439,N_29643,N_29072);
nand UO_1440 (O_1440,N_29936,N_29489);
xnor UO_1441 (O_1441,N_29269,N_29897);
and UO_1442 (O_1442,N_29560,N_29601);
and UO_1443 (O_1443,N_29271,N_29410);
nand UO_1444 (O_1444,N_29343,N_29355);
or UO_1445 (O_1445,N_29548,N_29663);
nor UO_1446 (O_1446,N_29021,N_29164);
nor UO_1447 (O_1447,N_29902,N_29747);
or UO_1448 (O_1448,N_29680,N_29166);
xnor UO_1449 (O_1449,N_29694,N_29718);
nor UO_1450 (O_1450,N_29742,N_29892);
and UO_1451 (O_1451,N_29093,N_29711);
nand UO_1452 (O_1452,N_29780,N_29416);
nor UO_1453 (O_1453,N_29857,N_29614);
or UO_1454 (O_1454,N_29876,N_29449);
and UO_1455 (O_1455,N_29447,N_29277);
nor UO_1456 (O_1456,N_29150,N_29838);
or UO_1457 (O_1457,N_29056,N_29525);
nand UO_1458 (O_1458,N_29919,N_29413);
xnor UO_1459 (O_1459,N_29092,N_29168);
or UO_1460 (O_1460,N_29385,N_29503);
or UO_1461 (O_1461,N_29553,N_29500);
xnor UO_1462 (O_1462,N_29127,N_29608);
nor UO_1463 (O_1463,N_29159,N_29328);
nor UO_1464 (O_1464,N_29103,N_29386);
or UO_1465 (O_1465,N_29941,N_29958);
xnor UO_1466 (O_1466,N_29402,N_29992);
or UO_1467 (O_1467,N_29129,N_29014);
nand UO_1468 (O_1468,N_29498,N_29874);
and UO_1469 (O_1469,N_29043,N_29482);
xnor UO_1470 (O_1470,N_29624,N_29772);
nor UO_1471 (O_1471,N_29578,N_29021);
xor UO_1472 (O_1472,N_29478,N_29145);
and UO_1473 (O_1473,N_29545,N_29966);
nor UO_1474 (O_1474,N_29179,N_29376);
xnor UO_1475 (O_1475,N_29110,N_29994);
xor UO_1476 (O_1476,N_29181,N_29728);
nor UO_1477 (O_1477,N_29420,N_29765);
xnor UO_1478 (O_1478,N_29458,N_29534);
nand UO_1479 (O_1479,N_29779,N_29669);
xor UO_1480 (O_1480,N_29553,N_29914);
xnor UO_1481 (O_1481,N_29111,N_29114);
and UO_1482 (O_1482,N_29586,N_29785);
nor UO_1483 (O_1483,N_29092,N_29020);
and UO_1484 (O_1484,N_29098,N_29453);
or UO_1485 (O_1485,N_29231,N_29585);
nor UO_1486 (O_1486,N_29904,N_29128);
xnor UO_1487 (O_1487,N_29232,N_29231);
xor UO_1488 (O_1488,N_29015,N_29086);
nand UO_1489 (O_1489,N_29352,N_29356);
xnor UO_1490 (O_1490,N_29359,N_29543);
and UO_1491 (O_1491,N_29044,N_29013);
nor UO_1492 (O_1492,N_29804,N_29307);
and UO_1493 (O_1493,N_29991,N_29725);
nor UO_1494 (O_1494,N_29147,N_29393);
and UO_1495 (O_1495,N_29763,N_29383);
and UO_1496 (O_1496,N_29658,N_29700);
and UO_1497 (O_1497,N_29791,N_29605);
or UO_1498 (O_1498,N_29478,N_29284);
nand UO_1499 (O_1499,N_29167,N_29344);
xor UO_1500 (O_1500,N_29046,N_29252);
or UO_1501 (O_1501,N_29295,N_29433);
and UO_1502 (O_1502,N_29968,N_29104);
and UO_1503 (O_1503,N_29218,N_29473);
or UO_1504 (O_1504,N_29109,N_29346);
nor UO_1505 (O_1505,N_29537,N_29285);
and UO_1506 (O_1506,N_29586,N_29242);
and UO_1507 (O_1507,N_29614,N_29358);
nor UO_1508 (O_1508,N_29579,N_29905);
nand UO_1509 (O_1509,N_29323,N_29756);
nand UO_1510 (O_1510,N_29967,N_29782);
xnor UO_1511 (O_1511,N_29110,N_29777);
xnor UO_1512 (O_1512,N_29583,N_29802);
and UO_1513 (O_1513,N_29140,N_29203);
and UO_1514 (O_1514,N_29887,N_29478);
or UO_1515 (O_1515,N_29379,N_29115);
and UO_1516 (O_1516,N_29199,N_29521);
nand UO_1517 (O_1517,N_29134,N_29327);
xnor UO_1518 (O_1518,N_29501,N_29596);
xnor UO_1519 (O_1519,N_29752,N_29519);
and UO_1520 (O_1520,N_29923,N_29619);
xor UO_1521 (O_1521,N_29970,N_29266);
nor UO_1522 (O_1522,N_29332,N_29225);
nor UO_1523 (O_1523,N_29277,N_29735);
xnor UO_1524 (O_1524,N_29586,N_29022);
or UO_1525 (O_1525,N_29992,N_29601);
or UO_1526 (O_1526,N_29640,N_29948);
nand UO_1527 (O_1527,N_29290,N_29870);
xor UO_1528 (O_1528,N_29079,N_29604);
nand UO_1529 (O_1529,N_29095,N_29027);
and UO_1530 (O_1530,N_29684,N_29839);
xor UO_1531 (O_1531,N_29367,N_29410);
nand UO_1532 (O_1532,N_29982,N_29968);
nor UO_1533 (O_1533,N_29092,N_29019);
or UO_1534 (O_1534,N_29894,N_29128);
xnor UO_1535 (O_1535,N_29783,N_29183);
nor UO_1536 (O_1536,N_29356,N_29969);
and UO_1537 (O_1537,N_29903,N_29847);
and UO_1538 (O_1538,N_29550,N_29658);
and UO_1539 (O_1539,N_29500,N_29322);
and UO_1540 (O_1540,N_29742,N_29379);
and UO_1541 (O_1541,N_29442,N_29932);
nor UO_1542 (O_1542,N_29247,N_29609);
and UO_1543 (O_1543,N_29431,N_29627);
or UO_1544 (O_1544,N_29981,N_29159);
xnor UO_1545 (O_1545,N_29456,N_29500);
and UO_1546 (O_1546,N_29463,N_29211);
nand UO_1547 (O_1547,N_29775,N_29822);
nor UO_1548 (O_1548,N_29412,N_29078);
xor UO_1549 (O_1549,N_29618,N_29105);
nor UO_1550 (O_1550,N_29739,N_29529);
nor UO_1551 (O_1551,N_29784,N_29823);
nor UO_1552 (O_1552,N_29850,N_29473);
or UO_1553 (O_1553,N_29497,N_29958);
nand UO_1554 (O_1554,N_29130,N_29439);
xor UO_1555 (O_1555,N_29155,N_29872);
and UO_1556 (O_1556,N_29850,N_29221);
and UO_1557 (O_1557,N_29878,N_29905);
xnor UO_1558 (O_1558,N_29718,N_29707);
nand UO_1559 (O_1559,N_29210,N_29581);
nand UO_1560 (O_1560,N_29154,N_29657);
nor UO_1561 (O_1561,N_29124,N_29903);
or UO_1562 (O_1562,N_29109,N_29131);
xor UO_1563 (O_1563,N_29239,N_29380);
and UO_1564 (O_1564,N_29724,N_29105);
xor UO_1565 (O_1565,N_29071,N_29670);
or UO_1566 (O_1566,N_29455,N_29048);
xnor UO_1567 (O_1567,N_29194,N_29129);
and UO_1568 (O_1568,N_29836,N_29834);
xor UO_1569 (O_1569,N_29655,N_29714);
xnor UO_1570 (O_1570,N_29324,N_29298);
or UO_1571 (O_1571,N_29394,N_29127);
nor UO_1572 (O_1572,N_29570,N_29789);
xor UO_1573 (O_1573,N_29304,N_29808);
xnor UO_1574 (O_1574,N_29367,N_29504);
and UO_1575 (O_1575,N_29585,N_29964);
and UO_1576 (O_1576,N_29273,N_29551);
xnor UO_1577 (O_1577,N_29247,N_29997);
nor UO_1578 (O_1578,N_29850,N_29276);
xnor UO_1579 (O_1579,N_29354,N_29652);
and UO_1580 (O_1580,N_29087,N_29128);
and UO_1581 (O_1581,N_29104,N_29566);
nor UO_1582 (O_1582,N_29262,N_29621);
or UO_1583 (O_1583,N_29090,N_29524);
xor UO_1584 (O_1584,N_29784,N_29124);
and UO_1585 (O_1585,N_29454,N_29848);
or UO_1586 (O_1586,N_29170,N_29188);
or UO_1587 (O_1587,N_29843,N_29553);
and UO_1588 (O_1588,N_29331,N_29613);
nand UO_1589 (O_1589,N_29836,N_29744);
or UO_1590 (O_1590,N_29029,N_29960);
and UO_1591 (O_1591,N_29452,N_29802);
and UO_1592 (O_1592,N_29429,N_29974);
nand UO_1593 (O_1593,N_29511,N_29399);
and UO_1594 (O_1594,N_29295,N_29566);
nor UO_1595 (O_1595,N_29071,N_29813);
xor UO_1596 (O_1596,N_29272,N_29114);
nand UO_1597 (O_1597,N_29726,N_29041);
nand UO_1598 (O_1598,N_29307,N_29099);
or UO_1599 (O_1599,N_29008,N_29757);
and UO_1600 (O_1600,N_29707,N_29105);
nor UO_1601 (O_1601,N_29221,N_29068);
xor UO_1602 (O_1602,N_29379,N_29156);
and UO_1603 (O_1603,N_29870,N_29362);
xnor UO_1604 (O_1604,N_29746,N_29243);
nand UO_1605 (O_1605,N_29809,N_29507);
xor UO_1606 (O_1606,N_29967,N_29119);
nor UO_1607 (O_1607,N_29038,N_29534);
and UO_1608 (O_1608,N_29419,N_29426);
and UO_1609 (O_1609,N_29765,N_29296);
and UO_1610 (O_1610,N_29760,N_29357);
nand UO_1611 (O_1611,N_29596,N_29789);
and UO_1612 (O_1612,N_29181,N_29127);
or UO_1613 (O_1613,N_29352,N_29663);
nor UO_1614 (O_1614,N_29808,N_29676);
or UO_1615 (O_1615,N_29176,N_29502);
xor UO_1616 (O_1616,N_29181,N_29096);
nor UO_1617 (O_1617,N_29903,N_29716);
nand UO_1618 (O_1618,N_29679,N_29618);
and UO_1619 (O_1619,N_29869,N_29829);
xnor UO_1620 (O_1620,N_29675,N_29730);
xor UO_1621 (O_1621,N_29994,N_29745);
nand UO_1622 (O_1622,N_29578,N_29181);
or UO_1623 (O_1623,N_29408,N_29633);
xnor UO_1624 (O_1624,N_29520,N_29776);
and UO_1625 (O_1625,N_29925,N_29637);
and UO_1626 (O_1626,N_29180,N_29265);
xor UO_1627 (O_1627,N_29454,N_29489);
xnor UO_1628 (O_1628,N_29022,N_29776);
or UO_1629 (O_1629,N_29844,N_29185);
and UO_1630 (O_1630,N_29012,N_29122);
xnor UO_1631 (O_1631,N_29988,N_29152);
nand UO_1632 (O_1632,N_29276,N_29190);
nor UO_1633 (O_1633,N_29716,N_29819);
nand UO_1634 (O_1634,N_29243,N_29493);
nand UO_1635 (O_1635,N_29845,N_29654);
or UO_1636 (O_1636,N_29663,N_29283);
xor UO_1637 (O_1637,N_29046,N_29692);
and UO_1638 (O_1638,N_29173,N_29037);
nor UO_1639 (O_1639,N_29360,N_29459);
nand UO_1640 (O_1640,N_29052,N_29569);
nand UO_1641 (O_1641,N_29970,N_29500);
xnor UO_1642 (O_1642,N_29937,N_29668);
or UO_1643 (O_1643,N_29284,N_29127);
and UO_1644 (O_1644,N_29923,N_29318);
or UO_1645 (O_1645,N_29448,N_29145);
and UO_1646 (O_1646,N_29866,N_29065);
and UO_1647 (O_1647,N_29531,N_29885);
or UO_1648 (O_1648,N_29631,N_29944);
or UO_1649 (O_1649,N_29821,N_29997);
nor UO_1650 (O_1650,N_29676,N_29641);
nor UO_1651 (O_1651,N_29605,N_29033);
nand UO_1652 (O_1652,N_29419,N_29899);
or UO_1653 (O_1653,N_29308,N_29563);
and UO_1654 (O_1654,N_29078,N_29648);
or UO_1655 (O_1655,N_29545,N_29943);
nand UO_1656 (O_1656,N_29795,N_29109);
nand UO_1657 (O_1657,N_29245,N_29503);
xnor UO_1658 (O_1658,N_29748,N_29271);
nand UO_1659 (O_1659,N_29089,N_29168);
and UO_1660 (O_1660,N_29955,N_29374);
or UO_1661 (O_1661,N_29570,N_29946);
xor UO_1662 (O_1662,N_29659,N_29698);
nor UO_1663 (O_1663,N_29107,N_29223);
nor UO_1664 (O_1664,N_29469,N_29426);
xor UO_1665 (O_1665,N_29944,N_29418);
nor UO_1666 (O_1666,N_29133,N_29970);
and UO_1667 (O_1667,N_29397,N_29408);
nand UO_1668 (O_1668,N_29241,N_29318);
xor UO_1669 (O_1669,N_29818,N_29584);
nor UO_1670 (O_1670,N_29916,N_29153);
xor UO_1671 (O_1671,N_29410,N_29057);
or UO_1672 (O_1672,N_29510,N_29841);
or UO_1673 (O_1673,N_29265,N_29185);
nor UO_1674 (O_1674,N_29067,N_29279);
nand UO_1675 (O_1675,N_29576,N_29297);
and UO_1676 (O_1676,N_29410,N_29953);
or UO_1677 (O_1677,N_29948,N_29371);
xor UO_1678 (O_1678,N_29557,N_29523);
nand UO_1679 (O_1679,N_29544,N_29623);
nand UO_1680 (O_1680,N_29524,N_29891);
and UO_1681 (O_1681,N_29538,N_29499);
nand UO_1682 (O_1682,N_29038,N_29184);
xor UO_1683 (O_1683,N_29536,N_29001);
xor UO_1684 (O_1684,N_29127,N_29114);
nor UO_1685 (O_1685,N_29970,N_29969);
xor UO_1686 (O_1686,N_29832,N_29210);
xor UO_1687 (O_1687,N_29474,N_29235);
xnor UO_1688 (O_1688,N_29979,N_29366);
or UO_1689 (O_1689,N_29215,N_29922);
xor UO_1690 (O_1690,N_29390,N_29136);
xnor UO_1691 (O_1691,N_29893,N_29310);
and UO_1692 (O_1692,N_29490,N_29577);
or UO_1693 (O_1693,N_29643,N_29350);
or UO_1694 (O_1694,N_29475,N_29241);
xnor UO_1695 (O_1695,N_29378,N_29441);
xnor UO_1696 (O_1696,N_29227,N_29303);
nor UO_1697 (O_1697,N_29462,N_29615);
and UO_1698 (O_1698,N_29920,N_29796);
or UO_1699 (O_1699,N_29524,N_29072);
or UO_1700 (O_1700,N_29216,N_29867);
and UO_1701 (O_1701,N_29917,N_29334);
xnor UO_1702 (O_1702,N_29406,N_29117);
nor UO_1703 (O_1703,N_29081,N_29630);
xor UO_1704 (O_1704,N_29229,N_29637);
nor UO_1705 (O_1705,N_29609,N_29197);
or UO_1706 (O_1706,N_29226,N_29775);
and UO_1707 (O_1707,N_29570,N_29718);
xnor UO_1708 (O_1708,N_29526,N_29944);
xor UO_1709 (O_1709,N_29859,N_29088);
and UO_1710 (O_1710,N_29455,N_29284);
nand UO_1711 (O_1711,N_29234,N_29355);
nand UO_1712 (O_1712,N_29245,N_29108);
xnor UO_1713 (O_1713,N_29479,N_29455);
nand UO_1714 (O_1714,N_29164,N_29056);
or UO_1715 (O_1715,N_29368,N_29703);
nand UO_1716 (O_1716,N_29194,N_29349);
or UO_1717 (O_1717,N_29851,N_29435);
xor UO_1718 (O_1718,N_29009,N_29244);
nand UO_1719 (O_1719,N_29790,N_29505);
and UO_1720 (O_1720,N_29063,N_29604);
xor UO_1721 (O_1721,N_29508,N_29694);
nand UO_1722 (O_1722,N_29260,N_29469);
and UO_1723 (O_1723,N_29449,N_29476);
xnor UO_1724 (O_1724,N_29974,N_29578);
xor UO_1725 (O_1725,N_29081,N_29851);
nand UO_1726 (O_1726,N_29088,N_29821);
xnor UO_1727 (O_1727,N_29615,N_29237);
xor UO_1728 (O_1728,N_29585,N_29643);
nand UO_1729 (O_1729,N_29549,N_29607);
nand UO_1730 (O_1730,N_29203,N_29292);
and UO_1731 (O_1731,N_29382,N_29495);
nand UO_1732 (O_1732,N_29123,N_29862);
xnor UO_1733 (O_1733,N_29590,N_29820);
or UO_1734 (O_1734,N_29316,N_29477);
xnor UO_1735 (O_1735,N_29604,N_29171);
and UO_1736 (O_1736,N_29476,N_29810);
nor UO_1737 (O_1737,N_29529,N_29434);
nor UO_1738 (O_1738,N_29022,N_29905);
or UO_1739 (O_1739,N_29953,N_29087);
and UO_1740 (O_1740,N_29635,N_29456);
nand UO_1741 (O_1741,N_29039,N_29932);
and UO_1742 (O_1742,N_29073,N_29374);
xor UO_1743 (O_1743,N_29441,N_29613);
or UO_1744 (O_1744,N_29854,N_29084);
or UO_1745 (O_1745,N_29616,N_29407);
and UO_1746 (O_1746,N_29614,N_29523);
and UO_1747 (O_1747,N_29385,N_29648);
or UO_1748 (O_1748,N_29092,N_29941);
and UO_1749 (O_1749,N_29175,N_29181);
and UO_1750 (O_1750,N_29982,N_29575);
and UO_1751 (O_1751,N_29388,N_29459);
and UO_1752 (O_1752,N_29339,N_29753);
xnor UO_1753 (O_1753,N_29779,N_29712);
nor UO_1754 (O_1754,N_29694,N_29700);
nor UO_1755 (O_1755,N_29823,N_29582);
and UO_1756 (O_1756,N_29089,N_29348);
nor UO_1757 (O_1757,N_29895,N_29849);
xor UO_1758 (O_1758,N_29429,N_29947);
or UO_1759 (O_1759,N_29957,N_29347);
xnor UO_1760 (O_1760,N_29719,N_29677);
nor UO_1761 (O_1761,N_29429,N_29775);
nor UO_1762 (O_1762,N_29756,N_29206);
nand UO_1763 (O_1763,N_29126,N_29764);
nand UO_1764 (O_1764,N_29966,N_29624);
nand UO_1765 (O_1765,N_29045,N_29967);
or UO_1766 (O_1766,N_29433,N_29083);
nor UO_1767 (O_1767,N_29642,N_29981);
xor UO_1768 (O_1768,N_29455,N_29214);
or UO_1769 (O_1769,N_29046,N_29851);
xnor UO_1770 (O_1770,N_29762,N_29904);
nor UO_1771 (O_1771,N_29980,N_29847);
or UO_1772 (O_1772,N_29273,N_29927);
nor UO_1773 (O_1773,N_29164,N_29036);
nand UO_1774 (O_1774,N_29083,N_29516);
nand UO_1775 (O_1775,N_29177,N_29334);
nand UO_1776 (O_1776,N_29516,N_29212);
nand UO_1777 (O_1777,N_29113,N_29667);
or UO_1778 (O_1778,N_29501,N_29132);
xor UO_1779 (O_1779,N_29462,N_29665);
nor UO_1780 (O_1780,N_29317,N_29847);
nor UO_1781 (O_1781,N_29953,N_29801);
or UO_1782 (O_1782,N_29187,N_29916);
nand UO_1783 (O_1783,N_29754,N_29578);
nand UO_1784 (O_1784,N_29798,N_29179);
nand UO_1785 (O_1785,N_29188,N_29206);
nor UO_1786 (O_1786,N_29790,N_29202);
nor UO_1787 (O_1787,N_29091,N_29710);
nor UO_1788 (O_1788,N_29288,N_29212);
and UO_1789 (O_1789,N_29816,N_29180);
nand UO_1790 (O_1790,N_29050,N_29715);
xnor UO_1791 (O_1791,N_29230,N_29034);
nor UO_1792 (O_1792,N_29673,N_29733);
or UO_1793 (O_1793,N_29821,N_29949);
xnor UO_1794 (O_1794,N_29163,N_29168);
nor UO_1795 (O_1795,N_29174,N_29436);
or UO_1796 (O_1796,N_29942,N_29457);
or UO_1797 (O_1797,N_29420,N_29417);
nand UO_1798 (O_1798,N_29851,N_29840);
xnor UO_1799 (O_1799,N_29105,N_29419);
xnor UO_1800 (O_1800,N_29296,N_29401);
and UO_1801 (O_1801,N_29509,N_29932);
nand UO_1802 (O_1802,N_29325,N_29822);
or UO_1803 (O_1803,N_29831,N_29569);
xor UO_1804 (O_1804,N_29056,N_29727);
nand UO_1805 (O_1805,N_29673,N_29928);
and UO_1806 (O_1806,N_29170,N_29898);
nand UO_1807 (O_1807,N_29022,N_29991);
nand UO_1808 (O_1808,N_29345,N_29662);
or UO_1809 (O_1809,N_29321,N_29144);
nand UO_1810 (O_1810,N_29453,N_29948);
xnor UO_1811 (O_1811,N_29078,N_29500);
or UO_1812 (O_1812,N_29405,N_29915);
nand UO_1813 (O_1813,N_29741,N_29841);
nand UO_1814 (O_1814,N_29191,N_29940);
and UO_1815 (O_1815,N_29325,N_29222);
and UO_1816 (O_1816,N_29771,N_29109);
nor UO_1817 (O_1817,N_29702,N_29406);
and UO_1818 (O_1818,N_29075,N_29062);
and UO_1819 (O_1819,N_29270,N_29507);
xor UO_1820 (O_1820,N_29257,N_29871);
nand UO_1821 (O_1821,N_29871,N_29505);
or UO_1822 (O_1822,N_29125,N_29519);
or UO_1823 (O_1823,N_29552,N_29875);
nor UO_1824 (O_1824,N_29955,N_29186);
and UO_1825 (O_1825,N_29653,N_29130);
and UO_1826 (O_1826,N_29476,N_29311);
nor UO_1827 (O_1827,N_29177,N_29354);
nor UO_1828 (O_1828,N_29156,N_29052);
nand UO_1829 (O_1829,N_29371,N_29119);
or UO_1830 (O_1830,N_29273,N_29315);
nor UO_1831 (O_1831,N_29804,N_29002);
nor UO_1832 (O_1832,N_29254,N_29656);
and UO_1833 (O_1833,N_29946,N_29931);
or UO_1834 (O_1834,N_29985,N_29101);
nor UO_1835 (O_1835,N_29846,N_29903);
nor UO_1836 (O_1836,N_29063,N_29941);
nand UO_1837 (O_1837,N_29393,N_29717);
or UO_1838 (O_1838,N_29890,N_29703);
and UO_1839 (O_1839,N_29122,N_29472);
or UO_1840 (O_1840,N_29913,N_29051);
nand UO_1841 (O_1841,N_29199,N_29948);
and UO_1842 (O_1842,N_29359,N_29600);
nand UO_1843 (O_1843,N_29870,N_29426);
or UO_1844 (O_1844,N_29780,N_29298);
nand UO_1845 (O_1845,N_29461,N_29164);
or UO_1846 (O_1846,N_29734,N_29149);
and UO_1847 (O_1847,N_29116,N_29474);
nor UO_1848 (O_1848,N_29933,N_29047);
or UO_1849 (O_1849,N_29786,N_29759);
nor UO_1850 (O_1850,N_29255,N_29218);
xor UO_1851 (O_1851,N_29369,N_29024);
or UO_1852 (O_1852,N_29958,N_29052);
nor UO_1853 (O_1853,N_29503,N_29053);
nor UO_1854 (O_1854,N_29688,N_29415);
or UO_1855 (O_1855,N_29314,N_29450);
and UO_1856 (O_1856,N_29203,N_29856);
nand UO_1857 (O_1857,N_29274,N_29715);
or UO_1858 (O_1858,N_29904,N_29141);
nor UO_1859 (O_1859,N_29577,N_29328);
and UO_1860 (O_1860,N_29405,N_29889);
or UO_1861 (O_1861,N_29401,N_29953);
xor UO_1862 (O_1862,N_29457,N_29978);
or UO_1863 (O_1863,N_29084,N_29052);
or UO_1864 (O_1864,N_29876,N_29501);
nand UO_1865 (O_1865,N_29794,N_29153);
nor UO_1866 (O_1866,N_29352,N_29708);
nor UO_1867 (O_1867,N_29350,N_29613);
xnor UO_1868 (O_1868,N_29659,N_29000);
nor UO_1869 (O_1869,N_29211,N_29413);
or UO_1870 (O_1870,N_29965,N_29190);
and UO_1871 (O_1871,N_29269,N_29999);
or UO_1872 (O_1872,N_29430,N_29010);
xor UO_1873 (O_1873,N_29191,N_29406);
nor UO_1874 (O_1874,N_29435,N_29052);
xor UO_1875 (O_1875,N_29444,N_29157);
nand UO_1876 (O_1876,N_29017,N_29997);
nand UO_1877 (O_1877,N_29966,N_29625);
nand UO_1878 (O_1878,N_29730,N_29290);
nor UO_1879 (O_1879,N_29633,N_29559);
nand UO_1880 (O_1880,N_29555,N_29337);
nor UO_1881 (O_1881,N_29908,N_29095);
xor UO_1882 (O_1882,N_29688,N_29051);
or UO_1883 (O_1883,N_29719,N_29032);
or UO_1884 (O_1884,N_29937,N_29532);
and UO_1885 (O_1885,N_29927,N_29628);
and UO_1886 (O_1886,N_29197,N_29477);
nand UO_1887 (O_1887,N_29589,N_29147);
and UO_1888 (O_1888,N_29516,N_29747);
nor UO_1889 (O_1889,N_29917,N_29570);
xnor UO_1890 (O_1890,N_29974,N_29378);
nand UO_1891 (O_1891,N_29068,N_29413);
and UO_1892 (O_1892,N_29952,N_29934);
or UO_1893 (O_1893,N_29259,N_29122);
nor UO_1894 (O_1894,N_29151,N_29999);
nand UO_1895 (O_1895,N_29124,N_29895);
nand UO_1896 (O_1896,N_29801,N_29149);
and UO_1897 (O_1897,N_29379,N_29914);
xor UO_1898 (O_1898,N_29701,N_29918);
xnor UO_1899 (O_1899,N_29775,N_29074);
or UO_1900 (O_1900,N_29205,N_29769);
xnor UO_1901 (O_1901,N_29737,N_29706);
nor UO_1902 (O_1902,N_29908,N_29315);
or UO_1903 (O_1903,N_29225,N_29897);
or UO_1904 (O_1904,N_29046,N_29795);
nor UO_1905 (O_1905,N_29258,N_29644);
or UO_1906 (O_1906,N_29620,N_29228);
nor UO_1907 (O_1907,N_29228,N_29769);
xnor UO_1908 (O_1908,N_29831,N_29830);
xor UO_1909 (O_1909,N_29130,N_29078);
xor UO_1910 (O_1910,N_29317,N_29809);
or UO_1911 (O_1911,N_29258,N_29399);
nand UO_1912 (O_1912,N_29273,N_29346);
or UO_1913 (O_1913,N_29108,N_29748);
nand UO_1914 (O_1914,N_29400,N_29201);
nor UO_1915 (O_1915,N_29397,N_29388);
xnor UO_1916 (O_1916,N_29108,N_29887);
and UO_1917 (O_1917,N_29626,N_29209);
and UO_1918 (O_1918,N_29891,N_29070);
nor UO_1919 (O_1919,N_29932,N_29103);
nor UO_1920 (O_1920,N_29910,N_29264);
and UO_1921 (O_1921,N_29605,N_29706);
nor UO_1922 (O_1922,N_29505,N_29563);
or UO_1923 (O_1923,N_29608,N_29023);
and UO_1924 (O_1924,N_29313,N_29164);
nand UO_1925 (O_1925,N_29365,N_29280);
nor UO_1926 (O_1926,N_29349,N_29900);
nor UO_1927 (O_1927,N_29655,N_29281);
or UO_1928 (O_1928,N_29070,N_29686);
and UO_1929 (O_1929,N_29026,N_29825);
xor UO_1930 (O_1930,N_29841,N_29329);
or UO_1931 (O_1931,N_29922,N_29594);
xnor UO_1932 (O_1932,N_29562,N_29204);
nand UO_1933 (O_1933,N_29143,N_29079);
xnor UO_1934 (O_1934,N_29021,N_29437);
xor UO_1935 (O_1935,N_29128,N_29093);
or UO_1936 (O_1936,N_29914,N_29630);
nor UO_1937 (O_1937,N_29134,N_29140);
nor UO_1938 (O_1938,N_29594,N_29755);
and UO_1939 (O_1939,N_29216,N_29554);
and UO_1940 (O_1940,N_29552,N_29526);
nand UO_1941 (O_1941,N_29155,N_29196);
nand UO_1942 (O_1942,N_29636,N_29357);
or UO_1943 (O_1943,N_29366,N_29320);
xnor UO_1944 (O_1944,N_29964,N_29913);
and UO_1945 (O_1945,N_29692,N_29852);
xnor UO_1946 (O_1946,N_29824,N_29745);
nor UO_1947 (O_1947,N_29852,N_29593);
or UO_1948 (O_1948,N_29182,N_29580);
nand UO_1949 (O_1949,N_29898,N_29390);
nand UO_1950 (O_1950,N_29869,N_29079);
xor UO_1951 (O_1951,N_29745,N_29982);
xor UO_1952 (O_1952,N_29159,N_29107);
or UO_1953 (O_1953,N_29639,N_29255);
nor UO_1954 (O_1954,N_29764,N_29186);
nor UO_1955 (O_1955,N_29602,N_29453);
nor UO_1956 (O_1956,N_29073,N_29232);
or UO_1957 (O_1957,N_29269,N_29069);
xnor UO_1958 (O_1958,N_29913,N_29795);
nor UO_1959 (O_1959,N_29059,N_29512);
nor UO_1960 (O_1960,N_29356,N_29381);
xnor UO_1961 (O_1961,N_29355,N_29508);
nor UO_1962 (O_1962,N_29052,N_29619);
or UO_1963 (O_1963,N_29984,N_29908);
or UO_1964 (O_1964,N_29990,N_29712);
xnor UO_1965 (O_1965,N_29039,N_29212);
xor UO_1966 (O_1966,N_29869,N_29813);
xor UO_1967 (O_1967,N_29614,N_29464);
xor UO_1968 (O_1968,N_29724,N_29671);
nand UO_1969 (O_1969,N_29439,N_29009);
xor UO_1970 (O_1970,N_29300,N_29522);
or UO_1971 (O_1971,N_29277,N_29517);
nand UO_1972 (O_1972,N_29486,N_29525);
xnor UO_1973 (O_1973,N_29781,N_29055);
nor UO_1974 (O_1974,N_29484,N_29027);
nand UO_1975 (O_1975,N_29376,N_29334);
nand UO_1976 (O_1976,N_29299,N_29354);
xnor UO_1977 (O_1977,N_29986,N_29299);
xor UO_1978 (O_1978,N_29643,N_29480);
or UO_1979 (O_1979,N_29357,N_29451);
or UO_1980 (O_1980,N_29716,N_29844);
nor UO_1981 (O_1981,N_29847,N_29194);
and UO_1982 (O_1982,N_29288,N_29068);
or UO_1983 (O_1983,N_29136,N_29584);
xor UO_1984 (O_1984,N_29256,N_29944);
or UO_1985 (O_1985,N_29610,N_29232);
and UO_1986 (O_1986,N_29606,N_29022);
and UO_1987 (O_1987,N_29287,N_29044);
xor UO_1988 (O_1988,N_29218,N_29381);
xor UO_1989 (O_1989,N_29191,N_29730);
or UO_1990 (O_1990,N_29544,N_29342);
xor UO_1991 (O_1991,N_29057,N_29061);
and UO_1992 (O_1992,N_29027,N_29946);
or UO_1993 (O_1993,N_29364,N_29704);
nor UO_1994 (O_1994,N_29068,N_29074);
xor UO_1995 (O_1995,N_29725,N_29962);
and UO_1996 (O_1996,N_29783,N_29288);
xnor UO_1997 (O_1997,N_29331,N_29891);
nor UO_1998 (O_1998,N_29324,N_29701);
and UO_1999 (O_1999,N_29234,N_29491);
nand UO_2000 (O_2000,N_29755,N_29530);
or UO_2001 (O_2001,N_29849,N_29792);
and UO_2002 (O_2002,N_29199,N_29252);
nand UO_2003 (O_2003,N_29518,N_29656);
nor UO_2004 (O_2004,N_29221,N_29681);
nand UO_2005 (O_2005,N_29402,N_29765);
and UO_2006 (O_2006,N_29316,N_29790);
and UO_2007 (O_2007,N_29325,N_29583);
and UO_2008 (O_2008,N_29462,N_29494);
xnor UO_2009 (O_2009,N_29338,N_29299);
nand UO_2010 (O_2010,N_29395,N_29618);
and UO_2011 (O_2011,N_29044,N_29800);
or UO_2012 (O_2012,N_29753,N_29055);
xor UO_2013 (O_2013,N_29277,N_29186);
nand UO_2014 (O_2014,N_29605,N_29919);
and UO_2015 (O_2015,N_29682,N_29872);
xor UO_2016 (O_2016,N_29682,N_29359);
or UO_2017 (O_2017,N_29581,N_29738);
xor UO_2018 (O_2018,N_29681,N_29202);
or UO_2019 (O_2019,N_29160,N_29830);
xnor UO_2020 (O_2020,N_29512,N_29126);
xor UO_2021 (O_2021,N_29352,N_29674);
nor UO_2022 (O_2022,N_29386,N_29461);
nand UO_2023 (O_2023,N_29453,N_29073);
xnor UO_2024 (O_2024,N_29236,N_29147);
or UO_2025 (O_2025,N_29645,N_29027);
nor UO_2026 (O_2026,N_29973,N_29141);
nand UO_2027 (O_2027,N_29474,N_29534);
nand UO_2028 (O_2028,N_29182,N_29914);
nand UO_2029 (O_2029,N_29295,N_29365);
and UO_2030 (O_2030,N_29757,N_29598);
nor UO_2031 (O_2031,N_29068,N_29437);
or UO_2032 (O_2032,N_29227,N_29300);
or UO_2033 (O_2033,N_29327,N_29580);
nor UO_2034 (O_2034,N_29720,N_29674);
nor UO_2035 (O_2035,N_29192,N_29991);
xnor UO_2036 (O_2036,N_29687,N_29727);
and UO_2037 (O_2037,N_29748,N_29281);
xnor UO_2038 (O_2038,N_29679,N_29889);
nor UO_2039 (O_2039,N_29102,N_29479);
xnor UO_2040 (O_2040,N_29434,N_29428);
nor UO_2041 (O_2041,N_29997,N_29924);
xnor UO_2042 (O_2042,N_29938,N_29252);
xor UO_2043 (O_2043,N_29154,N_29195);
and UO_2044 (O_2044,N_29710,N_29026);
and UO_2045 (O_2045,N_29349,N_29937);
and UO_2046 (O_2046,N_29573,N_29586);
and UO_2047 (O_2047,N_29776,N_29438);
and UO_2048 (O_2048,N_29851,N_29192);
xor UO_2049 (O_2049,N_29162,N_29066);
xnor UO_2050 (O_2050,N_29260,N_29826);
nor UO_2051 (O_2051,N_29251,N_29315);
xnor UO_2052 (O_2052,N_29360,N_29045);
xnor UO_2053 (O_2053,N_29957,N_29190);
xnor UO_2054 (O_2054,N_29262,N_29463);
or UO_2055 (O_2055,N_29933,N_29156);
nor UO_2056 (O_2056,N_29296,N_29414);
nor UO_2057 (O_2057,N_29960,N_29873);
or UO_2058 (O_2058,N_29223,N_29568);
nor UO_2059 (O_2059,N_29493,N_29604);
or UO_2060 (O_2060,N_29087,N_29003);
or UO_2061 (O_2061,N_29142,N_29109);
and UO_2062 (O_2062,N_29381,N_29192);
xnor UO_2063 (O_2063,N_29162,N_29087);
xnor UO_2064 (O_2064,N_29061,N_29403);
nand UO_2065 (O_2065,N_29377,N_29680);
and UO_2066 (O_2066,N_29312,N_29110);
and UO_2067 (O_2067,N_29111,N_29355);
nor UO_2068 (O_2068,N_29204,N_29298);
xor UO_2069 (O_2069,N_29172,N_29634);
nand UO_2070 (O_2070,N_29062,N_29243);
and UO_2071 (O_2071,N_29080,N_29755);
or UO_2072 (O_2072,N_29879,N_29931);
nor UO_2073 (O_2073,N_29040,N_29177);
nand UO_2074 (O_2074,N_29657,N_29583);
or UO_2075 (O_2075,N_29605,N_29381);
nand UO_2076 (O_2076,N_29519,N_29196);
and UO_2077 (O_2077,N_29470,N_29332);
xnor UO_2078 (O_2078,N_29197,N_29864);
or UO_2079 (O_2079,N_29098,N_29123);
and UO_2080 (O_2080,N_29532,N_29807);
or UO_2081 (O_2081,N_29177,N_29906);
nor UO_2082 (O_2082,N_29939,N_29136);
nor UO_2083 (O_2083,N_29545,N_29989);
or UO_2084 (O_2084,N_29800,N_29731);
or UO_2085 (O_2085,N_29506,N_29143);
and UO_2086 (O_2086,N_29189,N_29419);
and UO_2087 (O_2087,N_29014,N_29568);
and UO_2088 (O_2088,N_29875,N_29585);
nor UO_2089 (O_2089,N_29196,N_29048);
nand UO_2090 (O_2090,N_29987,N_29483);
nand UO_2091 (O_2091,N_29694,N_29199);
and UO_2092 (O_2092,N_29587,N_29718);
or UO_2093 (O_2093,N_29753,N_29655);
nor UO_2094 (O_2094,N_29132,N_29339);
xor UO_2095 (O_2095,N_29877,N_29928);
or UO_2096 (O_2096,N_29312,N_29391);
xor UO_2097 (O_2097,N_29954,N_29391);
xnor UO_2098 (O_2098,N_29542,N_29749);
nand UO_2099 (O_2099,N_29988,N_29484);
or UO_2100 (O_2100,N_29994,N_29178);
nand UO_2101 (O_2101,N_29353,N_29026);
xnor UO_2102 (O_2102,N_29265,N_29977);
nand UO_2103 (O_2103,N_29713,N_29859);
or UO_2104 (O_2104,N_29779,N_29794);
nor UO_2105 (O_2105,N_29481,N_29202);
and UO_2106 (O_2106,N_29613,N_29273);
xnor UO_2107 (O_2107,N_29613,N_29237);
nand UO_2108 (O_2108,N_29645,N_29183);
nor UO_2109 (O_2109,N_29039,N_29692);
xnor UO_2110 (O_2110,N_29628,N_29780);
and UO_2111 (O_2111,N_29811,N_29909);
nand UO_2112 (O_2112,N_29499,N_29429);
nand UO_2113 (O_2113,N_29380,N_29976);
and UO_2114 (O_2114,N_29963,N_29979);
nor UO_2115 (O_2115,N_29357,N_29135);
and UO_2116 (O_2116,N_29207,N_29784);
and UO_2117 (O_2117,N_29569,N_29092);
xor UO_2118 (O_2118,N_29914,N_29426);
or UO_2119 (O_2119,N_29215,N_29932);
nor UO_2120 (O_2120,N_29285,N_29610);
or UO_2121 (O_2121,N_29416,N_29415);
xnor UO_2122 (O_2122,N_29402,N_29751);
and UO_2123 (O_2123,N_29545,N_29844);
or UO_2124 (O_2124,N_29676,N_29028);
or UO_2125 (O_2125,N_29384,N_29189);
nor UO_2126 (O_2126,N_29346,N_29480);
nand UO_2127 (O_2127,N_29000,N_29328);
xor UO_2128 (O_2128,N_29328,N_29858);
nand UO_2129 (O_2129,N_29743,N_29051);
xnor UO_2130 (O_2130,N_29385,N_29366);
xor UO_2131 (O_2131,N_29285,N_29280);
and UO_2132 (O_2132,N_29951,N_29976);
nor UO_2133 (O_2133,N_29964,N_29726);
and UO_2134 (O_2134,N_29467,N_29409);
and UO_2135 (O_2135,N_29864,N_29439);
or UO_2136 (O_2136,N_29860,N_29964);
xnor UO_2137 (O_2137,N_29705,N_29034);
or UO_2138 (O_2138,N_29480,N_29299);
and UO_2139 (O_2139,N_29162,N_29539);
nor UO_2140 (O_2140,N_29864,N_29775);
xor UO_2141 (O_2141,N_29034,N_29318);
or UO_2142 (O_2142,N_29340,N_29091);
and UO_2143 (O_2143,N_29336,N_29878);
nand UO_2144 (O_2144,N_29084,N_29220);
and UO_2145 (O_2145,N_29300,N_29697);
nand UO_2146 (O_2146,N_29506,N_29720);
nor UO_2147 (O_2147,N_29552,N_29495);
xnor UO_2148 (O_2148,N_29994,N_29691);
and UO_2149 (O_2149,N_29468,N_29214);
xor UO_2150 (O_2150,N_29943,N_29313);
nor UO_2151 (O_2151,N_29101,N_29571);
or UO_2152 (O_2152,N_29511,N_29591);
nor UO_2153 (O_2153,N_29939,N_29378);
nand UO_2154 (O_2154,N_29048,N_29951);
and UO_2155 (O_2155,N_29589,N_29884);
nand UO_2156 (O_2156,N_29331,N_29791);
or UO_2157 (O_2157,N_29962,N_29633);
xor UO_2158 (O_2158,N_29421,N_29307);
nor UO_2159 (O_2159,N_29899,N_29103);
or UO_2160 (O_2160,N_29149,N_29684);
and UO_2161 (O_2161,N_29879,N_29280);
or UO_2162 (O_2162,N_29464,N_29656);
and UO_2163 (O_2163,N_29210,N_29995);
nand UO_2164 (O_2164,N_29804,N_29485);
or UO_2165 (O_2165,N_29938,N_29411);
or UO_2166 (O_2166,N_29981,N_29507);
and UO_2167 (O_2167,N_29030,N_29701);
nor UO_2168 (O_2168,N_29975,N_29224);
nand UO_2169 (O_2169,N_29893,N_29448);
and UO_2170 (O_2170,N_29936,N_29990);
or UO_2171 (O_2171,N_29432,N_29373);
nand UO_2172 (O_2172,N_29676,N_29968);
and UO_2173 (O_2173,N_29578,N_29941);
nand UO_2174 (O_2174,N_29175,N_29685);
and UO_2175 (O_2175,N_29562,N_29890);
or UO_2176 (O_2176,N_29768,N_29790);
and UO_2177 (O_2177,N_29318,N_29176);
xnor UO_2178 (O_2178,N_29159,N_29576);
xnor UO_2179 (O_2179,N_29967,N_29581);
xnor UO_2180 (O_2180,N_29151,N_29186);
nor UO_2181 (O_2181,N_29541,N_29308);
xor UO_2182 (O_2182,N_29134,N_29747);
nand UO_2183 (O_2183,N_29637,N_29600);
and UO_2184 (O_2184,N_29416,N_29466);
or UO_2185 (O_2185,N_29994,N_29506);
nor UO_2186 (O_2186,N_29585,N_29974);
or UO_2187 (O_2187,N_29908,N_29107);
nor UO_2188 (O_2188,N_29110,N_29239);
xor UO_2189 (O_2189,N_29421,N_29398);
or UO_2190 (O_2190,N_29100,N_29930);
and UO_2191 (O_2191,N_29611,N_29939);
or UO_2192 (O_2192,N_29488,N_29535);
nand UO_2193 (O_2193,N_29532,N_29901);
nand UO_2194 (O_2194,N_29238,N_29266);
and UO_2195 (O_2195,N_29766,N_29134);
or UO_2196 (O_2196,N_29284,N_29567);
and UO_2197 (O_2197,N_29906,N_29675);
nand UO_2198 (O_2198,N_29939,N_29639);
nor UO_2199 (O_2199,N_29513,N_29118);
nand UO_2200 (O_2200,N_29471,N_29403);
or UO_2201 (O_2201,N_29066,N_29799);
nor UO_2202 (O_2202,N_29299,N_29035);
nand UO_2203 (O_2203,N_29388,N_29957);
nand UO_2204 (O_2204,N_29901,N_29862);
xnor UO_2205 (O_2205,N_29660,N_29135);
nand UO_2206 (O_2206,N_29581,N_29509);
nor UO_2207 (O_2207,N_29966,N_29836);
or UO_2208 (O_2208,N_29166,N_29064);
nor UO_2209 (O_2209,N_29374,N_29632);
or UO_2210 (O_2210,N_29422,N_29680);
or UO_2211 (O_2211,N_29634,N_29282);
or UO_2212 (O_2212,N_29914,N_29804);
nand UO_2213 (O_2213,N_29057,N_29029);
nand UO_2214 (O_2214,N_29949,N_29680);
xor UO_2215 (O_2215,N_29107,N_29743);
and UO_2216 (O_2216,N_29159,N_29422);
nor UO_2217 (O_2217,N_29993,N_29864);
and UO_2218 (O_2218,N_29422,N_29834);
or UO_2219 (O_2219,N_29815,N_29807);
xor UO_2220 (O_2220,N_29356,N_29593);
nand UO_2221 (O_2221,N_29244,N_29105);
nor UO_2222 (O_2222,N_29946,N_29949);
or UO_2223 (O_2223,N_29918,N_29482);
xnor UO_2224 (O_2224,N_29871,N_29048);
xor UO_2225 (O_2225,N_29518,N_29870);
nand UO_2226 (O_2226,N_29106,N_29483);
xnor UO_2227 (O_2227,N_29748,N_29058);
and UO_2228 (O_2228,N_29027,N_29452);
xor UO_2229 (O_2229,N_29335,N_29697);
nand UO_2230 (O_2230,N_29910,N_29510);
xnor UO_2231 (O_2231,N_29284,N_29015);
xor UO_2232 (O_2232,N_29538,N_29721);
nand UO_2233 (O_2233,N_29787,N_29377);
nor UO_2234 (O_2234,N_29751,N_29765);
nand UO_2235 (O_2235,N_29154,N_29532);
nand UO_2236 (O_2236,N_29258,N_29946);
and UO_2237 (O_2237,N_29483,N_29477);
or UO_2238 (O_2238,N_29175,N_29515);
or UO_2239 (O_2239,N_29683,N_29494);
xor UO_2240 (O_2240,N_29719,N_29017);
or UO_2241 (O_2241,N_29112,N_29691);
nor UO_2242 (O_2242,N_29217,N_29110);
or UO_2243 (O_2243,N_29240,N_29579);
and UO_2244 (O_2244,N_29824,N_29258);
or UO_2245 (O_2245,N_29457,N_29867);
or UO_2246 (O_2246,N_29406,N_29441);
nand UO_2247 (O_2247,N_29734,N_29687);
nand UO_2248 (O_2248,N_29205,N_29617);
nand UO_2249 (O_2249,N_29794,N_29240);
nor UO_2250 (O_2250,N_29953,N_29898);
or UO_2251 (O_2251,N_29556,N_29952);
and UO_2252 (O_2252,N_29743,N_29605);
nand UO_2253 (O_2253,N_29641,N_29599);
nand UO_2254 (O_2254,N_29909,N_29403);
and UO_2255 (O_2255,N_29646,N_29126);
or UO_2256 (O_2256,N_29502,N_29193);
and UO_2257 (O_2257,N_29285,N_29602);
nand UO_2258 (O_2258,N_29547,N_29822);
or UO_2259 (O_2259,N_29838,N_29826);
xnor UO_2260 (O_2260,N_29449,N_29543);
xnor UO_2261 (O_2261,N_29913,N_29452);
and UO_2262 (O_2262,N_29764,N_29069);
or UO_2263 (O_2263,N_29449,N_29362);
xor UO_2264 (O_2264,N_29532,N_29782);
xnor UO_2265 (O_2265,N_29252,N_29928);
and UO_2266 (O_2266,N_29066,N_29051);
xor UO_2267 (O_2267,N_29362,N_29091);
nand UO_2268 (O_2268,N_29165,N_29054);
or UO_2269 (O_2269,N_29401,N_29785);
and UO_2270 (O_2270,N_29002,N_29379);
and UO_2271 (O_2271,N_29973,N_29767);
nor UO_2272 (O_2272,N_29850,N_29777);
or UO_2273 (O_2273,N_29039,N_29733);
and UO_2274 (O_2274,N_29350,N_29862);
or UO_2275 (O_2275,N_29182,N_29179);
or UO_2276 (O_2276,N_29182,N_29002);
nand UO_2277 (O_2277,N_29424,N_29732);
xor UO_2278 (O_2278,N_29331,N_29517);
or UO_2279 (O_2279,N_29385,N_29941);
xnor UO_2280 (O_2280,N_29970,N_29092);
xor UO_2281 (O_2281,N_29416,N_29359);
nor UO_2282 (O_2282,N_29702,N_29812);
and UO_2283 (O_2283,N_29305,N_29139);
nand UO_2284 (O_2284,N_29999,N_29466);
and UO_2285 (O_2285,N_29053,N_29273);
nor UO_2286 (O_2286,N_29740,N_29488);
or UO_2287 (O_2287,N_29554,N_29627);
or UO_2288 (O_2288,N_29836,N_29690);
or UO_2289 (O_2289,N_29047,N_29438);
nor UO_2290 (O_2290,N_29975,N_29063);
nor UO_2291 (O_2291,N_29257,N_29612);
nand UO_2292 (O_2292,N_29499,N_29279);
nand UO_2293 (O_2293,N_29668,N_29923);
xnor UO_2294 (O_2294,N_29876,N_29763);
or UO_2295 (O_2295,N_29025,N_29189);
and UO_2296 (O_2296,N_29164,N_29858);
nor UO_2297 (O_2297,N_29906,N_29877);
or UO_2298 (O_2298,N_29040,N_29527);
or UO_2299 (O_2299,N_29430,N_29592);
or UO_2300 (O_2300,N_29049,N_29573);
nand UO_2301 (O_2301,N_29162,N_29023);
nand UO_2302 (O_2302,N_29353,N_29598);
and UO_2303 (O_2303,N_29756,N_29702);
xnor UO_2304 (O_2304,N_29251,N_29689);
xnor UO_2305 (O_2305,N_29165,N_29435);
xor UO_2306 (O_2306,N_29768,N_29919);
xnor UO_2307 (O_2307,N_29084,N_29544);
nand UO_2308 (O_2308,N_29074,N_29647);
or UO_2309 (O_2309,N_29947,N_29989);
xnor UO_2310 (O_2310,N_29782,N_29775);
xnor UO_2311 (O_2311,N_29424,N_29697);
and UO_2312 (O_2312,N_29736,N_29291);
xnor UO_2313 (O_2313,N_29871,N_29636);
nor UO_2314 (O_2314,N_29781,N_29692);
and UO_2315 (O_2315,N_29908,N_29868);
xnor UO_2316 (O_2316,N_29837,N_29523);
and UO_2317 (O_2317,N_29942,N_29730);
xnor UO_2318 (O_2318,N_29082,N_29342);
or UO_2319 (O_2319,N_29951,N_29561);
nand UO_2320 (O_2320,N_29694,N_29749);
and UO_2321 (O_2321,N_29193,N_29827);
nor UO_2322 (O_2322,N_29763,N_29573);
or UO_2323 (O_2323,N_29682,N_29317);
xnor UO_2324 (O_2324,N_29321,N_29980);
and UO_2325 (O_2325,N_29910,N_29100);
nor UO_2326 (O_2326,N_29183,N_29858);
and UO_2327 (O_2327,N_29760,N_29081);
or UO_2328 (O_2328,N_29504,N_29640);
and UO_2329 (O_2329,N_29688,N_29969);
and UO_2330 (O_2330,N_29767,N_29289);
nor UO_2331 (O_2331,N_29121,N_29324);
nand UO_2332 (O_2332,N_29765,N_29636);
nor UO_2333 (O_2333,N_29771,N_29806);
and UO_2334 (O_2334,N_29602,N_29629);
nor UO_2335 (O_2335,N_29488,N_29275);
or UO_2336 (O_2336,N_29707,N_29616);
or UO_2337 (O_2337,N_29679,N_29691);
and UO_2338 (O_2338,N_29742,N_29866);
nor UO_2339 (O_2339,N_29501,N_29881);
xor UO_2340 (O_2340,N_29555,N_29357);
and UO_2341 (O_2341,N_29324,N_29412);
xor UO_2342 (O_2342,N_29882,N_29801);
xnor UO_2343 (O_2343,N_29005,N_29173);
xor UO_2344 (O_2344,N_29908,N_29753);
nand UO_2345 (O_2345,N_29615,N_29173);
xnor UO_2346 (O_2346,N_29216,N_29486);
nor UO_2347 (O_2347,N_29817,N_29657);
or UO_2348 (O_2348,N_29450,N_29449);
nor UO_2349 (O_2349,N_29624,N_29679);
or UO_2350 (O_2350,N_29858,N_29576);
nor UO_2351 (O_2351,N_29455,N_29069);
nor UO_2352 (O_2352,N_29243,N_29344);
and UO_2353 (O_2353,N_29935,N_29187);
or UO_2354 (O_2354,N_29556,N_29186);
and UO_2355 (O_2355,N_29630,N_29194);
xnor UO_2356 (O_2356,N_29606,N_29402);
nor UO_2357 (O_2357,N_29844,N_29816);
nor UO_2358 (O_2358,N_29552,N_29137);
or UO_2359 (O_2359,N_29942,N_29072);
or UO_2360 (O_2360,N_29704,N_29327);
and UO_2361 (O_2361,N_29587,N_29068);
nand UO_2362 (O_2362,N_29259,N_29204);
nand UO_2363 (O_2363,N_29162,N_29006);
and UO_2364 (O_2364,N_29663,N_29233);
nor UO_2365 (O_2365,N_29961,N_29167);
and UO_2366 (O_2366,N_29154,N_29394);
or UO_2367 (O_2367,N_29864,N_29634);
nand UO_2368 (O_2368,N_29899,N_29721);
nand UO_2369 (O_2369,N_29498,N_29222);
xnor UO_2370 (O_2370,N_29579,N_29785);
nor UO_2371 (O_2371,N_29729,N_29942);
xor UO_2372 (O_2372,N_29485,N_29494);
xnor UO_2373 (O_2373,N_29981,N_29600);
nor UO_2374 (O_2374,N_29718,N_29177);
nand UO_2375 (O_2375,N_29663,N_29208);
xor UO_2376 (O_2376,N_29483,N_29225);
nand UO_2377 (O_2377,N_29866,N_29240);
xor UO_2378 (O_2378,N_29551,N_29394);
and UO_2379 (O_2379,N_29657,N_29184);
or UO_2380 (O_2380,N_29158,N_29938);
and UO_2381 (O_2381,N_29427,N_29737);
or UO_2382 (O_2382,N_29278,N_29785);
nor UO_2383 (O_2383,N_29085,N_29105);
nand UO_2384 (O_2384,N_29125,N_29900);
and UO_2385 (O_2385,N_29919,N_29552);
nand UO_2386 (O_2386,N_29091,N_29178);
xnor UO_2387 (O_2387,N_29189,N_29182);
xor UO_2388 (O_2388,N_29174,N_29011);
nand UO_2389 (O_2389,N_29016,N_29460);
and UO_2390 (O_2390,N_29691,N_29594);
and UO_2391 (O_2391,N_29990,N_29191);
nor UO_2392 (O_2392,N_29897,N_29980);
xor UO_2393 (O_2393,N_29409,N_29259);
and UO_2394 (O_2394,N_29413,N_29872);
and UO_2395 (O_2395,N_29803,N_29396);
nor UO_2396 (O_2396,N_29134,N_29256);
nor UO_2397 (O_2397,N_29001,N_29061);
or UO_2398 (O_2398,N_29388,N_29758);
xnor UO_2399 (O_2399,N_29043,N_29506);
nor UO_2400 (O_2400,N_29367,N_29952);
nand UO_2401 (O_2401,N_29157,N_29194);
and UO_2402 (O_2402,N_29216,N_29368);
and UO_2403 (O_2403,N_29745,N_29156);
xor UO_2404 (O_2404,N_29193,N_29643);
or UO_2405 (O_2405,N_29656,N_29945);
and UO_2406 (O_2406,N_29412,N_29082);
xor UO_2407 (O_2407,N_29573,N_29823);
nor UO_2408 (O_2408,N_29570,N_29520);
or UO_2409 (O_2409,N_29732,N_29011);
nor UO_2410 (O_2410,N_29823,N_29463);
nor UO_2411 (O_2411,N_29839,N_29579);
and UO_2412 (O_2412,N_29887,N_29267);
or UO_2413 (O_2413,N_29918,N_29420);
or UO_2414 (O_2414,N_29297,N_29738);
xnor UO_2415 (O_2415,N_29104,N_29549);
nor UO_2416 (O_2416,N_29680,N_29854);
xor UO_2417 (O_2417,N_29476,N_29126);
nand UO_2418 (O_2418,N_29990,N_29567);
nor UO_2419 (O_2419,N_29198,N_29895);
or UO_2420 (O_2420,N_29951,N_29851);
xnor UO_2421 (O_2421,N_29618,N_29961);
nor UO_2422 (O_2422,N_29828,N_29087);
nand UO_2423 (O_2423,N_29302,N_29050);
xnor UO_2424 (O_2424,N_29817,N_29406);
nor UO_2425 (O_2425,N_29125,N_29299);
or UO_2426 (O_2426,N_29110,N_29067);
nand UO_2427 (O_2427,N_29477,N_29789);
xor UO_2428 (O_2428,N_29529,N_29335);
nand UO_2429 (O_2429,N_29980,N_29948);
nor UO_2430 (O_2430,N_29646,N_29743);
and UO_2431 (O_2431,N_29897,N_29948);
or UO_2432 (O_2432,N_29177,N_29321);
nand UO_2433 (O_2433,N_29409,N_29630);
nand UO_2434 (O_2434,N_29294,N_29027);
xnor UO_2435 (O_2435,N_29638,N_29234);
nor UO_2436 (O_2436,N_29700,N_29498);
nor UO_2437 (O_2437,N_29710,N_29553);
nor UO_2438 (O_2438,N_29382,N_29856);
and UO_2439 (O_2439,N_29724,N_29382);
or UO_2440 (O_2440,N_29016,N_29272);
nand UO_2441 (O_2441,N_29926,N_29465);
or UO_2442 (O_2442,N_29562,N_29250);
xor UO_2443 (O_2443,N_29323,N_29770);
xnor UO_2444 (O_2444,N_29734,N_29859);
nor UO_2445 (O_2445,N_29086,N_29278);
or UO_2446 (O_2446,N_29495,N_29412);
xnor UO_2447 (O_2447,N_29635,N_29889);
and UO_2448 (O_2448,N_29508,N_29640);
or UO_2449 (O_2449,N_29683,N_29643);
nand UO_2450 (O_2450,N_29276,N_29803);
or UO_2451 (O_2451,N_29798,N_29950);
xor UO_2452 (O_2452,N_29907,N_29883);
xnor UO_2453 (O_2453,N_29620,N_29432);
xor UO_2454 (O_2454,N_29327,N_29681);
nor UO_2455 (O_2455,N_29869,N_29416);
nor UO_2456 (O_2456,N_29216,N_29384);
or UO_2457 (O_2457,N_29687,N_29940);
xor UO_2458 (O_2458,N_29335,N_29615);
or UO_2459 (O_2459,N_29554,N_29103);
and UO_2460 (O_2460,N_29374,N_29987);
and UO_2461 (O_2461,N_29533,N_29767);
and UO_2462 (O_2462,N_29733,N_29792);
nand UO_2463 (O_2463,N_29533,N_29106);
or UO_2464 (O_2464,N_29589,N_29042);
xnor UO_2465 (O_2465,N_29551,N_29759);
and UO_2466 (O_2466,N_29547,N_29186);
or UO_2467 (O_2467,N_29474,N_29149);
xnor UO_2468 (O_2468,N_29839,N_29909);
nand UO_2469 (O_2469,N_29527,N_29274);
nand UO_2470 (O_2470,N_29604,N_29364);
nand UO_2471 (O_2471,N_29525,N_29650);
nor UO_2472 (O_2472,N_29623,N_29604);
nand UO_2473 (O_2473,N_29597,N_29826);
and UO_2474 (O_2474,N_29967,N_29897);
nor UO_2475 (O_2475,N_29601,N_29411);
and UO_2476 (O_2476,N_29597,N_29383);
nand UO_2477 (O_2477,N_29950,N_29373);
xor UO_2478 (O_2478,N_29138,N_29765);
nor UO_2479 (O_2479,N_29535,N_29177);
xor UO_2480 (O_2480,N_29324,N_29925);
or UO_2481 (O_2481,N_29822,N_29541);
and UO_2482 (O_2482,N_29253,N_29489);
nor UO_2483 (O_2483,N_29126,N_29441);
and UO_2484 (O_2484,N_29953,N_29840);
nor UO_2485 (O_2485,N_29321,N_29948);
and UO_2486 (O_2486,N_29578,N_29229);
and UO_2487 (O_2487,N_29612,N_29323);
or UO_2488 (O_2488,N_29973,N_29282);
nor UO_2489 (O_2489,N_29602,N_29576);
nand UO_2490 (O_2490,N_29996,N_29962);
or UO_2491 (O_2491,N_29023,N_29239);
xnor UO_2492 (O_2492,N_29588,N_29359);
nand UO_2493 (O_2493,N_29972,N_29942);
and UO_2494 (O_2494,N_29729,N_29768);
or UO_2495 (O_2495,N_29088,N_29284);
nand UO_2496 (O_2496,N_29940,N_29753);
xnor UO_2497 (O_2497,N_29530,N_29179);
or UO_2498 (O_2498,N_29938,N_29792);
nand UO_2499 (O_2499,N_29853,N_29354);
and UO_2500 (O_2500,N_29478,N_29761);
and UO_2501 (O_2501,N_29558,N_29613);
xnor UO_2502 (O_2502,N_29593,N_29974);
or UO_2503 (O_2503,N_29158,N_29799);
nor UO_2504 (O_2504,N_29684,N_29217);
or UO_2505 (O_2505,N_29229,N_29844);
or UO_2506 (O_2506,N_29511,N_29810);
nor UO_2507 (O_2507,N_29332,N_29699);
nand UO_2508 (O_2508,N_29010,N_29452);
xnor UO_2509 (O_2509,N_29904,N_29328);
or UO_2510 (O_2510,N_29242,N_29571);
or UO_2511 (O_2511,N_29349,N_29298);
or UO_2512 (O_2512,N_29415,N_29466);
nand UO_2513 (O_2513,N_29296,N_29363);
or UO_2514 (O_2514,N_29662,N_29321);
nor UO_2515 (O_2515,N_29310,N_29070);
nand UO_2516 (O_2516,N_29594,N_29018);
and UO_2517 (O_2517,N_29980,N_29540);
nand UO_2518 (O_2518,N_29000,N_29297);
nand UO_2519 (O_2519,N_29207,N_29197);
xnor UO_2520 (O_2520,N_29827,N_29249);
and UO_2521 (O_2521,N_29122,N_29059);
xnor UO_2522 (O_2522,N_29523,N_29550);
or UO_2523 (O_2523,N_29106,N_29846);
xnor UO_2524 (O_2524,N_29608,N_29274);
and UO_2525 (O_2525,N_29943,N_29431);
nand UO_2526 (O_2526,N_29747,N_29147);
nor UO_2527 (O_2527,N_29509,N_29927);
xor UO_2528 (O_2528,N_29529,N_29242);
xor UO_2529 (O_2529,N_29023,N_29025);
nand UO_2530 (O_2530,N_29017,N_29545);
nand UO_2531 (O_2531,N_29541,N_29756);
xnor UO_2532 (O_2532,N_29036,N_29343);
xor UO_2533 (O_2533,N_29526,N_29342);
and UO_2534 (O_2534,N_29444,N_29717);
xnor UO_2535 (O_2535,N_29115,N_29236);
xor UO_2536 (O_2536,N_29148,N_29404);
xnor UO_2537 (O_2537,N_29064,N_29164);
xnor UO_2538 (O_2538,N_29111,N_29569);
or UO_2539 (O_2539,N_29682,N_29290);
nor UO_2540 (O_2540,N_29170,N_29886);
nor UO_2541 (O_2541,N_29023,N_29233);
and UO_2542 (O_2542,N_29674,N_29764);
and UO_2543 (O_2543,N_29739,N_29760);
nor UO_2544 (O_2544,N_29224,N_29529);
xnor UO_2545 (O_2545,N_29866,N_29382);
nor UO_2546 (O_2546,N_29927,N_29351);
xnor UO_2547 (O_2547,N_29311,N_29559);
nor UO_2548 (O_2548,N_29986,N_29750);
or UO_2549 (O_2549,N_29995,N_29401);
or UO_2550 (O_2550,N_29767,N_29916);
and UO_2551 (O_2551,N_29174,N_29859);
or UO_2552 (O_2552,N_29998,N_29807);
nand UO_2553 (O_2553,N_29955,N_29978);
xor UO_2554 (O_2554,N_29571,N_29929);
or UO_2555 (O_2555,N_29208,N_29550);
nand UO_2556 (O_2556,N_29533,N_29372);
and UO_2557 (O_2557,N_29097,N_29396);
nand UO_2558 (O_2558,N_29882,N_29314);
or UO_2559 (O_2559,N_29325,N_29843);
nand UO_2560 (O_2560,N_29777,N_29693);
nand UO_2561 (O_2561,N_29280,N_29789);
or UO_2562 (O_2562,N_29060,N_29356);
nand UO_2563 (O_2563,N_29257,N_29750);
and UO_2564 (O_2564,N_29417,N_29481);
xnor UO_2565 (O_2565,N_29984,N_29622);
nor UO_2566 (O_2566,N_29943,N_29822);
nand UO_2567 (O_2567,N_29183,N_29990);
nor UO_2568 (O_2568,N_29515,N_29454);
or UO_2569 (O_2569,N_29711,N_29913);
nor UO_2570 (O_2570,N_29882,N_29107);
and UO_2571 (O_2571,N_29503,N_29815);
nand UO_2572 (O_2572,N_29284,N_29009);
xor UO_2573 (O_2573,N_29001,N_29400);
or UO_2574 (O_2574,N_29225,N_29912);
or UO_2575 (O_2575,N_29371,N_29905);
nor UO_2576 (O_2576,N_29739,N_29807);
and UO_2577 (O_2577,N_29784,N_29100);
and UO_2578 (O_2578,N_29977,N_29149);
nand UO_2579 (O_2579,N_29386,N_29127);
nor UO_2580 (O_2580,N_29258,N_29547);
or UO_2581 (O_2581,N_29684,N_29964);
or UO_2582 (O_2582,N_29885,N_29108);
nor UO_2583 (O_2583,N_29764,N_29292);
and UO_2584 (O_2584,N_29018,N_29392);
nand UO_2585 (O_2585,N_29121,N_29646);
nor UO_2586 (O_2586,N_29716,N_29029);
nand UO_2587 (O_2587,N_29200,N_29953);
or UO_2588 (O_2588,N_29660,N_29178);
and UO_2589 (O_2589,N_29907,N_29486);
xnor UO_2590 (O_2590,N_29174,N_29645);
or UO_2591 (O_2591,N_29393,N_29235);
nand UO_2592 (O_2592,N_29697,N_29196);
nor UO_2593 (O_2593,N_29245,N_29683);
xnor UO_2594 (O_2594,N_29416,N_29867);
or UO_2595 (O_2595,N_29170,N_29427);
nor UO_2596 (O_2596,N_29457,N_29817);
or UO_2597 (O_2597,N_29279,N_29409);
nor UO_2598 (O_2598,N_29671,N_29160);
and UO_2599 (O_2599,N_29731,N_29583);
nor UO_2600 (O_2600,N_29385,N_29712);
or UO_2601 (O_2601,N_29413,N_29870);
xnor UO_2602 (O_2602,N_29365,N_29225);
nand UO_2603 (O_2603,N_29154,N_29143);
and UO_2604 (O_2604,N_29900,N_29075);
xnor UO_2605 (O_2605,N_29789,N_29571);
xnor UO_2606 (O_2606,N_29811,N_29346);
or UO_2607 (O_2607,N_29328,N_29103);
nor UO_2608 (O_2608,N_29940,N_29870);
or UO_2609 (O_2609,N_29192,N_29157);
xor UO_2610 (O_2610,N_29113,N_29731);
and UO_2611 (O_2611,N_29788,N_29698);
and UO_2612 (O_2612,N_29713,N_29120);
nand UO_2613 (O_2613,N_29519,N_29947);
xnor UO_2614 (O_2614,N_29296,N_29634);
nor UO_2615 (O_2615,N_29977,N_29365);
or UO_2616 (O_2616,N_29669,N_29994);
or UO_2617 (O_2617,N_29993,N_29767);
nand UO_2618 (O_2618,N_29248,N_29971);
nand UO_2619 (O_2619,N_29242,N_29123);
xor UO_2620 (O_2620,N_29632,N_29878);
nand UO_2621 (O_2621,N_29596,N_29630);
nor UO_2622 (O_2622,N_29813,N_29659);
nand UO_2623 (O_2623,N_29723,N_29129);
nor UO_2624 (O_2624,N_29225,N_29812);
or UO_2625 (O_2625,N_29743,N_29364);
or UO_2626 (O_2626,N_29734,N_29235);
and UO_2627 (O_2627,N_29769,N_29361);
or UO_2628 (O_2628,N_29437,N_29134);
or UO_2629 (O_2629,N_29134,N_29402);
nand UO_2630 (O_2630,N_29728,N_29789);
or UO_2631 (O_2631,N_29454,N_29035);
and UO_2632 (O_2632,N_29858,N_29206);
nand UO_2633 (O_2633,N_29917,N_29709);
or UO_2634 (O_2634,N_29709,N_29984);
nand UO_2635 (O_2635,N_29252,N_29072);
or UO_2636 (O_2636,N_29745,N_29133);
and UO_2637 (O_2637,N_29850,N_29016);
nor UO_2638 (O_2638,N_29937,N_29766);
nand UO_2639 (O_2639,N_29082,N_29665);
nor UO_2640 (O_2640,N_29550,N_29128);
and UO_2641 (O_2641,N_29458,N_29834);
or UO_2642 (O_2642,N_29002,N_29447);
nor UO_2643 (O_2643,N_29614,N_29885);
xor UO_2644 (O_2644,N_29533,N_29360);
xnor UO_2645 (O_2645,N_29128,N_29098);
nand UO_2646 (O_2646,N_29436,N_29851);
nand UO_2647 (O_2647,N_29582,N_29895);
or UO_2648 (O_2648,N_29873,N_29344);
xor UO_2649 (O_2649,N_29408,N_29990);
or UO_2650 (O_2650,N_29411,N_29686);
nor UO_2651 (O_2651,N_29494,N_29841);
or UO_2652 (O_2652,N_29149,N_29838);
xor UO_2653 (O_2653,N_29555,N_29447);
and UO_2654 (O_2654,N_29909,N_29609);
nor UO_2655 (O_2655,N_29003,N_29708);
xnor UO_2656 (O_2656,N_29467,N_29717);
xor UO_2657 (O_2657,N_29227,N_29178);
nand UO_2658 (O_2658,N_29863,N_29934);
or UO_2659 (O_2659,N_29153,N_29903);
and UO_2660 (O_2660,N_29289,N_29862);
xnor UO_2661 (O_2661,N_29503,N_29336);
nor UO_2662 (O_2662,N_29688,N_29128);
nand UO_2663 (O_2663,N_29748,N_29077);
nor UO_2664 (O_2664,N_29294,N_29377);
and UO_2665 (O_2665,N_29515,N_29613);
nand UO_2666 (O_2666,N_29975,N_29938);
or UO_2667 (O_2667,N_29235,N_29019);
xor UO_2668 (O_2668,N_29659,N_29194);
nand UO_2669 (O_2669,N_29377,N_29238);
nor UO_2670 (O_2670,N_29703,N_29153);
xor UO_2671 (O_2671,N_29861,N_29707);
and UO_2672 (O_2672,N_29661,N_29400);
nor UO_2673 (O_2673,N_29042,N_29567);
and UO_2674 (O_2674,N_29790,N_29331);
or UO_2675 (O_2675,N_29278,N_29578);
nand UO_2676 (O_2676,N_29032,N_29704);
and UO_2677 (O_2677,N_29285,N_29752);
xnor UO_2678 (O_2678,N_29417,N_29283);
nor UO_2679 (O_2679,N_29453,N_29622);
or UO_2680 (O_2680,N_29511,N_29871);
nand UO_2681 (O_2681,N_29116,N_29141);
and UO_2682 (O_2682,N_29249,N_29977);
xnor UO_2683 (O_2683,N_29241,N_29471);
nand UO_2684 (O_2684,N_29425,N_29880);
nor UO_2685 (O_2685,N_29967,N_29369);
nor UO_2686 (O_2686,N_29837,N_29746);
or UO_2687 (O_2687,N_29139,N_29467);
or UO_2688 (O_2688,N_29096,N_29072);
nor UO_2689 (O_2689,N_29804,N_29960);
and UO_2690 (O_2690,N_29511,N_29610);
nand UO_2691 (O_2691,N_29456,N_29220);
nor UO_2692 (O_2692,N_29161,N_29999);
or UO_2693 (O_2693,N_29079,N_29460);
or UO_2694 (O_2694,N_29603,N_29810);
nor UO_2695 (O_2695,N_29880,N_29538);
and UO_2696 (O_2696,N_29097,N_29607);
or UO_2697 (O_2697,N_29092,N_29768);
and UO_2698 (O_2698,N_29239,N_29141);
or UO_2699 (O_2699,N_29156,N_29137);
nand UO_2700 (O_2700,N_29469,N_29461);
and UO_2701 (O_2701,N_29152,N_29441);
or UO_2702 (O_2702,N_29503,N_29893);
and UO_2703 (O_2703,N_29349,N_29328);
xnor UO_2704 (O_2704,N_29444,N_29121);
xor UO_2705 (O_2705,N_29144,N_29379);
nor UO_2706 (O_2706,N_29336,N_29234);
or UO_2707 (O_2707,N_29424,N_29870);
nor UO_2708 (O_2708,N_29595,N_29311);
nand UO_2709 (O_2709,N_29175,N_29876);
and UO_2710 (O_2710,N_29037,N_29534);
nand UO_2711 (O_2711,N_29322,N_29854);
or UO_2712 (O_2712,N_29828,N_29654);
nand UO_2713 (O_2713,N_29407,N_29204);
nand UO_2714 (O_2714,N_29061,N_29477);
and UO_2715 (O_2715,N_29974,N_29916);
and UO_2716 (O_2716,N_29748,N_29219);
and UO_2717 (O_2717,N_29182,N_29598);
nand UO_2718 (O_2718,N_29551,N_29077);
and UO_2719 (O_2719,N_29002,N_29113);
or UO_2720 (O_2720,N_29724,N_29777);
or UO_2721 (O_2721,N_29876,N_29960);
or UO_2722 (O_2722,N_29052,N_29533);
nor UO_2723 (O_2723,N_29310,N_29717);
and UO_2724 (O_2724,N_29380,N_29423);
nand UO_2725 (O_2725,N_29907,N_29650);
or UO_2726 (O_2726,N_29800,N_29201);
or UO_2727 (O_2727,N_29064,N_29001);
nand UO_2728 (O_2728,N_29824,N_29995);
nor UO_2729 (O_2729,N_29586,N_29420);
nand UO_2730 (O_2730,N_29501,N_29475);
and UO_2731 (O_2731,N_29780,N_29331);
or UO_2732 (O_2732,N_29121,N_29706);
xnor UO_2733 (O_2733,N_29494,N_29514);
nor UO_2734 (O_2734,N_29472,N_29474);
nor UO_2735 (O_2735,N_29018,N_29861);
nor UO_2736 (O_2736,N_29936,N_29218);
and UO_2737 (O_2737,N_29876,N_29332);
and UO_2738 (O_2738,N_29144,N_29544);
and UO_2739 (O_2739,N_29779,N_29064);
and UO_2740 (O_2740,N_29321,N_29514);
xnor UO_2741 (O_2741,N_29645,N_29433);
nor UO_2742 (O_2742,N_29144,N_29223);
nand UO_2743 (O_2743,N_29735,N_29211);
xor UO_2744 (O_2744,N_29704,N_29393);
and UO_2745 (O_2745,N_29642,N_29937);
xnor UO_2746 (O_2746,N_29435,N_29941);
nor UO_2747 (O_2747,N_29175,N_29153);
xor UO_2748 (O_2748,N_29304,N_29612);
nand UO_2749 (O_2749,N_29769,N_29974);
or UO_2750 (O_2750,N_29279,N_29459);
xor UO_2751 (O_2751,N_29915,N_29847);
or UO_2752 (O_2752,N_29400,N_29867);
nand UO_2753 (O_2753,N_29055,N_29885);
nand UO_2754 (O_2754,N_29765,N_29704);
and UO_2755 (O_2755,N_29244,N_29172);
or UO_2756 (O_2756,N_29922,N_29624);
xor UO_2757 (O_2757,N_29626,N_29663);
nor UO_2758 (O_2758,N_29699,N_29959);
or UO_2759 (O_2759,N_29012,N_29296);
xnor UO_2760 (O_2760,N_29847,N_29134);
nand UO_2761 (O_2761,N_29520,N_29353);
or UO_2762 (O_2762,N_29941,N_29005);
or UO_2763 (O_2763,N_29427,N_29117);
nand UO_2764 (O_2764,N_29253,N_29512);
nand UO_2765 (O_2765,N_29010,N_29143);
nor UO_2766 (O_2766,N_29000,N_29592);
nor UO_2767 (O_2767,N_29319,N_29399);
xor UO_2768 (O_2768,N_29224,N_29910);
nand UO_2769 (O_2769,N_29740,N_29577);
and UO_2770 (O_2770,N_29835,N_29643);
xnor UO_2771 (O_2771,N_29671,N_29365);
or UO_2772 (O_2772,N_29929,N_29517);
or UO_2773 (O_2773,N_29736,N_29917);
and UO_2774 (O_2774,N_29972,N_29375);
nor UO_2775 (O_2775,N_29981,N_29578);
or UO_2776 (O_2776,N_29196,N_29040);
or UO_2777 (O_2777,N_29696,N_29522);
xnor UO_2778 (O_2778,N_29633,N_29366);
nand UO_2779 (O_2779,N_29921,N_29235);
xor UO_2780 (O_2780,N_29800,N_29854);
and UO_2781 (O_2781,N_29784,N_29422);
and UO_2782 (O_2782,N_29600,N_29855);
and UO_2783 (O_2783,N_29604,N_29711);
nand UO_2784 (O_2784,N_29885,N_29554);
xor UO_2785 (O_2785,N_29499,N_29856);
nor UO_2786 (O_2786,N_29634,N_29397);
and UO_2787 (O_2787,N_29882,N_29673);
nor UO_2788 (O_2788,N_29448,N_29193);
nand UO_2789 (O_2789,N_29183,N_29845);
or UO_2790 (O_2790,N_29344,N_29785);
or UO_2791 (O_2791,N_29969,N_29610);
and UO_2792 (O_2792,N_29252,N_29959);
or UO_2793 (O_2793,N_29168,N_29969);
and UO_2794 (O_2794,N_29168,N_29029);
nand UO_2795 (O_2795,N_29326,N_29371);
and UO_2796 (O_2796,N_29391,N_29511);
nor UO_2797 (O_2797,N_29414,N_29926);
nand UO_2798 (O_2798,N_29908,N_29240);
xnor UO_2799 (O_2799,N_29073,N_29857);
or UO_2800 (O_2800,N_29434,N_29074);
xor UO_2801 (O_2801,N_29381,N_29477);
nand UO_2802 (O_2802,N_29338,N_29181);
nand UO_2803 (O_2803,N_29638,N_29696);
and UO_2804 (O_2804,N_29816,N_29593);
xnor UO_2805 (O_2805,N_29897,N_29430);
nand UO_2806 (O_2806,N_29593,N_29577);
and UO_2807 (O_2807,N_29101,N_29580);
and UO_2808 (O_2808,N_29355,N_29683);
xor UO_2809 (O_2809,N_29177,N_29379);
and UO_2810 (O_2810,N_29647,N_29691);
xnor UO_2811 (O_2811,N_29736,N_29547);
nand UO_2812 (O_2812,N_29653,N_29112);
nand UO_2813 (O_2813,N_29487,N_29920);
or UO_2814 (O_2814,N_29785,N_29854);
and UO_2815 (O_2815,N_29729,N_29641);
or UO_2816 (O_2816,N_29313,N_29016);
nor UO_2817 (O_2817,N_29877,N_29007);
and UO_2818 (O_2818,N_29476,N_29875);
xnor UO_2819 (O_2819,N_29403,N_29611);
or UO_2820 (O_2820,N_29052,N_29767);
nor UO_2821 (O_2821,N_29174,N_29526);
xor UO_2822 (O_2822,N_29478,N_29732);
and UO_2823 (O_2823,N_29446,N_29022);
nand UO_2824 (O_2824,N_29885,N_29188);
and UO_2825 (O_2825,N_29011,N_29322);
and UO_2826 (O_2826,N_29423,N_29299);
xnor UO_2827 (O_2827,N_29349,N_29757);
nor UO_2828 (O_2828,N_29601,N_29533);
nand UO_2829 (O_2829,N_29002,N_29894);
xnor UO_2830 (O_2830,N_29377,N_29808);
xor UO_2831 (O_2831,N_29184,N_29438);
nand UO_2832 (O_2832,N_29312,N_29324);
xnor UO_2833 (O_2833,N_29154,N_29029);
and UO_2834 (O_2834,N_29132,N_29201);
nor UO_2835 (O_2835,N_29616,N_29928);
xnor UO_2836 (O_2836,N_29583,N_29981);
nand UO_2837 (O_2837,N_29326,N_29101);
and UO_2838 (O_2838,N_29546,N_29402);
and UO_2839 (O_2839,N_29198,N_29233);
nand UO_2840 (O_2840,N_29280,N_29910);
nor UO_2841 (O_2841,N_29605,N_29025);
nand UO_2842 (O_2842,N_29520,N_29235);
or UO_2843 (O_2843,N_29064,N_29162);
and UO_2844 (O_2844,N_29234,N_29958);
or UO_2845 (O_2845,N_29817,N_29343);
nand UO_2846 (O_2846,N_29374,N_29033);
xnor UO_2847 (O_2847,N_29684,N_29813);
xnor UO_2848 (O_2848,N_29539,N_29683);
and UO_2849 (O_2849,N_29056,N_29139);
and UO_2850 (O_2850,N_29572,N_29771);
nand UO_2851 (O_2851,N_29159,N_29626);
nor UO_2852 (O_2852,N_29023,N_29042);
xnor UO_2853 (O_2853,N_29691,N_29252);
xnor UO_2854 (O_2854,N_29487,N_29870);
and UO_2855 (O_2855,N_29568,N_29744);
nor UO_2856 (O_2856,N_29178,N_29145);
nor UO_2857 (O_2857,N_29631,N_29142);
nand UO_2858 (O_2858,N_29733,N_29376);
xor UO_2859 (O_2859,N_29955,N_29571);
nor UO_2860 (O_2860,N_29319,N_29314);
or UO_2861 (O_2861,N_29225,N_29795);
or UO_2862 (O_2862,N_29572,N_29441);
nor UO_2863 (O_2863,N_29440,N_29448);
nand UO_2864 (O_2864,N_29681,N_29586);
nor UO_2865 (O_2865,N_29427,N_29984);
nor UO_2866 (O_2866,N_29621,N_29040);
and UO_2867 (O_2867,N_29948,N_29066);
xnor UO_2868 (O_2868,N_29647,N_29648);
xnor UO_2869 (O_2869,N_29013,N_29758);
xor UO_2870 (O_2870,N_29261,N_29919);
or UO_2871 (O_2871,N_29667,N_29481);
xor UO_2872 (O_2872,N_29964,N_29497);
xor UO_2873 (O_2873,N_29480,N_29142);
nand UO_2874 (O_2874,N_29836,N_29088);
nand UO_2875 (O_2875,N_29752,N_29253);
and UO_2876 (O_2876,N_29759,N_29812);
nor UO_2877 (O_2877,N_29965,N_29432);
nor UO_2878 (O_2878,N_29995,N_29230);
or UO_2879 (O_2879,N_29563,N_29346);
and UO_2880 (O_2880,N_29734,N_29933);
xnor UO_2881 (O_2881,N_29708,N_29238);
xor UO_2882 (O_2882,N_29379,N_29532);
nor UO_2883 (O_2883,N_29738,N_29463);
and UO_2884 (O_2884,N_29305,N_29904);
or UO_2885 (O_2885,N_29033,N_29187);
nand UO_2886 (O_2886,N_29125,N_29607);
or UO_2887 (O_2887,N_29704,N_29218);
xnor UO_2888 (O_2888,N_29838,N_29890);
nand UO_2889 (O_2889,N_29036,N_29151);
xor UO_2890 (O_2890,N_29470,N_29287);
and UO_2891 (O_2891,N_29399,N_29270);
nand UO_2892 (O_2892,N_29068,N_29749);
and UO_2893 (O_2893,N_29615,N_29177);
and UO_2894 (O_2894,N_29645,N_29115);
or UO_2895 (O_2895,N_29788,N_29340);
or UO_2896 (O_2896,N_29567,N_29357);
nand UO_2897 (O_2897,N_29943,N_29354);
xnor UO_2898 (O_2898,N_29163,N_29715);
nand UO_2899 (O_2899,N_29668,N_29256);
and UO_2900 (O_2900,N_29057,N_29183);
and UO_2901 (O_2901,N_29433,N_29007);
nand UO_2902 (O_2902,N_29960,N_29785);
and UO_2903 (O_2903,N_29104,N_29427);
nand UO_2904 (O_2904,N_29920,N_29425);
xor UO_2905 (O_2905,N_29521,N_29431);
nand UO_2906 (O_2906,N_29771,N_29551);
nand UO_2907 (O_2907,N_29745,N_29121);
or UO_2908 (O_2908,N_29281,N_29536);
or UO_2909 (O_2909,N_29978,N_29222);
nand UO_2910 (O_2910,N_29581,N_29931);
nor UO_2911 (O_2911,N_29529,N_29284);
and UO_2912 (O_2912,N_29929,N_29416);
or UO_2913 (O_2913,N_29843,N_29875);
xnor UO_2914 (O_2914,N_29233,N_29012);
and UO_2915 (O_2915,N_29309,N_29725);
and UO_2916 (O_2916,N_29296,N_29477);
nor UO_2917 (O_2917,N_29209,N_29595);
or UO_2918 (O_2918,N_29274,N_29250);
and UO_2919 (O_2919,N_29093,N_29447);
and UO_2920 (O_2920,N_29296,N_29701);
and UO_2921 (O_2921,N_29295,N_29167);
or UO_2922 (O_2922,N_29055,N_29638);
and UO_2923 (O_2923,N_29544,N_29600);
xnor UO_2924 (O_2924,N_29226,N_29129);
or UO_2925 (O_2925,N_29885,N_29615);
nor UO_2926 (O_2926,N_29779,N_29289);
or UO_2927 (O_2927,N_29542,N_29752);
nand UO_2928 (O_2928,N_29471,N_29768);
xor UO_2929 (O_2929,N_29835,N_29161);
nor UO_2930 (O_2930,N_29802,N_29184);
or UO_2931 (O_2931,N_29896,N_29367);
xnor UO_2932 (O_2932,N_29383,N_29729);
nor UO_2933 (O_2933,N_29956,N_29396);
nand UO_2934 (O_2934,N_29510,N_29893);
nor UO_2935 (O_2935,N_29531,N_29000);
nand UO_2936 (O_2936,N_29773,N_29356);
or UO_2937 (O_2937,N_29893,N_29505);
xnor UO_2938 (O_2938,N_29255,N_29230);
and UO_2939 (O_2939,N_29490,N_29881);
or UO_2940 (O_2940,N_29294,N_29135);
nor UO_2941 (O_2941,N_29668,N_29118);
nor UO_2942 (O_2942,N_29917,N_29032);
xor UO_2943 (O_2943,N_29255,N_29765);
and UO_2944 (O_2944,N_29508,N_29765);
xnor UO_2945 (O_2945,N_29042,N_29147);
and UO_2946 (O_2946,N_29285,N_29811);
or UO_2947 (O_2947,N_29455,N_29146);
or UO_2948 (O_2948,N_29869,N_29323);
xor UO_2949 (O_2949,N_29782,N_29324);
and UO_2950 (O_2950,N_29957,N_29984);
xnor UO_2951 (O_2951,N_29229,N_29945);
nand UO_2952 (O_2952,N_29271,N_29444);
nand UO_2953 (O_2953,N_29333,N_29190);
and UO_2954 (O_2954,N_29915,N_29663);
nand UO_2955 (O_2955,N_29998,N_29366);
nand UO_2956 (O_2956,N_29270,N_29299);
nand UO_2957 (O_2957,N_29013,N_29017);
nor UO_2958 (O_2958,N_29633,N_29321);
nor UO_2959 (O_2959,N_29411,N_29464);
nand UO_2960 (O_2960,N_29057,N_29120);
or UO_2961 (O_2961,N_29413,N_29168);
or UO_2962 (O_2962,N_29728,N_29573);
and UO_2963 (O_2963,N_29353,N_29132);
or UO_2964 (O_2964,N_29000,N_29861);
or UO_2965 (O_2965,N_29315,N_29664);
xnor UO_2966 (O_2966,N_29223,N_29196);
nor UO_2967 (O_2967,N_29284,N_29129);
and UO_2968 (O_2968,N_29358,N_29272);
nand UO_2969 (O_2969,N_29117,N_29396);
and UO_2970 (O_2970,N_29423,N_29124);
xnor UO_2971 (O_2971,N_29143,N_29916);
nor UO_2972 (O_2972,N_29863,N_29071);
and UO_2973 (O_2973,N_29597,N_29427);
nor UO_2974 (O_2974,N_29725,N_29439);
xnor UO_2975 (O_2975,N_29335,N_29490);
or UO_2976 (O_2976,N_29025,N_29014);
nand UO_2977 (O_2977,N_29746,N_29780);
nand UO_2978 (O_2978,N_29515,N_29254);
nand UO_2979 (O_2979,N_29402,N_29638);
nor UO_2980 (O_2980,N_29438,N_29070);
and UO_2981 (O_2981,N_29846,N_29863);
nor UO_2982 (O_2982,N_29684,N_29347);
nor UO_2983 (O_2983,N_29490,N_29207);
or UO_2984 (O_2984,N_29890,N_29646);
xor UO_2985 (O_2985,N_29322,N_29863);
nor UO_2986 (O_2986,N_29393,N_29180);
or UO_2987 (O_2987,N_29879,N_29881);
nor UO_2988 (O_2988,N_29284,N_29489);
nor UO_2989 (O_2989,N_29607,N_29925);
or UO_2990 (O_2990,N_29349,N_29072);
nor UO_2991 (O_2991,N_29452,N_29582);
or UO_2992 (O_2992,N_29235,N_29401);
nand UO_2993 (O_2993,N_29806,N_29208);
nand UO_2994 (O_2994,N_29052,N_29815);
or UO_2995 (O_2995,N_29011,N_29692);
nor UO_2996 (O_2996,N_29010,N_29546);
or UO_2997 (O_2997,N_29112,N_29004);
nor UO_2998 (O_2998,N_29447,N_29809);
and UO_2999 (O_2999,N_29003,N_29719);
and UO_3000 (O_3000,N_29527,N_29116);
or UO_3001 (O_3001,N_29177,N_29948);
and UO_3002 (O_3002,N_29724,N_29352);
nor UO_3003 (O_3003,N_29811,N_29051);
and UO_3004 (O_3004,N_29290,N_29417);
and UO_3005 (O_3005,N_29348,N_29297);
and UO_3006 (O_3006,N_29656,N_29450);
and UO_3007 (O_3007,N_29061,N_29818);
and UO_3008 (O_3008,N_29627,N_29704);
nand UO_3009 (O_3009,N_29315,N_29502);
and UO_3010 (O_3010,N_29864,N_29911);
nand UO_3011 (O_3011,N_29199,N_29619);
and UO_3012 (O_3012,N_29866,N_29518);
or UO_3013 (O_3013,N_29513,N_29881);
nand UO_3014 (O_3014,N_29315,N_29524);
or UO_3015 (O_3015,N_29581,N_29053);
nand UO_3016 (O_3016,N_29004,N_29662);
xor UO_3017 (O_3017,N_29332,N_29579);
xor UO_3018 (O_3018,N_29126,N_29794);
xor UO_3019 (O_3019,N_29223,N_29733);
nand UO_3020 (O_3020,N_29794,N_29147);
or UO_3021 (O_3021,N_29383,N_29940);
or UO_3022 (O_3022,N_29400,N_29699);
and UO_3023 (O_3023,N_29713,N_29856);
xor UO_3024 (O_3024,N_29144,N_29432);
nor UO_3025 (O_3025,N_29261,N_29390);
nor UO_3026 (O_3026,N_29479,N_29954);
nand UO_3027 (O_3027,N_29662,N_29397);
or UO_3028 (O_3028,N_29766,N_29607);
nand UO_3029 (O_3029,N_29938,N_29275);
nand UO_3030 (O_3030,N_29916,N_29793);
nor UO_3031 (O_3031,N_29684,N_29788);
xor UO_3032 (O_3032,N_29055,N_29356);
or UO_3033 (O_3033,N_29578,N_29337);
and UO_3034 (O_3034,N_29862,N_29020);
or UO_3035 (O_3035,N_29972,N_29566);
xnor UO_3036 (O_3036,N_29802,N_29308);
and UO_3037 (O_3037,N_29254,N_29968);
nor UO_3038 (O_3038,N_29815,N_29864);
or UO_3039 (O_3039,N_29508,N_29942);
and UO_3040 (O_3040,N_29891,N_29038);
nand UO_3041 (O_3041,N_29045,N_29285);
xnor UO_3042 (O_3042,N_29319,N_29542);
or UO_3043 (O_3043,N_29732,N_29901);
nor UO_3044 (O_3044,N_29480,N_29973);
nor UO_3045 (O_3045,N_29878,N_29133);
and UO_3046 (O_3046,N_29177,N_29009);
or UO_3047 (O_3047,N_29511,N_29748);
and UO_3048 (O_3048,N_29774,N_29225);
xnor UO_3049 (O_3049,N_29749,N_29405);
and UO_3050 (O_3050,N_29382,N_29427);
nand UO_3051 (O_3051,N_29499,N_29313);
nor UO_3052 (O_3052,N_29702,N_29416);
or UO_3053 (O_3053,N_29251,N_29686);
or UO_3054 (O_3054,N_29864,N_29495);
nor UO_3055 (O_3055,N_29018,N_29626);
nor UO_3056 (O_3056,N_29327,N_29969);
xor UO_3057 (O_3057,N_29615,N_29779);
xnor UO_3058 (O_3058,N_29584,N_29337);
xor UO_3059 (O_3059,N_29768,N_29509);
or UO_3060 (O_3060,N_29944,N_29166);
nor UO_3061 (O_3061,N_29096,N_29044);
and UO_3062 (O_3062,N_29741,N_29243);
nor UO_3063 (O_3063,N_29626,N_29036);
xor UO_3064 (O_3064,N_29143,N_29973);
nor UO_3065 (O_3065,N_29720,N_29613);
nor UO_3066 (O_3066,N_29821,N_29967);
nand UO_3067 (O_3067,N_29475,N_29487);
or UO_3068 (O_3068,N_29428,N_29912);
and UO_3069 (O_3069,N_29736,N_29016);
xnor UO_3070 (O_3070,N_29374,N_29310);
nor UO_3071 (O_3071,N_29807,N_29477);
and UO_3072 (O_3072,N_29697,N_29796);
xor UO_3073 (O_3073,N_29698,N_29492);
nand UO_3074 (O_3074,N_29739,N_29800);
or UO_3075 (O_3075,N_29842,N_29998);
nand UO_3076 (O_3076,N_29932,N_29812);
or UO_3077 (O_3077,N_29828,N_29454);
and UO_3078 (O_3078,N_29024,N_29040);
xor UO_3079 (O_3079,N_29205,N_29030);
nand UO_3080 (O_3080,N_29902,N_29307);
or UO_3081 (O_3081,N_29353,N_29879);
xnor UO_3082 (O_3082,N_29300,N_29575);
and UO_3083 (O_3083,N_29048,N_29192);
or UO_3084 (O_3084,N_29261,N_29711);
or UO_3085 (O_3085,N_29442,N_29142);
nor UO_3086 (O_3086,N_29882,N_29499);
and UO_3087 (O_3087,N_29840,N_29683);
and UO_3088 (O_3088,N_29312,N_29909);
nor UO_3089 (O_3089,N_29631,N_29841);
or UO_3090 (O_3090,N_29315,N_29855);
nand UO_3091 (O_3091,N_29038,N_29957);
nand UO_3092 (O_3092,N_29194,N_29617);
or UO_3093 (O_3093,N_29501,N_29651);
nor UO_3094 (O_3094,N_29436,N_29283);
and UO_3095 (O_3095,N_29893,N_29700);
or UO_3096 (O_3096,N_29664,N_29674);
nor UO_3097 (O_3097,N_29085,N_29873);
nand UO_3098 (O_3098,N_29226,N_29220);
xnor UO_3099 (O_3099,N_29461,N_29643);
or UO_3100 (O_3100,N_29603,N_29027);
nor UO_3101 (O_3101,N_29840,N_29566);
or UO_3102 (O_3102,N_29472,N_29388);
and UO_3103 (O_3103,N_29031,N_29890);
and UO_3104 (O_3104,N_29027,N_29577);
nor UO_3105 (O_3105,N_29326,N_29998);
or UO_3106 (O_3106,N_29782,N_29353);
nor UO_3107 (O_3107,N_29634,N_29709);
nor UO_3108 (O_3108,N_29198,N_29846);
or UO_3109 (O_3109,N_29809,N_29628);
and UO_3110 (O_3110,N_29838,N_29002);
nor UO_3111 (O_3111,N_29212,N_29426);
nand UO_3112 (O_3112,N_29888,N_29307);
xor UO_3113 (O_3113,N_29583,N_29126);
and UO_3114 (O_3114,N_29947,N_29563);
or UO_3115 (O_3115,N_29040,N_29488);
xnor UO_3116 (O_3116,N_29077,N_29706);
nor UO_3117 (O_3117,N_29229,N_29115);
and UO_3118 (O_3118,N_29381,N_29134);
xor UO_3119 (O_3119,N_29526,N_29216);
or UO_3120 (O_3120,N_29153,N_29160);
nor UO_3121 (O_3121,N_29846,N_29373);
or UO_3122 (O_3122,N_29701,N_29730);
or UO_3123 (O_3123,N_29887,N_29964);
nor UO_3124 (O_3124,N_29097,N_29268);
xor UO_3125 (O_3125,N_29985,N_29695);
nand UO_3126 (O_3126,N_29526,N_29824);
and UO_3127 (O_3127,N_29877,N_29656);
or UO_3128 (O_3128,N_29734,N_29607);
nand UO_3129 (O_3129,N_29666,N_29843);
nand UO_3130 (O_3130,N_29923,N_29181);
and UO_3131 (O_3131,N_29342,N_29187);
nand UO_3132 (O_3132,N_29074,N_29491);
or UO_3133 (O_3133,N_29380,N_29501);
xor UO_3134 (O_3134,N_29509,N_29879);
or UO_3135 (O_3135,N_29262,N_29415);
and UO_3136 (O_3136,N_29684,N_29991);
xnor UO_3137 (O_3137,N_29422,N_29731);
nor UO_3138 (O_3138,N_29534,N_29314);
nor UO_3139 (O_3139,N_29940,N_29495);
and UO_3140 (O_3140,N_29366,N_29204);
and UO_3141 (O_3141,N_29118,N_29708);
nand UO_3142 (O_3142,N_29932,N_29806);
nor UO_3143 (O_3143,N_29212,N_29413);
nand UO_3144 (O_3144,N_29545,N_29709);
and UO_3145 (O_3145,N_29947,N_29839);
and UO_3146 (O_3146,N_29511,N_29333);
nand UO_3147 (O_3147,N_29060,N_29015);
nand UO_3148 (O_3148,N_29110,N_29730);
xnor UO_3149 (O_3149,N_29388,N_29086);
nand UO_3150 (O_3150,N_29535,N_29452);
nand UO_3151 (O_3151,N_29283,N_29037);
xnor UO_3152 (O_3152,N_29330,N_29293);
nor UO_3153 (O_3153,N_29587,N_29314);
nand UO_3154 (O_3154,N_29904,N_29579);
xor UO_3155 (O_3155,N_29320,N_29628);
nand UO_3156 (O_3156,N_29274,N_29979);
and UO_3157 (O_3157,N_29473,N_29045);
or UO_3158 (O_3158,N_29917,N_29127);
and UO_3159 (O_3159,N_29482,N_29625);
nand UO_3160 (O_3160,N_29469,N_29394);
and UO_3161 (O_3161,N_29068,N_29460);
nor UO_3162 (O_3162,N_29465,N_29308);
nor UO_3163 (O_3163,N_29117,N_29401);
and UO_3164 (O_3164,N_29661,N_29926);
or UO_3165 (O_3165,N_29907,N_29164);
and UO_3166 (O_3166,N_29042,N_29701);
or UO_3167 (O_3167,N_29573,N_29579);
and UO_3168 (O_3168,N_29589,N_29089);
and UO_3169 (O_3169,N_29195,N_29393);
or UO_3170 (O_3170,N_29235,N_29689);
nand UO_3171 (O_3171,N_29494,N_29303);
nand UO_3172 (O_3172,N_29917,N_29954);
nand UO_3173 (O_3173,N_29791,N_29656);
and UO_3174 (O_3174,N_29848,N_29832);
and UO_3175 (O_3175,N_29119,N_29719);
and UO_3176 (O_3176,N_29921,N_29341);
xor UO_3177 (O_3177,N_29846,N_29515);
or UO_3178 (O_3178,N_29894,N_29462);
and UO_3179 (O_3179,N_29534,N_29558);
or UO_3180 (O_3180,N_29241,N_29146);
xor UO_3181 (O_3181,N_29867,N_29713);
nor UO_3182 (O_3182,N_29255,N_29544);
xor UO_3183 (O_3183,N_29203,N_29676);
xnor UO_3184 (O_3184,N_29674,N_29517);
nand UO_3185 (O_3185,N_29877,N_29964);
or UO_3186 (O_3186,N_29182,N_29484);
nand UO_3187 (O_3187,N_29915,N_29337);
nand UO_3188 (O_3188,N_29310,N_29077);
nand UO_3189 (O_3189,N_29997,N_29102);
xnor UO_3190 (O_3190,N_29229,N_29208);
and UO_3191 (O_3191,N_29910,N_29314);
nor UO_3192 (O_3192,N_29179,N_29928);
and UO_3193 (O_3193,N_29227,N_29410);
or UO_3194 (O_3194,N_29670,N_29513);
and UO_3195 (O_3195,N_29098,N_29600);
xnor UO_3196 (O_3196,N_29327,N_29850);
xnor UO_3197 (O_3197,N_29625,N_29129);
nand UO_3198 (O_3198,N_29086,N_29869);
nand UO_3199 (O_3199,N_29079,N_29641);
nand UO_3200 (O_3200,N_29120,N_29526);
and UO_3201 (O_3201,N_29803,N_29983);
or UO_3202 (O_3202,N_29983,N_29072);
and UO_3203 (O_3203,N_29138,N_29051);
xnor UO_3204 (O_3204,N_29186,N_29288);
xnor UO_3205 (O_3205,N_29213,N_29690);
and UO_3206 (O_3206,N_29822,N_29705);
nand UO_3207 (O_3207,N_29755,N_29209);
nand UO_3208 (O_3208,N_29836,N_29524);
and UO_3209 (O_3209,N_29311,N_29820);
xnor UO_3210 (O_3210,N_29184,N_29535);
xor UO_3211 (O_3211,N_29597,N_29962);
nor UO_3212 (O_3212,N_29559,N_29659);
and UO_3213 (O_3213,N_29103,N_29629);
nand UO_3214 (O_3214,N_29336,N_29851);
or UO_3215 (O_3215,N_29866,N_29731);
or UO_3216 (O_3216,N_29243,N_29693);
or UO_3217 (O_3217,N_29673,N_29213);
or UO_3218 (O_3218,N_29541,N_29636);
and UO_3219 (O_3219,N_29289,N_29471);
nor UO_3220 (O_3220,N_29899,N_29509);
xnor UO_3221 (O_3221,N_29086,N_29885);
or UO_3222 (O_3222,N_29520,N_29636);
xnor UO_3223 (O_3223,N_29833,N_29109);
nand UO_3224 (O_3224,N_29176,N_29205);
or UO_3225 (O_3225,N_29590,N_29838);
xnor UO_3226 (O_3226,N_29312,N_29534);
nor UO_3227 (O_3227,N_29829,N_29306);
nor UO_3228 (O_3228,N_29524,N_29537);
or UO_3229 (O_3229,N_29474,N_29731);
xor UO_3230 (O_3230,N_29777,N_29895);
or UO_3231 (O_3231,N_29375,N_29203);
and UO_3232 (O_3232,N_29282,N_29738);
and UO_3233 (O_3233,N_29127,N_29904);
xor UO_3234 (O_3234,N_29766,N_29938);
and UO_3235 (O_3235,N_29682,N_29568);
xnor UO_3236 (O_3236,N_29814,N_29231);
and UO_3237 (O_3237,N_29996,N_29427);
nand UO_3238 (O_3238,N_29889,N_29303);
xor UO_3239 (O_3239,N_29474,N_29793);
and UO_3240 (O_3240,N_29671,N_29063);
xnor UO_3241 (O_3241,N_29817,N_29661);
and UO_3242 (O_3242,N_29313,N_29804);
and UO_3243 (O_3243,N_29036,N_29322);
xnor UO_3244 (O_3244,N_29554,N_29028);
nor UO_3245 (O_3245,N_29051,N_29091);
xor UO_3246 (O_3246,N_29676,N_29085);
and UO_3247 (O_3247,N_29121,N_29076);
nor UO_3248 (O_3248,N_29226,N_29726);
or UO_3249 (O_3249,N_29432,N_29443);
or UO_3250 (O_3250,N_29055,N_29288);
and UO_3251 (O_3251,N_29694,N_29931);
and UO_3252 (O_3252,N_29347,N_29828);
or UO_3253 (O_3253,N_29744,N_29543);
or UO_3254 (O_3254,N_29215,N_29486);
xnor UO_3255 (O_3255,N_29500,N_29368);
nor UO_3256 (O_3256,N_29263,N_29605);
or UO_3257 (O_3257,N_29538,N_29031);
xor UO_3258 (O_3258,N_29360,N_29262);
or UO_3259 (O_3259,N_29384,N_29713);
nand UO_3260 (O_3260,N_29368,N_29670);
and UO_3261 (O_3261,N_29748,N_29785);
or UO_3262 (O_3262,N_29102,N_29006);
nand UO_3263 (O_3263,N_29837,N_29497);
and UO_3264 (O_3264,N_29843,N_29931);
xor UO_3265 (O_3265,N_29939,N_29515);
or UO_3266 (O_3266,N_29275,N_29907);
and UO_3267 (O_3267,N_29813,N_29228);
nand UO_3268 (O_3268,N_29951,N_29669);
nor UO_3269 (O_3269,N_29542,N_29443);
xnor UO_3270 (O_3270,N_29720,N_29287);
xor UO_3271 (O_3271,N_29519,N_29152);
nor UO_3272 (O_3272,N_29240,N_29463);
and UO_3273 (O_3273,N_29531,N_29491);
nor UO_3274 (O_3274,N_29601,N_29169);
nand UO_3275 (O_3275,N_29900,N_29566);
xnor UO_3276 (O_3276,N_29484,N_29158);
or UO_3277 (O_3277,N_29924,N_29019);
or UO_3278 (O_3278,N_29795,N_29360);
or UO_3279 (O_3279,N_29925,N_29759);
nand UO_3280 (O_3280,N_29561,N_29271);
xnor UO_3281 (O_3281,N_29321,N_29518);
or UO_3282 (O_3282,N_29045,N_29513);
or UO_3283 (O_3283,N_29950,N_29236);
xor UO_3284 (O_3284,N_29030,N_29718);
or UO_3285 (O_3285,N_29154,N_29156);
nand UO_3286 (O_3286,N_29720,N_29298);
nor UO_3287 (O_3287,N_29774,N_29612);
xnor UO_3288 (O_3288,N_29835,N_29824);
xor UO_3289 (O_3289,N_29342,N_29419);
nand UO_3290 (O_3290,N_29856,N_29824);
and UO_3291 (O_3291,N_29850,N_29299);
and UO_3292 (O_3292,N_29007,N_29131);
nand UO_3293 (O_3293,N_29437,N_29730);
nand UO_3294 (O_3294,N_29549,N_29292);
or UO_3295 (O_3295,N_29321,N_29468);
nand UO_3296 (O_3296,N_29878,N_29843);
nor UO_3297 (O_3297,N_29523,N_29118);
and UO_3298 (O_3298,N_29876,N_29102);
nor UO_3299 (O_3299,N_29401,N_29626);
xor UO_3300 (O_3300,N_29208,N_29898);
and UO_3301 (O_3301,N_29014,N_29472);
and UO_3302 (O_3302,N_29156,N_29311);
and UO_3303 (O_3303,N_29004,N_29019);
nand UO_3304 (O_3304,N_29298,N_29384);
or UO_3305 (O_3305,N_29941,N_29690);
nor UO_3306 (O_3306,N_29864,N_29706);
or UO_3307 (O_3307,N_29307,N_29394);
xor UO_3308 (O_3308,N_29343,N_29752);
xnor UO_3309 (O_3309,N_29062,N_29494);
nor UO_3310 (O_3310,N_29618,N_29488);
nand UO_3311 (O_3311,N_29746,N_29874);
and UO_3312 (O_3312,N_29275,N_29918);
and UO_3313 (O_3313,N_29319,N_29270);
and UO_3314 (O_3314,N_29109,N_29744);
nand UO_3315 (O_3315,N_29637,N_29385);
xor UO_3316 (O_3316,N_29599,N_29388);
or UO_3317 (O_3317,N_29657,N_29253);
nor UO_3318 (O_3318,N_29161,N_29308);
nor UO_3319 (O_3319,N_29373,N_29670);
and UO_3320 (O_3320,N_29747,N_29856);
nand UO_3321 (O_3321,N_29187,N_29882);
nor UO_3322 (O_3322,N_29637,N_29513);
or UO_3323 (O_3323,N_29316,N_29902);
or UO_3324 (O_3324,N_29347,N_29624);
and UO_3325 (O_3325,N_29669,N_29164);
nand UO_3326 (O_3326,N_29684,N_29059);
and UO_3327 (O_3327,N_29717,N_29983);
xor UO_3328 (O_3328,N_29546,N_29235);
or UO_3329 (O_3329,N_29993,N_29482);
nand UO_3330 (O_3330,N_29833,N_29370);
or UO_3331 (O_3331,N_29905,N_29880);
and UO_3332 (O_3332,N_29977,N_29218);
xor UO_3333 (O_3333,N_29798,N_29516);
nand UO_3334 (O_3334,N_29692,N_29849);
nor UO_3335 (O_3335,N_29176,N_29771);
or UO_3336 (O_3336,N_29334,N_29459);
and UO_3337 (O_3337,N_29766,N_29297);
xor UO_3338 (O_3338,N_29319,N_29726);
or UO_3339 (O_3339,N_29522,N_29253);
and UO_3340 (O_3340,N_29073,N_29887);
and UO_3341 (O_3341,N_29306,N_29198);
and UO_3342 (O_3342,N_29552,N_29171);
xnor UO_3343 (O_3343,N_29055,N_29451);
or UO_3344 (O_3344,N_29142,N_29000);
nor UO_3345 (O_3345,N_29913,N_29891);
or UO_3346 (O_3346,N_29096,N_29926);
or UO_3347 (O_3347,N_29340,N_29485);
nor UO_3348 (O_3348,N_29150,N_29649);
nor UO_3349 (O_3349,N_29209,N_29294);
xnor UO_3350 (O_3350,N_29822,N_29037);
nand UO_3351 (O_3351,N_29284,N_29598);
xor UO_3352 (O_3352,N_29630,N_29139);
xor UO_3353 (O_3353,N_29682,N_29124);
or UO_3354 (O_3354,N_29406,N_29299);
and UO_3355 (O_3355,N_29592,N_29482);
and UO_3356 (O_3356,N_29156,N_29133);
or UO_3357 (O_3357,N_29599,N_29127);
nand UO_3358 (O_3358,N_29678,N_29993);
or UO_3359 (O_3359,N_29696,N_29281);
and UO_3360 (O_3360,N_29802,N_29425);
and UO_3361 (O_3361,N_29468,N_29081);
and UO_3362 (O_3362,N_29710,N_29396);
xnor UO_3363 (O_3363,N_29028,N_29510);
xnor UO_3364 (O_3364,N_29818,N_29422);
or UO_3365 (O_3365,N_29460,N_29797);
and UO_3366 (O_3366,N_29027,N_29730);
and UO_3367 (O_3367,N_29505,N_29808);
nor UO_3368 (O_3368,N_29980,N_29290);
and UO_3369 (O_3369,N_29133,N_29915);
and UO_3370 (O_3370,N_29537,N_29133);
and UO_3371 (O_3371,N_29318,N_29221);
xnor UO_3372 (O_3372,N_29861,N_29326);
and UO_3373 (O_3373,N_29667,N_29375);
xor UO_3374 (O_3374,N_29107,N_29201);
xnor UO_3375 (O_3375,N_29433,N_29602);
nand UO_3376 (O_3376,N_29845,N_29588);
nand UO_3377 (O_3377,N_29597,N_29960);
nand UO_3378 (O_3378,N_29771,N_29738);
nand UO_3379 (O_3379,N_29373,N_29192);
xnor UO_3380 (O_3380,N_29583,N_29740);
or UO_3381 (O_3381,N_29991,N_29706);
nand UO_3382 (O_3382,N_29497,N_29344);
xor UO_3383 (O_3383,N_29079,N_29105);
and UO_3384 (O_3384,N_29266,N_29536);
or UO_3385 (O_3385,N_29681,N_29625);
and UO_3386 (O_3386,N_29172,N_29698);
and UO_3387 (O_3387,N_29417,N_29814);
xor UO_3388 (O_3388,N_29433,N_29399);
and UO_3389 (O_3389,N_29394,N_29025);
nor UO_3390 (O_3390,N_29144,N_29387);
xnor UO_3391 (O_3391,N_29014,N_29060);
nor UO_3392 (O_3392,N_29744,N_29525);
or UO_3393 (O_3393,N_29546,N_29595);
xnor UO_3394 (O_3394,N_29070,N_29380);
nand UO_3395 (O_3395,N_29994,N_29855);
nand UO_3396 (O_3396,N_29428,N_29708);
and UO_3397 (O_3397,N_29049,N_29999);
nand UO_3398 (O_3398,N_29245,N_29306);
nor UO_3399 (O_3399,N_29164,N_29447);
or UO_3400 (O_3400,N_29290,N_29598);
xor UO_3401 (O_3401,N_29607,N_29202);
nor UO_3402 (O_3402,N_29181,N_29367);
and UO_3403 (O_3403,N_29809,N_29245);
xor UO_3404 (O_3404,N_29187,N_29936);
and UO_3405 (O_3405,N_29760,N_29259);
nand UO_3406 (O_3406,N_29696,N_29115);
xor UO_3407 (O_3407,N_29256,N_29820);
or UO_3408 (O_3408,N_29275,N_29948);
nor UO_3409 (O_3409,N_29386,N_29512);
nand UO_3410 (O_3410,N_29348,N_29774);
xor UO_3411 (O_3411,N_29376,N_29805);
or UO_3412 (O_3412,N_29990,N_29389);
and UO_3413 (O_3413,N_29771,N_29168);
nor UO_3414 (O_3414,N_29459,N_29977);
xnor UO_3415 (O_3415,N_29770,N_29486);
and UO_3416 (O_3416,N_29649,N_29862);
or UO_3417 (O_3417,N_29150,N_29809);
nand UO_3418 (O_3418,N_29496,N_29695);
or UO_3419 (O_3419,N_29589,N_29496);
nor UO_3420 (O_3420,N_29680,N_29836);
xnor UO_3421 (O_3421,N_29904,N_29892);
xor UO_3422 (O_3422,N_29156,N_29746);
and UO_3423 (O_3423,N_29975,N_29366);
or UO_3424 (O_3424,N_29494,N_29616);
nand UO_3425 (O_3425,N_29815,N_29542);
and UO_3426 (O_3426,N_29197,N_29702);
xnor UO_3427 (O_3427,N_29374,N_29535);
xnor UO_3428 (O_3428,N_29089,N_29532);
xnor UO_3429 (O_3429,N_29433,N_29226);
xnor UO_3430 (O_3430,N_29639,N_29574);
or UO_3431 (O_3431,N_29113,N_29989);
and UO_3432 (O_3432,N_29678,N_29297);
and UO_3433 (O_3433,N_29868,N_29837);
and UO_3434 (O_3434,N_29748,N_29199);
nor UO_3435 (O_3435,N_29365,N_29540);
and UO_3436 (O_3436,N_29522,N_29189);
nor UO_3437 (O_3437,N_29060,N_29942);
nand UO_3438 (O_3438,N_29764,N_29525);
nor UO_3439 (O_3439,N_29462,N_29022);
nor UO_3440 (O_3440,N_29038,N_29982);
xor UO_3441 (O_3441,N_29897,N_29917);
nor UO_3442 (O_3442,N_29114,N_29619);
nor UO_3443 (O_3443,N_29952,N_29753);
or UO_3444 (O_3444,N_29575,N_29394);
nand UO_3445 (O_3445,N_29568,N_29902);
xor UO_3446 (O_3446,N_29841,N_29944);
and UO_3447 (O_3447,N_29622,N_29736);
and UO_3448 (O_3448,N_29092,N_29435);
nor UO_3449 (O_3449,N_29968,N_29883);
nand UO_3450 (O_3450,N_29649,N_29156);
nand UO_3451 (O_3451,N_29299,N_29160);
nand UO_3452 (O_3452,N_29516,N_29667);
nand UO_3453 (O_3453,N_29195,N_29561);
xnor UO_3454 (O_3454,N_29266,N_29336);
and UO_3455 (O_3455,N_29458,N_29223);
and UO_3456 (O_3456,N_29518,N_29166);
or UO_3457 (O_3457,N_29187,N_29635);
and UO_3458 (O_3458,N_29934,N_29113);
nor UO_3459 (O_3459,N_29497,N_29451);
or UO_3460 (O_3460,N_29343,N_29704);
nand UO_3461 (O_3461,N_29899,N_29855);
and UO_3462 (O_3462,N_29767,N_29795);
or UO_3463 (O_3463,N_29961,N_29181);
xnor UO_3464 (O_3464,N_29087,N_29507);
nor UO_3465 (O_3465,N_29555,N_29953);
xnor UO_3466 (O_3466,N_29631,N_29368);
and UO_3467 (O_3467,N_29192,N_29367);
and UO_3468 (O_3468,N_29841,N_29518);
or UO_3469 (O_3469,N_29473,N_29471);
xnor UO_3470 (O_3470,N_29073,N_29116);
nor UO_3471 (O_3471,N_29576,N_29996);
nor UO_3472 (O_3472,N_29730,N_29788);
nor UO_3473 (O_3473,N_29523,N_29640);
nor UO_3474 (O_3474,N_29944,N_29775);
and UO_3475 (O_3475,N_29872,N_29398);
or UO_3476 (O_3476,N_29843,N_29575);
and UO_3477 (O_3477,N_29425,N_29333);
and UO_3478 (O_3478,N_29276,N_29932);
xor UO_3479 (O_3479,N_29662,N_29494);
and UO_3480 (O_3480,N_29709,N_29784);
and UO_3481 (O_3481,N_29198,N_29366);
or UO_3482 (O_3482,N_29399,N_29253);
or UO_3483 (O_3483,N_29789,N_29981);
xor UO_3484 (O_3484,N_29658,N_29745);
xor UO_3485 (O_3485,N_29569,N_29794);
or UO_3486 (O_3486,N_29699,N_29284);
xor UO_3487 (O_3487,N_29079,N_29808);
xnor UO_3488 (O_3488,N_29312,N_29703);
and UO_3489 (O_3489,N_29959,N_29847);
xor UO_3490 (O_3490,N_29528,N_29300);
or UO_3491 (O_3491,N_29416,N_29680);
and UO_3492 (O_3492,N_29143,N_29384);
xnor UO_3493 (O_3493,N_29183,N_29911);
nand UO_3494 (O_3494,N_29982,N_29401);
xor UO_3495 (O_3495,N_29005,N_29463);
nand UO_3496 (O_3496,N_29519,N_29643);
nand UO_3497 (O_3497,N_29709,N_29453);
nor UO_3498 (O_3498,N_29831,N_29611);
and UO_3499 (O_3499,N_29883,N_29043);
endmodule