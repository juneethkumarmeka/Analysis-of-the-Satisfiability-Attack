module basic_500_3000_500_50_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_0,In_269);
or U1 (N_1,In_312,In_437);
xnor U2 (N_2,In_204,In_205);
and U3 (N_3,In_348,In_111);
or U4 (N_4,In_404,In_30);
and U5 (N_5,In_153,In_243);
nor U6 (N_6,In_471,In_159);
or U7 (N_7,In_11,In_350);
and U8 (N_8,In_440,In_89);
nor U9 (N_9,In_161,In_163);
or U10 (N_10,In_219,In_317);
and U11 (N_11,In_424,In_379);
and U12 (N_12,In_18,In_431);
nand U13 (N_13,In_29,In_355);
and U14 (N_14,In_233,In_104);
or U15 (N_15,In_494,In_178);
nor U16 (N_16,In_232,In_194);
xnor U17 (N_17,In_22,In_248);
and U18 (N_18,In_287,In_139);
or U19 (N_19,In_293,In_66);
nor U20 (N_20,In_121,In_131);
nand U21 (N_21,In_419,In_462);
or U22 (N_22,In_414,In_145);
and U23 (N_23,In_127,In_260);
and U24 (N_24,In_192,In_353);
and U25 (N_25,In_169,In_439);
xor U26 (N_26,In_388,In_133);
nand U27 (N_27,In_280,In_108);
xor U28 (N_28,In_375,In_14);
nor U29 (N_29,In_210,In_25);
or U30 (N_30,In_349,In_137);
or U31 (N_31,In_92,In_495);
nand U32 (N_32,In_142,In_24);
and U33 (N_33,In_203,In_428);
or U34 (N_34,In_463,In_472);
xnor U35 (N_35,In_197,In_213);
nand U36 (N_36,In_473,In_126);
xor U37 (N_37,In_129,In_106);
or U38 (N_38,In_412,In_402);
or U39 (N_39,In_374,In_368);
nand U40 (N_40,In_271,In_228);
and U41 (N_41,In_393,In_120);
and U42 (N_42,In_32,In_158);
or U43 (N_43,In_426,In_199);
nand U44 (N_44,In_469,In_239);
nor U45 (N_45,In_125,In_427);
or U46 (N_46,In_123,In_183);
nor U47 (N_47,In_115,In_272);
or U48 (N_48,In_164,In_313);
xor U49 (N_49,In_258,In_436);
and U50 (N_50,In_324,In_267);
or U51 (N_51,In_481,In_179);
or U52 (N_52,In_52,In_177);
xnor U53 (N_53,In_377,In_144);
or U54 (N_54,In_378,In_311);
and U55 (N_55,In_67,In_300);
and U56 (N_56,In_208,In_250);
nor U57 (N_57,In_189,In_434);
nor U58 (N_58,In_284,In_455);
nand U59 (N_59,In_227,In_396);
xnor U60 (N_60,In_44,In_405);
and U61 (N_61,N_55,N_36);
or U62 (N_62,N_43,N_11);
and U63 (N_63,N_41,In_403);
nor U64 (N_64,In_61,In_279);
nand U65 (N_65,In_215,In_338);
nor U66 (N_66,In_399,In_225);
and U67 (N_67,In_372,In_451);
nor U68 (N_68,In_351,In_238);
or U69 (N_69,In_314,In_435);
or U70 (N_70,In_334,In_170);
and U71 (N_71,In_282,In_28);
nand U72 (N_72,N_23,In_480);
nand U73 (N_73,In_229,In_152);
or U74 (N_74,In_201,In_395);
nand U75 (N_75,In_217,In_460);
or U76 (N_76,In_51,N_46);
nand U77 (N_77,In_342,In_485);
nand U78 (N_78,N_50,In_397);
or U79 (N_79,In_488,In_187);
nor U80 (N_80,In_408,In_134);
nor U81 (N_81,In_332,In_9);
or U82 (N_82,In_63,N_19);
or U83 (N_83,In_482,In_200);
nand U84 (N_84,In_140,In_257);
and U85 (N_85,In_46,N_44);
or U86 (N_86,In_7,In_58);
or U87 (N_87,In_454,N_14);
nor U88 (N_88,In_291,In_433);
or U89 (N_89,In_319,In_94);
and U90 (N_90,In_222,In_336);
xor U91 (N_91,In_156,N_52);
nand U92 (N_92,In_341,In_497);
nor U93 (N_93,In_425,In_83);
nand U94 (N_94,In_172,In_162);
or U95 (N_95,In_306,In_429);
or U96 (N_96,In_268,In_36);
nand U97 (N_97,In_392,N_15);
nand U98 (N_98,In_376,In_154);
nor U99 (N_99,In_4,In_80);
or U100 (N_100,In_251,In_160);
xor U101 (N_101,In_363,In_445);
nand U102 (N_102,N_53,In_305);
and U103 (N_103,N_0,In_235);
and U104 (N_104,In_323,In_99);
nor U105 (N_105,In_68,In_491);
nand U106 (N_106,In_343,In_149);
or U107 (N_107,In_246,In_138);
xnor U108 (N_108,N_13,In_303);
or U109 (N_109,In_422,In_223);
nor U110 (N_110,In_263,N_56);
nor U111 (N_111,In_171,In_496);
or U112 (N_112,In_17,In_86);
and U113 (N_113,In_371,N_31);
and U114 (N_114,In_132,In_309);
and U115 (N_115,In_489,In_432);
nand U116 (N_116,In_413,In_55);
and U117 (N_117,In_340,In_185);
or U118 (N_118,In_347,In_96);
nor U119 (N_119,In_245,In_265);
and U120 (N_120,N_118,In_304);
and U121 (N_121,In_212,In_382);
nand U122 (N_122,In_274,In_289);
and U123 (N_123,In_110,N_106);
or U124 (N_124,In_155,In_452);
or U125 (N_125,In_236,N_12);
xor U126 (N_126,N_105,In_486);
nand U127 (N_127,N_99,In_2);
nand U128 (N_128,N_25,In_195);
nand U129 (N_129,N_3,In_448);
or U130 (N_130,In_56,In_146);
and U131 (N_131,In_418,In_33);
nor U132 (N_132,N_21,N_77);
and U133 (N_133,In_483,In_38);
nand U134 (N_134,N_116,N_119);
and U135 (N_135,In_13,In_499);
and U136 (N_136,N_16,N_27);
or U137 (N_137,In_430,N_45);
nand U138 (N_138,N_72,In_254);
and U139 (N_139,In_176,N_39);
or U140 (N_140,N_61,In_47);
nand U141 (N_141,N_96,In_103);
or U142 (N_142,N_6,In_286);
or U143 (N_143,In_262,In_492);
nor U144 (N_144,N_103,In_302);
or U145 (N_145,In_385,In_400);
nand U146 (N_146,In_37,In_459);
nor U147 (N_147,In_296,In_109);
and U148 (N_148,In_321,In_143);
nand U149 (N_149,N_117,In_87);
or U150 (N_150,In_124,In_113);
or U151 (N_151,N_30,In_389);
nor U152 (N_152,N_97,N_68);
xnor U153 (N_153,In_1,N_79);
nand U154 (N_154,In_415,In_288);
nand U155 (N_155,N_7,In_490);
nor U156 (N_156,In_224,In_468);
or U157 (N_157,N_113,In_76);
nand U158 (N_158,N_92,N_51);
and U159 (N_159,In_456,In_361);
or U160 (N_160,In_64,In_394);
nand U161 (N_161,In_450,In_357);
and U162 (N_162,In_34,N_63);
or U163 (N_163,N_33,In_270);
or U164 (N_164,N_83,In_420);
or U165 (N_165,In_277,In_114);
or U166 (N_166,In_181,In_97);
nand U167 (N_167,In_476,In_26);
and U168 (N_168,In_417,In_100);
nand U169 (N_169,In_331,N_2);
and U170 (N_170,In_441,In_479);
xor U171 (N_171,In_40,In_220);
nor U172 (N_172,N_115,In_328);
and U173 (N_173,N_95,N_38);
nand U174 (N_174,In_180,In_453);
and U175 (N_175,N_71,N_94);
nand U176 (N_176,In_88,In_449);
nand U177 (N_177,N_22,In_256);
nand U178 (N_178,N_4,In_358);
or U179 (N_179,In_310,N_59);
and U180 (N_180,In_364,In_186);
nand U181 (N_181,In_19,In_211);
and U182 (N_182,In_42,In_493);
or U183 (N_183,N_114,N_84);
or U184 (N_184,In_117,N_58);
or U185 (N_185,In_470,N_74);
nand U186 (N_186,N_160,In_327);
nor U187 (N_187,In_90,N_18);
or U188 (N_188,In_370,In_406);
and U189 (N_189,In_387,In_95);
or U190 (N_190,In_242,In_249);
nor U191 (N_191,In_118,In_226);
and U192 (N_192,N_131,In_206);
nor U193 (N_193,In_330,In_21);
nand U194 (N_194,In_380,In_301);
and U195 (N_195,In_157,In_184);
nor U196 (N_196,In_352,In_315);
nor U197 (N_197,N_133,In_384);
nand U198 (N_198,In_136,In_105);
nor U199 (N_199,N_149,N_32);
nor U200 (N_200,In_174,In_231);
nor U201 (N_201,N_132,N_124);
nor U202 (N_202,In_12,In_74);
or U203 (N_203,N_57,N_148);
and U204 (N_204,N_80,In_16);
or U205 (N_205,N_67,N_47);
and U206 (N_206,In_78,In_381);
nand U207 (N_207,In_41,N_128);
xnor U208 (N_208,In_168,N_136);
and U209 (N_209,In_356,In_31);
or U210 (N_210,In_423,N_111);
nand U211 (N_211,In_446,In_50);
nand U212 (N_212,In_72,N_100);
or U213 (N_213,N_120,In_365);
or U214 (N_214,N_122,In_45);
and U215 (N_215,In_458,N_166);
nand U216 (N_216,In_234,N_171);
or U217 (N_217,In_166,N_112);
xnor U218 (N_218,In_278,In_255);
nor U219 (N_219,In_57,N_42);
nor U220 (N_220,In_60,In_15);
or U221 (N_221,In_173,In_318);
nand U222 (N_222,In_266,N_48);
or U223 (N_223,In_107,N_140);
nor U224 (N_224,In_218,In_297);
or U225 (N_225,In_326,In_438);
nand U226 (N_226,N_162,In_299);
nand U227 (N_227,N_134,In_175);
nor U228 (N_228,In_292,In_112);
xnor U229 (N_229,In_81,In_190);
nor U230 (N_230,N_179,N_64);
nand U231 (N_231,In_461,In_322);
nor U232 (N_232,In_261,N_121);
xnor U233 (N_233,In_410,N_62);
or U234 (N_234,N_138,N_35);
xor U235 (N_235,N_129,In_191);
nor U236 (N_236,In_91,N_29);
and U237 (N_237,N_170,In_335);
and U238 (N_238,N_70,In_421);
nand U239 (N_239,N_127,In_165);
nor U240 (N_240,N_146,N_223);
and U241 (N_241,In_75,N_222);
nand U242 (N_242,In_244,N_161);
nor U243 (N_243,In_230,In_198);
and U244 (N_244,N_139,N_8);
nor U245 (N_245,In_241,N_190);
and U246 (N_246,N_191,In_135);
xor U247 (N_247,In_457,N_209);
and U248 (N_248,In_116,In_151);
nand U249 (N_249,N_125,In_39);
and U250 (N_250,In_122,In_283);
nand U251 (N_251,N_37,N_234);
and U252 (N_252,In_307,N_182);
and U253 (N_253,In_337,N_193);
and U254 (N_254,In_3,In_130);
and U255 (N_255,N_225,In_484);
nand U256 (N_256,In_98,N_205);
nand U257 (N_257,N_204,In_247);
nand U258 (N_258,In_101,In_498);
nand U259 (N_259,N_232,In_10);
or U260 (N_260,N_152,In_339);
or U261 (N_261,N_93,In_391);
xnor U262 (N_262,N_20,In_102);
nor U263 (N_263,In_464,N_229);
and U264 (N_264,N_88,In_62);
or U265 (N_265,N_230,In_320);
or U266 (N_266,In_65,In_325);
and U267 (N_267,In_202,N_206);
xor U268 (N_268,In_443,N_173);
nor U269 (N_269,N_10,N_216);
and U270 (N_270,In_275,N_224);
nor U271 (N_271,N_208,N_195);
nor U272 (N_272,N_239,N_215);
nand U273 (N_273,In_196,N_156);
and U274 (N_274,In_93,N_157);
xnor U275 (N_275,In_285,In_150);
nor U276 (N_276,In_316,N_167);
nor U277 (N_277,In_290,N_189);
or U278 (N_278,N_181,In_209);
or U279 (N_279,In_333,In_214);
nand U280 (N_280,In_70,N_187);
nand U281 (N_281,N_90,N_228);
nand U282 (N_282,N_227,N_185);
or U283 (N_283,In_119,In_444);
nor U284 (N_284,In_466,In_79);
xnor U285 (N_285,In_182,N_213);
or U286 (N_286,In_411,N_143);
xnor U287 (N_287,In_407,N_89);
or U288 (N_288,N_26,In_383);
or U289 (N_289,N_17,In_148);
nor U290 (N_290,N_85,In_477);
and U291 (N_291,In_373,N_210);
nand U292 (N_292,In_167,N_65);
nand U293 (N_293,N_186,N_145);
and U294 (N_294,N_212,N_75);
and U295 (N_295,N_34,N_177);
nor U296 (N_296,In_27,In_281);
and U297 (N_297,N_28,N_98);
or U298 (N_298,N_60,In_467);
and U299 (N_299,N_126,N_192);
nand U300 (N_300,N_284,N_169);
and U301 (N_301,N_293,In_59);
and U302 (N_302,In_237,N_249);
or U303 (N_303,N_295,In_221);
xor U304 (N_304,N_1,In_49);
nand U305 (N_305,N_87,In_401);
nor U306 (N_306,N_123,N_231);
and U307 (N_307,N_130,N_196);
xnor U308 (N_308,In_346,N_141);
xor U309 (N_309,In_362,N_144);
nor U310 (N_310,N_247,N_242);
and U311 (N_311,In_216,N_275);
or U312 (N_312,N_164,In_367);
and U313 (N_313,N_110,In_366);
or U314 (N_314,N_236,In_82);
nand U315 (N_315,N_194,N_252);
and U316 (N_316,N_266,In_53);
and U317 (N_317,N_261,N_76);
and U318 (N_318,In_442,In_147);
or U319 (N_319,N_286,In_474);
and U320 (N_320,In_252,In_253);
and U321 (N_321,In_273,In_193);
or U322 (N_322,In_416,In_386);
nor U323 (N_323,In_141,N_176);
nor U324 (N_324,In_48,In_128);
and U325 (N_325,N_86,N_220);
or U326 (N_326,N_262,N_135);
and U327 (N_327,In_487,N_292);
nor U328 (N_328,In_398,N_282);
and U329 (N_329,N_277,N_200);
xor U330 (N_330,In_6,N_298);
and U331 (N_331,In_465,N_168);
nor U332 (N_332,N_276,N_278);
and U333 (N_333,In_409,N_155);
or U334 (N_334,In_354,N_287);
xor U335 (N_335,N_108,N_279);
nor U336 (N_336,In_259,N_73);
nand U337 (N_337,N_244,N_203);
xnor U338 (N_338,In_329,N_259);
nand U339 (N_339,In_478,N_251);
or U340 (N_340,N_246,In_188);
and U341 (N_341,N_271,N_24);
nor U342 (N_342,N_264,N_294);
or U343 (N_343,N_233,N_165);
or U344 (N_344,N_268,N_285);
and U345 (N_345,N_40,N_5);
nand U346 (N_346,N_214,In_294);
nor U347 (N_347,N_260,N_66);
nor U348 (N_348,N_270,N_291);
or U349 (N_349,In_308,N_297);
and U350 (N_350,N_243,N_273);
or U351 (N_351,N_54,N_202);
nor U352 (N_352,N_107,N_221);
nand U353 (N_353,N_255,N_218);
nor U354 (N_354,N_254,N_248);
nand U355 (N_355,N_263,N_153);
nor U356 (N_356,In_84,In_240);
and U357 (N_357,N_250,N_211);
nand U358 (N_358,N_137,N_283);
nor U359 (N_359,N_235,In_298);
or U360 (N_360,N_304,N_241);
nor U361 (N_361,N_350,In_264);
nor U362 (N_362,N_356,In_344);
and U363 (N_363,N_109,N_150);
nor U364 (N_364,N_180,N_328);
nor U365 (N_365,N_272,N_318);
nand U366 (N_366,N_82,N_310);
nor U367 (N_367,N_353,In_54);
xnor U368 (N_368,N_269,N_330);
xnor U369 (N_369,N_154,N_102);
nor U370 (N_370,In_369,N_296);
or U371 (N_371,N_207,N_309);
or U372 (N_372,In_69,N_151);
nor U373 (N_373,N_336,In_77);
nor U374 (N_374,N_352,N_312);
and U375 (N_375,N_338,N_81);
nand U376 (N_376,N_78,N_327);
nand U377 (N_377,In_276,In_43);
nor U378 (N_378,N_323,N_69);
nor U379 (N_379,N_349,N_359);
or U380 (N_380,N_326,N_238);
or U381 (N_381,N_147,N_253);
nand U382 (N_382,N_307,N_142);
nand U383 (N_383,N_217,N_340);
or U384 (N_384,In_71,In_35);
nand U385 (N_385,N_301,N_300);
nor U386 (N_386,N_281,N_315);
or U387 (N_387,N_348,N_290);
and U388 (N_388,N_329,N_197);
nor U389 (N_389,N_267,N_101);
nand U390 (N_390,N_354,In_73);
or U391 (N_391,N_178,N_303);
nor U392 (N_392,In_85,N_219);
nor U393 (N_393,N_104,N_357);
nor U394 (N_394,N_226,N_308);
nor U395 (N_395,N_322,In_447);
or U396 (N_396,N_302,In_475);
or U397 (N_397,N_332,N_274);
and U398 (N_398,N_347,N_237);
xnor U399 (N_399,In_23,N_158);
nand U400 (N_400,N_240,N_341);
nand U401 (N_401,In_295,N_199);
nand U402 (N_402,N_9,N_245);
and U403 (N_403,N_345,N_351);
and U404 (N_404,In_207,N_333);
or U405 (N_405,N_288,N_314);
nor U406 (N_406,N_339,N_289);
and U407 (N_407,In_390,N_334);
nor U408 (N_408,N_305,N_342);
or U409 (N_409,N_265,N_320);
xor U410 (N_410,N_355,N_319);
nor U411 (N_411,N_325,N_163);
nand U412 (N_412,N_257,In_5);
or U413 (N_413,N_280,N_91);
or U414 (N_414,In_20,N_343);
xnor U415 (N_415,N_337,N_299);
or U416 (N_416,N_184,N_198);
nor U417 (N_417,N_256,N_324);
and U418 (N_418,N_344,N_175);
and U419 (N_419,N_346,N_159);
nor U420 (N_420,N_360,N_400);
or U421 (N_421,N_407,N_358);
and U422 (N_422,N_372,N_183);
nor U423 (N_423,N_402,N_394);
nand U424 (N_424,In_345,N_316);
nor U425 (N_425,N_362,N_395);
or U426 (N_426,N_387,N_317);
and U427 (N_427,N_393,N_406);
nand U428 (N_428,N_414,N_365);
and U429 (N_429,N_335,N_408);
nor U430 (N_430,N_398,N_370);
nor U431 (N_431,N_410,N_201);
or U432 (N_432,N_401,N_172);
and U433 (N_433,N_367,N_405);
nor U434 (N_434,N_368,N_419);
nand U435 (N_435,N_369,N_413);
nand U436 (N_436,N_376,N_363);
xnor U437 (N_437,In_359,N_412);
and U438 (N_438,N_409,N_377);
xor U439 (N_439,N_306,N_397);
xnor U440 (N_440,N_371,N_391);
nor U441 (N_441,N_331,N_374);
nor U442 (N_442,N_399,N_382);
nand U443 (N_443,In_8,In_360);
nand U444 (N_444,N_174,N_389);
nor U445 (N_445,N_384,N_390);
xor U446 (N_446,N_385,N_188);
and U447 (N_447,N_383,N_416);
nand U448 (N_448,N_49,N_321);
nor U449 (N_449,N_378,N_364);
nor U450 (N_450,N_411,N_386);
or U451 (N_451,N_380,N_379);
nor U452 (N_452,N_258,N_311);
nand U453 (N_453,N_404,N_392);
xor U454 (N_454,N_373,N_375);
or U455 (N_455,N_403,N_418);
and U456 (N_456,N_417,N_381);
nand U457 (N_457,N_313,N_388);
nand U458 (N_458,N_396,N_366);
nand U459 (N_459,N_415,N_361);
and U460 (N_460,N_367,N_414);
or U461 (N_461,N_401,N_374);
nor U462 (N_462,N_418,N_361);
and U463 (N_463,N_369,N_370);
or U464 (N_464,N_368,N_376);
nand U465 (N_465,N_49,In_8);
nand U466 (N_466,N_413,N_385);
and U467 (N_467,N_396,N_387);
or U468 (N_468,N_394,N_389);
nor U469 (N_469,N_390,N_364);
and U470 (N_470,N_394,N_388);
nor U471 (N_471,N_313,N_401);
and U472 (N_472,N_419,N_367);
nand U473 (N_473,N_368,N_366);
or U474 (N_474,In_345,N_321);
nor U475 (N_475,N_172,N_382);
or U476 (N_476,N_413,N_172);
nand U477 (N_477,N_399,N_258);
nand U478 (N_478,N_188,N_410);
nor U479 (N_479,N_370,N_360);
or U480 (N_480,N_465,N_447);
and U481 (N_481,N_446,N_450);
or U482 (N_482,N_427,N_454);
nand U483 (N_483,N_457,N_438);
nand U484 (N_484,N_440,N_432);
and U485 (N_485,N_470,N_476);
or U486 (N_486,N_472,N_477);
nor U487 (N_487,N_421,N_435);
nor U488 (N_488,N_462,N_431);
or U489 (N_489,N_461,N_455);
nand U490 (N_490,N_430,N_453);
xnor U491 (N_491,N_437,N_425);
or U492 (N_492,N_464,N_467);
nor U493 (N_493,N_433,N_471);
nand U494 (N_494,N_463,N_460);
nand U495 (N_495,N_456,N_459);
and U496 (N_496,N_452,N_449);
or U497 (N_497,N_429,N_443);
or U498 (N_498,N_426,N_478);
and U499 (N_499,N_473,N_466);
and U500 (N_500,N_474,N_458);
nand U501 (N_501,N_441,N_469);
and U502 (N_502,N_422,N_451);
or U503 (N_503,N_424,N_448);
nor U504 (N_504,N_468,N_442);
nand U505 (N_505,N_434,N_445);
or U506 (N_506,N_475,N_428);
and U507 (N_507,N_423,N_439);
xor U508 (N_508,N_479,N_436);
or U509 (N_509,N_420,N_444);
or U510 (N_510,N_439,N_452);
or U511 (N_511,N_426,N_451);
nand U512 (N_512,N_462,N_456);
nand U513 (N_513,N_430,N_473);
and U514 (N_514,N_472,N_429);
or U515 (N_515,N_459,N_463);
xor U516 (N_516,N_463,N_470);
or U517 (N_517,N_442,N_452);
xor U518 (N_518,N_473,N_474);
and U519 (N_519,N_428,N_447);
nor U520 (N_520,N_476,N_473);
or U521 (N_521,N_475,N_460);
and U522 (N_522,N_424,N_450);
nand U523 (N_523,N_423,N_463);
or U524 (N_524,N_429,N_450);
or U525 (N_525,N_449,N_440);
nor U526 (N_526,N_442,N_466);
and U527 (N_527,N_473,N_432);
nand U528 (N_528,N_444,N_465);
nor U529 (N_529,N_462,N_473);
nor U530 (N_530,N_436,N_446);
nand U531 (N_531,N_459,N_428);
or U532 (N_532,N_432,N_427);
nor U533 (N_533,N_450,N_437);
and U534 (N_534,N_450,N_455);
nand U535 (N_535,N_454,N_421);
nor U536 (N_536,N_430,N_432);
nand U537 (N_537,N_443,N_432);
nand U538 (N_538,N_443,N_441);
and U539 (N_539,N_465,N_428);
xor U540 (N_540,N_494,N_486);
xnor U541 (N_541,N_513,N_485);
or U542 (N_542,N_528,N_508);
or U543 (N_543,N_529,N_531);
or U544 (N_544,N_522,N_527);
nand U545 (N_545,N_495,N_532);
or U546 (N_546,N_539,N_481);
or U547 (N_547,N_505,N_517);
and U548 (N_548,N_491,N_483);
or U549 (N_549,N_493,N_534);
nor U550 (N_550,N_502,N_487);
or U551 (N_551,N_500,N_523);
and U552 (N_552,N_538,N_514);
nor U553 (N_553,N_511,N_524);
or U554 (N_554,N_519,N_504);
and U555 (N_555,N_484,N_530);
nor U556 (N_556,N_512,N_537);
and U557 (N_557,N_499,N_501);
xnor U558 (N_558,N_482,N_489);
xnor U559 (N_559,N_492,N_488);
and U560 (N_560,N_521,N_533);
and U561 (N_561,N_507,N_518);
nand U562 (N_562,N_525,N_506);
nand U563 (N_563,N_480,N_510);
and U564 (N_564,N_516,N_526);
nor U565 (N_565,N_498,N_496);
and U566 (N_566,N_515,N_490);
or U567 (N_567,N_497,N_509);
xor U568 (N_568,N_503,N_535);
nand U569 (N_569,N_536,N_520);
nand U570 (N_570,N_526,N_533);
and U571 (N_571,N_495,N_487);
xnor U572 (N_572,N_534,N_488);
nor U573 (N_573,N_537,N_509);
and U574 (N_574,N_510,N_495);
nand U575 (N_575,N_504,N_482);
nand U576 (N_576,N_533,N_484);
xor U577 (N_577,N_522,N_490);
nor U578 (N_578,N_486,N_512);
nand U579 (N_579,N_512,N_511);
nand U580 (N_580,N_516,N_512);
and U581 (N_581,N_495,N_505);
nor U582 (N_582,N_522,N_497);
or U583 (N_583,N_505,N_533);
nor U584 (N_584,N_498,N_495);
and U585 (N_585,N_510,N_538);
nand U586 (N_586,N_503,N_536);
xnor U587 (N_587,N_481,N_509);
xor U588 (N_588,N_519,N_528);
or U589 (N_589,N_484,N_508);
and U590 (N_590,N_481,N_523);
and U591 (N_591,N_531,N_535);
nand U592 (N_592,N_504,N_535);
nor U593 (N_593,N_494,N_508);
xnor U594 (N_594,N_515,N_505);
nand U595 (N_595,N_512,N_498);
nor U596 (N_596,N_538,N_526);
nor U597 (N_597,N_524,N_494);
and U598 (N_598,N_504,N_499);
or U599 (N_599,N_496,N_517);
nor U600 (N_600,N_542,N_555);
nand U601 (N_601,N_574,N_583);
or U602 (N_602,N_598,N_591);
xor U603 (N_603,N_569,N_577);
or U604 (N_604,N_540,N_546);
or U605 (N_605,N_566,N_585);
or U606 (N_606,N_589,N_590);
nor U607 (N_607,N_551,N_573);
nor U608 (N_608,N_541,N_549);
and U609 (N_609,N_584,N_582);
or U610 (N_610,N_544,N_561);
and U611 (N_611,N_568,N_553);
nand U612 (N_612,N_575,N_565);
xnor U613 (N_613,N_563,N_554);
nand U614 (N_614,N_550,N_559);
and U615 (N_615,N_548,N_572);
or U616 (N_616,N_557,N_562);
nand U617 (N_617,N_543,N_547);
or U618 (N_618,N_592,N_597);
nor U619 (N_619,N_593,N_545);
and U620 (N_620,N_571,N_588);
or U621 (N_621,N_587,N_578);
or U622 (N_622,N_596,N_599);
and U623 (N_623,N_594,N_558);
nand U624 (N_624,N_580,N_595);
xor U625 (N_625,N_567,N_570);
nand U626 (N_626,N_586,N_564);
nand U627 (N_627,N_560,N_556);
xnor U628 (N_628,N_579,N_581);
xor U629 (N_629,N_552,N_576);
or U630 (N_630,N_586,N_550);
nor U631 (N_631,N_554,N_598);
or U632 (N_632,N_591,N_548);
or U633 (N_633,N_552,N_584);
and U634 (N_634,N_588,N_548);
and U635 (N_635,N_564,N_572);
nor U636 (N_636,N_567,N_555);
or U637 (N_637,N_592,N_548);
nor U638 (N_638,N_554,N_573);
nor U639 (N_639,N_582,N_568);
and U640 (N_640,N_591,N_562);
nand U641 (N_641,N_595,N_540);
and U642 (N_642,N_546,N_555);
xnor U643 (N_643,N_585,N_577);
nand U644 (N_644,N_563,N_588);
nor U645 (N_645,N_578,N_581);
and U646 (N_646,N_558,N_541);
nor U647 (N_647,N_590,N_554);
or U648 (N_648,N_559,N_564);
or U649 (N_649,N_568,N_562);
nor U650 (N_650,N_591,N_550);
nand U651 (N_651,N_596,N_580);
and U652 (N_652,N_572,N_581);
nor U653 (N_653,N_583,N_551);
and U654 (N_654,N_588,N_542);
nor U655 (N_655,N_575,N_544);
nor U656 (N_656,N_566,N_561);
nor U657 (N_657,N_569,N_553);
nand U658 (N_658,N_543,N_573);
and U659 (N_659,N_546,N_558);
xor U660 (N_660,N_608,N_635);
or U661 (N_661,N_618,N_617);
or U662 (N_662,N_654,N_637);
nor U663 (N_663,N_603,N_613);
or U664 (N_664,N_610,N_657);
xor U665 (N_665,N_646,N_607);
nor U666 (N_666,N_655,N_642);
nand U667 (N_667,N_652,N_606);
xor U668 (N_668,N_653,N_658);
nand U669 (N_669,N_624,N_611);
and U670 (N_670,N_612,N_649);
or U671 (N_671,N_604,N_621);
nor U672 (N_672,N_629,N_647);
and U673 (N_673,N_639,N_631);
nor U674 (N_674,N_616,N_638);
or U675 (N_675,N_645,N_626);
nor U676 (N_676,N_628,N_601);
or U677 (N_677,N_625,N_622);
and U678 (N_678,N_632,N_651);
and U679 (N_679,N_627,N_650);
and U680 (N_680,N_656,N_605);
nand U681 (N_681,N_615,N_640);
nand U682 (N_682,N_641,N_644);
or U683 (N_683,N_623,N_609);
or U684 (N_684,N_643,N_659);
xnor U685 (N_685,N_600,N_619);
and U686 (N_686,N_630,N_648);
nand U687 (N_687,N_602,N_633);
or U688 (N_688,N_636,N_634);
nor U689 (N_689,N_614,N_620);
and U690 (N_690,N_654,N_650);
nand U691 (N_691,N_652,N_630);
and U692 (N_692,N_613,N_608);
nor U693 (N_693,N_652,N_620);
nand U694 (N_694,N_637,N_650);
and U695 (N_695,N_640,N_611);
nand U696 (N_696,N_640,N_655);
nand U697 (N_697,N_654,N_659);
or U698 (N_698,N_628,N_631);
and U699 (N_699,N_609,N_625);
nand U700 (N_700,N_602,N_628);
and U701 (N_701,N_617,N_641);
nor U702 (N_702,N_602,N_619);
nand U703 (N_703,N_618,N_636);
nand U704 (N_704,N_658,N_606);
and U705 (N_705,N_615,N_605);
nand U706 (N_706,N_639,N_656);
or U707 (N_707,N_632,N_649);
and U708 (N_708,N_614,N_640);
and U709 (N_709,N_659,N_627);
nand U710 (N_710,N_650,N_624);
and U711 (N_711,N_636,N_646);
and U712 (N_712,N_637,N_625);
and U713 (N_713,N_608,N_659);
nand U714 (N_714,N_642,N_624);
and U715 (N_715,N_614,N_630);
or U716 (N_716,N_608,N_634);
and U717 (N_717,N_627,N_644);
nand U718 (N_718,N_621,N_657);
and U719 (N_719,N_614,N_642);
or U720 (N_720,N_705,N_668);
or U721 (N_721,N_680,N_664);
or U722 (N_722,N_715,N_696);
or U723 (N_723,N_682,N_671);
or U724 (N_724,N_694,N_695);
and U725 (N_725,N_676,N_661);
and U726 (N_726,N_688,N_708);
and U727 (N_727,N_683,N_717);
nor U728 (N_728,N_686,N_697);
nand U729 (N_729,N_674,N_678);
and U730 (N_730,N_707,N_700);
xor U731 (N_731,N_663,N_690);
and U732 (N_732,N_687,N_679);
nor U733 (N_733,N_689,N_672);
and U734 (N_734,N_692,N_703);
or U735 (N_735,N_716,N_677);
nand U736 (N_736,N_667,N_699);
xor U737 (N_737,N_719,N_704);
nor U738 (N_738,N_662,N_712);
and U739 (N_739,N_718,N_710);
nand U740 (N_740,N_684,N_711);
or U741 (N_741,N_698,N_681);
nand U742 (N_742,N_714,N_665);
or U743 (N_743,N_675,N_691);
and U744 (N_744,N_666,N_673);
nand U745 (N_745,N_701,N_669);
and U746 (N_746,N_702,N_709);
nor U747 (N_747,N_706,N_693);
nor U748 (N_748,N_685,N_670);
or U749 (N_749,N_660,N_713);
xor U750 (N_750,N_687,N_717);
nand U751 (N_751,N_714,N_670);
or U752 (N_752,N_669,N_685);
or U753 (N_753,N_668,N_682);
xor U754 (N_754,N_694,N_708);
nor U755 (N_755,N_693,N_715);
nor U756 (N_756,N_716,N_667);
and U757 (N_757,N_668,N_712);
nor U758 (N_758,N_694,N_701);
nor U759 (N_759,N_663,N_677);
or U760 (N_760,N_688,N_683);
or U761 (N_761,N_669,N_693);
nand U762 (N_762,N_676,N_669);
or U763 (N_763,N_697,N_705);
xnor U764 (N_764,N_703,N_693);
nor U765 (N_765,N_686,N_678);
and U766 (N_766,N_687,N_670);
xor U767 (N_767,N_709,N_696);
nand U768 (N_768,N_679,N_702);
nor U769 (N_769,N_692,N_700);
nor U770 (N_770,N_679,N_664);
xnor U771 (N_771,N_679,N_706);
or U772 (N_772,N_679,N_709);
nand U773 (N_773,N_672,N_703);
and U774 (N_774,N_661,N_700);
xnor U775 (N_775,N_695,N_677);
and U776 (N_776,N_669,N_698);
nand U777 (N_777,N_673,N_719);
nor U778 (N_778,N_717,N_667);
or U779 (N_779,N_672,N_679);
nand U780 (N_780,N_744,N_743);
nor U781 (N_781,N_765,N_733);
xor U782 (N_782,N_732,N_769);
or U783 (N_783,N_764,N_729);
and U784 (N_784,N_754,N_726);
and U785 (N_785,N_761,N_755);
nand U786 (N_786,N_770,N_735);
and U787 (N_787,N_753,N_772);
xnor U788 (N_788,N_759,N_763);
nand U789 (N_789,N_760,N_767);
xnor U790 (N_790,N_775,N_741);
and U791 (N_791,N_748,N_725);
xor U792 (N_792,N_762,N_751);
nand U793 (N_793,N_720,N_771);
nand U794 (N_794,N_777,N_723);
and U795 (N_795,N_758,N_728);
or U796 (N_796,N_742,N_737);
or U797 (N_797,N_745,N_749);
and U798 (N_798,N_739,N_731);
nand U799 (N_799,N_757,N_746);
or U800 (N_800,N_747,N_774);
nor U801 (N_801,N_734,N_740);
and U802 (N_802,N_722,N_727);
nor U803 (N_803,N_776,N_730);
nand U804 (N_804,N_721,N_738);
or U805 (N_805,N_750,N_779);
or U806 (N_806,N_768,N_752);
and U807 (N_807,N_724,N_773);
and U808 (N_808,N_736,N_766);
nor U809 (N_809,N_778,N_756);
or U810 (N_810,N_764,N_754);
or U811 (N_811,N_744,N_739);
nand U812 (N_812,N_768,N_724);
nor U813 (N_813,N_765,N_773);
nand U814 (N_814,N_724,N_774);
and U815 (N_815,N_737,N_753);
or U816 (N_816,N_764,N_751);
or U817 (N_817,N_761,N_769);
or U818 (N_818,N_742,N_770);
nand U819 (N_819,N_726,N_765);
nor U820 (N_820,N_727,N_724);
nor U821 (N_821,N_762,N_756);
and U822 (N_822,N_756,N_738);
or U823 (N_823,N_736,N_769);
or U824 (N_824,N_774,N_778);
nand U825 (N_825,N_734,N_775);
or U826 (N_826,N_744,N_760);
or U827 (N_827,N_729,N_722);
and U828 (N_828,N_744,N_779);
nand U829 (N_829,N_740,N_753);
xnor U830 (N_830,N_743,N_720);
nand U831 (N_831,N_755,N_724);
xnor U832 (N_832,N_748,N_731);
nand U833 (N_833,N_768,N_758);
and U834 (N_834,N_728,N_768);
and U835 (N_835,N_746,N_745);
or U836 (N_836,N_772,N_743);
and U837 (N_837,N_720,N_751);
and U838 (N_838,N_721,N_773);
or U839 (N_839,N_720,N_772);
xor U840 (N_840,N_799,N_793);
and U841 (N_841,N_809,N_789);
or U842 (N_842,N_786,N_780);
or U843 (N_843,N_790,N_800);
nor U844 (N_844,N_781,N_823);
xor U845 (N_845,N_819,N_804);
nand U846 (N_846,N_838,N_837);
or U847 (N_847,N_826,N_782);
nand U848 (N_848,N_792,N_808);
or U849 (N_849,N_834,N_810);
nor U850 (N_850,N_836,N_794);
nand U851 (N_851,N_813,N_820);
and U852 (N_852,N_821,N_822);
nand U853 (N_853,N_797,N_788);
and U854 (N_854,N_832,N_830);
and U855 (N_855,N_796,N_807);
nor U856 (N_856,N_783,N_828);
and U857 (N_857,N_806,N_833);
and U858 (N_858,N_816,N_812);
or U859 (N_859,N_825,N_805);
xnor U860 (N_860,N_815,N_839);
nand U861 (N_861,N_787,N_829);
nand U862 (N_862,N_801,N_817);
and U863 (N_863,N_814,N_784);
nand U864 (N_864,N_818,N_824);
nor U865 (N_865,N_802,N_791);
or U866 (N_866,N_831,N_827);
or U867 (N_867,N_798,N_811);
xnor U868 (N_868,N_785,N_795);
nand U869 (N_869,N_803,N_835);
nand U870 (N_870,N_831,N_820);
xnor U871 (N_871,N_825,N_816);
and U872 (N_872,N_803,N_806);
nor U873 (N_873,N_834,N_793);
and U874 (N_874,N_780,N_793);
or U875 (N_875,N_781,N_793);
nand U876 (N_876,N_811,N_807);
nand U877 (N_877,N_818,N_834);
or U878 (N_878,N_784,N_805);
nand U879 (N_879,N_826,N_780);
nand U880 (N_880,N_828,N_799);
nand U881 (N_881,N_790,N_819);
nand U882 (N_882,N_825,N_792);
and U883 (N_883,N_792,N_818);
and U884 (N_884,N_809,N_784);
or U885 (N_885,N_800,N_836);
and U886 (N_886,N_800,N_785);
nand U887 (N_887,N_825,N_826);
nand U888 (N_888,N_798,N_782);
and U889 (N_889,N_810,N_808);
or U890 (N_890,N_802,N_817);
nand U891 (N_891,N_838,N_812);
and U892 (N_892,N_819,N_800);
and U893 (N_893,N_839,N_819);
or U894 (N_894,N_783,N_794);
and U895 (N_895,N_825,N_798);
or U896 (N_896,N_828,N_833);
and U897 (N_897,N_809,N_798);
and U898 (N_898,N_786,N_784);
and U899 (N_899,N_818,N_806);
nand U900 (N_900,N_851,N_894);
nor U901 (N_901,N_846,N_858);
or U902 (N_902,N_860,N_886);
and U903 (N_903,N_892,N_888);
or U904 (N_904,N_879,N_893);
xor U905 (N_905,N_859,N_869);
nand U906 (N_906,N_874,N_863);
or U907 (N_907,N_882,N_862);
nor U908 (N_908,N_897,N_889);
nand U909 (N_909,N_857,N_855);
or U910 (N_910,N_865,N_895);
nand U911 (N_911,N_847,N_852);
and U912 (N_912,N_871,N_866);
or U913 (N_913,N_878,N_880);
or U914 (N_914,N_842,N_884);
and U915 (N_915,N_864,N_890);
or U916 (N_916,N_841,N_845);
and U917 (N_917,N_898,N_853);
or U918 (N_918,N_868,N_875);
xor U919 (N_919,N_843,N_899);
nor U920 (N_920,N_840,N_872);
nand U921 (N_921,N_854,N_881);
or U922 (N_922,N_873,N_849);
or U923 (N_923,N_891,N_844);
xnor U924 (N_924,N_885,N_883);
nor U925 (N_925,N_867,N_877);
and U926 (N_926,N_876,N_870);
nand U927 (N_927,N_850,N_856);
nor U928 (N_928,N_848,N_896);
or U929 (N_929,N_861,N_887);
nand U930 (N_930,N_873,N_886);
xnor U931 (N_931,N_891,N_876);
nand U932 (N_932,N_880,N_873);
and U933 (N_933,N_845,N_854);
or U934 (N_934,N_845,N_875);
nand U935 (N_935,N_875,N_847);
nand U936 (N_936,N_843,N_892);
nor U937 (N_937,N_856,N_852);
xnor U938 (N_938,N_851,N_853);
nand U939 (N_939,N_882,N_841);
nand U940 (N_940,N_888,N_857);
nor U941 (N_941,N_872,N_891);
and U942 (N_942,N_880,N_898);
or U943 (N_943,N_873,N_860);
nand U944 (N_944,N_887,N_882);
nand U945 (N_945,N_846,N_885);
xor U946 (N_946,N_854,N_886);
and U947 (N_947,N_855,N_871);
nand U948 (N_948,N_867,N_843);
nor U949 (N_949,N_898,N_864);
nor U950 (N_950,N_872,N_858);
nand U951 (N_951,N_869,N_861);
and U952 (N_952,N_857,N_841);
nor U953 (N_953,N_877,N_871);
and U954 (N_954,N_869,N_885);
or U955 (N_955,N_841,N_868);
or U956 (N_956,N_878,N_864);
nor U957 (N_957,N_851,N_859);
and U958 (N_958,N_871,N_842);
or U959 (N_959,N_890,N_858);
and U960 (N_960,N_932,N_902);
nand U961 (N_961,N_944,N_908);
xor U962 (N_962,N_946,N_917);
and U963 (N_963,N_927,N_950);
and U964 (N_964,N_913,N_910);
nor U965 (N_965,N_907,N_916);
nor U966 (N_966,N_935,N_912);
nor U967 (N_967,N_911,N_952);
or U968 (N_968,N_905,N_928);
or U969 (N_969,N_936,N_930);
or U970 (N_970,N_933,N_958);
xor U971 (N_971,N_914,N_918);
nor U972 (N_972,N_906,N_922);
nand U973 (N_973,N_925,N_909);
and U974 (N_974,N_941,N_903);
or U975 (N_975,N_943,N_901);
or U976 (N_976,N_937,N_926);
xnor U977 (N_977,N_956,N_924);
and U978 (N_978,N_954,N_929);
nor U979 (N_979,N_919,N_949);
and U980 (N_980,N_951,N_953);
or U981 (N_981,N_942,N_938);
or U982 (N_982,N_904,N_915);
and U983 (N_983,N_947,N_940);
or U984 (N_984,N_945,N_957);
nand U985 (N_985,N_948,N_931);
nand U986 (N_986,N_939,N_959);
nor U987 (N_987,N_921,N_900);
and U988 (N_988,N_920,N_923);
or U989 (N_989,N_955,N_934);
xnor U990 (N_990,N_948,N_923);
nand U991 (N_991,N_945,N_941);
and U992 (N_992,N_946,N_958);
and U993 (N_993,N_904,N_930);
nand U994 (N_994,N_940,N_918);
or U995 (N_995,N_910,N_932);
nand U996 (N_996,N_933,N_952);
and U997 (N_997,N_951,N_923);
nor U998 (N_998,N_929,N_913);
nand U999 (N_999,N_957,N_905);
nor U1000 (N_1000,N_959,N_914);
and U1001 (N_1001,N_939,N_936);
nor U1002 (N_1002,N_953,N_935);
or U1003 (N_1003,N_951,N_930);
and U1004 (N_1004,N_944,N_926);
nor U1005 (N_1005,N_927,N_931);
and U1006 (N_1006,N_917,N_951);
nor U1007 (N_1007,N_903,N_907);
nand U1008 (N_1008,N_918,N_915);
nor U1009 (N_1009,N_939,N_913);
nand U1010 (N_1010,N_945,N_958);
nor U1011 (N_1011,N_932,N_913);
or U1012 (N_1012,N_933,N_932);
nand U1013 (N_1013,N_930,N_901);
and U1014 (N_1014,N_942,N_901);
xor U1015 (N_1015,N_918,N_909);
and U1016 (N_1016,N_950,N_959);
or U1017 (N_1017,N_907,N_909);
nor U1018 (N_1018,N_902,N_940);
or U1019 (N_1019,N_948,N_935);
nand U1020 (N_1020,N_998,N_990);
or U1021 (N_1021,N_1005,N_974);
nand U1022 (N_1022,N_972,N_1002);
and U1023 (N_1023,N_1000,N_1008);
and U1024 (N_1024,N_986,N_984);
or U1025 (N_1025,N_979,N_996);
or U1026 (N_1026,N_1013,N_1009);
and U1027 (N_1027,N_1015,N_983);
xnor U1028 (N_1028,N_993,N_1016);
and U1029 (N_1029,N_1001,N_995);
nor U1030 (N_1030,N_1019,N_976);
or U1031 (N_1031,N_977,N_1010);
nor U1032 (N_1032,N_971,N_1014);
nand U1033 (N_1033,N_980,N_1006);
nor U1034 (N_1034,N_988,N_962);
nand U1035 (N_1035,N_992,N_1012);
xnor U1036 (N_1036,N_1018,N_997);
and U1037 (N_1037,N_978,N_987);
or U1038 (N_1038,N_966,N_1011);
nand U1039 (N_1039,N_1017,N_965);
nand U1040 (N_1040,N_967,N_975);
nor U1041 (N_1041,N_994,N_981);
or U1042 (N_1042,N_968,N_991);
or U1043 (N_1043,N_970,N_964);
xnor U1044 (N_1044,N_960,N_985);
nor U1045 (N_1045,N_982,N_989);
and U1046 (N_1046,N_1003,N_1004);
nand U1047 (N_1047,N_963,N_969);
or U1048 (N_1048,N_1007,N_973);
nor U1049 (N_1049,N_961,N_999);
nor U1050 (N_1050,N_984,N_981);
or U1051 (N_1051,N_1007,N_968);
or U1052 (N_1052,N_977,N_979);
nor U1053 (N_1053,N_962,N_968);
nand U1054 (N_1054,N_998,N_965);
and U1055 (N_1055,N_1008,N_990);
or U1056 (N_1056,N_1002,N_969);
or U1057 (N_1057,N_971,N_985);
nor U1058 (N_1058,N_1014,N_963);
xor U1059 (N_1059,N_1010,N_1001);
and U1060 (N_1060,N_1008,N_1006);
nor U1061 (N_1061,N_976,N_989);
and U1062 (N_1062,N_960,N_975);
nor U1063 (N_1063,N_988,N_986);
or U1064 (N_1064,N_973,N_963);
nand U1065 (N_1065,N_989,N_997);
and U1066 (N_1066,N_963,N_1012);
nor U1067 (N_1067,N_969,N_1008);
nor U1068 (N_1068,N_981,N_979);
nor U1069 (N_1069,N_985,N_986);
xor U1070 (N_1070,N_964,N_987);
or U1071 (N_1071,N_1010,N_982);
nand U1072 (N_1072,N_993,N_1004);
or U1073 (N_1073,N_992,N_1001);
or U1074 (N_1074,N_967,N_993);
nand U1075 (N_1075,N_976,N_1002);
and U1076 (N_1076,N_1014,N_1001);
nand U1077 (N_1077,N_1015,N_963);
or U1078 (N_1078,N_988,N_991);
and U1079 (N_1079,N_979,N_1017);
or U1080 (N_1080,N_1048,N_1045);
and U1081 (N_1081,N_1054,N_1038);
or U1082 (N_1082,N_1057,N_1075);
or U1083 (N_1083,N_1050,N_1077);
nor U1084 (N_1084,N_1040,N_1034);
nor U1085 (N_1085,N_1036,N_1027);
and U1086 (N_1086,N_1049,N_1079);
nor U1087 (N_1087,N_1047,N_1046);
nor U1088 (N_1088,N_1032,N_1065);
xor U1089 (N_1089,N_1074,N_1066);
and U1090 (N_1090,N_1060,N_1044);
xor U1091 (N_1091,N_1063,N_1069);
nor U1092 (N_1092,N_1062,N_1056);
nand U1093 (N_1093,N_1023,N_1035);
nor U1094 (N_1094,N_1043,N_1055);
or U1095 (N_1095,N_1025,N_1067);
and U1096 (N_1096,N_1033,N_1026);
or U1097 (N_1097,N_1052,N_1076);
nand U1098 (N_1098,N_1061,N_1042);
or U1099 (N_1099,N_1037,N_1020);
xnor U1100 (N_1100,N_1022,N_1072);
nand U1101 (N_1101,N_1051,N_1078);
and U1102 (N_1102,N_1059,N_1029);
and U1103 (N_1103,N_1031,N_1024);
nor U1104 (N_1104,N_1068,N_1058);
or U1105 (N_1105,N_1028,N_1021);
nor U1106 (N_1106,N_1071,N_1073);
and U1107 (N_1107,N_1053,N_1041);
nand U1108 (N_1108,N_1039,N_1070);
and U1109 (N_1109,N_1030,N_1064);
and U1110 (N_1110,N_1051,N_1034);
or U1111 (N_1111,N_1036,N_1069);
or U1112 (N_1112,N_1048,N_1032);
nor U1113 (N_1113,N_1075,N_1026);
xnor U1114 (N_1114,N_1048,N_1064);
nor U1115 (N_1115,N_1045,N_1047);
or U1116 (N_1116,N_1057,N_1040);
nand U1117 (N_1117,N_1044,N_1036);
or U1118 (N_1118,N_1054,N_1074);
or U1119 (N_1119,N_1071,N_1034);
nand U1120 (N_1120,N_1032,N_1068);
nor U1121 (N_1121,N_1059,N_1051);
or U1122 (N_1122,N_1037,N_1045);
or U1123 (N_1123,N_1078,N_1069);
nand U1124 (N_1124,N_1024,N_1067);
nand U1125 (N_1125,N_1030,N_1043);
xor U1126 (N_1126,N_1029,N_1031);
or U1127 (N_1127,N_1022,N_1039);
nor U1128 (N_1128,N_1039,N_1049);
or U1129 (N_1129,N_1051,N_1043);
and U1130 (N_1130,N_1027,N_1062);
nand U1131 (N_1131,N_1029,N_1020);
nand U1132 (N_1132,N_1063,N_1070);
nor U1133 (N_1133,N_1071,N_1078);
and U1134 (N_1134,N_1020,N_1068);
nand U1135 (N_1135,N_1042,N_1070);
nand U1136 (N_1136,N_1021,N_1030);
or U1137 (N_1137,N_1076,N_1059);
or U1138 (N_1138,N_1044,N_1040);
xor U1139 (N_1139,N_1035,N_1067);
nand U1140 (N_1140,N_1081,N_1104);
and U1141 (N_1141,N_1113,N_1135);
or U1142 (N_1142,N_1119,N_1103);
and U1143 (N_1143,N_1111,N_1080);
nor U1144 (N_1144,N_1110,N_1122);
or U1145 (N_1145,N_1116,N_1115);
nand U1146 (N_1146,N_1124,N_1117);
nand U1147 (N_1147,N_1137,N_1127);
xor U1148 (N_1148,N_1107,N_1132);
or U1149 (N_1149,N_1130,N_1126);
and U1150 (N_1150,N_1121,N_1108);
nor U1151 (N_1151,N_1097,N_1085);
or U1152 (N_1152,N_1138,N_1093);
xor U1153 (N_1153,N_1106,N_1090);
or U1154 (N_1154,N_1131,N_1084);
nor U1155 (N_1155,N_1123,N_1088);
or U1156 (N_1156,N_1083,N_1101);
nor U1157 (N_1157,N_1094,N_1105);
nand U1158 (N_1158,N_1099,N_1095);
nand U1159 (N_1159,N_1133,N_1098);
nand U1160 (N_1160,N_1092,N_1087);
nor U1161 (N_1161,N_1129,N_1134);
nor U1162 (N_1162,N_1112,N_1120);
and U1163 (N_1163,N_1096,N_1089);
and U1164 (N_1164,N_1109,N_1136);
nor U1165 (N_1165,N_1100,N_1091);
nand U1166 (N_1166,N_1125,N_1086);
nand U1167 (N_1167,N_1118,N_1102);
and U1168 (N_1168,N_1139,N_1082);
or U1169 (N_1169,N_1114,N_1128);
and U1170 (N_1170,N_1128,N_1080);
nor U1171 (N_1171,N_1132,N_1085);
or U1172 (N_1172,N_1087,N_1109);
or U1173 (N_1173,N_1127,N_1130);
and U1174 (N_1174,N_1094,N_1100);
nand U1175 (N_1175,N_1137,N_1120);
nor U1176 (N_1176,N_1081,N_1114);
or U1177 (N_1177,N_1115,N_1136);
or U1178 (N_1178,N_1123,N_1089);
and U1179 (N_1179,N_1091,N_1114);
nand U1180 (N_1180,N_1083,N_1102);
and U1181 (N_1181,N_1110,N_1130);
nor U1182 (N_1182,N_1138,N_1127);
xnor U1183 (N_1183,N_1138,N_1091);
and U1184 (N_1184,N_1104,N_1113);
nand U1185 (N_1185,N_1131,N_1106);
and U1186 (N_1186,N_1103,N_1123);
nand U1187 (N_1187,N_1125,N_1117);
nand U1188 (N_1188,N_1088,N_1092);
or U1189 (N_1189,N_1135,N_1131);
and U1190 (N_1190,N_1113,N_1103);
or U1191 (N_1191,N_1127,N_1090);
nand U1192 (N_1192,N_1135,N_1098);
nand U1193 (N_1193,N_1129,N_1084);
xor U1194 (N_1194,N_1105,N_1131);
nor U1195 (N_1195,N_1094,N_1113);
nor U1196 (N_1196,N_1085,N_1119);
xor U1197 (N_1197,N_1105,N_1133);
nand U1198 (N_1198,N_1131,N_1128);
or U1199 (N_1199,N_1121,N_1114);
or U1200 (N_1200,N_1147,N_1177);
nand U1201 (N_1201,N_1161,N_1151);
or U1202 (N_1202,N_1144,N_1167);
nand U1203 (N_1203,N_1141,N_1170);
and U1204 (N_1204,N_1186,N_1179);
nand U1205 (N_1205,N_1164,N_1146);
or U1206 (N_1206,N_1158,N_1183);
and U1207 (N_1207,N_1163,N_1182);
nor U1208 (N_1208,N_1140,N_1198);
and U1209 (N_1209,N_1172,N_1153);
nor U1210 (N_1210,N_1142,N_1152);
nor U1211 (N_1211,N_1185,N_1181);
nor U1212 (N_1212,N_1178,N_1184);
nor U1213 (N_1213,N_1168,N_1173);
xor U1214 (N_1214,N_1197,N_1193);
and U1215 (N_1215,N_1191,N_1159);
and U1216 (N_1216,N_1199,N_1192);
or U1217 (N_1217,N_1188,N_1180);
nor U1218 (N_1218,N_1143,N_1149);
nor U1219 (N_1219,N_1165,N_1187);
and U1220 (N_1220,N_1145,N_1194);
nand U1221 (N_1221,N_1155,N_1154);
nor U1222 (N_1222,N_1189,N_1195);
or U1223 (N_1223,N_1175,N_1148);
nor U1224 (N_1224,N_1169,N_1160);
or U1225 (N_1225,N_1162,N_1157);
nor U1226 (N_1226,N_1190,N_1176);
nor U1227 (N_1227,N_1166,N_1150);
and U1228 (N_1228,N_1196,N_1171);
nand U1229 (N_1229,N_1174,N_1156);
nand U1230 (N_1230,N_1158,N_1167);
nor U1231 (N_1231,N_1153,N_1148);
nor U1232 (N_1232,N_1175,N_1181);
nor U1233 (N_1233,N_1168,N_1151);
nor U1234 (N_1234,N_1145,N_1187);
xnor U1235 (N_1235,N_1171,N_1151);
or U1236 (N_1236,N_1163,N_1175);
or U1237 (N_1237,N_1169,N_1140);
nand U1238 (N_1238,N_1194,N_1156);
and U1239 (N_1239,N_1188,N_1153);
or U1240 (N_1240,N_1154,N_1141);
and U1241 (N_1241,N_1179,N_1197);
or U1242 (N_1242,N_1164,N_1180);
nand U1243 (N_1243,N_1157,N_1141);
or U1244 (N_1244,N_1197,N_1148);
or U1245 (N_1245,N_1175,N_1190);
nor U1246 (N_1246,N_1166,N_1165);
nand U1247 (N_1247,N_1183,N_1172);
and U1248 (N_1248,N_1150,N_1141);
nand U1249 (N_1249,N_1186,N_1197);
nand U1250 (N_1250,N_1182,N_1149);
or U1251 (N_1251,N_1192,N_1189);
or U1252 (N_1252,N_1189,N_1185);
or U1253 (N_1253,N_1155,N_1153);
nor U1254 (N_1254,N_1148,N_1176);
nor U1255 (N_1255,N_1142,N_1153);
xor U1256 (N_1256,N_1179,N_1184);
nor U1257 (N_1257,N_1198,N_1170);
or U1258 (N_1258,N_1198,N_1171);
or U1259 (N_1259,N_1173,N_1140);
or U1260 (N_1260,N_1227,N_1246);
and U1261 (N_1261,N_1210,N_1255);
and U1262 (N_1262,N_1248,N_1239);
nor U1263 (N_1263,N_1213,N_1201);
nand U1264 (N_1264,N_1224,N_1230);
nand U1265 (N_1265,N_1214,N_1204);
and U1266 (N_1266,N_1244,N_1247);
or U1267 (N_1267,N_1217,N_1245);
xor U1268 (N_1268,N_1241,N_1205);
or U1269 (N_1269,N_1231,N_1215);
or U1270 (N_1270,N_1218,N_1254);
nand U1271 (N_1271,N_1236,N_1238);
or U1272 (N_1272,N_1259,N_1200);
and U1273 (N_1273,N_1226,N_1233);
or U1274 (N_1274,N_1209,N_1220);
and U1275 (N_1275,N_1207,N_1240);
nand U1276 (N_1276,N_1212,N_1216);
nand U1277 (N_1277,N_1232,N_1203);
and U1278 (N_1278,N_1219,N_1256);
or U1279 (N_1279,N_1237,N_1253);
xnor U1280 (N_1280,N_1223,N_1221);
or U1281 (N_1281,N_1252,N_1242);
nor U1282 (N_1282,N_1251,N_1257);
nand U1283 (N_1283,N_1229,N_1222);
and U1284 (N_1284,N_1235,N_1208);
nor U1285 (N_1285,N_1206,N_1228);
nor U1286 (N_1286,N_1234,N_1225);
or U1287 (N_1287,N_1211,N_1258);
nand U1288 (N_1288,N_1202,N_1249);
and U1289 (N_1289,N_1250,N_1243);
nor U1290 (N_1290,N_1210,N_1248);
or U1291 (N_1291,N_1222,N_1210);
xnor U1292 (N_1292,N_1219,N_1253);
nor U1293 (N_1293,N_1249,N_1239);
and U1294 (N_1294,N_1235,N_1239);
and U1295 (N_1295,N_1219,N_1234);
nand U1296 (N_1296,N_1205,N_1245);
and U1297 (N_1297,N_1210,N_1203);
xor U1298 (N_1298,N_1255,N_1229);
and U1299 (N_1299,N_1251,N_1258);
nor U1300 (N_1300,N_1202,N_1252);
and U1301 (N_1301,N_1257,N_1224);
nor U1302 (N_1302,N_1244,N_1245);
and U1303 (N_1303,N_1215,N_1258);
and U1304 (N_1304,N_1249,N_1207);
or U1305 (N_1305,N_1219,N_1259);
nand U1306 (N_1306,N_1234,N_1212);
or U1307 (N_1307,N_1226,N_1213);
and U1308 (N_1308,N_1210,N_1244);
nor U1309 (N_1309,N_1240,N_1236);
nor U1310 (N_1310,N_1224,N_1219);
or U1311 (N_1311,N_1244,N_1203);
or U1312 (N_1312,N_1223,N_1203);
or U1313 (N_1313,N_1217,N_1226);
or U1314 (N_1314,N_1249,N_1255);
xnor U1315 (N_1315,N_1213,N_1257);
nand U1316 (N_1316,N_1227,N_1233);
or U1317 (N_1317,N_1217,N_1234);
or U1318 (N_1318,N_1238,N_1251);
nor U1319 (N_1319,N_1209,N_1223);
nand U1320 (N_1320,N_1263,N_1265);
or U1321 (N_1321,N_1319,N_1308);
nor U1322 (N_1322,N_1301,N_1289);
nand U1323 (N_1323,N_1281,N_1288);
xor U1324 (N_1324,N_1272,N_1300);
nand U1325 (N_1325,N_1275,N_1271);
or U1326 (N_1326,N_1311,N_1282);
nand U1327 (N_1327,N_1269,N_1273);
nand U1328 (N_1328,N_1266,N_1262);
nor U1329 (N_1329,N_1280,N_1317);
and U1330 (N_1330,N_1314,N_1310);
nand U1331 (N_1331,N_1302,N_1292);
nand U1332 (N_1332,N_1290,N_1284);
and U1333 (N_1333,N_1261,N_1315);
nor U1334 (N_1334,N_1287,N_1295);
nor U1335 (N_1335,N_1276,N_1278);
nand U1336 (N_1336,N_1299,N_1313);
and U1337 (N_1337,N_1316,N_1294);
or U1338 (N_1338,N_1293,N_1260);
nand U1339 (N_1339,N_1277,N_1279);
nand U1340 (N_1340,N_1267,N_1291);
or U1341 (N_1341,N_1303,N_1318);
nand U1342 (N_1342,N_1309,N_1312);
nor U1343 (N_1343,N_1306,N_1297);
nand U1344 (N_1344,N_1270,N_1305);
and U1345 (N_1345,N_1296,N_1268);
and U1346 (N_1346,N_1307,N_1283);
nand U1347 (N_1347,N_1285,N_1286);
or U1348 (N_1348,N_1264,N_1298);
nor U1349 (N_1349,N_1274,N_1304);
nor U1350 (N_1350,N_1286,N_1280);
and U1351 (N_1351,N_1267,N_1294);
nand U1352 (N_1352,N_1268,N_1308);
nor U1353 (N_1353,N_1289,N_1304);
and U1354 (N_1354,N_1317,N_1299);
nor U1355 (N_1355,N_1314,N_1268);
nor U1356 (N_1356,N_1298,N_1294);
nor U1357 (N_1357,N_1285,N_1306);
and U1358 (N_1358,N_1297,N_1260);
and U1359 (N_1359,N_1296,N_1265);
or U1360 (N_1360,N_1305,N_1282);
or U1361 (N_1361,N_1290,N_1274);
nor U1362 (N_1362,N_1261,N_1275);
or U1363 (N_1363,N_1289,N_1270);
and U1364 (N_1364,N_1302,N_1316);
nor U1365 (N_1365,N_1299,N_1307);
nor U1366 (N_1366,N_1262,N_1261);
and U1367 (N_1367,N_1305,N_1290);
nand U1368 (N_1368,N_1296,N_1297);
nand U1369 (N_1369,N_1261,N_1303);
and U1370 (N_1370,N_1273,N_1291);
xnor U1371 (N_1371,N_1292,N_1312);
nor U1372 (N_1372,N_1281,N_1271);
nor U1373 (N_1373,N_1301,N_1311);
and U1374 (N_1374,N_1317,N_1266);
nor U1375 (N_1375,N_1266,N_1290);
nor U1376 (N_1376,N_1315,N_1281);
nor U1377 (N_1377,N_1261,N_1316);
xnor U1378 (N_1378,N_1308,N_1285);
and U1379 (N_1379,N_1279,N_1300);
and U1380 (N_1380,N_1339,N_1370);
nor U1381 (N_1381,N_1360,N_1354);
nand U1382 (N_1382,N_1371,N_1373);
nor U1383 (N_1383,N_1372,N_1351);
nand U1384 (N_1384,N_1336,N_1357);
and U1385 (N_1385,N_1376,N_1347);
nand U1386 (N_1386,N_1374,N_1328);
nor U1387 (N_1387,N_1326,N_1355);
and U1388 (N_1388,N_1329,N_1353);
nand U1389 (N_1389,N_1356,N_1366);
nor U1390 (N_1390,N_1324,N_1332);
nand U1391 (N_1391,N_1358,N_1342);
nand U1392 (N_1392,N_1338,N_1335);
nor U1393 (N_1393,N_1337,N_1341);
and U1394 (N_1394,N_1348,N_1361);
nand U1395 (N_1395,N_1346,N_1344);
nand U1396 (N_1396,N_1379,N_1377);
and U1397 (N_1397,N_1345,N_1343);
xor U1398 (N_1398,N_1325,N_1327);
nor U1399 (N_1399,N_1333,N_1378);
or U1400 (N_1400,N_1331,N_1321);
xnor U1401 (N_1401,N_1368,N_1369);
nand U1402 (N_1402,N_1349,N_1359);
nand U1403 (N_1403,N_1350,N_1323);
nor U1404 (N_1404,N_1375,N_1367);
nand U1405 (N_1405,N_1334,N_1363);
nor U1406 (N_1406,N_1364,N_1340);
nand U1407 (N_1407,N_1320,N_1365);
and U1408 (N_1408,N_1322,N_1352);
or U1409 (N_1409,N_1362,N_1330);
nor U1410 (N_1410,N_1354,N_1353);
and U1411 (N_1411,N_1330,N_1331);
nor U1412 (N_1412,N_1343,N_1340);
nand U1413 (N_1413,N_1370,N_1359);
xor U1414 (N_1414,N_1328,N_1361);
and U1415 (N_1415,N_1361,N_1364);
nand U1416 (N_1416,N_1335,N_1343);
nor U1417 (N_1417,N_1357,N_1351);
xnor U1418 (N_1418,N_1326,N_1349);
and U1419 (N_1419,N_1332,N_1344);
and U1420 (N_1420,N_1377,N_1346);
or U1421 (N_1421,N_1353,N_1367);
or U1422 (N_1422,N_1330,N_1352);
nor U1423 (N_1423,N_1347,N_1323);
nand U1424 (N_1424,N_1362,N_1372);
nand U1425 (N_1425,N_1321,N_1333);
xor U1426 (N_1426,N_1350,N_1331);
nand U1427 (N_1427,N_1348,N_1350);
and U1428 (N_1428,N_1330,N_1333);
and U1429 (N_1429,N_1340,N_1323);
and U1430 (N_1430,N_1364,N_1365);
nor U1431 (N_1431,N_1363,N_1329);
and U1432 (N_1432,N_1370,N_1361);
and U1433 (N_1433,N_1362,N_1338);
or U1434 (N_1434,N_1332,N_1327);
or U1435 (N_1435,N_1329,N_1342);
nor U1436 (N_1436,N_1379,N_1359);
xor U1437 (N_1437,N_1354,N_1336);
nor U1438 (N_1438,N_1376,N_1379);
or U1439 (N_1439,N_1334,N_1371);
and U1440 (N_1440,N_1421,N_1428);
nand U1441 (N_1441,N_1433,N_1425);
xor U1442 (N_1442,N_1435,N_1437);
or U1443 (N_1443,N_1429,N_1394);
or U1444 (N_1444,N_1407,N_1424);
or U1445 (N_1445,N_1410,N_1418);
or U1446 (N_1446,N_1380,N_1420);
and U1447 (N_1447,N_1434,N_1395);
nand U1448 (N_1448,N_1393,N_1427);
or U1449 (N_1449,N_1438,N_1386);
xnor U1450 (N_1450,N_1423,N_1381);
nand U1451 (N_1451,N_1413,N_1432);
and U1452 (N_1452,N_1388,N_1426);
nand U1453 (N_1453,N_1422,N_1389);
or U1454 (N_1454,N_1439,N_1397);
and U1455 (N_1455,N_1401,N_1436);
and U1456 (N_1456,N_1416,N_1404);
nand U1457 (N_1457,N_1399,N_1403);
and U1458 (N_1458,N_1391,N_1387);
nor U1459 (N_1459,N_1390,N_1411);
xnor U1460 (N_1460,N_1384,N_1430);
or U1461 (N_1461,N_1419,N_1400);
nand U1462 (N_1462,N_1405,N_1402);
or U1463 (N_1463,N_1406,N_1408);
or U1464 (N_1464,N_1382,N_1396);
nor U1465 (N_1465,N_1431,N_1414);
nand U1466 (N_1466,N_1385,N_1417);
or U1467 (N_1467,N_1383,N_1392);
xnor U1468 (N_1468,N_1412,N_1415);
nor U1469 (N_1469,N_1409,N_1398);
nand U1470 (N_1470,N_1423,N_1416);
nor U1471 (N_1471,N_1439,N_1420);
nor U1472 (N_1472,N_1408,N_1409);
nor U1473 (N_1473,N_1424,N_1406);
nor U1474 (N_1474,N_1437,N_1415);
nand U1475 (N_1475,N_1382,N_1384);
nand U1476 (N_1476,N_1425,N_1427);
or U1477 (N_1477,N_1422,N_1382);
or U1478 (N_1478,N_1434,N_1415);
nor U1479 (N_1479,N_1403,N_1429);
or U1480 (N_1480,N_1384,N_1435);
nor U1481 (N_1481,N_1413,N_1421);
nand U1482 (N_1482,N_1424,N_1381);
and U1483 (N_1483,N_1407,N_1431);
and U1484 (N_1484,N_1398,N_1388);
or U1485 (N_1485,N_1399,N_1391);
and U1486 (N_1486,N_1434,N_1424);
nor U1487 (N_1487,N_1403,N_1414);
and U1488 (N_1488,N_1419,N_1417);
nand U1489 (N_1489,N_1410,N_1437);
nor U1490 (N_1490,N_1380,N_1395);
xnor U1491 (N_1491,N_1386,N_1433);
nor U1492 (N_1492,N_1423,N_1388);
or U1493 (N_1493,N_1384,N_1424);
nor U1494 (N_1494,N_1435,N_1399);
nand U1495 (N_1495,N_1439,N_1425);
nand U1496 (N_1496,N_1389,N_1388);
or U1497 (N_1497,N_1414,N_1391);
or U1498 (N_1498,N_1406,N_1415);
and U1499 (N_1499,N_1382,N_1416);
xnor U1500 (N_1500,N_1486,N_1490);
nor U1501 (N_1501,N_1458,N_1480);
and U1502 (N_1502,N_1489,N_1454);
xnor U1503 (N_1503,N_1455,N_1444);
or U1504 (N_1504,N_1466,N_1461);
nor U1505 (N_1505,N_1471,N_1484);
xnor U1506 (N_1506,N_1469,N_1482);
nand U1507 (N_1507,N_1445,N_1459);
nand U1508 (N_1508,N_1440,N_1457);
nand U1509 (N_1509,N_1460,N_1448);
or U1510 (N_1510,N_1449,N_1494);
xor U1511 (N_1511,N_1465,N_1452);
and U1512 (N_1512,N_1447,N_1498);
xnor U1513 (N_1513,N_1479,N_1474);
or U1514 (N_1514,N_1481,N_1451);
and U1515 (N_1515,N_1488,N_1487);
nand U1516 (N_1516,N_1473,N_1456);
or U1517 (N_1517,N_1496,N_1495);
nor U1518 (N_1518,N_1442,N_1462);
and U1519 (N_1519,N_1441,N_1464);
and U1520 (N_1520,N_1485,N_1467);
and U1521 (N_1521,N_1497,N_1443);
nor U1522 (N_1522,N_1475,N_1472);
nor U1523 (N_1523,N_1477,N_1493);
nand U1524 (N_1524,N_1470,N_1450);
or U1525 (N_1525,N_1468,N_1446);
nand U1526 (N_1526,N_1483,N_1478);
and U1527 (N_1527,N_1453,N_1492);
xor U1528 (N_1528,N_1476,N_1463);
nor U1529 (N_1529,N_1491,N_1499);
nor U1530 (N_1530,N_1494,N_1475);
or U1531 (N_1531,N_1497,N_1461);
nand U1532 (N_1532,N_1471,N_1442);
nand U1533 (N_1533,N_1479,N_1440);
nor U1534 (N_1534,N_1455,N_1471);
nand U1535 (N_1535,N_1454,N_1459);
nand U1536 (N_1536,N_1459,N_1443);
or U1537 (N_1537,N_1455,N_1462);
and U1538 (N_1538,N_1473,N_1453);
or U1539 (N_1539,N_1460,N_1481);
nor U1540 (N_1540,N_1468,N_1498);
nand U1541 (N_1541,N_1469,N_1441);
or U1542 (N_1542,N_1462,N_1475);
and U1543 (N_1543,N_1497,N_1493);
xor U1544 (N_1544,N_1451,N_1454);
or U1545 (N_1545,N_1462,N_1463);
xnor U1546 (N_1546,N_1478,N_1443);
nand U1547 (N_1547,N_1446,N_1491);
xnor U1548 (N_1548,N_1442,N_1470);
and U1549 (N_1549,N_1491,N_1479);
nand U1550 (N_1550,N_1466,N_1445);
and U1551 (N_1551,N_1460,N_1449);
or U1552 (N_1552,N_1451,N_1496);
nand U1553 (N_1553,N_1479,N_1488);
nor U1554 (N_1554,N_1448,N_1468);
and U1555 (N_1555,N_1465,N_1458);
nand U1556 (N_1556,N_1486,N_1451);
and U1557 (N_1557,N_1495,N_1465);
nor U1558 (N_1558,N_1472,N_1455);
nor U1559 (N_1559,N_1458,N_1497);
nand U1560 (N_1560,N_1554,N_1544);
nor U1561 (N_1561,N_1526,N_1513);
nor U1562 (N_1562,N_1517,N_1551);
and U1563 (N_1563,N_1545,N_1539);
xnor U1564 (N_1564,N_1549,N_1557);
nor U1565 (N_1565,N_1523,N_1558);
and U1566 (N_1566,N_1502,N_1522);
nand U1567 (N_1567,N_1542,N_1503);
nand U1568 (N_1568,N_1536,N_1506);
nand U1569 (N_1569,N_1518,N_1507);
or U1570 (N_1570,N_1528,N_1556);
nand U1571 (N_1571,N_1519,N_1538);
and U1572 (N_1572,N_1541,N_1512);
nor U1573 (N_1573,N_1547,N_1555);
xnor U1574 (N_1574,N_1500,N_1552);
nor U1575 (N_1575,N_1509,N_1505);
nand U1576 (N_1576,N_1527,N_1520);
nor U1577 (N_1577,N_1543,N_1548);
nand U1578 (N_1578,N_1550,N_1532);
nor U1579 (N_1579,N_1537,N_1525);
and U1580 (N_1580,N_1529,N_1535);
nand U1581 (N_1581,N_1514,N_1508);
nor U1582 (N_1582,N_1533,N_1521);
and U1583 (N_1583,N_1511,N_1515);
xnor U1584 (N_1584,N_1530,N_1516);
xor U1585 (N_1585,N_1546,N_1534);
nor U1586 (N_1586,N_1559,N_1531);
or U1587 (N_1587,N_1553,N_1524);
nor U1588 (N_1588,N_1504,N_1501);
and U1589 (N_1589,N_1510,N_1540);
nor U1590 (N_1590,N_1524,N_1505);
nor U1591 (N_1591,N_1547,N_1513);
nand U1592 (N_1592,N_1558,N_1522);
or U1593 (N_1593,N_1503,N_1527);
nand U1594 (N_1594,N_1544,N_1536);
or U1595 (N_1595,N_1529,N_1500);
and U1596 (N_1596,N_1548,N_1505);
and U1597 (N_1597,N_1513,N_1541);
or U1598 (N_1598,N_1527,N_1518);
or U1599 (N_1599,N_1552,N_1505);
nand U1600 (N_1600,N_1531,N_1548);
nor U1601 (N_1601,N_1551,N_1536);
nor U1602 (N_1602,N_1508,N_1557);
or U1603 (N_1603,N_1545,N_1548);
nand U1604 (N_1604,N_1536,N_1524);
and U1605 (N_1605,N_1513,N_1511);
xnor U1606 (N_1606,N_1516,N_1557);
nor U1607 (N_1607,N_1532,N_1531);
and U1608 (N_1608,N_1556,N_1518);
or U1609 (N_1609,N_1537,N_1536);
or U1610 (N_1610,N_1520,N_1523);
nor U1611 (N_1611,N_1554,N_1531);
nor U1612 (N_1612,N_1523,N_1514);
nor U1613 (N_1613,N_1555,N_1545);
nand U1614 (N_1614,N_1556,N_1527);
or U1615 (N_1615,N_1540,N_1501);
nor U1616 (N_1616,N_1536,N_1557);
nor U1617 (N_1617,N_1503,N_1517);
nand U1618 (N_1618,N_1513,N_1535);
nand U1619 (N_1619,N_1500,N_1539);
or U1620 (N_1620,N_1598,N_1575);
nor U1621 (N_1621,N_1589,N_1577);
and U1622 (N_1622,N_1572,N_1586);
or U1623 (N_1623,N_1588,N_1585);
xnor U1624 (N_1624,N_1565,N_1580);
nor U1625 (N_1625,N_1578,N_1560);
nand U1626 (N_1626,N_1596,N_1566);
and U1627 (N_1627,N_1615,N_1617);
nand U1628 (N_1628,N_1576,N_1571);
nor U1629 (N_1629,N_1616,N_1603);
or U1630 (N_1630,N_1600,N_1574);
and U1631 (N_1631,N_1591,N_1602);
or U1632 (N_1632,N_1610,N_1579);
nor U1633 (N_1633,N_1593,N_1581);
xnor U1634 (N_1634,N_1599,N_1607);
nand U1635 (N_1635,N_1570,N_1594);
or U1636 (N_1636,N_1618,N_1613);
xor U1637 (N_1637,N_1601,N_1573);
xor U1638 (N_1638,N_1609,N_1564);
or U1639 (N_1639,N_1563,N_1562);
xor U1640 (N_1640,N_1608,N_1567);
nor U1641 (N_1641,N_1606,N_1614);
and U1642 (N_1642,N_1597,N_1619);
nor U1643 (N_1643,N_1582,N_1587);
nand U1644 (N_1644,N_1561,N_1590);
nor U1645 (N_1645,N_1611,N_1584);
xor U1646 (N_1646,N_1612,N_1569);
xnor U1647 (N_1647,N_1583,N_1568);
nor U1648 (N_1648,N_1595,N_1604);
nand U1649 (N_1649,N_1605,N_1592);
nor U1650 (N_1650,N_1579,N_1571);
nand U1651 (N_1651,N_1595,N_1614);
or U1652 (N_1652,N_1618,N_1570);
xnor U1653 (N_1653,N_1619,N_1574);
or U1654 (N_1654,N_1573,N_1586);
and U1655 (N_1655,N_1596,N_1582);
nor U1656 (N_1656,N_1570,N_1564);
nand U1657 (N_1657,N_1567,N_1591);
nand U1658 (N_1658,N_1616,N_1573);
nor U1659 (N_1659,N_1568,N_1612);
and U1660 (N_1660,N_1602,N_1604);
or U1661 (N_1661,N_1614,N_1569);
or U1662 (N_1662,N_1604,N_1573);
nor U1663 (N_1663,N_1587,N_1608);
or U1664 (N_1664,N_1615,N_1607);
or U1665 (N_1665,N_1573,N_1570);
xor U1666 (N_1666,N_1593,N_1588);
and U1667 (N_1667,N_1607,N_1610);
and U1668 (N_1668,N_1578,N_1607);
and U1669 (N_1669,N_1567,N_1595);
xnor U1670 (N_1670,N_1601,N_1576);
or U1671 (N_1671,N_1589,N_1619);
nor U1672 (N_1672,N_1611,N_1581);
and U1673 (N_1673,N_1617,N_1597);
nand U1674 (N_1674,N_1596,N_1570);
or U1675 (N_1675,N_1618,N_1575);
nor U1676 (N_1676,N_1598,N_1618);
or U1677 (N_1677,N_1573,N_1587);
nand U1678 (N_1678,N_1600,N_1610);
nand U1679 (N_1679,N_1566,N_1603);
nor U1680 (N_1680,N_1675,N_1676);
or U1681 (N_1681,N_1649,N_1660);
nand U1682 (N_1682,N_1643,N_1669);
nor U1683 (N_1683,N_1646,N_1678);
nand U1684 (N_1684,N_1629,N_1647);
or U1685 (N_1685,N_1664,N_1638);
nand U1686 (N_1686,N_1628,N_1621);
nand U1687 (N_1687,N_1671,N_1656);
xnor U1688 (N_1688,N_1650,N_1659);
and U1689 (N_1689,N_1654,N_1623);
xnor U1690 (N_1690,N_1667,N_1624);
nand U1691 (N_1691,N_1634,N_1627);
xnor U1692 (N_1692,N_1639,N_1652);
nor U1693 (N_1693,N_1625,N_1672);
xor U1694 (N_1694,N_1653,N_1679);
and U1695 (N_1695,N_1640,N_1674);
nand U1696 (N_1696,N_1670,N_1632);
xnor U1697 (N_1697,N_1631,N_1665);
or U1698 (N_1698,N_1663,N_1644);
or U1699 (N_1699,N_1648,N_1651);
or U1700 (N_1700,N_1668,N_1633);
nor U1701 (N_1701,N_1630,N_1645);
or U1702 (N_1702,N_1637,N_1626);
nor U1703 (N_1703,N_1642,N_1655);
nand U1704 (N_1704,N_1677,N_1673);
nand U1705 (N_1705,N_1658,N_1636);
nor U1706 (N_1706,N_1635,N_1661);
xor U1707 (N_1707,N_1662,N_1666);
xor U1708 (N_1708,N_1657,N_1620);
or U1709 (N_1709,N_1641,N_1622);
nor U1710 (N_1710,N_1622,N_1658);
and U1711 (N_1711,N_1659,N_1658);
and U1712 (N_1712,N_1624,N_1676);
nor U1713 (N_1713,N_1649,N_1665);
nor U1714 (N_1714,N_1629,N_1641);
nor U1715 (N_1715,N_1654,N_1647);
or U1716 (N_1716,N_1639,N_1637);
nor U1717 (N_1717,N_1672,N_1671);
or U1718 (N_1718,N_1657,N_1642);
and U1719 (N_1719,N_1635,N_1641);
nor U1720 (N_1720,N_1663,N_1620);
nor U1721 (N_1721,N_1661,N_1659);
or U1722 (N_1722,N_1640,N_1675);
xor U1723 (N_1723,N_1656,N_1661);
and U1724 (N_1724,N_1675,N_1674);
and U1725 (N_1725,N_1642,N_1645);
and U1726 (N_1726,N_1626,N_1651);
nor U1727 (N_1727,N_1675,N_1667);
nand U1728 (N_1728,N_1678,N_1651);
nand U1729 (N_1729,N_1667,N_1671);
nor U1730 (N_1730,N_1644,N_1630);
or U1731 (N_1731,N_1666,N_1640);
xor U1732 (N_1732,N_1635,N_1629);
or U1733 (N_1733,N_1666,N_1639);
nor U1734 (N_1734,N_1645,N_1675);
nand U1735 (N_1735,N_1646,N_1663);
or U1736 (N_1736,N_1623,N_1678);
nand U1737 (N_1737,N_1671,N_1632);
nor U1738 (N_1738,N_1635,N_1632);
and U1739 (N_1739,N_1650,N_1660);
nor U1740 (N_1740,N_1711,N_1734);
nand U1741 (N_1741,N_1686,N_1737);
and U1742 (N_1742,N_1703,N_1729);
nor U1743 (N_1743,N_1722,N_1715);
xnor U1744 (N_1744,N_1698,N_1733);
and U1745 (N_1745,N_1732,N_1738);
nand U1746 (N_1746,N_1714,N_1697);
or U1747 (N_1747,N_1702,N_1706);
or U1748 (N_1748,N_1723,N_1688);
or U1749 (N_1749,N_1689,N_1685);
nand U1750 (N_1750,N_1708,N_1719);
xor U1751 (N_1751,N_1713,N_1728);
and U1752 (N_1752,N_1700,N_1682);
and U1753 (N_1753,N_1687,N_1680);
nand U1754 (N_1754,N_1699,N_1730);
nand U1755 (N_1755,N_1727,N_1712);
and U1756 (N_1756,N_1695,N_1683);
nor U1757 (N_1757,N_1693,N_1718);
and U1758 (N_1758,N_1701,N_1731);
or U1759 (N_1759,N_1690,N_1696);
or U1760 (N_1760,N_1720,N_1709);
and U1761 (N_1761,N_1704,N_1707);
nand U1762 (N_1762,N_1705,N_1717);
xor U1763 (N_1763,N_1716,N_1694);
or U1764 (N_1764,N_1725,N_1739);
or U1765 (N_1765,N_1681,N_1721);
nand U1766 (N_1766,N_1692,N_1710);
xnor U1767 (N_1767,N_1724,N_1691);
xnor U1768 (N_1768,N_1726,N_1735);
and U1769 (N_1769,N_1684,N_1736);
and U1770 (N_1770,N_1694,N_1715);
or U1771 (N_1771,N_1717,N_1725);
xnor U1772 (N_1772,N_1695,N_1687);
and U1773 (N_1773,N_1700,N_1734);
nand U1774 (N_1774,N_1695,N_1705);
or U1775 (N_1775,N_1731,N_1712);
or U1776 (N_1776,N_1717,N_1727);
and U1777 (N_1777,N_1700,N_1712);
nand U1778 (N_1778,N_1681,N_1732);
or U1779 (N_1779,N_1716,N_1719);
and U1780 (N_1780,N_1680,N_1691);
xor U1781 (N_1781,N_1718,N_1735);
nand U1782 (N_1782,N_1733,N_1680);
and U1783 (N_1783,N_1683,N_1730);
and U1784 (N_1784,N_1699,N_1721);
and U1785 (N_1785,N_1697,N_1719);
and U1786 (N_1786,N_1729,N_1739);
nor U1787 (N_1787,N_1705,N_1681);
nor U1788 (N_1788,N_1721,N_1687);
nand U1789 (N_1789,N_1711,N_1681);
and U1790 (N_1790,N_1694,N_1724);
and U1791 (N_1791,N_1694,N_1729);
and U1792 (N_1792,N_1697,N_1693);
nor U1793 (N_1793,N_1718,N_1707);
nand U1794 (N_1794,N_1703,N_1682);
and U1795 (N_1795,N_1690,N_1716);
or U1796 (N_1796,N_1697,N_1712);
nor U1797 (N_1797,N_1688,N_1712);
or U1798 (N_1798,N_1703,N_1688);
nand U1799 (N_1799,N_1739,N_1738);
xnor U1800 (N_1800,N_1757,N_1741);
nand U1801 (N_1801,N_1797,N_1762);
xor U1802 (N_1802,N_1747,N_1792);
or U1803 (N_1803,N_1796,N_1758);
nand U1804 (N_1804,N_1787,N_1780);
xnor U1805 (N_1805,N_1759,N_1771);
and U1806 (N_1806,N_1786,N_1773);
nor U1807 (N_1807,N_1768,N_1798);
xor U1808 (N_1808,N_1751,N_1745);
nor U1809 (N_1809,N_1761,N_1777);
and U1810 (N_1810,N_1770,N_1775);
nor U1811 (N_1811,N_1779,N_1794);
xor U1812 (N_1812,N_1750,N_1799);
nor U1813 (N_1813,N_1756,N_1767);
xor U1814 (N_1814,N_1785,N_1760);
and U1815 (N_1815,N_1763,N_1766);
nand U1816 (N_1816,N_1784,N_1748);
and U1817 (N_1817,N_1776,N_1769);
nor U1818 (N_1818,N_1742,N_1778);
and U1819 (N_1819,N_1783,N_1765);
or U1820 (N_1820,N_1791,N_1782);
and U1821 (N_1821,N_1743,N_1793);
nor U1822 (N_1822,N_1772,N_1795);
or U1823 (N_1823,N_1752,N_1749);
and U1824 (N_1824,N_1754,N_1746);
or U1825 (N_1825,N_1744,N_1781);
and U1826 (N_1826,N_1764,N_1753);
nor U1827 (N_1827,N_1790,N_1788);
nand U1828 (N_1828,N_1740,N_1755);
nand U1829 (N_1829,N_1774,N_1789);
xor U1830 (N_1830,N_1756,N_1752);
or U1831 (N_1831,N_1745,N_1762);
or U1832 (N_1832,N_1755,N_1752);
xor U1833 (N_1833,N_1756,N_1797);
nor U1834 (N_1834,N_1742,N_1777);
and U1835 (N_1835,N_1752,N_1776);
and U1836 (N_1836,N_1793,N_1790);
xnor U1837 (N_1837,N_1746,N_1786);
xnor U1838 (N_1838,N_1755,N_1789);
nand U1839 (N_1839,N_1774,N_1778);
or U1840 (N_1840,N_1744,N_1759);
nor U1841 (N_1841,N_1758,N_1748);
nand U1842 (N_1842,N_1761,N_1748);
or U1843 (N_1843,N_1768,N_1771);
nor U1844 (N_1844,N_1790,N_1775);
nand U1845 (N_1845,N_1796,N_1743);
or U1846 (N_1846,N_1744,N_1778);
or U1847 (N_1847,N_1763,N_1783);
and U1848 (N_1848,N_1786,N_1749);
nor U1849 (N_1849,N_1746,N_1767);
nor U1850 (N_1850,N_1764,N_1744);
nand U1851 (N_1851,N_1793,N_1781);
nand U1852 (N_1852,N_1748,N_1756);
nor U1853 (N_1853,N_1758,N_1745);
nand U1854 (N_1854,N_1772,N_1786);
nand U1855 (N_1855,N_1762,N_1741);
nand U1856 (N_1856,N_1749,N_1747);
xnor U1857 (N_1857,N_1766,N_1785);
xnor U1858 (N_1858,N_1764,N_1773);
and U1859 (N_1859,N_1783,N_1761);
and U1860 (N_1860,N_1819,N_1822);
and U1861 (N_1861,N_1821,N_1832);
xor U1862 (N_1862,N_1820,N_1825);
or U1863 (N_1863,N_1836,N_1818);
nand U1864 (N_1864,N_1817,N_1829);
and U1865 (N_1865,N_1846,N_1856);
nand U1866 (N_1866,N_1813,N_1838);
nor U1867 (N_1867,N_1844,N_1851);
xnor U1868 (N_1868,N_1839,N_1808);
or U1869 (N_1869,N_1833,N_1824);
and U1870 (N_1870,N_1811,N_1831);
or U1871 (N_1871,N_1853,N_1827);
nor U1872 (N_1872,N_1852,N_1828);
nor U1873 (N_1873,N_1850,N_1843);
xnor U1874 (N_1874,N_1823,N_1830);
xor U1875 (N_1875,N_1801,N_1815);
nor U1876 (N_1876,N_1841,N_1849);
or U1877 (N_1877,N_1847,N_1859);
nand U1878 (N_1878,N_1855,N_1848);
and U1879 (N_1879,N_1840,N_1854);
nor U1880 (N_1880,N_1804,N_1816);
nand U1881 (N_1881,N_1842,N_1857);
nand U1882 (N_1882,N_1806,N_1834);
and U1883 (N_1883,N_1826,N_1835);
nand U1884 (N_1884,N_1810,N_1809);
or U1885 (N_1885,N_1837,N_1805);
nor U1886 (N_1886,N_1803,N_1802);
nor U1887 (N_1887,N_1807,N_1845);
nand U1888 (N_1888,N_1812,N_1858);
and U1889 (N_1889,N_1800,N_1814);
nand U1890 (N_1890,N_1853,N_1811);
and U1891 (N_1891,N_1853,N_1801);
or U1892 (N_1892,N_1805,N_1851);
or U1893 (N_1893,N_1836,N_1820);
nor U1894 (N_1894,N_1814,N_1804);
and U1895 (N_1895,N_1853,N_1835);
nor U1896 (N_1896,N_1858,N_1832);
or U1897 (N_1897,N_1815,N_1851);
nand U1898 (N_1898,N_1852,N_1842);
or U1899 (N_1899,N_1815,N_1854);
nor U1900 (N_1900,N_1821,N_1833);
nand U1901 (N_1901,N_1813,N_1832);
nor U1902 (N_1902,N_1813,N_1839);
nand U1903 (N_1903,N_1850,N_1819);
and U1904 (N_1904,N_1812,N_1841);
and U1905 (N_1905,N_1801,N_1839);
xnor U1906 (N_1906,N_1847,N_1855);
xor U1907 (N_1907,N_1822,N_1839);
and U1908 (N_1908,N_1838,N_1804);
and U1909 (N_1909,N_1830,N_1810);
nor U1910 (N_1910,N_1821,N_1819);
and U1911 (N_1911,N_1823,N_1802);
and U1912 (N_1912,N_1825,N_1827);
nand U1913 (N_1913,N_1825,N_1837);
nand U1914 (N_1914,N_1815,N_1805);
nor U1915 (N_1915,N_1833,N_1830);
or U1916 (N_1916,N_1809,N_1858);
nor U1917 (N_1917,N_1823,N_1828);
nand U1918 (N_1918,N_1801,N_1859);
or U1919 (N_1919,N_1838,N_1859);
xnor U1920 (N_1920,N_1899,N_1879);
or U1921 (N_1921,N_1910,N_1919);
or U1922 (N_1922,N_1864,N_1878);
and U1923 (N_1923,N_1907,N_1904);
or U1924 (N_1924,N_1862,N_1860);
or U1925 (N_1925,N_1898,N_1888);
or U1926 (N_1926,N_1918,N_1915);
and U1927 (N_1927,N_1886,N_1874);
nor U1928 (N_1928,N_1877,N_1909);
and U1929 (N_1929,N_1885,N_1913);
nand U1930 (N_1930,N_1865,N_1916);
or U1931 (N_1931,N_1914,N_1901);
nand U1932 (N_1932,N_1917,N_1883);
nor U1933 (N_1933,N_1897,N_1892);
nor U1934 (N_1934,N_1871,N_1896);
or U1935 (N_1935,N_1880,N_1867);
and U1936 (N_1936,N_1873,N_1881);
or U1937 (N_1937,N_1895,N_1905);
and U1938 (N_1938,N_1876,N_1866);
nor U1939 (N_1939,N_1893,N_1882);
or U1940 (N_1940,N_1887,N_1912);
nand U1941 (N_1941,N_1869,N_1908);
nor U1942 (N_1942,N_1902,N_1875);
and U1943 (N_1943,N_1906,N_1890);
xnor U1944 (N_1944,N_1900,N_1863);
nor U1945 (N_1945,N_1868,N_1870);
nor U1946 (N_1946,N_1861,N_1891);
or U1947 (N_1947,N_1872,N_1894);
or U1948 (N_1948,N_1911,N_1889);
nor U1949 (N_1949,N_1884,N_1903);
nand U1950 (N_1950,N_1870,N_1863);
xor U1951 (N_1951,N_1863,N_1860);
and U1952 (N_1952,N_1868,N_1874);
nand U1953 (N_1953,N_1882,N_1908);
nor U1954 (N_1954,N_1886,N_1876);
nor U1955 (N_1955,N_1919,N_1884);
nand U1956 (N_1956,N_1902,N_1890);
xnor U1957 (N_1957,N_1903,N_1914);
and U1958 (N_1958,N_1883,N_1888);
nor U1959 (N_1959,N_1879,N_1904);
and U1960 (N_1960,N_1869,N_1862);
or U1961 (N_1961,N_1897,N_1874);
nor U1962 (N_1962,N_1879,N_1902);
or U1963 (N_1963,N_1867,N_1874);
nand U1964 (N_1964,N_1872,N_1896);
or U1965 (N_1965,N_1865,N_1893);
nor U1966 (N_1966,N_1918,N_1878);
nand U1967 (N_1967,N_1889,N_1894);
and U1968 (N_1968,N_1875,N_1897);
and U1969 (N_1969,N_1878,N_1866);
nand U1970 (N_1970,N_1884,N_1911);
nand U1971 (N_1971,N_1892,N_1902);
nand U1972 (N_1972,N_1862,N_1909);
and U1973 (N_1973,N_1918,N_1906);
and U1974 (N_1974,N_1899,N_1906);
nand U1975 (N_1975,N_1882,N_1867);
or U1976 (N_1976,N_1891,N_1902);
nor U1977 (N_1977,N_1871,N_1881);
xor U1978 (N_1978,N_1902,N_1889);
nand U1979 (N_1979,N_1917,N_1899);
xnor U1980 (N_1980,N_1920,N_1959);
and U1981 (N_1981,N_1949,N_1968);
or U1982 (N_1982,N_1958,N_1940);
xor U1983 (N_1983,N_1939,N_1977);
or U1984 (N_1984,N_1957,N_1924);
and U1985 (N_1985,N_1974,N_1976);
or U1986 (N_1986,N_1925,N_1944);
or U1987 (N_1987,N_1946,N_1954);
nor U1988 (N_1988,N_1978,N_1937);
and U1989 (N_1989,N_1969,N_1966);
nand U1990 (N_1990,N_1960,N_1934);
and U1991 (N_1991,N_1930,N_1956);
and U1992 (N_1992,N_1971,N_1942);
and U1993 (N_1993,N_1947,N_1941);
or U1994 (N_1994,N_1928,N_1975);
and U1995 (N_1995,N_1936,N_1933);
xor U1996 (N_1996,N_1931,N_1955);
nand U1997 (N_1997,N_1923,N_1965);
nor U1998 (N_1998,N_1979,N_1945);
nor U1999 (N_1999,N_1926,N_1935);
and U2000 (N_2000,N_1952,N_1932);
or U2001 (N_2001,N_1921,N_1972);
nand U2002 (N_2002,N_1953,N_1948);
or U2003 (N_2003,N_1938,N_1973);
nor U2004 (N_2004,N_1964,N_1963);
and U2005 (N_2005,N_1922,N_1950);
and U2006 (N_2006,N_1962,N_1927);
and U2007 (N_2007,N_1951,N_1970);
nand U2008 (N_2008,N_1929,N_1943);
and U2009 (N_2009,N_1967,N_1961);
nand U2010 (N_2010,N_1937,N_1920);
nor U2011 (N_2011,N_1947,N_1968);
nor U2012 (N_2012,N_1968,N_1922);
or U2013 (N_2013,N_1977,N_1946);
nand U2014 (N_2014,N_1947,N_1963);
nor U2015 (N_2015,N_1960,N_1930);
or U2016 (N_2016,N_1951,N_1926);
or U2017 (N_2017,N_1948,N_1943);
and U2018 (N_2018,N_1957,N_1967);
nand U2019 (N_2019,N_1922,N_1965);
xnor U2020 (N_2020,N_1950,N_1941);
nor U2021 (N_2021,N_1948,N_1946);
or U2022 (N_2022,N_1971,N_1948);
nand U2023 (N_2023,N_1946,N_1925);
nand U2024 (N_2024,N_1969,N_1934);
nand U2025 (N_2025,N_1979,N_1946);
and U2026 (N_2026,N_1964,N_1930);
or U2027 (N_2027,N_1970,N_1958);
and U2028 (N_2028,N_1949,N_1953);
xnor U2029 (N_2029,N_1979,N_1950);
and U2030 (N_2030,N_1922,N_1941);
nor U2031 (N_2031,N_1954,N_1957);
or U2032 (N_2032,N_1940,N_1949);
or U2033 (N_2033,N_1931,N_1926);
or U2034 (N_2034,N_1933,N_1976);
nand U2035 (N_2035,N_1971,N_1977);
nand U2036 (N_2036,N_1948,N_1966);
nor U2037 (N_2037,N_1948,N_1956);
and U2038 (N_2038,N_1931,N_1929);
xor U2039 (N_2039,N_1923,N_1953);
and U2040 (N_2040,N_1987,N_2032);
and U2041 (N_2041,N_2010,N_1990);
nand U2042 (N_2042,N_1998,N_2026);
xnor U2043 (N_2043,N_2012,N_2011);
and U2044 (N_2044,N_1997,N_1991);
and U2045 (N_2045,N_2016,N_1993);
nand U2046 (N_2046,N_2003,N_2007);
nor U2047 (N_2047,N_2014,N_2006);
nand U2048 (N_2048,N_2039,N_1985);
nor U2049 (N_2049,N_1981,N_2015);
xor U2050 (N_2050,N_1994,N_2028);
nand U2051 (N_2051,N_1983,N_1999);
nor U2052 (N_2052,N_2029,N_2004);
nor U2053 (N_2053,N_2027,N_2019);
nor U2054 (N_2054,N_2020,N_2013);
and U2055 (N_2055,N_2034,N_2024);
nand U2056 (N_2056,N_2009,N_2001);
and U2057 (N_2057,N_1992,N_2036);
nand U2058 (N_2058,N_2033,N_1996);
or U2059 (N_2059,N_1988,N_2008);
nand U2060 (N_2060,N_2018,N_2021);
xnor U2061 (N_2061,N_1982,N_2037);
or U2062 (N_2062,N_2038,N_2023);
and U2063 (N_2063,N_2002,N_1980);
nand U2064 (N_2064,N_2031,N_1995);
nand U2065 (N_2065,N_2005,N_2025);
and U2066 (N_2066,N_2000,N_2017);
nand U2067 (N_2067,N_2030,N_1984);
and U2068 (N_2068,N_1986,N_1989);
nor U2069 (N_2069,N_2035,N_2022);
xnor U2070 (N_2070,N_2025,N_1982);
and U2071 (N_2071,N_2023,N_1998);
xor U2072 (N_2072,N_1988,N_2027);
nor U2073 (N_2073,N_1998,N_2017);
and U2074 (N_2074,N_2006,N_1998);
nand U2075 (N_2075,N_2029,N_2008);
or U2076 (N_2076,N_2001,N_2000);
nor U2077 (N_2077,N_1983,N_1982);
or U2078 (N_2078,N_1988,N_2033);
nand U2079 (N_2079,N_2035,N_2028);
nor U2080 (N_2080,N_2017,N_1989);
xor U2081 (N_2081,N_1995,N_2014);
nor U2082 (N_2082,N_2022,N_1998);
xnor U2083 (N_2083,N_2029,N_2031);
nand U2084 (N_2084,N_2031,N_1994);
xnor U2085 (N_2085,N_1996,N_2039);
nor U2086 (N_2086,N_2017,N_2015);
nand U2087 (N_2087,N_1989,N_2011);
or U2088 (N_2088,N_1985,N_2017);
and U2089 (N_2089,N_2035,N_1992);
and U2090 (N_2090,N_1991,N_1985);
and U2091 (N_2091,N_2031,N_2026);
nand U2092 (N_2092,N_2014,N_2035);
nand U2093 (N_2093,N_1986,N_2023);
nor U2094 (N_2094,N_1994,N_2037);
and U2095 (N_2095,N_2020,N_2001);
or U2096 (N_2096,N_2002,N_2017);
or U2097 (N_2097,N_2002,N_1993);
and U2098 (N_2098,N_1997,N_2006);
or U2099 (N_2099,N_2026,N_2005);
nor U2100 (N_2100,N_2090,N_2092);
nor U2101 (N_2101,N_2042,N_2057);
xnor U2102 (N_2102,N_2062,N_2072);
or U2103 (N_2103,N_2081,N_2048);
xor U2104 (N_2104,N_2096,N_2055);
nand U2105 (N_2105,N_2051,N_2095);
nand U2106 (N_2106,N_2066,N_2063);
xor U2107 (N_2107,N_2074,N_2068);
or U2108 (N_2108,N_2086,N_2098);
nand U2109 (N_2109,N_2044,N_2041);
nor U2110 (N_2110,N_2078,N_2084);
xnor U2111 (N_2111,N_2060,N_2064);
nor U2112 (N_2112,N_2085,N_2099);
and U2113 (N_2113,N_2091,N_2056);
nand U2114 (N_2114,N_2075,N_2069);
and U2115 (N_2115,N_2061,N_2070);
and U2116 (N_2116,N_2058,N_2049);
nand U2117 (N_2117,N_2054,N_2077);
or U2118 (N_2118,N_2047,N_2094);
nor U2119 (N_2119,N_2045,N_2065);
nor U2120 (N_2120,N_2059,N_2046);
nand U2121 (N_2121,N_2076,N_2087);
and U2122 (N_2122,N_2093,N_2097);
nor U2123 (N_2123,N_2050,N_2071);
and U2124 (N_2124,N_2083,N_2088);
nand U2125 (N_2125,N_2089,N_2052);
and U2126 (N_2126,N_2079,N_2080);
nand U2127 (N_2127,N_2082,N_2053);
or U2128 (N_2128,N_2040,N_2073);
nor U2129 (N_2129,N_2067,N_2043);
and U2130 (N_2130,N_2094,N_2078);
or U2131 (N_2131,N_2056,N_2052);
and U2132 (N_2132,N_2046,N_2092);
or U2133 (N_2133,N_2048,N_2072);
and U2134 (N_2134,N_2072,N_2056);
and U2135 (N_2135,N_2056,N_2066);
nand U2136 (N_2136,N_2063,N_2052);
or U2137 (N_2137,N_2050,N_2058);
nand U2138 (N_2138,N_2089,N_2057);
or U2139 (N_2139,N_2082,N_2058);
and U2140 (N_2140,N_2069,N_2044);
and U2141 (N_2141,N_2086,N_2048);
or U2142 (N_2142,N_2074,N_2066);
and U2143 (N_2143,N_2071,N_2081);
or U2144 (N_2144,N_2093,N_2067);
and U2145 (N_2145,N_2046,N_2054);
or U2146 (N_2146,N_2091,N_2092);
nand U2147 (N_2147,N_2078,N_2091);
xnor U2148 (N_2148,N_2078,N_2082);
or U2149 (N_2149,N_2044,N_2097);
nor U2150 (N_2150,N_2047,N_2063);
and U2151 (N_2151,N_2088,N_2068);
or U2152 (N_2152,N_2088,N_2080);
and U2153 (N_2153,N_2065,N_2095);
or U2154 (N_2154,N_2070,N_2055);
or U2155 (N_2155,N_2077,N_2068);
nand U2156 (N_2156,N_2042,N_2079);
nand U2157 (N_2157,N_2075,N_2066);
nor U2158 (N_2158,N_2055,N_2091);
nor U2159 (N_2159,N_2062,N_2098);
nand U2160 (N_2160,N_2102,N_2139);
xor U2161 (N_2161,N_2135,N_2124);
xnor U2162 (N_2162,N_2159,N_2152);
xnor U2163 (N_2163,N_2157,N_2141);
and U2164 (N_2164,N_2132,N_2133);
nand U2165 (N_2165,N_2111,N_2105);
nor U2166 (N_2166,N_2110,N_2113);
or U2167 (N_2167,N_2137,N_2146);
or U2168 (N_2168,N_2158,N_2115);
nand U2169 (N_2169,N_2140,N_2126);
or U2170 (N_2170,N_2117,N_2119);
nor U2171 (N_2171,N_2109,N_2130);
nand U2172 (N_2172,N_2143,N_2122);
and U2173 (N_2173,N_2101,N_2149);
nor U2174 (N_2174,N_2120,N_2144);
or U2175 (N_2175,N_2108,N_2153);
or U2176 (N_2176,N_2134,N_2145);
and U2177 (N_2177,N_2106,N_2121);
or U2178 (N_2178,N_2154,N_2123);
or U2179 (N_2179,N_2138,N_2103);
or U2180 (N_2180,N_2114,N_2148);
or U2181 (N_2181,N_2125,N_2136);
and U2182 (N_2182,N_2147,N_2116);
nor U2183 (N_2183,N_2104,N_2127);
and U2184 (N_2184,N_2128,N_2150);
xnor U2185 (N_2185,N_2155,N_2107);
or U2186 (N_2186,N_2142,N_2100);
nor U2187 (N_2187,N_2129,N_2156);
or U2188 (N_2188,N_2118,N_2112);
or U2189 (N_2189,N_2151,N_2131);
xnor U2190 (N_2190,N_2130,N_2155);
nand U2191 (N_2191,N_2138,N_2128);
xnor U2192 (N_2192,N_2103,N_2117);
and U2193 (N_2193,N_2111,N_2113);
nor U2194 (N_2194,N_2141,N_2107);
or U2195 (N_2195,N_2100,N_2107);
nor U2196 (N_2196,N_2125,N_2143);
nor U2197 (N_2197,N_2148,N_2154);
nor U2198 (N_2198,N_2146,N_2101);
nand U2199 (N_2199,N_2144,N_2143);
nand U2200 (N_2200,N_2142,N_2130);
nor U2201 (N_2201,N_2156,N_2130);
xor U2202 (N_2202,N_2102,N_2106);
and U2203 (N_2203,N_2157,N_2119);
nor U2204 (N_2204,N_2131,N_2122);
and U2205 (N_2205,N_2111,N_2152);
nor U2206 (N_2206,N_2144,N_2147);
or U2207 (N_2207,N_2109,N_2145);
or U2208 (N_2208,N_2112,N_2107);
or U2209 (N_2209,N_2119,N_2149);
or U2210 (N_2210,N_2111,N_2149);
nor U2211 (N_2211,N_2132,N_2151);
nor U2212 (N_2212,N_2144,N_2106);
or U2213 (N_2213,N_2151,N_2137);
nand U2214 (N_2214,N_2158,N_2113);
nand U2215 (N_2215,N_2104,N_2110);
or U2216 (N_2216,N_2159,N_2102);
and U2217 (N_2217,N_2117,N_2101);
nor U2218 (N_2218,N_2136,N_2140);
nor U2219 (N_2219,N_2103,N_2121);
or U2220 (N_2220,N_2216,N_2218);
xnor U2221 (N_2221,N_2162,N_2207);
or U2222 (N_2222,N_2172,N_2202);
and U2223 (N_2223,N_2176,N_2199);
and U2224 (N_2224,N_2210,N_2164);
or U2225 (N_2225,N_2219,N_2203);
xor U2226 (N_2226,N_2166,N_2188);
nor U2227 (N_2227,N_2195,N_2169);
and U2228 (N_2228,N_2167,N_2198);
or U2229 (N_2229,N_2175,N_2171);
nor U2230 (N_2230,N_2180,N_2205);
and U2231 (N_2231,N_2212,N_2168);
nand U2232 (N_2232,N_2174,N_2213);
nand U2233 (N_2233,N_2170,N_2178);
xnor U2234 (N_2234,N_2190,N_2182);
xnor U2235 (N_2235,N_2217,N_2208);
nor U2236 (N_2236,N_2193,N_2184);
or U2237 (N_2237,N_2192,N_2191);
xnor U2238 (N_2238,N_2160,N_2200);
nor U2239 (N_2239,N_2179,N_2185);
nand U2240 (N_2240,N_2173,N_2183);
nand U2241 (N_2241,N_2201,N_2163);
and U2242 (N_2242,N_2204,N_2197);
and U2243 (N_2243,N_2211,N_2161);
and U2244 (N_2244,N_2177,N_2215);
nor U2245 (N_2245,N_2181,N_2187);
nor U2246 (N_2246,N_2196,N_2206);
nor U2247 (N_2247,N_2214,N_2194);
or U2248 (N_2248,N_2209,N_2186);
nor U2249 (N_2249,N_2189,N_2165);
nor U2250 (N_2250,N_2189,N_2201);
xnor U2251 (N_2251,N_2169,N_2199);
nand U2252 (N_2252,N_2189,N_2214);
nor U2253 (N_2253,N_2162,N_2187);
or U2254 (N_2254,N_2200,N_2182);
nand U2255 (N_2255,N_2178,N_2200);
nand U2256 (N_2256,N_2174,N_2204);
and U2257 (N_2257,N_2200,N_2189);
or U2258 (N_2258,N_2191,N_2172);
or U2259 (N_2259,N_2161,N_2216);
and U2260 (N_2260,N_2201,N_2193);
nor U2261 (N_2261,N_2162,N_2189);
nand U2262 (N_2262,N_2182,N_2205);
and U2263 (N_2263,N_2201,N_2172);
nand U2264 (N_2264,N_2164,N_2205);
or U2265 (N_2265,N_2162,N_2169);
nand U2266 (N_2266,N_2210,N_2217);
nor U2267 (N_2267,N_2177,N_2174);
or U2268 (N_2268,N_2217,N_2175);
or U2269 (N_2269,N_2166,N_2161);
nand U2270 (N_2270,N_2164,N_2208);
nor U2271 (N_2271,N_2161,N_2178);
nand U2272 (N_2272,N_2183,N_2196);
or U2273 (N_2273,N_2209,N_2163);
xnor U2274 (N_2274,N_2184,N_2211);
nand U2275 (N_2275,N_2173,N_2200);
nand U2276 (N_2276,N_2201,N_2179);
nor U2277 (N_2277,N_2173,N_2193);
nor U2278 (N_2278,N_2171,N_2160);
nand U2279 (N_2279,N_2211,N_2160);
nor U2280 (N_2280,N_2230,N_2251);
or U2281 (N_2281,N_2241,N_2277);
nor U2282 (N_2282,N_2271,N_2260);
nor U2283 (N_2283,N_2265,N_2222);
and U2284 (N_2284,N_2262,N_2247);
nand U2285 (N_2285,N_2267,N_2276);
xor U2286 (N_2286,N_2226,N_2254);
nor U2287 (N_2287,N_2231,N_2257);
and U2288 (N_2288,N_2272,N_2255);
nand U2289 (N_2289,N_2263,N_2279);
and U2290 (N_2290,N_2261,N_2238);
xnor U2291 (N_2291,N_2269,N_2259);
nor U2292 (N_2292,N_2268,N_2234);
nand U2293 (N_2293,N_2275,N_2227);
nor U2294 (N_2294,N_2246,N_2252);
and U2295 (N_2295,N_2274,N_2244);
or U2296 (N_2296,N_2228,N_2236);
nand U2297 (N_2297,N_2240,N_2253);
or U2298 (N_2298,N_2245,N_2264);
or U2299 (N_2299,N_2229,N_2221);
nor U2300 (N_2300,N_2250,N_2248);
nor U2301 (N_2301,N_2220,N_2270);
nor U2302 (N_2302,N_2237,N_2239);
nor U2303 (N_2303,N_2242,N_2223);
nand U2304 (N_2304,N_2266,N_2225);
xnor U2305 (N_2305,N_2243,N_2278);
or U2306 (N_2306,N_2249,N_2224);
and U2307 (N_2307,N_2258,N_2273);
xor U2308 (N_2308,N_2233,N_2232);
xnor U2309 (N_2309,N_2235,N_2256);
nand U2310 (N_2310,N_2256,N_2226);
and U2311 (N_2311,N_2279,N_2260);
nor U2312 (N_2312,N_2226,N_2262);
or U2313 (N_2313,N_2235,N_2226);
nor U2314 (N_2314,N_2228,N_2234);
or U2315 (N_2315,N_2269,N_2258);
xnor U2316 (N_2316,N_2266,N_2240);
nand U2317 (N_2317,N_2265,N_2228);
nor U2318 (N_2318,N_2238,N_2229);
or U2319 (N_2319,N_2275,N_2246);
and U2320 (N_2320,N_2223,N_2268);
nor U2321 (N_2321,N_2271,N_2239);
nand U2322 (N_2322,N_2222,N_2234);
and U2323 (N_2323,N_2240,N_2247);
nand U2324 (N_2324,N_2263,N_2268);
or U2325 (N_2325,N_2235,N_2222);
or U2326 (N_2326,N_2264,N_2231);
nor U2327 (N_2327,N_2228,N_2248);
nand U2328 (N_2328,N_2263,N_2270);
nand U2329 (N_2329,N_2238,N_2259);
and U2330 (N_2330,N_2235,N_2246);
nor U2331 (N_2331,N_2262,N_2258);
or U2332 (N_2332,N_2266,N_2246);
nand U2333 (N_2333,N_2277,N_2261);
or U2334 (N_2334,N_2279,N_2257);
or U2335 (N_2335,N_2232,N_2262);
and U2336 (N_2336,N_2239,N_2257);
or U2337 (N_2337,N_2228,N_2220);
nor U2338 (N_2338,N_2239,N_2266);
nor U2339 (N_2339,N_2242,N_2246);
nor U2340 (N_2340,N_2287,N_2295);
nor U2341 (N_2341,N_2298,N_2331);
xnor U2342 (N_2342,N_2315,N_2300);
nand U2343 (N_2343,N_2321,N_2312);
and U2344 (N_2344,N_2339,N_2283);
nor U2345 (N_2345,N_2280,N_2292);
or U2346 (N_2346,N_2304,N_2325);
nand U2347 (N_2347,N_2324,N_2286);
and U2348 (N_2348,N_2294,N_2301);
xnor U2349 (N_2349,N_2285,N_2316);
xnor U2350 (N_2350,N_2307,N_2313);
and U2351 (N_2351,N_2322,N_2333);
or U2352 (N_2352,N_2335,N_2308);
or U2353 (N_2353,N_2337,N_2332);
xnor U2354 (N_2354,N_2297,N_2302);
or U2355 (N_2355,N_2296,N_2291);
and U2356 (N_2356,N_2310,N_2327);
xor U2357 (N_2357,N_2320,N_2293);
and U2358 (N_2358,N_2290,N_2336);
nor U2359 (N_2359,N_2314,N_2282);
and U2360 (N_2360,N_2328,N_2323);
or U2361 (N_2361,N_2288,N_2281);
xor U2362 (N_2362,N_2338,N_2326);
nor U2363 (N_2363,N_2330,N_2311);
and U2364 (N_2364,N_2309,N_2306);
and U2365 (N_2365,N_2319,N_2289);
or U2366 (N_2366,N_2318,N_2303);
nor U2367 (N_2367,N_2329,N_2284);
or U2368 (N_2368,N_2305,N_2334);
nor U2369 (N_2369,N_2299,N_2317);
and U2370 (N_2370,N_2317,N_2296);
and U2371 (N_2371,N_2291,N_2302);
or U2372 (N_2372,N_2315,N_2303);
nor U2373 (N_2373,N_2318,N_2317);
nor U2374 (N_2374,N_2289,N_2301);
and U2375 (N_2375,N_2304,N_2314);
or U2376 (N_2376,N_2335,N_2311);
nor U2377 (N_2377,N_2305,N_2315);
xnor U2378 (N_2378,N_2314,N_2281);
and U2379 (N_2379,N_2330,N_2284);
nand U2380 (N_2380,N_2337,N_2301);
or U2381 (N_2381,N_2306,N_2288);
xor U2382 (N_2382,N_2335,N_2316);
or U2383 (N_2383,N_2337,N_2286);
nor U2384 (N_2384,N_2323,N_2325);
or U2385 (N_2385,N_2316,N_2288);
and U2386 (N_2386,N_2308,N_2329);
or U2387 (N_2387,N_2319,N_2335);
or U2388 (N_2388,N_2325,N_2317);
and U2389 (N_2389,N_2280,N_2325);
and U2390 (N_2390,N_2320,N_2282);
nand U2391 (N_2391,N_2324,N_2283);
and U2392 (N_2392,N_2322,N_2325);
and U2393 (N_2393,N_2312,N_2330);
xor U2394 (N_2394,N_2310,N_2309);
nor U2395 (N_2395,N_2312,N_2304);
or U2396 (N_2396,N_2283,N_2322);
and U2397 (N_2397,N_2323,N_2300);
or U2398 (N_2398,N_2329,N_2328);
and U2399 (N_2399,N_2319,N_2328);
nor U2400 (N_2400,N_2393,N_2356);
nor U2401 (N_2401,N_2380,N_2397);
nor U2402 (N_2402,N_2371,N_2350);
and U2403 (N_2403,N_2369,N_2365);
nor U2404 (N_2404,N_2383,N_2375);
xor U2405 (N_2405,N_2394,N_2392);
and U2406 (N_2406,N_2346,N_2376);
xnor U2407 (N_2407,N_2395,N_2391);
xor U2408 (N_2408,N_2368,N_2358);
nor U2409 (N_2409,N_2344,N_2367);
and U2410 (N_2410,N_2372,N_2370);
or U2411 (N_2411,N_2341,N_2353);
or U2412 (N_2412,N_2387,N_2352);
nand U2413 (N_2413,N_2382,N_2378);
nand U2414 (N_2414,N_2363,N_2357);
and U2415 (N_2415,N_2374,N_2362);
nand U2416 (N_2416,N_2340,N_2396);
and U2417 (N_2417,N_2381,N_2384);
and U2418 (N_2418,N_2359,N_2347);
nand U2419 (N_2419,N_2351,N_2385);
nor U2420 (N_2420,N_2364,N_2354);
nand U2421 (N_2421,N_2390,N_2355);
and U2422 (N_2422,N_2398,N_2345);
xor U2423 (N_2423,N_2342,N_2386);
or U2424 (N_2424,N_2343,N_2349);
nand U2425 (N_2425,N_2373,N_2388);
or U2426 (N_2426,N_2399,N_2389);
or U2427 (N_2427,N_2360,N_2348);
nand U2428 (N_2428,N_2361,N_2366);
nand U2429 (N_2429,N_2379,N_2377);
or U2430 (N_2430,N_2383,N_2374);
nand U2431 (N_2431,N_2399,N_2348);
and U2432 (N_2432,N_2386,N_2349);
nor U2433 (N_2433,N_2361,N_2390);
xnor U2434 (N_2434,N_2342,N_2397);
xor U2435 (N_2435,N_2370,N_2375);
or U2436 (N_2436,N_2363,N_2399);
nor U2437 (N_2437,N_2351,N_2377);
nand U2438 (N_2438,N_2362,N_2360);
nor U2439 (N_2439,N_2373,N_2341);
xor U2440 (N_2440,N_2387,N_2344);
and U2441 (N_2441,N_2387,N_2342);
and U2442 (N_2442,N_2392,N_2385);
xor U2443 (N_2443,N_2380,N_2359);
and U2444 (N_2444,N_2343,N_2340);
nand U2445 (N_2445,N_2368,N_2380);
and U2446 (N_2446,N_2355,N_2354);
and U2447 (N_2447,N_2340,N_2358);
xnor U2448 (N_2448,N_2355,N_2375);
nand U2449 (N_2449,N_2394,N_2340);
and U2450 (N_2450,N_2388,N_2385);
nand U2451 (N_2451,N_2341,N_2389);
nor U2452 (N_2452,N_2361,N_2371);
nand U2453 (N_2453,N_2371,N_2383);
or U2454 (N_2454,N_2390,N_2354);
nor U2455 (N_2455,N_2362,N_2342);
and U2456 (N_2456,N_2372,N_2345);
or U2457 (N_2457,N_2380,N_2381);
nand U2458 (N_2458,N_2341,N_2377);
xor U2459 (N_2459,N_2384,N_2367);
or U2460 (N_2460,N_2402,N_2432);
xor U2461 (N_2461,N_2418,N_2445);
and U2462 (N_2462,N_2452,N_2416);
nor U2463 (N_2463,N_2414,N_2449);
and U2464 (N_2464,N_2408,N_2441);
nor U2465 (N_2465,N_2437,N_2458);
nor U2466 (N_2466,N_2409,N_2407);
nor U2467 (N_2467,N_2442,N_2413);
nand U2468 (N_2468,N_2406,N_2425);
xnor U2469 (N_2469,N_2411,N_2435);
nand U2470 (N_2470,N_2446,N_2405);
or U2471 (N_2471,N_2434,N_2428);
and U2472 (N_2472,N_2422,N_2412);
nand U2473 (N_2473,N_2424,N_2415);
nand U2474 (N_2474,N_2451,N_2450);
or U2475 (N_2475,N_2401,N_2420);
or U2476 (N_2476,N_2455,N_2429);
nand U2477 (N_2477,N_2448,N_2459);
nand U2478 (N_2478,N_2404,N_2421);
xor U2479 (N_2479,N_2443,N_2433);
nor U2480 (N_2480,N_2453,N_2400);
nor U2481 (N_2481,N_2427,N_2410);
nand U2482 (N_2482,N_2447,N_2444);
nor U2483 (N_2483,N_2456,N_2438);
or U2484 (N_2484,N_2454,N_2457);
and U2485 (N_2485,N_2436,N_2430);
xor U2486 (N_2486,N_2439,N_2426);
xnor U2487 (N_2487,N_2440,N_2419);
and U2488 (N_2488,N_2417,N_2423);
or U2489 (N_2489,N_2431,N_2403);
nand U2490 (N_2490,N_2431,N_2444);
nand U2491 (N_2491,N_2416,N_2424);
nand U2492 (N_2492,N_2434,N_2416);
and U2493 (N_2493,N_2426,N_2429);
and U2494 (N_2494,N_2446,N_2436);
xor U2495 (N_2495,N_2435,N_2419);
nand U2496 (N_2496,N_2439,N_2405);
nand U2497 (N_2497,N_2420,N_2428);
or U2498 (N_2498,N_2440,N_2453);
xnor U2499 (N_2499,N_2401,N_2429);
xnor U2500 (N_2500,N_2421,N_2456);
and U2501 (N_2501,N_2404,N_2456);
and U2502 (N_2502,N_2455,N_2430);
and U2503 (N_2503,N_2402,N_2457);
and U2504 (N_2504,N_2421,N_2436);
nor U2505 (N_2505,N_2441,N_2454);
and U2506 (N_2506,N_2438,N_2454);
or U2507 (N_2507,N_2457,N_2453);
or U2508 (N_2508,N_2457,N_2459);
and U2509 (N_2509,N_2418,N_2406);
and U2510 (N_2510,N_2406,N_2404);
xor U2511 (N_2511,N_2429,N_2435);
nand U2512 (N_2512,N_2445,N_2436);
and U2513 (N_2513,N_2431,N_2405);
nor U2514 (N_2514,N_2418,N_2437);
and U2515 (N_2515,N_2425,N_2436);
nand U2516 (N_2516,N_2404,N_2455);
or U2517 (N_2517,N_2447,N_2446);
or U2518 (N_2518,N_2436,N_2419);
nand U2519 (N_2519,N_2416,N_2429);
nand U2520 (N_2520,N_2503,N_2487);
or U2521 (N_2521,N_2515,N_2475);
nor U2522 (N_2522,N_2513,N_2463);
and U2523 (N_2523,N_2502,N_2486);
nand U2524 (N_2524,N_2473,N_2471);
and U2525 (N_2525,N_2465,N_2494);
and U2526 (N_2526,N_2490,N_2491);
nor U2527 (N_2527,N_2467,N_2483);
nand U2528 (N_2528,N_2466,N_2499);
xnor U2529 (N_2529,N_2495,N_2505);
nand U2530 (N_2530,N_2511,N_2477);
nand U2531 (N_2531,N_2461,N_2492);
or U2532 (N_2532,N_2517,N_2509);
and U2533 (N_2533,N_2510,N_2508);
or U2534 (N_2534,N_2500,N_2498);
and U2535 (N_2535,N_2518,N_2469);
or U2536 (N_2536,N_2476,N_2497);
nand U2537 (N_2537,N_2474,N_2462);
or U2538 (N_2538,N_2501,N_2460);
nand U2539 (N_2539,N_2507,N_2481);
nand U2540 (N_2540,N_2489,N_2519);
or U2541 (N_2541,N_2470,N_2512);
or U2542 (N_2542,N_2478,N_2488);
and U2543 (N_2543,N_2496,N_2504);
or U2544 (N_2544,N_2479,N_2484);
and U2545 (N_2545,N_2464,N_2480);
or U2546 (N_2546,N_2468,N_2506);
nand U2547 (N_2547,N_2485,N_2514);
and U2548 (N_2548,N_2472,N_2493);
nand U2549 (N_2549,N_2482,N_2516);
and U2550 (N_2550,N_2513,N_2475);
nor U2551 (N_2551,N_2484,N_2493);
and U2552 (N_2552,N_2478,N_2474);
nor U2553 (N_2553,N_2516,N_2490);
nand U2554 (N_2554,N_2493,N_2511);
xnor U2555 (N_2555,N_2500,N_2516);
and U2556 (N_2556,N_2493,N_2512);
or U2557 (N_2557,N_2477,N_2491);
or U2558 (N_2558,N_2472,N_2499);
and U2559 (N_2559,N_2484,N_2476);
or U2560 (N_2560,N_2500,N_2472);
and U2561 (N_2561,N_2491,N_2487);
and U2562 (N_2562,N_2516,N_2504);
nor U2563 (N_2563,N_2460,N_2481);
xor U2564 (N_2564,N_2492,N_2509);
and U2565 (N_2565,N_2480,N_2510);
or U2566 (N_2566,N_2477,N_2516);
or U2567 (N_2567,N_2480,N_2499);
nand U2568 (N_2568,N_2485,N_2517);
nor U2569 (N_2569,N_2515,N_2491);
and U2570 (N_2570,N_2469,N_2463);
nand U2571 (N_2571,N_2475,N_2471);
nand U2572 (N_2572,N_2516,N_2476);
nor U2573 (N_2573,N_2505,N_2477);
and U2574 (N_2574,N_2510,N_2496);
nand U2575 (N_2575,N_2478,N_2516);
and U2576 (N_2576,N_2460,N_2468);
nand U2577 (N_2577,N_2467,N_2461);
nor U2578 (N_2578,N_2460,N_2477);
or U2579 (N_2579,N_2501,N_2477);
xor U2580 (N_2580,N_2575,N_2528);
nand U2581 (N_2581,N_2546,N_2542);
nand U2582 (N_2582,N_2524,N_2552);
nand U2583 (N_2583,N_2559,N_2566);
nor U2584 (N_2584,N_2521,N_2526);
nand U2585 (N_2585,N_2549,N_2544);
nor U2586 (N_2586,N_2569,N_2579);
or U2587 (N_2587,N_2563,N_2547);
or U2588 (N_2588,N_2520,N_2576);
nand U2589 (N_2589,N_2531,N_2555);
nor U2590 (N_2590,N_2570,N_2572);
nor U2591 (N_2591,N_2541,N_2557);
and U2592 (N_2592,N_2558,N_2561);
xor U2593 (N_2593,N_2574,N_2534);
or U2594 (N_2594,N_2556,N_2529);
and U2595 (N_2595,N_2577,N_2565);
or U2596 (N_2596,N_2571,N_2562);
nor U2597 (N_2597,N_2522,N_2545);
xnor U2598 (N_2598,N_2539,N_2535);
nor U2599 (N_2599,N_2553,N_2573);
nand U2600 (N_2600,N_2533,N_2550);
nand U2601 (N_2601,N_2543,N_2540);
nor U2602 (N_2602,N_2564,N_2567);
and U2603 (N_2603,N_2551,N_2578);
and U2604 (N_2604,N_2527,N_2530);
or U2605 (N_2605,N_2525,N_2554);
nor U2606 (N_2606,N_2523,N_2560);
or U2607 (N_2607,N_2538,N_2537);
nor U2608 (N_2608,N_2532,N_2536);
nor U2609 (N_2609,N_2548,N_2568);
nor U2610 (N_2610,N_2553,N_2527);
and U2611 (N_2611,N_2554,N_2565);
nor U2612 (N_2612,N_2559,N_2537);
or U2613 (N_2613,N_2530,N_2569);
nor U2614 (N_2614,N_2576,N_2551);
nor U2615 (N_2615,N_2542,N_2547);
or U2616 (N_2616,N_2522,N_2559);
and U2617 (N_2617,N_2570,N_2520);
nand U2618 (N_2618,N_2572,N_2529);
nand U2619 (N_2619,N_2549,N_2577);
and U2620 (N_2620,N_2522,N_2557);
and U2621 (N_2621,N_2565,N_2557);
and U2622 (N_2622,N_2566,N_2538);
nor U2623 (N_2623,N_2568,N_2579);
and U2624 (N_2624,N_2546,N_2570);
nor U2625 (N_2625,N_2540,N_2520);
or U2626 (N_2626,N_2562,N_2529);
or U2627 (N_2627,N_2521,N_2576);
nand U2628 (N_2628,N_2545,N_2576);
xnor U2629 (N_2629,N_2566,N_2567);
nand U2630 (N_2630,N_2543,N_2549);
or U2631 (N_2631,N_2546,N_2549);
and U2632 (N_2632,N_2553,N_2521);
or U2633 (N_2633,N_2575,N_2556);
and U2634 (N_2634,N_2562,N_2534);
or U2635 (N_2635,N_2533,N_2535);
nand U2636 (N_2636,N_2554,N_2576);
or U2637 (N_2637,N_2574,N_2577);
nand U2638 (N_2638,N_2540,N_2546);
or U2639 (N_2639,N_2532,N_2546);
nor U2640 (N_2640,N_2592,N_2639);
nor U2641 (N_2641,N_2616,N_2617);
or U2642 (N_2642,N_2589,N_2590);
and U2643 (N_2643,N_2634,N_2636);
nand U2644 (N_2644,N_2600,N_2614);
or U2645 (N_2645,N_2620,N_2587);
and U2646 (N_2646,N_2618,N_2612);
or U2647 (N_2647,N_2597,N_2591);
nor U2648 (N_2648,N_2601,N_2585);
and U2649 (N_2649,N_2588,N_2622);
and U2650 (N_2650,N_2631,N_2594);
nor U2651 (N_2651,N_2596,N_2629);
nor U2652 (N_2652,N_2627,N_2637);
and U2653 (N_2653,N_2638,N_2609);
or U2654 (N_2654,N_2632,N_2595);
xnor U2655 (N_2655,N_2605,N_2586);
and U2656 (N_2656,N_2608,N_2611);
nor U2657 (N_2657,N_2624,N_2621);
or U2658 (N_2658,N_2603,N_2613);
nor U2659 (N_2659,N_2580,N_2610);
nor U2660 (N_2660,N_2623,N_2606);
or U2661 (N_2661,N_2607,N_2615);
or U2662 (N_2662,N_2602,N_2619);
nand U2663 (N_2663,N_2599,N_2581);
or U2664 (N_2664,N_2635,N_2582);
and U2665 (N_2665,N_2604,N_2625);
xnor U2666 (N_2666,N_2633,N_2628);
xor U2667 (N_2667,N_2630,N_2583);
or U2668 (N_2668,N_2593,N_2626);
or U2669 (N_2669,N_2584,N_2598);
or U2670 (N_2670,N_2599,N_2638);
nand U2671 (N_2671,N_2620,N_2599);
nor U2672 (N_2672,N_2586,N_2607);
nand U2673 (N_2673,N_2624,N_2627);
nand U2674 (N_2674,N_2616,N_2584);
or U2675 (N_2675,N_2583,N_2587);
or U2676 (N_2676,N_2596,N_2608);
xor U2677 (N_2677,N_2583,N_2636);
and U2678 (N_2678,N_2628,N_2622);
nand U2679 (N_2679,N_2602,N_2592);
nor U2680 (N_2680,N_2613,N_2581);
and U2681 (N_2681,N_2632,N_2615);
nand U2682 (N_2682,N_2628,N_2585);
nor U2683 (N_2683,N_2620,N_2616);
nand U2684 (N_2684,N_2636,N_2638);
xnor U2685 (N_2685,N_2617,N_2591);
or U2686 (N_2686,N_2594,N_2601);
nand U2687 (N_2687,N_2636,N_2629);
nor U2688 (N_2688,N_2623,N_2584);
xnor U2689 (N_2689,N_2583,N_2614);
xnor U2690 (N_2690,N_2592,N_2635);
nor U2691 (N_2691,N_2581,N_2624);
nor U2692 (N_2692,N_2607,N_2581);
nand U2693 (N_2693,N_2599,N_2589);
nor U2694 (N_2694,N_2591,N_2615);
and U2695 (N_2695,N_2611,N_2632);
xnor U2696 (N_2696,N_2590,N_2600);
nand U2697 (N_2697,N_2619,N_2584);
or U2698 (N_2698,N_2592,N_2597);
nor U2699 (N_2699,N_2603,N_2630);
xnor U2700 (N_2700,N_2669,N_2695);
nor U2701 (N_2701,N_2654,N_2681);
and U2702 (N_2702,N_2655,N_2668);
or U2703 (N_2703,N_2696,N_2658);
nand U2704 (N_2704,N_2667,N_2640);
nor U2705 (N_2705,N_2652,N_2680);
or U2706 (N_2706,N_2694,N_2697);
or U2707 (N_2707,N_2648,N_2671);
xor U2708 (N_2708,N_2683,N_2674);
and U2709 (N_2709,N_2688,N_2699);
and U2710 (N_2710,N_2686,N_2644);
and U2711 (N_2711,N_2656,N_2650);
or U2712 (N_2712,N_2645,N_2692);
nand U2713 (N_2713,N_2685,N_2643);
and U2714 (N_2714,N_2641,N_2647);
nand U2715 (N_2715,N_2677,N_2684);
nand U2716 (N_2716,N_2657,N_2642);
xnor U2717 (N_2717,N_2698,N_2653);
and U2718 (N_2718,N_2664,N_2663);
and U2719 (N_2719,N_2678,N_2676);
nor U2720 (N_2720,N_2675,N_2693);
or U2721 (N_2721,N_2646,N_2682);
or U2722 (N_2722,N_2649,N_2691);
or U2723 (N_2723,N_2662,N_2666);
and U2724 (N_2724,N_2672,N_2687);
nand U2725 (N_2725,N_2690,N_2670);
or U2726 (N_2726,N_2661,N_2673);
and U2727 (N_2727,N_2660,N_2689);
nor U2728 (N_2728,N_2665,N_2651);
and U2729 (N_2729,N_2679,N_2659);
and U2730 (N_2730,N_2698,N_2688);
nor U2731 (N_2731,N_2688,N_2669);
nand U2732 (N_2732,N_2696,N_2669);
and U2733 (N_2733,N_2697,N_2657);
or U2734 (N_2734,N_2690,N_2647);
nor U2735 (N_2735,N_2677,N_2680);
nand U2736 (N_2736,N_2656,N_2671);
xnor U2737 (N_2737,N_2658,N_2677);
or U2738 (N_2738,N_2689,N_2667);
nor U2739 (N_2739,N_2667,N_2644);
nor U2740 (N_2740,N_2646,N_2681);
nand U2741 (N_2741,N_2667,N_2649);
and U2742 (N_2742,N_2640,N_2674);
nand U2743 (N_2743,N_2684,N_2694);
nand U2744 (N_2744,N_2668,N_2660);
nor U2745 (N_2745,N_2670,N_2655);
nand U2746 (N_2746,N_2654,N_2668);
nor U2747 (N_2747,N_2640,N_2692);
nor U2748 (N_2748,N_2652,N_2645);
or U2749 (N_2749,N_2674,N_2653);
and U2750 (N_2750,N_2689,N_2694);
nor U2751 (N_2751,N_2665,N_2649);
nand U2752 (N_2752,N_2671,N_2698);
nor U2753 (N_2753,N_2647,N_2685);
nor U2754 (N_2754,N_2645,N_2670);
xnor U2755 (N_2755,N_2686,N_2687);
nand U2756 (N_2756,N_2687,N_2657);
and U2757 (N_2757,N_2664,N_2654);
and U2758 (N_2758,N_2687,N_2668);
or U2759 (N_2759,N_2667,N_2670);
xnor U2760 (N_2760,N_2726,N_2721);
or U2761 (N_2761,N_2719,N_2744);
xor U2762 (N_2762,N_2739,N_2701);
and U2763 (N_2763,N_2731,N_2732);
or U2764 (N_2764,N_2705,N_2710);
or U2765 (N_2765,N_2741,N_2704);
nor U2766 (N_2766,N_2722,N_2750);
xor U2767 (N_2767,N_2708,N_2700);
nand U2768 (N_2768,N_2725,N_2755);
or U2769 (N_2769,N_2733,N_2734);
nand U2770 (N_2770,N_2757,N_2728);
and U2771 (N_2771,N_2743,N_2735);
nand U2772 (N_2772,N_2753,N_2707);
or U2773 (N_2773,N_2752,N_2715);
nand U2774 (N_2774,N_2723,N_2759);
nor U2775 (N_2775,N_2730,N_2709);
nand U2776 (N_2776,N_2716,N_2751);
or U2777 (N_2777,N_2706,N_2711);
and U2778 (N_2778,N_2714,N_2712);
and U2779 (N_2779,N_2748,N_2724);
and U2780 (N_2780,N_2729,N_2737);
nand U2781 (N_2781,N_2717,N_2742);
or U2782 (N_2782,N_2727,N_2756);
nor U2783 (N_2783,N_2749,N_2736);
xor U2784 (N_2784,N_2745,N_2718);
and U2785 (N_2785,N_2720,N_2702);
xnor U2786 (N_2786,N_2754,N_2747);
nor U2787 (N_2787,N_2738,N_2740);
or U2788 (N_2788,N_2713,N_2703);
nor U2789 (N_2789,N_2746,N_2758);
xnor U2790 (N_2790,N_2743,N_2732);
or U2791 (N_2791,N_2753,N_2747);
and U2792 (N_2792,N_2749,N_2705);
or U2793 (N_2793,N_2710,N_2700);
and U2794 (N_2794,N_2705,N_2719);
nand U2795 (N_2795,N_2731,N_2726);
nor U2796 (N_2796,N_2753,N_2728);
and U2797 (N_2797,N_2723,N_2725);
xnor U2798 (N_2798,N_2739,N_2709);
nand U2799 (N_2799,N_2709,N_2710);
nand U2800 (N_2800,N_2723,N_2718);
or U2801 (N_2801,N_2729,N_2743);
and U2802 (N_2802,N_2747,N_2739);
or U2803 (N_2803,N_2759,N_2745);
nor U2804 (N_2804,N_2748,N_2757);
or U2805 (N_2805,N_2720,N_2744);
nor U2806 (N_2806,N_2750,N_2705);
or U2807 (N_2807,N_2730,N_2701);
and U2808 (N_2808,N_2724,N_2736);
nor U2809 (N_2809,N_2752,N_2749);
or U2810 (N_2810,N_2705,N_2701);
nand U2811 (N_2811,N_2728,N_2743);
xnor U2812 (N_2812,N_2710,N_2707);
nand U2813 (N_2813,N_2754,N_2739);
xnor U2814 (N_2814,N_2743,N_2725);
nand U2815 (N_2815,N_2727,N_2742);
or U2816 (N_2816,N_2742,N_2738);
or U2817 (N_2817,N_2736,N_2750);
and U2818 (N_2818,N_2734,N_2746);
and U2819 (N_2819,N_2717,N_2752);
nand U2820 (N_2820,N_2774,N_2767);
nor U2821 (N_2821,N_2809,N_2771);
or U2822 (N_2822,N_2764,N_2816);
xnor U2823 (N_2823,N_2787,N_2795);
or U2824 (N_2824,N_2766,N_2761);
and U2825 (N_2825,N_2812,N_2768);
xor U2826 (N_2826,N_2817,N_2813);
nor U2827 (N_2827,N_2807,N_2796);
nor U2828 (N_2828,N_2784,N_2804);
nand U2829 (N_2829,N_2793,N_2762);
and U2830 (N_2830,N_2806,N_2785);
nor U2831 (N_2831,N_2786,N_2776);
nor U2832 (N_2832,N_2808,N_2781);
nand U2833 (N_2833,N_2798,N_2783);
or U2834 (N_2834,N_2775,N_2770);
nand U2835 (N_2835,N_2769,N_2803);
or U2836 (N_2836,N_2811,N_2779);
nand U2837 (N_2837,N_2791,N_2763);
or U2838 (N_2838,N_2818,N_2801);
or U2839 (N_2839,N_2789,N_2815);
nor U2840 (N_2840,N_2782,N_2810);
nand U2841 (N_2841,N_2788,N_2765);
and U2842 (N_2842,N_2802,N_2792);
nand U2843 (N_2843,N_2814,N_2777);
or U2844 (N_2844,N_2819,N_2778);
and U2845 (N_2845,N_2805,N_2760);
nor U2846 (N_2846,N_2799,N_2800);
nand U2847 (N_2847,N_2794,N_2790);
and U2848 (N_2848,N_2780,N_2773);
nor U2849 (N_2849,N_2797,N_2772);
xnor U2850 (N_2850,N_2794,N_2813);
nand U2851 (N_2851,N_2795,N_2810);
nor U2852 (N_2852,N_2816,N_2800);
nor U2853 (N_2853,N_2765,N_2809);
nor U2854 (N_2854,N_2777,N_2798);
and U2855 (N_2855,N_2772,N_2815);
nand U2856 (N_2856,N_2808,N_2799);
or U2857 (N_2857,N_2813,N_2811);
or U2858 (N_2858,N_2762,N_2784);
nand U2859 (N_2859,N_2768,N_2791);
and U2860 (N_2860,N_2770,N_2806);
nand U2861 (N_2861,N_2774,N_2815);
and U2862 (N_2862,N_2802,N_2800);
and U2863 (N_2863,N_2807,N_2798);
and U2864 (N_2864,N_2789,N_2808);
xnor U2865 (N_2865,N_2775,N_2818);
or U2866 (N_2866,N_2796,N_2794);
and U2867 (N_2867,N_2813,N_2772);
and U2868 (N_2868,N_2774,N_2801);
xor U2869 (N_2869,N_2799,N_2774);
nand U2870 (N_2870,N_2760,N_2809);
xnor U2871 (N_2871,N_2794,N_2805);
and U2872 (N_2872,N_2805,N_2780);
nand U2873 (N_2873,N_2771,N_2778);
or U2874 (N_2874,N_2781,N_2806);
nor U2875 (N_2875,N_2817,N_2773);
or U2876 (N_2876,N_2802,N_2782);
and U2877 (N_2877,N_2815,N_2800);
or U2878 (N_2878,N_2773,N_2815);
nor U2879 (N_2879,N_2760,N_2775);
nor U2880 (N_2880,N_2844,N_2836);
xnor U2881 (N_2881,N_2831,N_2842);
nand U2882 (N_2882,N_2853,N_2868);
nand U2883 (N_2883,N_2854,N_2837);
xor U2884 (N_2884,N_2845,N_2835);
or U2885 (N_2885,N_2848,N_2823);
or U2886 (N_2886,N_2828,N_2850);
and U2887 (N_2887,N_2822,N_2866);
or U2888 (N_2888,N_2861,N_2855);
nor U2889 (N_2889,N_2852,N_2865);
nor U2890 (N_2890,N_2846,N_2871);
or U2891 (N_2891,N_2873,N_2840);
and U2892 (N_2892,N_2847,N_2841);
and U2893 (N_2893,N_2851,N_2870);
or U2894 (N_2894,N_2877,N_2872);
nor U2895 (N_2895,N_2856,N_2833);
nor U2896 (N_2896,N_2839,N_2875);
nand U2897 (N_2897,N_2869,N_2838);
xor U2898 (N_2898,N_2830,N_2879);
nor U2899 (N_2899,N_2826,N_2874);
or U2900 (N_2900,N_2867,N_2860);
nor U2901 (N_2901,N_2849,N_2863);
and U2902 (N_2902,N_2862,N_2827);
nor U2903 (N_2903,N_2820,N_2857);
nand U2904 (N_2904,N_2821,N_2829);
or U2905 (N_2905,N_2859,N_2858);
nand U2906 (N_2906,N_2843,N_2825);
or U2907 (N_2907,N_2834,N_2876);
nor U2908 (N_2908,N_2864,N_2824);
and U2909 (N_2909,N_2878,N_2832);
nor U2910 (N_2910,N_2854,N_2871);
nand U2911 (N_2911,N_2855,N_2847);
and U2912 (N_2912,N_2850,N_2824);
and U2913 (N_2913,N_2873,N_2831);
or U2914 (N_2914,N_2840,N_2857);
xnor U2915 (N_2915,N_2855,N_2858);
nor U2916 (N_2916,N_2828,N_2825);
and U2917 (N_2917,N_2845,N_2834);
nand U2918 (N_2918,N_2865,N_2873);
xnor U2919 (N_2919,N_2872,N_2832);
nor U2920 (N_2920,N_2854,N_2855);
or U2921 (N_2921,N_2877,N_2879);
nand U2922 (N_2922,N_2879,N_2872);
nand U2923 (N_2923,N_2842,N_2821);
nor U2924 (N_2924,N_2847,N_2823);
xnor U2925 (N_2925,N_2839,N_2847);
nor U2926 (N_2926,N_2866,N_2841);
nand U2927 (N_2927,N_2860,N_2854);
nor U2928 (N_2928,N_2845,N_2849);
or U2929 (N_2929,N_2826,N_2824);
nor U2930 (N_2930,N_2834,N_2839);
xor U2931 (N_2931,N_2842,N_2859);
nand U2932 (N_2932,N_2867,N_2849);
and U2933 (N_2933,N_2825,N_2858);
and U2934 (N_2934,N_2853,N_2822);
nand U2935 (N_2935,N_2877,N_2820);
or U2936 (N_2936,N_2855,N_2829);
xnor U2937 (N_2937,N_2829,N_2846);
or U2938 (N_2938,N_2831,N_2851);
nor U2939 (N_2939,N_2866,N_2827);
nor U2940 (N_2940,N_2922,N_2925);
nand U2941 (N_2941,N_2912,N_2932);
and U2942 (N_2942,N_2899,N_2903);
and U2943 (N_2943,N_2896,N_2885);
nand U2944 (N_2944,N_2881,N_2937);
and U2945 (N_2945,N_2935,N_2898);
and U2946 (N_2946,N_2904,N_2920);
and U2947 (N_2947,N_2929,N_2934);
nor U2948 (N_2948,N_2907,N_2921);
or U2949 (N_2949,N_2918,N_2897);
and U2950 (N_2950,N_2926,N_2916);
nand U2951 (N_2951,N_2880,N_2882);
or U2952 (N_2952,N_2906,N_2917);
nor U2953 (N_2953,N_2939,N_2887);
nand U2954 (N_2954,N_2893,N_2886);
nor U2955 (N_2955,N_2890,N_2883);
and U2956 (N_2956,N_2900,N_2914);
and U2957 (N_2957,N_2938,N_2888);
or U2958 (N_2958,N_2902,N_2884);
nand U2959 (N_2959,N_2909,N_2895);
or U2960 (N_2960,N_2931,N_2933);
nor U2961 (N_2961,N_2915,N_2913);
or U2962 (N_2962,N_2930,N_2927);
nand U2963 (N_2963,N_2911,N_2924);
xor U2964 (N_2964,N_2908,N_2936);
and U2965 (N_2965,N_2923,N_2891);
nand U2966 (N_2966,N_2928,N_2894);
nor U2967 (N_2967,N_2892,N_2889);
nor U2968 (N_2968,N_2910,N_2905);
nor U2969 (N_2969,N_2901,N_2919);
and U2970 (N_2970,N_2909,N_2935);
and U2971 (N_2971,N_2934,N_2914);
or U2972 (N_2972,N_2894,N_2936);
nand U2973 (N_2973,N_2895,N_2936);
nor U2974 (N_2974,N_2931,N_2881);
and U2975 (N_2975,N_2908,N_2911);
xnor U2976 (N_2976,N_2928,N_2932);
or U2977 (N_2977,N_2893,N_2925);
xor U2978 (N_2978,N_2905,N_2932);
nor U2979 (N_2979,N_2890,N_2915);
nand U2980 (N_2980,N_2939,N_2907);
or U2981 (N_2981,N_2928,N_2938);
nand U2982 (N_2982,N_2900,N_2924);
nor U2983 (N_2983,N_2884,N_2908);
nand U2984 (N_2984,N_2885,N_2898);
and U2985 (N_2985,N_2937,N_2930);
and U2986 (N_2986,N_2938,N_2893);
nand U2987 (N_2987,N_2889,N_2939);
and U2988 (N_2988,N_2930,N_2883);
and U2989 (N_2989,N_2923,N_2897);
or U2990 (N_2990,N_2924,N_2936);
and U2991 (N_2991,N_2889,N_2907);
nand U2992 (N_2992,N_2888,N_2925);
nand U2993 (N_2993,N_2886,N_2938);
or U2994 (N_2994,N_2889,N_2912);
or U2995 (N_2995,N_2883,N_2901);
xnor U2996 (N_2996,N_2898,N_2919);
nor U2997 (N_2997,N_2934,N_2921);
or U2998 (N_2998,N_2881,N_2903);
nor U2999 (N_2999,N_2900,N_2919);
nand UO_0 (O_0,N_2964,N_2970);
and UO_1 (O_1,N_2981,N_2998);
nor UO_2 (O_2,N_2950,N_2948);
and UO_3 (O_3,N_2972,N_2968);
or UO_4 (O_4,N_2952,N_2973);
nand UO_5 (O_5,N_2945,N_2965);
xor UO_6 (O_6,N_2963,N_2986);
nor UO_7 (O_7,N_2991,N_2956);
or UO_8 (O_8,N_2955,N_2940);
and UO_9 (O_9,N_2947,N_2957);
nor UO_10 (O_10,N_2975,N_2960);
or UO_11 (O_11,N_2983,N_2978);
nand UO_12 (O_12,N_2989,N_2946);
nor UO_13 (O_13,N_2996,N_2942);
nand UO_14 (O_14,N_2992,N_2999);
xnor UO_15 (O_15,N_2969,N_2990);
nor UO_16 (O_16,N_2997,N_2984);
nor UO_17 (O_17,N_2994,N_2987);
or UO_18 (O_18,N_2982,N_2954);
or UO_19 (O_19,N_2959,N_2943);
nor UO_20 (O_20,N_2941,N_2951);
nand UO_21 (O_21,N_2988,N_2961);
nand UO_22 (O_22,N_2985,N_2977);
nand UO_23 (O_23,N_2967,N_2958);
nand UO_24 (O_24,N_2976,N_2949);
or UO_25 (O_25,N_2993,N_2953);
or UO_26 (O_26,N_2944,N_2980);
nor UO_27 (O_27,N_2962,N_2979);
xor UO_28 (O_28,N_2974,N_2995);
nor UO_29 (O_29,N_2966,N_2971);
nor UO_30 (O_30,N_2987,N_2978);
nor UO_31 (O_31,N_2974,N_2955);
nand UO_32 (O_32,N_2947,N_2958);
nand UO_33 (O_33,N_2980,N_2999);
nor UO_34 (O_34,N_2958,N_2945);
or UO_35 (O_35,N_2996,N_2998);
nand UO_36 (O_36,N_2955,N_2947);
and UO_37 (O_37,N_2943,N_2978);
and UO_38 (O_38,N_2941,N_2999);
nand UO_39 (O_39,N_2970,N_2962);
or UO_40 (O_40,N_2953,N_2983);
nand UO_41 (O_41,N_2942,N_2964);
and UO_42 (O_42,N_2947,N_2997);
or UO_43 (O_43,N_2991,N_2965);
or UO_44 (O_44,N_2972,N_2962);
nor UO_45 (O_45,N_2958,N_2952);
nand UO_46 (O_46,N_2990,N_2986);
and UO_47 (O_47,N_2953,N_2942);
nand UO_48 (O_48,N_2976,N_2940);
xnor UO_49 (O_49,N_2978,N_2974);
nor UO_50 (O_50,N_2974,N_2998);
and UO_51 (O_51,N_2996,N_2979);
nand UO_52 (O_52,N_2954,N_2977);
nor UO_53 (O_53,N_2985,N_2988);
xor UO_54 (O_54,N_2997,N_2983);
or UO_55 (O_55,N_2979,N_2958);
or UO_56 (O_56,N_2958,N_2956);
and UO_57 (O_57,N_2960,N_2995);
or UO_58 (O_58,N_2988,N_2975);
xor UO_59 (O_59,N_2976,N_2945);
or UO_60 (O_60,N_2942,N_2944);
and UO_61 (O_61,N_2995,N_2952);
nand UO_62 (O_62,N_2946,N_2958);
xor UO_63 (O_63,N_2941,N_2953);
and UO_64 (O_64,N_2987,N_2997);
or UO_65 (O_65,N_2986,N_2987);
nor UO_66 (O_66,N_2976,N_2978);
and UO_67 (O_67,N_2957,N_2964);
and UO_68 (O_68,N_2943,N_2968);
and UO_69 (O_69,N_2979,N_2982);
nor UO_70 (O_70,N_2940,N_2999);
xor UO_71 (O_71,N_2973,N_2981);
and UO_72 (O_72,N_2952,N_2941);
or UO_73 (O_73,N_2994,N_2951);
or UO_74 (O_74,N_2975,N_2955);
or UO_75 (O_75,N_2991,N_2977);
xor UO_76 (O_76,N_2997,N_2968);
or UO_77 (O_77,N_2954,N_2992);
and UO_78 (O_78,N_2945,N_2974);
or UO_79 (O_79,N_2975,N_2964);
nand UO_80 (O_80,N_2966,N_2996);
or UO_81 (O_81,N_2987,N_2953);
nor UO_82 (O_82,N_2974,N_2976);
or UO_83 (O_83,N_2941,N_2971);
and UO_84 (O_84,N_2943,N_2940);
nor UO_85 (O_85,N_2968,N_2994);
and UO_86 (O_86,N_2940,N_2945);
or UO_87 (O_87,N_2946,N_2969);
nand UO_88 (O_88,N_2990,N_2951);
and UO_89 (O_89,N_2951,N_2970);
or UO_90 (O_90,N_2981,N_2982);
xor UO_91 (O_91,N_2959,N_2993);
and UO_92 (O_92,N_2972,N_2985);
and UO_93 (O_93,N_2988,N_2940);
nand UO_94 (O_94,N_2962,N_2941);
or UO_95 (O_95,N_2958,N_2961);
nand UO_96 (O_96,N_2975,N_2947);
nor UO_97 (O_97,N_2971,N_2973);
xnor UO_98 (O_98,N_2954,N_2966);
and UO_99 (O_99,N_2981,N_2945);
and UO_100 (O_100,N_2968,N_2971);
or UO_101 (O_101,N_2998,N_2952);
nor UO_102 (O_102,N_2944,N_2951);
and UO_103 (O_103,N_2966,N_2941);
and UO_104 (O_104,N_2972,N_2996);
and UO_105 (O_105,N_2946,N_2980);
or UO_106 (O_106,N_2964,N_2952);
nor UO_107 (O_107,N_2943,N_2962);
xnor UO_108 (O_108,N_2945,N_2956);
or UO_109 (O_109,N_2972,N_2941);
and UO_110 (O_110,N_2985,N_2989);
or UO_111 (O_111,N_2996,N_2987);
nor UO_112 (O_112,N_2998,N_2945);
or UO_113 (O_113,N_2990,N_2988);
nand UO_114 (O_114,N_2990,N_2976);
or UO_115 (O_115,N_2965,N_2961);
or UO_116 (O_116,N_2949,N_2960);
xor UO_117 (O_117,N_2995,N_2977);
nor UO_118 (O_118,N_2993,N_2971);
or UO_119 (O_119,N_2952,N_2984);
xor UO_120 (O_120,N_2999,N_2983);
nand UO_121 (O_121,N_2965,N_2953);
nand UO_122 (O_122,N_2997,N_2960);
nor UO_123 (O_123,N_2983,N_2971);
or UO_124 (O_124,N_2993,N_2982);
nor UO_125 (O_125,N_2953,N_2991);
nor UO_126 (O_126,N_2974,N_2988);
nand UO_127 (O_127,N_2948,N_2949);
nand UO_128 (O_128,N_2970,N_2982);
or UO_129 (O_129,N_2968,N_2969);
and UO_130 (O_130,N_2989,N_2982);
or UO_131 (O_131,N_2958,N_2988);
nand UO_132 (O_132,N_2964,N_2988);
or UO_133 (O_133,N_2966,N_2957);
xor UO_134 (O_134,N_2990,N_2994);
xor UO_135 (O_135,N_2941,N_2963);
or UO_136 (O_136,N_2986,N_2975);
and UO_137 (O_137,N_2962,N_2977);
or UO_138 (O_138,N_2948,N_2958);
and UO_139 (O_139,N_2975,N_2942);
nor UO_140 (O_140,N_2972,N_2953);
or UO_141 (O_141,N_2992,N_2990);
or UO_142 (O_142,N_2961,N_2967);
nand UO_143 (O_143,N_2987,N_2955);
xnor UO_144 (O_144,N_2994,N_2972);
and UO_145 (O_145,N_2944,N_2983);
xnor UO_146 (O_146,N_2964,N_2951);
and UO_147 (O_147,N_2981,N_2944);
or UO_148 (O_148,N_2956,N_2993);
xor UO_149 (O_149,N_2945,N_2983);
nand UO_150 (O_150,N_2946,N_2949);
xnor UO_151 (O_151,N_2988,N_2962);
and UO_152 (O_152,N_2989,N_2963);
or UO_153 (O_153,N_2993,N_2979);
nor UO_154 (O_154,N_2978,N_2991);
nor UO_155 (O_155,N_2949,N_2975);
nand UO_156 (O_156,N_2988,N_2973);
nor UO_157 (O_157,N_2995,N_2967);
and UO_158 (O_158,N_2976,N_2959);
or UO_159 (O_159,N_2960,N_2964);
nor UO_160 (O_160,N_2979,N_2952);
nor UO_161 (O_161,N_2976,N_2981);
and UO_162 (O_162,N_2983,N_2994);
and UO_163 (O_163,N_2961,N_2981);
nor UO_164 (O_164,N_2945,N_2960);
nand UO_165 (O_165,N_2980,N_2949);
nor UO_166 (O_166,N_2960,N_2951);
and UO_167 (O_167,N_2980,N_2995);
nor UO_168 (O_168,N_2995,N_2976);
nand UO_169 (O_169,N_2998,N_2967);
or UO_170 (O_170,N_2984,N_2995);
nand UO_171 (O_171,N_2951,N_2975);
or UO_172 (O_172,N_2986,N_2992);
and UO_173 (O_173,N_2951,N_2969);
nor UO_174 (O_174,N_2946,N_2979);
nor UO_175 (O_175,N_2976,N_2948);
or UO_176 (O_176,N_2979,N_2971);
and UO_177 (O_177,N_2949,N_2958);
nor UO_178 (O_178,N_2968,N_2973);
and UO_179 (O_179,N_2946,N_2951);
nand UO_180 (O_180,N_2998,N_2976);
nand UO_181 (O_181,N_2979,N_2978);
and UO_182 (O_182,N_2946,N_2950);
or UO_183 (O_183,N_2967,N_2973);
or UO_184 (O_184,N_2989,N_2940);
nand UO_185 (O_185,N_2995,N_2953);
nor UO_186 (O_186,N_2977,N_2970);
and UO_187 (O_187,N_2974,N_2972);
and UO_188 (O_188,N_2998,N_2978);
and UO_189 (O_189,N_2975,N_2965);
nand UO_190 (O_190,N_2975,N_2953);
and UO_191 (O_191,N_2973,N_2976);
and UO_192 (O_192,N_2962,N_2993);
nor UO_193 (O_193,N_2994,N_2960);
and UO_194 (O_194,N_2974,N_2990);
nand UO_195 (O_195,N_2940,N_2968);
or UO_196 (O_196,N_2957,N_2996);
and UO_197 (O_197,N_2967,N_2993);
nor UO_198 (O_198,N_2997,N_2993);
nand UO_199 (O_199,N_2976,N_2954);
or UO_200 (O_200,N_2971,N_2975);
nand UO_201 (O_201,N_2983,N_2989);
or UO_202 (O_202,N_2950,N_2989);
or UO_203 (O_203,N_2990,N_2942);
xor UO_204 (O_204,N_2992,N_2959);
nand UO_205 (O_205,N_2990,N_2947);
or UO_206 (O_206,N_2956,N_2979);
xor UO_207 (O_207,N_2951,N_2973);
nor UO_208 (O_208,N_2955,N_2971);
or UO_209 (O_209,N_2968,N_2957);
nand UO_210 (O_210,N_2955,N_2992);
and UO_211 (O_211,N_2959,N_2980);
nor UO_212 (O_212,N_2963,N_2960);
or UO_213 (O_213,N_2953,N_2943);
nand UO_214 (O_214,N_2983,N_2987);
nor UO_215 (O_215,N_2969,N_2950);
or UO_216 (O_216,N_2957,N_2940);
xor UO_217 (O_217,N_2965,N_2984);
nor UO_218 (O_218,N_2984,N_2940);
nor UO_219 (O_219,N_2950,N_2992);
nor UO_220 (O_220,N_2976,N_2999);
xnor UO_221 (O_221,N_2981,N_2948);
or UO_222 (O_222,N_2968,N_2995);
or UO_223 (O_223,N_2970,N_2976);
nand UO_224 (O_224,N_2947,N_2948);
or UO_225 (O_225,N_2969,N_2964);
nand UO_226 (O_226,N_2962,N_2999);
nor UO_227 (O_227,N_2993,N_2963);
and UO_228 (O_228,N_2964,N_2999);
or UO_229 (O_229,N_2959,N_2979);
xnor UO_230 (O_230,N_2972,N_2979);
and UO_231 (O_231,N_2990,N_2978);
and UO_232 (O_232,N_2997,N_2954);
nand UO_233 (O_233,N_2947,N_2984);
or UO_234 (O_234,N_2992,N_2949);
nor UO_235 (O_235,N_2950,N_2952);
and UO_236 (O_236,N_2985,N_2996);
and UO_237 (O_237,N_2976,N_2980);
nand UO_238 (O_238,N_2961,N_2980);
and UO_239 (O_239,N_2953,N_2977);
and UO_240 (O_240,N_2994,N_2996);
or UO_241 (O_241,N_2982,N_2974);
and UO_242 (O_242,N_2968,N_2962);
or UO_243 (O_243,N_2943,N_2980);
nor UO_244 (O_244,N_2977,N_2966);
and UO_245 (O_245,N_2961,N_2971);
nor UO_246 (O_246,N_2981,N_2952);
nand UO_247 (O_247,N_2997,N_2971);
or UO_248 (O_248,N_2977,N_2982);
and UO_249 (O_249,N_2968,N_2953);
nor UO_250 (O_250,N_2953,N_2951);
and UO_251 (O_251,N_2990,N_2982);
and UO_252 (O_252,N_2949,N_2950);
nor UO_253 (O_253,N_2946,N_2960);
nor UO_254 (O_254,N_2954,N_2958);
nand UO_255 (O_255,N_2993,N_2966);
nor UO_256 (O_256,N_2942,N_2994);
nand UO_257 (O_257,N_2953,N_2960);
or UO_258 (O_258,N_2987,N_2992);
nor UO_259 (O_259,N_2951,N_2963);
and UO_260 (O_260,N_2940,N_2951);
nand UO_261 (O_261,N_2974,N_2999);
nand UO_262 (O_262,N_2945,N_2979);
nor UO_263 (O_263,N_2948,N_2957);
or UO_264 (O_264,N_2976,N_2966);
nor UO_265 (O_265,N_2982,N_2959);
xor UO_266 (O_266,N_2959,N_2994);
xnor UO_267 (O_267,N_2996,N_2995);
nand UO_268 (O_268,N_2998,N_2985);
nor UO_269 (O_269,N_2954,N_2955);
nand UO_270 (O_270,N_2975,N_2944);
nor UO_271 (O_271,N_2955,N_2943);
nand UO_272 (O_272,N_2945,N_2961);
nand UO_273 (O_273,N_2990,N_2996);
nor UO_274 (O_274,N_2967,N_2944);
or UO_275 (O_275,N_2965,N_2962);
nand UO_276 (O_276,N_2992,N_2953);
nor UO_277 (O_277,N_2967,N_2983);
nor UO_278 (O_278,N_2982,N_2980);
nor UO_279 (O_279,N_2978,N_2971);
and UO_280 (O_280,N_2942,N_2955);
nand UO_281 (O_281,N_2980,N_2955);
or UO_282 (O_282,N_2994,N_2949);
nand UO_283 (O_283,N_2940,N_2983);
nand UO_284 (O_284,N_2941,N_2994);
nand UO_285 (O_285,N_2995,N_2989);
nor UO_286 (O_286,N_2970,N_2991);
or UO_287 (O_287,N_2984,N_2975);
or UO_288 (O_288,N_2975,N_2948);
nand UO_289 (O_289,N_2960,N_2952);
nand UO_290 (O_290,N_2946,N_2977);
or UO_291 (O_291,N_2983,N_2976);
and UO_292 (O_292,N_2941,N_2996);
or UO_293 (O_293,N_2966,N_2963);
nand UO_294 (O_294,N_2999,N_2994);
nand UO_295 (O_295,N_2947,N_2972);
nor UO_296 (O_296,N_2962,N_2953);
or UO_297 (O_297,N_2949,N_2945);
and UO_298 (O_298,N_2985,N_2973);
or UO_299 (O_299,N_2999,N_2952);
nand UO_300 (O_300,N_2959,N_2970);
nor UO_301 (O_301,N_2995,N_2956);
nand UO_302 (O_302,N_2961,N_2942);
or UO_303 (O_303,N_2940,N_2944);
and UO_304 (O_304,N_2975,N_2962);
nand UO_305 (O_305,N_2956,N_2970);
and UO_306 (O_306,N_2985,N_2971);
nor UO_307 (O_307,N_2993,N_2985);
nand UO_308 (O_308,N_2987,N_2954);
and UO_309 (O_309,N_2956,N_2980);
or UO_310 (O_310,N_2966,N_2943);
nor UO_311 (O_311,N_2991,N_2948);
or UO_312 (O_312,N_2968,N_2951);
nor UO_313 (O_313,N_2941,N_2981);
nand UO_314 (O_314,N_2952,N_2985);
xnor UO_315 (O_315,N_2974,N_2991);
xnor UO_316 (O_316,N_2997,N_2988);
nand UO_317 (O_317,N_2971,N_2940);
or UO_318 (O_318,N_2954,N_2969);
nor UO_319 (O_319,N_2958,N_2998);
xor UO_320 (O_320,N_2965,N_2992);
or UO_321 (O_321,N_2968,N_2946);
nor UO_322 (O_322,N_2945,N_2978);
and UO_323 (O_323,N_2963,N_2994);
nand UO_324 (O_324,N_2998,N_2959);
nor UO_325 (O_325,N_2994,N_2986);
nand UO_326 (O_326,N_2995,N_2971);
nor UO_327 (O_327,N_2940,N_2973);
and UO_328 (O_328,N_2974,N_2979);
and UO_329 (O_329,N_2963,N_2984);
or UO_330 (O_330,N_2948,N_2997);
and UO_331 (O_331,N_2955,N_2998);
nor UO_332 (O_332,N_2996,N_2992);
xor UO_333 (O_333,N_2974,N_2953);
nand UO_334 (O_334,N_2989,N_2966);
or UO_335 (O_335,N_2964,N_2995);
nor UO_336 (O_336,N_2975,N_2978);
and UO_337 (O_337,N_2990,N_2964);
nor UO_338 (O_338,N_2955,N_2984);
and UO_339 (O_339,N_2968,N_2947);
or UO_340 (O_340,N_2948,N_2972);
nor UO_341 (O_341,N_2954,N_2945);
nand UO_342 (O_342,N_2972,N_2975);
or UO_343 (O_343,N_2986,N_2999);
nor UO_344 (O_344,N_2987,N_2944);
nor UO_345 (O_345,N_2975,N_2946);
nor UO_346 (O_346,N_2991,N_2987);
and UO_347 (O_347,N_2958,N_2957);
or UO_348 (O_348,N_2993,N_2952);
nor UO_349 (O_349,N_2995,N_2998);
and UO_350 (O_350,N_2950,N_2966);
and UO_351 (O_351,N_2951,N_2977);
nand UO_352 (O_352,N_2956,N_2981);
nand UO_353 (O_353,N_2996,N_2969);
or UO_354 (O_354,N_2979,N_2955);
and UO_355 (O_355,N_2976,N_2957);
nand UO_356 (O_356,N_2981,N_2977);
nand UO_357 (O_357,N_2969,N_2994);
nand UO_358 (O_358,N_2976,N_2968);
and UO_359 (O_359,N_2988,N_2999);
nor UO_360 (O_360,N_2944,N_2948);
xor UO_361 (O_361,N_2945,N_2941);
and UO_362 (O_362,N_2997,N_2965);
xor UO_363 (O_363,N_2984,N_2961);
and UO_364 (O_364,N_2990,N_2963);
and UO_365 (O_365,N_2960,N_2948);
and UO_366 (O_366,N_2963,N_2964);
nand UO_367 (O_367,N_2984,N_2979);
or UO_368 (O_368,N_2956,N_2971);
or UO_369 (O_369,N_2970,N_2945);
xnor UO_370 (O_370,N_2958,N_2986);
nor UO_371 (O_371,N_2965,N_2976);
nor UO_372 (O_372,N_2942,N_2960);
nand UO_373 (O_373,N_2995,N_2975);
nand UO_374 (O_374,N_2996,N_2945);
xor UO_375 (O_375,N_2988,N_2967);
and UO_376 (O_376,N_2960,N_2988);
nor UO_377 (O_377,N_2986,N_2993);
nand UO_378 (O_378,N_2949,N_2953);
and UO_379 (O_379,N_2996,N_2963);
nand UO_380 (O_380,N_2994,N_2943);
nor UO_381 (O_381,N_2942,N_2982);
and UO_382 (O_382,N_2940,N_2995);
and UO_383 (O_383,N_2958,N_2940);
or UO_384 (O_384,N_2954,N_2967);
nor UO_385 (O_385,N_2971,N_2981);
and UO_386 (O_386,N_2965,N_2968);
nor UO_387 (O_387,N_2975,N_2997);
and UO_388 (O_388,N_2984,N_2974);
and UO_389 (O_389,N_2940,N_2980);
nor UO_390 (O_390,N_2991,N_2951);
or UO_391 (O_391,N_2991,N_2968);
xor UO_392 (O_392,N_2981,N_2996);
nor UO_393 (O_393,N_2966,N_2997);
nand UO_394 (O_394,N_2946,N_2961);
nor UO_395 (O_395,N_2993,N_2964);
nor UO_396 (O_396,N_2957,N_2963);
nor UO_397 (O_397,N_2986,N_2976);
and UO_398 (O_398,N_2965,N_2964);
nor UO_399 (O_399,N_2964,N_2966);
xnor UO_400 (O_400,N_2947,N_2962);
nor UO_401 (O_401,N_2951,N_2947);
or UO_402 (O_402,N_2979,N_2949);
and UO_403 (O_403,N_2960,N_2956);
nor UO_404 (O_404,N_2980,N_2967);
nor UO_405 (O_405,N_2949,N_2977);
nor UO_406 (O_406,N_2987,N_2960);
nor UO_407 (O_407,N_2980,N_2947);
nor UO_408 (O_408,N_2952,N_2970);
nor UO_409 (O_409,N_2956,N_2944);
xnor UO_410 (O_410,N_2945,N_2967);
nand UO_411 (O_411,N_2967,N_2960);
nand UO_412 (O_412,N_2983,N_2958);
nand UO_413 (O_413,N_2968,N_2941);
nand UO_414 (O_414,N_2948,N_2999);
nand UO_415 (O_415,N_2963,N_2974);
or UO_416 (O_416,N_2962,N_2958);
nand UO_417 (O_417,N_2943,N_2961);
or UO_418 (O_418,N_2969,N_2952);
nor UO_419 (O_419,N_2957,N_2952);
nor UO_420 (O_420,N_2959,N_2957);
nor UO_421 (O_421,N_2969,N_2953);
and UO_422 (O_422,N_2979,N_2944);
and UO_423 (O_423,N_2990,N_2948);
nor UO_424 (O_424,N_2967,N_2953);
or UO_425 (O_425,N_2995,N_2992);
xnor UO_426 (O_426,N_2979,N_2986);
nand UO_427 (O_427,N_2943,N_2989);
nor UO_428 (O_428,N_2940,N_2992);
and UO_429 (O_429,N_2967,N_2984);
xnor UO_430 (O_430,N_2974,N_2944);
nor UO_431 (O_431,N_2990,N_2949);
or UO_432 (O_432,N_2953,N_2970);
and UO_433 (O_433,N_2948,N_2943);
or UO_434 (O_434,N_2979,N_2997);
or UO_435 (O_435,N_2967,N_2979);
xor UO_436 (O_436,N_2984,N_2957);
and UO_437 (O_437,N_2955,N_2969);
nor UO_438 (O_438,N_2992,N_2977);
xor UO_439 (O_439,N_2983,N_2951);
nor UO_440 (O_440,N_2974,N_2996);
or UO_441 (O_441,N_2955,N_2949);
nand UO_442 (O_442,N_2974,N_2942);
xor UO_443 (O_443,N_2975,N_2961);
and UO_444 (O_444,N_2996,N_2964);
nand UO_445 (O_445,N_2966,N_2968);
nand UO_446 (O_446,N_2955,N_2967);
xnor UO_447 (O_447,N_2962,N_2940);
nor UO_448 (O_448,N_2977,N_2983);
nor UO_449 (O_449,N_2957,N_2961);
or UO_450 (O_450,N_2957,N_2983);
and UO_451 (O_451,N_2983,N_2970);
and UO_452 (O_452,N_2969,N_2948);
and UO_453 (O_453,N_2942,N_2970);
or UO_454 (O_454,N_2951,N_2945);
nor UO_455 (O_455,N_2960,N_2989);
nand UO_456 (O_456,N_2942,N_2949);
or UO_457 (O_457,N_2950,N_2947);
nand UO_458 (O_458,N_2980,N_2997);
or UO_459 (O_459,N_2991,N_2984);
or UO_460 (O_460,N_2964,N_2974);
nand UO_461 (O_461,N_2991,N_2946);
xnor UO_462 (O_462,N_2986,N_2967);
nand UO_463 (O_463,N_2961,N_2972);
nand UO_464 (O_464,N_2969,N_2975);
or UO_465 (O_465,N_2985,N_2978);
nor UO_466 (O_466,N_2962,N_2961);
nand UO_467 (O_467,N_2988,N_2952);
and UO_468 (O_468,N_2997,N_2994);
nor UO_469 (O_469,N_2950,N_2980);
or UO_470 (O_470,N_2984,N_2988);
or UO_471 (O_471,N_2968,N_2950);
nor UO_472 (O_472,N_2973,N_2992);
and UO_473 (O_473,N_2959,N_2952);
or UO_474 (O_474,N_2997,N_2985);
or UO_475 (O_475,N_2970,N_2974);
or UO_476 (O_476,N_2950,N_2974);
nand UO_477 (O_477,N_2951,N_2950);
nor UO_478 (O_478,N_2991,N_2949);
nor UO_479 (O_479,N_2982,N_2971);
nor UO_480 (O_480,N_2950,N_2973);
or UO_481 (O_481,N_2996,N_2986);
nor UO_482 (O_482,N_2949,N_2987);
and UO_483 (O_483,N_2973,N_2999);
nand UO_484 (O_484,N_2945,N_2948);
nor UO_485 (O_485,N_2983,N_2959);
nand UO_486 (O_486,N_2943,N_2990);
and UO_487 (O_487,N_2972,N_2991);
and UO_488 (O_488,N_2977,N_2974);
or UO_489 (O_489,N_2974,N_2952);
nor UO_490 (O_490,N_2942,N_2984);
nand UO_491 (O_491,N_2979,N_2941);
nor UO_492 (O_492,N_2940,N_2948);
nor UO_493 (O_493,N_2998,N_2954);
nor UO_494 (O_494,N_2997,N_2957);
nand UO_495 (O_495,N_2992,N_2948);
nand UO_496 (O_496,N_2940,N_2947);
nand UO_497 (O_497,N_2973,N_2961);
xor UO_498 (O_498,N_2963,N_2981);
nand UO_499 (O_499,N_2956,N_2990);
endmodule