module basic_750_5000_1000_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_285,In_303);
or U1 (N_1,In_455,In_18);
and U2 (N_2,In_571,In_528);
and U3 (N_3,In_515,In_79);
and U4 (N_4,In_342,In_129);
and U5 (N_5,In_340,In_211);
and U6 (N_6,In_167,In_563);
and U7 (N_7,In_514,In_505);
or U8 (N_8,In_556,In_492);
nor U9 (N_9,In_678,In_623);
and U10 (N_10,In_404,In_479);
xnor U11 (N_11,In_363,In_95);
xor U12 (N_12,In_605,In_546);
and U13 (N_13,In_629,In_341);
or U14 (N_14,In_88,In_581);
xnor U15 (N_15,In_651,In_734);
or U16 (N_16,In_742,In_36);
nand U17 (N_17,In_162,In_390);
nand U18 (N_18,In_133,In_686);
xnor U19 (N_19,In_447,In_714);
nor U20 (N_20,In_444,In_520);
and U21 (N_21,In_206,In_466);
and U22 (N_22,In_712,In_674);
nor U23 (N_23,In_319,In_335);
and U24 (N_24,In_534,In_663);
nor U25 (N_25,In_609,In_282);
and U26 (N_26,In_433,In_398);
or U27 (N_27,In_707,In_576);
nor U28 (N_28,In_442,In_747);
nor U29 (N_29,In_10,In_439);
nor U30 (N_30,In_62,In_566);
nor U31 (N_31,In_538,In_558);
nand U32 (N_32,In_382,In_236);
nor U33 (N_33,In_407,In_715);
xor U34 (N_34,In_680,In_483);
or U35 (N_35,In_308,In_684);
nor U36 (N_36,In_147,In_251);
xnor U37 (N_37,In_224,In_70);
nor U38 (N_38,In_194,In_395);
xor U39 (N_39,In_735,In_518);
nand U40 (N_40,In_393,In_354);
nand U41 (N_41,In_591,In_328);
nor U42 (N_42,In_107,In_170);
or U43 (N_43,In_608,In_628);
xor U44 (N_44,In_344,In_427);
xor U45 (N_45,In_625,In_215);
nor U46 (N_46,In_358,In_740);
nor U47 (N_47,In_137,In_499);
and U48 (N_48,In_667,In_347);
nand U49 (N_49,In_592,In_66);
xor U50 (N_50,In_695,In_662);
or U51 (N_51,In_117,In_293);
and U52 (N_52,In_384,In_68);
nor U53 (N_53,In_148,In_507);
or U54 (N_54,In_632,In_336);
nand U55 (N_55,In_54,In_337);
nand U56 (N_56,In_230,In_713);
and U57 (N_57,In_74,In_654);
or U58 (N_58,In_530,In_265);
or U59 (N_59,In_50,In_590);
nand U60 (N_60,In_484,In_250);
nor U61 (N_61,In_212,In_537);
xor U62 (N_62,In_639,In_633);
nor U63 (N_63,In_216,In_535);
and U64 (N_64,In_562,In_696);
or U65 (N_65,In_233,In_600);
or U66 (N_66,In_7,In_367);
and U67 (N_67,In_320,In_174);
or U68 (N_68,In_288,In_524);
or U69 (N_69,In_136,In_181);
nand U70 (N_70,In_247,In_128);
nand U71 (N_71,In_708,In_267);
nor U72 (N_72,In_432,In_89);
xnor U73 (N_73,In_205,In_24);
and U74 (N_74,In_657,In_94);
nand U75 (N_75,In_47,In_145);
nor U76 (N_76,In_109,In_301);
and U77 (N_77,In_445,In_653);
nor U78 (N_78,In_176,In_679);
and U79 (N_79,In_182,In_346);
and U80 (N_80,In_324,In_85);
nor U81 (N_81,In_33,In_57);
and U82 (N_82,In_177,In_144);
nor U83 (N_83,In_339,In_245);
nand U84 (N_84,In_589,In_273);
nand U85 (N_85,In_456,In_417);
nor U86 (N_86,In_533,In_310);
or U87 (N_87,In_171,In_370);
or U88 (N_88,In_682,In_87);
nor U89 (N_89,In_683,In_497);
or U90 (N_90,In_116,In_65);
and U91 (N_91,In_744,In_588);
or U92 (N_92,In_98,In_688);
nor U93 (N_93,In_292,In_333);
nand U94 (N_94,In_553,In_480);
and U95 (N_95,In_32,In_501);
nand U96 (N_96,In_75,In_272);
or U97 (N_97,In_254,In_25);
or U98 (N_98,In_733,In_406);
nor U99 (N_99,In_737,In_86);
or U100 (N_100,In_352,In_257);
or U101 (N_101,In_675,In_502);
nor U102 (N_102,In_697,In_401);
xor U103 (N_103,In_329,In_659);
or U104 (N_104,In_504,In_77);
nand U105 (N_105,In_702,In_710);
and U106 (N_106,In_540,In_369);
or U107 (N_107,In_371,In_214);
nor U108 (N_108,In_193,In_631);
or U109 (N_109,In_299,In_49);
and U110 (N_110,In_490,In_378);
and U111 (N_111,In_192,In_284);
and U112 (N_112,In_616,In_749);
and U113 (N_113,In_529,In_289);
and U114 (N_114,In_186,In_727);
and U115 (N_115,In_513,In_113);
or U116 (N_116,In_29,In_721);
and U117 (N_117,In_200,In_380);
or U118 (N_118,In_239,In_154);
nor U119 (N_119,In_157,In_687);
nor U120 (N_120,In_190,In_309);
nor U121 (N_121,In_374,In_90);
or U122 (N_122,In_559,In_699);
nand U123 (N_123,In_332,In_315);
nor U124 (N_124,In_579,In_151);
and U125 (N_125,In_392,In_55);
nor U126 (N_126,In_231,In_641);
and U127 (N_127,In_138,In_468);
nor U128 (N_128,In_306,In_652);
nand U129 (N_129,In_495,In_718);
and U130 (N_130,In_202,In_656);
or U131 (N_131,In_408,In_620);
nand U132 (N_132,In_263,In_135);
and U133 (N_133,In_115,In_464);
nor U134 (N_134,In_40,In_743);
or U135 (N_135,In_436,In_291);
or U136 (N_136,In_6,In_467);
or U137 (N_137,In_706,In_201);
xor U138 (N_138,In_410,In_331);
xor U139 (N_139,In_12,In_615);
and U140 (N_140,In_711,In_361);
or U141 (N_141,In_368,In_585);
nand U142 (N_142,In_573,In_475);
or U143 (N_143,In_720,In_409);
or U144 (N_144,In_732,In_372);
or U145 (N_145,In_584,In_305);
nor U146 (N_146,In_44,In_15);
and U147 (N_147,In_106,In_21);
nand U148 (N_148,In_671,In_416);
nand U149 (N_149,In_478,In_644);
nor U150 (N_150,In_635,In_353);
or U151 (N_151,In_220,In_122);
nand U152 (N_152,In_156,In_208);
nand U153 (N_153,In_326,In_618);
and U154 (N_154,In_286,In_541);
nand U155 (N_155,In_121,In_100);
or U156 (N_156,In_27,In_542);
or U157 (N_157,In_195,In_709);
and U158 (N_158,In_161,In_738);
nand U159 (N_159,In_745,In_362);
nand U160 (N_160,In_31,In_124);
nand U161 (N_161,In_716,In_448);
nand U162 (N_162,In_681,In_460);
nor U163 (N_163,In_249,In_229);
nor U164 (N_164,In_638,In_626);
and U165 (N_165,In_330,In_237);
nor U166 (N_166,In_334,In_165);
or U167 (N_167,In_351,In_627);
or U168 (N_168,In_511,In_343);
nor U169 (N_169,In_80,In_314);
or U170 (N_170,In_127,In_350);
nand U171 (N_171,In_473,In_73);
nor U172 (N_172,In_422,In_204);
and U173 (N_173,In_96,In_166);
nor U174 (N_174,In_321,In_381);
nand U175 (N_175,In_338,In_489);
or U176 (N_176,In_131,In_421);
and U177 (N_177,In_169,In_72);
nand U178 (N_178,In_580,In_345);
xnor U179 (N_179,In_457,In_210);
nand U180 (N_180,In_42,In_424);
nand U181 (N_181,In_736,In_377);
xor U182 (N_182,In_664,In_59);
nor U183 (N_183,In_454,In_405);
nand U184 (N_184,In_287,In_394);
and U185 (N_185,In_522,In_598);
and U186 (N_186,In_403,In_112);
xor U187 (N_187,In_385,In_595);
or U188 (N_188,In_28,In_673);
and U189 (N_189,In_209,In_586);
nand U190 (N_190,In_411,In_188);
or U191 (N_191,In_748,In_389);
and U192 (N_192,In_35,In_640);
nor U193 (N_193,In_300,In_105);
and U194 (N_194,In_423,In_82);
nand U195 (N_195,In_143,In_415);
xor U196 (N_196,In_92,In_271);
nor U197 (N_197,In_649,In_431);
and U198 (N_198,In_213,In_283);
nand U199 (N_199,In_276,In_104);
and U200 (N_200,In_700,In_2);
or U201 (N_201,In_14,In_185);
nor U202 (N_202,In_426,In_601);
nand U203 (N_203,In_463,In_593);
nand U204 (N_204,In_731,In_160);
and U205 (N_205,In_471,In_232);
or U206 (N_206,In_689,In_270);
nor U207 (N_207,In_741,In_525);
or U208 (N_208,In_302,In_587);
or U209 (N_209,In_459,In_567);
or U210 (N_210,In_120,In_577);
nand U211 (N_211,In_693,In_516);
nor U212 (N_212,In_258,In_611);
xnor U213 (N_213,In_583,In_668);
nor U214 (N_214,In_677,In_304);
or U215 (N_215,In_596,In_103);
nand U216 (N_216,In_602,In_67);
and U217 (N_217,In_565,In_560);
or U218 (N_218,In_41,In_704);
or U219 (N_219,In_461,In_110);
and U220 (N_220,In_399,In_199);
nor U221 (N_221,In_730,In_114);
or U222 (N_222,In_477,In_22);
and U223 (N_223,In_387,In_56);
nor U224 (N_224,In_221,In_150);
and U225 (N_225,In_278,In_617);
or U226 (N_226,In_163,In_634);
nor U227 (N_227,In_146,In_261);
and U228 (N_228,In_3,In_451);
xor U229 (N_229,In_16,In_536);
and U230 (N_230,In_97,In_81);
xor U231 (N_231,In_313,In_544);
nand U232 (N_232,In_307,In_512);
nor U233 (N_233,In_48,In_327);
and U234 (N_234,In_400,In_207);
and U235 (N_235,In_187,In_685);
nor U236 (N_236,In_295,In_547);
nand U237 (N_237,In_597,In_246);
nor U238 (N_238,In_11,In_125);
and U239 (N_239,In_172,In_142);
xor U240 (N_240,In_219,In_509);
and U241 (N_241,In_531,In_108);
nand U242 (N_242,In_223,In_578);
nor U243 (N_243,In_256,In_443);
nor U244 (N_244,In_349,In_39);
and U245 (N_245,In_434,In_462);
nor U246 (N_246,In_366,In_99);
or U247 (N_247,In_419,In_672);
nand U248 (N_248,In_189,In_373);
or U249 (N_249,In_348,In_435);
and U250 (N_250,In_365,In_391);
nand U251 (N_251,In_506,In_84);
or U252 (N_252,In_260,In_38);
and U253 (N_253,In_676,In_452);
and U254 (N_254,In_413,In_521);
xor U255 (N_255,In_101,In_575);
nor U256 (N_256,In_388,In_312);
and U257 (N_257,In_102,In_690);
and U258 (N_258,In_17,In_5);
or U259 (N_259,In_123,In_13);
nand U260 (N_260,In_76,In_294);
nand U261 (N_261,In_396,In_316);
xor U262 (N_262,In_482,In_164);
or U263 (N_263,In_496,In_594);
nand U264 (N_264,In_179,In_43);
xnor U265 (N_265,In_621,In_655);
or U266 (N_266,In_83,In_572);
or U267 (N_267,In_545,In_63);
and U268 (N_268,In_666,In_375);
xnor U269 (N_269,In_527,In_45);
nand U270 (N_270,In_607,In_397);
nor U271 (N_271,In_158,In_141);
and U272 (N_272,In_196,In_93);
or U273 (N_273,In_60,In_425);
or U274 (N_274,In_551,In_357);
nand U275 (N_275,In_429,In_268);
nor U276 (N_276,In_152,In_637);
or U277 (N_277,In_203,In_485);
or U278 (N_278,In_379,In_23);
or U279 (N_279,In_487,In_446);
nor U280 (N_280,In_494,In_184);
nor U281 (N_281,In_266,In_488);
or U282 (N_282,In_61,In_183);
nor U283 (N_283,In_437,In_222);
nand U284 (N_284,In_134,In_722);
and U285 (N_285,In_8,In_554);
and U286 (N_286,In_225,In_360);
and U287 (N_287,In_500,In_604);
nor U288 (N_288,In_111,In_280);
and U289 (N_289,In_610,In_642);
and U290 (N_290,In_481,In_275);
nor U291 (N_291,In_561,In_178);
and U292 (N_292,In_726,In_472);
or U293 (N_293,In_168,In_78);
xnor U294 (N_294,In_139,In_355);
and U295 (N_295,In_614,In_318);
nand U296 (N_296,In_240,In_549);
nand U297 (N_297,In_255,In_430);
and U298 (N_298,In_235,In_130);
or U299 (N_299,In_119,In_498);
nor U300 (N_300,In_149,In_218);
nor U301 (N_301,In_570,In_645);
and U302 (N_302,In_636,In_91);
nand U303 (N_303,In_4,In_317);
nand U304 (N_304,In_648,In_717);
and U305 (N_305,In_465,In_725);
and U306 (N_306,In_650,In_550);
nand U307 (N_307,In_582,In_274);
nand U308 (N_308,In_26,In_19);
or U309 (N_309,In_386,In_281);
or U310 (N_310,In_647,In_724);
or U311 (N_311,In_269,In_30);
and U312 (N_312,In_476,In_691);
or U313 (N_313,In_418,In_552);
nor U314 (N_314,In_248,In_264);
or U315 (N_315,In_729,In_69);
or U316 (N_316,In_450,In_428);
and U317 (N_317,In_526,In_624);
xnor U318 (N_318,In_491,In_440);
nor U319 (N_319,In_180,In_118);
or U320 (N_320,In_252,In_279);
and U321 (N_321,In_458,In_197);
nand U322 (N_322,In_420,In_242);
or U323 (N_323,In_414,In_568);
and U324 (N_324,In_52,In_723);
nand U325 (N_325,In_493,In_503);
and U326 (N_326,In_159,In_34);
and U327 (N_327,In_630,In_132);
nor U328 (N_328,In_297,In_262);
nand U329 (N_329,In_259,In_217);
nand U330 (N_330,In_539,In_606);
or U331 (N_331,In_441,In_728);
and U332 (N_332,In_449,In_64);
nor U333 (N_333,In_228,In_453);
xnor U334 (N_334,In_198,In_277);
nand U335 (N_335,In_719,In_569);
nor U336 (N_336,In_508,In_701);
and U337 (N_337,In_140,In_519);
and U338 (N_338,In_227,In_705);
or U339 (N_339,In_244,In_1);
xor U340 (N_340,In_322,In_746);
and U341 (N_341,In_323,In_665);
nor U342 (N_342,In_486,In_234);
nor U343 (N_343,In_226,In_37);
or U344 (N_344,In_613,In_243);
nand U345 (N_345,In_356,In_155);
and U346 (N_346,In_692,In_469);
nand U347 (N_347,In_9,In_470);
or U348 (N_348,In_574,In_298);
or U349 (N_349,In_660,In_646);
xor U350 (N_350,In_612,In_622);
nor U351 (N_351,In_661,In_643);
nand U352 (N_352,In_253,In_694);
nor U353 (N_353,In_175,In_543);
nor U354 (N_354,In_698,In_739);
nand U355 (N_355,In_670,In_703);
xnor U356 (N_356,In_548,In_412);
and U357 (N_357,In_53,In_126);
or U358 (N_358,In_71,In_658);
xnor U359 (N_359,In_517,In_438);
xor U360 (N_360,In_58,In_619);
and U361 (N_361,In_296,In_523);
and U362 (N_362,In_46,In_290);
nand U363 (N_363,In_383,In_153);
nor U364 (N_364,In_599,In_20);
nand U365 (N_365,In_325,In_173);
xnor U366 (N_366,In_474,In_557);
nor U367 (N_367,In_311,In_510);
or U368 (N_368,In_376,In_555);
and U369 (N_369,In_402,In_564);
nand U370 (N_370,In_603,In_669);
nand U371 (N_371,In_359,In_191);
and U372 (N_372,In_532,In_241);
nor U373 (N_373,In_0,In_364);
or U374 (N_374,In_238,In_51);
nor U375 (N_375,In_556,In_639);
or U376 (N_376,In_540,In_658);
nor U377 (N_377,In_436,In_297);
xnor U378 (N_378,In_394,In_512);
and U379 (N_379,In_311,In_100);
or U380 (N_380,In_24,In_492);
and U381 (N_381,In_417,In_363);
nor U382 (N_382,In_412,In_319);
nand U383 (N_383,In_5,In_562);
and U384 (N_384,In_607,In_654);
nand U385 (N_385,In_136,In_382);
xor U386 (N_386,In_607,In_22);
and U387 (N_387,In_387,In_683);
xor U388 (N_388,In_670,In_33);
nand U389 (N_389,In_572,In_254);
nor U390 (N_390,In_657,In_373);
nor U391 (N_391,In_294,In_456);
or U392 (N_392,In_135,In_83);
nand U393 (N_393,In_276,In_148);
nand U394 (N_394,In_384,In_369);
nand U395 (N_395,In_129,In_422);
and U396 (N_396,In_43,In_294);
xnor U397 (N_397,In_535,In_258);
nand U398 (N_398,In_735,In_122);
and U399 (N_399,In_357,In_194);
xnor U400 (N_400,In_175,In_489);
xnor U401 (N_401,In_159,In_535);
nor U402 (N_402,In_254,In_119);
and U403 (N_403,In_572,In_564);
or U404 (N_404,In_696,In_547);
and U405 (N_405,In_283,In_458);
or U406 (N_406,In_315,In_537);
or U407 (N_407,In_5,In_330);
and U408 (N_408,In_302,In_272);
and U409 (N_409,In_332,In_664);
nor U410 (N_410,In_464,In_365);
or U411 (N_411,In_161,In_387);
xnor U412 (N_412,In_453,In_555);
or U413 (N_413,In_416,In_488);
xor U414 (N_414,In_494,In_375);
nand U415 (N_415,In_532,In_337);
nand U416 (N_416,In_46,In_347);
or U417 (N_417,In_719,In_348);
nor U418 (N_418,In_471,In_610);
or U419 (N_419,In_612,In_236);
nor U420 (N_420,In_416,In_277);
nand U421 (N_421,In_227,In_224);
nor U422 (N_422,In_341,In_420);
nand U423 (N_423,In_460,In_128);
xnor U424 (N_424,In_190,In_289);
or U425 (N_425,In_663,In_361);
nor U426 (N_426,In_439,In_128);
nand U427 (N_427,In_75,In_715);
xnor U428 (N_428,In_403,In_58);
nor U429 (N_429,In_125,In_40);
nand U430 (N_430,In_610,In_497);
nor U431 (N_431,In_68,In_529);
and U432 (N_432,In_402,In_526);
xnor U433 (N_433,In_579,In_20);
and U434 (N_434,In_571,In_428);
nor U435 (N_435,In_683,In_630);
or U436 (N_436,In_414,In_492);
nor U437 (N_437,In_643,In_594);
nor U438 (N_438,In_686,In_379);
nand U439 (N_439,In_202,In_565);
nand U440 (N_440,In_599,In_643);
nand U441 (N_441,In_456,In_21);
nor U442 (N_442,In_490,In_312);
nor U443 (N_443,In_498,In_51);
and U444 (N_444,In_243,In_494);
or U445 (N_445,In_96,In_297);
xnor U446 (N_446,In_44,In_116);
nor U447 (N_447,In_171,In_741);
or U448 (N_448,In_70,In_84);
nor U449 (N_449,In_603,In_487);
and U450 (N_450,In_304,In_324);
xnor U451 (N_451,In_677,In_29);
or U452 (N_452,In_603,In_175);
or U453 (N_453,In_149,In_151);
nand U454 (N_454,In_718,In_262);
nor U455 (N_455,In_21,In_348);
nor U456 (N_456,In_575,In_465);
nand U457 (N_457,In_607,In_655);
nand U458 (N_458,In_301,In_112);
nand U459 (N_459,In_10,In_719);
and U460 (N_460,In_11,In_136);
nor U461 (N_461,In_331,In_339);
or U462 (N_462,In_626,In_671);
nand U463 (N_463,In_437,In_291);
or U464 (N_464,In_440,In_71);
nor U465 (N_465,In_282,In_177);
nor U466 (N_466,In_730,In_120);
or U467 (N_467,In_574,In_101);
or U468 (N_468,In_656,In_555);
and U469 (N_469,In_564,In_299);
nor U470 (N_470,In_564,In_14);
or U471 (N_471,In_76,In_680);
and U472 (N_472,In_510,In_583);
nor U473 (N_473,In_593,In_186);
nor U474 (N_474,In_704,In_180);
nor U475 (N_475,In_120,In_569);
nor U476 (N_476,In_741,In_307);
nor U477 (N_477,In_291,In_642);
nor U478 (N_478,In_169,In_45);
or U479 (N_479,In_503,In_403);
or U480 (N_480,In_682,In_16);
and U481 (N_481,In_356,In_674);
xnor U482 (N_482,In_595,In_89);
nand U483 (N_483,In_487,In_459);
and U484 (N_484,In_368,In_702);
or U485 (N_485,In_524,In_592);
or U486 (N_486,In_271,In_264);
or U487 (N_487,In_276,In_487);
nand U488 (N_488,In_723,In_264);
xor U489 (N_489,In_194,In_122);
and U490 (N_490,In_570,In_170);
nor U491 (N_491,In_406,In_565);
nor U492 (N_492,In_673,In_639);
and U493 (N_493,In_748,In_593);
nand U494 (N_494,In_393,In_123);
nand U495 (N_495,In_57,In_711);
xor U496 (N_496,In_87,In_168);
nand U497 (N_497,In_557,In_401);
and U498 (N_498,In_127,In_437);
or U499 (N_499,In_286,In_90);
nor U500 (N_500,N_104,N_92);
nand U501 (N_501,N_354,N_296);
xnor U502 (N_502,N_139,N_345);
and U503 (N_503,N_51,N_118);
nor U504 (N_504,N_88,N_406);
nor U505 (N_505,N_372,N_281);
or U506 (N_506,N_140,N_400);
nor U507 (N_507,N_379,N_63);
or U508 (N_508,N_324,N_55);
nor U509 (N_509,N_327,N_457);
and U510 (N_510,N_13,N_87);
xor U511 (N_511,N_267,N_276);
or U512 (N_512,N_444,N_52);
nand U513 (N_513,N_393,N_154);
nor U514 (N_514,N_263,N_355);
and U515 (N_515,N_259,N_65);
nor U516 (N_516,N_349,N_423);
nand U517 (N_517,N_223,N_28);
nor U518 (N_518,N_152,N_231);
nand U519 (N_519,N_463,N_269);
and U520 (N_520,N_472,N_19);
nor U521 (N_521,N_342,N_71);
and U522 (N_522,N_204,N_486);
nor U523 (N_523,N_390,N_435);
and U524 (N_524,N_209,N_405);
nor U525 (N_525,N_326,N_158);
and U526 (N_526,N_16,N_280);
and U527 (N_527,N_262,N_432);
nor U528 (N_528,N_242,N_471);
nor U529 (N_529,N_235,N_311);
nor U530 (N_530,N_145,N_381);
nor U531 (N_531,N_184,N_344);
and U532 (N_532,N_214,N_144);
nand U533 (N_533,N_50,N_308);
nor U534 (N_534,N_243,N_39);
and U535 (N_535,N_226,N_234);
nand U536 (N_536,N_285,N_80);
nor U537 (N_537,N_377,N_93);
or U538 (N_538,N_389,N_112);
nor U539 (N_539,N_241,N_388);
xor U540 (N_540,N_356,N_272);
nand U541 (N_541,N_45,N_199);
nor U542 (N_542,N_190,N_75);
nor U543 (N_543,N_481,N_477);
nor U544 (N_544,N_206,N_341);
nor U545 (N_545,N_462,N_96);
and U546 (N_546,N_394,N_153);
and U547 (N_547,N_11,N_361);
nor U548 (N_548,N_443,N_76);
nand U549 (N_549,N_44,N_362);
and U550 (N_550,N_32,N_151);
and U551 (N_551,N_286,N_191);
nor U552 (N_552,N_358,N_165);
nor U553 (N_553,N_168,N_319);
nand U554 (N_554,N_136,N_9);
or U555 (N_555,N_34,N_429);
or U556 (N_556,N_53,N_447);
xnor U557 (N_557,N_498,N_185);
and U558 (N_558,N_0,N_363);
xnor U559 (N_559,N_428,N_111);
xor U560 (N_560,N_227,N_255);
nand U561 (N_561,N_284,N_279);
xor U562 (N_562,N_146,N_245);
xor U563 (N_563,N_219,N_137);
nand U564 (N_564,N_6,N_431);
and U565 (N_565,N_480,N_120);
and U566 (N_566,N_407,N_375);
nand U567 (N_567,N_482,N_192);
nor U568 (N_568,N_290,N_339);
nand U569 (N_569,N_367,N_395);
nor U570 (N_570,N_312,N_304);
nand U571 (N_571,N_86,N_261);
nand U572 (N_572,N_173,N_494);
xnor U573 (N_573,N_236,N_2);
or U574 (N_574,N_205,N_133);
nor U575 (N_575,N_91,N_313);
and U576 (N_576,N_253,N_40);
and U577 (N_577,N_15,N_217);
and U578 (N_578,N_222,N_239);
nor U579 (N_579,N_195,N_66);
nand U580 (N_580,N_121,N_484);
nand U581 (N_581,N_371,N_427);
nand U582 (N_582,N_413,N_3);
xor U583 (N_583,N_161,N_456);
or U584 (N_584,N_335,N_421);
or U585 (N_585,N_257,N_115);
and U586 (N_586,N_433,N_424);
xnor U587 (N_587,N_113,N_249);
nor U588 (N_588,N_17,N_186);
and U589 (N_589,N_454,N_174);
or U590 (N_590,N_418,N_159);
xnor U591 (N_591,N_221,N_399);
and U592 (N_592,N_141,N_126);
nand U593 (N_593,N_365,N_175);
nand U594 (N_594,N_46,N_114);
and U595 (N_595,N_301,N_321);
and U596 (N_596,N_378,N_440);
and U597 (N_597,N_7,N_69);
or U598 (N_598,N_26,N_387);
and U599 (N_599,N_232,N_189);
nor U600 (N_600,N_446,N_216);
and U601 (N_601,N_207,N_305);
xor U602 (N_602,N_202,N_396);
nor U603 (N_603,N_41,N_420);
xnor U604 (N_604,N_260,N_122);
and U605 (N_605,N_167,N_169);
and U606 (N_606,N_451,N_62);
xor U607 (N_607,N_374,N_442);
and U608 (N_608,N_397,N_64);
nor U609 (N_609,N_156,N_176);
or U610 (N_610,N_439,N_47);
and U611 (N_611,N_54,N_282);
xnor U612 (N_612,N_36,N_128);
or U613 (N_613,N_49,N_203);
or U614 (N_614,N_225,N_148);
or U615 (N_615,N_157,N_437);
nand U616 (N_616,N_270,N_409);
nor U617 (N_617,N_359,N_74);
nand U618 (N_618,N_376,N_380);
nor U619 (N_619,N_14,N_89);
or U620 (N_620,N_67,N_455);
or U621 (N_621,N_487,N_132);
and U622 (N_622,N_97,N_177);
or U623 (N_623,N_228,N_470);
nand U624 (N_624,N_287,N_127);
and U625 (N_625,N_33,N_322);
or U626 (N_626,N_331,N_1);
nand U627 (N_627,N_254,N_201);
nor U628 (N_628,N_27,N_70);
xnor U629 (N_629,N_213,N_138);
and U630 (N_630,N_338,N_103);
or U631 (N_631,N_419,N_237);
nand U632 (N_632,N_408,N_283);
or U633 (N_633,N_117,N_197);
nand U634 (N_634,N_317,N_398);
nand U635 (N_635,N_271,N_266);
and U636 (N_636,N_252,N_179);
or U637 (N_637,N_12,N_476);
nor U638 (N_638,N_277,N_58);
nor U639 (N_639,N_323,N_330);
or U640 (N_640,N_496,N_320);
nand U641 (N_641,N_109,N_475);
and U642 (N_642,N_57,N_85);
nand U643 (N_643,N_465,N_188);
or U644 (N_644,N_315,N_61);
nor U645 (N_645,N_495,N_147);
nand U646 (N_646,N_134,N_43);
or U647 (N_647,N_404,N_488);
nor U648 (N_648,N_81,N_450);
nor U649 (N_649,N_79,N_302);
or U650 (N_650,N_460,N_499);
xor U651 (N_651,N_247,N_461);
and U652 (N_652,N_170,N_83);
and U653 (N_653,N_23,N_108);
and U654 (N_654,N_212,N_211);
nand U655 (N_655,N_278,N_178);
nor U656 (N_656,N_448,N_384);
and U657 (N_657,N_306,N_401);
nor U658 (N_658,N_422,N_493);
nand U659 (N_659,N_392,N_351);
and U660 (N_660,N_265,N_68);
or U661 (N_661,N_467,N_402);
nand U662 (N_662,N_386,N_100);
nand U663 (N_663,N_329,N_491);
or U664 (N_664,N_347,N_468);
and U665 (N_665,N_171,N_105);
nor U666 (N_666,N_18,N_123);
and U667 (N_667,N_56,N_38);
or U668 (N_668,N_72,N_426);
xor U669 (N_669,N_198,N_416);
xnor U670 (N_670,N_452,N_60);
nor U671 (N_671,N_8,N_303);
nor U672 (N_672,N_98,N_293);
or U673 (N_673,N_129,N_314);
and U674 (N_674,N_233,N_230);
nand U675 (N_675,N_357,N_258);
nor U676 (N_676,N_194,N_383);
nand U677 (N_677,N_441,N_430);
or U678 (N_678,N_490,N_385);
nor U679 (N_679,N_200,N_5);
nor U680 (N_680,N_343,N_110);
nand U681 (N_681,N_298,N_350);
and U682 (N_682,N_164,N_410);
xnor U683 (N_683,N_309,N_155);
and U684 (N_684,N_334,N_474);
and U685 (N_685,N_59,N_336);
nand U686 (N_686,N_248,N_31);
xnor U687 (N_687,N_149,N_166);
nor U688 (N_688,N_469,N_391);
and U689 (N_689,N_143,N_288);
or U690 (N_690,N_22,N_449);
nor U691 (N_691,N_412,N_292);
or U692 (N_692,N_483,N_160);
nand U693 (N_693,N_492,N_37);
or U694 (N_694,N_466,N_150);
or U695 (N_695,N_220,N_182);
nand U696 (N_696,N_42,N_251);
nand U697 (N_697,N_473,N_415);
nor U698 (N_698,N_135,N_82);
and U699 (N_699,N_130,N_464);
and U700 (N_700,N_453,N_4);
xnor U701 (N_701,N_180,N_163);
and U702 (N_702,N_90,N_21);
nor U703 (N_703,N_224,N_116);
or U704 (N_704,N_268,N_196);
xor U705 (N_705,N_94,N_310);
nand U706 (N_706,N_346,N_240);
or U707 (N_707,N_333,N_478);
xor U708 (N_708,N_438,N_99);
or U709 (N_709,N_295,N_337);
and U710 (N_710,N_183,N_497);
or U711 (N_711,N_10,N_294);
nor U712 (N_712,N_291,N_48);
and U713 (N_713,N_364,N_25);
or U714 (N_714,N_373,N_300);
and U715 (N_715,N_238,N_172);
nand U716 (N_716,N_30,N_325);
nand U717 (N_717,N_425,N_95);
and U718 (N_718,N_368,N_414);
nor U719 (N_719,N_193,N_250);
and U720 (N_720,N_35,N_289);
nor U721 (N_721,N_417,N_218);
or U722 (N_722,N_229,N_299);
or U723 (N_723,N_479,N_256);
nand U724 (N_724,N_352,N_125);
nand U725 (N_725,N_107,N_370);
and U726 (N_726,N_29,N_181);
and U727 (N_727,N_489,N_318);
and U728 (N_728,N_459,N_131);
and U729 (N_729,N_24,N_332);
and U730 (N_730,N_275,N_101);
nand U731 (N_731,N_124,N_297);
xnor U732 (N_732,N_210,N_340);
or U733 (N_733,N_434,N_328);
or U734 (N_734,N_162,N_458);
and U735 (N_735,N_77,N_316);
or U736 (N_736,N_353,N_436);
xor U737 (N_737,N_273,N_360);
or U738 (N_738,N_485,N_208);
nor U739 (N_739,N_403,N_411);
and U740 (N_740,N_369,N_244);
xor U741 (N_741,N_246,N_348);
nand U742 (N_742,N_187,N_106);
and U743 (N_743,N_382,N_102);
or U744 (N_744,N_366,N_78);
and U745 (N_745,N_142,N_215);
and U746 (N_746,N_73,N_84);
or U747 (N_747,N_20,N_274);
nand U748 (N_748,N_264,N_307);
nor U749 (N_749,N_445,N_119);
and U750 (N_750,N_289,N_214);
nand U751 (N_751,N_434,N_400);
and U752 (N_752,N_18,N_153);
xor U753 (N_753,N_370,N_7);
nand U754 (N_754,N_22,N_137);
or U755 (N_755,N_166,N_380);
or U756 (N_756,N_200,N_165);
and U757 (N_757,N_75,N_266);
nor U758 (N_758,N_374,N_269);
nor U759 (N_759,N_455,N_159);
or U760 (N_760,N_345,N_384);
or U761 (N_761,N_312,N_475);
nor U762 (N_762,N_162,N_466);
nand U763 (N_763,N_448,N_285);
xnor U764 (N_764,N_288,N_265);
and U765 (N_765,N_302,N_27);
and U766 (N_766,N_79,N_238);
or U767 (N_767,N_331,N_14);
or U768 (N_768,N_246,N_382);
nand U769 (N_769,N_254,N_347);
xor U770 (N_770,N_375,N_266);
nand U771 (N_771,N_314,N_249);
nor U772 (N_772,N_80,N_189);
xnor U773 (N_773,N_343,N_283);
and U774 (N_774,N_348,N_51);
or U775 (N_775,N_497,N_490);
or U776 (N_776,N_287,N_167);
or U777 (N_777,N_331,N_191);
nor U778 (N_778,N_33,N_363);
nor U779 (N_779,N_236,N_348);
nand U780 (N_780,N_462,N_10);
nor U781 (N_781,N_285,N_238);
xor U782 (N_782,N_120,N_229);
nor U783 (N_783,N_296,N_300);
or U784 (N_784,N_80,N_259);
nand U785 (N_785,N_171,N_434);
and U786 (N_786,N_431,N_78);
nor U787 (N_787,N_11,N_324);
nor U788 (N_788,N_174,N_59);
xor U789 (N_789,N_183,N_3);
and U790 (N_790,N_373,N_479);
nand U791 (N_791,N_476,N_404);
nor U792 (N_792,N_279,N_429);
nor U793 (N_793,N_464,N_105);
or U794 (N_794,N_231,N_321);
and U795 (N_795,N_433,N_33);
nor U796 (N_796,N_25,N_30);
nor U797 (N_797,N_218,N_336);
nand U798 (N_798,N_108,N_314);
nand U799 (N_799,N_429,N_173);
nor U800 (N_800,N_340,N_90);
nor U801 (N_801,N_280,N_236);
or U802 (N_802,N_227,N_75);
or U803 (N_803,N_63,N_472);
or U804 (N_804,N_141,N_358);
nor U805 (N_805,N_51,N_262);
nor U806 (N_806,N_256,N_182);
xor U807 (N_807,N_126,N_455);
xnor U808 (N_808,N_61,N_45);
nor U809 (N_809,N_110,N_464);
nand U810 (N_810,N_304,N_234);
nor U811 (N_811,N_66,N_17);
nor U812 (N_812,N_441,N_76);
nor U813 (N_813,N_134,N_413);
and U814 (N_814,N_296,N_57);
nor U815 (N_815,N_192,N_326);
or U816 (N_816,N_322,N_234);
nor U817 (N_817,N_13,N_495);
nand U818 (N_818,N_312,N_462);
nand U819 (N_819,N_210,N_31);
nor U820 (N_820,N_84,N_109);
nor U821 (N_821,N_457,N_63);
nand U822 (N_822,N_69,N_199);
nand U823 (N_823,N_275,N_233);
nor U824 (N_824,N_363,N_78);
nand U825 (N_825,N_290,N_19);
or U826 (N_826,N_403,N_192);
nand U827 (N_827,N_371,N_266);
xor U828 (N_828,N_157,N_401);
or U829 (N_829,N_485,N_479);
or U830 (N_830,N_450,N_184);
nor U831 (N_831,N_166,N_122);
xor U832 (N_832,N_278,N_124);
nor U833 (N_833,N_266,N_439);
xor U834 (N_834,N_495,N_26);
nor U835 (N_835,N_372,N_66);
and U836 (N_836,N_332,N_159);
nor U837 (N_837,N_234,N_175);
xor U838 (N_838,N_412,N_191);
and U839 (N_839,N_251,N_215);
nor U840 (N_840,N_177,N_94);
or U841 (N_841,N_312,N_1);
or U842 (N_842,N_395,N_465);
xnor U843 (N_843,N_263,N_42);
nand U844 (N_844,N_265,N_477);
nor U845 (N_845,N_217,N_32);
nand U846 (N_846,N_487,N_473);
and U847 (N_847,N_413,N_471);
or U848 (N_848,N_238,N_388);
nor U849 (N_849,N_409,N_212);
and U850 (N_850,N_298,N_293);
nor U851 (N_851,N_306,N_104);
nand U852 (N_852,N_208,N_298);
nand U853 (N_853,N_378,N_135);
or U854 (N_854,N_387,N_243);
and U855 (N_855,N_339,N_58);
or U856 (N_856,N_493,N_402);
and U857 (N_857,N_163,N_452);
or U858 (N_858,N_204,N_344);
or U859 (N_859,N_92,N_50);
nor U860 (N_860,N_21,N_275);
or U861 (N_861,N_224,N_274);
nand U862 (N_862,N_466,N_152);
nor U863 (N_863,N_430,N_69);
nand U864 (N_864,N_460,N_29);
nand U865 (N_865,N_362,N_344);
nor U866 (N_866,N_471,N_144);
xor U867 (N_867,N_432,N_314);
and U868 (N_868,N_123,N_474);
or U869 (N_869,N_452,N_171);
nand U870 (N_870,N_76,N_482);
or U871 (N_871,N_201,N_386);
or U872 (N_872,N_224,N_227);
nor U873 (N_873,N_117,N_211);
and U874 (N_874,N_91,N_352);
xnor U875 (N_875,N_374,N_365);
nor U876 (N_876,N_64,N_233);
xnor U877 (N_877,N_401,N_177);
nor U878 (N_878,N_143,N_487);
nand U879 (N_879,N_368,N_236);
or U880 (N_880,N_430,N_95);
xnor U881 (N_881,N_126,N_459);
xnor U882 (N_882,N_90,N_62);
nor U883 (N_883,N_35,N_216);
nor U884 (N_884,N_305,N_326);
xnor U885 (N_885,N_329,N_478);
and U886 (N_886,N_201,N_97);
and U887 (N_887,N_347,N_180);
nand U888 (N_888,N_237,N_167);
and U889 (N_889,N_43,N_315);
or U890 (N_890,N_465,N_223);
and U891 (N_891,N_473,N_70);
and U892 (N_892,N_14,N_48);
and U893 (N_893,N_316,N_432);
nand U894 (N_894,N_313,N_169);
or U895 (N_895,N_450,N_349);
nand U896 (N_896,N_351,N_407);
or U897 (N_897,N_288,N_280);
or U898 (N_898,N_187,N_296);
nand U899 (N_899,N_476,N_316);
nor U900 (N_900,N_215,N_28);
and U901 (N_901,N_430,N_212);
nand U902 (N_902,N_7,N_228);
nand U903 (N_903,N_325,N_399);
nand U904 (N_904,N_389,N_71);
nand U905 (N_905,N_458,N_6);
and U906 (N_906,N_59,N_479);
nand U907 (N_907,N_17,N_167);
nor U908 (N_908,N_140,N_131);
xor U909 (N_909,N_427,N_109);
and U910 (N_910,N_181,N_9);
or U911 (N_911,N_95,N_32);
or U912 (N_912,N_450,N_96);
nor U913 (N_913,N_429,N_404);
nand U914 (N_914,N_378,N_271);
nor U915 (N_915,N_287,N_269);
and U916 (N_916,N_153,N_353);
and U917 (N_917,N_364,N_316);
or U918 (N_918,N_122,N_201);
nand U919 (N_919,N_344,N_319);
nand U920 (N_920,N_2,N_345);
and U921 (N_921,N_258,N_24);
or U922 (N_922,N_464,N_278);
or U923 (N_923,N_330,N_499);
nand U924 (N_924,N_165,N_245);
xnor U925 (N_925,N_9,N_156);
or U926 (N_926,N_431,N_169);
nor U927 (N_927,N_425,N_443);
nor U928 (N_928,N_421,N_419);
nor U929 (N_929,N_149,N_172);
and U930 (N_930,N_384,N_299);
nand U931 (N_931,N_384,N_52);
nand U932 (N_932,N_366,N_464);
nand U933 (N_933,N_60,N_478);
or U934 (N_934,N_70,N_21);
nor U935 (N_935,N_447,N_424);
and U936 (N_936,N_332,N_95);
nor U937 (N_937,N_405,N_425);
or U938 (N_938,N_323,N_171);
nand U939 (N_939,N_491,N_271);
or U940 (N_940,N_454,N_211);
nor U941 (N_941,N_61,N_179);
nor U942 (N_942,N_48,N_345);
and U943 (N_943,N_90,N_122);
xnor U944 (N_944,N_340,N_441);
and U945 (N_945,N_319,N_273);
and U946 (N_946,N_434,N_182);
or U947 (N_947,N_14,N_434);
nor U948 (N_948,N_94,N_135);
nor U949 (N_949,N_292,N_116);
or U950 (N_950,N_53,N_319);
nand U951 (N_951,N_2,N_244);
nand U952 (N_952,N_207,N_239);
nand U953 (N_953,N_70,N_486);
or U954 (N_954,N_141,N_11);
and U955 (N_955,N_163,N_211);
and U956 (N_956,N_226,N_380);
nor U957 (N_957,N_36,N_298);
nor U958 (N_958,N_130,N_283);
nor U959 (N_959,N_460,N_46);
nor U960 (N_960,N_433,N_409);
or U961 (N_961,N_114,N_38);
nor U962 (N_962,N_24,N_200);
xnor U963 (N_963,N_374,N_182);
nor U964 (N_964,N_161,N_74);
and U965 (N_965,N_444,N_295);
or U966 (N_966,N_309,N_266);
xnor U967 (N_967,N_279,N_272);
nand U968 (N_968,N_208,N_452);
or U969 (N_969,N_349,N_319);
nor U970 (N_970,N_442,N_201);
nor U971 (N_971,N_44,N_206);
nand U972 (N_972,N_321,N_309);
and U973 (N_973,N_154,N_485);
and U974 (N_974,N_86,N_293);
nand U975 (N_975,N_439,N_103);
or U976 (N_976,N_84,N_123);
nand U977 (N_977,N_221,N_441);
and U978 (N_978,N_66,N_36);
or U979 (N_979,N_258,N_370);
nand U980 (N_980,N_489,N_6);
or U981 (N_981,N_119,N_35);
and U982 (N_982,N_122,N_374);
nand U983 (N_983,N_465,N_382);
xor U984 (N_984,N_21,N_376);
and U985 (N_985,N_356,N_326);
and U986 (N_986,N_291,N_14);
nor U987 (N_987,N_165,N_143);
and U988 (N_988,N_218,N_421);
nor U989 (N_989,N_67,N_32);
and U990 (N_990,N_177,N_485);
or U991 (N_991,N_97,N_451);
and U992 (N_992,N_328,N_150);
and U993 (N_993,N_256,N_197);
nor U994 (N_994,N_265,N_262);
and U995 (N_995,N_403,N_292);
nor U996 (N_996,N_491,N_394);
or U997 (N_997,N_84,N_13);
or U998 (N_998,N_246,N_153);
and U999 (N_999,N_397,N_90);
and U1000 (N_1000,N_972,N_589);
or U1001 (N_1001,N_593,N_629);
nand U1002 (N_1002,N_640,N_663);
nor U1003 (N_1003,N_917,N_509);
or U1004 (N_1004,N_909,N_967);
nor U1005 (N_1005,N_694,N_821);
nor U1006 (N_1006,N_881,N_591);
or U1007 (N_1007,N_634,N_770);
or U1008 (N_1008,N_583,N_944);
nand U1009 (N_1009,N_928,N_960);
or U1010 (N_1010,N_708,N_735);
or U1011 (N_1011,N_789,N_991);
xnor U1012 (N_1012,N_807,N_810);
nor U1013 (N_1013,N_752,N_938);
nor U1014 (N_1014,N_986,N_844);
and U1015 (N_1015,N_984,N_706);
or U1016 (N_1016,N_685,N_876);
nand U1017 (N_1017,N_519,N_504);
nor U1018 (N_1018,N_673,N_966);
and U1019 (N_1019,N_920,N_771);
nand U1020 (N_1020,N_571,N_666);
or U1021 (N_1021,N_647,N_761);
nor U1022 (N_1022,N_992,N_786);
nand U1023 (N_1023,N_719,N_897);
or U1024 (N_1024,N_563,N_850);
and U1025 (N_1025,N_532,N_644);
nand U1026 (N_1026,N_689,N_621);
or U1027 (N_1027,N_934,N_747);
and U1028 (N_1028,N_985,N_699);
nor U1029 (N_1029,N_787,N_904);
and U1030 (N_1030,N_603,N_531);
and U1031 (N_1031,N_683,N_562);
or U1032 (N_1032,N_641,N_868);
nor U1033 (N_1033,N_619,N_534);
nand U1034 (N_1034,N_742,N_906);
nor U1035 (N_1035,N_746,N_713);
nor U1036 (N_1036,N_880,N_614);
nor U1037 (N_1037,N_919,N_801);
or U1038 (N_1038,N_542,N_628);
and U1039 (N_1039,N_592,N_914);
nor U1040 (N_1040,N_611,N_602);
and U1041 (N_1041,N_744,N_768);
or U1042 (N_1042,N_971,N_533);
or U1043 (N_1043,N_775,N_808);
or U1044 (N_1044,N_882,N_740);
or U1045 (N_1045,N_861,N_728);
and U1046 (N_1046,N_760,N_849);
nand U1047 (N_1047,N_525,N_726);
nor U1048 (N_1048,N_669,N_825);
nand U1049 (N_1049,N_851,N_766);
or U1050 (N_1050,N_942,N_837);
nand U1051 (N_1051,N_951,N_998);
and U1052 (N_1052,N_530,N_921);
nor U1053 (N_1053,N_668,N_645);
or U1054 (N_1054,N_975,N_551);
or U1055 (N_1055,N_968,N_883);
and U1056 (N_1056,N_983,N_774);
nor U1057 (N_1057,N_935,N_756);
nor U1058 (N_1058,N_510,N_762);
and U1059 (N_1059,N_853,N_556);
nor U1060 (N_1060,N_675,N_651);
xnor U1061 (N_1061,N_863,N_721);
and U1062 (N_1062,N_702,N_627);
nand U1063 (N_1063,N_577,N_950);
nand U1064 (N_1064,N_930,N_672);
and U1065 (N_1065,N_833,N_703);
or U1066 (N_1066,N_979,N_654);
or U1067 (N_1067,N_576,N_748);
nand U1068 (N_1068,N_587,N_598);
xor U1069 (N_1069,N_506,N_847);
nor U1070 (N_1070,N_658,N_927);
nand U1071 (N_1071,N_759,N_639);
nand U1072 (N_1072,N_829,N_918);
nor U1073 (N_1073,N_554,N_780);
and U1074 (N_1074,N_581,N_965);
and U1075 (N_1075,N_862,N_945);
nand U1076 (N_1076,N_933,N_501);
nand U1077 (N_1077,N_815,N_676);
and U1078 (N_1078,N_846,N_769);
nor U1079 (N_1079,N_867,N_575);
and U1080 (N_1080,N_782,N_947);
nand U1081 (N_1081,N_600,N_606);
nand U1082 (N_1082,N_548,N_535);
xnor U1083 (N_1083,N_503,N_572);
and U1084 (N_1084,N_677,N_910);
and U1085 (N_1085,N_637,N_860);
or U1086 (N_1086,N_670,N_843);
xnor U1087 (N_1087,N_750,N_795);
nor U1088 (N_1088,N_870,N_646);
nand U1089 (N_1089,N_630,N_660);
nand U1090 (N_1090,N_717,N_517);
nand U1091 (N_1091,N_565,N_537);
nor U1092 (N_1092,N_999,N_693);
and U1093 (N_1093,N_659,N_974);
or U1094 (N_1094,N_802,N_733);
nor U1095 (N_1095,N_890,N_635);
or U1096 (N_1096,N_835,N_874);
or U1097 (N_1097,N_757,N_539);
and U1098 (N_1098,N_538,N_697);
and U1099 (N_1099,N_811,N_963);
xnor U1100 (N_1100,N_596,N_764);
or U1101 (N_1101,N_544,N_731);
nand U1102 (N_1102,N_633,N_625);
and U1103 (N_1103,N_579,N_936);
or U1104 (N_1104,N_671,N_734);
nand U1105 (N_1105,N_657,N_573);
nor U1106 (N_1106,N_969,N_831);
or U1107 (N_1107,N_569,N_872);
nor U1108 (N_1108,N_711,N_956);
xor U1109 (N_1109,N_973,N_604);
nor U1110 (N_1110,N_680,N_878);
or U1111 (N_1111,N_566,N_824);
nor U1112 (N_1112,N_805,N_700);
nand U1113 (N_1113,N_737,N_873);
nand U1114 (N_1114,N_858,N_559);
nor U1115 (N_1115,N_922,N_692);
and U1116 (N_1116,N_987,N_946);
nor U1117 (N_1117,N_799,N_594);
and U1118 (N_1118,N_836,N_926);
xnor U1119 (N_1119,N_638,N_642);
and U1120 (N_1120,N_798,N_588);
nor U1121 (N_1121,N_949,N_546);
nor U1122 (N_1122,N_653,N_816);
nand U1123 (N_1123,N_570,N_901);
xnor U1124 (N_1124,N_839,N_655);
or U1125 (N_1125,N_515,N_608);
xnor U1126 (N_1126,N_679,N_781);
nor U1127 (N_1127,N_527,N_988);
and U1128 (N_1128,N_648,N_560);
and U1129 (N_1129,N_743,N_652);
nor U1130 (N_1130,N_989,N_714);
nor U1131 (N_1131,N_557,N_540);
or U1132 (N_1132,N_777,N_955);
nor U1133 (N_1133,N_605,N_932);
or U1134 (N_1134,N_895,N_518);
or U1135 (N_1135,N_553,N_736);
nand U1136 (N_1136,N_864,N_613);
xnor U1137 (N_1137,N_716,N_845);
nor U1138 (N_1138,N_848,N_662);
nor U1139 (N_1139,N_886,N_940);
and U1140 (N_1140,N_552,N_529);
or U1141 (N_1141,N_511,N_856);
nor U1142 (N_1142,N_615,N_695);
xnor U1143 (N_1143,N_674,N_751);
or U1144 (N_1144,N_871,N_943);
and U1145 (N_1145,N_767,N_586);
or U1146 (N_1146,N_822,N_543);
nand U1147 (N_1147,N_819,N_954);
and U1148 (N_1148,N_970,N_607);
nor U1149 (N_1149,N_792,N_892);
and U1150 (N_1150,N_500,N_727);
and U1151 (N_1151,N_724,N_541);
xnor U1152 (N_1152,N_574,N_791);
and U1153 (N_1153,N_643,N_661);
nand U1154 (N_1154,N_939,N_650);
nor U1155 (N_1155,N_888,N_884);
or U1156 (N_1156,N_961,N_686);
nor U1157 (N_1157,N_597,N_937);
and U1158 (N_1158,N_514,N_712);
or U1159 (N_1159,N_809,N_665);
nor U1160 (N_1160,N_564,N_948);
or U1161 (N_1161,N_827,N_705);
nand U1162 (N_1162,N_977,N_701);
and U1163 (N_1163,N_924,N_707);
nor U1164 (N_1164,N_723,N_753);
and U1165 (N_1165,N_842,N_855);
or U1166 (N_1166,N_567,N_929);
xor U1167 (N_1167,N_745,N_996);
and U1168 (N_1168,N_820,N_907);
or U1169 (N_1169,N_722,N_558);
or U1170 (N_1170,N_818,N_763);
and U1171 (N_1171,N_520,N_632);
and U1172 (N_1172,N_796,N_620);
nand U1173 (N_1173,N_585,N_964);
nand U1174 (N_1174,N_980,N_841);
and U1175 (N_1175,N_832,N_905);
nand U1176 (N_1176,N_691,N_730);
and U1177 (N_1177,N_698,N_528);
or U1178 (N_1178,N_704,N_899);
and U1179 (N_1179,N_636,N_958);
nand U1180 (N_1180,N_755,N_526);
nor U1181 (N_1181,N_793,N_840);
nand U1182 (N_1182,N_838,N_649);
nor U1183 (N_1183,N_976,N_854);
nand U1184 (N_1184,N_779,N_814);
or U1185 (N_1185,N_941,N_507);
nor U1186 (N_1186,N_952,N_813);
or U1187 (N_1187,N_729,N_664);
or U1188 (N_1188,N_885,N_990);
or U1189 (N_1189,N_582,N_561);
or U1190 (N_1190,N_690,N_797);
nand U1191 (N_1191,N_612,N_513);
and U1192 (N_1192,N_590,N_826);
xor U1193 (N_1193,N_994,N_812);
and U1194 (N_1194,N_720,N_869);
nor U1195 (N_1195,N_800,N_523);
xor U1196 (N_1196,N_681,N_617);
or U1197 (N_1197,N_912,N_725);
and U1198 (N_1198,N_696,N_978);
or U1199 (N_1199,N_790,N_718);
and U1200 (N_1200,N_889,N_715);
xnor U1201 (N_1201,N_902,N_788);
xnor U1202 (N_1202,N_754,N_891);
nand U1203 (N_1203,N_738,N_893);
or U1204 (N_1204,N_817,N_982);
and U1205 (N_1205,N_773,N_555);
and U1206 (N_1206,N_522,N_898);
and U1207 (N_1207,N_524,N_828);
nand U1208 (N_1208,N_916,N_732);
or U1209 (N_1209,N_626,N_682);
nor U1210 (N_1210,N_896,N_758);
or U1211 (N_1211,N_962,N_997);
nand U1212 (N_1212,N_580,N_521);
and U1213 (N_1213,N_741,N_595);
xnor U1214 (N_1214,N_887,N_953);
or U1215 (N_1215,N_687,N_622);
nand U1216 (N_1216,N_857,N_508);
nand U1217 (N_1217,N_894,N_900);
nor U1218 (N_1218,N_624,N_877);
nand U1219 (N_1219,N_834,N_778);
xnor U1220 (N_1220,N_710,N_776);
or U1221 (N_1221,N_785,N_806);
nor U1222 (N_1222,N_739,N_688);
or U1223 (N_1223,N_631,N_830);
nand U1224 (N_1224,N_875,N_505);
nor U1225 (N_1225,N_550,N_879);
and U1226 (N_1226,N_601,N_623);
nor U1227 (N_1227,N_709,N_993);
nand U1228 (N_1228,N_923,N_866);
nor U1229 (N_1229,N_549,N_859);
nand U1230 (N_1230,N_545,N_616);
and U1231 (N_1231,N_765,N_959);
or U1232 (N_1232,N_578,N_599);
nor U1233 (N_1233,N_865,N_547);
nand U1234 (N_1234,N_536,N_783);
or U1235 (N_1235,N_684,N_981);
and U1236 (N_1236,N_995,N_925);
nor U1237 (N_1237,N_913,N_931);
xnor U1238 (N_1238,N_957,N_784);
or U1239 (N_1239,N_609,N_911);
nor U1240 (N_1240,N_584,N_667);
or U1241 (N_1241,N_804,N_803);
nand U1242 (N_1242,N_915,N_794);
xnor U1243 (N_1243,N_568,N_749);
nand U1244 (N_1244,N_610,N_516);
xor U1245 (N_1245,N_512,N_772);
nor U1246 (N_1246,N_903,N_618);
nor U1247 (N_1247,N_908,N_823);
and U1248 (N_1248,N_852,N_656);
nand U1249 (N_1249,N_678,N_502);
nand U1250 (N_1250,N_980,N_800);
and U1251 (N_1251,N_685,N_599);
or U1252 (N_1252,N_983,N_672);
nand U1253 (N_1253,N_771,N_722);
and U1254 (N_1254,N_525,N_845);
nor U1255 (N_1255,N_694,N_701);
and U1256 (N_1256,N_723,N_669);
nor U1257 (N_1257,N_556,N_625);
and U1258 (N_1258,N_979,N_786);
or U1259 (N_1259,N_678,N_551);
or U1260 (N_1260,N_803,N_770);
nor U1261 (N_1261,N_905,N_638);
or U1262 (N_1262,N_855,N_802);
and U1263 (N_1263,N_610,N_543);
or U1264 (N_1264,N_614,N_864);
and U1265 (N_1265,N_970,N_688);
or U1266 (N_1266,N_817,N_723);
xnor U1267 (N_1267,N_541,N_736);
and U1268 (N_1268,N_717,N_753);
or U1269 (N_1269,N_567,N_788);
nor U1270 (N_1270,N_968,N_613);
xor U1271 (N_1271,N_894,N_744);
or U1272 (N_1272,N_511,N_939);
or U1273 (N_1273,N_712,N_509);
or U1274 (N_1274,N_623,N_966);
xor U1275 (N_1275,N_940,N_760);
xnor U1276 (N_1276,N_926,N_604);
nor U1277 (N_1277,N_517,N_546);
nor U1278 (N_1278,N_784,N_949);
and U1279 (N_1279,N_877,N_645);
or U1280 (N_1280,N_500,N_868);
and U1281 (N_1281,N_795,N_545);
nor U1282 (N_1282,N_901,N_527);
and U1283 (N_1283,N_808,N_610);
or U1284 (N_1284,N_733,N_904);
nand U1285 (N_1285,N_738,N_901);
and U1286 (N_1286,N_765,N_733);
or U1287 (N_1287,N_978,N_849);
and U1288 (N_1288,N_531,N_790);
or U1289 (N_1289,N_829,N_857);
and U1290 (N_1290,N_875,N_850);
nand U1291 (N_1291,N_988,N_829);
or U1292 (N_1292,N_785,N_852);
and U1293 (N_1293,N_816,N_557);
nand U1294 (N_1294,N_624,N_508);
xnor U1295 (N_1295,N_856,N_547);
nor U1296 (N_1296,N_689,N_914);
nor U1297 (N_1297,N_774,N_601);
nor U1298 (N_1298,N_770,N_912);
nor U1299 (N_1299,N_944,N_501);
nand U1300 (N_1300,N_582,N_675);
and U1301 (N_1301,N_694,N_581);
xor U1302 (N_1302,N_540,N_946);
nand U1303 (N_1303,N_687,N_681);
nand U1304 (N_1304,N_947,N_868);
and U1305 (N_1305,N_578,N_648);
nor U1306 (N_1306,N_832,N_771);
or U1307 (N_1307,N_655,N_660);
or U1308 (N_1308,N_950,N_835);
or U1309 (N_1309,N_813,N_627);
or U1310 (N_1310,N_677,N_706);
nor U1311 (N_1311,N_928,N_582);
nand U1312 (N_1312,N_624,N_534);
and U1313 (N_1313,N_831,N_838);
and U1314 (N_1314,N_817,N_865);
nor U1315 (N_1315,N_983,N_862);
and U1316 (N_1316,N_740,N_947);
or U1317 (N_1317,N_848,N_937);
and U1318 (N_1318,N_523,N_758);
and U1319 (N_1319,N_552,N_786);
nor U1320 (N_1320,N_702,N_911);
nor U1321 (N_1321,N_502,N_772);
nor U1322 (N_1322,N_892,N_606);
or U1323 (N_1323,N_524,N_706);
xor U1324 (N_1324,N_751,N_581);
or U1325 (N_1325,N_558,N_871);
and U1326 (N_1326,N_789,N_919);
or U1327 (N_1327,N_589,N_976);
nand U1328 (N_1328,N_542,N_580);
or U1329 (N_1329,N_950,N_871);
and U1330 (N_1330,N_675,N_507);
nand U1331 (N_1331,N_994,N_899);
or U1332 (N_1332,N_632,N_620);
and U1333 (N_1333,N_994,N_763);
xnor U1334 (N_1334,N_672,N_971);
and U1335 (N_1335,N_882,N_869);
xor U1336 (N_1336,N_512,N_791);
and U1337 (N_1337,N_858,N_705);
and U1338 (N_1338,N_594,N_868);
nand U1339 (N_1339,N_810,N_962);
and U1340 (N_1340,N_885,N_642);
nand U1341 (N_1341,N_610,N_600);
and U1342 (N_1342,N_990,N_505);
or U1343 (N_1343,N_878,N_641);
or U1344 (N_1344,N_800,N_848);
xor U1345 (N_1345,N_687,N_662);
nand U1346 (N_1346,N_824,N_764);
and U1347 (N_1347,N_843,N_569);
nand U1348 (N_1348,N_816,N_554);
nand U1349 (N_1349,N_780,N_698);
xnor U1350 (N_1350,N_548,N_774);
xnor U1351 (N_1351,N_904,N_698);
or U1352 (N_1352,N_777,N_638);
nand U1353 (N_1353,N_878,N_964);
nor U1354 (N_1354,N_942,N_695);
and U1355 (N_1355,N_787,N_744);
or U1356 (N_1356,N_861,N_608);
nor U1357 (N_1357,N_680,N_651);
nor U1358 (N_1358,N_696,N_610);
nand U1359 (N_1359,N_807,N_675);
and U1360 (N_1360,N_657,N_805);
or U1361 (N_1361,N_955,N_519);
nand U1362 (N_1362,N_887,N_986);
nand U1363 (N_1363,N_792,N_551);
nor U1364 (N_1364,N_938,N_522);
or U1365 (N_1365,N_813,N_743);
and U1366 (N_1366,N_884,N_828);
nor U1367 (N_1367,N_988,N_901);
nor U1368 (N_1368,N_869,N_793);
or U1369 (N_1369,N_906,N_763);
nor U1370 (N_1370,N_652,N_547);
and U1371 (N_1371,N_994,N_609);
or U1372 (N_1372,N_627,N_922);
and U1373 (N_1373,N_866,N_766);
or U1374 (N_1374,N_733,N_986);
and U1375 (N_1375,N_943,N_898);
nand U1376 (N_1376,N_611,N_995);
or U1377 (N_1377,N_791,N_675);
nand U1378 (N_1378,N_890,N_818);
nand U1379 (N_1379,N_812,N_888);
and U1380 (N_1380,N_896,N_829);
nor U1381 (N_1381,N_985,N_768);
and U1382 (N_1382,N_695,N_765);
nor U1383 (N_1383,N_858,N_766);
or U1384 (N_1384,N_945,N_511);
or U1385 (N_1385,N_598,N_519);
or U1386 (N_1386,N_684,N_908);
nand U1387 (N_1387,N_965,N_682);
and U1388 (N_1388,N_604,N_771);
xor U1389 (N_1389,N_967,N_507);
and U1390 (N_1390,N_651,N_892);
xor U1391 (N_1391,N_621,N_886);
nor U1392 (N_1392,N_928,N_793);
or U1393 (N_1393,N_663,N_610);
or U1394 (N_1394,N_678,N_973);
nor U1395 (N_1395,N_816,N_779);
or U1396 (N_1396,N_850,N_614);
or U1397 (N_1397,N_968,N_771);
nor U1398 (N_1398,N_914,N_590);
nor U1399 (N_1399,N_650,N_968);
nor U1400 (N_1400,N_523,N_560);
nand U1401 (N_1401,N_702,N_574);
nand U1402 (N_1402,N_842,N_646);
and U1403 (N_1403,N_739,N_635);
and U1404 (N_1404,N_558,N_940);
nand U1405 (N_1405,N_530,N_911);
and U1406 (N_1406,N_518,N_745);
nand U1407 (N_1407,N_686,N_517);
nand U1408 (N_1408,N_693,N_818);
nand U1409 (N_1409,N_905,N_643);
nor U1410 (N_1410,N_589,N_749);
or U1411 (N_1411,N_715,N_834);
and U1412 (N_1412,N_842,N_760);
xnor U1413 (N_1413,N_625,N_863);
and U1414 (N_1414,N_965,N_743);
xnor U1415 (N_1415,N_682,N_554);
nand U1416 (N_1416,N_755,N_938);
nor U1417 (N_1417,N_545,N_687);
xor U1418 (N_1418,N_536,N_742);
and U1419 (N_1419,N_817,N_584);
nand U1420 (N_1420,N_771,N_869);
and U1421 (N_1421,N_606,N_508);
nand U1422 (N_1422,N_908,N_596);
nand U1423 (N_1423,N_664,N_735);
or U1424 (N_1424,N_836,N_545);
nor U1425 (N_1425,N_904,N_884);
xnor U1426 (N_1426,N_911,N_699);
nand U1427 (N_1427,N_905,N_535);
and U1428 (N_1428,N_788,N_735);
xnor U1429 (N_1429,N_786,N_532);
or U1430 (N_1430,N_579,N_637);
and U1431 (N_1431,N_871,N_772);
nand U1432 (N_1432,N_557,N_802);
nor U1433 (N_1433,N_781,N_682);
and U1434 (N_1434,N_808,N_733);
and U1435 (N_1435,N_900,N_715);
nor U1436 (N_1436,N_547,N_686);
and U1437 (N_1437,N_946,N_900);
nand U1438 (N_1438,N_562,N_761);
and U1439 (N_1439,N_788,N_819);
nand U1440 (N_1440,N_667,N_960);
and U1441 (N_1441,N_567,N_999);
nand U1442 (N_1442,N_615,N_988);
and U1443 (N_1443,N_628,N_796);
nand U1444 (N_1444,N_773,N_910);
xnor U1445 (N_1445,N_550,N_547);
or U1446 (N_1446,N_807,N_828);
nor U1447 (N_1447,N_821,N_839);
or U1448 (N_1448,N_945,N_618);
nand U1449 (N_1449,N_729,N_988);
or U1450 (N_1450,N_720,N_724);
nor U1451 (N_1451,N_947,N_842);
nand U1452 (N_1452,N_608,N_684);
nor U1453 (N_1453,N_576,N_682);
xnor U1454 (N_1454,N_683,N_903);
or U1455 (N_1455,N_813,N_912);
nand U1456 (N_1456,N_540,N_858);
nand U1457 (N_1457,N_563,N_626);
nand U1458 (N_1458,N_813,N_983);
and U1459 (N_1459,N_874,N_729);
nor U1460 (N_1460,N_732,N_663);
nor U1461 (N_1461,N_726,N_584);
xnor U1462 (N_1462,N_830,N_867);
nor U1463 (N_1463,N_506,N_592);
nand U1464 (N_1464,N_726,N_524);
nand U1465 (N_1465,N_846,N_631);
nand U1466 (N_1466,N_593,N_731);
or U1467 (N_1467,N_851,N_779);
or U1468 (N_1468,N_845,N_674);
xor U1469 (N_1469,N_617,N_604);
nor U1470 (N_1470,N_501,N_540);
nand U1471 (N_1471,N_636,N_730);
or U1472 (N_1472,N_785,N_828);
nor U1473 (N_1473,N_798,N_538);
nand U1474 (N_1474,N_945,N_541);
nand U1475 (N_1475,N_727,N_864);
xor U1476 (N_1476,N_669,N_545);
nor U1477 (N_1477,N_536,N_502);
nor U1478 (N_1478,N_700,N_554);
xnor U1479 (N_1479,N_818,N_976);
nand U1480 (N_1480,N_591,N_681);
or U1481 (N_1481,N_602,N_709);
and U1482 (N_1482,N_893,N_841);
and U1483 (N_1483,N_503,N_917);
nor U1484 (N_1484,N_711,N_836);
and U1485 (N_1485,N_817,N_591);
or U1486 (N_1486,N_552,N_871);
or U1487 (N_1487,N_610,N_592);
or U1488 (N_1488,N_946,N_807);
or U1489 (N_1489,N_741,N_754);
and U1490 (N_1490,N_744,N_838);
or U1491 (N_1491,N_819,N_554);
or U1492 (N_1492,N_522,N_562);
and U1493 (N_1493,N_625,N_844);
and U1494 (N_1494,N_764,N_531);
nand U1495 (N_1495,N_875,N_996);
nor U1496 (N_1496,N_618,N_968);
and U1497 (N_1497,N_969,N_525);
or U1498 (N_1498,N_582,N_709);
nand U1499 (N_1499,N_988,N_617);
or U1500 (N_1500,N_1042,N_1378);
nor U1501 (N_1501,N_1390,N_1293);
xor U1502 (N_1502,N_1387,N_1000);
or U1503 (N_1503,N_1284,N_1489);
or U1504 (N_1504,N_1356,N_1246);
and U1505 (N_1505,N_1324,N_1287);
xor U1506 (N_1506,N_1054,N_1288);
and U1507 (N_1507,N_1447,N_1277);
nand U1508 (N_1508,N_1100,N_1337);
nand U1509 (N_1509,N_1112,N_1001);
nor U1510 (N_1510,N_1189,N_1087);
and U1511 (N_1511,N_1104,N_1401);
nand U1512 (N_1512,N_1304,N_1197);
and U1513 (N_1513,N_1340,N_1279);
nand U1514 (N_1514,N_1400,N_1116);
nor U1515 (N_1515,N_1039,N_1363);
or U1516 (N_1516,N_1011,N_1081);
and U1517 (N_1517,N_1017,N_1265);
nand U1518 (N_1518,N_1088,N_1498);
and U1519 (N_1519,N_1089,N_1052);
nor U1520 (N_1520,N_1426,N_1470);
nand U1521 (N_1521,N_1151,N_1394);
or U1522 (N_1522,N_1022,N_1380);
or U1523 (N_1523,N_1172,N_1347);
nor U1524 (N_1524,N_1077,N_1484);
or U1525 (N_1525,N_1275,N_1407);
or U1526 (N_1526,N_1019,N_1259);
nand U1527 (N_1527,N_1384,N_1434);
or U1528 (N_1528,N_1360,N_1067);
nand U1529 (N_1529,N_1374,N_1111);
and U1530 (N_1530,N_1469,N_1428);
xnor U1531 (N_1531,N_1243,N_1226);
xor U1532 (N_1532,N_1136,N_1405);
and U1533 (N_1533,N_1313,N_1154);
or U1534 (N_1534,N_1205,N_1063);
xnor U1535 (N_1535,N_1494,N_1131);
nor U1536 (N_1536,N_1412,N_1015);
nand U1537 (N_1537,N_1072,N_1093);
xnor U1538 (N_1538,N_1451,N_1429);
or U1539 (N_1539,N_1149,N_1179);
nor U1540 (N_1540,N_1106,N_1186);
xor U1541 (N_1541,N_1200,N_1033);
nor U1542 (N_1542,N_1289,N_1075);
nand U1543 (N_1543,N_1098,N_1233);
nand U1544 (N_1544,N_1472,N_1268);
xor U1545 (N_1545,N_1158,N_1252);
nor U1546 (N_1546,N_1345,N_1209);
and U1547 (N_1547,N_1457,N_1124);
xor U1548 (N_1548,N_1182,N_1016);
and U1549 (N_1549,N_1148,N_1406);
nand U1550 (N_1550,N_1397,N_1121);
nor U1551 (N_1551,N_1109,N_1296);
nand U1552 (N_1552,N_1456,N_1485);
nand U1553 (N_1553,N_1163,N_1481);
or U1554 (N_1554,N_1291,N_1257);
and U1555 (N_1555,N_1091,N_1160);
nand U1556 (N_1556,N_1239,N_1222);
nor U1557 (N_1557,N_1278,N_1329);
or U1558 (N_1558,N_1495,N_1213);
nand U1559 (N_1559,N_1008,N_1351);
or U1560 (N_1560,N_1312,N_1263);
nor U1561 (N_1561,N_1006,N_1129);
and U1562 (N_1562,N_1343,N_1333);
nand U1563 (N_1563,N_1143,N_1388);
nand U1564 (N_1564,N_1079,N_1188);
nand U1565 (N_1565,N_1009,N_1013);
nor U1566 (N_1566,N_1153,N_1332);
or U1567 (N_1567,N_1235,N_1286);
or U1568 (N_1568,N_1492,N_1310);
nor U1569 (N_1569,N_1432,N_1454);
nor U1570 (N_1570,N_1027,N_1326);
xnor U1571 (N_1571,N_1038,N_1414);
and U1572 (N_1572,N_1021,N_1114);
nor U1573 (N_1573,N_1375,N_1377);
or U1574 (N_1574,N_1224,N_1024);
and U1575 (N_1575,N_1411,N_1191);
nand U1576 (N_1576,N_1193,N_1463);
nand U1577 (N_1577,N_1364,N_1036);
and U1578 (N_1578,N_1371,N_1146);
xor U1579 (N_1579,N_1105,N_1295);
xor U1580 (N_1580,N_1242,N_1167);
and U1581 (N_1581,N_1330,N_1493);
or U1582 (N_1582,N_1315,N_1477);
and U1583 (N_1583,N_1344,N_1141);
and U1584 (N_1584,N_1491,N_1165);
or U1585 (N_1585,N_1464,N_1073);
or U1586 (N_1586,N_1236,N_1095);
or U1587 (N_1587,N_1183,N_1399);
xor U1588 (N_1588,N_1455,N_1386);
and U1589 (N_1589,N_1218,N_1458);
and U1590 (N_1590,N_1176,N_1338);
nand U1591 (N_1591,N_1264,N_1096);
xor U1592 (N_1592,N_1012,N_1497);
nand U1593 (N_1593,N_1444,N_1061);
or U1594 (N_1594,N_1418,N_1297);
or U1595 (N_1595,N_1474,N_1299);
nor U1596 (N_1596,N_1083,N_1427);
and U1597 (N_1597,N_1478,N_1415);
and U1598 (N_1598,N_1194,N_1108);
and U1599 (N_1599,N_1119,N_1357);
xor U1600 (N_1600,N_1408,N_1228);
or U1601 (N_1601,N_1223,N_1225);
and U1602 (N_1602,N_1334,N_1281);
and U1603 (N_1603,N_1342,N_1068);
nor U1604 (N_1604,N_1180,N_1041);
nand U1605 (N_1605,N_1385,N_1331);
or U1606 (N_1606,N_1328,N_1206);
xnor U1607 (N_1607,N_1247,N_1169);
or U1608 (N_1608,N_1102,N_1272);
nand U1609 (N_1609,N_1483,N_1271);
xnor U1610 (N_1610,N_1241,N_1441);
nand U1611 (N_1611,N_1320,N_1175);
or U1612 (N_1612,N_1488,N_1060);
or U1613 (N_1613,N_1285,N_1190);
or U1614 (N_1614,N_1227,N_1035);
nand U1615 (N_1615,N_1306,N_1361);
or U1616 (N_1616,N_1202,N_1322);
xnor U1617 (N_1617,N_1048,N_1201);
xnor U1618 (N_1618,N_1379,N_1362);
or U1619 (N_1619,N_1250,N_1499);
nor U1620 (N_1620,N_1448,N_1480);
and U1621 (N_1621,N_1311,N_1181);
or U1622 (N_1622,N_1398,N_1443);
nand U1623 (N_1623,N_1391,N_1425);
or U1624 (N_1624,N_1350,N_1062);
and U1625 (N_1625,N_1014,N_1269);
nor U1626 (N_1626,N_1486,N_1309);
nand U1627 (N_1627,N_1402,N_1118);
and U1628 (N_1628,N_1128,N_1099);
xnor U1629 (N_1629,N_1382,N_1107);
nor U1630 (N_1630,N_1438,N_1171);
nand U1631 (N_1631,N_1248,N_1487);
nand U1632 (N_1632,N_1335,N_1249);
nor U1633 (N_1633,N_1450,N_1198);
nor U1634 (N_1634,N_1221,N_1260);
and U1635 (N_1635,N_1170,N_1300);
and U1636 (N_1636,N_1086,N_1056);
nand U1637 (N_1637,N_1040,N_1092);
nor U1638 (N_1638,N_1349,N_1409);
and U1639 (N_1639,N_1173,N_1307);
nand U1640 (N_1640,N_1126,N_1254);
nand U1641 (N_1641,N_1471,N_1396);
xor U1642 (N_1642,N_1220,N_1135);
or U1643 (N_1643,N_1211,N_1025);
nand U1644 (N_1644,N_1032,N_1234);
or U1645 (N_1645,N_1103,N_1034);
or U1646 (N_1646,N_1381,N_1187);
nand U1647 (N_1647,N_1047,N_1436);
or U1648 (N_1648,N_1231,N_1274);
and U1649 (N_1649,N_1256,N_1403);
or U1650 (N_1650,N_1080,N_1139);
nor U1651 (N_1651,N_1157,N_1317);
and U1652 (N_1652,N_1442,N_1431);
xnor U1653 (N_1653,N_1479,N_1413);
nor U1654 (N_1654,N_1301,N_1440);
or U1655 (N_1655,N_1207,N_1159);
nor U1656 (N_1656,N_1298,N_1290);
or U1657 (N_1657,N_1185,N_1475);
nand U1658 (N_1658,N_1057,N_1461);
or U1659 (N_1659,N_1162,N_1476);
nand U1660 (N_1660,N_1430,N_1245);
and U1661 (N_1661,N_1283,N_1370);
nand U1662 (N_1662,N_1417,N_1294);
nand U1663 (N_1663,N_1037,N_1420);
nand U1664 (N_1664,N_1076,N_1150);
nand U1665 (N_1665,N_1416,N_1123);
nand U1666 (N_1666,N_1184,N_1002);
nand U1667 (N_1667,N_1439,N_1134);
and U1668 (N_1668,N_1028,N_1168);
and U1669 (N_1669,N_1318,N_1467);
nor U1670 (N_1670,N_1051,N_1145);
nand U1671 (N_1671,N_1140,N_1496);
or U1672 (N_1672,N_1459,N_1064);
and U1673 (N_1673,N_1059,N_1266);
nand U1674 (N_1674,N_1152,N_1353);
nor U1675 (N_1675,N_1452,N_1043);
or U1676 (N_1676,N_1336,N_1237);
xor U1677 (N_1677,N_1422,N_1070);
xor U1678 (N_1678,N_1346,N_1280);
nand U1679 (N_1679,N_1319,N_1367);
or U1680 (N_1680,N_1466,N_1262);
and U1681 (N_1681,N_1214,N_1462);
nor U1682 (N_1682,N_1066,N_1195);
or U1683 (N_1683,N_1004,N_1046);
nor U1684 (N_1684,N_1435,N_1327);
xor U1685 (N_1685,N_1174,N_1437);
nor U1686 (N_1686,N_1069,N_1449);
and U1687 (N_1687,N_1473,N_1115);
nand U1688 (N_1688,N_1164,N_1065);
or U1689 (N_1689,N_1208,N_1389);
nand U1690 (N_1690,N_1058,N_1196);
nor U1691 (N_1691,N_1270,N_1120);
and U1692 (N_1692,N_1210,N_1354);
or U1693 (N_1693,N_1085,N_1003);
nand U1694 (N_1694,N_1192,N_1352);
nor U1695 (N_1695,N_1005,N_1433);
nand U1696 (N_1696,N_1465,N_1314);
xnor U1697 (N_1697,N_1078,N_1240);
nand U1698 (N_1698,N_1468,N_1122);
and U1699 (N_1699,N_1178,N_1097);
nand U1700 (N_1700,N_1177,N_1445);
nand U1701 (N_1701,N_1010,N_1339);
and U1702 (N_1702,N_1216,N_1359);
nand U1703 (N_1703,N_1018,N_1316);
nand U1704 (N_1704,N_1090,N_1023);
nand U1705 (N_1705,N_1204,N_1212);
or U1706 (N_1706,N_1215,N_1376);
nand U1707 (N_1707,N_1082,N_1421);
xor U1708 (N_1708,N_1155,N_1253);
nor U1709 (N_1709,N_1026,N_1020);
nor U1710 (N_1710,N_1302,N_1325);
nand U1711 (N_1711,N_1138,N_1045);
nand U1712 (N_1712,N_1094,N_1238);
xor U1713 (N_1713,N_1273,N_1303);
or U1714 (N_1714,N_1460,N_1229);
xor U1715 (N_1715,N_1244,N_1282);
xor U1716 (N_1716,N_1410,N_1232);
nand U1717 (N_1717,N_1292,N_1369);
nand U1718 (N_1718,N_1419,N_1117);
nor U1719 (N_1719,N_1358,N_1323);
and U1720 (N_1720,N_1161,N_1084);
xnor U1721 (N_1721,N_1276,N_1137);
nor U1722 (N_1722,N_1044,N_1258);
nand U1723 (N_1723,N_1393,N_1395);
and U1724 (N_1724,N_1490,N_1203);
or U1725 (N_1725,N_1130,N_1365);
or U1726 (N_1726,N_1255,N_1308);
xnor U1727 (N_1727,N_1341,N_1132);
and U1728 (N_1728,N_1368,N_1142);
or U1729 (N_1729,N_1113,N_1219);
or U1730 (N_1730,N_1404,N_1348);
nor U1731 (N_1731,N_1355,N_1007);
and U1732 (N_1732,N_1049,N_1446);
or U1733 (N_1733,N_1031,N_1030);
nand U1734 (N_1734,N_1424,N_1392);
nor U1735 (N_1735,N_1321,N_1110);
nand U1736 (N_1736,N_1053,N_1230);
nand U1737 (N_1737,N_1125,N_1050);
and U1738 (N_1738,N_1156,N_1029);
nor U1739 (N_1739,N_1482,N_1366);
nor U1740 (N_1740,N_1217,N_1133);
nand U1741 (N_1741,N_1101,N_1372);
or U1742 (N_1742,N_1127,N_1074);
nor U1743 (N_1743,N_1251,N_1261);
nand U1744 (N_1744,N_1144,N_1453);
or U1745 (N_1745,N_1055,N_1305);
and U1746 (N_1746,N_1166,N_1267);
nand U1747 (N_1747,N_1423,N_1071);
nand U1748 (N_1748,N_1147,N_1383);
or U1749 (N_1749,N_1373,N_1199);
xor U1750 (N_1750,N_1093,N_1245);
nor U1751 (N_1751,N_1282,N_1298);
or U1752 (N_1752,N_1340,N_1261);
and U1753 (N_1753,N_1485,N_1165);
nand U1754 (N_1754,N_1365,N_1183);
or U1755 (N_1755,N_1245,N_1330);
or U1756 (N_1756,N_1354,N_1398);
nor U1757 (N_1757,N_1381,N_1380);
nand U1758 (N_1758,N_1111,N_1461);
or U1759 (N_1759,N_1149,N_1001);
nand U1760 (N_1760,N_1310,N_1251);
xnor U1761 (N_1761,N_1470,N_1408);
nor U1762 (N_1762,N_1450,N_1184);
or U1763 (N_1763,N_1117,N_1142);
xnor U1764 (N_1764,N_1420,N_1246);
and U1765 (N_1765,N_1368,N_1216);
and U1766 (N_1766,N_1384,N_1389);
nand U1767 (N_1767,N_1280,N_1037);
and U1768 (N_1768,N_1201,N_1250);
nand U1769 (N_1769,N_1429,N_1456);
nor U1770 (N_1770,N_1316,N_1466);
or U1771 (N_1771,N_1389,N_1110);
or U1772 (N_1772,N_1452,N_1156);
nand U1773 (N_1773,N_1456,N_1038);
and U1774 (N_1774,N_1401,N_1105);
or U1775 (N_1775,N_1131,N_1065);
xor U1776 (N_1776,N_1155,N_1165);
nand U1777 (N_1777,N_1408,N_1426);
nor U1778 (N_1778,N_1349,N_1249);
and U1779 (N_1779,N_1133,N_1235);
or U1780 (N_1780,N_1271,N_1085);
xnor U1781 (N_1781,N_1279,N_1446);
and U1782 (N_1782,N_1394,N_1385);
xor U1783 (N_1783,N_1460,N_1209);
nand U1784 (N_1784,N_1306,N_1330);
and U1785 (N_1785,N_1063,N_1198);
or U1786 (N_1786,N_1236,N_1255);
or U1787 (N_1787,N_1412,N_1182);
and U1788 (N_1788,N_1126,N_1263);
nor U1789 (N_1789,N_1288,N_1210);
and U1790 (N_1790,N_1370,N_1281);
nor U1791 (N_1791,N_1400,N_1396);
nand U1792 (N_1792,N_1092,N_1065);
nor U1793 (N_1793,N_1357,N_1309);
and U1794 (N_1794,N_1471,N_1065);
and U1795 (N_1795,N_1345,N_1088);
xor U1796 (N_1796,N_1466,N_1260);
nor U1797 (N_1797,N_1268,N_1025);
nand U1798 (N_1798,N_1471,N_1462);
nand U1799 (N_1799,N_1216,N_1296);
or U1800 (N_1800,N_1138,N_1422);
nand U1801 (N_1801,N_1376,N_1494);
nand U1802 (N_1802,N_1318,N_1026);
or U1803 (N_1803,N_1281,N_1449);
nand U1804 (N_1804,N_1115,N_1065);
nand U1805 (N_1805,N_1077,N_1215);
nor U1806 (N_1806,N_1347,N_1462);
or U1807 (N_1807,N_1349,N_1222);
nor U1808 (N_1808,N_1259,N_1027);
or U1809 (N_1809,N_1345,N_1025);
and U1810 (N_1810,N_1425,N_1098);
nor U1811 (N_1811,N_1356,N_1063);
or U1812 (N_1812,N_1475,N_1323);
nand U1813 (N_1813,N_1045,N_1306);
xor U1814 (N_1814,N_1430,N_1126);
xnor U1815 (N_1815,N_1043,N_1479);
xnor U1816 (N_1816,N_1344,N_1382);
or U1817 (N_1817,N_1360,N_1386);
nor U1818 (N_1818,N_1358,N_1134);
nand U1819 (N_1819,N_1177,N_1418);
or U1820 (N_1820,N_1195,N_1406);
or U1821 (N_1821,N_1057,N_1013);
or U1822 (N_1822,N_1275,N_1208);
nand U1823 (N_1823,N_1333,N_1429);
nand U1824 (N_1824,N_1410,N_1443);
and U1825 (N_1825,N_1049,N_1494);
nand U1826 (N_1826,N_1360,N_1117);
or U1827 (N_1827,N_1479,N_1213);
nor U1828 (N_1828,N_1112,N_1416);
xor U1829 (N_1829,N_1333,N_1021);
nor U1830 (N_1830,N_1497,N_1211);
and U1831 (N_1831,N_1249,N_1324);
and U1832 (N_1832,N_1377,N_1136);
or U1833 (N_1833,N_1156,N_1458);
nor U1834 (N_1834,N_1338,N_1392);
and U1835 (N_1835,N_1480,N_1196);
or U1836 (N_1836,N_1036,N_1039);
nor U1837 (N_1837,N_1124,N_1127);
and U1838 (N_1838,N_1444,N_1071);
nor U1839 (N_1839,N_1255,N_1453);
and U1840 (N_1840,N_1040,N_1214);
nand U1841 (N_1841,N_1450,N_1460);
nor U1842 (N_1842,N_1171,N_1136);
and U1843 (N_1843,N_1435,N_1300);
xor U1844 (N_1844,N_1470,N_1070);
and U1845 (N_1845,N_1435,N_1460);
or U1846 (N_1846,N_1098,N_1463);
or U1847 (N_1847,N_1478,N_1118);
and U1848 (N_1848,N_1259,N_1070);
and U1849 (N_1849,N_1043,N_1388);
or U1850 (N_1850,N_1357,N_1122);
and U1851 (N_1851,N_1151,N_1153);
or U1852 (N_1852,N_1042,N_1349);
nor U1853 (N_1853,N_1467,N_1052);
nor U1854 (N_1854,N_1053,N_1253);
and U1855 (N_1855,N_1439,N_1393);
or U1856 (N_1856,N_1115,N_1248);
xnor U1857 (N_1857,N_1332,N_1497);
nor U1858 (N_1858,N_1217,N_1130);
nand U1859 (N_1859,N_1285,N_1483);
or U1860 (N_1860,N_1144,N_1130);
nand U1861 (N_1861,N_1456,N_1281);
nand U1862 (N_1862,N_1150,N_1128);
and U1863 (N_1863,N_1475,N_1042);
and U1864 (N_1864,N_1231,N_1212);
or U1865 (N_1865,N_1243,N_1394);
or U1866 (N_1866,N_1164,N_1237);
or U1867 (N_1867,N_1464,N_1453);
nor U1868 (N_1868,N_1055,N_1008);
nand U1869 (N_1869,N_1494,N_1211);
or U1870 (N_1870,N_1385,N_1283);
nor U1871 (N_1871,N_1281,N_1199);
nand U1872 (N_1872,N_1175,N_1444);
nand U1873 (N_1873,N_1184,N_1253);
nand U1874 (N_1874,N_1185,N_1369);
nor U1875 (N_1875,N_1385,N_1461);
and U1876 (N_1876,N_1046,N_1201);
or U1877 (N_1877,N_1075,N_1046);
or U1878 (N_1878,N_1302,N_1018);
nor U1879 (N_1879,N_1256,N_1481);
or U1880 (N_1880,N_1294,N_1012);
or U1881 (N_1881,N_1244,N_1168);
xnor U1882 (N_1882,N_1147,N_1211);
nand U1883 (N_1883,N_1245,N_1293);
nor U1884 (N_1884,N_1457,N_1224);
or U1885 (N_1885,N_1306,N_1010);
xor U1886 (N_1886,N_1253,N_1137);
and U1887 (N_1887,N_1386,N_1218);
nor U1888 (N_1888,N_1092,N_1204);
xor U1889 (N_1889,N_1340,N_1262);
xor U1890 (N_1890,N_1015,N_1142);
or U1891 (N_1891,N_1308,N_1331);
nand U1892 (N_1892,N_1298,N_1463);
nand U1893 (N_1893,N_1361,N_1093);
nor U1894 (N_1894,N_1241,N_1427);
and U1895 (N_1895,N_1242,N_1440);
nand U1896 (N_1896,N_1255,N_1089);
nor U1897 (N_1897,N_1471,N_1289);
and U1898 (N_1898,N_1291,N_1288);
or U1899 (N_1899,N_1420,N_1228);
and U1900 (N_1900,N_1031,N_1449);
xor U1901 (N_1901,N_1391,N_1075);
and U1902 (N_1902,N_1324,N_1152);
and U1903 (N_1903,N_1057,N_1429);
or U1904 (N_1904,N_1183,N_1274);
or U1905 (N_1905,N_1367,N_1128);
or U1906 (N_1906,N_1369,N_1446);
nand U1907 (N_1907,N_1032,N_1405);
nand U1908 (N_1908,N_1146,N_1002);
or U1909 (N_1909,N_1083,N_1478);
nor U1910 (N_1910,N_1395,N_1384);
nor U1911 (N_1911,N_1134,N_1086);
nor U1912 (N_1912,N_1178,N_1154);
and U1913 (N_1913,N_1357,N_1469);
or U1914 (N_1914,N_1381,N_1499);
and U1915 (N_1915,N_1436,N_1182);
nand U1916 (N_1916,N_1092,N_1404);
or U1917 (N_1917,N_1423,N_1486);
xor U1918 (N_1918,N_1485,N_1152);
and U1919 (N_1919,N_1408,N_1274);
or U1920 (N_1920,N_1257,N_1194);
nand U1921 (N_1921,N_1265,N_1131);
xor U1922 (N_1922,N_1404,N_1151);
or U1923 (N_1923,N_1266,N_1495);
or U1924 (N_1924,N_1380,N_1326);
and U1925 (N_1925,N_1218,N_1318);
nand U1926 (N_1926,N_1010,N_1359);
nand U1927 (N_1927,N_1159,N_1196);
xnor U1928 (N_1928,N_1229,N_1191);
nor U1929 (N_1929,N_1098,N_1134);
nand U1930 (N_1930,N_1270,N_1195);
or U1931 (N_1931,N_1140,N_1108);
xor U1932 (N_1932,N_1337,N_1446);
nand U1933 (N_1933,N_1443,N_1257);
or U1934 (N_1934,N_1347,N_1129);
and U1935 (N_1935,N_1436,N_1126);
and U1936 (N_1936,N_1403,N_1425);
nand U1937 (N_1937,N_1250,N_1401);
or U1938 (N_1938,N_1036,N_1356);
and U1939 (N_1939,N_1007,N_1468);
and U1940 (N_1940,N_1469,N_1376);
nor U1941 (N_1941,N_1334,N_1144);
xor U1942 (N_1942,N_1471,N_1183);
and U1943 (N_1943,N_1169,N_1174);
and U1944 (N_1944,N_1134,N_1381);
nand U1945 (N_1945,N_1334,N_1459);
nand U1946 (N_1946,N_1043,N_1360);
nand U1947 (N_1947,N_1231,N_1227);
or U1948 (N_1948,N_1402,N_1454);
and U1949 (N_1949,N_1018,N_1391);
and U1950 (N_1950,N_1307,N_1162);
or U1951 (N_1951,N_1406,N_1096);
nand U1952 (N_1952,N_1472,N_1115);
nand U1953 (N_1953,N_1158,N_1281);
or U1954 (N_1954,N_1320,N_1439);
and U1955 (N_1955,N_1112,N_1240);
xor U1956 (N_1956,N_1428,N_1082);
nand U1957 (N_1957,N_1156,N_1406);
or U1958 (N_1958,N_1147,N_1269);
nor U1959 (N_1959,N_1252,N_1178);
or U1960 (N_1960,N_1023,N_1095);
nand U1961 (N_1961,N_1020,N_1411);
nand U1962 (N_1962,N_1061,N_1176);
or U1963 (N_1963,N_1185,N_1008);
or U1964 (N_1964,N_1481,N_1470);
and U1965 (N_1965,N_1320,N_1096);
nor U1966 (N_1966,N_1402,N_1327);
nand U1967 (N_1967,N_1157,N_1353);
xnor U1968 (N_1968,N_1003,N_1070);
nand U1969 (N_1969,N_1023,N_1136);
nor U1970 (N_1970,N_1342,N_1258);
nor U1971 (N_1971,N_1154,N_1465);
nor U1972 (N_1972,N_1008,N_1027);
xor U1973 (N_1973,N_1020,N_1395);
or U1974 (N_1974,N_1234,N_1463);
nand U1975 (N_1975,N_1321,N_1418);
nand U1976 (N_1976,N_1065,N_1287);
nor U1977 (N_1977,N_1431,N_1495);
or U1978 (N_1978,N_1307,N_1155);
xnor U1979 (N_1979,N_1193,N_1236);
xor U1980 (N_1980,N_1485,N_1449);
nor U1981 (N_1981,N_1459,N_1095);
nand U1982 (N_1982,N_1484,N_1141);
nand U1983 (N_1983,N_1040,N_1010);
or U1984 (N_1984,N_1016,N_1442);
and U1985 (N_1985,N_1043,N_1353);
or U1986 (N_1986,N_1494,N_1330);
or U1987 (N_1987,N_1291,N_1134);
and U1988 (N_1988,N_1287,N_1124);
and U1989 (N_1989,N_1131,N_1431);
nand U1990 (N_1990,N_1442,N_1186);
nor U1991 (N_1991,N_1407,N_1497);
nand U1992 (N_1992,N_1173,N_1245);
or U1993 (N_1993,N_1476,N_1313);
and U1994 (N_1994,N_1186,N_1359);
nor U1995 (N_1995,N_1295,N_1190);
nand U1996 (N_1996,N_1019,N_1271);
nand U1997 (N_1997,N_1422,N_1068);
or U1998 (N_1998,N_1248,N_1482);
nor U1999 (N_1999,N_1376,N_1307);
and U2000 (N_2000,N_1725,N_1893);
nor U2001 (N_2001,N_1779,N_1941);
nand U2002 (N_2002,N_1559,N_1795);
and U2003 (N_2003,N_1561,N_1562);
or U2004 (N_2004,N_1550,N_1657);
and U2005 (N_2005,N_1669,N_1913);
or U2006 (N_2006,N_1504,N_1810);
nand U2007 (N_2007,N_1843,N_1639);
and U2008 (N_2008,N_1993,N_1822);
nand U2009 (N_2009,N_1633,N_1876);
nand U2010 (N_2010,N_1741,N_1646);
nand U2011 (N_2011,N_1812,N_1645);
or U2012 (N_2012,N_1923,N_1611);
xnor U2013 (N_2013,N_1512,N_1994);
and U2014 (N_2014,N_1790,N_1684);
or U2015 (N_2015,N_1865,N_1794);
nand U2016 (N_2016,N_1612,N_1547);
nand U2017 (N_2017,N_1807,N_1863);
xnor U2018 (N_2018,N_1882,N_1797);
and U2019 (N_2019,N_1915,N_1723);
or U2020 (N_2020,N_1598,N_1596);
nor U2021 (N_2021,N_1903,N_1543);
and U2022 (N_2022,N_1511,N_1827);
or U2023 (N_2023,N_1638,N_1803);
nor U2024 (N_2024,N_1768,N_1883);
nor U2025 (N_2025,N_1658,N_1692);
nor U2026 (N_2026,N_1948,N_1837);
nor U2027 (N_2027,N_1718,N_1715);
and U2028 (N_2028,N_1744,N_1593);
or U2029 (N_2029,N_1588,N_1628);
and U2030 (N_2030,N_1592,N_1885);
xor U2031 (N_2031,N_1789,N_1686);
nand U2032 (N_2032,N_1517,N_1800);
nand U2033 (N_2033,N_1976,N_1866);
xor U2034 (N_2034,N_1745,N_1660);
nor U2035 (N_2035,N_1955,N_1548);
nor U2036 (N_2036,N_1506,N_1602);
or U2037 (N_2037,N_1533,N_1814);
and U2038 (N_2038,N_1652,N_1867);
or U2039 (N_2039,N_1960,N_1566);
or U2040 (N_2040,N_1930,N_1792);
or U2041 (N_2041,N_1966,N_1530);
nor U2042 (N_2042,N_1701,N_1653);
nand U2043 (N_2043,N_1514,N_1921);
nor U2044 (N_2044,N_1555,N_1574);
and U2045 (N_2045,N_1722,N_1809);
and U2046 (N_2046,N_1911,N_1989);
or U2047 (N_2047,N_1610,N_1580);
xor U2048 (N_2048,N_1661,N_1651);
nor U2049 (N_2049,N_1733,N_1697);
or U2050 (N_2050,N_1627,N_1799);
or U2051 (N_2051,N_1896,N_1900);
and U2052 (N_2052,N_1852,N_1636);
nor U2053 (N_2053,N_1939,N_1886);
or U2054 (N_2054,N_1750,N_1862);
and U2055 (N_2055,N_1920,N_1617);
or U2056 (N_2056,N_1600,N_1500);
nand U2057 (N_2057,N_1502,N_1683);
and U2058 (N_2058,N_1791,N_1844);
and U2059 (N_2059,N_1774,N_1678);
nand U2060 (N_2060,N_1631,N_1972);
and U2061 (N_2061,N_1990,N_1680);
nand U2062 (N_2062,N_1808,N_1614);
xnor U2063 (N_2063,N_1712,N_1772);
nand U2064 (N_2064,N_1674,N_1667);
or U2065 (N_2065,N_1553,N_1591);
nor U2066 (N_2066,N_1541,N_1713);
and U2067 (N_2067,N_1933,N_1594);
nor U2068 (N_2068,N_1938,N_1936);
nor U2069 (N_2069,N_1988,N_1520);
and U2070 (N_2070,N_1927,N_1558);
nor U2071 (N_2071,N_1872,N_1981);
nand U2072 (N_2072,N_1877,N_1889);
nor U2073 (N_2073,N_1606,N_1902);
nor U2074 (N_2074,N_1884,N_1782);
nand U2075 (N_2075,N_1690,N_1572);
nor U2076 (N_2076,N_1663,N_1507);
or U2077 (N_2077,N_1724,N_1695);
nand U2078 (N_2078,N_1780,N_1564);
and U2079 (N_2079,N_1853,N_1630);
nand U2080 (N_2080,N_1526,N_1919);
nor U2081 (N_2081,N_1912,N_1519);
or U2082 (N_2082,N_1529,N_1735);
nand U2083 (N_2083,N_1626,N_1621);
and U2084 (N_2084,N_1585,N_1505);
nand U2085 (N_2085,N_1601,N_1605);
and U2086 (N_2086,N_1648,N_1687);
or U2087 (N_2087,N_1859,N_1751);
and U2088 (N_2088,N_1576,N_1549);
nor U2089 (N_2089,N_1855,N_1878);
nand U2090 (N_2090,N_1828,N_1620);
xnor U2091 (N_2091,N_1757,N_1958);
xnor U2092 (N_2092,N_1523,N_1760);
and U2093 (N_2093,N_1624,N_1673);
and U2094 (N_2094,N_1894,N_1573);
and U2095 (N_2095,N_1534,N_1714);
xor U2096 (N_2096,N_1699,N_1986);
and U2097 (N_2097,N_1644,N_1858);
nand U2098 (N_2098,N_1603,N_1682);
or U2099 (N_2099,N_1829,N_1609);
or U2100 (N_2100,N_1542,N_1879);
nand U2101 (N_2101,N_1937,N_1521);
or U2102 (N_2102,N_1607,N_1796);
or U2103 (N_2103,N_1640,N_1964);
xor U2104 (N_2104,N_1934,N_1999);
or U2105 (N_2105,N_1615,N_1545);
nand U2106 (N_2106,N_1887,N_1525);
or U2107 (N_2107,N_1704,N_1554);
xnor U2108 (N_2108,N_1556,N_1579);
or U2109 (N_2109,N_1581,N_1702);
xor U2110 (N_2110,N_1775,N_1965);
nor U2111 (N_2111,N_1875,N_1975);
nand U2112 (N_2112,N_1643,N_1916);
xnor U2113 (N_2113,N_1719,N_1959);
nand U2114 (N_2114,N_1873,N_1590);
or U2115 (N_2115,N_1629,N_1732);
and U2116 (N_2116,N_1688,N_1717);
nor U2117 (N_2117,N_1785,N_1871);
or U2118 (N_2118,N_1953,N_1929);
nand U2119 (N_2119,N_1618,N_1944);
or U2120 (N_2120,N_1842,N_1928);
nor U2121 (N_2121,N_1671,N_1954);
nand U2122 (N_2122,N_1868,N_1584);
nand U2123 (N_2123,N_1968,N_1535);
nor U2124 (N_2124,N_1995,N_1734);
nor U2125 (N_2125,N_1942,N_1851);
xor U2126 (N_2126,N_1753,N_1703);
or U2127 (N_2127,N_1991,N_1501);
nor U2128 (N_2128,N_1761,N_1767);
or U2129 (N_2129,N_1532,N_1721);
xor U2130 (N_2130,N_1546,N_1992);
xor U2131 (N_2131,N_1974,N_1950);
nand U2132 (N_2132,N_1905,N_1895);
or U2133 (N_2133,N_1848,N_1765);
and U2134 (N_2134,N_1890,N_1743);
and U2135 (N_2135,N_1727,N_1552);
nor U2136 (N_2136,N_1996,N_1908);
or U2137 (N_2137,N_1962,N_1613);
xnor U2138 (N_2138,N_1931,N_1777);
or U2139 (N_2139,N_1659,N_1946);
nand U2140 (N_2140,N_1971,N_1811);
and U2141 (N_2141,N_1802,N_1823);
and U2142 (N_2142,N_1710,N_1847);
xor U2143 (N_2143,N_1957,N_1728);
and U2144 (N_2144,N_1746,N_1625);
or U2145 (N_2145,N_1917,N_1677);
nand U2146 (N_2146,N_1635,N_1516);
or U2147 (N_2147,N_1557,N_1838);
nor U2148 (N_2148,N_1864,N_1676);
xnor U2149 (N_2149,N_1764,N_1694);
or U2150 (N_2150,N_1577,N_1604);
or U2151 (N_2151,N_1565,N_1531);
or U2152 (N_2152,N_1935,N_1826);
or U2153 (N_2153,N_1539,N_1909);
xnor U2154 (N_2154,N_1696,N_1984);
xnor U2155 (N_2155,N_1589,N_1632);
nand U2156 (N_2156,N_1874,N_1716);
or U2157 (N_2157,N_1708,N_1693);
or U2158 (N_2158,N_1787,N_1771);
nor U2159 (N_2159,N_1738,N_1980);
nor U2160 (N_2160,N_1897,N_1821);
or U2161 (N_2161,N_1608,N_1773);
xor U2162 (N_2162,N_1570,N_1706);
and U2163 (N_2163,N_1595,N_1776);
nand U2164 (N_2164,N_1527,N_1675);
nand U2165 (N_2165,N_1982,N_1849);
xor U2166 (N_2166,N_1970,N_1681);
and U2167 (N_2167,N_1813,N_1736);
nand U2168 (N_2168,N_1985,N_1833);
or U2169 (N_2169,N_1622,N_1845);
or U2170 (N_2170,N_1711,N_1825);
and U2171 (N_2171,N_1508,N_1892);
and U2172 (N_2172,N_1540,N_1518);
and U2173 (N_2173,N_1947,N_1762);
or U2174 (N_2174,N_1544,N_1705);
nor U2175 (N_2175,N_1850,N_1956);
or U2176 (N_2176,N_1698,N_1707);
or U2177 (N_2177,N_1815,N_1551);
nand U2178 (N_2178,N_1784,N_1740);
nand U2179 (N_2179,N_1569,N_1730);
or U2180 (N_2180,N_1649,N_1769);
nand U2181 (N_2181,N_1729,N_1709);
nor U2182 (N_2182,N_1830,N_1922);
nor U2183 (N_2183,N_1571,N_1563);
nor U2184 (N_2184,N_1839,N_1515);
nand U2185 (N_2185,N_1650,N_1578);
and U2186 (N_2186,N_1891,N_1888);
nand U2187 (N_2187,N_1538,N_1689);
nor U2188 (N_2188,N_1616,N_1781);
nor U2189 (N_2189,N_1925,N_1739);
and U2190 (N_2190,N_1820,N_1513);
and U2191 (N_2191,N_1528,N_1623);
and U2192 (N_2192,N_1906,N_1910);
nand U2193 (N_2193,N_1914,N_1932);
xnor U2194 (N_2194,N_1759,N_1666);
xor U2195 (N_2195,N_1869,N_1587);
nand U2196 (N_2196,N_1700,N_1841);
or U2197 (N_2197,N_1881,N_1963);
nor U2198 (N_2198,N_1793,N_1856);
and U2199 (N_2199,N_1656,N_1834);
nor U2200 (N_2200,N_1619,N_1798);
nand U2201 (N_2201,N_1749,N_1951);
nand U2202 (N_2202,N_1537,N_1998);
or U2203 (N_2203,N_1817,N_1918);
or U2204 (N_2204,N_1818,N_1763);
and U2205 (N_2205,N_1898,N_1961);
nor U2206 (N_2206,N_1503,N_1586);
nand U2207 (N_2207,N_1840,N_1854);
nor U2208 (N_2208,N_1536,N_1665);
and U2209 (N_2209,N_1804,N_1655);
nand U2210 (N_2210,N_1664,N_1668);
and U2211 (N_2211,N_1766,N_1987);
xnor U2212 (N_2212,N_1997,N_1510);
nand U2213 (N_2213,N_1597,N_1901);
nor U2214 (N_2214,N_1924,N_1634);
nor U2215 (N_2215,N_1748,N_1949);
or U2216 (N_2216,N_1786,N_1788);
and U2217 (N_2217,N_1742,N_1969);
and U2218 (N_2218,N_1756,N_1806);
nor U2219 (N_2219,N_1755,N_1654);
and U2220 (N_2220,N_1835,N_1846);
nor U2221 (N_2221,N_1836,N_1582);
nor U2222 (N_2222,N_1726,N_1860);
and U2223 (N_2223,N_1567,N_1637);
nor U2224 (N_2224,N_1778,N_1752);
nor U2225 (N_2225,N_1642,N_1870);
and U2226 (N_2226,N_1568,N_1880);
and U2227 (N_2227,N_1575,N_1819);
xnor U2228 (N_2228,N_1770,N_1945);
or U2229 (N_2229,N_1754,N_1691);
nand U2230 (N_2230,N_1685,N_1662);
and U2231 (N_2231,N_1979,N_1977);
and U2232 (N_2232,N_1783,N_1904);
and U2233 (N_2233,N_1670,N_1940);
nor U2234 (N_2234,N_1899,N_1967);
and U2235 (N_2235,N_1983,N_1560);
xnor U2236 (N_2236,N_1737,N_1599);
nand U2237 (N_2237,N_1832,N_1801);
xnor U2238 (N_2238,N_1907,N_1824);
nor U2239 (N_2239,N_1758,N_1816);
nand U2240 (N_2240,N_1861,N_1943);
or U2241 (N_2241,N_1647,N_1522);
or U2242 (N_2242,N_1747,N_1720);
nor U2243 (N_2243,N_1857,N_1831);
or U2244 (N_2244,N_1679,N_1641);
nand U2245 (N_2245,N_1952,N_1524);
and U2246 (N_2246,N_1973,N_1731);
nor U2247 (N_2247,N_1672,N_1509);
xor U2248 (N_2248,N_1926,N_1583);
and U2249 (N_2249,N_1805,N_1978);
and U2250 (N_2250,N_1500,N_1834);
and U2251 (N_2251,N_1506,N_1590);
and U2252 (N_2252,N_1787,N_1708);
nor U2253 (N_2253,N_1858,N_1696);
nand U2254 (N_2254,N_1522,N_1560);
or U2255 (N_2255,N_1962,N_1788);
nand U2256 (N_2256,N_1807,N_1763);
nand U2257 (N_2257,N_1784,N_1820);
nor U2258 (N_2258,N_1972,N_1963);
or U2259 (N_2259,N_1883,N_1698);
nor U2260 (N_2260,N_1513,N_1691);
or U2261 (N_2261,N_1972,N_1997);
and U2262 (N_2262,N_1981,N_1930);
and U2263 (N_2263,N_1693,N_1590);
and U2264 (N_2264,N_1952,N_1651);
and U2265 (N_2265,N_1899,N_1854);
nor U2266 (N_2266,N_1766,N_1951);
or U2267 (N_2267,N_1856,N_1561);
nand U2268 (N_2268,N_1679,N_1593);
or U2269 (N_2269,N_1614,N_1548);
nand U2270 (N_2270,N_1908,N_1816);
nor U2271 (N_2271,N_1998,N_1894);
and U2272 (N_2272,N_1764,N_1573);
or U2273 (N_2273,N_1852,N_1560);
nor U2274 (N_2274,N_1922,N_1611);
or U2275 (N_2275,N_1735,N_1975);
or U2276 (N_2276,N_1789,N_1741);
and U2277 (N_2277,N_1545,N_1786);
xor U2278 (N_2278,N_1615,N_1715);
nor U2279 (N_2279,N_1553,N_1624);
or U2280 (N_2280,N_1853,N_1860);
or U2281 (N_2281,N_1749,N_1769);
and U2282 (N_2282,N_1639,N_1621);
and U2283 (N_2283,N_1546,N_1644);
xor U2284 (N_2284,N_1975,N_1609);
or U2285 (N_2285,N_1502,N_1747);
nand U2286 (N_2286,N_1951,N_1690);
nand U2287 (N_2287,N_1534,N_1941);
nor U2288 (N_2288,N_1848,N_1857);
xnor U2289 (N_2289,N_1692,N_1975);
nor U2290 (N_2290,N_1945,N_1691);
nor U2291 (N_2291,N_1661,N_1915);
or U2292 (N_2292,N_1733,N_1868);
or U2293 (N_2293,N_1528,N_1647);
or U2294 (N_2294,N_1991,N_1638);
nand U2295 (N_2295,N_1759,N_1949);
or U2296 (N_2296,N_1697,N_1599);
nor U2297 (N_2297,N_1537,N_1933);
nor U2298 (N_2298,N_1929,N_1613);
and U2299 (N_2299,N_1613,N_1596);
and U2300 (N_2300,N_1669,N_1724);
nand U2301 (N_2301,N_1701,N_1840);
and U2302 (N_2302,N_1961,N_1893);
nand U2303 (N_2303,N_1827,N_1931);
nor U2304 (N_2304,N_1835,N_1681);
and U2305 (N_2305,N_1880,N_1985);
nor U2306 (N_2306,N_1530,N_1565);
and U2307 (N_2307,N_1561,N_1830);
and U2308 (N_2308,N_1909,N_1619);
nand U2309 (N_2309,N_1945,N_1804);
and U2310 (N_2310,N_1782,N_1763);
nand U2311 (N_2311,N_1967,N_1557);
nand U2312 (N_2312,N_1875,N_1619);
and U2313 (N_2313,N_1589,N_1509);
or U2314 (N_2314,N_1896,N_1566);
or U2315 (N_2315,N_1876,N_1850);
nor U2316 (N_2316,N_1876,N_1584);
xor U2317 (N_2317,N_1528,N_1774);
or U2318 (N_2318,N_1671,N_1700);
nand U2319 (N_2319,N_1761,N_1981);
and U2320 (N_2320,N_1574,N_1635);
and U2321 (N_2321,N_1551,N_1813);
nand U2322 (N_2322,N_1753,N_1767);
nand U2323 (N_2323,N_1611,N_1840);
nor U2324 (N_2324,N_1502,N_1543);
or U2325 (N_2325,N_1829,N_1998);
nor U2326 (N_2326,N_1566,N_1990);
nor U2327 (N_2327,N_1626,N_1957);
nor U2328 (N_2328,N_1596,N_1600);
nand U2329 (N_2329,N_1512,N_1709);
nand U2330 (N_2330,N_1591,N_1838);
nor U2331 (N_2331,N_1902,N_1769);
and U2332 (N_2332,N_1733,N_1966);
nor U2333 (N_2333,N_1573,N_1533);
nand U2334 (N_2334,N_1752,N_1574);
nand U2335 (N_2335,N_1803,N_1597);
nor U2336 (N_2336,N_1783,N_1980);
or U2337 (N_2337,N_1529,N_1623);
nand U2338 (N_2338,N_1530,N_1636);
or U2339 (N_2339,N_1509,N_1536);
and U2340 (N_2340,N_1797,N_1814);
nor U2341 (N_2341,N_1821,N_1730);
nor U2342 (N_2342,N_1581,N_1886);
and U2343 (N_2343,N_1762,N_1873);
nand U2344 (N_2344,N_1675,N_1740);
nand U2345 (N_2345,N_1654,N_1565);
or U2346 (N_2346,N_1815,N_1895);
nor U2347 (N_2347,N_1766,N_1676);
or U2348 (N_2348,N_1921,N_1723);
nand U2349 (N_2349,N_1633,N_1956);
and U2350 (N_2350,N_1617,N_1956);
nor U2351 (N_2351,N_1705,N_1931);
and U2352 (N_2352,N_1923,N_1592);
nor U2353 (N_2353,N_1949,N_1879);
or U2354 (N_2354,N_1767,N_1947);
xnor U2355 (N_2355,N_1985,N_1883);
and U2356 (N_2356,N_1649,N_1555);
or U2357 (N_2357,N_1994,N_1770);
or U2358 (N_2358,N_1568,N_1702);
and U2359 (N_2359,N_1706,N_1638);
and U2360 (N_2360,N_1950,N_1646);
nand U2361 (N_2361,N_1996,N_1664);
nand U2362 (N_2362,N_1886,N_1689);
nand U2363 (N_2363,N_1902,N_1568);
nand U2364 (N_2364,N_1668,N_1803);
and U2365 (N_2365,N_1911,N_1843);
nor U2366 (N_2366,N_1757,N_1777);
nand U2367 (N_2367,N_1605,N_1654);
and U2368 (N_2368,N_1641,N_1702);
or U2369 (N_2369,N_1950,N_1798);
or U2370 (N_2370,N_1607,N_1765);
xnor U2371 (N_2371,N_1919,N_1938);
nor U2372 (N_2372,N_1657,N_1649);
or U2373 (N_2373,N_1813,N_1951);
nand U2374 (N_2374,N_1783,N_1641);
nor U2375 (N_2375,N_1627,N_1810);
nand U2376 (N_2376,N_1893,N_1599);
xor U2377 (N_2377,N_1657,N_1653);
and U2378 (N_2378,N_1872,N_1684);
nor U2379 (N_2379,N_1507,N_1842);
or U2380 (N_2380,N_1514,N_1542);
or U2381 (N_2381,N_1717,N_1965);
and U2382 (N_2382,N_1733,N_1523);
or U2383 (N_2383,N_1964,N_1683);
nor U2384 (N_2384,N_1901,N_1750);
nand U2385 (N_2385,N_1897,N_1504);
or U2386 (N_2386,N_1956,N_1780);
xnor U2387 (N_2387,N_1970,N_1539);
and U2388 (N_2388,N_1677,N_1685);
and U2389 (N_2389,N_1564,N_1539);
or U2390 (N_2390,N_1543,N_1775);
and U2391 (N_2391,N_1555,N_1583);
xor U2392 (N_2392,N_1516,N_1716);
nor U2393 (N_2393,N_1897,N_1916);
xnor U2394 (N_2394,N_1582,N_1871);
nor U2395 (N_2395,N_1785,N_1818);
nand U2396 (N_2396,N_1690,N_1571);
nor U2397 (N_2397,N_1720,N_1598);
nor U2398 (N_2398,N_1659,N_1671);
or U2399 (N_2399,N_1963,N_1592);
nor U2400 (N_2400,N_1890,N_1574);
or U2401 (N_2401,N_1795,N_1634);
nand U2402 (N_2402,N_1594,N_1910);
or U2403 (N_2403,N_1838,N_1721);
nand U2404 (N_2404,N_1701,N_1632);
nor U2405 (N_2405,N_1892,N_1909);
xor U2406 (N_2406,N_1856,N_1953);
xor U2407 (N_2407,N_1817,N_1574);
and U2408 (N_2408,N_1710,N_1884);
nor U2409 (N_2409,N_1588,N_1658);
nor U2410 (N_2410,N_1715,N_1703);
or U2411 (N_2411,N_1560,N_1561);
or U2412 (N_2412,N_1524,N_1753);
nand U2413 (N_2413,N_1654,N_1713);
nor U2414 (N_2414,N_1654,N_1511);
nand U2415 (N_2415,N_1938,N_1661);
or U2416 (N_2416,N_1583,N_1903);
and U2417 (N_2417,N_1524,N_1767);
nor U2418 (N_2418,N_1978,N_1604);
nand U2419 (N_2419,N_1577,N_1629);
and U2420 (N_2420,N_1708,N_1839);
and U2421 (N_2421,N_1763,N_1862);
nand U2422 (N_2422,N_1621,N_1503);
or U2423 (N_2423,N_1526,N_1604);
xor U2424 (N_2424,N_1869,N_1582);
or U2425 (N_2425,N_1569,N_1685);
nor U2426 (N_2426,N_1950,N_1959);
or U2427 (N_2427,N_1732,N_1567);
or U2428 (N_2428,N_1641,N_1514);
and U2429 (N_2429,N_1549,N_1726);
and U2430 (N_2430,N_1747,N_1530);
and U2431 (N_2431,N_1851,N_1826);
nand U2432 (N_2432,N_1695,N_1881);
or U2433 (N_2433,N_1821,N_1836);
xor U2434 (N_2434,N_1909,N_1525);
nor U2435 (N_2435,N_1932,N_1805);
nor U2436 (N_2436,N_1695,N_1537);
nand U2437 (N_2437,N_1982,N_1910);
nand U2438 (N_2438,N_1717,N_1919);
nand U2439 (N_2439,N_1794,N_1864);
nor U2440 (N_2440,N_1934,N_1731);
nand U2441 (N_2441,N_1920,N_1848);
xor U2442 (N_2442,N_1650,N_1786);
nand U2443 (N_2443,N_1580,N_1584);
nor U2444 (N_2444,N_1963,N_1608);
nor U2445 (N_2445,N_1654,N_1899);
nand U2446 (N_2446,N_1974,N_1680);
nor U2447 (N_2447,N_1599,N_1690);
nand U2448 (N_2448,N_1513,N_1585);
nand U2449 (N_2449,N_1914,N_1900);
nand U2450 (N_2450,N_1924,N_1745);
and U2451 (N_2451,N_1932,N_1887);
nand U2452 (N_2452,N_1777,N_1953);
and U2453 (N_2453,N_1802,N_1777);
nor U2454 (N_2454,N_1850,N_1628);
nand U2455 (N_2455,N_1619,N_1979);
nand U2456 (N_2456,N_1605,N_1730);
nor U2457 (N_2457,N_1724,N_1665);
nor U2458 (N_2458,N_1646,N_1817);
and U2459 (N_2459,N_1819,N_1731);
nor U2460 (N_2460,N_1904,N_1683);
nor U2461 (N_2461,N_1964,N_1734);
xor U2462 (N_2462,N_1929,N_1826);
or U2463 (N_2463,N_1914,N_1670);
and U2464 (N_2464,N_1862,N_1683);
or U2465 (N_2465,N_1878,N_1857);
nand U2466 (N_2466,N_1923,N_1860);
xnor U2467 (N_2467,N_1505,N_1682);
and U2468 (N_2468,N_1713,N_1954);
or U2469 (N_2469,N_1925,N_1589);
nand U2470 (N_2470,N_1939,N_1933);
or U2471 (N_2471,N_1768,N_1666);
xor U2472 (N_2472,N_1970,N_1976);
or U2473 (N_2473,N_1686,N_1771);
nand U2474 (N_2474,N_1920,N_1715);
xnor U2475 (N_2475,N_1912,N_1909);
and U2476 (N_2476,N_1988,N_1514);
and U2477 (N_2477,N_1831,N_1878);
nand U2478 (N_2478,N_1768,N_1788);
nand U2479 (N_2479,N_1538,N_1587);
and U2480 (N_2480,N_1637,N_1910);
xor U2481 (N_2481,N_1537,N_1560);
nand U2482 (N_2482,N_1532,N_1876);
and U2483 (N_2483,N_1851,N_1721);
or U2484 (N_2484,N_1960,N_1882);
nor U2485 (N_2485,N_1959,N_1698);
nand U2486 (N_2486,N_1898,N_1817);
nand U2487 (N_2487,N_1726,N_1666);
nand U2488 (N_2488,N_1511,N_1691);
or U2489 (N_2489,N_1641,N_1912);
or U2490 (N_2490,N_1818,N_1522);
xnor U2491 (N_2491,N_1999,N_1766);
nor U2492 (N_2492,N_1578,N_1890);
and U2493 (N_2493,N_1840,N_1715);
or U2494 (N_2494,N_1769,N_1597);
nand U2495 (N_2495,N_1831,N_1798);
nand U2496 (N_2496,N_1716,N_1619);
nor U2497 (N_2497,N_1776,N_1580);
nor U2498 (N_2498,N_1806,N_1939);
or U2499 (N_2499,N_1781,N_1797);
nand U2500 (N_2500,N_2117,N_2394);
or U2501 (N_2501,N_2030,N_2225);
nand U2502 (N_2502,N_2297,N_2427);
and U2503 (N_2503,N_2392,N_2376);
nand U2504 (N_2504,N_2323,N_2306);
or U2505 (N_2505,N_2152,N_2230);
xnor U2506 (N_2506,N_2118,N_2383);
or U2507 (N_2507,N_2484,N_2217);
or U2508 (N_2508,N_2182,N_2411);
nand U2509 (N_2509,N_2005,N_2114);
or U2510 (N_2510,N_2069,N_2280);
and U2511 (N_2511,N_2378,N_2149);
nand U2512 (N_2512,N_2399,N_2325);
nand U2513 (N_2513,N_2400,N_2129);
and U2514 (N_2514,N_2353,N_2082);
nand U2515 (N_2515,N_2140,N_2252);
nand U2516 (N_2516,N_2019,N_2169);
nand U2517 (N_2517,N_2421,N_2491);
nor U2518 (N_2518,N_2216,N_2115);
nand U2519 (N_2519,N_2458,N_2103);
nand U2520 (N_2520,N_2262,N_2255);
nor U2521 (N_2521,N_2402,N_2076);
nor U2522 (N_2522,N_2309,N_2305);
nand U2523 (N_2523,N_2112,N_2497);
or U2524 (N_2524,N_2151,N_2153);
or U2525 (N_2525,N_2355,N_2104);
or U2526 (N_2526,N_2126,N_2063);
nand U2527 (N_2527,N_2450,N_2443);
nand U2528 (N_2528,N_2227,N_2423);
and U2529 (N_2529,N_2131,N_2270);
nor U2530 (N_2530,N_2177,N_2037);
nor U2531 (N_2531,N_2387,N_2106);
nand U2532 (N_2532,N_2286,N_2381);
nand U2533 (N_2533,N_2245,N_2235);
nand U2534 (N_2534,N_2460,N_2490);
nand U2535 (N_2535,N_2320,N_2284);
or U2536 (N_2536,N_2304,N_2397);
nand U2537 (N_2537,N_2467,N_2193);
nand U2538 (N_2538,N_2471,N_2242);
nor U2539 (N_2539,N_2477,N_2271);
nor U2540 (N_2540,N_2081,N_2483);
and U2541 (N_2541,N_2016,N_2053);
and U2542 (N_2542,N_2420,N_2260);
nand U2543 (N_2543,N_2318,N_2253);
nand U2544 (N_2544,N_2334,N_2111);
or U2545 (N_2545,N_2316,N_2208);
or U2546 (N_2546,N_2178,N_2027);
nand U2547 (N_2547,N_2404,N_2487);
or U2548 (N_2548,N_2370,N_2422);
or U2549 (N_2549,N_2246,N_2154);
or U2550 (N_2550,N_2220,N_2125);
nor U2551 (N_2551,N_2345,N_2453);
xor U2552 (N_2552,N_2377,N_2013);
nor U2553 (N_2553,N_2061,N_2384);
nor U2554 (N_2554,N_2303,N_2007);
and U2555 (N_2555,N_2444,N_2045);
nand U2556 (N_2556,N_2464,N_2113);
and U2557 (N_2557,N_2031,N_2446);
xnor U2558 (N_2558,N_2163,N_2101);
nand U2559 (N_2559,N_2040,N_2386);
and U2560 (N_2560,N_2447,N_2424);
and U2561 (N_2561,N_2202,N_2234);
or U2562 (N_2562,N_2176,N_2186);
nand U2563 (N_2563,N_2184,N_2134);
nor U2564 (N_2564,N_2480,N_2469);
nor U2565 (N_2565,N_2011,N_2344);
or U2566 (N_2566,N_2493,N_2046);
nand U2567 (N_2567,N_2089,N_2431);
xnor U2568 (N_2568,N_2072,N_2332);
and U2569 (N_2569,N_2142,N_2433);
nor U2570 (N_2570,N_2358,N_2416);
nand U2571 (N_2571,N_2375,N_2247);
nor U2572 (N_2572,N_2071,N_2489);
and U2573 (N_2573,N_2298,N_2165);
xor U2574 (N_2574,N_2024,N_2192);
xnor U2575 (N_2575,N_2273,N_2293);
or U2576 (N_2576,N_2048,N_2197);
or U2577 (N_2577,N_2343,N_2313);
and U2578 (N_2578,N_2002,N_2494);
and U2579 (N_2579,N_2406,N_2495);
and U2580 (N_2580,N_2212,N_2287);
and U2581 (N_2581,N_2060,N_2364);
nand U2582 (N_2582,N_2035,N_2440);
and U2583 (N_2583,N_2354,N_2020);
nand U2584 (N_2584,N_2466,N_2417);
nor U2585 (N_2585,N_2437,N_2401);
and U2586 (N_2586,N_2156,N_2105);
nand U2587 (N_2587,N_2229,N_2055);
or U2588 (N_2588,N_2233,N_2175);
and U2589 (N_2589,N_2391,N_2094);
nor U2590 (N_2590,N_2223,N_2144);
xnor U2591 (N_2591,N_2499,N_2008);
and U2592 (N_2592,N_2419,N_2302);
nand U2593 (N_2593,N_2413,N_2425);
nand U2594 (N_2594,N_2181,N_2241);
nor U2595 (N_2595,N_2108,N_2215);
nor U2596 (N_2596,N_2438,N_2461);
and U2597 (N_2597,N_2341,N_2338);
nor U2598 (N_2598,N_2240,N_2078);
or U2599 (N_2599,N_2064,N_2161);
or U2600 (N_2600,N_2171,N_2195);
and U2601 (N_2601,N_2371,N_2315);
and U2602 (N_2602,N_2412,N_2022);
nand U2603 (N_2603,N_2395,N_2127);
or U2604 (N_2604,N_2367,N_2374);
nand U2605 (N_2605,N_2349,N_2137);
or U2606 (N_2606,N_2026,N_2025);
and U2607 (N_2607,N_2166,N_2258);
nor U2608 (N_2608,N_2362,N_2018);
nor U2609 (N_2609,N_2257,N_2319);
nor U2610 (N_2610,N_2244,N_2167);
or U2611 (N_2611,N_2079,N_2277);
and U2612 (N_2612,N_2296,N_2058);
and U2613 (N_2613,N_2158,N_2199);
or U2614 (N_2614,N_2122,N_2451);
and U2615 (N_2615,N_2096,N_2232);
nand U2616 (N_2616,N_2299,N_2050);
nor U2617 (N_2617,N_2333,N_2256);
and U2618 (N_2618,N_2003,N_2476);
xor U2619 (N_2619,N_2428,N_2357);
and U2620 (N_2620,N_2097,N_2219);
or U2621 (N_2621,N_2363,N_2389);
or U2622 (N_2622,N_2179,N_2472);
and U2623 (N_2623,N_2084,N_2074);
or U2624 (N_2624,N_2164,N_2368);
or U2625 (N_2625,N_2066,N_2330);
nand U2626 (N_2626,N_2100,N_2205);
or U2627 (N_2627,N_2481,N_2265);
nand U2628 (N_2628,N_2017,N_2004);
and U2629 (N_2629,N_2077,N_2174);
or U2630 (N_2630,N_2301,N_2143);
and U2631 (N_2631,N_2308,N_2128);
nor U2632 (N_2632,N_2311,N_2373);
nand U2633 (N_2633,N_2052,N_2398);
or U2634 (N_2634,N_2238,N_2000);
nor U2635 (N_2635,N_2196,N_2148);
nand U2636 (N_2636,N_2083,N_2214);
nand U2637 (N_2637,N_2136,N_2200);
nand U2638 (N_2638,N_2462,N_2041);
or U2639 (N_2639,N_2183,N_2056);
nand U2640 (N_2640,N_2327,N_2087);
nand U2641 (N_2641,N_2021,N_2292);
xnor U2642 (N_2642,N_2231,N_2410);
nand U2643 (N_2643,N_2426,N_2051);
and U2644 (N_2644,N_2390,N_2075);
or U2645 (N_2645,N_2326,N_2057);
or U2646 (N_2646,N_2157,N_2088);
nor U2647 (N_2647,N_2285,N_2123);
nand U2648 (N_2648,N_2482,N_2014);
nand U2649 (N_2649,N_2283,N_2028);
nor U2650 (N_2650,N_2248,N_2243);
and U2651 (N_2651,N_2457,N_2150);
nor U2652 (N_2652,N_2147,N_2145);
or U2653 (N_2653,N_2415,N_2409);
or U2654 (N_2654,N_2172,N_2328);
nor U2655 (N_2655,N_2249,N_2190);
and U2656 (N_2656,N_2359,N_2209);
nand U2657 (N_2657,N_2307,N_2294);
nand U2658 (N_2658,N_2369,N_2288);
nor U2659 (N_2659,N_2485,N_2356);
nor U2660 (N_2660,N_2086,N_2213);
nand U2661 (N_2661,N_2264,N_2237);
and U2662 (N_2662,N_2194,N_2160);
and U2663 (N_2663,N_2073,N_2159);
nand U2664 (N_2664,N_2099,N_2116);
xor U2665 (N_2665,N_2454,N_2130);
or U2666 (N_2666,N_2430,N_2091);
or U2667 (N_2667,N_2329,N_2155);
nand U2668 (N_2668,N_2185,N_2445);
nand U2669 (N_2669,N_2168,N_2351);
nor U2670 (N_2670,N_2488,N_2382);
nand U2671 (N_2671,N_2281,N_2414);
nand U2672 (N_2672,N_2439,N_2203);
nand U2673 (N_2673,N_2442,N_2342);
nand U2674 (N_2674,N_2322,N_2210);
nand U2675 (N_2675,N_2336,N_2317);
nor U2676 (N_2676,N_2204,N_2380);
or U2677 (N_2677,N_2054,N_2366);
and U2678 (N_2678,N_2361,N_2272);
and U2679 (N_2679,N_2173,N_2033);
nor U2680 (N_2680,N_2448,N_2012);
or U2681 (N_2681,N_2043,N_2059);
nor U2682 (N_2682,N_2279,N_2034);
xor U2683 (N_2683,N_2224,N_2095);
and U2684 (N_2684,N_2236,N_2379);
xor U2685 (N_2685,N_2405,N_2070);
nor U2686 (N_2686,N_2119,N_2092);
xnor U2687 (N_2687,N_2010,N_2435);
and U2688 (N_2688,N_2042,N_2463);
nor U2689 (N_2689,N_2352,N_2492);
and U2690 (N_2690,N_2314,N_2187);
and U2691 (N_2691,N_2044,N_2282);
nand U2692 (N_2692,N_2455,N_2062);
nand U2693 (N_2693,N_2408,N_2310);
and U2694 (N_2694,N_2312,N_2189);
nor U2695 (N_2695,N_2407,N_2432);
nor U2696 (N_2696,N_2009,N_2276);
xnor U2697 (N_2697,N_2188,N_2267);
nand U2698 (N_2698,N_2133,N_2218);
nand U2699 (N_2699,N_2478,N_2023);
nor U2700 (N_2700,N_2347,N_2459);
nand U2701 (N_2701,N_2429,N_2486);
nor U2702 (N_2702,N_2228,N_2346);
and U2703 (N_2703,N_2396,N_2139);
nand U2704 (N_2704,N_2001,N_2350);
or U2705 (N_2705,N_2120,N_2065);
nand U2706 (N_2706,N_2449,N_2269);
nand U2707 (N_2707,N_2274,N_2337);
and U2708 (N_2708,N_2470,N_2226);
or U2709 (N_2709,N_2372,N_2268);
nor U2710 (N_2710,N_2465,N_2393);
nand U2711 (N_2711,N_2250,N_2032);
nand U2712 (N_2712,N_2254,N_2475);
nand U2713 (N_2713,N_2290,N_2222);
or U2714 (N_2714,N_2335,N_2038);
or U2715 (N_2715,N_2295,N_2085);
or U2716 (N_2716,N_2047,N_2121);
nor U2717 (N_2717,N_2289,N_2080);
and U2718 (N_2718,N_2110,N_2434);
nor U2719 (N_2719,N_2479,N_2259);
nor U2720 (N_2720,N_2340,N_2365);
and U2721 (N_2721,N_2275,N_2141);
and U2722 (N_2722,N_2263,N_2339);
or U2723 (N_2723,N_2291,N_2029);
nand U2724 (N_2724,N_2221,N_2132);
nand U2725 (N_2725,N_2191,N_2170);
nor U2726 (N_2726,N_2124,N_2403);
and U2727 (N_2727,N_2039,N_2456);
and U2728 (N_2728,N_2049,N_2090);
xnor U2729 (N_2729,N_2107,N_2441);
nor U2730 (N_2730,N_2474,N_2473);
nor U2731 (N_2731,N_2015,N_2206);
and U2732 (N_2732,N_2321,N_2162);
nand U2733 (N_2733,N_2102,N_2201);
and U2734 (N_2734,N_2067,N_2452);
and U2735 (N_2735,N_2251,N_2278);
nand U2736 (N_2736,N_2006,N_2261);
nand U2737 (N_2737,N_2385,N_2135);
nor U2738 (N_2738,N_2498,N_2239);
nand U2739 (N_2739,N_2098,N_2436);
nor U2740 (N_2740,N_2266,N_2388);
xor U2741 (N_2741,N_2324,N_2138);
or U2742 (N_2742,N_2348,N_2468);
and U2743 (N_2743,N_2109,N_2146);
and U2744 (N_2744,N_2331,N_2068);
xnor U2745 (N_2745,N_2496,N_2211);
and U2746 (N_2746,N_2093,N_2300);
nand U2747 (N_2747,N_2418,N_2180);
and U2748 (N_2748,N_2207,N_2036);
or U2749 (N_2749,N_2198,N_2360);
xnor U2750 (N_2750,N_2027,N_2125);
xnor U2751 (N_2751,N_2015,N_2408);
and U2752 (N_2752,N_2340,N_2082);
or U2753 (N_2753,N_2323,N_2187);
and U2754 (N_2754,N_2125,N_2456);
nor U2755 (N_2755,N_2455,N_2273);
nor U2756 (N_2756,N_2173,N_2397);
nand U2757 (N_2757,N_2031,N_2196);
or U2758 (N_2758,N_2201,N_2034);
and U2759 (N_2759,N_2306,N_2468);
and U2760 (N_2760,N_2328,N_2188);
and U2761 (N_2761,N_2362,N_2241);
and U2762 (N_2762,N_2453,N_2012);
and U2763 (N_2763,N_2099,N_2299);
nand U2764 (N_2764,N_2097,N_2403);
nand U2765 (N_2765,N_2413,N_2103);
or U2766 (N_2766,N_2276,N_2023);
and U2767 (N_2767,N_2373,N_2345);
xor U2768 (N_2768,N_2092,N_2401);
or U2769 (N_2769,N_2192,N_2034);
or U2770 (N_2770,N_2173,N_2425);
nor U2771 (N_2771,N_2199,N_2433);
or U2772 (N_2772,N_2414,N_2314);
nand U2773 (N_2773,N_2118,N_2099);
nor U2774 (N_2774,N_2490,N_2459);
xnor U2775 (N_2775,N_2448,N_2108);
and U2776 (N_2776,N_2154,N_2206);
and U2777 (N_2777,N_2392,N_2228);
or U2778 (N_2778,N_2424,N_2013);
nor U2779 (N_2779,N_2251,N_2107);
and U2780 (N_2780,N_2069,N_2109);
or U2781 (N_2781,N_2117,N_2219);
nand U2782 (N_2782,N_2260,N_2399);
nor U2783 (N_2783,N_2045,N_2422);
nor U2784 (N_2784,N_2201,N_2146);
and U2785 (N_2785,N_2091,N_2388);
nand U2786 (N_2786,N_2290,N_2052);
and U2787 (N_2787,N_2008,N_2265);
nand U2788 (N_2788,N_2409,N_2266);
or U2789 (N_2789,N_2400,N_2334);
or U2790 (N_2790,N_2081,N_2102);
nand U2791 (N_2791,N_2004,N_2198);
or U2792 (N_2792,N_2473,N_2288);
and U2793 (N_2793,N_2131,N_2364);
nor U2794 (N_2794,N_2184,N_2351);
or U2795 (N_2795,N_2254,N_2037);
and U2796 (N_2796,N_2086,N_2047);
nand U2797 (N_2797,N_2056,N_2405);
or U2798 (N_2798,N_2456,N_2296);
xor U2799 (N_2799,N_2353,N_2417);
or U2800 (N_2800,N_2061,N_2497);
nor U2801 (N_2801,N_2259,N_2384);
nor U2802 (N_2802,N_2363,N_2182);
and U2803 (N_2803,N_2267,N_2321);
or U2804 (N_2804,N_2470,N_2436);
xor U2805 (N_2805,N_2355,N_2021);
or U2806 (N_2806,N_2153,N_2180);
and U2807 (N_2807,N_2114,N_2452);
nor U2808 (N_2808,N_2036,N_2354);
nand U2809 (N_2809,N_2071,N_2144);
or U2810 (N_2810,N_2044,N_2434);
nand U2811 (N_2811,N_2107,N_2493);
or U2812 (N_2812,N_2484,N_2282);
nand U2813 (N_2813,N_2472,N_2255);
or U2814 (N_2814,N_2008,N_2064);
nand U2815 (N_2815,N_2077,N_2072);
and U2816 (N_2816,N_2126,N_2043);
or U2817 (N_2817,N_2310,N_2376);
nand U2818 (N_2818,N_2118,N_2114);
nand U2819 (N_2819,N_2106,N_2147);
and U2820 (N_2820,N_2433,N_2212);
or U2821 (N_2821,N_2274,N_2052);
nand U2822 (N_2822,N_2101,N_2389);
nor U2823 (N_2823,N_2364,N_2194);
nand U2824 (N_2824,N_2471,N_2199);
nor U2825 (N_2825,N_2078,N_2129);
and U2826 (N_2826,N_2380,N_2270);
or U2827 (N_2827,N_2196,N_2474);
or U2828 (N_2828,N_2243,N_2356);
nor U2829 (N_2829,N_2431,N_2111);
or U2830 (N_2830,N_2124,N_2106);
xnor U2831 (N_2831,N_2379,N_2148);
nor U2832 (N_2832,N_2046,N_2264);
nor U2833 (N_2833,N_2246,N_2181);
and U2834 (N_2834,N_2051,N_2121);
nor U2835 (N_2835,N_2051,N_2280);
xor U2836 (N_2836,N_2474,N_2364);
nand U2837 (N_2837,N_2118,N_2096);
nor U2838 (N_2838,N_2028,N_2261);
nor U2839 (N_2839,N_2451,N_2114);
or U2840 (N_2840,N_2176,N_2244);
or U2841 (N_2841,N_2045,N_2323);
nand U2842 (N_2842,N_2236,N_2026);
or U2843 (N_2843,N_2354,N_2203);
nand U2844 (N_2844,N_2372,N_2178);
and U2845 (N_2845,N_2204,N_2327);
and U2846 (N_2846,N_2280,N_2452);
nor U2847 (N_2847,N_2317,N_2176);
and U2848 (N_2848,N_2396,N_2287);
nand U2849 (N_2849,N_2147,N_2217);
nand U2850 (N_2850,N_2103,N_2213);
and U2851 (N_2851,N_2281,N_2120);
nor U2852 (N_2852,N_2448,N_2124);
and U2853 (N_2853,N_2007,N_2000);
or U2854 (N_2854,N_2390,N_2232);
nand U2855 (N_2855,N_2192,N_2011);
and U2856 (N_2856,N_2155,N_2159);
or U2857 (N_2857,N_2394,N_2404);
and U2858 (N_2858,N_2485,N_2213);
or U2859 (N_2859,N_2442,N_2005);
or U2860 (N_2860,N_2189,N_2148);
xor U2861 (N_2861,N_2361,N_2452);
nor U2862 (N_2862,N_2236,N_2142);
nand U2863 (N_2863,N_2287,N_2305);
or U2864 (N_2864,N_2298,N_2346);
and U2865 (N_2865,N_2374,N_2094);
and U2866 (N_2866,N_2386,N_2472);
nand U2867 (N_2867,N_2385,N_2213);
xor U2868 (N_2868,N_2071,N_2038);
nor U2869 (N_2869,N_2226,N_2402);
and U2870 (N_2870,N_2495,N_2135);
nand U2871 (N_2871,N_2209,N_2224);
or U2872 (N_2872,N_2195,N_2201);
nand U2873 (N_2873,N_2374,N_2370);
nor U2874 (N_2874,N_2433,N_2341);
and U2875 (N_2875,N_2318,N_2404);
or U2876 (N_2876,N_2281,N_2007);
and U2877 (N_2877,N_2347,N_2478);
and U2878 (N_2878,N_2316,N_2308);
and U2879 (N_2879,N_2022,N_2069);
nand U2880 (N_2880,N_2302,N_2476);
nor U2881 (N_2881,N_2314,N_2295);
xor U2882 (N_2882,N_2492,N_2428);
nor U2883 (N_2883,N_2296,N_2067);
nand U2884 (N_2884,N_2100,N_2165);
nor U2885 (N_2885,N_2396,N_2134);
or U2886 (N_2886,N_2032,N_2389);
or U2887 (N_2887,N_2375,N_2484);
nor U2888 (N_2888,N_2288,N_2296);
nor U2889 (N_2889,N_2353,N_2252);
nand U2890 (N_2890,N_2490,N_2190);
nand U2891 (N_2891,N_2018,N_2151);
nor U2892 (N_2892,N_2310,N_2364);
and U2893 (N_2893,N_2377,N_2186);
xnor U2894 (N_2894,N_2438,N_2443);
nor U2895 (N_2895,N_2186,N_2406);
nand U2896 (N_2896,N_2107,N_2457);
nand U2897 (N_2897,N_2238,N_2002);
nor U2898 (N_2898,N_2408,N_2106);
xnor U2899 (N_2899,N_2187,N_2409);
or U2900 (N_2900,N_2018,N_2078);
or U2901 (N_2901,N_2419,N_2418);
and U2902 (N_2902,N_2173,N_2307);
or U2903 (N_2903,N_2027,N_2226);
nor U2904 (N_2904,N_2015,N_2212);
nand U2905 (N_2905,N_2265,N_2369);
or U2906 (N_2906,N_2251,N_2482);
nand U2907 (N_2907,N_2010,N_2232);
xor U2908 (N_2908,N_2252,N_2049);
xor U2909 (N_2909,N_2431,N_2223);
or U2910 (N_2910,N_2347,N_2201);
xnor U2911 (N_2911,N_2244,N_2072);
nor U2912 (N_2912,N_2484,N_2255);
nand U2913 (N_2913,N_2293,N_2010);
or U2914 (N_2914,N_2250,N_2094);
or U2915 (N_2915,N_2462,N_2416);
and U2916 (N_2916,N_2095,N_2065);
or U2917 (N_2917,N_2413,N_2192);
nor U2918 (N_2918,N_2150,N_2250);
and U2919 (N_2919,N_2174,N_2159);
nor U2920 (N_2920,N_2159,N_2429);
or U2921 (N_2921,N_2297,N_2419);
nor U2922 (N_2922,N_2214,N_2044);
and U2923 (N_2923,N_2411,N_2308);
or U2924 (N_2924,N_2158,N_2313);
or U2925 (N_2925,N_2012,N_2133);
nand U2926 (N_2926,N_2223,N_2435);
and U2927 (N_2927,N_2128,N_2468);
and U2928 (N_2928,N_2302,N_2147);
nand U2929 (N_2929,N_2079,N_2064);
nor U2930 (N_2930,N_2410,N_2383);
or U2931 (N_2931,N_2476,N_2362);
or U2932 (N_2932,N_2370,N_2477);
nand U2933 (N_2933,N_2089,N_2265);
xnor U2934 (N_2934,N_2072,N_2251);
nand U2935 (N_2935,N_2470,N_2014);
nand U2936 (N_2936,N_2359,N_2322);
or U2937 (N_2937,N_2269,N_2295);
nand U2938 (N_2938,N_2450,N_2053);
and U2939 (N_2939,N_2310,N_2480);
and U2940 (N_2940,N_2219,N_2193);
and U2941 (N_2941,N_2343,N_2363);
or U2942 (N_2942,N_2046,N_2087);
xor U2943 (N_2943,N_2119,N_2417);
or U2944 (N_2944,N_2000,N_2432);
nor U2945 (N_2945,N_2351,N_2107);
and U2946 (N_2946,N_2111,N_2020);
xor U2947 (N_2947,N_2229,N_2020);
nand U2948 (N_2948,N_2005,N_2137);
nor U2949 (N_2949,N_2042,N_2388);
and U2950 (N_2950,N_2257,N_2157);
or U2951 (N_2951,N_2047,N_2068);
or U2952 (N_2952,N_2145,N_2393);
nor U2953 (N_2953,N_2148,N_2333);
and U2954 (N_2954,N_2338,N_2089);
nand U2955 (N_2955,N_2031,N_2354);
nor U2956 (N_2956,N_2476,N_2019);
or U2957 (N_2957,N_2165,N_2095);
or U2958 (N_2958,N_2453,N_2225);
and U2959 (N_2959,N_2332,N_2465);
nor U2960 (N_2960,N_2028,N_2405);
or U2961 (N_2961,N_2366,N_2073);
nor U2962 (N_2962,N_2350,N_2426);
xnor U2963 (N_2963,N_2238,N_2266);
or U2964 (N_2964,N_2072,N_2050);
or U2965 (N_2965,N_2282,N_2353);
and U2966 (N_2966,N_2497,N_2367);
nand U2967 (N_2967,N_2451,N_2118);
and U2968 (N_2968,N_2438,N_2349);
nor U2969 (N_2969,N_2273,N_2307);
nor U2970 (N_2970,N_2055,N_2050);
nand U2971 (N_2971,N_2490,N_2266);
nor U2972 (N_2972,N_2005,N_2379);
nand U2973 (N_2973,N_2088,N_2481);
nand U2974 (N_2974,N_2407,N_2261);
nor U2975 (N_2975,N_2300,N_2396);
nor U2976 (N_2976,N_2071,N_2033);
or U2977 (N_2977,N_2067,N_2421);
or U2978 (N_2978,N_2414,N_2266);
and U2979 (N_2979,N_2428,N_2412);
nand U2980 (N_2980,N_2173,N_2010);
and U2981 (N_2981,N_2192,N_2366);
nand U2982 (N_2982,N_2009,N_2055);
nand U2983 (N_2983,N_2457,N_2092);
nand U2984 (N_2984,N_2007,N_2492);
xor U2985 (N_2985,N_2462,N_2118);
or U2986 (N_2986,N_2053,N_2367);
and U2987 (N_2987,N_2341,N_2428);
nor U2988 (N_2988,N_2284,N_2286);
or U2989 (N_2989,N_2080,N_2276);
nand U2990 (N_2990,N_2174,N_2444);
and U2991 (N_2991,N_2064,N_2222);
and U2992 (N_2992,N_2159,N_2355);
nor U2993 (N_2993,N_2443,N_2177);
or U2994 (N_2994,N_2348,N_2061);
nor U2995 (N_2995,N_2146,N_2288);
and U2996 (N_2996,N_2169,N_2275);
and U2997 (N_2997,N_2187,N_2285);
or U2998 (N_2998,N_2373,N_2443);
and U2999 (N_2999,N_2185,N_2418);
and U3000 (N_3000,N_2849,N_2851);
nand U3001 (N_3001,N_2758,N_2918);
and U3002 (N_3002,N_2947,N_2940);
or U3003 (N_3003,N_2829,N_2696);
nor U3004 (N_3004,N_2846,N_2586);
nand U3005 (N_3005,N_2527,N_2782);
and U3006 (N_3006,N_2732,N_2518);
xor U3007 (N_3007,N_2894,N_2889);
nor U3008 (N_3008,N_2835,N_2797);
xor U3009 (N_3009,N_2517,N_2890);
nand U3010 (N_3010,N_2552,N_2824);
nor U3011 (N_3011,N_2999,N_2744);
and U3012 (N_3012,N_2583,N_2653);
nand U3013 (N_3013,N_2925,N_2861);
or U3014 (N_3014,N_2743,N_2862);
xnor U3015 (N_3015,N_2562,N_2981);
and U3016 (N_3016,N_2612,N_2971);
xnor U3017 (N_3017,N_2593,N_2860);
and U3018 (N_3018,N_2854,N_2775);
nand U3019 (N_3019,N_2974,N_2932);
xnor U3020 (N_3020,N_2572,N_2872);
nor U3021 (N_3021,N_2560,N_2605);
nand U3022 (N_3022,N_2624,N_2539);
nand U3023 (N_3023,N_2810,N_2841);
and U3024 (N_3024,N_2815,N_2937);
xor U3025 (N_3025,N_2858,N_2968);
or U3026 (N_3026,N_2659,N_2726);
or U3027 (N_3027,N_2965,N_2707);
nand U3028 (N_3028,N_2542,N_2808);
and U3029 (N_3029,N_2695,N_2551);
nor U3030 (N_3030,N_2781,N_2504);
nor U3031 (N_3031,N_2864,N_2511);
and U3032 (N_3032,N_2859,N_2961);
nor U3033 (N_3033,N_2746,N_2591);
or U3034 (N_3034,N_2990,N_2959);
nand U3035 (N_3035,N_2803,N_2789);
xor U3036 (N_3036,N_2745,N_2665);
or U3037 (N_3037,N_2727,N_2700);
and U3038 (N_3038,N_2784,N_2523);
nand U3039 (N_3039,N_2931,N_2589);
and U3040 (N_3040,N_2888,N_2832);
or U3041 (N_3041,N_2577,N_2655);
nor U3042 (N_3042,N_2935,N_2924);
or U3043 (N_3043,N_2647,N_2760);
nor U3044 (N_3044,N_2598,N_2666);
and U3045 (N_3045,N_2934,N_2801);
and U3046 (N_3046,N_2923,N_2609);
nand U3047 (N_3047,N_2541,N_2530);
nor U3048 (N_3048,N_2713,N_2709);
and U3049 (N_3049,N_2876,N_2607);
and U3050 (N_3050,N_2857,N_2712);
nand U3051 (N_3051,N_2936,N_2692);
or U3052 (N_3052,N_2818,N_2989);
nand U3053 (N_3053,N_2617,N_2926);
nand U3054 (N_3054,N_2730,N_2564);
nor U3055 (N_3055,N_2606,N_2930);
or U3056 (N_3056,N_2597,N_2515);
or U3057 (N_3057,N_2718,N_2741);
and U3058 (N_3058,N_2643,N_2977);
nor U3059 (N_3059,N_2626,N_2793);
and U3060 (N_3060,N_2948,N_2615);
nor U3061 (N_3061,N_2637,N_2817);
nor U3062 (N_3062,N_2919,N_2717);
or U3063 (N_3063,N_2529,N_2688);
and U3064 (N_3064,N_2522,N_2806);
xor U3065 (N_3065,N_2650,N_2594);
and U3066 (N_3066,N_2933,N_2544);
nand U3067 (N_3067,N_2502,N_2619);
xnor U3068 (N_3068,N_2865,N_2507);
nand U3069 (N_3069,N_2673,N_2592);
or U3070 (N_3070,N_2847,N_2869);
or U3071 (N_3071,N_2773,N_2769);
nand U3072 (N_3072,N_2599,N_2505);
and U3073 (N_3073,N_2979,N_2702);
or U3074 (N_3074,N_2677,N_2831);
and U3075 (N_3075,N_2680,N_2553);
or U3076 (N_3076,N_2545,N_2761);
and U3077 (N_3077,N_2557,N_2568);
and U3078 (N_3078,N_2994,N_2570);
and U3079 (N_3079,N_2852,N_2682);
xor U3080 (N_3080,N_2500,N_2833);
nand U3081 (N_3081,N_2715,N_2516);
and U3082 (N_3082,N_2903,N_2799);
nor U3083 (N_3083,N_2873,N_2770);
and U3084 (N_3084,N_2705,N_2762);
or U3085 (N_3085,N_2842,N_2674);
nand U3086 (N_3086,N_2883,N_2764);
or U3087 (N_3087,N_2565,N_2547);
nand U3088 (N_3088,N_2897,N_2588);
or U3089 (N_3089,N_2834,N_2640);
or U3090 (N_3090,N_2519,N_2942);
xor U3091 (N_3091,N_2644,N_2687);
nand U3092 (N_3092,N_2711,N_2955);
xor U3093 (N_3093,N_2976,N_2549);
nand U3094 (N_3094,N_2967,N_2885);
and U3095 (N_3095,N_2988,N_2941);
xnor U3096 (N_3096,N_2657,N_2649);
and U3097 (N_3097,N_2908,N_2870);
and U3098 (N_3098,N_2953,N_2578);
nor U3099 (N_3099,N_2735,N_2914);
nand U3100 (N_3100,N_2874,N_2658);
nand U3101 (N_3101,N_2752,N_2907);
or U3102 (N_3102,N_2652,N_2915);
nor U3103 (N_3103,N_2526,N_2997);
and U3104 (N_3104,N_2962,N_2664);
nor U3105 (N_3105,N_2618,N_2710);
xor U3106 (N_3106,N_2689,N_2729);
or U3107 (N_3107,N_2813,N_2899);
and U3108 (N_3108,N_2563,N_2699);
nand U3109 (N_3109,N_2748,N_2638);
nor U3110 (N_3110,N_2683,N_2843);
nand U3111 (N_3111,N_2807,N_2678);
nand U3112 (N_3112,N_2958,N_2755);
or U3113 (N_3113,N_2927,N_2540);
and U3114 (N_3114,N_2508,N_2736);
xnor U3115 (N_3115,N_2534,N_2698);
nand U3116 (N_3116,N_2892,N_2716);
nand U3117 (N_3117,N_2884,N_2840);
nand U3118 (N_3118,N_2660,N_2998);
and U3119 (N_3119,N_2567,N_2654);
and U3120 (N_3120,N_2603,N_2632);
xnor U3121 (N_3121,N_2800,N_2796);
nand U3122 (N_3122,N_2561,N_2641);
and U3123 (N_3123,N_2697,N_2728);
xnor U3124 (N_3124,N_2780,N_2992);
nor U3125 (N_3125,N_2996,N_2573);
nor U3126 (N_3126,N_2929,N_2628);
nand U3127 (N_3127,N_2521,N_2820);
nor U3128 (N_3128,N_2763,N_2610);
nand U3129 (N_3129,N_2809,N_2646);
nand U3130 (N_3130,N_2821,N_2811);
and U3131 (N_3131,N_2566,N_2853);
nand U3132 (N_3132,N_2768,N_2771);
xor U3133 (N_3133,N_2531,N_2604);
nor U3134 (N_3134,N_2537,N_2788);
xnor U3135 (N_3135,N_2951,N_2737);
nand U3136 (N_3136,N_2751,N_2895);
xor U3137 (N_3137,N_2957,N_2816);
and U3138 (N_3138,N_2661,N_2920);
xnor U3139 (N_3139,N_2804,N_2891);
and U3140 (N_3140,N_2669,N_2532);
or U3141 (N_3141,N_2886,N_2651);
nand U3142 (N_3142,N_2946,N_2798);
xnor U3143 (N_3143,N_2635,N_2837);
nand U3144 (N_3144,N_2765,N_2670);
nand U3145 (N_3145,N_2686,N_2571);
xor U3146 (N_3146,N_2645,N_2533);
xor U3147 (N_3147,N_2587,N_2877);
and U3148 (N_3148,N_2916,N_2772);
or U3149 (N_3149,N_2738,N_2595);
xor U3150 (N_3150,N_2912,N_2528);
nand U3151 (N_3151,N_2778,N_2671);
or U3152 (N_3152,N_2574,N_2792);
nor U3153 (N_3153,N_2921,N_2902);
nand U3154 (N_3154,N_2911,N_2719);
nand U3155 (N_3155,N_2830,N_2882);
and U3156 (N_3156,N_2721,N_2950);
nand U3157 (N_3157,N_2945,N_2724);
and U3158 (N_3158,N_2867,N_2938);
and U3159 (N_3159,N_2706,N_2900);
or U3160 (N_3160,N_2787,N_2759);
nor U3161 (N_3161,N_2734,N_2575);
and U3162 (N_3162,N_2939,N_2856);
nor U3163 (N_3163,N_2960,N_2753);
or U3164 (N_3164,N_2579,N_2723);
or U3165 (N_3165,N_2648,N_2703);
or U3166 (N_3166,N_2693,N_2836);
or U3167 (N_3167,N_2898,N_2613);
or U3168 (N_3168,N_2827,N_2621);
and U3169 (N_3169,N_2868,N_2584);
or U3170 (N_3170,N_2986,N_2987);
and U3171 (N_3171,N_2656,N_2554);
nand U3172 (N_3172,N_2733,N_2905);
or U3173 (N_3173,N_2614,N_2576);
or U3174 (N_3174,N_2754,N_2558);
or U3175 (N_3175,N_2616,N_2995);
nand U3176 (N_3176,N_2582,N_2909);
nor U3177 (N_3177,N_2879,N_2904);
nor U3178 (N_3178,N_2520,N_2863);
nand U3179 (N_3179,N_2783,N_2910);
and U3180 (N_3180,N_2684,N_2952);
or U3181 (N_3181,N_2602,N_2901);
nor U3182 (N_3182,N_2708,N_2963);
or U3183 (N_3183,N_2625,N_2601);
nor U3184 (N_3184,N_2510,N_2585);
nand U3185 (N_3185,N_2631,N_2720);
nor U3186 (N_3186,N_2819,N_2668);
nand U3187 (N_3187,N_2893,N_2675);
and U3188 (N_3188,N_2949,N_2636);
nand U3189 (N_3189,N_2805,N_2972);
or U3190 (N_3190,N_2690,N_2917);
nor U3191 (N_3191,N_2747,N_2774);
nand U3192 (N_3192,N_2633,N_2506);
or U3193 (N_3193,N_2590,N_2524);
or U3194 (N_3194,N_2913,N_2548);
and U3195 (N_3195,N_2828,N_2786);
or U3196 (N_3196,N_2975,N_2725);
or U3197 (N_3197,N_2581,N_2826);
and U3198 (N_3198,N_2731,N_2676);
or U3199 (N_3199,N_2823,N_2922);
or U3200 (N_3200,N_2559,N_2878);
and U3201 (N_3201,N_2896,N_2756);
nor U3202 (N_3202,N_2982,N_2662);
or U3203 (N_3203,N_2776,N_2825);
nor U3204 (N_3204,N_2866,N_2642);
nor U3205 (N_3205,N_2794,N_2546);
nor U3206 (N_3206,N_2964,N_2634);
or U3207 (N_3207,N_2501,N_2795);
and U3208 (N_3208,N_2956,N_2875);
or U3209 (N_3209,N_2749,N_2694);
or U3210 (N_3210,N_2538,N_2844);
nand U3211 (N_3211,N_2750,N_2779);
nand U3212 (N_3212,N_2685,N_2740);
nor U3213 (N_3213,N_2639,N_2627);
or U3214 (N_3214,N_2785,N_2993);
or U3215 (N_3215,N_2535,N_2681);
nand U3216 (N_3216,N_2679,N_2556);
and U3217 (N_3217,N_2767,N_2611);
xnor U3218 (N_3218,N_2944,N_2871);
nor U3219 (N_3219,N_2701,N_2814);
and U3220 (N_3220,N_2943,N_2973);
nor U3221 (N_3221,N_2822,N_2954);
nor U3222 (N_3222,N_2848,N_2691);
nor U3223 (N_3223,N_2629,N_2600);
or U3224 (N_3224,N_2881,N_2791);
nand U3225 (N_3225,N_2622,N_2980);
and U3226 (N_3226,N_2580,N_2623);
nand U3227 (N_3227,N_2536,N_2969);
and U3228 (N_3228,N_2596,N_2984);
nor U3229 (N_3229,N_2555,N_2714);
nand U3230 (N_3230,N_2790,N_2887);
nand U3231 (N_3231,N_2757,N_2667);
nand U3232 (N_3232,N_2742,N_2991);
nor U3233 (N_3233,N_2928,N_2970);
nand U3234 (N_3234,N_2802,N_2630);
or U3235 (N_3235,N_2543,N_2550);
xor U3236 (N_3236,N_2608,N_2509);
nand U3237 (N_3237,N_2839,N_2503);
nand U3238 (N_3238,N_2966,N_2525);
xnor U3239 (N_3239,N_2722,N_2978);
nor U3240 (N_3240,N_2620,N_2985);
nand U3241 (N_3241,N_2777,N_2739);
nor U3242 (N_3242,N_2855,N_2704);
nand U3243 (N_3243,N_2663,N_2812);
or U3244 (N_3244,N_2838,N_2850);
nor U3245 (N_3245,N_2845,N_2514);
or U3246 (N_3246,N_2983,N_2513);
or U3247 (N_3247,N_2569,N_2880);
or U3248 (N_3248,N_2766,N_2672);
nor U3249 (N_3249,N_2512,N_2906);
or U3250 (N_3250,N_2623,N_2720);
and U3251 (N_3251,N_2722,N_2544);
nor U3252 (N_3252,N_2782,N_2822);
or U3253 (N_3253,N_2607,N_2703);
and U3254 (N_3254,N_2627,N_2807);
or U3255 (N_3255,N_2670,N_2907);
or U3256 (N_3256,N_2968,N_2737);
or U3257 (N_3257,N_2917,N_2544);
or U3258 (N_3258,N_2960,N_2633);
or U3259 (N_3259,N_2945,N_2866);
nand U3260 (N_3260,N_2956,N_2656);
nor U3261 (N_3261,N_2885,N_2593);
nor U3262 (N_3262,N_2597,N_2760);
nand U3263 (N_3263,N_2581,N_2930);
nand U3264 (N_3264,N_2757,N_2944);
or U3265 (N_3265,N_2676,N_2944);
or U3266 (N_3266,N_2809,N_2651);
nor U3267 (N_3267,N_2997,N_2853);
or U3268 (N_3268,N_2806,N_2708);
nor U3269 (N_3269,N_2582,N_2798);
and U3270 (N_3270,N_2729,N_2945);
nor U3271 (N_3271,N_2692,N_2758);
xor U3272 (N_3272,N_2500,N_2576);
nor U3273 (N_3273,N_2598,N_2541);
or U3274 (N_3274,N_2506,N_2839);
nor U3275 (N_3275,N_2876,N_2827);
nand U3276 (N_3276,N_2895,N_2586);
and U3277 (N_3277,N_2542,N_2837);
xor U3278 (N_3278,N_2564,N_2961);
nand U3279 (N_3279,N_2923,N_2518);
and U3280 (N_3280,N_2603,N_2948);
nor U3281 (N_3281,N_2995,N_2946);
and U3282 (N_3282,N_2713,N_2975);
nand U3283 (N_3283,N_2793,N_2862);
nor U3284 (N_3284,N_2758,N_2805);
or U3285 (N_3285,N_2835,N_2606);
nand U3286 (N_3286,N_2936,N_2950);
nand U3287 (N_3287,N_2901,N_2763);
nor U3288 (N_3288,N_2959,N_2522);
and U3289 (N_3289,N_2511,N_2825);
xor U3290 (N_3290,N_2737,N_2915);
nand U3291 (N_3291,N_2539,N_2723);
nor U3292 (N_3292,N_2689,N_2529);
and U3293 (N_3293,N_2604,N_2949);
or U3294 (N_3294,N_2613,N_2894);
xor U3295 (N_3295,N_2662,N_2685);
and U3296 (N_3296,N_2926,N_2521);
or U3297 (N_3297,N_2608,N_2585);
nor U3298 (N_3298,N_2604,N_2860);
nand U3299 (N_3299,N_2973,N_2561);
and U3300 (N_3300,N_2501,N_2757);
or U3301 (N_3301,N_2630,N_2936);
or U3302 (N_3302,N_2851,N_2565);
xor U3303 (N_3303,N_2945,N_2737);
nor U3304 (N_3304,N_2631,N_2535);
nor U3305 (N_3305,N_2650,N_2748);
nand U3306 (N_3306,N_2869,N_2751);
nor U3307 (N_3307,N_2766,N_2967);
nand U3308 (N_3308,N_2976,N_2587);
or U3309 (N_3309,N_2605,N_2892);
and U3310 (N_3310,N_2826,N_2871);
and U3311 (N_3311,N_2802,N_2642);
or U3312 (N_3312,N_2966,N_2993);
and U3313 (N_3313,N_2794,N_2908);
or U3314 (N_3314,N_2571,N_2624);
or U3315 (N_3315,N_2755,N_2655);
nor U3316 (N_3316,N_2610,N_2928);
nor U3317 (N_3317,N_2559,N_2916);
or U3318 (N_3318,N_2997,N_2844);
nor U3319 (N_3319,N_2963,N_2927);
nor U3320 (N_3320,N_2850,N_2902);
xor U3321 (N_3321,N_2642,N_2751);
nand U3322 (N_3322,N_2838,N_2817);
xnor U3323 (N_3323,N_2742,N_2573);
or U3324 (N_3324,N_2771,N_2688);
and U3325 (N_3325,N_2735,N_2912);
xor U3326 (N_3326,N_2791,N_2640);
nor U3327 (N_3327,N_2777,N_2582);
xor U3328 (N_3328,N_2583,N_2987);
or U3329 (N_3329,N_2599,N_2652);
nor U3330 (N_3330,N_2618,N_2578);
nor U3331 (N_3331,N_2974,N_2897);
and U3332 (N_3332,N_2720,N_2777);
nor U3333 (N_3333,N_2712,N_2566);
nor U3334 (N_3334,N_2940,N_2776);
and U3335 (N_3335,N_2912,N_2823);
xnor U3336 (N_3336,N_2511,N_2547);
nand U3337 (N_3337,N_2720,N_2672);
and U3338 (N_3338,N_2681,N_2987);
xnor U3339 (N_3339,N_2808,N_2511);
and U3340 (N_3340,N_2832,N_2564);
nand U3341 (N_3341,N_2762,N_2801);
or U3342 (N_3342,N_2932,N_2814);
and U3343 (N_3343,N_2971,N_2562);
and U3344 (N_3344,N_2947,N_2781);
or U3345 (N_3345,N_2740,N_2816);
and U3346 (N_3346,N_2574,N_2738);
nand U3347 (N_3347,N_2677,N_2864);
or U3348 (N_3348,N_2705,N_2504);
nand U3349 (N_3349,N_2585,N_2773);
nor U3350 (N_3350,N_2517,N_2925);
or U3351 (N_3351,N_2928,N_2513);
and U3352 (N_3352,N_2623,N_2537);
and U3353 (N_3353,N_2797,N_2530);
xor U3354 (N_3354,N_2976,N_2915);
xor U3355 (N_3355,N_2694,N_2513);
nor U3356 (N_3356,N_2697,N_2627);
nor U3357 (N_3357,N_2658,N_2782);
or U3358 (N_3358,N_2706,N_2915);
and U3359 (N_3359,N_2941,N_2626);
nor U3360 (N_3360,N_2846,N_2501);
nor U3361 (N_3361,N_2753,N_2982);
and U3362 (N_3362,N_2627,N_2555);
or U3363 (N_3363,N_2875,N_2580);
nor U3364 (N_3364,N_2933,N_2501);
nor U3365 (N_3365,N_2939,N_2592);
xor U3366 (N_3366,N_2572,N_2679);
or U3367 (N_3367,N_2551,N_2617);
and U3368 (N_3368,N_2942,N_2777);
or U3369 (N_3369,N_2848,N_2972);
nand U3370 (N_3370,N_2771,N_2794);
or U3371 (N_3371,N_2525,N_2872);
and U3372 (N_3372,N_2740,N_2731);
nor U3373 (N_3373,N_2673,N_2710);
xnor U3374 (N_3374,N_2931,N_2808);
or U3375 (N_3375,N_2687,N_2688);
nand U3376 (N_3376,N_2881,N_2783);
nand U3377 (N_3377,N_2872,N_2640);
xor U3378 (N_3378,N_2650,N_2530);
nor U3379 (N_3379,N_2879,N_2538);
and U3380 (N_3380,N_2975,N_2706);
nor U3381 (N_3381,N_2894,N_2595);
nand U3382 (N_3382,N_2580,N_2688);
nor U3383 (N_3383,N_2732,N_2730);
and U3384 (N_3384,N_2805,N_2723);
nand U3385 (N_3385,N_2746,N_2912);
nor U3386 (N_3386,N_2999,N_2929);
nor U3387 (N_3387,N_2894,N_2920);
and U3388 (N_3388,N_2969,N_2750);
nor U3389 (N_3389,N_2940,N_2699);
nor U3390 (N_3390,N_2573,N_2966);
nor U3391 (N_3391,N_2855,N_2944);
xnor U3392 (N_3392,N_2824,N_2516);
nor U3393 (N_3393,N_2574,N_2845);
nand U3394 (N_3394,N_2553,N_2536);
nand U3395 (N_3395,N_2749,N_2996);
nor U3396 (N_3396,N_2879,N_2650);
nand U3397 (N_3397,N_2959,N_2993);
or U3398 (N_3398,N_2864,N_2760);
or U3399 (N_3399,N_2903,N_2885);
nor U3400 (N_3400,N_2647,N_2833);
xnor U3401 (N_3401,N_2930,N_2757);
nor U3402 (N_3402,N_2973,N_2667);
and U3403 (N_3403,N_2643,N_2889);
nand U3404 (N_3404,N_2853,N_2749);
xnor U3405 (N_3405,N_2874,N_2618);
and U3406 (N_3406,N_2872,N_2900);
and U3407 (N_3407,N_2621,N_2826);
or U3408 (N_3408,N_2859,N_2881);
nor U3409 (N_3409,N_2988,N_2779);
or U3410 (N_3410,N_2667,N_2825);
and U3411 (N_3411,N_2728,N_2950);
nand U3412 (N_3412,N_2703,N_2911);
nor U3413 (N_3413,N_2685,N_2833);
and U3414 (N_3414,N_2710,N_2989);
nand U3415 (N_3415,N_2861,N_2686);
or U3416 (N_3416,N_2657,N_2788);
nor U3417 (N_3417,N_2827,N_2540);
and U3418 (N_3418,N_2896,N_2780);
and U3419 (N_3419,N_2682,N_2726);
nor U3420 (N_3420,N_2827,N_2728);
nand U3421 (N_3421,N_2607,N_2622);
nor U3422 (N_3422,N_2696,N_2977);
nor U3423 (N_3423,N_2618,N_2511);
nand U3424 (N_3424,N_2670,N_2783);
nor U3425 (N_3425,N_2774,N_2657);
or U3426 (N_3426,N_2984,N_2884);
nor U3427 (N_3427,N_2815,N_2807);
or U3428 (N_3428,N_2920,N_2922);
nand U3429 (N_3429,N_2715,N_2846);
nor U3430 (N_3430,N_2839,N_2638);
nor U3431 (N_3431,N_2603,N_2983);
nor U3432 (N_3432,N_2993,N_2550);
nand U3433 (N_3433,N_2883,N_2553);
nand U3434 (N_3434,N_2584,N_2582);
nor U3435 (N_3435,N_2691,N_2519);
nand U3436 (N_3436,N_2970,N_2587);
nor U3437 (N_3437,N_2898,N_2915);
nand U3438 (N_3438,N_2842,N_2507);
xnor U3439 (N_3439,N_2827,N_2845);
nor U3440 (N_3440,N_2671,N_2565);
and U3441 (N_3441,N_2948,N_2688);
and U3442 (N_3442,N_2599,N_2759);
or U3443 (N_3443,N_2967,N_2595);
nor U3444 (N_3444,N_2920,N_2995);
or U3445 (N_3445,N_2718,N_2786);
nor U3446 (N_3446,N_2840,N_2969);
nor U3447 (N_3447,N_2627,N_2885);
nand U3448 (N_3448,N_2821,N_2586);
nor U3449 (N_3449,N_2763,N_2801);
nor U3450 (N_3450,N_2815,N_2795);
nand U3451 (N_3451,N_2892,N_2778);
nand U3452 (N_3452,N_2950,N_2705);
nor U3453 (N_3453,N_2634,N_2993);
and U3454 (N_3454,N_2765,N_2757);
and U3455 (N_3455,N_2507,N_2795);
and U3456 (N_3456,N_2989,N_2877);
nor U3457 (N_3457,N_2707,N_2816);
nand U3458 (N_3458,N_2967,N_2605);
nor U3459 (N_3459,N_2594,N_2702);
nor U3460 (N_3460,N_2882,N_2967);
xnor U3461 (N_3461,N_2517,N_2934);
xnor U3462 (N_3462,N_2621,N_2525);
and U3463 (N_3463,N_2515,N_2524);
nand U3464 (N_3464,N_2701,N_2862);
nor U3465 (N_3465,N_2605,N_2511);
and U3466 (N_3466,N_2843,N_2622);
or U3467 (N_3467,N_2825,N_2639);
or U3468 (N_3468,N_2666,N_2708);
nand U3469 (N_3469,N_2890,N_2818);
and U3470 (N_3470,N_2635,N_2769);
nor U3471 (N_3471,N_2978,N_2802);
nor U3472 (N_3472,N_2507,N_2726);
nand U3473 (N_3473,N_2565,N_2931);
and U3474 (N_3474,N_2921,N_2661);
or U3475 (N_3475,N_2916,N_2928);
and U3476 (N_3476,N_2732,N_2870);
xor U3477 (N_3477,N_2505,N_2774);
nand U3478 (N_3478,N_2923,N_2695);
xor U3479 (N_3479,N_2726,N_2926);
or U3480 (N_3480,N_2521,N_2725);
nor U3481 (N_3481,N_2919,N_2960);
nand U3482 (N_3482,N_2562,N_2891);
xnor U3483 (N_3483,N_2597,N_2537);
or U3484 (N_3484,N_2943,N_2822);
nor U3485 (N_3485,N_2778,N_2719);
and U3486 (N_3486,N_2500,N_2788);
nor U3487 (N_3487,N_2647,N_2778);
nand U3488 (N_3488,N_2829,N_2677);
nand U3489 (N_3489,N_2503,N_2687);
nor U3490 (N_3490,N_2825,N_2948);
nor U3491 (N_3491,N_2881,N_2504);
nor U3492 (N_3492,N_2746,N_2917);
or U3493 (N_3493,N_2956,N_2887);
and U3494 (N_3494,N_2937,N_2804);
nand U3495 (N_3495,N_2736,N_2833);
nand U3496 (N_3496,N_2787,N_2723);
nand U3497 (N_3497,N_2768,N_2512);
nand U3498 (N_3498,N_2936,N_2744);
and U3499 (N_3499,N_2683,N_2690);
nand U3500 (N_3500,N_3449,N_3324);
nor U3501 (N_3501,N_3327,N_3121);
and U3502 (N_3502,N_3369,N_3013);
nor U3503 (N_3503,N_3409,N_3275);
xnor U3504 (N_3504,N_3082,N_3021);
nand U3505 (N_3505,N_3264,N_3471);
or U3506 (N_3506,N_3341,N_3134);
nand U3507 (N_3507,N_3367,N_3095);
nand U3508 (N_3508,N_3238,N_3180);
or U3509 (N_3509,N_3041,N_3287);
nor U3510 (N_3510,N_3486,N_3417);
or U3511 (N_3511,N_3453,N_3339);
and U3512 (N_3512,N_3211,N_3196);
or U3513 (N_3513,N_3476,N_3316);
and U3514 (N_3514,N_3089,N_3252);
and U3515 (N_3515,N_3458,N_3485);
and U3516 (N_3516,N_3009,N_3189);
nand U3517 (N_3517,N_3410,N_3257);
nand U3518 (N_3518,N_3097,N_3260);
or U3519 (N_3519,N_3040,N_3002);
and U3520 (N_3520,N_3229,N_3261);
or U3521 (N_3521,N_3142,N_3487);
nor U3522 (N_3522,N_3284,N_3499);
nand U3523 (N_3523,N_3343,N_3191);
or U3524 (N_3524,N_3143,N_3396);
and U3525 (N_3525,N_3025,N_3430);
or U3526 (N_3526,N_3333,N_3187);
nand U3527 (N_3527,N_3387,N_3311);
nor U3528 (N_3528,N_3220,N_3145);
nand U3529 (N_3529,N_3256,N_3477);
xnor U3530 (N_3530,N_3161,N_3394);
and U3531 (N_3531,N_3182,N_3156);
or U3532 (N_3532,N_3210,N_3338);
nor U3533 (N_3533,N_3456,N_3470);
nand U3534 (N_3534,N_3459,N_3170);
or U3535 (N_3535,N_3087,N_3299);
or U3536 (N_3536,N_3362,N_3282);
and U3537 (N_3537,N_3030,N_3378);
xor U3538 (N_3538,N_3231,N_3199);
nor U3539 (N_3539,N_3334,N_3043);
and U3540 (N_3540,N_3463,N_3461);
nor U3541 (N_3541,N_3026,N_3281);
or U3542 (N_3542,N_3490,N_3091);
or U3543 (N_3543,N_3246,N_3320);
nor U3544 (N_3544,N_3107,N_3350);
or U3545 (N_3545,N_3366,N_3222);
and U3546 (N_3546,N_3176,N_3444);
nor U3547 (N_3547,N_3441,N_3266);
nand U3548 (N_3548,N_3179,N_3307);
nor U3549 (N_3549,N_3137,N_3169);
and U3550 (N_3550,N_3272,N_3151);
nand U3551 (N_3551,N_3290,N_3200);
and U3552 (N_3552,N_3186,N_3240);
and U3553 (N_3553,N_3308,N_3271);
or U3554 (N_3554,N_3132,N_3157);
nor U3555 (N_3555,N_3291,N_3072);
and U3556 (N_3556,N_3105,N_3401);
xor U3557 (N_3557,N_3206,N_3054);
and U3558 (N_3558,N_3439,N_3322);
and U3559 (N_3559,N_3152,N_3429);
nand U3560 (N_3560,N_3058,N_3475);
xnor U3561 (N_3561,N_3244,N_3276);
nor U3562 (N_3562,N_3216,N_3245);
nand U3563 (N_3563,N_3201,N_3028);
nand U3564 (N_3564,N_3313,N_3125);
nand U3565 (N_3565,N_3113,N_3269);
or U3566 (N_3566,N_3069,N_3305);
and U3567 (N_3567,N_3106,N_3076);
and U3568 (N_3568,N_3144,N_3140);
nor U3569 (N_3569,N_3436,N_3223);
nand U3570 (N_3570,N_3258,N_3138);
and U3571 (N_3571,N_3473,N_3412);
nand U3572 (N_3572,N_3133,N_3012);
and U3573 (N_3573,N_3045,N_3177);
nand U3574 (N_3574,N_3194,N_3032);
or U3575 (N_3575,N_3184,N_3359);
and U3576 (N_3576,N_3468,N_3348);
xor U3577 (N_3577,N_3329,N_3039);
and U3578 (N_3578,N_3209,N_3004);
nor U3579 (N_3579,N_3388,N_3406);
nand U3580 (N_3580,N_3024,N_3445);
xor U3581 (N_3581,N_3285,N_3126);
or U3582 (N_3582,N_3128,N_3064);
nand U3583 (N_3583,N_3168,N_3005);
nor U3584 (N_3584,N_3361,N_3314);
and U3585 (N_3585,N_3407,N_3086);
or U3586 (N_3586,N_3434,N_3044);
or U3587 (N_3587,N_3347,N_3037);
nand U3588 (N_3588,N_3047,N_3204);
xnor U3589 (N_3589,N_3131,N_3389);
nand U3590 (N_3590,N_3321,N_3274);
nand U3591 (N_3591,N_3426,N_3385);
or U3592 (N_3592,N_3268,N_3421);
nor U3593 (N_3593,N_3059,N_3093);
or U3594 (N_3594,N_3353,N_3018);
nand U3595 (N_3595,N_3263,N_3312);
xor U3596 (N_3596,N_3242,N_3014);
xor U3597 (N_3597,N_3304,N_3262);
or U3598 (N_3598,N_3099,N_3382);
nand U3599 (N_3599,N_3297,N_3249);
nand U3600 (N_3600,N_3165,N_3150);
nor U3601 (N_3601,N_3428,N_3035);
xnor U3602 (N_3602,N_3214,N_3247);
nor U3603 (N_3603,N_3104,N_3001);
nor U3604 (N_3604,N_3202,N_3413);
and U3605 (N_3605,N_3224,N_3474);
nand U3606 (N_3606,N_3363,N_3063);
and U3607 (N_3607,N_3323,N_3080);
nor U3608 (N_3608,N_3265,N_3042);
xnor U3609 (N_3609,N_3115,N_3301);
or U3610 (N_3610,N_3164,N_3495);
xor U3611 (N_3611,N_3460,N_3195);
and U3612 (N_3612,N_3478,N_3218);
and U3613 (N_3613,N_3377,N_3052);
or U3614 (N_3614,N_3055,N_3172);
and U3615 (N_3615,N_3386,N_3255);
and U3616 (N_3616,N_3491,N_3100);
and U3617 (N_3617,N_3136,N_3141);
or U3618 (N_3618,N_3267,N_3392);
nor U3619 (N_3619,N_3067,N_3494);
and U3620 (N_3620,N_3008,N_3368);
and U3621 (N_3621,N_3365,N_3425);
or U3622 (N_3622,N_3454,N_3130);
and U3623 (N_3623,N_3212,N_3090);
xnor U3624 (N_3624,N_3110,N_3102);
nand U3625 (N_3625,N_3469,N_3084);
or U3626 (N_3626,N_3124,N_3457);
nand U3627 (N_3627,N_3003,N_3451);
nor U3628 (N_3628,N_3357,N_3437);
or U3629 (N_3629,N_3480,N_3250);
or U3630 (N_3630,N_3390,N_3081);
or U3631 (N_3631,N_3167,N_3198);
nand U3632 (N_3632,N_3455,N_3158);
and U3633 (N_3633,N_3472,N_3007);
nor U3634 (N_3634,N_3162,N_3112);
or U3635 (N_3635,N_3057,N_3315);
or U3636 (N_3636,N_3411,N_3029);
and U3637 (N_3637,N_3402,N_3356);
nand U3638 (N_3638,N_3225,N_3354);
and U3639 (N_3639,N_3330,N_3020);
nor U3640 (N_3640,N_3497,N_3479);
or U3641 (N_3641,N_3062,N_3006);
and U3642 (N_3642,N_3336,N_3375);
or U3643 (N_3643,N_3424,N_3217);
and U3644 (N_3644,N_3318,N_3443);
nand U3645 (N_3645,N_3283,N_3419);
or U3646 (N_3646,N_3160,N_3237);
or U3647 (N_3647,N_3109,N_3228);
nand U3648 (N_3648,N_3418,N_3060);
nor U3649 (N_3649,N_3450,N_3391);
nor U3650 (N_3650,N_3482,N_3071);
nand U3651 (N_3651,N_3015,N_3226);
and U3652 (N_3652,N_3349,N_3023);
xnor U3653 (N_3653,N_3203,N_3061);
or U3654 (N_3654,N_3483,N_3163);
or U3655 (N_3655,N_3467,N_3351);
nor U3656 (N_3656,N_3033,N_3292);
and U3657 (N_3657,N_3075,N_3118);
nand U3658 (N_3658,N_3448,N_3493);
or U3659 (N_3659,N_3383,N_3416);
and U3660 (N_3660,N_3066,N_3098);
and U3661 (N_3661,N_3345,N_3219);
nor U3662 (N_3662,N_3122,N_3384);
and U3663 (N_3663,N_3337,N_3233);
nor U3664 (N_3664,N_3079,N_3360);
and U3665 (N_3665,N_3358,N_3155);
and U3666 (N_3666,N_3447,N_3254);
or U3667 (N_3667,N_3481,N_3036);
and U3668 (N_3668,N_3300,N_3465);
xnor U3669 (N_3669,N_3031,N_3498);
or U3670 (N_3670,N_3193,N_3174);
xnor U3671 (N_3671,N_3440,N_3153);
and U3672 (N_3672,N_3293,N_3022);
nand U3673 (N_3673,N_3395,N_3294);
nor U3674 (N_3674,N_3248,N_3065);
nand U3675 (N_3675,N_3046,N_3011);
nor U3676 (N_3676,N_3068,N_3146);
xnor U3677 (N_3677,N_3302,N_3352);
nand U3678 (N_3678,N_3114,N_3370);
and U3679 (N_3679,N_3096,N_3074);
and U3680 (N_3680,N_3148,N_3117);
or U3681 (N_3681,N_3403,N_3317);
and U3682 (N_3682,N_3295,N_3178);
nor U3683 (N_3683,N_3017,N_3000);
nand U3684 (N_3684,N_3446,N_3078);
nand U3685 (N_3685,N_3306,N_3408);
nor U3686 (N_3686,N_3108,N_3332);
and U3687 (N_3687,N_3135,N_3119);
and U3688 (N_3688,N_3423,N_3371);
nor U3689 (N_3689,N_3346,N_3259);
and U3690 (N_3690,N_3123,N_3380);
and U3691 (N_3691,N_3038,N_3056);
or U3692 (N_3692,N_3192,N_3239);
or U3693 (N_3693,N_3175,N_3399);
or U3694 (N_3694,N_3373,N_3232);
nand U3695 (N_3695,N_3234,N_3432);
xnor U3696 (N_3696,N_3435,N_3207);
or U3697 (N_3697,N_3205,N_3414);
nand U3698 (N_3698,N_3221,N_3235);
xor U3699 (N_3699,N_3464,N_3325);
nand U3700 (N_3700,N_3073,N_3438);
nand U3701 (N_3701,N_3111,N_3227);
or U3702 (N_3702,N_3376,N_3273);
nand U3703 (N_3703,N_3088,N_3083);
nand U3704 (N_3704,N_3364,N_3215);
nor U3705 (N_3705,N_3277,N_3070);
nand U3706 (N_3706,N_3326,N_3303);
or U3707 (N_3707,N_3094,N_3253);
or U3708 (N_3708,N_3050,N_3027);
and U3709 (N_3709,N_3496,N_3053);
nand U3710 (N_3710,N_3484,N_3236);
and U3711 (N_3711,N_3101,N_3185);
or U3712 (N_3712,N_3181,N_3335);
xnor U3713 (N_3713,N_3139,N_3116);
or U3714 (N_3714,N_3188,N_3309);
and U3715 (N_3715,N_3280,N_3298);
nor U3716 (N_3716,N_3420,N_3466);
nand U3717 (N_3717,N_3149,N_3415);
nand U3718 (N_3718,N_3288,N_3379);
and U3719 (N_3719,N_3173,N_3230);
and U3720 (N_3720,N_3278,N_3279);
nand U3721 (N_3721,N_3492,N_3355);
and U3722 (N_3722,N_3400,N_3286);
nor U3723 (N_3723,N_3019,N_3374);
nor U3724 (N_3724,N_3340,N_3296);
nand U3725 (N_3725,N_3289,N_3489);
xnor U3726 (N_3726,N_3010,N_3422);
xnor U3727 (N_3727,N_3452,N_3344);
and U3728 (N_3728,N_3319,N_3120);
or U3729 (N_3729,N_3251,N_3433);
or U3730 (N_3730,N_3398,N_3016);
nor U3731 (N_3731,N_3488,N_3183);
nand U3732 (N_3732,N_3310,N_3328);
and U3733 (N_3733,N_3034,N_3342);
nand U3734 (N_3734,N_3243,N_3190);
or U3735 (N_3735,N_3171,N_3213);
and U3736 (N_3736,N_3208,N_3372);
nand U3737 (N_3737,N_3159,N_3381);
and U3738 (N_3738,N_3462,N_3154);
nor U3739 (N_3739,N_3241,N_3127);
nand U3740 (N_3740,N_3431,N_3051);
xnor U3741 (N_3741,N_3393,N_3397);
or U3742 (N_3742,N_3442,N_3331);
and U3743 (N_3743,N_3049,N_3103);
xor U3744 (N_3744,N_3166,N_3270);
or U3745 (N_3745,N_3147,N_3129);
nand U3746 (N_3746,N_3197,N_3048);
and U3747 (N_3747,N_3427,N_3077);
xor U3748 (N_3748,N_3092,N_3404);
nand U3749 (N_3749,N_3085,N_3405);
nor U3750 (N_3750,N_3194,N_3415);
and U3751 (N_3751,N_3236,N_3377);
or U3752 (N_3752,N_3413,N_3264);
nand U3753 (N_3753,N_3491,N_3121);
nand U3754 (N_3754,N_3317,N_3322);
nand U3755 (N_3755,N_3266,N_3052);
nand U3756 (N_3756,N_3471,N_3177);
xor U3757 (N_3757,N_3146,N_3057);
xor U3758 (N_3758,N_3090,N_3305);
or U3759 (N_3759,N_3487,N_3337);
and U3760 (N_3760,N_3462,N_3417);
and U3761 (N_3761,N_3388,N_3195);
or U3762 (N_3762,N_3454,N_3318);
nand U3763 (N_3763,N_3260,N_3356);
and U3764 (N_3764,N_3094,N_3129);
and U3765 (N_3765,N_3409,N_3332);
or U3766 (N_3766,N_3218,N_3107);
or U3767 (N_3767,N_3459,N_3439);
and U3768 (N_3768,N_3458,N_3370);
or U3769 (N_3769,N_3126,N_3358);
nand U3770 (N_3770,N_3044,N_3413);
or U3771 (N_3771,N_3159,N_3163);
xnor U3772 (N_3772,N_3061,N_3040);
xor U3773 (N_3773,N_3474,N_3068);
nand U3774 (N_3774,N_3004,N_3061);
or U3775 (N_3775,N_3113,N_3323);
or U3776 (N_3776,N_3293,N_3124);
or U3777 (N_3777,N_3470,N_3009);
or U3778 (N_3778,N_3492,N_3212);
or U3779 (N_3779,N_3270,N_3402);
xor U3780 (N_3780,N_3490,N_3332);
and U3781 (N_3781,N_3426,N_3230);
nor U3782 (N_3782,N_3019,N_3368);
or U3783 (N_3783,N_3120,N_3307);
or U3784 (N_3784,N_3493,N_3449);
nor U3785 (N_3785,N_3278,N_3018);
xor U3786 (N_3786,N_3205,N_3335);
and U3787 (N_3787,N_3413,N_3330);
and U3788 (N_3788,N_3413,N_3144);
nor U3789 (N_3789,N_3107,N_3276);
nor U3790 (N_3790,N_3017,N_3348);
and U3791 (N_3791,N_3406,N_3109);
nor U3792 (N_3792,N_3216,N_3139);
or U3793 (N_3793,N_3294,N_3114);
and U3794 (N_3794,N_3294,N_3388);
nor U3795 (N_3795,N_3047,N_3259);
nor U3796 (N_3796,N_3045,N_3038);
nor U3797 (N_3797,N_3340,N_3349);
xor U3798 (N_3798,N_3124,N_3248);
nor U3799 (N_3799,N_3185,N_3305);
nor U3800 (N_3800,N_3322,N_3031);
nor U3801 (N_3801,N_3377,N_3319);
nand U3802 (N_3802,N_3295,N_3433);
xnor U3803 (N_3803,N_3222,N_3324);
nor U3804 (N_3804,N_3064,N_3332);
nand U3805 (N_3805,N_3364,N_3204);
nand U3806 (N_3806,N_3404,N_3486);
nand U3807 (N_3807,N_3281,N_3452);
nand U3808 (N_3808,N_3464,N_3193);
or U3809 (N_3809,N_3252,N_3021);
xnor U3810 (N_3810,N_3184,N_3478);
or U3811 (N_3811,N_3025,N_3371);
nand U3812 (N_3812,N_3104,N_3455);
or U3813 (N_3813,N_3179,N_3193);
nand U3814 (N_3814,N_3396,N_3493);
and U3815 (N_3815,N_3009,N_3144);
nand U3816 (N_3816,N_3026,N_3158);
or U3817 (N_3817,N_3324,N_3321);
nor U3818 (N_3818,N_3283,N_3111);
and U3819 (N_3819,N_3247,N_3317);
and U3820 (N_3820,N_3339,N_3099);
and U3821 (N_3821,N_3431,N_3059);
nand U3822 (N_3822,N_3480,N_3434);
or U3823 (N_3823,N_3486,N_3406);
and U3824 (N_3824,N_3339,N_3363);
and U3825 (N_3825,N_3405,N_3421);
xor U3826 (N_3826,N_3114,N_3364);
nor U3827 (N_3827,N_3179,N_3249);
nand U3828 (N_3828,N_3057,N_3183);
nor U3829 (N_3829,N_3100,N_3066);
nand U3830 (N_3830,N_3248,N_3307);
and U3831 (N_3831,N_3182,N_3439);
nor U3832 (N_3832,N_3081,N_3067);
and U3833 (N_3833,N_3112,N_3471);
nand U3834 (N_3834,N_3337,N_3364);
nor U3835 (N_3835,N_3240,N_3161);
nand U3836 (N_3836,N_3412,N_3213);
nand U3837 (N_3837,N_3093,N_3052);
nand U3838 (N_3838,N_3265,N_3244);
or U3839 (N_3839,N_3339,N_3224);
nand U3840 (N_3840,N_3274,N_3471);
xor U3841 (N_3841,N_3192,N_3111);
nand U3842 (N_3842,N_3002,N_3452);
or U3843 (N_3843,N_3302,N_3038);
xnor U3844 (N_3844,N_3248,N_3050);
xor U3845 (N_3845,N_3416,N_3040);
nand U3846 (N_3846,N_3490,N_3219);
or U3847 (N_3847,N_3228,N_3468);
nor U3848 (N_3848,N_3337,N_3457);
or U3849 (N_3849,N_3222,N_3094);
nor U3850 (N_3850,N_3119,N_3301);
and U3851 (N_3851,N_3109,N_3121);
or U3852 (N_3852,N_3262,N_3231);
nor U3853 (N_3853,N_3237,N_3268);
nand U3854 (N_3854,N_3346,N_3250);
nand U3855 (N_3855,N_3379,N_3327);
nor U3856 (N_3856,N_3174,N_3444);
and U3857 (N_3857,N_3055,N_3103);
nor U3858 (N_3858,N_3481,N_3338);
or U3859 (N_3859,N_3304,N_3457);
nor U3860 (N_3860,N_3087,N_3352);
or U3861 (N_3861,N_3163,N_3472);
and U3862 (N_3862,N_3364,N_3349);
nand U3863 (N_3863,N_3211,N_3181);
nand U3864 (N_3864,N_3289,N_3334);
and U3865 (N_3865,N_3322,N_3303);
or U3866 (N_3866,N_3213,N_3015);
and U3867 (N_3867,N_3109,N_3105);
nor U3868 (N_3868,N_3402,N_3380);
nand U3869 (N_3869,N_3426,N_3177);
nor U3870 (N_3870,N_3417,N_3473);
nor U3871 (N_3871,N_3294,N_3110);
and U3872 (N_3872,N_3023,N_3330);
nand U3873 (N_3873,N_3488,N_3265);
and U3874 (N_3874,N_3292,N_3313);
and U3875 (N_3875,N_3010,N_3037);
or U3876 (N_3876,N_3117,N_3449);
and U3877 (N_3877,N_3323,N_3437);
nand U3878 (N_3878,N_3301,N_3017);
and U3879 (N_3879,N_3297,N_3472);
nand U3880 (N_3880,N_3134,N_3057);
or U3881 (N_3881,N_3308,N_3310);
and U3882 (N_3882,N_3074,N_3448);
nor U3883 (N_3883,N_3452,N_3339);
nand U3884 (N_3884,N_3399,N_3112);
nand U3885 (N_3885,N_3430,N_3008);
and U3886 (N_3886,N_3340,N_3148);
nor U3887 (N_3887,N_3331,N_3202);
and U3888 (N_3888,N_3211,N_3339);
nand U3889 (N_3889,N_3047,N_3494);
nand U3890 (N_3890,N_3095,N_3057);
nor U3891 (N_3891,N_3163,N_3305);
or U3892 (N_3892,N_3417,N_3322);
nor U3893 (N_3893,N_3426,N_3192);
nor U3894 (N_3894,N_3383,N_3059);
and U3895 (N_3895,N_3368,N_3326);
xnor U3896 (N_3896,N_3465,N_3247);
nor U3897 (N_3897,N_3207,N_3043);
xnor U3898 (N_3898,N_3181,N_3134);
nand U3899 (N_3899,N_3279,N_3395);
or U3900 (N_3900,N_3479,N_3037);
and U3901 (N_3901,N_3425,N_3179);
and U3902 (N_3902,N_3098,N_3331);
nor U3903 (N_3903,N_3358,N_3298);
or U3904 (N_3904,N_3337,N_3093);
nor U3905 (N_3905,N_3258,N_3158);
nor U3906 (N_3906,N_3427,N_3079);
and U3907 (N_3907,N_3019,N_3159);
or U3908 (N_3908,N_3444,N_3255);
nor U3909 (N_3909,N_3007,N_3017);
and U3910 (N_3910,N_3281,N_3190);
nand U3911 (N_3911,N_3446,N_3332);
and U3912 (N_3912,N_3082,N_3004);
nor U3913 (N_3913,N_3116,N_3343);
or U3914 (N_3914,N_3440,N_3141);
or U3915 (N_3915,N_3472,N_3185);
and U3916 (N_3916,N_3226,N_3377);
or U3917 (N_3917,N_3322,N_3402);
xnor U3918 (N_3918,N_3489,N_3100);
or U3919 (N_3919,N_3072,N_3227);
and U3920 (N_3920,N_3294,N_3025);
or U3921 (N_3921,N_3128,N_3206);
nor U3922 (N_3922,N_3462,N_3287);
and U3923 (N_3923,N_3358,N_3156);
nor U3924 (N_3924,N_3038,N_3058);
nor U3925 (N_3925,N_3211,N_3124);
or U3926 (N_3926,N_3087,N_3434);
or U3927 (N_3927,N_3177,N_3318);
nor U3928 (N_3928,N_3296,N_3353);
nor U3929 (N_3929,N_3145,N_3080);
nor U3930 (N_3930,N_3007,N_3191);
xor U3931 (N_3931,N_3360,N_3347);
and U3932 (N_3932,N_3162,N_3387);
xor U3933 (N_3933,N_3419,N_3480);
nor U3934 (N_3934,N_3207,N_3208);
nand U3935 (N_3935,N_3470,N_3127);
and U3936 (N_3936,N_3442,N_3348);
or U3937 (N_3937,N_3076,N_3406);
nor U3938 (N_3938,N_3120,N_3114);
and U3939 (N_3939,N_3471,N_3020);
nand U3940 (N_3940,N_3243,N_3290);
nor U3941 (N_3941,N_3286,N_3385);
xor U3942 (N_3942,N_3246,N_3374);
nor U3943 (N_3943,N_3326,N_3030);
or U3944 (N_3944,N_3221,N_3319);
or U3945 (N_3945,N_3275,N_3090);
nor U3946 (N_3946,N_3271,N_3103);
nor U3947 (N_3947,N_3415,N_3483);
and U3948 (N_3948,N_3215,N_3476);
nand U3949 (N_3949,N_3253,N_3106);
xnor U3950 (N_3950,N_3130,N_3453);
nor U3951 (N_3951,N_3458,N_3363);
or U3952 (N_3952,N_3075,N_3256);
and U3953 (N_3953,N_3106,N_3236);
or U3954 (N_3954,N_3311,N_3102);
or U3955 (N_3955,N_3082,N_3195);
nand U3956 (N_3956,N_3177,N_3411);
nand U3957 (N_3957,N_3076,N_3428);
nand U3958 (N_3958,N_3317,N_3121);
and U3959 (N_3959,N_3356,N_3330);
nand U3960 (N_3960,N_3140,N_3175);
nor U3961 (N_3961,N_3087,N_3353);
and U3962 (N_3962,N_3389,N_3430);
and U3963 (N_3963,N_3005,N_3416);
and U3964 (N_3964,N_3052,N_3000);
nor U3965 (N_3965,N_3358,N_3102);
xor U3966 (N_3966,N_3453,N_3389);
nor U3967 (N_3967,N_3328,N_3332);
and U3968 (N_3968,N_3043,N_3402);
nor U3969 (N_3969,N_3420,N_3281);
nand U3970 (N_3970,N_3484,N_3474);
or U3971 (N_3971,N_3258,N_3124);
and U3972 (N_3972,N_3466,N_3110);
xnor U3973 (N_3973,N_3294,N_3422);
nor U3974 (N_3974,N_3163,N_3086);
or U3975 (N_3975,N_3113,N_3103);
and U3976 (N_3976,N_3087,N_3392);
or U3977 (N_3977,N_3147,N_3440);
nand U3978 (N_3978,N_3323,N_3124);
and U3979 (N_3979,N_3170,N_3134);
nand U3980 (N_3980,N_3124,N_3253);
or U3981 (N_3981,N_3042,N_3069);
nor U3982 (N_3982,N_3133,N_3342);
nor U3983 (N_3983,N_3382,N_3136);
nand U3984 (N_3984,N_3076,N_3088);
and U3985 (N_3985,N_3029,N_3413);
xnor U3986 (N_3986,N_3273,N_3380);
and U3987 (N_3987,N_3082,N_3094);
nand U3988 (N_3988,N_3371,N_3120);
or U3989 (N_3989,N_3411,N_3125);
nand U3990 (N_3990,N_3405,N_3038);
nand U3991 (N_3991,N_3307,N_3353);
nor U3992 (N_3992,N_3463,N_3340);
or U3993 (N_3993,N_3205,N_3407);
nand U3994 (N_3994,N_3217,N_3463);
and U3995 (N_3995,N_3388,N_3472);
nor U3996 (N_3996,N_3211,N_3388);
xor U3997 (N_3997,N_3322,N_3345);
nand U3998 (N_3998,N_3387,N_3189);
xor U3999 (N_3999,N_3246,N_3214);
nor U4000 (N_4000,N_3993,N_3572);
or U4001 (N_4001,N_3650,N_3913);
or U4002 (N_4002,N_3938,N_3796);
or U4003 (N_4003,N_3700,N_3826);
xnor U4004 (N_4004,N_3897,N_3620);
nand U4005 (N_4005,N_3995,N_3561);
xnor U4006 (N_4006,N_3854,N_3887);
and U4007 (N_4007,N_3668,N_3847);
or U4008 (N_4008,N_3922,N_3708);
nor U4009 (N_4009,N_3767,N_3905);
and U4010 (N_4010,N_3698,N_3825);
nand U4011 (N_4011,N_3912,N_3657);
nor U4012 (N_4012,N_3630,N_3602);
nand U4013 (N_4013,N_3859,N_3762);
nand U4014 (N_4014,N_3637,N_3635);
nand U4015 (N_4015,N_3643,N_3879);
xnor U4016 (N_4016,N_3516,N_3975);
nor U4017 (N_4017,N_3638,N_3576);
nand U4018 (N_4018,N_3895,N_3678);
or U4019 (N_4019,N_3838,N_3794);
nor U4020 (N_4020,N_3896,N_3935);
nand U4021 (N_4021,N_3866,N_3661);
nand U4022 (N_4022,N_3961,N_3660);
or U4023 (N_4023,N_3687,N_3501);
nor U4024 (N_4024,N_3754,N_3998);
or U4025 (N_4025,N_3969,N_3776);
nor U4026 (N_4026,N_3758,N_3565);
nand U4027 (N_4027,N_3505,N_3552);
xnor U4028 (N_4028,N_3985,N_3503);
nand U4029 (N_4029,N_3590,N_3931);
and U4030 (N_4030,N_3760,N_3679);
xor U4031 (N_4031,N_3894,N_3682);
nand U4032 (N_4032,N_3528,N_3514);
nand U4033 (N_4033,N_3622,N_3951);
nand U4034 (N_4034,N_3560,N_3535);
nand U4035 (N_4035,N_3783,N_3818);
nor U4036 (N_4036,N_3915,N_3612);
nor U4037 (N_4037,N_3671,N_3792);
or U4038 (N_4038,N_3753,N_3672);
nand U4039 (N_4039,N_3613,N_3833);
nand U4040 (N_4040,N_3828,N_3936);
xnor U4041 (N_4041,N_3947,N_3869);
nand U4042 (N_4042,N_3717,N_3569);
nor U4043 (N_4043,N_3997,N_3734);
nand U4044 (N_4044,N_3556,N_3709);
nand U4045 (N_4045,N_3846,N_3524);
or U4046 (N_4046,N_3750,N_3759);
and U4047 (N_4047,N_3621,N_3581);
nor U4048 (N_4048,N_3730,N_3903);
or U4049 (N_4049,N_3521,N_3566);
and U4050 (N_4050,N_3604,N_3674);
xnor U4051 (N_4051,N_3761,N_3603);
or U4052 (N_4052,N_3600,N_3864);
nor U4053 (N_4053,N_3536,N_3523);
nor U4054 (N_4054,N_3970,N_3712);
nor U4055 (N_4055,N_3964,N_3858);
nand U4056 (N_4056,N_3878,N_3738);
and U4057 (N_4057,N_3551,N_3898);
nor U4058 (N_4058,N_3723,N_3929);
or U4059 (N_4059,N_3800,N_3808);
nand U4060 (N_4060,N_3959,N_3667);
and U4061 (N_4061,N_3704,N_3763);
xor U4062 (N_4062,N_3651,N_3865);
and U4063 (N_4063,N_3525,N_3824);
and U4064 (N_4064,N_3507,N_3699);
and U4065 (N_4065,N_3795,N_3706);
nand U4066 (N_4066,N_3876,N_3749);
xnor U4067 (N_4067,N_3948,N_3537);
nor U4068 (N_4068,N_3790,N_3954);
xor U4069 (N_4069,N_3670,N_3862);
xnor U4070 (N_4070,N_3733,N_3740);
and U4071 (N_4071,N_3798,N_3558);
and U4072 (N_4072,N_3557,N_3930);
or U4073 (N_4073,N_3748,N_3933);
nand U4074 (N_4074,N_3583,N_3577);
and U4075 (N_4075,N_3914,N_3520);
and U4076 (N_4076,N_3909,N_3618);
and U4077 (N_4077,N_3889,N_3665);
nand U4078 (N_4078,N_3570,N_3724);
and U4079 (N_4079,N_3703,N_3980);
nor U4080 (N_4080,N_3873,N_3967);
and U4081 (N_4081,N_3949,N_3982);
nand U4082 (N_4082,N_3787,N_3739);
or U4083 (N_4083,N_3777,N_3968);
nand U4084 (N_4084,N_3647,N_3844);
nor U4085 (N_4085,N_3908,N_3564);
nor U4086 (N_4086,N_3764,N_3628);
nor U4087 (N_4087,N_3918,N_3868);
and U4088 (N_4088,N_3882,N_3591);
and U4089 (N_4089,N_3770,N_3606);
nor U4090 (N_4090,N_3685,N_3953);
or U4091 (N_4091,N_3680,N_3751);
nand U4092 (N_4092,N_3715,N_3927);
nand U4093 (N_4093,N_3956,N_3546);
and U4094 (N_4094,N_3595,N_3994);
and U4095 (N_4095,N_3735,N_3654);
nor U4096 (N_4096,N_3957,N_3626);
and U4097 (N_4097,N_3989,N_3928);
nand U4098 (N_4098,N_3834,N_3966);
and U4099 (N_4099,N_3639,N_3642);
nand U4100 (N_4100,N_3999,N_3852);
or U4101 (N_4101,N_3599,N_3744);
or U4102 (N_4102,N_3702,N_3554);
or U4103 (N_4103,N_3863,N_3568);
or U4104 (N_4104,N_3973,N_3526);
or U4105 (N_4105,N_3979,N_3944);
nand U4106 (N_4106,N_3529,N_3555);
and U4107 (N_4107,N_3977,N_3900);
xnor U4108 (N_4108,N_3511,N_3815);
or U4109 (N_4109,N_3644,N_3745);
and U4110 (N_4110,N_3666,N_3904);
nand U4111 (N_4111,N_3884,N_3585);
nor U4112 (N_4112,N_3856,N_3901);
and U4113 (N_4113,N_3534,N_3769);
and U4114 (N_4114,N_3669,N_3710);
nor U4115 (N_4115,N_3885,N_3640);
nor U4116 (N_4116,N_3544,N_3788);
nor U4117 (N_4117,N_3586,N_3701);
or U4118 (N_4118,N_3713,N_3648);
and U4119 (N_4119,N_3737,N_3881);
and U4120 (N_4120,N_3874,N_3832);
nor U4121 (N_4121,N_3519,N_3821);
or U4122 (N_4122,N_3504,N_3579);
or U4123 (N_4123,N_3725,N_3593);
and U4124 (N_4124,N_3742,N_3939);
nand U4125 (N_4125,N_3906,N_3571);
or U4126 (N_4126,N_3624,N_3976);
xnor U4127 (N_4127,N_3728,N_3786);
or U4128 (N_4128,N_3817,N_3924);
nor U4129 (N_4129,N_3890,N_3587);
nand U4130 (N_4130,N_3752,N_3946);
xnor U4131 (N_4131,N_3731,N_3765);
and U4132 (N_4132,N_3594,N_3871);
nand U4133 (N_4133,N_3925,N_3988);
nand U4134 (N_4134,N_3664,N_3515);
or U4135 (N_4135,N_3950,N_3646);
xor U4136 (N_4136,N_3848,N_3797);
nor U4137 (N_4137,N_3598,N_3681);
nor U4138 (N_4138,N_3697,N_3799);
and U4139 (N_4139,N_3517,N_3827);
or U4140 (N_4140,N_3958,N_3610);
nor U4141 (N_4141,N_3553,N_3992);
nand U4142 (N_4142,N_3645,N_3836);
or U4143 (N_4143,N_3839,N_3690);
nor U4144 (N_4144,N_3575,N_3766);
and U4145 (N_4145,N_3996,N_3963);
and U4146 (N_4146,N_3527,N_3789);
or U4147 (N_4147,N_3867,N_3907);
or U4148 (N_4148,N_3563,N_3542);
and U4149 (N_4149,N_3804,N_3607);
nor U4150 (N_4150,N_3711,N_3778);
xnor U4151 (N_4151,N_3716,N_3849);
or U4152 (N_4152,N_3893,N_3960);
nor U4153 (N_4153,N_3802,N_3853);
or U4154 (N_4154,N_3965,N_3722);
nand U4155 (N_4155,N_3589,N_3781);
and U4156 (N_4156,N_3785,N_3978);
or U4157 (N_4157,N_3616,N_3549);
nor U4158 (N_4158,N_3746,N_3851);
nand U4159 (N_4159,N_3676,N_3793);
or U4160 (N_4160,N_3509,N_3510);
nand U4161 (N_4161,N_3803,N_3806);
or U4162 (N_4162,N_3580,N_3653);
and U4163 (N_4163,N_3972,N_3810);
nor U4164 (N_4164,N_3574,N_3983);
nor U4165 (N_4165,N_3842,N_3513);
and U4166 (N_4166,N_3736,N_3823);
xnor U4167 (N_4167,N_3943,N_3771);
nor U4168 (N_4168,N_3926,N_3531);
and U4169 (N_4169,N_3741,N_3633);
nor U4170 (N_4170,N_3855,N_3619);
nand U4171 (N_4171,N_3605,N_3693);
nor U4172 (N_4172,N_3608,N_3872);
nand U4173 (N_4173,N_3518,N_3780);
nand U4174 (N_4174,N_3691,N_3615);
or U4175 (N_4175,N_3902,N_3541);
nor U4176 (N_4176,N_3841,N_3923);
or U4177 (N_4177,N_3756,N_3934);
and U4178 (N_4178,N_3952,N_3910);
nor U4179 (N_4179,N_3562,N_3782);
nor U4180 (N_4180,N_3784,N_3632);
nor U4181 (N_4181,N_3625,N_3942);
nor U4182 (N_4182,N_3683,N_3719);
nand U4183 (N_4183,N_3811,N_3636);
and U4184 (N_4184,N_3677,N_3870);
nand U4185 (N_4185,N_3688,N_3547);
and U4186 (N_4186,N_3631,N_3920);
xnor U4187 (N_4187,N_3649,N_3861);
or U4188 (N_4188,N_3837,N_3512);
or U4189 (N_4189,N_3888,N_3659);
and U4190 (N_4190,N_3538,N_3533);
and U4191 (N_4191,N_3500,N_3506);
xnor U4192 (N_4192,N_3831,N_3860);
or U4193 (N_4193,N_3609,N_3582);
and U4194 (N_4194,N_3601,N_3981);
nor U4195 (N_4195,N_3816,N_3508);
nor U4196 (N_4196,N_3809,N_3641);
nand U4197 (N_4197,N_3550,N_3886);
nand U4198 (N_4198,N_3791,N_3774);
and U4199 (N_4199,N_3768,N_3692);
or U4200 (N_4200,N_3921,N_3658);
nor U4201 (N_4201,N_3592,N_3801);
and U4202 (N_4202,N_3718,N_3617);
nand U4203 (N_4203,N_3892,N_3974);
or U4204 (N_4204,N_3614,N_3578);
or U4205 (N_4205,N_3727,N_3689);
nand U4206 (N_4206,N_3757,N_3559);
nand U4207 (N_4207,N_3911,N_3629);
nor U4208 (N_4208,N_3850,N_3627);
or U4209 (N_4209,N_3655,N_3813);
or U4210 (N_4210,N_3819,N_3812);
xor U4211 (N_4211,N_3991,N_3721);
and U4212 (N_4212,N_3597,N_3880);
or U4213 (N_4213,N_3729,N_3843);
or U4214 (N_4214,N_3707,N_3984);
nand U4215 (N_4215,N_3623,N_3845);
or U4216 (N_4216,N_3945,N_3899);
nor U4217 (N_4217,N_3772,N_3596);
nand U4218 (N_4218,N_3540,N_3611);
nand U4219 (N_4219,N_3805,N_3696);
and U4220 (N_4220,N_3971,N_3675);
nor U4221 (N_4221,N_3726,N_3916);
and U4222 (N_4222,N_3877,N_3705);
and U4223 (N_4223,N_3530,N_3932);
nor U4224 (N_4224,N_3857,N_3941);
or U4225 (N_4225,N_3955,N_3673);
xnor U4226 (N_4226,N_3695,N_3652);
and U4227 (N_4227,N_3714,N_3990);
nor U4228 (N_4228,N_3743,N_3584);
nand U4229 (N_4229,N_3662,N_3684);
or U4230 (N_4230,N_3835,N_3891);
nand U4231 (N_4231,N_3875,N_3548);
nand U4232 (N_4232,N_3775,N_3694);
or U4233 (N_4233,N_3634,N_3807);
nor U4234 (N_4234,N_3883,N_3573);
xnor U4235 (N_4235,N_3522,N_3937);
or U4236 (N_4236,N_3940,N_3830);
xor U4237 (N_4237,N_3539,N_3543);
and U4238 (N_4238,N_3567,N_3656);
or U4239 (N_4239,N_3773,N_3917);
nand U4240 (N_4240,N_3502,N_3820);
nor U4241 (N_4241,N_3732,N_3663);
xor U4242 (N_4242,N_3919,N_3686);
nand U4243 (N_4243,N_3814,N_3840);
nand U4244 (N_4244,N_3986,N_3779);
xnor U4245 (N_4245,N_3755,N_3822);
nand U4246 (N_4246,N_3987,N_3532);
nor U4247 (N_4247,N_3720,N_3829);
nand U4248 (N_4248,N_3545,N_3747);
xnor U4249 (N_4249,N_3588,N_3962);
or U4250 (N_4250,N_3593,N_3738);
nor U4251 (N_4251,N_3571,N_3749);
nand U4252 (N_4252,N_3687,N_3904);
or U4253 (N_4253,N_3594,N_3838);
nand U4254 (N_4254,N_3603,N_3938);
or U4255 (N_4255,N_3512,N_3606);
nor U4256 (N_4256,N_3658,N_3996);
and U4257 (N_4257,N_3587,N_3782);
or U4258 (N_4258,N_3549,N_3553);
and U4259 (N_4259,N_3994,N_3696);
or U4260 (N_4260,N_3784,N_3562);
nor U4261 (N_4261,N_3802,N_3640);
nand U4262 (N_4262,N_3989,N_3746);
or U4263 (N_4263,N_3982,N_3945);
nand U4264 (N_4264,N_3790,N_3528);
and U4265 (N_4265,N_3571,N_3648);
nand U4266 (N_4266,N_3987,N_3518);
or U4267 (N_4267,N_3518,N_3623);
or U4268 (N_4268,N_3989,N_3901);
nand U4269 (N_4269,N_3961,N_3511);
or U4270 (N_4270,N_3681,N_3553);
and U4271 (N_4271,N_3950,N_3783);
or U4272 (N_4272,N_3907,N_3753);
xnor U4273 (N_4273,N_3773,N_3953);
or U4274 (N_4274,N_3807,N_3893);
and U4275 (N_4275,N_3579,N_3852);
nand U4276 (N_4276,N_3764,N_3983);
nand U4277 (N_4277,N_3755,N_3624);
or U4278 (N_4278,N_3553,N_3647);
nor U4279 (N_4279,N_3788,N_3976);
xnor U4280 (N_4280,N_3891,N_3700);
nor U4281 (N_4281,N_3704,N_3555);
and U4282 (N_4282,N_3850,N_3653);
nor U4283 (N_4283,N_3578,N_3739);
and U4284 (N_4284,N_3843,N_3967);
nand U4285 (N_4285,N_3580,N_3750);
nand U4286 (N_4286,N_3714,N_3735);
nand U4287 (N_4287,N_3867,N_3589);
nand U4288 (N_4288,N_3606,N_3824);
nand U4289 (N_4289,N_3853,N_3941);
nand U4290 (N_4290,N_3765,N_3993);
nand U4291 (N_4291,N_3584,N_3720);
nand U4292 (N_4292,N_3584,N_3645);
nor U4293 (N_4293,N_3785,N_3716);
and U4294 (N_4294,N_3789,N_3926);
nor U4295 (N_4295,N_3827,N_3857);
nand U4296 (N_4296,N_3687,N_3629);
nor U4297 (N_4297,N_3809,N_3814);
nand U4298 (N_4298,N_3605,N_3986);
nand U4299 (N_4299,N_3529,N_3895);
or U4300 (N_4300,N_3605,N_3671);
and U4301 (N_4301,N_3951,N_3957);
xor U4302 (N_4302,N_3980,N_3992);
or U4303 (N_4303,N_3672,N_3679);
or U4304 (N_4304,N_3747,N_3562);
or U4305 (N_4305,N_3931,N_3963);
nand U4306 (N_4306,N_3533,N_3556);
nand U4307 (N_4307,N_3675,N_3842);
and U4308 (N_4308,N_3550,N_3855);
or U4309 (N_4309,N_3502,N_3971);
nand U4310 (N_4310,N_3596,N_3714);
nor U4311 (N_4311,N_3700,N_3978);
and U4312 (N_4312,N_3638,N_3599);
xnor U4313 (N_4313,N_3701,N_3904);
and U4314 (N_4314,N_3617,N_3937);
or U4315 (N_4315,N_3803,N_3593);
or U4316 (N_4316,N_3996,N_3853);
and U4317 (N_4317,N_3907,N_3786);
nand U4318 (N_4318,N_3928,N_3798);
xor U4319 (N_4319,N_3585,N_3847);
nand U4320 (N_4320,N_3959,N_3885);
nor U4321 (N_4321,N_3955,N_3755);
nor U4322 (N_4322,N_3794,N_3964);
nor U4323 (N_4323,N_3574,N_3938);
nor U4324 (N_4324,N_3874,N_3736);
nand U4325 (N_4325,N_3720,N_3655);
nor U4326 (N_4326,N_3569,N_3699);
xnor U4327 (N_4327,N_3621,N_3555);
nand U4328 (N_4328,N_3903,N_3580);
or U4329 (N_4329,N_3772,N_3685);
xor U4330 (N_4330,N_3878,N_3605);
or U4331 (N_4331,N_3677,N_3822);
nor U4332 (N_4332,N_3758,N_3725);
nand U4333 (N_4333,N_3634,N_3897);
xor U4334 (N_4334,N_3721,N_3920);
or U4335 (N_4335,N_3977,N_3733);
nand U4336 (N_4336,N_3716,N_3525);
or U4337 (N_4337,N_3587,N_3700);
nand U4338 (N_4338,N_3826,N_3783);
xnor U4339 (N_4339,N_3849,N_3804);
nor U4340 (N_4340,N_3575,N_3982);
nor U4341 (N_4341,N_3820,N_3737);
xnor U4342 (N_4342,N_3599,N_3595);
or U4343 (N_4343,N_3615,N_3905);
and U4344 (N_4344,N_3724,N_3579);
or U4345 (N_4345,N_3508,N_3842);
or U4346 (N_4346,N_3865,N_3863);
or U4347 (N_4347,N_3755,N_3558);
and U4348 (N_4348,N_3544,N_3683);
xor U4349 (N_4349,N_3754,N_3626);
nor U4350 (N_4350,N_3765,N_3581);
xnor U4351 (N_4351,N_3850,N_3623);
or U4352 (N_4352,N_3736,N_3692);
and U4353 (N_4353,N_3758,N_3505);
and U4354 (N_4354,N_3850,N_3833);
and U4355 (N_4355,N_3601,N_3936);
and U4356 (N_4356,N_3648,N_3665);
nand U4357 (N_4357,N_3505,N_3586);
and U4358 (N_4358,N_3792,N_3597);
or U4359 (N_4359,N_3649,N_3979);
nor U4360 (N_4360,N_3852,N_3648);
and U4361 (N_4361,N_3790,N_3717);
nor U4362 (N_4362,N_3826,N_3975);
nand U4363 (N_4363,N_3886,N_3560);
nand U4364 (N_4364,N_3967,N_3832);
and U4365 (N_4365,N_3718,N_3625);
nor U4366 (N_4366,N_3550,N_3947);
and U4367 (N_4367,N_3870,N_3901);
xor U4368 (N_4368,N_3779,N_3952);
nor U4369 (N_4369,N_3780,N_3728);
xnor U4370 (N_4370,N_3651,N_3878);
and U4371 (N_4371,N_3885,N_3884);
nand U4372 (N_4372,N_3846,N_3597);
nor U4373 (N_4373,N_3510,N_3772);
and U4374 (N_4374,N_3993,N_3928);
and U4375 (N_4375,N_3913,N_3865);
nand U4376 (N_4376,N_3774,N_3684);
nand U4377 (N_4377,N_3863,N_3908);
nand U4378 (N_4378,N_3724,N_3960);
nand U4379 (N_4379,N_3557,N_3968);
nand U4380 (N_4380,N_3635,N_3757);
nand U4381 (N_4381,N_3817,N_3841);
nand U4382 (N_4382,N_3919,N_3614);
and U4383 (N_4383,N_3856,N_3914);
nand U4384 (N_4384,N_3561,N_3931);
nand U4385 (N_4385,N_3563,N_3910);
nand U4386 (N_4386,N_3646,N_3603);
and U4387 (N_4387,N_3941,N_3838);
nor U4388 (N_4388,N_3893,N_3810);
nor U4389 (N_4389,N_3912,N_3582);
and U4390 (N_4390,N_3953,N_3602);
nor U4391 (N_4391,N_3959,N_3747);
and U4392 (N_4392,N_3916,N_3514);
or U4393 (N_4393,N_3740,N_3695);
or U4394 (N_4394,N_3632,N_3679);
xor U4395 (N_4395,N_3854,N_3865);
and U4396 (N_4396,N_3530,N_3983);
nand U4397 (N_4397,N_3762,N_3589);
nor U4398 (N_4398,N_3558,N_3719);
nor U4399 (N_4399,N_3519,N_3812);
or U4400 (N_4400,N_3837,N_3752);
and U4401 (N_4401,N_3675,N_3587);
nor U4402 (N_4402,N_3523,N_3500);
nor U4403 (N_4403,N_3656,N_3955);
or U4404 (N_4404,N_3632,N_3704);
or U4405 (N_4405,N_3654,N_3853);
nor U4406 (N_4406,N_3723,N_3571);
or U4407 (N_4407,N_3791,N_3649);
nor U4408 (N_4408,N_3962,N_3854);
nor U4409 (N_4409,N_3797,N_3582);
and U4410 (N_4410,N_3522,N_3546);
nor U4411 (N_4411,N_3573,N_3576);
xnor U4412 (N_4412,N_3858,N_3536);
and U4413 (N_4413,N_3761,N_3693);
nand U4414 (N_4414,N_3560,N_3748);
and U4415 (N_4415,N_3860,N_3674);
and U4416 (N_4416,N_3711,N_3959);
or U4417 (N_4417,N_3740,N_3646);
nand U4418 (N_4418,N_3608,N_3973);
nor U4419 (N_4419,N_3969,N_3613);
or U4420 (N_4420,N_3790,N_3927);
nor U4421 (N_4421,N_3648,N_3784);
xnor U4422 (N_4422,N_3751,N_3515);
and U4423 (N_4423,N_3680,N_3654);
nand U4424 (N_4424,N_3643,N_3591);
or U4425 (N_4425,N_3685,N_3782);
nor U4426 (N_4426,N_3782,N_3939);
and U4427 (N_4427,N_3904,N_3524);
or U4428 (N_4428,N_3604,N_3608);
nor U4429 (N_4429,N_3613,N_3743);
nand U4430 (N_4430,N_3647,N_3689);
nand U4431 (N_4431,N_3857,N_3685);
nor U4432 (N_4432,N_3950,N_3981);
nand U4433 (N_4433,N_3777,N_3725);
or U4434 (N_4434,N_3676,N_3728);
nand U4435 (N_4435,N_3944,N_3594);
and U4436 (N_4436,N_3820,N_3569);
nor U4437 (N_4437,N_3678,N_3867);
nand U4438 (N_4438,N_3852,N_3608);
and U4439 (N_4439,N_3928,N_3834);
nand U4440 (N_4440,N_3918,N_3976);
or U4441 (N_4441,N_3692,N_3720);
and U4442 (N_4442,N_3533,N_3748);
and U4443 (N_4443,N_3657,N_3875);
and U4444 (N_4444,N_3863,N_3972);
and U4445 (N_4445,N_3841,N_3601);
nor U4446 (N_4446,N_3795,N_3516);
nand U4447 (N_4447,N_3701,N_3960);
and U4448 (N_4448,N_3793,N_3664);
xnor U4449 (N_4449,N_3590,N_3923);
nand U4450 (N_4450,N_3632,N_3665);
and U4451 (N_4451,N_3974,N_3657);
nor U4452 (N_4452,N_3768,N_3626);
and U4453 (N_4453,N_3702,N_3767);
or U4454 (N_4454,N_3763,N_3827);
nand U4455 (N_4455,N_3859,N_3819);
xor U4456 (N_4456,N_3686,N_3775);
xnor U4457 (N_4457,N_3668,N_3964);
or U4458 (N_4458,N_3646,N_3606);
nand U4459 (N_4459,N_3651,N_3985);
and U4460 (N_4460,N_3561,N_3926);
or U4461 (N_4461,N_3742,N_3752);
or U4462 (N_4462,N_3848,N_3901);
and U4463 (N_4463,N_3948,N_3640);
nand U4464 (N_4464,N_3688,N_3723);
nor U4465 (N_4465,N_3869,N_3632);
nor U4466 (N_4466,N_3816,N_3583);
and U4467 (N_4467,N_3723,N_3928);
nand U4468 (N_4468,N_3641,N_3857);
xnor U4469 (N_4469,N_3539,N_3682);
xor U4470 (N_4470,N_3880,N_3828);
or U4471 (N_4471,N_3719,N_3697);
nor U4472 (N_4472,N_3569,N_3747);
xor U4473 (N_4473,N_3538,N_3895);
nand U4474 (N_4474,N_3706,N_3715);
xor U4475 (N_4475,N_3885,N_3794);
or U4476 (N_4476,N_3766,N_3866);
and U4477 (N_4477,N_3512,N_3862);
and U4478 (N_4478,N_3717,N_3825);
xor U4479 (N_4479,N_3925,N_3811);
or U4480 (N_4480,N_3921,N_3828);
and U4481 (N_4481,N_3818,N_3848);
or U4482 (N_4482,N_3656,N_3711);
and U4483 (N_4483,N_3780,N_3743);
nand U4484 (N_4484,N_3860,N_3534);
nor U4485 (N_4485,N_3899,N_3803);
or U4486 (N_4486,N_3630,N_3703);
nand U4487 (N_4487,N_3811,N_3530);
or U4488 (N_4488,N_3547,N_3607);
nand U4489 (N_4489,N_3547,N_3779);
nor U4490 (N_4490,N_3976,N_3742);
and U4491 (N_4491,N_3868,N_3595);
nor U4492 (N_4492,N_3745,N_3922);
or U4493 (N_4493,N_3863,N_3617);
or U4494 (N_4494,N_3814,N_3925);
nand U4495 (N_4495,N_3567,N_3657);
and U4496 (N_4496,N_3544,N_3588);
and U4497 (N_4497,N_3995,N_3900);
and U4498 (N_4498,N_3612,N_3952);
and U4499 (N_4499,N_3940,N_3820);
and U4500 (N_4500,N_4089,N_4426);
nand U4501 (N_4501,N_4220,N_4321);
nand U4502 (N_4502,N_4392,N_4249);
or U4503 (N_4503,N_4276,N_4326);
xor U4504 (N_4504,N_4064,N_4479);
and U4505 (N_4505,N_4011,N_4128);
and U4506 (N_4506,N_4232,N_4308);
xor U4507 (N_4507,N_4238,N_4202);
and U4508 (N_4508,N_4384,N_4218);
and U4509 (N_4509,N_4059,N_4250);
nand U4510 (N_4510,N_4325,N_4465);
xor U4511 (N_4511,N_4228,N_4283);
or U4512 (N_4512,N_4241,N_4034);
or U4513 (N_4513,N_4138,N_4285);
nor U4514 (N_4514,N_4083,N_4313);
nor U4515 (N_4515,N_4445,N_4247);
xnor U4516 (N_4516,N_4466,N_4018);
nor U4517 (N_4517,N_4448,N_4193);
nor U4518 (N_4518,N_4364,N_4158);
nand U4519 (N_4519,N_4009,N_4294);
nor U4520 (N_4520,N_4168,N_4171);
and U4521 (N_4521,N_4380,N_4396);
and U4522 (N_4522,N_4177,N_4292);
or U4523 (N_4523,N_4328,N_4097);
or U4524 (N_4524,N_4441,N_4290);
or U4525 (N_4525,N_4414,N_4116);
nor U4526 (N_4526,N_4015,N_4181);
and U4527 (N_4527,N_4067,N_4062);
or U4528 (N_4528,N_4470,N_4301);
and U4529 (N_4529,N_4192,N_4302);
nand U4530 (N_4530,N_4147,N_4230);
nand U4531 (N_4531,N_4222,N_4201);
nor U4532 (N_4532,N_4262,N_4494);
and U4533 (N_4533,N_4022,N_4439);
or U4534 (N_4534,N_4284,N_4005);
nand U4535 (N_4535,N_4454,N_4440);
or U4536 (N_4536,N_4031,N_4182);
nand U4537 (N_4537,N_4281,N_4280);
and U4538 (N_4538,N_4274,N_4122);
nor U4539 (N_4539,N_4449,N_4299);
and U4540 (N_4540,N_4170,N_4038);
nand U4541 (N_4541,N_4113,N_4189);
or U4542 (N_4542,N_4112,N_4119);
or U4543 (N_4543,N_4322,N_4333);
nand U4544 (N_4544,N_4106,N_4300);
and U4545 (N_4545,N_4279,N_4307);
nor U4546 (N_4546,N_4371,N_4408);
nor U4547 (N_4547,N_4187,N_4446);
xnor U4548 (N_4548,N_4125,N_4073);
nand U4549 (N_4549,N_4331,N_4190);
nor U4550 (N_4550,N_4431,N_4288);
nor U4551 (N_4551,N_4224,N_4462);
and U4552 (N_4552,N_4374,N_4376);
xnor U4553 (N_4553,N_4099,N_4235);
and U4554 (N_4554,N_4207,N_4378);
xnor U4555 (N_4555,N_4443,N_4151);
nand U4556 (N_4556,N_4404,N_4039);
nand U4557 (N_4557,N_4107,N_4499);
nor U4558 (N_4558,N_4155,N_4037);
or U4559 (N_4559,N_4358,N_4256);
nor U4560 (N_4560,N_4475,N_4251);
nand U4561 (N_4561,N_4141,N_4156);
nor U4562 (N_4562,N_4263,N_4267);
and U4563 (N_4563,N_4338,N_4336);
nand U4564 (N_4564,N_4355,N_4381);
and U4565 (N_4565,N_4058,N_4487);
nand U4566 (N_4566,N_4061,N_4101);
nand U4567 (N_4567,N_4486,N_4117);
xnor U4568 (N_4568,N_4016,N_4471);
xor U4569 (N_4569,N_4407,N_4135);
nor U4570 (N_4570,N_4260,N_4076);
or U4571 (N_4571,N_4273,N_4161);
and U4572 (N_4572,N_4140,N_4103);
and U4573 (N_4573,N_4143,N_4272);
and U4574 (N_4574,N_4060,N_4052);
nor U4575 (N_4575,N_4390,N_4409);
xor U4576 (N_4576,N_4210,N_4341);
nand U4577 (N_4577,N_4229,N_4007);
and U4578 (N_4578,N_4367,N_4463);
nor U4579 (N_4579,N_4054,N_4360);
nand U4580 (N_4580,N_4199,N_4315);
and U4581 (N_4581,N_4419,N_4402);
xor U4582 (N_4582,N_4478,N_4043);
and U4583 (N_4583,N_4417,N_4354);
or U4584 (N_4584,N_4468,N_4040);
or U4585 (N_4585,N_4342,N_4123);
and U4586 (N_4586,N_4204,N_4436);
xor U4587 (N_4587,N_4361,N_4314);
nand U4588 (N_4588,N_4447,N_4346);
nand U4589 (N_4589,N_4359,N_4074);
and U4590 (N_4590,N_4191,N_4254);
and U4591 (N_4591,N_4093,N_4421);
nor U4592 (N_4592,N_4226,N_4277);
and U4593 (N_4593,N_4065,N_4266);
nor U4594 (N_4594,N_4066,N_4169);
xnor U4595 (N_4595,N_4146,N_4027);
nand U4596 (N_4596,N_4438,N_4053);
or U4597 (N_4597,N_4287,N_4227);
or U4598 (N_4598,N_4176,N_4002);
and U4599 (N_4599,N_4236,N_4096);
or U4600 (N_4600,N_4063,N_4023);
and U4601 (N_4601,N_4351,N_4049);
nand U4602 (N_4602,N_4424,N_4377);
or U4603 (N_4603,N_4091,N_4282);
or U4604 (N_4604,N_4382,N_4186);
nor U4605 (N_4605,N_4363,N_4042);
xnor U4606 (N_4606,N_4148,N_4026);
or U4607 (N_4607,N_4188,N_4370);
and U4608 (N_4608,N_4434,N_4435);
or U4609 (N_4609,N_4464,N_4339);
or U4610 (N_4610,N_4388,N_4221);
and U4611 (N_4611,N_4303,N_4057);
xnor U4612 (N_4612,N_4418,N_4327);
nand U4613 (N_4613,N_4369,N_4410);
nand U4614 (N_4614,N_4102,N_4337);
nor U4615 (N_4615,N_4304,N_4179);
or U4616 (N_4616,N_4350,N_4139);
xor U4617 (N_4617,N_4244,N_4312);
nor U4618 (N_4618,N_4457,N_4114);
or U4619 (N_4619,N_4041,N_4162);
nor U4620 (N_4620,N_4269,N_4003);
nor U4621 (N_4621,N_4134,N_4398);
nand U4622 (N_4622,N_4021,N_4180);
and U4623 (N_4623,N_4278,N_4142);
and U4624 (N_4624,N_4121,N_4437);
xor U4625 (N_4625,N_4233,N_4197);
nor U4626 (N_4626,N_4387,N_4298);
or U4627 (N_4627,N_4335,N_4217);
or U4628 (N_4628,N_4271,N_4024);
xor U4629 (N_4629,N_4131,N_4391);
and U4630 (N_4630,N_4077,N_4356);
nor U4631 (N_4631,N_4020,N_4483);
nand U4632 (N_4632,N_4324,N_4045);
and U4633 (N_4633,N_4496,N_4344);
nor U4634 (N_4634,N_4401,N_4240);
nor U4635 (N_4635,N_4100,N_4033);
and U4636 (N_4636,N_4212,N_4195);
or U4637 (N_4637,N_4000,N_4019);
and U4638 (N_4638,N_4050,N_4451);
and U4639 (N_4639,N_4366,N_4084);
and U4640 (N_4640,N_4268,N_4025);
or U4641 (N_4641,N_4044,N_4166);
nand U4642 (N_4642,N_4194,N_4072);
nand U4643 (N_4643,N_4329,N_4476);
nand U4644 (N_4644,N_4094,N_4126);
and U4645 (N_4645,N_4425,N_4118);
nor U4646 (N_4646,N_4458,N_4352);
nand U4647 (N_4647,N_4444,N_4498);
nand U4648 (N_4648,N_4085,N_4320);
nand U4649 (N_4649,N_4423,N_4348);
and U4650 (N_4650,N_4129,N_4428);
nor U4651 (N_4651,N_4453,N_4413);
nand U4652 (N_4652,N_4490,N_4252);
nand U4653 (N_4653,N_4332,N_4270);
xnor U4654 (N_4654,N_4185,N_4157);
nor U4655 (N_4655,N_4017,N_4014);
xor U4656 (N_4656,N_4255,N_4460);
nor U4657 (N_4657,N_4372,N_4133);
and U4658 (N_4658,N_4048,N_4368);
nor U4659 (N_4659,N_4461,N_4450);
and U4660 (N_4660,N_4253,N_4137);
nand U4661 (N_4661,N_4154,N_4485);
and U4662 (N_4662,N_4264,N_4205);
nand U4663 (N_4663,N_4245,N_4365);
and U4664 (N_4664,N_4160,N_4412);
and U4665 (N_4665,N_4415,N_4297);
nand U4666 (N_4666,N_4257,N_4400);
nand U4667 (N_4667,N_4343,N_4200);
nor U4668 (N_4668,N_4152,N_4130);
nor U4669 (N_4669,N_4068,N_4008);
or U4670 (N_4670,N_4203,N_4079);
and U4671 (N_4671,N_4196,N_4234);
nor U4672 (N_4672,N_4237,N_4353);
xor U4673 (N_4673,N_4075,N_4318);
xnor U4674 (N_4674,N_4108,N_4088);
nor U4675 (N_4675,N_4144,N_4167);
or U4676 (N_4676,N_4150,N_4459);
or U4677 (N_4677,N_4178,N_4422);
nor U4678 (N_4678,N_4149,N_4484);
xor U4679 (N_4679,N_4416,N_4373);
nor U4680 (N_4680,N_4296,N_4482);
and U4681 (N_4681,N_4124,N_4051);
nor U4682 (N_4682,N_4006,N_4491);
nand U4683 (N_4683,N_4399,N_4206);
and U4684 (N_4684,N_4397,N_4375);
or U4685 (N_4685,N_4334,N_4243);
or U4686 (N_4686,N_4291,N_4165);
or U4687 (N_4687,N_4488,N_4163);
xnor U4688 (N_4688,N_4455,N_4078);
or U4689 (N_4689,N_4469,N_4120);
or U4690 (N_4690,N_4242,N_4001);
nor U4691 (N_4691,N_4136,N_4497);
xnor U4692 (N_4692,N_4183,N_4319);
nor U4693 (N_4693,N_4411,N_4208);
and U4694 (N_4694,N_4216,N_4098);
nor U4695 (N_4695,N_4092,N_4474);
and U4696 (N_4696,N_4082,N_4010);
and U4697 (N_4697,N_4070,N_4013);
or U4698 (N_4698,N_4071,N_4473);
or U4699 (N_4699,N_4105,N_4115);
or U4700 (N_4700,N_4214,N_4164);
nand U4701 (N_4701,N_4132,N_4261);
or U4702 (N_4702,N_4225,N_4111);
nand U4703 (N_4703,N_4184,N_4442);
nand U4704 (N_4704,N_4047,N_4393);
nor U4705 (N_4705,N_4090,N_4386);
nand U4706 (N_4706,N_4258,N_4055);
nand U4707 (N_4707,N_4309,N_4036);
xor U4708 (N_4708,N_4323,N_4427);
and U4709 (N_4709,N_4175,N_4056);
or U4710 (N_4710,N_4403,N_4104);
nand U4711 (N_4711,N_4383,N_4467);
or U4712 (N_4712,N_4480,N_4306);
nor U4713 (N_4713,N_4275,N_4347);
nor U4714 (N_4714,N_4456,N_4223);
and U4715 (N_4715,N_4035,N_4211);
or U4716 (N_4716,N_4265,N_4305);
nand U4717 (N_4717,N_4430,N_4493);
and U4718 (N_4718,N_4420,N_4429);
or U4719 (N_4719,N_4215,N_4012);
nor U4720 (N_4720,N_4030,N_4289);
nand U4721 (N_4721,N_4330,N_4213);
or U4722 (N_4722,N_4173,N_4174);
nand U4723 (N_4723,N_4310,N_4248);
nor U4724 (N_4724,N_4357,N_4159);
nand U4725 (N_4725,N_4127,N_4246);
nand U4726 (N_4726,N_4345,N_4069);
and U4727 (N_4727,N_4406,N_4395);
nor U4728 (N_4728,N_4153,N_4145);
or U4729 (N_4729,N_4209,N_4295);
nor U4730 (N_4730,N_4086,N_4080);
nand U4731 (N_4731,N_4492,N_4286);
or U4732 (N_4732,N_4004,N_4477);
xor U4733 (N_4733,N_4379,N_4046);
or U4734 (N_4734,N_4489,N_4032);
nor U4735 (N_4735,N_4259,N_4087);
or U4736 (N_4736,N_4389,N_4028);
or U4737 (N_4737,N_4495,N_4172);
nor U4738 (N_4738,N_4349,N_4311);
or U4739 (N_4739,N_4198,N_4095);
or U4740 (N_4740,N_4029,N_4394);
or U4741 (N_4741,N_4452,N_4109);
and U4742 (N_4742,N_4316,N_4081);
nor U4743 (N_4743,N_4219,N_4432);
and U4744 (N_4744,N_4405,N_4385);
xor U4745 (N_4745,N_4293,N_4239);
nand U4746 (N_4746,N_4472,N_4481);
nor U4747 (N_4747,N_4433,N_4231);
nor U4748 (N_4748,N_4362,N_4110);
or U4749 (N_4749,N_4340,N_4317);
and U4750 (N_4750,N_4267,N_4179);
or U4751 (N_4751,N_4251,N_4030);
and U4752 (N_4752,N_4119,N_4433);
and U4753 (N_4753,N_4127,N_4289);
and U4754 (N_4754,N_4070,N_4220);
or U4755 (N_4755,N_4143,N_4325);
and U4756 (N_4756,N_4136,N_4426);
or U4757 (N_4757,N_4222,N_4303);
xnor U4758 (N_4758,N_4120,N_4299);
xor U4759 (N_4759,N_4295,N_4181);
nand U4760 (N_4760,N_4270,N_4311);
and U4761 (N_4761,N_4429,N_4417);
and U4762 (N_4762,N_4107,N_4079);
or U4763 (N_4763,N_4314,N_4319);
and U4764 (N_4764,N_4160,N_4396);
and U4765 (N_4765,N_4176,N_4360);
xor U4766 (N_4766,N_4392,N_4451);
nand U4767 (N_4767,N_4157,N_4384);
or U4768 (N_4768,N_4237,N_4255);
nor U4769 (N_4769,N_4391,N_4004);
and U4770 (N_4770,N_4446,N_4111);
nand U4771 (N_4771,N_4335,N_4254);
nor U4772 (N_4772,N_4423,N_4409);
or U4773 (N_4773,N_4476,N_4308);
nor U4774 (N_4774,N_4332,N_4427);
nand U4775 (N_4775,N_4499,N_4471);
nand U4776 (N_4776,N_4193,N_4476);
nand U4777 (N_4777,N_4190,N_4333);
or U4778 (N_4778,N_4096,N_4468);
xor U4779 (N_4779,N_4281,N_4415);
nand U4780 (N_4780,N_4212,N_4364);
or U4781 (N_4781,N_4114,N_4295);
nand U4782 (N_4782,N_4299,N_4321);
and U4783 (N_4783,N_4303,N_4017);
nor U4784 (N_4784,N_4476,N_4246);
or U4785 (N_4785,N_4264,N_4079);
and U4786 (N_4786,N_4446,N_4295);
and U4787 (N_4787,N_4186,N_4315);
or U4788 (N_4788,N_4006,N_4024);
nand U4789 (N_4789,N_4414,N_4239);
nor U4790 (N_4790,N_4254,N_4376);
nor U4791 (N_4791,N_4095,N_4125);
nor U4792 (N_4792,N_4214,N_4107);
and U4793 (N_4793,N_4414,N_4332);
and U4794 (N_4794,N_4118,N_4435);
or U4795 (N_4795,N_4066,N_4044);
and U4796 (N_4796,N_4064,N_4155);
and U4797 (N_4797,N_4153,N_4220);
nand U4798 (N_4798,N_4318,N_4214);
and U4799 (N_4799,N_4465,N_4210);
or U4800 (N_4800,N_4333,N_4213);
or U4801 (N_4801,N_4300,N_4263);
xnor U4802 (N_4802,N_4415,N_4144);
and U4803 (N_4803,N_4228,N_4077);
nor U4804 (N_4804,N_4257,N_4181);
nor U4805 (N_4805,N_4120,N_4040);
and U4806 (N_4806,N_4029,N_4184);
or U4807 (N_4807,N_4039,N_4319);
nand U4808 (N_4808,N_4266,N_4176);
nand U4809 (N_4809,N_4273,N_4379);
and U4810 (N_4810,N_4491,N_4208);
nor U4811 (N_4811,N_4301,N_4288);
nor U4812 (N_4812,N_4381,N_4334);
nor U4813 (N_4813,N_4269,N_4324);
xnor U4814 (N_4814,N_4166,N_4229);
nand U4815 (N_4815,N_4301,N_4225);
nor U4816 (N_4816,N_4388,N_4096);
nor U4817 (N_4817,N_4275,N_4089);
nor U4818 (N_4818,N_4278,N_4086);
nor U4819 (N_4819,N_4193,N_4018);
or U4820 (N_4820,N_4092,N_4345);
xor U4821 (N_4821,N_4176,N_4472);
nand U4822 (N_4822,N_4057,N_4420);
xnor U4823 (N_4823,N_4236,N_4295);
or U4824 (N_4824,N_4467,N_4099);
and U4825 (N_4825,N_4354,N_4088);
nand U4826 (N_4826,N_4259,N_4461);
or U4827 (N_4827,N_4195,N_4257);
or U4828 (N_4828,N_4456,N_4412);
nor U4829 (N_4829,N_4341,N_4398);
nand U4830 (N_4830,N_4053,N_4231);
and U4831 (N_4831,N_4469,N_4305);
nand U4832 (N_4832,N_4307,N_4191);
xnor U4833 (N_4833,N_4163,N_4150);
nand U4834 (N_4834,N_4207,N_4226);
or U4835 (N_4835,N_4467,N_4090);
or U4836 (N_4836,N_4161,N_4304);
or U4837 (N_4837,N_4358,N_4215);
nand U4838 (N_4838,N_4219,N_4287);
nor U4839 (N_4839,N_4193,N_4105);
or U4840 (N_4840,N_4172,N_4134);
nor U4841 (N_4841,N_4086,N_4304);
and U4842 (N_4842,N_4139,N_4225);
and U4843 (N_4843,N_4477,N_4300);
nand U4844 (N_4844,N_4159,N_4484);
nor U4845 (N_4845,N_4452,N_4448);
nand U4846 (N_4846,N_4389,N_4218);
nor U4847 (N_4847,N_4178,N_4327);
nand U4848 (N_4848,N_4324,N_4206);
and U4849 (N_4849,N_4380,N_4316);
nand U4850 (N_4850,N_4378,N_4350);
nor U4851 (N_4851,N_4468,N_4192);
or U4852 (N_4852,N_4109,N_4119);
and U4853 (N_4853,N_4416,N_4186);
nand U4854 (N_4854,N_4383,N_4299);
nand U4855 (N_4855,N_4322,N_4368);
nand U4856 (N_4856,N_4386,N_4406);
or U4857 (N_4857,N_4069,N_4374);
or U4858 (N_4858,N_4420,N_4264);
or U4859 (N_4859,N_4128,N_4335);
or U4860 (N_4860,N_4150,N_4157);
xor U4861 (N_4861,N_4161,N_4032);
nand U4862 (N_4862,N_4271,N_4219);
and U4863 (N_4863,N_4408,N_4279);
or U4864 (N_4864,N_4321,N_4219);
xnor U4865 (N_4865,N_4236,N_4228);
nor U4866 (N_4866,N_4314,N_4368);
xnor U4867 (N_4867,N_4332,N_4136);
nor U4868 (N_4868,N_4126,N_4092);
nand U4869 (N_4869,N_4040,N_4245);
xnor U4870 (N_4870,N_4227,N_4329);
or U4871 (N_4871,N_4024,N_4484);
nand U4872 (N_4872,N_4075,N_4289);
or U4873 (N_4873,N_4387,N_4447);
and U4874 (N_4874,N_4351,N_4121);
or U4875 (N_4875,N_4265,N_4276);
nor U4876 (N_4876,N_4460,N_4089);
nor U4877 (N_4877,N_4465,N_4149);
or U4878 (N_4878,N_4012,N_4430);
and U4879 (N_4879,N_4201,N_4033);
and U4880 (N_4880,N_4252,N_4423);
nor U4881 (N_4881,N_4139,N_4320);
or U4882 (N_4882,N_4240,N_4237);
and U4883 (N_4883,N_4405,N_4099);
nor U4884 (N_4884,N_4055,N_4244);
or U4885 (N_4885,N_4348,N_4404);
nor U4886 (N_4886,N_4192,N_4442);
and U4887 (N_4887,N_4292,N_4483);
nor U4888 (N_4888,N_4431,N_4387);
nor U4889 (N_4889,N_4293,N_4263);
xor U4890 (N_4890,N_4098,N_4450);
xor U4891 (N_4891,N_4361,N_4322);
nor U4892 (N_4892,N_4143,N_4383);
xnor U4893 (N_4893,N_4084,N_4469);
xnor U4894 (N_4894,N_4036,N_4123);
nor U4895 (N_4895,N_4266,N_4070);
or U4896 (N_4896,N_4102,N_4455);
and U4897 (N_4897,N_4345,N_4018);
nor U4898 (N_4898,N_4311,N_4470);
and U4899 (N_4899,N_4392,N_4282);
and U4900 (N_4900,N_4149,N_4180);
nor U4901 (N_4901,N_4227,N_4411);
nor U4902 (N_4902,N_4035,N_4015);
nand U4903 (N_4903,N_4439,N_4253);
and U4904 (N_4904,N_4270,N_4324);
or U4905 (N_4905,N_4114,N_4402);
nand U4906 (N_4906,N_4466,N_4122);
and U4907 (N_4907,N_4169,N_4492);
and U4908 (N_4908,N_4322,N_4031);
nand U4909 (N_4909,N_4346,N_4192);
nand U4910 (N_4910,N_4324,N_4103);
xor U4911 (N_4911,N_4092,N_4185);
and U4912 (N_4912,N_4483,N_4211);
nand U4913 (N_4913,N_4498,N_4176);
and U4914 (N_4914,N_4185,N_4413);
and U4915 (N_4915,N_4462,N_4036);
nand U4916 (N_4916,N_4485,N_4235);
nand U4917 (N_4917,N_4236,N_4453);
nor U4918 (N_4918,N_4206,N_4418);
nor U4919 (N_4919,N_4337,N_4421);
and U4920 (N_4920,N_4104,N_4034);
or U4921 (N_4921,N_4145,N_4474);
and U4922 (N_4922,N_4255,N_4225);
and U4923 (N_4923,N_4179,N_4414);
and U4924 (N_4924,N_4372,N_4127);
nor U4925 (N_4925,N_4032,N_4245);
and U4926 (N_4926,N_4005,N_4053);
or U4927 (N_4927,N_4415,N_4003);
nor U4928 (N_4928,N_4146,N_4386);
or U4929 (N_4929,N_4497,N_4093);
nor U4930 (N_4930,N_4037,N_4358);
nor U4931 (N_4931,N_4452,N_4354);
and U4932 (N_4932,N_4332,N_4093);
and U4933 (N_4933,N_4342,N_4250);
or U4934 (N_4934,N_4159,N_4247);
nand U4935 (N_4935,N_4042,N_4011);
or U4936 (N_4936,N_4096,N_4209);
and U4937 (N_4937,N_4339,N_4076);
or U4938 (N_4938,N_4273,N_4239);
nand U4939 (N_4939,N_4471,N_4278);
and U4940 (N_4940,N_4170,N_4207);
nor U4941 (N_4941,N_4213,N_4482);
and U4942 (N_4942,N_4250,N_4002);
nor U4943 (N_4943,N_4236,N_4280);
and U4944 (N_4944,N_4154,N_4133);
or U4945 (N_4945,N_4156,N_4001);
xnor U4946 (N_4946,N_4299,N_4180);
and U4947 (N_4947,N_4207,N_4470);
nand U4948 (N_4948,N_4395,N_4320);
and U4949 (N_4949,N_4210,N_4048);
nand U4950 (N_4950,N_4153,N_4421);
nand U4951 (N_4951,N_4201,N_4156);
nor U4952 (N_4952,N_4249,N_4304);
nand U4953 (N_4953,N_4249,N_4420);
nor U4954 (N_4954,N_4485,N_4293);
xnor U4955 (N_4955,N_4086,N_4287);
and U4956 (N_4956,N_4154,N_4025);
nand U4957 (N_4957,N_4101,N_4306);
nor U4958 (N_4958,N_4001,N_4478);
xor U4959 (N_4959,N_4479,N_4392);
or U4960 (N_4960,N_4241,N_4284);
xor U4961 (N_4961,N_4435,N_4241);
or U4962 (N_4962,N_4071,N_4111);
nor U4963 (N_4963,N_4409,N_4108);
nand U4964 (N_4964,N_4463,N_4272);
or U4965 (N_4965,N_4334,N_4464);
nor U4966 (N_4966,N_4262,N_4497);
xnor U4967 (N_4967,N_4168,N_4407);
or U4968 (N_4968,N_4103,N_4044);
and U4969 (N_4969,N_4303,N_4023);
or U4970 (N_4970,N_4076,N_4253);
and U4971 (N_4971,N_4036,N_4481);
nand U4972 (N_4972,N_4343,N_4264);
or U4973 (N_4973,N_4266,N_4303);
and U4974 (N_4974,N_4187,N_4130);
nor U4975 (N_4975,N_4202,N_4084);
and U4976 (N_4976,N_4152,N_4498);
nand U4977 (N_4977,N_4109,N_4397);
or U4978 (N_4978,N_4189,N_4464);
xnor U4979 (N_4979,N_4237,N_4460);
nor U4980 (N_4980,N_4204,N_4300);
xnor U4981 (N_4981,N_4309,N_4222);
xnor U4982 (N_4982,N_4083,N_4192);
or U4983 (N_4983,N_4115,N_4174);
or U4984 (N_4984,N_4348,N_4424);
nand U4985 (N_4985,N_4442,N_4063);
nor U4986 (N_4986,N_4370,N_4051);
xnor U4987 (N_4987,N_4426,N_4466);
or U4988 (N_4988,N_4059,N_4273);
nand U4989 (N_4989,N_4262,N_4245);
and U4990 (N_4990,N_4048,N_4359);
or U4991 (N_4991,N_4421,N_4165);
and U4992 (N_4992,N_4365,N_4190);
nand U4993 (N_4993,N_4458,N_4207);
nor U4994 (N_4994,N_4285,N_4223);
xor U4995 (N_4995,N_4107,N_4234);
nor U4996 (N_4996,N_4400,N_4322);
nor U4997 (N_4997,N_4028,N_4396);
nor U4998 (N_4998,N_4214,N_4007);
nor U4999 (N_4999,N_4301,N_4368);
nor UO_0 (O_0,N_4619,N_4900);
nor UO_1 (O_1,N_4665,N_4845);
nand UO_2 (O_2,N_4676,N_4592);
nor UO_3 (O_3,N_4680,N_4581);
or UO_4 (O_4,N_4746,N_4636);
nor UO_5 (O_5,N_4600,N_4921);
nor UO_6 (O_6,N_4591,N_4730);
or UO_7 (O_7,N_4578,N_4882);
or UO_8 (O_8,N_4951,N_4723);
nor UO_9 (O_9,N_4797,N_4962);
and UO_10 (O_10,N_4806,N_4749);
nand UO_11 (O_11,N_4594,N_4731);
nand UO_12 (O_12,N_4769,N_4656);
and UO_13 (O_13,N_4979,N_4599);
and UO_14 (O_14,N_4791,N_4673);
nor UO_15 (O_15,N_4865,N_4885);
or UO_16 (O_16,N_4847,N_4950);
nor UO_17 (O_17,N_4706,N_4641);
nand UO_18 (O_18,N_4884,N_4721);
and UO_19 (O_19,N_4707,N_4938);
nor UO_20 (O_20,N_4898,N_4501);
and UO_21 (O_21,N_4576,N_4633);
nand UO_22 (O_22,N_4798,N_4887);
and UO_23 (O_23,N_4651,N_4539);
nand UO_24 (O_24,N_4700,N_4844);
or UO_25 (O_25,N_4519,N_4699);
nor UO_26 (O_26,N_4760,N_4854);
nand UO_27 (O_27,N_4992,N_4792);
nor UO_28 (O_28,N_4763,N_4856);
and UO_29 (O_29,N_4892,N_4925);
xnor UO_30 (O_30,N_4508,N_4929);
nor UO_31 (O_31,N_4561,N_4981);
nor UO_32 (O_32,N_4575,N_4766);
or UO_33 (O_33,N_4704,N_4523);
nand UO_34 (O_34,N_4796,N_4531);
nand UO_35 (O_35,N_4756,N_4642);
and UO_36 (O_36,N_4615,N_4790);
or UO_37 (O_37,N_4907,N_4819);
nand UO_38 (O_38,N_4928,N_4776);
or UO_39 (O_39,N_4978,N_4540);
nor UO_40 (O_40,N_4744,N_4794);
or UO_41 (O_41,N_4852,N_4698);
and UO_42 (O_42,N_4529,N_4692);
and UO_43 (O_43,N_4520,N_4954);
or UO_44 (O_44,N_4653,N_4977);
nor UO_45 (O_45,N_4917,N_4754);
or UO_46 (O_46,N_4714,N_4574);
nand UO_47 (O_47,N_4638,N_4683);
and UO_48 (O_48,N_4565,N_4691);
nor UO_49 (O_49,N_4621,N_4681);
and UO_50 (O_50,N_4555,N_4660);
nand UO_51 (O_51,N_4982,N_4687);
or UO_52 (O_52,N_4940,N_4635);
nand UO_53 (O_53,N_4828,N_4500);
nor UO_54 (O_54,N_4858,N_4504);
nand UO_55 (O_55,N_4963,N_4972);
and UO_56 (O_56,N_4617,N_4886);
nor UO_57 (O_57,N_4780,N_4814);
or UO_58 (O_58,N_4643,N_4778);
and UO_59 (O_59,N_4842,N_4710);
nand UO_60 (O_60,N_4622,N_4559);
nand UO_61 (O_61,N_4703,N_4611);
or UO_62 (O_62,N_4804,N_4840);
and UO_63 (O_63,N_4663,N_4807);
nor UO_64 (O_64,N_4813,N_4782);
nor UO_65 (O_65,N_4659,N_4906);
and UO_66 (O_66,N_4616,N_4602);
nand UO_67 (O_67,N_4739,N_4815);
nand UO_68 (O_68,N_4625,N_4672);
and UO_69 (O_69,N_4866,N_4601);
and UO_70 (O_70,N_4878,N_4969);
nor UO_71 (O_71,N_4914,N_4585);
and UO_72 (O_72,N_4715,N_4697);
nand UO_73 (O_73,N_4548,N_4944);
nor UO_74 (O_74,N_4932,N_4553);
and UO_75 (O_75,N_4912,N_4996);
or UO_76 (O_76,N_4831,N_4855);
or UO_77 (O_77,N_4696,N_4899);
or UO_78 (O_78,N_4666,N_4607);
or UO_79 (O_79,N_4830,N_4544);
or UO_80 (O_80,N_4862,N_4597);
and UO_81 (O_81,N_4598,N_4727);
nand UO_82 (O_82,N_4631,N_4875);
xnor UO_83 (O_83,N_4571,N_4765);
or UO_84 (O_84,N_4521,N_4684);
or UO_85 (O_85,N_4927,N_4772);
or UO_86 (O_86,N_4793,N_4915);
or UO_87 (O_87,N_4573,N_4717);
or UO_88 (O_88,N_4580,N_4564);
and UO_89 (O_89,N_4848,N_4516);
nand UO_90 (O_90,N_4771,N_4670);
or UO_91 (O_91,N_4933,N_4708);
nand UO_92 (O_92,N_4527,N_4628);
nor UO_93 (O_93,N_4869,N_4720);
or UO_94 (O_94,N_4836,N_4911);
nor UO_95 (O_95,N_4664,N_4980);
xor UO_96 (O_96,N_4624,N_4901);
nand UO_97 (O_97,N_4952,N_4546);
or UO_98 (O_98,N_4510,N_4986);
and UO_99 (O_99,N_4736,N_4604);
nor UO_100 (O_100,N_4974,N_4550);
or UO_101 (O_101,N_4511,N_4957);
nand UO_102 (O_102,N_4705,N_4505);
and UO_103 (O_103,N_4733,N_4652);
and UO_104 (O_104,N_4823,N_4737);
nand UO_105 (O_105,N_4669,N_4909);
xor UO_106 (O_106,N_4997,N_4947);
xnor UO_107 (O_107,N_4724,N_4729);
nor UO_108 (O_108,N_4542,N_4945);
nor UO_109 (O_109,N_4515,N_4816);
nor UO_110 (O_110,N_4777,N_4820);
and UO_111 (O_111,N_4563,N_4964);
or UO_112 (O_112,N_4870,N_4570);
and UO_113 (O_113,N_4541,N_4606);
nor UO_114 (O_114,N_4758,N_4863);
and UO_115 (O_115,N_4655,N_4747);
nor UO_116 (O_116,N_4965,N_4554);
or UO_117 (O_117,N_4716,N_4904);
nor UO_118 (O_118,N_4608,N_4779);
or UO_119 (O_119,N_4567,N_4536);
or UO_120 (O_120,N_4586,N_4572);
xor UO_121 (O_121,N_4877,N_4627);
nand UO_122 (O_122,N_4818,N_4867);
nor UO_123 (O_123,N_4623,N_4789);
nand UO_124 (O_124,N_4924,N_4719);
nor UO_125 (O_125,N_4787,N_4662);
nor UO_126 (O_126,N_4868,N_4695);
xor UO_127 (O_127,N_4538,N_4506);
nor UO_128 (O_128,N_4752,N_4654);
nor UO_129 (O_129,N_4658,N_4639);
nor UO_130 (O_130,N_4690,N_4509);
or UO_131 (O_131,N_4674,N_4713);
nand UO_132 (O_132,N_4937,N_4552);
nor UO_133 (O_133,N_4799,N_4908);
nand UO_134 (O_134,N_4577,N_4883);
xor UO_135 (O_135,N_4893,N_4872);
and UO_136 (O_136,N_4750,N_4991);
and UO_137 (O_137,N_4603,N_4835);
or UO_138 (O_138,N_4851,N_4593);
and UO_139 (O_139,N_4566,N_4678);
nand UO_140 (O_140,N_4846,N_4989);
or UO_141 (O_141,N_4725,N_4918);
and UO_142 (O_142,N_4795,N_4745);
xnor UO_143 (O_143,N_4873,N_4988);
or UO_144 (O_144,N_4537,N_4612);
and UO_145 (O_145,N_4742,N_4800);
or UO_146 (O_146,N_4613,N_4524);
nor UO_147 (O_147,N_4919,N_4949);
or UO_148 (O_148,N_4941,N_4589);
or UO_149 (O_149,N_4595,N_4701);
and UO_150 (O_150,N_4502,N_4528);
nand UO_151 (O_151,N_4668,N_4817);
or UO_152 (O_152,N_4518,N_4618);
or UO_153 (O_153,N_4960,N_4811);
nor UO_154 (O_154,N_4667,N_4740);
xnor UO_155 (O_155,N_4838,N_4913);
nor UO_156 (O_156,N_4936,N_4786);
xor UO_157 (O_157,N_4530,N_4990);
nor UO_158 (O_158,N_4590,N_4547);
nor UO_159 (O_159,N_4810,N_4897);
and UO_160 (O_160,N_4543,N_4788);
and UO_161 (O_161,N_4558,N_4751);
and UO_162 (O_162,N_4525,N_4757);
nand UO_163 (O_163,N_4822,N_4946);
and UO_164 (O_164,N_4916,N_4959);
or UO_165 (O_165,N_4920,N_4970);
and UO_166 (O_166,N_4998,N_4976);
or UO_167 (O_167,N_4930,N_4943);
or UO_168 (O_168,N_4896,N_4614);
nand UO_169 (O_169,N_4588,N_4995);
nor UO_170 (O_170,N_4839,N_4753);
nand UO_171 (O_171,N_4584,N_4532);
nand UO_172 (O_172,N_4514,N_4709);
nor UO_173 (O_173,N_4999,N_4881);
nand UO_174 (O_174,N_4735,N_4985);
or UO_175 (O_175,N_4626,N_4809);
and UO_176 (O_176,N_4910,N_4994);
and UO_177 (O_177,N_4903,N_4876);
or UO_178 (O_178,N_4637,N_4812);
nor UO_179 (O_179,N_4583,N_4738);
nand UO_180 (O_180,N_4645,N_4890);
nor UO_181 (O_181,N_4843,N_4826);
and UO_182 (O_182,N_4644,N_4993);
xor UO_183 (O_183,N_4609,N_4634);
or UO_184 (O_184,N_4694,N_4834);
nor UO_185 (O_185,N_4685,N_4650);
and UO_186 (O_186,N_4891,N_4871);
or UO_187 (O_187,N_4512,N_4551);
or UO_188 (O_188,N_4773,N_4905);
xor UO_189 (O_189,N_4850,N_4712);
or UO_190 (O_190,N_4961,N_4732);
or UO_191 (O_191,N_4775,N_4702);
or UO_192 (O_192,N_4889,N_4770);
and UO_193 (O_193,N_4827,N_4726);
nand UO_194 (O_194,N_4649,N_4734);
nor UO_195 (O_195,N_4675,N_4569);
nor UO_196 (O_196,N_4967,N_4805);
and UO_197 (O_197,N_4534,N_4934);
and UO_198 (O_198,N_4507,N_4973);
nand UO_199 (O_199,N_4728,N_4833);
and UO_200 (O_200,N_4722,N_4802);
or UO_201 (O_201,N_4966,N_4864);
nor UO_202 (O_202,N_4661,N_4513);
xor UO_203 (O_203,N_4861,N_4688);
nand UO_204 (O_204,N_4557,N_4517);
nor UO_205 (O_205,N_4568,N_4596);
or UO_206 (O_206,N_4939,N_4556);
or UO_207 (O_207,N_4849,N_4647);
nor UO_208 (O_208,N_4748,N_4879);
and UO_209 (O_209,N_4888,N_4689);
nor UO_210 (O_210,N_4503,N_4931);
or UO_211 (O_211,N_4774,N_4923);
and UO_212 (O_212,N_4821,N_4987);
nor UO_213 (O_213,N_4686,N_4526);
nand UO_214 (O_214,N_4579,N_4743);
nor UO_215 (O_215,N_4693,N_4837);
and UO_216 (O_216,N_4860,N_4935);
xor UO_217 (O_217,N_4630,N_4582);
and UO_218 (O_218,N_4880,N_4562);
nand UO_219 (O_219,N_4956,N_4620);
or UO_220 (O_220,N_4968,N_4741);
or UO_221 (O_221,N_4767,N_4829);
nand UO_222 (O_222,N_4768,N_4825);
and UO_223 (O_223,N_4975,N_4533);
nand UO_224 (O_224,N_4857,N_4955);
nand UO_225 (O_225,N_4958,N_4711);
nand UO_226 (O_226,N_4942,N_4560);
nand UO_227 (O_227,N_4922,N_4648);
and UO_228 (O_228,N_4832,N_4953);
or UO_229 (O_229,N_4984,N_4785);
nor UO_230 (O_230,N_4948,N_4610);
or UO_231 (O_231,N_4646,N_4761);
and UO_232 (O_232,N_4640,N_4679);
and UO_233 (O_233,N_4759,N_4605);
nor UO_234 (O_234,N_4632,N_4971);
or UO_235 (O_235,N_4801,N_4549);
or UO_236 (O_236,N_4657,N_4803);
xor UO_237 (O_237,N_4522,N_4824);
and UO_238 (O_238,N_4894,N_4545);
nor UO_239 (O_239,N_4535,N_4853);
nor UO_240 (O_240,N_4718,N_4629);
nor UO_241 (O_241,N_4587,N_4682);
nand UO_242 (O_242,N_4755,N_4762);
or UO_243 (O_243,N_4671,N_4859);
and UO_244 (O_244,N_4902,N_4841);
xnor UO_245 (O_245,N_4983,N_4874);
xor UO_246 (O_246,N_4895,N_4808);
xor UO_247 (O_247,N_4781,N_4764);
nand UO_248 (O_248,N_4784,N_4926);
or UO_249 (O_249,N_4783,N_4677);
nor UO_250 (O_250,N_4889,N_4861);
nand UO_251 (O_251,N_4615,N_4957);
nand UO_252 (O_252,N_4925,N_4861);
and UO_253 (O_253,N_4913,N_4784);
and UO_254 (O_254,N_4812,N_4852);
or UO_255 (O_255,N_4788,N_4887);
and UO_256 (O_256,N_4679,N_4977);
or UO_257 (O_257,N_4685,N_4569);
nand UO_258 (O_258,N_4908,N_4724);
and UO_259 (O_259,N_4939,N_4819);
or UO_260 (O_260,N_4641,N_4988);
and UO_261 (O_261,N_4560,N_4529);
nand UO_262 (O_262,N_4731,N_4818);
or UO_263 (O_263,N_4709,N_4944);
or UO_264 (O_264,N_4856,N_4787);
or UO_265 (O_265,N_4501,N_4814);
and UO_266 (O_266,N_4874,N_4596);
xnor UO_267 (O_267,N_4776,N_4828);
nand UO_268 (O_268,N_4604,N_4893);
and UO_269 (O_269,N_4841,N_4822);
nand UO_270 (O_270,N_4574,N_4848);
nand UO_271 (O_271,N_4937,N_4839);
and UO_272 (O_272,N_4557,N_4621);
nand UO_273 (O_273,N_4558,N_4570);
or UO_274 (O_274,N_4625,N_4633);
nor UO_275 (O_275,N_4868,N_4638);
or UO_276 (O_276,N_4582,N_4881);
nand UO_277 (O_277,N_4709,N_4549);
xor UO_278 (O_278,N_4707,N_4592);
and UO_279 (O_279,N_4885,N_4908);
nand UO_280 (O_280,N_4929,N_4739);
nand UO_281 (O_281,N_4691,N_4562);
nand UO_282 (O_282,N_4658,N_4986);
nor UO_283 (O_283,N_4932,N_4984);
and UO_284 (O_284,N_4596,N_4527);
nor UO_285 (O_285,N_4817,N_4725);
or UO_286 (O_286,N_4524,N_4930);
and UO_287 (O_287,N_4773,N_4749);
nand UO_288 (O_288,N_4973,N_4716);
or UO_289 (O_289,N_4970,N_4561);
nand UO_290 (O_290,N_4581,N_4511);
and UO_291 (O_291,N_4812,N_4644);
or UO_292 (O_292,N_4704,N_4950);
nor UO_293 (O_293,N_4772,N_4888);
or UO_294 (O_294,N_4971,N_4761);
xor UO_295 (O_295,N_4931,N_4783);
nor UO_296 (O_296,N_4582,N_4664);
nand UO_297 (O_297,N_4671,N_4640);
xnor UO_298 (O_298,N_4778,N_4731);
nand UO_299 (O_299,N_4716,N_4886);
and UO_300 (O_300,N_4706,N_4574);
and UO_301 (O_301,N_4942,N_4591);
and UO_302 (O_302,N_4886,N_4984);
nor UO_303 (O_303,N_4980,N_4811);
or UO_304 (O_304,N_4921,N_4526);
nand UO_305 (O_305,N_4564,N_4546);
and UO_306 (O_306,N_4967,N_4667);
nand UO_307 (O_307,N_4967,N_4670);
nand UO_308 (O_308,N_4883,N_4522);
or UO_309 (O_309,N_4555,N_4713);
nor UO_310 (O_310,N_4585,N_4837);
nor UO_311 (O_311,N_4949,N_4603);
nand UO_312 (O_312,N_4564,N_4555);
or UO_313 (O_313,N_4787,N_4544);
or UO_314 (O_314,N_4652,N_4628);
or UO_315 (O_315,N_4769,N_4817);
nor UO_316 (O_316,N_4555,N_4687);
nand UO_317 (O_317,N_4601,N_4850);
xnor UO_318 (O_318,N_4878,N_4569);
and UO_319 (O_319,N_4773,N_4676);
nand UO_320 (O_320,N_4854,N_4637);
nor UO_321 (O_321,N_4766,N_4765);
and UO_322 (O_322,N_4652,N_4952);
nand UO_323 (O_323,N_4799,N_4683);
nor UO_324 (O_324,N_4734,N_4780);
xor UO_325 (O_325,N_4594,N_4672);
nand UO_326 (O_326,N_4683,N_4898);
nand UO_327 (O_327,N_4703,N_4518);
and UO_328 (O_328,N_4677,N_4503);
or UO_329 (O_329,N_4571,N_4695);
nor UO_330 (O_330,N_4991,N_4504);
or UO_331 (O_331,N_4828,N_4873);
xor UO_332 (O_332,N_4979,N_4834);
or UO_333 (O_333,N_4653,N_4914);
or UO_334 (O_334,N_4976,N_4728);
or UO_335 (O_335,N_4756,N_4725);
or UO_336 (O_336,N_4706,N_4803);
nor UO_337 (O_337,N_4598,N_4823);
or UO_338 (O_338,N_4919,N_4728);
nand UO_339 (O_339,N_4780,N_4507);
nand UO_340 (O_340,N_4987,N_4783);
xnor UO_341 (O_341,N_4659,N_4838);
nor UO_342 (O_342,N_4906,N_4530);
and UO_343 (O_343,N_4559,N_4506);
xor UO_344 (O_344,N_4772,N_4806);
xor UO_345 (O_345,N_4562,N_4906);
or UO_346 (O_346,N_4892,N_4852);
nand UO_347 (O_347,N_4610,N_4667);
and UO_348 (O_348,N_4689,N_4980);
nand UO_349 (O_349,N_4727,N_4751);
nor UO_350 (O_350,N_4751,N_4965);
or UO_351 (O_351,N_4687,N_4822);
and UO_352 (O_352,N_4732,N_4956);
xnor UO_353 (O_353,N_4777,N_4730);
xnor UO_354 (O_354,N_4754,N_4872);
and UO_355 (O_355,N_4991,N_4744);
and UO_356 (O_356,N_4549,N_4725);
xnor UO_357 (O_357,N_4911,N_4549);
and UO_358 (O_358,N_4577,N_4876);
and UO_359 (O_359,N_4510,N_4872);
nor UO_360 (O_360,N_4571,N_4713);
or UO_361 (O_361,N_4985,N_4807);
nand UO_362 (O_362,N_4696,N_4958);
nor UO_363 (O_363,N_4798,N_4568);
nand UO_364 (O_364,N_4735,N_4708);
nand UO_365 (O_365,N_4666,N_4969);
and UO_366 (O_366,N_4862,N_4883);
or UO_367 (O_367,N_4814,N_4504);
nor UO_368 (O_368,N_4570,N_4680);
nor UO_369 (O_369,N_4730,N_4788);
nor UO_370 (O_370,N_4954,N_4696);
nor UO_371 (O_371,N_4666,N_4824);
and UO_372 (O_372,N_4982,N_4902);
or UO_373 (O_373,N_4847,N_4591);
nand UO_374 (O_374,N_4864,N_4568);
nor UO_375 (O_375,N_4664,N_4807);
and UO_376 (O_376,N_4883,N_4956);
nor UO_377 (O_377,N_4655,N_4674);
and UO_378 (O_378,N_4583,N_4900);
or UO_379 (O_379,N_4862,N_4839);
nand UO_380 (O_380,N_4863,N_4628);
or UO_381 (O_381,N_4784,N_4606);
nand UO_382 (O_382,N_4572,N_4557);
nand UO_383 (O_383,N_4958,N_4683);
nand UO_384 (O_384,N_4612,N_4554);
and UO_385 (O_385,N_4696,N_4512);
and UO_386 (O_386,N_4812,N_4670);
or UO_387 (O_387,N_4819,N_4775);
nand UO_388 (O_388,N_4603,N_4697);
and UO_389 (O_389,N_4529,N_4972);
and UO_390 (O_390,N_4969,N_4794);
nand UO_391 (O_391,N_4855,N_4761);
nand UO_392 (O_392,N_4897,N_4582);
nand UO_393 (O_393,N_4986,N_4560);
nor UO_394 (O_394,N_4968,N_4760);
xor UO_395 (O_395,N_4530,N_4520);
and UO_396 (O_396,N_4567,N_4755);
and UO_397 (O_397,N_4779,N_4960);
or UO_398 (O_398,N_4546,N_4509);
xor UO_399 (O_399,N_4733,N_4978);
nand UO_400 (O_400,N_4876,N_4870);
nand UO_401 (O_401,N_4683,N_4657);
nor UO_402 (O_402,N_4990,N_4771);
nor UO_403 (O_403,N_4613,N_4616);
nor UO_404 (O_404,N_4534,N_4708);
and UO_405 (O_405,N_4675,N_4580);
nor UO_406 (O_406,N_4693,N_4534);
or UO_407 (O_407,N_4515,N_4592);
or UO_408 (O_408,N_4986,N_4534);
nand UO_409 (O_409,N_4790,N_4950);
or UO_410 (O_410,N_4633,N_4583);
xnor UO_411 (O_411,N_4949,N_4932);
nand UO_412 (O_412,N_4605,N_4732);
nor UO_413 (O_413,N_4672,N_4563);
or UO_414 (O_414,N_4929,N_4506);
and UO_415 (O_415,N_4825,N_4690);
and UO_416 (O_416,N_4610,N_4725);
and UO_417 (O_417,N_4645,N_4613);
nor UO_418 (O_418,N_4539,N_4935);
nand UO_419 (O_419,N_4873,N_4552);
nand UO_420 (O_420,N_4504,N_4999);
nand UO_421 (O_421,N_4610,N_4831);
or UO_422 (O_422,N_4851,N_4915);
nand UO_423 (O_423,N_4993,N_4678);
nand UO_424 (O_424,N_4662,N_4665);
and UO_425 (O_425,N_4511,N_4902);
or UO_426 (O_426,N_4925,N_4559);
and UO_427 (O_427,N_4809,N_4970);
nand UO_428 (O_428,N_4535,N_4599);
or UO_429 (O_429,N_4692,N_4840);
and UO_430 (O_430,N_4733,N_4925);
or UO_431 (O_431,N_4658,N_4531);
and UO_432 (O_432,N_4993,N_4671);
nand UO_433 (O_433,N_4958,N_4509);
nand UO_434 (O_434,N_4949,N_4880);
nand UO_435 (O_435,N_4994,N_4547);
and UO_436 (O_436,N_4704,N_4820);
and UO_437 (O_437,N_4987,N_4577);
nand UO_438 (O_438,N_4927,N_4960);
or UO_439 (O_439,N_4984,N_4602);
xnor UO_440 (O_440,N_4827,N_4517);
xnor UO_441 (O_441,N_4605,N_4691);
nor UO_442 (O_442,N_4892,N_4974);
nor UO_443 (O_443,N_4765,N_4907);
xor UO_444 (O_444,N_4824,N_4965);
and UO_445 (O_445,N_4672,N_4968);
nor UO_446 (O_446,N_4670,N_4605);
xnor UO_447 (O_447,N_4533,N_4795);
or UO_448 (O_448,N_4503,N_4760);
and UO_449 (O_449,N_4885,N_4969);
or UO_450 (O_450,N_4791,N_4552);
or UO_451 (O_451,N_4786,N_4654);
and UO_452 (O_452,N_4831,N_4989);
nor UO_453 (O_453,N_4607,N_4654);
nor UO_454 (O_454,N_4790,N_4833);
and UO_455 (O_455,N_4725,N_4792);
nor UO_456 (O_456,N_4567,N_4917);
and UO_457 (O_457,N_4872,N_4975);
nand UO_458 (O_458,N_4826,N_4849);
nand UO_459 (O_459,N_4958,N_4731);
nand UO_460 (O_460,N_4637,N_4895);
or UO_461 (O_461,N_4937,N_4874);
nor UO_462 (O_462,N_4593,N_4883);
or UO_463 (O_463,N_4939,N_4620);
and UO_464 (O_464,N_4889,N_4841);
nand UO_465 (O_465,N_4832,N_4544);
and UO_466 (O_466,N_4966,N_4509);
and UO_467 (O_467,N_4553,N_4823);
nor UO_468 (O_468,N_4727,N_4935);
or UO_469 (O_469,N_4505,N_4858);
nor UO_470 (O_470,N_4699,N_4648);
and UO_471 (O_471,N_4702,N_4908);
xnor UO_472 (O_472,N_4760,N_4953);
nor UO_473 (O_473,N_4584,N_4691);
nand UO_474 (O_474,N_4959,N_4507);
nand UO_475 (O_475,N_4734,N_4546);
nand UO_476 (O_476,N_4899,N_4655);
or UO_477 (O_477,N_4878,N_4751);
or UO_478 (O_478,N_4601,N_4610);
xnor UO_479 (O_479,N_4851,N_4809);
and UO_480 (O_480,N_4838,N_4505);
nand UO_481 (O_481,N_4705,N_4756);
nor UO_482 (O_482,N_4994,N_4985);
and UO_483 (O_483,N_4518,N_4686);
or UO_484 (O_484,N_4975,N_4640);
nor UO_485 (O_485,N_4636,N_4848);
nand UO_486 (O_486,N_4615,N_4573);
nor UO_487 (O_487,N_4783,N_4660);
nor UO_488 (O_488,N_4705,N_4755);
or UO_489 (O_489,N_4559,N_4898);
or UO_490 (O_490,N_4531,N_4886);
nand UO_491 (O_491,N_4870,N_4625);
or UO_492 (O_492,N_4809,N_4817);
and UO_493 (O_493,N_4547,N_4618);
xor UO_494 (O_494,N_4509,N_4962);
or UO_495 (O_495,N_4928,N_4653);
nand UO_496 (O_496,N_4784,N_4772);
or UO_497 (O_497,N_4752,N_4739);
nand UO_498 (O_498,N_4817,N_4551);
and UO_499 (O_499,N_4725,N_4863);
or UO_500 (O_500,N_4796,N_4959);
or UO_501 (O_501,N_4947,N_4993);
or UO_502 (O_502,N_4955,N_4805);
or UO_503 (O_503,N_4866,N_4766);
or UO_504 (O_504,N_4608,N_4715);
nand UO_505 (O_505,N_4878,N_4675);
or UO_506 (O_506,N_4796,N_4934);
or UO_507 (O_507,N_4734,N_4607);
nor UO_508 (O_508,N_4639,N_4919);
nand UO_509 (O_509,N_4726,N_4541);
or UO_510 (O_510,N_4508,N_4807);
xor UO_511 (O_511,N_4747,N_4900);
or UO_512 (O_512,N_4694,N_4688);
or UO_513 (O_513,N_4643,N_4780);
nor UO_514 (O_514,N_4503,N_4727);
nor UO_515 (O_515,N_4802,N_4677);
or UO_516 (O_516,N_4800,N_4769);
nor UO_517 (O_517,N_4585,N_4519);
or UO_518 (O_518,N_4948,N_4648);
nand UO_519 (O_519,N_4749,N_4953);
nor UO_520 (O_520,N_4612,N_4936);
nand UO_521 (O_521,N_4507,N_4882);
nor UO_522 (O_522,N_4983,N_4802);
and UO_523 (O_523,N_4994,N_4861);
nor UO_524 (O_524,N_4821,N_4761);
nand UO_525 (O_525,N_4894,N_4827);
nand UO_526 (O_526,N_4635,N_4691);
or UO_527 (O_527,N_4749,N_4835);
and UO_528 (O_528,N_4918,N_4582);
and UO_529 (O_529,N_4558,N_4920);
and UO_530 (O_530,N_4515,N_4630);
and UO_531 (O_531,N_4592,N_4552);
nand UO_532 (O_532,N_4679,N_4686);
nor UO_533 (O_533,N_4834,N_4889);
nor UO_534 (O_534,N_4678,N_4631);
nand UO_535 (O_535,N_4888,N_4626);
nor UO_536 (O_536,N_4827,N_4957);
and UO_537 (O_537,N_4611,N_4535);
nor UO_538 (O_538,N_4629,N_4759);
or UO_539 (O_539,N_4743,N_4756);
and UO_540 (O_540,N_4617,N_4648);
or UO_541 (O_541,N_4652,N_4643);
nand UO_542 (O_542,N_4671,N_4856);
and UO_543 (O_543,N_4940,N_4945);
nand UO_544 (O_544,N_4875,N_4890);
xor UO_545 (O_545,N_4948,N_4923);
and UO_546 (O_546,N_4846,N_4684);
xor UO_547 (O_547,N_4931,N_4766);
or UO_548 (O_548,N_4573,N_4782);
and UO_549 (O_549,N_4763,N_4963);
and UO_550 (O_550,N_4768,N_4740);
nand UO_551 (O_551,N_4571,N_4832);
or UO_552 (O_552,N_4510,N_4624);
nand UO_553 (O_553,N_4667,N_4992);
nand UO_554 (O_554,N_4605,N_4919);
or UO_555 (O_555,N_4610,N_4720);
nor UO_556 (O_556,N_4861,N_4943);
nand UO_557 (O_557,N_4776,N_4650);
or UO_558 (O_558,N_4555,N_4545);
nand UO_559 (O_559,N_4534,N_4825);
xnor UO_560 (O_560,N_4724,N_4698);
or UO_561 (O_561,N_4508,N_4819);
or UO_562 (O_562,N_4575,N_4550);
nor UO_563 (O_563,N_4659,N_4626);
nand UO_564 (O_564,N_4538,N_4546);
nand UO_565 (O_565,N_4588,N_4660);
nand UO_566 (O_566,N_4973,N_4930);
or UO_567 (O_567,N_4790,N_4872);
nor UO_568 (O_568,N_4997,N_4755);
or UO_569 (O_569,N_4506,N_4803);
and UO_570 (O_570,N_4935,N_4982);
nand UO_571 (O_571,N_4568,N_4587);
or UO_572 (O_572,N_4965,N_4820);
or UO_573 (O_573,N_4994,N_4741);
and UO_574 (O_574,N_4941,N_4822);
nor UO_575 (O_575,N_4799,N_4512);
nor UO_576 (O_576,N_4898,N_4557);
nor UO_577 (O_577,N_4595,N_4642);
and UO_578 (O_578,N_4968,N_4827);
nor UO_579 (O_579,N_4791,N_4693);
or UO_580 (O_580,N_4601,N_4512);
or UO_581 (O_581,N_4887,N_4682);
nor UO_582 (O_582,N_4930,N_4608);
nand UO_583 (O_583,N_4544,N_4874);
nand UO_584 (O_584,N_4516,N_4989);
nand UO_585 (O_585,N_4729,N_4543);
or UO_586 (O_586,N_4691,N_4760);
or UO_587 (O_587,N_4562,N_4761);
or UO_588 (O_588,N_4714,N_4943);
nand UO_589 (O_589,N_4617,N_4719);
or UO_590 (O_590,N_4825,N_4890);
xnor UO_591 (O_591,N_4791,N_4599);
nor UO_592 (O_592,N_4638,N_4590);
nand UO_593 (O_593,N_4603,N_4850);
nor UO_594 (O_594,N_4983,N_4857);
or UO_595 (O_595,N_4932,N_4896);
nor UO_596 (O_596,N_4826,N_4763);
or UO_597 (O_597,N_4954,N_4582);
nor UO_598 (O_598,N_4691,N_4572);
nor UO_599 (O_599,N_4660,N_4685);
xor UO_600 (O_600,N_4979,N_4823);
or UO_601 (O_601,N_4915,N_4583);
or UO_602 (O_602,N_4798,N_4727);
xnor UO_603 (O_603,N_4666,N_4843);
nor UO_604 (O_604,N_4698,N_4894);
and UO_605 (O_605,N_4754,N_4887);
nand UO_606 (O_606,N_4921,N_4824);
or UO_607 (O_607,N_4861,N_4838);
or UO_608 (O_608,N_4943,N_4880);
nor UO_609 (O_609,N_4990,N_4794);
xnor UO_610 (O_610,N_4516,N_4787);
nand UO_611 (O_611,N_4734,N_4786);
nand UO_612 (O_612,N_4740,N_4636);
nand UO_613 (O_613,N_4680,N_4819);
or UO_614 (O_614,N_4570,N_4702);
or UO_615 (O_615,N_4952,N_4589);
nor UO_616 (O_616,N_4669,N_4601);
and UO_617 (O_617,N_4749,N_4811);
and UO_618 (O_618,N_4520,N_4784);
nand UO_619 (O_619,N_4514,N_4964);
xnor UO_620 (O_620,N_4591,N_4616);
xnor UO_621 (O_621,N_4695,N_4795);
nand UO_622 (O_622,N_4724,N_4699);
nand UO_623 (O_623,N_4500,N_4644);
and UO_624 (O_624,N_4532,N_4696);
xor UO_625 (O_625,N_4513,N_4669);
or UO_626 (O_626,N_4799,N_4541);
and UO_627 (O_627,N_4773,N_4770);
and UO_628 (O_628,N_4806,N_4600);
nor UO_629 (O_629,N_4910,N_4622);
nor UO_630 (O_630,N_4741,N_4970);
nor UO_631 (O_631,N_4928,N_4652);
nand UO_632 (O_632,N_4708,N_4825);
or UO_633 (O_633,N_4906,N_4510);
nand UO_634 (O_634,N_4992,N_4594);
xnor UO_635 (O_635,N_4555,N_4827);
nand UO_636 (O_636,N_4758,N_4552);
or UO_637 (O_637,N_4595,N_4555);
xnor UO_638 (O_638,N_4806,N_4960);
nand UO_639 (O_639,N_4987,N_4683);
and UO_640 (O_640,N_4551,N_4998);
nand UO_641 (O_641,N_4598,N_4751);
and UO_642 (O_642,N_4835,N_4734);
nor UO_643 (O_643,N_4896,N_4599);
and UO_644 (O_644,N_4522,N_4842);
or UO_645 (O_645,N_4601,N_4622);
or UO_646 (O_646,N_4560,N_4977);
xor UO_647 (O_647,N_4908,N_4657);
and UO_648 (O_648,N_4717,N_4763);
nor UO_649 (O_649,N_4958,N_4751);
or UO_650 (O_650,N_4917,N_4938);
and UO_651 (O_651,N_4847,N_4599);
or UO_652 (O_652,N_4585,N_4726);
xor UO_653 (O_653,N_4733,N_4557);
or UO_654 (O_654,N_4857,N_4747);
nand UO_655 (O_655,N_4956,N_4579);
nor UO_656 (O_656,N_4635,N_4854);
and UO_657 (O_657,N_4983,N_4612);
or UO_658 (O_658,N_4877,N_4850);
and UO_659 (O_659,N_4675,N_4998);
nand UO_660 (O_660,N_4827,N_4831);
or UO_661 (O_661,N_4845,N_4620);
nand UO_662 (O_662,N_4663,N_4905);
xor UO_663 (O_663,N_4947,N_4827);
and UO_664 (O_664,N_4913,N_4749);
or UO_665 (O_665,N_4704,N_4854);
or UO_666 (O_666,N_4750,N_4541);
nor UO_667 (O_667,N_4722,N_4628);
and UO_668 (O_668,N_4836,N_4599);
or UO_669 (O_669,N_4834,N_4542);
nand UO_670 (O_670,N_4686,N_4726);
or UO_671 (O_671,N_4687,N_4700);
nor UO_672 (O_672,N_4804,N_4721);
and UO_673 (O_673,N_4591,N_4744);
nand UO_674 (O_674,N_4917,N_4642);
and UO_675 (O_675,N_4766,N_4895);
and UO_676 (O_676,N_4923,N_4934);
nor UO_677 (O_677,N_4676,N_4788);
or UO_678 (O_678,N_4899,N_4782);
nand UO_679 (O_679,N_4820,N_4863);
and UO_680 (O_680,N_4541,N_4585);
or UO_681 (O_681,N_4664,N_4741);
nor UO_682 (O_682,N_4563,N_4983);
or UO_683 (O_683,N_4951,N_4587);
or UO_684 (O_684,N_4850,N_4691);
and UO_685 (O_685,N_4621,N_4748);
nand UO_686 (O_686,N_4523,N_4510);
and UO_687 (O_687,N_4851,N_4933);
or UO_688 (O_688,N_4516,N_4663);
or UO_689 (O_689,N_4986,N_4985);
or UO_690 (O_690,N_4620,N_4832);
nor UO_691 (O_691,N_4784,N_4693);
nor UO_692 (O_692,N_4699,N_4800);
and UO_693 (O_693,N_4932,N_4567);
or UO_694 (O_694,N_4652,N_4511);
nand UO_695 (O_695,N_4749,N_4946);
nand UO_696 (O_696,N_4826,N_4985);
or UO_697 (O_697,N_4796,N_4747);
and UO_698 (O_698,N_4883,N_4832);
and UO_699 (O_699,N_4746,N_4942);
and UO_700 (O_700,N_4978,N_4813);
nand UO_701 (O_701,N_4557,N_4868);
nand UO_702 (O_702,N_4993,N_4841);
nor UO_703 (O_703,N_4713,N_4916);
and UO_704 (O_704,N_4600,N_4734);
xor UO_705 (O_705,N_4955,N_4681);
nor UO_706 (O_706,N_4880,N_4821);
nand UO_707 (O_707,N_4638,N_4893);
nor UO_708 (O_708,N_4975,N_4964);
nor UO_709 (O_709,N_4995,N_4926);
nor UO_710 (O_710,N_4630,N_4518);
and UO_711 (O_711,N_4861,N_4626);
nand UO_712 (O_712,N_4564,N_4961);
nand UO_713 (O_713,N_4639,N_4948);
xor UO_714 (O_714,N_4886,N_4553);
nor UO_715 (O_715,N_4551,N_4660);
nand UO_716 (O_716,N_4957,N_4618);
nand UO_717 (O_717,N_4904,N_4987);
nand UO_718 (O_718,N_4531,N_4743);
nand UO_719 (O_719,N_4536,N_4840);
or UO_720 (O_720,N_4550,N_4854);
or UO_721 (O_721,N_4953,N_4756);
or UO_722 (O_722,N_4638,N_4801);
or UO_723 (O_723,N_4879,N_4846);
or UO_724 (O_724,N_4897,N_4722);
and UO_725 (O_725,N_4515,N_4626);
xnor UO_726 (O_726,N_4973,N_4947);
or UO_727 (O_727,N_4918,N_4548);
or UO_728 (O_728,N_4671,N_4988);
nor UO_729 (O_729,N_4977,N_4633);
or UO_730 (O_730,N_4816,N_4525);
xor UO_731 (O_731,N_4990,N_4692);
nor UO_732 (O_732,N_4920,N_4771);
or UO_733 (O_733,N_4762,N_4864);
nand UO_734 (O_734,N_4669,N_4922);
or UO_735 (O_735,N_4668,N_4917);
nand UO_736 (O_736,N_4524,N_4672);
nor UO_737 (O_737,N_4889,N_4905);
or UO_738 (O_738,N_4952,N_4898);
nand UO_739 (O_739,N_4608,N_4884);
nor UO_740 (O_740,N_4546,N_4816);
or UO_741 (O_741,N_4988,N_4856);
or UO_742 (O_742,N_4601,N_4965);
xor UO_743 (O_743,N_4547,N_4835);
and UO_744 (O_744,N_4631,N_4793);
or UO_745 (O_745,N_4652,N_4558);
nand UO_746 (O_746,N_4660,N_4811);
and UO_747 (O_747,N_4930,N_4895);
and UO_748 (O_748,N_4914,N_4813);
and UO_749 (O_749,N_4960,N_4986);
and UO_750 (O_750,N_4526,N_4972);
or UO_751 (O_751,N_4505,N_4814);
and UO_752 (O_752,N_4615,N_4759);
or UO_753 (O_753,N_4741,N_4799);
nor UO_754 (O_754,N_4614,N_4500);
nand UO_755 (O_755,N_4752,N_4919);
xnor UO_756 (O_756,N_4853,N_4611);
and UO_757 (O_757,N_4738,N_4890);
and UO_758 (O_758,N_4743,N_4523);
nand UO_759 (O_759,N_4774,N_4967);
nor UO_760 (O_760,N_4520,N_4756);
or UO_761 (O_761,N_4844,N_4953);
and UO_762 (O_762,N_4593,N_4633);
and UO_763 (O_763,N_4741,N_4990);
nand UO_764 (O_764,N_4816,N_4757);
xor UO_765 (O_765,N_4545,N_4551);
nand UO_766 (O_766,N_4846,N_4822);
and UO_767 (O_767,N_4913,N_4796);
nor UO_768 (O_768,N_4913,N_4562);
nand UO_769 (O_769,N_4903,N_4877);
or UO_770 (O_770,N_4617,N_4867);
nand UO_771 (O_771,N_4946,N_4635);
and UO_772 (O_772,N_4821,N_4723);
nand UO_773 (O_773,N_4656,N_4655);
or UO_774 (O_774,N_4887,N_4696);
or UO_775 (O_775,N_4694,N_4712);
nor UO_776 (O_776,N_4878,N_4610);
and UO_777 (O_777,N_4693,N_4529);
nor UO_778 (O_778,N_4565,N_4793);
and UO_779 (O_779,N_4541,N_4601);
and UO_780 (O_780,N_4604,N_4668);
xnor UO_781 (O_781,N_4642,N_4988);
or UO_782 (O_782,N_4806,N_4704);
and UO_783 (O_783,N_4605,N_4772);
nor UO_784 (O_784,N_4874,N_4885);
nand UO_785 (O_785,N_4744,N_4571);
nor UO_786 (O_786,N_4800,N_4655);
or UO_787 (O_787,N_4982,N_4855);
or UO_788 (O_788,N_4950,N_4624);
and UO_789 (O_789,N_4647,N_4761);
nor UO_790 (O_790,N_4835,N_4534);
xnor UO_791 (O_791,N_4686,N_4837);
nor UO_792 (O_792,N_4529,N_4863);
nand UO_793 (O_793,N_4540,N_4620);
nor UO_794 (O_794,N_4833,N_4865);
and UO_795 (O_795,N_4923,N_4991);
or UO_796 (O_796,N_4554,N_4572);
or UO_797 (O_797,N_4855,N_4926);
or UO_798 (O_798,N_4727,N_4838);
and UO_799 (O_799,N_4618,N_4716);
and UO_800 (O_800,N_4926,N_4571);
xnor UO_801 (O_801,N_4501,N_4760);
and UO_802 (O_802,N_4950,N_4711);
and UO_803 (O_803,N_4566,N_4876);
nor UO_804 (O_804,N_4654,N_4766);
nand UO_805 (O_805,N_4534,N_4900);
xnor UO_806 (O_806,N_4523,N_4753);
nand UO_807 (O_807,N_4534,N_4812);
nor UO_808 (O_808,N_4546,N_4923);
nor UO_809 (O_809,N_4711,N_4525);
or UO_810 (O_810,N_4618,N_4610);
or UO_811 (O_811,N_4707,N_4565);
nor UO_812 (O_812,N_4623,N_4660);
or UO_813 (O_813,N_4710,N_4754);
and UO_814 (O_814,N_4761,N_4521);
nor UO_815 (O_815,N_4573,N_4622);
nand UO_816 (O_816,N_4677,N_4948);
nand UO_817 (O_817,N_4724,N_4986);
and UO_818 (O_818,N_4725,N_4885);
nor UO_819 (O_819,N_4890,N_4542);
nand UO_820 (O_820,N_4868,N_4859);
nand UO_821 (O_821,N_4832,N_4803);
nor UO_822 (O_822,N_4904,N_4636);
xnor UO_823 (O_823,N_4654,N_4952);
nand UO_824 (O_824,N_4944,N_4929);
or UO_825 (O_825,N_4797,N_4515);
xnor UO_826 (O_826,N_4836,N_4610);
nand UO_827 (O_827,N_4544,N_4987);
nand UO_828 (O_828,N_4998,N_4619);
xnor UO_829 (O_829,N_4666,N_4829);
nand UO_830 (O_830,N_4596,N_4697);
and UO_831 (O_831,N_4739,N_4935);
nand UO_832 (O_832,N_4731,N_4584);
and UO_833 (O_833,N_4878,N_4834);
nor UO_834 (O_834,N_4717,N_4621);
and UO_835 (O_835,N_4637,N_4747);
nor UO_836 (O_836,N_4892,N_4688);
nor UO_837 (O_837,N_4745,N_4724);
nor UO_838 (O_838,N_4551,N_4995);
and UO_839 (O_839,N_4845,N_4848);
and UO_840 (O_840,N_4904,N_4944);
nor UO_841 (O_841,N_4897,N_4688);
and UO_842 (O_842,N_4912,N_4678);
nor UO_843 (O_843,N_4885,N_4994);
xnor UO_844 (O_844,N_4612,N_4974);
and UO_845 (O_845,N_4971,N_4846);
nor UO_846 (O_846,N_4890,N_4909);
nand UO_847 (O_847,N_4989,N_4887);
and UO_848 (O_848,N_4871,N_4946);
or UO_849 (O_849,N_4661,N_4744);
or UO_850 (O_850,N_4696,N_4955);
and UO_851 (O_851,N_4758,N_4556);
or UO_852 (O_852,N_4824,N_4578);
or UO_853 (O_853,N_4900,N_4738);
xor UO_854 (O_854,N_4613,N_4982);
nor UO_855 (O_855,N_4534,N_4845);
nor UO_856 (O_856,N_4629,N_4664);
nand UO_857 (O_857,N_4517,N_4943);
nor UO_858 (O_858,N_4960,N_4886);
and UO_859 (O_859,N_4660,N_4836);
nand UO_860 (O_860,N_4699,N_4624);
nor UO_861 (O_861,N_4929,N_4846);
nor UO_862 (O_862,N_4925,N_4728);
and UO_863 (O_863,N_4833,N_4632);
or UO_864 (O_864,N_4554,N_4729);
nand UO_865 (O_865,N_4924,N_4558);
and UO_866 (O_866,N_4804,N_4748);
nor UO_867 (O_867,N_4995,N_4650);
xnor UO_868 (O_868,N_4794,N_4812);
nor UO_869 (O_869,N_4615,N_4839);
and UO_870 (O_870,N_4817,N_4747);
nand UO_871 (O_871,N_4647,N_4794);
nor UO_872 (O_872,N_4827,N_4792);
or UO_873 (O_873,N_4727,N_4847);
or UO_874 (O_874,N_4714,N_4743);
and UO_875 (O_875,N_4831,N_4824);
or UO_876 (O_876,N_4864,N_4720);
or UO_877 (O_877,N_4801,N_4959);
and UO_878 (O_878,N_4783,N_4965);
or UO_879 (O_879,N_4722,N_4727);
nand UO_880 (O_880,N_4726,N_4800);
nor UO_881 (O_881,N_4795,N_4607);
and UO_882 (O_882,N_4567,N_4547);
and UO_883 (O_883,N_4971,N_4653);
and UO_884 (O_884,N_4631,N_4783);
and UO_885 (O_885,N_4768,N_4737);
nand UO_886 (O_886,N_4620,N_4994);
or UO_887 (O_887,N_4819,N_4821);
and UO_888 (O_888,N_4609,N_4977);
nand UO_889 (O_889,N_4849,N_4638);
nor UO_890 (O_890,N_4580,N_4825);
and UO_891 (O_891,N_4565,N_4553);
or UO_892 (O_892,N_4502,N_4736);
and UO_893 (O_893,N_4870,N_4639);
or UO_894 (O_894,N_4758,N_4561);
nor UO_895 (O_895,N_4756,N_4817);
nor UO_896 (O_896,N_4719,N_4620);
and UO_897 (O_897,N_4616,N_4559);
nor UO_898 (O_898,N_4944,N_4956);
nor UO_899 (O_899,N_4898,N_4710);
nand UO_900 (O_900,N_4762,N_4625);
or UO_901 (O_901,N_4716,N_4594);
nand UO_902 (O_902,N_4888,N_4612);
and UO_903 (O_903,N_4728,N_4918);
nand UO_904 (O_904,N_4687,N_4739);
or UO_905 (O_905,N_4765,N_4989);
and UO_906 (O_906,N_4575,N_4617);
or UO_907 (O_907,N_4694,N_4678);
nand UO_908 (O_908,N_4748,N_4643);
nand UO_909 (O_909,N_4930,N_4939);
nand UO_910 (O_910,N_4757,N_4865);
or UO_911 (O_911,N_4894,N_4788);
or UO_912 (O_912,N_4594,N_4520);
and UO_913 (O_913,N_4902,N_4871);
and UO_914 (O_914,N_4656,N_4507);
nor UO_915 (O_915,N_4598,N_4807);
xor UO_916 (O_916,N_4594,N_4620);
xnor UO_917 (O_917,N_4620,N_4596);
or UO_918 (O_918,N_4558,N_4886);
xor UO_919 (O_919,N_4970,N_4750);
nor UO_920 (O_920,N_4865,N_4706);
nor UO_921 (O_921,N_4695,N_4689);
or UO_922 (O_922,N_4921,N_4508);
or UO_923 (O_923,N_4681,N_4947);
nand UO_924 (O_924,N_4999,N_4950);
nor UO_925 (O_925,N_4544,N_4793);
nor UO_926 (O_926,N_4808,N_4772);
nand UO_927 (O_927,N_4808,N_4665);
or UO_928 (O_928,N_4876,N_4900);
nor UO_929 (O_929,N_4892,N_4590);
and UO_930 (O_930,N_4707,N_4558);
nor UO_931 (O_931,N_4748,N_4942);
or UO_932 (O_932,N_4628,N_4867);
or UO_933 (O_933,N_4979,N_4581);
or UO_934 (O_934,N_4532,N_4743);
nor UO_935 (O_935,N_4873,N_4734);
or UO_936 (O_936,N_4517,N_4763);
or UO_937 (O_937,N_4991,N_4831);
xor UO_938 (O_938,N_4960,N_4965);
nor UO_939 (O_939,N_4840,N_4776);
and UO_940 (O_940,N_4617,N_4661);
xnor UO_941 (O_941,N_4962,N_4851);
nor UO_942 (O_942,N_4589,N_4578);
or UO_943 (O_943,N_4912,N_4795);
and UO_944 (O_944,N_4887,N_4927);
nor UO_945 (O_945,N_4616,N_4711);
nor UO_946 (O_946,N_4795,N_4859);
nand UO_947 (O_947,N_4911,N_4652);
nor UO_948 (O_948,N_4871,N_4760);
xnor UO_949 (O_949,N_4699,N_4982);
or UO_950 (O_950,N_4547,N_4719);
nor UO_951 (O_951,N_4579,N_4520);
and UO_952 (O_952,N_4551,N_4586);
nand UO_953 (O_953,N_4977,N_4635);
nor UO_954 (O_954,N_4966,N_4856);
or UO_955 (O_955,N_4689,N_4817);
or UO_956 (O_956,N_4767,N_4868);
nand UO_957 (O_957,N_4563,N_4892);
nand UO_958 (O_958,N_4780,N_4652);
nor UO_959 (O_959,N_4628,N_4904);
or UO_960 (O_960,N_4953,N_4858);
nand UO_961 (O_961,N_4813,N_4684);
nor UO_962 (O_962,N_4960,N_4503);
or UO_963 (O_963,N_4705,N_4604);
xor UO_964 (O_964,N_4963,N_4791);
nor UO_965 (O_965,N_4957,N_4933);
nand UO_966 (O_966,N_4904,N_4501);
nor UO_967 (O_967,N_4842,N_4817);
or UO_968 (O_968,N_4593,N_4578);
xnor UO_969 (O_969,N_4679,N_4938);
nor UO_970 (O_970,N_4708,N_4751);
and UO_971 (O_971,N_4530,N_4709);
nor UO_972 (O_972,N_4603,N_4537);
nand UO_973 (O_973,N_4751,N_4686);
or UO_974 (O_974,N_4578,N_4708);
nor UO_975 (O_975,N_4856,N_4774);
or UO_976 (O_976,N_4913,N_4631);
xnor UO_977 (O_977,N_4703,N_4513);
and UO_978 (O_978,N_4906,N_4502);
and UO_979 (O_979,N_4677,N_4768);
nand UO_980 (O_980,N_4865,N_4967);
and UO_981 (O_981,N_4561,N_4711);
and UO_982 (O_982,N_4515,N_4608);
and UO_983 (O_983,N_4906,N_4840);
or UO_984 (O_984,N_4610,N_4557);
and UO_985 (O_985,N_4526,N_4828);
and UO_986 (O_986,N_4930,N_4885);
or UO_987 (O_987,N_4554,N_4955);
nand UO_988 (O_988,N_4914,N_4796);
nand UO_989 (O_989,N_4850,N_4899);
nand UO_990 (O_990,N_4511,N_4593);
or UO_991 (O_991,N_4981,N_4797);
nor UO_992 (O_992,N_4536,N_4634);
or UO_993 (O_993,N_4929,N_4722);
nand UO_994 (O_994,N_4963,N_4728);
and UO_995 (O_995,N_4951,N_4832);
and UO_996 (O_996,N_4962,N_4956);
nand UO_997 (O_997,N_4788,N_4541);
and UO_998 (O_998,N_4662,N_4869);
and UO_999 (O_999,N_4558,N_4830);
endmodule