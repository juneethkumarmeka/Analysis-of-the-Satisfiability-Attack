module basic_500_3000_500_60_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_170,In_497);
nand U1 (N_1,In_141,In_225);
nand U2 (N_2,In_331,In_407);
nor U3 (N_3,In_334,In_479);
and U4 (N_4,In_483,In_143);
or U5 (N_5,In_60,In_104);
or U6 (N_6,In_159,In_464);
and U7 (N_7,In_498,In_97);
nor U8 (N_8,In_129,In_138);
nand U9 (N_9,In_163,In_108);
or U10 (N_10,In_357,In_128);
or U11 (N_11,In_8,In_297);
nand U12 (N_12,In_183,In_124);
or U13 (N_13,In_413,In_388);
and U14 (N_14,In_194,In_311);
or U15 (N_15,In_121,In_445);
nand U16 (N_16,In_385,In_476);
nand U17 (N_17,In_323,In_294);
or U18 (N_18,In_375,In_230);
and U19 (N_19,In_0,In_154);
nor U20 (N_20,In_342,In_283);
nor U21 (N_21,In_228,In_290);
or U22 (N_22,In_161,In_303);
nand U23 (N_23,In_463,In_231);
nor U24 (N_24,In_412,In_247);
nor U25 (N_25,In_343,In_282);
and U26 (N_26,In_434,In_68);
nand U27 (N_27,In_49,In_236);
or U28 (N_28,In_246,In_160);
and U29 (N_29,In_379,In_279);
nand U30 (N_30,In_115,In_269);
or U31 (N_31,In_111,In_245);
nand U32 (N_32,In_299,In_372);
nand U33 (N_33,In_140,In_196);
nor U34 (N_34,In_472,In_447);
nor U35 (N_35,In_75,In_201);
and U36 (N_36,In_190,In_178);
nor U37 (N_37,In_289,In_10);
nand U38 (N_38,In_244,In_376);
nand U39 (N_39,In_264,In_36);
nand U40 (N_40,In_136,In_329);
and U41 (N_41,In_287,In_112);
or U42 (N_42,In_38,In_274);
and U43 (N_43,In_281,In_81);
nand U44 (N_44,In_226,In_465);
and U45 (N_45,In_48,In_195);
xor U46 (N_46,In_370,In_355);
and U47 (N_47,In_489,In_448);
or U48 (N_48,In_272,In_318);
and U49 (N_49,In_17,In_53);
nor U50 (N_50,N_18,In_213);
and U51 (N_51,In_4,In_384);
and U52 (N_52,In_458,In_389);
nand U53 (N_53,In_198,In_18);
and U54 (N_54,In_87,In_471);
nand U55 (N_55,In_23,In_485);
nor U56 (N_56,N_35,In_452);
and U57 (N_57,In_100,In_52);
nor U58 (N_58,In_133,In_31);
or U59 (N_59,In_66,In_344);
and U60 (N_60,In_171,In_98);
nand U61 (N_61,In_59,In_250);
nor U62 (N_62,In_371,In_227);
or U63 (N_63,In_152,In_340);
nand U64 (N_64,In_150,In_401);
or U65 (N_65,N_24,In_260);
nor U66 (N_66,In_442,In_288);
nor U67 (N_67,In_267,N_41);
nor U68 (N_68,In_78,In_107);
or U69 (N_69,In_216,In_433);
and U70 (N_70,N_44,In_429);
and U71 (N_71,In_335,In_450);
nor U72 (N_72,In_238,In_324);
or U73 (N_73,In_271,In_117);
or U74 (N_74,In_494,In_220);
or U75 (N_75,In_45,In_223);
or U76 (N_76,In_263,In_35);
or U77 (N_77,In_469,In_16);
and U78 (N_78,In_113,In_417);
or U79 (N_79,In_387,In_364);
and U80 (N_80,In_421,In_484);
nand U81 (N_81,In_467,N_27);
or U82 (N_82,In_73,In_293);
and U83 (N_83,N_10,In_224);
nor U84 (N_84,In_253,In_7);
nor U85 (N_85,N_12,In_168);
nand U86 (N_86,In_395,In_317);
and U87 (N_87,In_90,In_427);
or U88 (N_88,N_25,In_425);
or U89 (N_89,In_5,In_431);
and U90 (N_90,In_22,In_188);
nand U91 (N_91,In_56,In_157);
or U92 (N_92,In_339,In_235);
nand U93 (N_93,In_208,In_306);
nand U94 (N_94,In_301,In_257);
and U95 (N_95,In_446,In_94);
nand U96 (N_96,In_30,In_424);
or U97 (N_97,N_14,In_74);
nor U98 (N_98,In_482,In_27);
or U99 (N_99,In_219,N_11);
xor U100 (N_100,In_34,N_78);
nand U101 (N_101,In_89,In_423);
and U102 (N_102,In_80,In_3);
or U103 (N_103,In_173,In_258);
and U104 (N_104,In_474,N_76);
or U105 (N_105,In_416,In_268);
or U106 (N_106,In_93,N_49);
nand U107 (N_107,In_391,N_45);
nor U108 (N_108,In_347,N_79);
nand U109 (N_109,In_346,In_459);
nor U110 (N_110,In_153,In_312);
nor U111 (N_111,In_480,In_41);
nor U112 (N_112,In_278,N_85);
and U113 (N_113,In_47,In_475);
or U114 (N_114,In_2,In_210);
or U115 (N_115,In_72,N_80);
or U116 (N_116,In_39,In_217);
or U117 (N_117,In_449,N_29);
or U118 (N_118,In_63,In_350);
nand U119 (N_119,In_135,In_266);
nor U120 (N_120,In_369,In_277);
nor U121 (N_121,In_396,In_300);
nor U122 (N_122,In_130,N_5);
nor U123 (N_123,In_13,In_46);
nor U124 (N_124,In_214,In_197);
nor U125 (N_125,In_358,In_50);
nand U126 (N_126,In_305,In_451);
or U127 (N_127,N_90,In_259);
and U128 (N_128,In_119,In_9);
nand U129 (N_129,In_79,In_116);
or U130 (N_130,In_187,N_57);
nor U131 (N_131,In_212,In_313);
xnor U132 (N_132,In_54,In_373);
and U133 (N_133,In_348,N_2);
nor U134 (N_134,In_462,N_20);
or U135 (N_135,N_92,In_256);
and U136 (N_136,In_106,N_47);
or U137 (N_137,In_105,In_356);
and U138 (N_138,In_304,In_182);
or U139 (N_139,N_13,In_310);
nor U140 (N_140,In_248,N_65);
nand U141 (N_141,N_33,In_67);
nor U142 (N_142,In_298,N_67);
or U143 (N_143,In_354,In_481);
nand U144 (N_144,In_363,In_207);
and U145 (N_145,In_125,N_23);
nand U146 (N_146,N_46,In_65);
or U147 (N_147,In_443,In_499);
nor U148 (N_148,In_349,In_408);
and U149 (N_149,In_493,N_38);
nand U150 (N_150,N_103,In_1);
or U151 (N_151,N_68,N_15);
and U152 (N_152,N_26,In_441);
and U153 (N_153,N_22,N_139);
nand U154 (N_154,In_490,N_94);
or U155 (N_155,In_166,In_209);
or U156 (N_156,N_34,In_205);
and U157 (N_157,In_418,In_134);
and U158 (N_158,N_148,In_333);
or U159 (N_159,N_8,In_14);
and U160 (N_160,In_162,In_202);
nand U161 (N_161,N_135,In_394);
xor U162 (N_162,N_127,N_66);
or U163 (N_163,In_176,In_234);
nor U164 (N_164,N_37,N_73);
and U165 (N_165,In_11,N_39);
and U166 (N_166,In_92,N_6);
and U167 (N_167,N_7,In_203);
nor U168 (N_168,In_148,In_437);
and U169 (N_169,In_167,N_123);
nand U170 (N_170,N_77,In_122);
nand U171 (N_171,In_237,In_273);
nor U172 (N_172,In_12,N_0);
nor U173 (N_173,In_88,In_345);
nand U174 (N_174,In_131,In_222);
nor U175 (N_175,In_142,In_383);
or U176 (N_176,In_316,N_43);
nand U177 (N_177,In_145,In_221);
or U178 (N_178,In_118,In_399);
nand U179 (N_179,In_478,N_98);
or U180 (N_180,In_460,In_57);
and U181 (N_181,N_70,In_366);
and U182 (N_182,In_398,In_326);
nor U183 (N_183,N_142,In_193);
nor U184 (N_184,In_26,In_314);
nand U185 (N_185,In_101,In_359);
nor U186 (N_186,In_496,In_155);
nor U187 (N_187,N_88,N_97);
nor U188 (N_188,In_428,In_19);
nor U189 (N_189,In_32,In_420);
nand U190 (N_190,In_491,In_454);
and U191 (N_191,In_432,N_87);
nand U192 (N_192,In_139,In_95);
nand U193 (N_193,In_6,In_204);
or U194 (N_194,N_115,N_64);
nor U195 (N_195,In_164,In_172);
or U196 (N_196,In_62,In_186);
and U197 (N_197,In_33,In_103);
and U198 (N_198,In_147,In_96);
nor U199 (N_199,In_200,In_189);
or U200 (N_200,In_422,In_365);
and U201 (N_201,N_21,N_102);
nand U202 (N_202,N_50,In_99);
nor U203 (N_203,N_156,N_143);
and U204 (N_204,N_188,In_308);
and U205 (N_205,In_495,In_243);
and U206 (N_206,N_93,N_178);
and U207 (N_207,N_164,In_319);
nand U208 (N_208,N_126,In_20);
nand U209 (N_209,N_128,N_175);
or U210 (N_210,In_120,In_165);
or U211 (N_211,In_492,N_72);
nand U212 (N_212,In_151,N_169);
or U213 (N_213,N_129,In_453);
and U214 (N_214,N_189,In_40);
or U215 (N_215,In_102,In_132);
and U216 (N_216,N_125,In_232);
and U217 (N_217,N_157,In_367);
nand U218 (N_218,In_240,N_160);
nor U219 (N_219,N_131,In_411);
and U220 (N_220,In_127,In_261);
and U221 (N_221,In_486,In_351);
nor U222 (N_222,In_21,In_175);
nand U223 (N_223,N_28,In_158);
or U224 (N_224,In_61,N_120);
xor U225 (N_225,N_161,N_190);
nand U226 (N_226,In_415,N_30);
nor U227 (N_227,N_81,In_206);
nand U228 (N_228,In_336,In_361);
or U229 (N_229,N_54,N_150);
nor U230 (N_230,In_402,N_60);
and U231 (N_231,In_114,In_77);
or U232 (N_232,In_332,In_380);
or U233 (N_233,In_275,In_215);
nand U234 (N_234,N_195,In_315);
nand U235 (N_235,In_262,In_320);
or U236 (N_236,N_113,In_382);
and U237 (N_237,N_153,N_184);
or U238 (N_238,In_286,In_252);
or U239 (N_239,N_144,N_179);
and U240 (N_240,N_105,N_36);
and U241 (N_241,In_397,In_179);
and U242 (N_242,In_409,In_28);
or U243 (N_243,In_330,In_322);
and U244 (N_244,In_341,N_199);
or U245 (N_245,N_114,In_487);
or U246 (N_246,In_470,In_42);
nand U247 (N_247,In_181,In_381);
and U248 (N_248,N_52,N_141);
and U249 (N_249,In_123,In_180);
nand U250 (N_250,In_430,In_468);
nand U251 (N_251,N_117,In_456);
nand U252 (N_252,N_136,In_126);
nor U253 (N_253,N_122,N_218);
and U254 (N_254,N_203,In_321);
or U255 (N_255,In_455,N_234);
or U256 (N_256,N_165,N_180);
nor U257 (N_257,In_184,In_360);
or U258 (N_258,In_192,In_440);
nor U259 (N_259,In_362,N_53);
or U260 (N_260,In_69,N_69);
or U261 (N_261,N_229,N_186);
nor U262 (N_262,N_167,In_292);
nand U263 (N_263,N_104,In_177);
nor U264 (N_264,N_83,In_174);
or U265 (N_265,In_403,In_390);
nand U266 (N_266,In_473,In_185);
nand U267 (N_267,N_166,In_25);
nand U268 (N_268,In_255,In_229);
nor U269 (N_269,N_183,N_152);
nor U270 (N_270,N_173,In_211);
nor U271 (N_271,In_436,N_200);
nand U272 (N_272,N_119,N_145);
nor U273 (N_273,In_325,In_352);
nand U274 (N_274,In_377,In_110);
nor U275 (N_275,In_58,In_24);
or U276 (N_276,N_111,N_9);
nand U277 (N_277,In_477,In_44);
nand U278 (N_278,N_101,N_196);
or U279 (N_279,In_83,N_215);
or U280 (N_280,N_59,N_216);
and U281 (N_281,N_162,N_86);
or U282 (N_282,N_155,In_438);
or U283 (N_283,N_112,N_147);
nand U284 (N_284,N_149,In_291);
or U285 (N_285,N_56,N_192);
nand U286 (N_286,N_71,In_43);
xor U287 (N_287,In_199,In_109);
or U288 (N_288,N_225,N_130);
nor U289 (N_289,N_17,In_353);
nor U290 (N_290,N_124,In_70);
nor U291 (N_291,N_230,N_187);
nand U292 (N_292,In_71,In_84);
and U293 (N_293,N_159,In_156);
or U294 (N_294,N_74,In_461);
nor U295 (N_295,In_368,N_219);
nor U296 (N_296,N_140,N_61);
or U297 (N_297,N_172,N_137);
nor U298 (N_298,In_378,N_171);
or U299 (N_299,In_392,In_419);
and U300 (N_300,N_191,N_31);
nand U301 (N_301,N_174,In_285);
or U302 (N_302,In_91,N_222);
or U303 (N_303,N_290,N_261);
and U304 (N_304,N_280,N_132);
and U305 (N_305,N_213,N_91);
nor U306 (N_306,In_280,N_244);
xnor U307 (N_307,N_193,In_406);
nor U308 (N_308,In_444,N_247);
or U309 (N_309,N_241,In_386);
or U310 (N_310,In_86,In_29);
or U311 (N_311,N_269,In_302);
and U312 (N_312,N_209,N_270);
and U313 (N_313,N_291,N_239);
and U314 (N_314,N_224,N_297);
or U315 (N_315,N_275,N_32);
and U316 (N_316,N_235,N_100);
and U317 (N_317,N_214,N_121);
or U318 (N_318,N_267,In_435);
nor U319 (N_319,N_282,N_233);
or U320 (N_320,N_63,N_177);
or U321 (N_321,N_246,In_488);
nand U322 (N_322,In_37,N_266);
nor U323 (N_323,N_255,N_133);
nand U324 (N_324,N_197,In_426);
nand U325 (N_325,N_257,N_201);
nor U326 (N_326,N_236,N_208);
and U327 (N_327,N_288,N_207);
nand U328 (N_328,N_154,In_337);
and U329 (N_329,N_55,N_245);
or U330 (N_330,N_271,N_293);
nand U331 (N_331,N_158,In_233);
nor U332 (N_332,N_108,N_227);
nor U333 (N_333,N_262,N_252);
nand U334 (N_334,In_393,N_260);
and U335 (N_335,N_283,In_218);
xnor U336 (N_336,N_204,N_277);
and U337 (N_337,N_168,N_221);
xnor U338 (N_338,N_294,N_170);
nand U339 (N_339,N_268,N_202);
nand U340 (N_340,N_75,N_182);
nand U341 (N_341,N_163,N_89);
nand U342 (N_342,N_256,N_286);
or U343 (N_343,In_307,In_64);
and U344 (N_344,N_237,In_137);
or U345 (N_345,N_273,In_82);
nor U346 (N_346,N_279,N_48);
nor U347 (N_347,In_242,In_239);
nor U348 (N_348,N_287,N_3);
nor U349 (N_349,In_241,In_55);
or U350 (N_350,N_110,In_404);
nand U351 (N_351,N_295,N_62);
and U352 (N_352,In_400,N_264);
nor U353 (N_353,N_339,N_242);
and U354 (N_354,In_146,In_338);
nor U355 (N_355,N_116,In_466);
nor U356 (N_356,N_329,In_457);
nor U357 (N_357,N_217,N_198);
and U358 (N_358,N_254,N_231);
nor U359 (N_359,N_300,N_332);
or U360 (N_360,In_191,N_194);
or U361 (N_361,N_314,N_211);
nand U362 (N_362,In_439,N_82);
nand U363 (N_363,N_299,N_176);
nand U364 (N_364,In_249,N_106);
nand U365 (N_365,N_220,N_210);
nor U366 (N_366,N_309,In_169);
and U367 (N_367,In_15,N_301);
or U368 (N_368,N_324,N_42);
or U369 (N_369,N_205,N_305);
or U370 (N_370,N_325,In_295);
and U371 (N_371,N_212,In_414);
and U372 (N_372,In_309,N_310);
and U373 (N_373,N_326,In_144);
and U374 (N_374,N_337,N_330);
and U375 (N_375,N_265,N_40);
and U376 (N_376,N_347,N_334);
or U377 (N_377,N_327,N_302);
nor U378 (N_378,In_85,N_321);
or U379 (N_379,N_272,In_374);
or U380 (N_380,N_281,N_331);
or U381 (N_381,N_296,N_344);
nor U382 (N_382,N_328,N_343);
nor U383 (N_383,N_248,N_4);
and U384 (N_384,N_274,In_251);
or U385 (N_385,N_316,N_232);
or U386 (N_386,N_151,N_51);
and U387 (N_387,In_296,N_251);
and U388 (N_388,N_276,N_284);
nor U389 (N_389,N_311,In_149);
and U390 (N_390,N_258,N_146);
or U391 (N_391,N_206,N_303);
or U392 (N_392,N_1,In_284);
or U393 (N_393,N_228,N_99);
nand U394 (N_394,N_313,N_307);
or U395 (N_395,N_278,N_58);
and U396 (N_396,N_84,N_19);
nand U397 (N_397,N_138,N_95);
nor U398 (N_398,N_240,In_327);
or U399 (N_399,N_322,In_254);
or U400 (N_400,N_263,N_351);
nand U401 (N_401,N_226,In_265);
and U402 (N_402,N_346,N_366);
nand U403 (N_403,N_238,N_398);
nand U404 (N_404,N_259,In_76);
and U405 (N_405,N_250,N_285);
and U406 (N_406,N_249,N_380);
and U407 (N_407,N_350,N_298);
nand U408 (N_408,N_253,N_185);
and U409 (N_409,In_276,N_368);
and U410 (N_410,N_394,N_317);
and U411 (N_411,N_320,N_359);
nor U412 (N_412,N_354,N_361);
nand U413 (N_413,N_312,N_181);
nor U414 (N_414,In_51,N_388);
nor U415 (N_415,N_397,N_349);
nand U416 (N_416,N_352,N_382);
or U417 (N_417,N_336,N_243);
or U418 (N_418,N_304,N_384);
nand U419 (N_419,N_348,N_355);
and U420 (N_420,N_371,N_333);
nor U421 (N_421,N_338,N_399);
and U422 (N_422,N_134,N_393);
or U423 (N_423,N_292,N_395);
nor U424 (N_424,N_315,N_340);
nand U425 (N_425,N_376,N_107);
nor U426 (N_426,N_365,N_385);
nand U427 (N_427,In_270,N_386);
nor U428 (N_428,N_345,N_367);
or U429 (N_429,N_306,N_364);
nand U430 (N_430,N_381,N_391);
nor U431 (N_431,N_392,N_375);
and U432 (N_432,In_405,N_378);
nor U433 (N_433,N_342,N_341);
and U434 (N_434,N_289,N_223);
or U435 (N_435,N_362,N_109);
or U436 (N_436,N_118,N_369);
or U437 (N_437,N_396,N_377);
and U438 (N_438,N_373,N_387);
nand U439 (N_439,N_390,N_318);
and U440 (N_440,N_308,N_370);
nor U441 (N_441,In_410,N_356);
or U442 (N_442,N_335,N_319);
or U443 (N_443,N_96,N_374);
and U444 (N_444,N_389,N_363);
or U445 (N_445,N_383,N_358);
and U446 (N_446,In_328,N_372);
nor U447 (N_447,N_16,N_323);
nand U448 (N_448,N_360,N_357);
nand U449 (N_449,N_379,N_353);
and U450 (N_450,N_429,N_412);
nand U451 (N_451,N_436,N_442);
or U452 (N_452,N_417,N_425);
or U453 (N_453,N_441,N_431);
nand U454 (N_454,N_440,N_400);
nor U455 (N_455,N_439,N_437);
nor U456 (N_456,N_401,N_408);
and U457 (N_457,N_420,N_423);
or U458 (N_458,N_402,N_426);
nor U459 (N_459,N_413,N_410);
nor U460 (N_460,N_418,N_422);
nand U461 (N_461,N_415,N_430);
nand U462 (N_462,N_432,N_406);
nor U463 (N_463,N_421,N_435);
nor U464 (N_464,N_405,N_447);
nor U465 (N_465,N_419,N_434);
nand U466 (N_466,N_414,N_411);
nand U467 (N_467,N_403,N_428);
or U468 (N_468,N_445,N_449);
and U469 (N_469,N_438,N_424);
nand U470 (N_470,N_427,N_433);
nand U471 (N_471,N_407,N_446);
xnor U472 (N_472,N_444,N_416);
nor U473 (N_473,N_448,N_404);
or U474 (N_474,N_443,N_409);
nand U475 (N_475,N_433,N_430);
and U476 (N_476,N_417,N_400);
or U477 (N_477,N_438,N_428);
nor U478 (N_478,N_419,N_449);
or U479 (N_479,N_435,N_446);
nor U480 (N_480,N_444,N_437);
and U481 (N_481,N_429,N_400);
and U482 (N_482,N_419,N_410);
and U483 (N_483,N_407,N_417);
nand U484 (N_484,N_418,N_417);
and U485 (N_485,N_422,N_404);
nand U486 (N_486,N_428,N_445);
or U487 (N_487,N_428,N_419);
and U488 (N_488,N_444,N_420);
nand U489 (N_489,N_408,N_402);
nor U490 (N_490,N_439,N_443);
and U491 (N_491,N_435,N_415);
xor U492 (N_492,N_428,N_441);
and U493 (N_493,N_441,N_444);
or U494 (N_494,N_426,N_429);
nand U495 (N_495,N_425,N_413);
or U496 (N_496,N_420,N_447);
nand U497 (N_497,N_442,N_438);
and U498 (N_498,N_437,N_423);
nand U499 (N_499,N_417,N_429);
nor U500 (N_500,N_463,N_470);
nor U501 (N_501,N_497,N_461);
and U502 (N_502,N_462,N_465);
or U503 (N_503,N_475,N_498);
and U504 (N_504,N_469,N_473);
nand U505 (N_505,N_482,N_471);
or U506 (N_506,N_492,N_456);
and U507 (N_507,N_457,N_499);
nor U508 (N_508,N_452,N_484);
or U509 (N_509,N_478,N_455);
and U510 (N_510,N_458,N_468);
nor U511 (N_511,N_464,N_487);
nor U512 (N_512,N_496,N_494);
nand U513 (N_513,N_459,N_486);
nand U514 (N_514,N_476,N_474);
or U515 (N_515,N_454,N_466);
nand U516 (N_516,N_493,N_483);
nand U517 (N_517,N_495,N_467);
nor U518 (N_518,N_488,N_480);
nand U519 (N_519,N_451,N_490);
nor U520 (N_520,N_485,N_477);
or U521 (N_521,N_481,N_472);
and U522 (N_522,N_460,N_489);
nor U523 (N_523,N_479,N_450);
or U524 (N_524,N_491,N_453);
nand U525 (N_525,N_488,N_459);
nor U526 (N_526,N_477,N_481);
nand U527 (N_527,N_470,N_457);
nand U528 (N_528,N_453,N_482);
nor U529 (N_529,N_475,N_495);
nand U530 (N_530,N_463,N_456);
nor U531 (N_531,N_492,N_452);
and U532 (N_532,N_458,N_481);
and U533 (N_533,N_492,N_459);
or U534 (N_534,N_459,N_476);
nor U535 (N_535,N_452,N_458);
nor U536 (N_536,N_490,N_494);
nand U537 (N_537,N_472,N_453);
nand U538 (N_538,N_469,N_493);
nand U539 (N_539,N_470,N_479);
and U540 (N_540,N_475,N_488);
and U541 (N_541,N_492,N_489);
nand U542 (N_542,N_479,N_484);
or U543 (N_543,N_478,N_495);
nor U544 (N_544,N_463,N_496);
nand U545 (N_545,N_481,N_455);
or U546 (N_546,N_470,N_494);
or U547 (N_547,N_461,N_494);
or U548 (N_548,N_496,N_470);
and U549 (N_549,N_498,N_462);
or U550 (N_550,N_532,N_505);
nor U551 (N_551,N_533,N_530);
and U552 (N_552,N_500,N_518);
nor U553 (N_553,N_542,N_506);
nor U554 (N_554,N_538,N_521);
nor U555 (N_555,N_548,N_549);
nor U556 (N_556,N_509,N_504);
or U557 (N_557,N_529,N_525);
nor U558 (N_558,N_526,N_516);
nand U559 (N_559,N_540,N_515);
nand U560 (N_560,N_511,N_517);
nor U561 (N_561,N_536,N_531);
or U562 (N_562,N_543,N_545);
or U563 (N_563,N_512,N_522);
and U564 (N_564,N_546,N_523);
nor U565 (N_565,N_547,N_501);
or U566 (N_566,N_507,N_519);
or U567 (N_567,N_528,N_524);
nor U568 (N_568,N_544,N_535);
and U569 (N_569,N_502,N_503);
and U570 (N_570,N_508,N_537);
and U571 (N_571,N_514,N_510);
and U572 (N_572,N_520,N_534);
and U573 (N_573,N_541,N_527);
nand U574 (N_574,N_513,N_539);
and U575 (N_575,N_544,N_504);
and U576 (N_576,N_515,N_530);
nor U577 (N_577,N_536,N_548);
nor U578 (N_578,N_530,N_540);
and U579 (N_579,N_532,N_519);
nand U580 (N_580,N_509,N_518);
or U581 (N_581,N_511,N_503);
nand U582 (N_582,N_549,N_525);
nand U583 (N_583,N_540,N_534);
and U584 (N_584,N_520,N_509);
and U585 (N_585,N_510,N_512);
or U586 (N_586,N_501,N_506);
and U587 (N_587,N_541,N_522);
or U588 (N_588,N_536,N_547);
nor U589 (N_589,N_503,N_519);
nand U590 (N_590,N_525,N_540);
or U591 (N_591,N_500,N_543);
nor U592 (N_592,N_518,N_545);
nor U593 (N_593,N_527,N_549);
and U594 (N_594,N_512,N_504);
nand U595 (N_595,N_531,N_532);
and U596 (N_596,N_522,N_516);
or U597 (N_597,N_536,N_538);
or U598 (N_598,N_541,N_512);
or U599 (N_599,N_543,N_509);
and U600 (N_600,N_563,N_562);
or U601 (N_601,N_597,N_555);
or U602 (N_602,N_581,N_586);
and U603 (N_603,N_572,N_587);
and U604 (N_604,N_594,N_599);
nor U605 (N_605,N_579,N_591);
and U606 (N_606,N_560,N_576);
and U607 (N_607,N_593,N_577);
or U608 (N_608,N_583,N_559);
and U609 (N_609,N_575,N_565);
or U610 (N_610,N_588,N_584);
nand U611 (N_611,N_589,N_558);
and U612 (N_612,N_551,N_557);
or U613 (N_613,N_552,N_569);
or U614 (N_614,N_556,N_568);
nor U615 (N_615,N_561,N_580);
and U616 (N_616,N_585,N_567);
nor U617 (N_617,N_570,N_550);
nor U618 (N_618,N_553,N_592);
nand U619 (N_619,N_564,N_598);
and U620 (N_620,N_595,N_578);
nand U621 (N_621,N_590,N_596);
and U622 (N_622,N_571,N_573);
nand U623 (N_623,N_574,N_582);
and U624 (N_624,N_554,N_566);
xor U625 (N_625,N_558,N_561);
nor U626 (N_626,N_594,N_592);
or U627 (N_627,N_597,N_581);
and U628 (N_628,N_551,N_567);
nor U629 (N_629,N_554,N_596);
and U630 (N_630,N_562,N_564);
and U631 (N_631,N_583,N_575);
and U632 (N_632,N_587,N_555);
or U633 (N_633,N_571,N_563);
nor U634 (N_634,N_579,N_558);
nand U635 (N_635,N_573,N_599);
nor U636 (N_636,N_560,N_565);
or U637 (N_637,N_586,N_562);
nand U638 (N_638,N_580,N_565);
nand U639 (N_639,N_582,N_598);
nand U640 (N_640,N_599,N_596);
nand U641 (N_641,N_564,N_570);
and U642 (N_642,N_582,N_595);
and U643 (N_643,N_554,N_597);
nand U644 (N_644,N_594,N_579);
or U645 (N_645,N_560,N_579);
nor U646 (N_646,N_568,N_565);
nand U647 (N_647,N_587,N_582);
nor U648 (N_648,N_561,N_555);
or U649 (N_649,N_579,N_575);
nor U650 (N_650,N_648,N_612);
nor U651 (N_651,N_625,N_642);
nand U652 (N_652,N_640,N_611);
or U653 (N_653,N_619,N_614);
or U654 (N_654,N_638,N_645);
and U655 (N_655,N_604,N_606);
nand U656 (N_656,N_644,N_618);
or U657 (N_657,N_610,N_627);
nand U658 (N_658,N_620,N_649);
nor U659 (N_659,N_635,N_631);
nor U660 (N_660,N_639,N_628);
nand U661 (N_661,N_646,N_623);
nor U662 (N_662,N_624,N_617);
nor U663 (N_663,N_615,N_643);
nand U664 (N_664,N_630,N_641);
and U665 (N_665,N_636,N_613);
or U666 (N_666,N_601,N_607);
or U667 (N_667,N_621,N_632);
and U668 (N_668,N_647,N_616);
nor U669 (N_669,N_605,N_603);
nor U670 (N_670,N_602,N_600);
or U671 (N_671,N_626,N_633);
nor U672 (N_672,N_629,N_637);
nor U673 (N_673,N_622,N_634);
or U674 (N_674,N_609,N_608);
nor U675 (N_675,N_628,N_602);
nor U676 (N_676,N_601,N_632);
nand U677 (N_677,N_603,N_613);
and U678 (N_678,N_639,N_627);
nor U679 (N_679,N_615,N_602);
or U680 (N_680,N_611,N_624);
and U681 (N_681,N_600,N_641);
nand U682 (N_682,N_640,N_620);
or U683 (N_683,N_616,N_622);
nor U684 (N_684,N_629,N_615);
or U685 (N_685,N_619,N_642);
xnor U686 (N_686,N_611,N_614);
or U687 (N_687,N_639,N_600);
nand U688 (N_688,N_602,N_627);
nand U689 (N_689,N_614,N_625);
nor U690 (N_690,N_646,N_638);
or U691 (N_691,N_643,N_600);
or U692 (N_692,N_627,N_601);
or U693 (N_693,N_621,N_615);
and U694 (N_694,N_627,N_613);
nor U695 (N_695,N_607,N_624);
nand U696 (N_696,N_612,N_641);
nand U697 (N_697,N_606,N_610);
and U698 (N_698,N_637,N_604);
and U699 (N_699,N_630,N_614);
nor U700 (N_700,N_679,N_676);
nor U701 (N_701,N_696,N_673);
nand U702 (N_702,N_681,N_694);
nor U703 (N_703,N_659,N_656);
nor U704 (N_704,N_699,N_698);
nand U705 (N_705,N_680,N_663);
and U706 (N_706,N_690,N_677);
or U707 (N_707,N_685,N_671);
nand U708 (N_708,N_684,N_664);
or U709 (N_709,N_666,N_669);
or U710 (N_710,N_674,N_672);
and U711 (N_711,N_655,N_697);
nand U712 (N_712,N_667,N_657);
nand U713 (N_713,N_660,N_683);
or U714 (N_714,N_650,N_692);
and U715 (N_715,N_682,N_661);
or U716 (N_716,N_665,N_662);
nor U717 (N_717,N_689,N_688);
nor U718 (N_718,N_670,N_653);
or U719 (N_719,N_654,N_687);
or U720 (N_720,N_658,N_652);
nand U721 (N_721,N_695,N_678);
nor U722 (N_722,N_668,N_693);
nor U723 (N_723,N_691,N_675);
and U724 (N_724,N_651,N_686);
or U725 (N_725,N_669,N_650);
nor U726 (N_726,N_670,N_685);
and U727 (N_727,N_656,N_675);
or U728 (N_728,N_681,N_651);
nand U729 (N_729,N_683,N_663);
and U730 (N_730,N_667,N_659);
and U731 (N_731,N_668,N_674);
or U732 (N_732,N_691,N_654);
nand U733 (N_733,N_656,N_679);
or U734 (N_734,N_671,N_699);
nand U735 (N_735,N_670,N_681);
nor U736 (N_736,N_661,N_664);
and U737 (N_737,N_689,N_661);
nand U738 (N_738,N_672,N_656);
nor U739 (N_739,N_695,N_698);
nand U740 (N_740,N_650,N_699);
nand U741 (N_741,N_676,N_689);
and U742 (N_742,N_672,N_682);
and U743 (N_743,N_668,N_672);
or U744 (N_744,N_671,N_656);
nor U745 (N_745,N_651,N_684);
and U746 (N_746,N_698,N_676);
nor U747 (N_747,N_690,N_667);
or U748 (N_748,N_688,N_694);
nand U749 (N_749,N_699,N_673);
nand U750 (N_750,N_704,N_703);
nor U751 (N_751,N_735,N_749);
nand U752 (N_752,N_714,N_729);
nand U753 (N_753,N_744,N_731);
and U754 (N_754,N_726,N_705);
nand U755 (N_755,N_728,N_722);
nand U756 (N_756,N_727,N_708);
or U757 (N_757,N_713,N_742);
or U758 (N_758,N_740,N_721);
xor U759 (N_759,N_730,N_711);
and U760 (N_760,N_743,N_736);
and U761 (N_761,N_725,N_700);
and U762 (N_762,N_718,N_702);
nand U763 (N_763,N_738,N_739);
nor U764 (N_764,N_715,N_710);
and U765 (N_765,N_707,N_723);
nor U766 (N_766,N_720,N_745);
nand U767 (N_767,N_737,N_701);
nor U768 (N_768,N_712,N_706);
or U769 (N_769,N_747,N_732);
and U770 (N_770,N_746,N_717);
and U771 (N_771,N_733,N_748);
nand U772 (N_772,N_719,N_724);
nor U773 (N_773,N_734,N_709);
and U774 (N_774,N_716,N_741);
and U775 (N_775,N_736,N_731);
or U776 (N_776,N_740,N_719);
nand U777 (N_777,N_741,N_707);
and U778 (N_778,N_722,N_737);
or U779 (N_779,N_736,N_727);
nor U780 (N_780,N_722,N_730);
and U781 (N_781,N_713,N_707);
and U782 (N_782,N_719,N_739);
nand U783 (N_783,N_736,N_719);
nor U784 (N_784,N_746,N_704);
or U785 (N_785,N_700,N_732);
and U786 (N_786,N_732,N_742);
nand U787 (N_787,N_707,N_725);
nand U788 (N_788,N_742,N_749);
or U789 (N_789,N_738,N_737);
nor U790 (N_790,N_705,N_748);
nor U791 (N_791,N_747,N_700);
or U792 (N_792,N_707,N_738);
or U793 (N_793,N_748,N_745);
xor U794 (N_794,N_709,N_730);
or U795 (N_795,N_708,N_738);
nor U796 (N_796,N_747,N_701);
nor U797 (N_797,N_713,N_711);
nor U798 (N_798,N_746,N_705);
nor U799 (N_799,N_702,N_739);
nor U800 (N_800,N_781,N_765);
and U801 (N_801,N_784,N_771);
nand U802 (N_802,N_768,N_783);
or U803 (N_803,N_756,N_762);
nor U804 (N_804,N_791,N_757);
nor U805 (N_805,N_775,N_773);
nor U806 (N_806,N_787,N_761);
nand U807 (N_807,N_777,N_792);
nand U808 (N_808,N_795,N_798);
nor U809 (N_809,N_780,N_785);
nor U810 (N_810,N_755,N_799);
or U811 (N_811,N_774,N_789);
nor U812 (N_812,N_760,N_793);
nor U813 (N_813,N_772,N_794);
and U814 (N_814,N_769,N_790);
nor U815 (N_815,N_754,N_764);
nor U816 (N_816,N_796,N_788);
nand U817 (N_817,N_770,N_797);
nand U818 (N_818,N_776,N_763);
or U819 (N_819,N_778,N_782);
nand U820 (N_820,N_766,N_759);
nor U821 (N_821,N_750,N_751);
and U822 (N_822,N_752,N_767);
nor U823 (N_823,N_758,N_786);
or U824 (N_824,N_753,N_779);
or U825 (N_825,N_761,N_790);
or U826 (N_826,N_765,N_764);
nor U827 (N_827,N_775,N_785);
and U828 (N_828,N_790,N_797);
nor U829 (N_829,N_773,N_782);
nor U830 (N_830,N_777,N_786);
nand U831 (N_831,N_785,N_773);
and U832 (N_832,N_791,N_756);
nor U833 (N_833,N_759,N_797);
nand U834 (N_834,N_782,N_755);
nand U835 (N_835,N_752,N_786);
and U836 (N_836,N_765,N_784);
or U837 (N_837,N_767,N_769);
nand U838 (N_838,N_765,N_753);
or U839 (N_839,N_758,N_776);
or U840 (N_840,N_787,N_755);
or U841 (N_841,N_775,N_784);
and U842 (N_842,N_777,N_764);
and U843 (N_843,N_798,N_766);
nand U844 (N_844,N_771,N_767);
nand U845 (N_845,N_759,N_778);
nand U846 (N_846,N_765,N_750);
nor U847 (N_847,N_787,N_779);
nor U848 (N_848,N_753,N_754);
nand U849 (N_849,N_765,N_756);
or U850 (N_850,N_849,N_830);
nor U851 (N_851,N_817,N_811);
nand U852 (N_852,N_827,N_803);
and U853 (N_853,N_846,N_820);
nand U854 (N_854,N_814,N_819);
and U855 (N_855,N_848,N_804);
or U856 (N_856,N_826,N_847);
and U857 (N_857,N_809,N_834);
nor U858 (N_858,N_822,N_838);
or U859 (N_859,N_840,N_824);
nand U860 (N_860,N_828,N_815);
or U861 (N_861,N_807,N_831);
or U862 (N_862,N_802,N_813);
or U863 (N_863,N_812,N_821);
nor U864 (N_864,N_825,N_829);
nand U865 (N_865,N_816,N_845);
nor U866 (N_866,N_810,N_805);
and U867 (N_867,N_818,N_800);
nand U868 (N_868,N_832,N_839);
and U869 (N_869,N_823,N_808);
nand U870 (N_870,N_806,N_835);
nand U871 (N_871,N_842,N_843);
nor U872 (N_872,N_844,N_841);
nor U873 (N_873,N_837,N_836);
nand U874 (N_874,N_801,N_833);
nor U875 (N_875,N_834,N_826);
nand U876 (N_876,N_818,N_838);
nor U877 (N_877,N_827,N_837);
and U878 (N_878,N_800,N_817);
and U879 (N_879,N_843,N_837);
nand U880 (N_880,N_801,N_846);
nor U881 (N_881,N_811,N_841);
and U882 (N_882,N_803,N_843);
and U883 (N_883,N_828,N_832);
and U884 (N_884,N_823,N_805);
or U885 (N_885,N_843,N_826);
nand U886 (N_886,N_841,N_837);
and U887 (N_887,N_819,N_847);
and U888 (N_888,N_806,N_800);
and U889 (N_889,N_837,N_801);
nor U890 (N_890,N_820,N_849);
and U891 (N_891,N_819,N_808);
or U892 (N_892,N_828,N_847);
nand U893 (N_893,N_827,N_832);
or U894 (N_894,N_837,N_842);
nand U895 (N_895,N_823,N_804);
and U896 (N_896,N_823,N_835);
nor U897 (N_897,N_836,N_806);
nor U898 (N_898,N_843,N_805);
xnor U899 (N_899,N_808,N_814);
or U900 (N_900,N_862,N_883);
or U901 (N_901,N_876,N_892);
or U902 (N_902,N_887,N_874);
nor U903 (N_903,N_872,N_891);
xor U904 (N_904,N_857,N_866);
or U905 (N_905,N_869,N_880);
or U906 (N_906,N_860,N_850);
or U907 (N_907,N_863,N_884);
nor U908 (N_908,N_853,N_865);
or U909 (N_909,N_898,N_897);
nor U910 (N_910,N_871,N_890);
nor U911 (N_911,N_864,N_877);
and U912 (N_912,N_859,N_894);
nor U913 (N_913,N_870,N_854);
or U914 (N_914,N_895,N_893);
and U915 (N_915,N_881,N_899);
and U916 (N_916,N_875,N_855);
or U917 (N_917,N_886,N_868);
nor U918 (N_918,N_885,N_867);
nand U919 (N_919,N_856,N_888);
nand U920 (N_920,N_861,N_896);
or U921 (N_921,N_889,N_878);
nand U922 (N_922,N_873,N_879);
nand U923 (N_923,N_852,N_851);
or U924 (N_924,N_882,N_858);
nand U925 (N_925,N_889,N_873);
nor U926 (N_926,N_879,N_891);
or U927 (N_927,N_879,N_870);
nand U928 (N_928,N_865,N_878);
nor U929 (N_929,N_874,N_854);
nor U930 (N_930,N_861,N_899);
or U931 (N_931,N_858,N_884);
and U932 (N_932,N_869,N_850);
nand U933 (N_933,N_879,N_859);
nand U934 (N_934,N_863,N_894);
nand U935 (N_935,N_886,N_856);
nor U936 (N_936,N_874,N_856);
nand U937 (N_937,N_898,N_899);
nand U938 (N_938,N_853,N_884);
and U939 (N_939,N_860,N_891);
nor U940 (N_940,N_871,N_889);
or U941 (N_941,N_867,N_853);
and U942 (N_942,N_859,N_868);
and U943 (N_943,N_862,N_877);
and U944 (N_944,N_871,N_884);
nand U945 (N_945,N_886,N_861);
nor U946 (N_946,N_858,N_875);
nand U947 (N_947,N_884,N_888);
nor U948 (N_948,N_887,N_858);
nand U949 (N_949,N_885,N_893);
nor U950 (N_950,N_920,N_942);
or U951 (N_951,N_912,N_921);
nand U952 (N_952,N_929,N_947);
nand U953 (N_953,N_923,N_946);
nand U954 (N_954,N_924,N_900);
or U955 (N_955,N_925,N_905);
and U956 (N_956,N_939,N_903);
nand U957 (N_957,N_915,N_932);
nand U958 (N_958,N_904,N_928);
and U959 (N_959,N_909,N_944);
and U960 (N_960,N_913,N_926);
nor U961 (N_961,N_930,N_937);
nor U962 (N_962,N_917,N_919);
nand U963 (N_963,N_922,N_906);
nor U964 (N_964,N_948,N_911);
nand U965 (N_965,N_933,N_941);
or U966 (N_966,N_916,N_943);
nand U967 (N_967,N_908,N_914);
or U968 (N_968,N_935,N_918);
nor U969 (N_969,N_927,N_936);
nor U970 (N_970,N_931,N_902);
and U971 (N_971,N_934,N_907);
or U972 (N_972,N_910,N_940);
nor U973 (N_973,N_949,N_938);
nand U974 (N_974,N_945,N_901);
and U975 (N_975,N_923,N_928);
nand U976 (N_976,N_923,N_911);
or U977 (N_977,N_909,N_918);
nor U978 (N_978,N_917,N_947);
nor U979 (N_979,N_917,N_930);
and U980 (N_980,N_927,N_900);
or U981 (N_981,N_913,N_917);
nand U982 (N_982,N_940,N_934);
or U983 (N_983,N_936,N_910);
or U984 (N_984,N_907,N_903);
nor U985 (N_985,N_949,N_939);
or U986 (N_986,N_913,N_905);
nor U987 (N_987,N_912,N_943);
nor U988 (N_988,N_944,N_920);
xnor U989 (N_989,N_934,N_930);
nand U990 (N_990,N_903,N_922);
nor U991 (N_991,N_911,N_941);
and U992 (N_992,N_934,N_947);
nand U993 (N_993,N_901,N_924);
xor U994 (N_994,N_938,N_921);
or U995 (N_995,N_908,N_919);
and U996 (N_996,N_924,N_911);
nand U997 (N_997,N_931,N_947);
nor U998 (N_998,N_911,N_903);
or U999 (N_999,N_930,N_926);
nor U1000 (N_1000,N_989,N_965);
or U1001 (N_1001,N_973,N_955);
and U1002 (N_1002,N_962,N_987);
nor U1003 (N_1003,N_983,N_952);
and U1004 (N_1004,N_999,N_960);
or U1005 (N_1005,N_951,N_996);
nor U1006 (N_1006,N_967,N_975);
nand U1007 (N_1007,N_997,N_974);
and U1008 (N_1008,N_990,N_971);
nor U1009 (N_1009,N_972,N_995);
and U1010 (N_1010,N_982,N_963);
nand U1011 (N_1011,N_966,N_980);
or U1012 (N_1012,N_977,N_969);
and U1013 (N_1013,N_970,N_986);
nand U1014 (N_1014,N_959,N_954);
and U1015 (N_1015,N_998,N_991);
nand U1016 (N_1016,N_950,N_979);
or U1017 (N_1017,N_976,N_978);
and U1018 (N_1018,N_985,N_994);
and U1019 (N_1019,N_984,N_988);
nor U1020 (N_1020,N_964,N_993);
nand U1021 (N_1021,N_981,N_953);
nor U1022 (N_1022,N_956,N_958);
or U1023 (N_1023,N_957,N_968);
nand U1024 (N_1024,N_992,N_961);
and U1025 (N_1025,N_970,N_971);
or U1026 (N_1026,N_995,N_991);
nand U1027 (N_1027,N_994,N_990);
or U1028 (N_1028,N_981,N_952);
and U1029 (N_1029,N_984,N_963);
and U1030 (N_1030,N_983,N_994);
and U1031 (N_1031,N_995,N_961);
or U1032 (N_1032,N_956,N_992);
and U1033 (N_1033,N_960,N_967);
nand U1034 (N_1034,N_990,N_987);
nor U1035 (N_1035,N_980,N_987);
nand U1036 (N_1036,N_972,N_990);
nor U1037 (N_1037,N_960,N_952);
nor U1038 (N_1038,N_960,N_998);
and U1039 (N_1039,N_961,N_988);
nand U1040 (N_1040,N_993,N_962);
nand U1041 (N_1041,N_963,N_960);
nor U1042 (N_1042,N_960,N_982);
nor U1043 (N_1043,N_984,N_999);
or U1044 (N_1044,N_982,N_978);
and U1045 (N_1045,N_963,N_988);
nor U1046 (N_1046,N_994,N_993);
nor U1047 (N_1047,N_954,N_965);
or U1048 (N_1048,N_989,N_963);
or U1049 (N_1049,N_970,N_964);
nand U1050 (N_1050,N_1012,N_1026);
or U1051 (N_1051,N_1000,N_1034);
and U1052 (N_1052,N_1031,N_1039);
nand U1053 (N_1053,N_1035,N_1023);
nand U1054 (N_1054,N_1042,N_1048);
or U1055 (N_1055,N_1019,N_1003);
and U1056 (N_1056,N_1014,N_1027);
and U1057 (N_1057,N_1025,N_1028);
and U1058 (N_1058,N_1001,N_1040);
and U1059 (N_1059,N_1022,N_1024);
nor U1060 (N_1060,N_1002,N_1013);
xnor U1061 (N_1061,N_1009,N_1037);
and U1062 (N_1062,N_1016,N_1021);
nor U1063 (N_1063,N_1045,N_1043);
xnor U1064 (N_1064,N_1038,N_1047);
nand U1065 (N_1065,N_1030,N_1007);
or U1066 (N_1066,N_1010,N_1044);
nor U1067 (N_1067,N_1033,N_1005);
or U1068 (N_1068,N_1029,N_1020);
or U1069 (N_1069,N_1011,N_1008);
or U1070 (N_1070,N_1018,N_1006);
nor U1071 (N_1071,N_1017,N_1046);
or U1072 (N_1072,N_1049,N_1015);
nor U1073 (N_1073,N_1041,N_1032);
and U1074 (N_1074,N_1036,N_1004);
and U1075 (N_1075,N_1048,N_1023);
nand U1076 (N_1076,N_1042,N_1032);
nor U1077 (N_1077,N_1045,N_1017);
nor U1078 (N_1078,N_1018,N_1013);
xor U1079 (N_1079,N_1041,N_1047);
or U1080 (N_1080,N_1049,N_1000);
and U1081 (N_1081,N_1006,N_1027);
and U1082 (N_1082,N_1011,N_1019);
nor U1083 (N_1083,N_1003,N_1013);
nand U1084 (N_1084,N_1010,N_1028);
nand U1085 (N_1085,N_1036,N_1010);
nand U1086 (N_1086,N_1009,N_1032);
or U1087 (N_1087,N_1021,N_1047);
and U1088 (N_1088,N_1041,N_1011);
or U1089 (N_1089,N_1045,N_1004);
nor U1090 (N_1090,N_1041,N_1044);
nand U1091 (N_1091,N_1004,N_1040);
nand U1092 (N_1092,N_1035,N_1036);
or U1093 (N_1093,N_1023,N_1044);
nand U1094 (N_1094,N_1041,N_1026);
and U1095 (N_1095,N_1036,N_1018);
nor U1096 (N_1096,N_1026,N_1016);
nand U1097 (N_1097,N_1026,N_1040);
nand U1098 (N_1098,N_1021,N_1018);
or U1099 (N_1099,N_1016,N_1013);
nor U1100 (N_1100,N_1072,N_1094);
or U1101 (N_1101,N_1098,N_1089);
or U1102 (N_1102,N_1059,N_1063);
or U1103 (N_1103,N_1079,N_1084);
nor U1104 (N_1104,N_1093,N_1057);
nor U1105 (N_1105,N_1076,N_1086);
nor U1106 (N_1106,N_1051,N_1090);
nand U1107 (N_1107,N_1065,N_1077);
and U1108 (N_1108,N_1099,N_1062);
or U1109 (N_1109,N_1081,N_1087);
nor U1110 (N_1110,N_1083,N_1092);
or U1111 (N_1111,N_1056,N_1095);
nor U1112 (N_1112,N_1069,N_1067);
and U1113 (N_1113,N_1064,N_1080);
nand U1114 (N_1114,N_1068,N_1075);
nand U1115 (N_1115,N_1066,N_1053);
and U1116 (N_1116,N_1071,N_1085);
and U1117 (N_1117,N_1058,N_1060);
and U1118 (N_1118,N_1050,N_1088);
nor U1119 (N_1119,N_1055,N_1091);
nor U1120 (N_1120,N_1078,N_1052);
and U1121 (N_1121,N_1096,N_1082);
nor U1122 (N_1122,N_1074,N_1070);
and U1123 (N_1123,N_1073,N_1061);
nor U1124 (N_1124,N_1054,N_1097);
or U1125 (N_1125,N_1053,N_1098);
or U1126 (N_1126,N_1089,N_1068);
nor U1127 (N_1127,N_1060,N_1096);
xnor U1128 (N_1128,N_1055,N_1054);
nand U1129 (N_1129,N_1077,N_1070);
nor U1130 (N_1130,N_1089,N_1073);
and U1131 (N_1131,N_1078,N_1073);
or U1132 (N_1132,N_1092,N_1091);
nand U1133 (N_1133,N_1094,N_1086);
nand U1134 (N_1134,N_1095,N_1074);
nor U1135 (N_1135,N_1056,N_1079);
and U1136 (N_1136,N_1075,N_1073);
nand U1137 (N_1137,N_1061,N_1085);
nor U1138 (N_1138,N_1098,N_1063);
or U1139 (N_1139,N_1082,N_1099);
nor U1140 (N_1140,N_1094,N_1067);
or U1141 (N_1141,N_1078,N_1057);
or U1142 (N_1142,N_1074,N_1061);
nand U1143 (N_1143,N_1088,N_1092);
and U1144 (N_1144,N_1052,N_1054);
and U1145 (N_1145,N_1060,N_1099);
or U1146 (N_1146,N_1063,N_1083);
nor U1147 (N_1147,N_1078,N_1063);
or U1148 (N_1148,N_1058,N_1084);
nor U1149 (N_1149,N_1056,N_1069);
or U1150 (N_1150,N_1133,N_1140);
nor U1151 (N_1151,N_1112,N_1117);
nor U1152 (N_1152,N_1102,N_1139);
nor U1153 (N_1153,N_1122,N_1123);
and U1154 (N_1154,N_1110,N_1118);
and U1155 (N_1155,N_1111,N_1100);
nand U1156 (N_1156,N_1144,N_1124);
nor U1157 (N_1157,N_1120,N_1137);
or U1158 (N_1158,N_1130,N_1107);
nor U1159 (N_1159,N_1114,N_1146);
nor U1160 (N_1160,N_1142,N_1141);
or U1161 (N_1161,N_1145,N_1129);
xor U1162 (N_1162,N_1113,N_1127);
and U1163 (N_1163,N_1105,N_1128);
or U1164 (N_1164,N_1149,N_1143);
nand U1165 (N_1165,N_1116,N_1131);
nor U1166 (N_1166,N_1148,N_1119);
nand U1167 (N_1167,N_1115,N_1109);
or U1168 (N_1168,N_1135,N_1108);
and U1169 (N_1169,N_1101,N_1136);
or U1170 (N_1170,N_1132,N_1106);
nor U1171 (N_1171,N_1121,N_1138);
and U1172 (N_1172,N_1104,N_1103);
nor U1173 (N_1173,N_1125,N_1126);
nand U1174 (N_1174,N_1147,N_1134);
nand U1175 (N_1175,N_1103,N_1105);
nand U1176 (N_1176,N_1119,N_1101);
nand U1177 (N_1177,N_1129,N_1139);
and U1178 (N_1178,N_1139,N_1120);
and U1179 (N_1179,N_1140,N_1120);
or U1180 (N_1180,N_1135,N_1120);
or U1181 (N_1181,N_1142,N_1119);
nand U1182 (N_1182,N_1130,N_1140);
and U1183 (N_1183,N_1117,N_1149);
or U1184 (N_1184,N_1125,N_1110);
and U1185 (N_1185,N_1105,N_1139);
nor U1186 (N_1186,N_1119,N_1149);
or U1187 (N_1187,N_1141,N_1111);
or U1188 (N_1188,N_1145,N_1113);
or U1189 (N_1189,N_1124,N_1139);
and U1190 (N_1190,N_1118,N_1119);
and U1191 (N_1191,N_1134,N_1132);
nand U1192 (N_1192,N_1120,N_1121);
nor U1193 (N_1193,N_1113,N_1112);
and U1194 (N_1194,N_1140,N_1100);
and U1195 (N_1195,N_1149,N_1135);
nand U1196 (N_1196,N_1107,N_1102);
and U1197 (N_1197,N_1101,N_1128);
or U1198 (N_1198,N_1112,N_1135);
and U1199 (N_1199,N_1149,N_1114);
or U1200 (N_1200,N_1173,N_1196);
and U1201 (N_1201,N_1171,N_1199);
nand U1202 (N_1202,N_1179,N_1165);
nand U1203 (N_1203,N_1194,N_1152);
or U1204 (N_1204,N_1183,N_1177);
nand U1205 (N_1205,N_1158,N_1188);
nand U1206 (N_1206,N_1191,N_1198);
nor U1207 (N_1207,N_1170,N_1189);
or U1208 (N_1208,N_1184,N_1186);
nor U1209 (N_1209,N_1172,N_1175);
and U1210 (N_1210,N_1195,N_1167);
nor U1211 (N_1211,N_1180,N_1185);
nor U1212 (N_1212,N_1190,N_1161);
nand U1213 (N_1213,N_1164,N_1169);
nand U1214 (N_1214,N_1157,N_1166);
nand U1215 (N_1215,N_1176,N_1178);
nor U1216 (N_1216,N_1156,N_1174);
nand U1217 (N_1217,N_1159,N_1162);
or U1218 (N_1218,N_1150,N_1182);
nor U1219 (N_1219,N_1160,N_1151);
nand U1220 (N_1220,N_1155,N_1153);
or U1221 (N_1221,N_1181,N_1197);
nor U1222 (N_1222,N_1192,N_1193);
or U1223 (N_1223,N_1168,N_1163);
nor U1224 (N_1224,N_1154,N_1187);
nor U1225 (N_1225,N_1183,N_1191);
and U1226 (N_1226,N_1151,N_1174);
nand U1227 (N_1227,N_1192,N_1197);
nand U1228 (N_1228,N_1182,N_1179);
nor U1229 (N_1229,N_1184,N_1166);
and U1230 (N_1230,N_1159,N_1179);
or U1231 (N_1231,N_1161,N_1176);
or U1232 (N_1232,N_1185,N_1164);
and U1233 (N_1233,N_1154,N_1196);
or U1234 (N_1234,N_1171,N_1150);
nor U1235 (N_1235,N_1163,N_1186);
nand U1236 (N_1236,N_1180,N_1187);
nor U1237 (N_1237,N_1193,N_1180);
nor U1238 (N_1238,N_1158,N_1176);
nand U1239 (N_1239,N_1168,N_1183);
and U1240 (N_1240,N_1188,N_1197);
or U1241 (N_1241,N_1160,N_1154);
nand U1242 (N_1242,N_1175,N_1150);
nor U1243 (N_1243,N_1155,N_1171);
and U1244 (N_1244,N_1199,N_1167);
nand U1245 (N_1245,N_1166,N_1178);
nand U1246 (N_1246,N_1154,N_1194);
and U1247 (N_1247,N_1156,N_1199);
nand U1248 (N_1248,N_1182,N_1191);
nand U1249 (N_1249,N_1177,N_1161);
nor U1250 (N_1250,N_1213,N_1233);
and U1251 (N_1251,N_1220,N_1245);
nand U1252 (N_1252,N_1222,N_1240);
or U1253 (N_1253,N_1235,N_1225);
and U1254 (N_1254,N_1218,N_1202);
and U1255 (N_1255,N_1217,N_1223);
xnor U1256 (N_1256,N_1228,N_1234);
and U1257 (N_1257,N_1241,N_1205);
or U1258 (N_1258,N_1243,N_1211);
and U1259 (N_1259,N_1236,N_1229);
nor U1260 (N_1260,N_1237,N_1208);
and U1261 (N_1261,N_1232,N_1200);
or U1262 (N_1262,N_1203,N_1210);
or U1263 (N_1263,N_1247,N_1212);
nor U1264 (N_1264,N_1239,N_1204);
and U1265 (N_1265,N_1216,N_1214);
and U1266 (N_1266,N_1224,N_1219);
nand U1267 (N_1267,N_1226,N_1215);
or U1268 (N_1268,N_1207,N_1238);
or U1269 (N_1269,N_1242,N_1221);
nand U1270 (N_1270,N_1230,N_1249);
nand U1271 (N_1271,N_1244,N_1201);
or U1272 (N_1272,N_1209,N_1231);
nand U1273 (N_1273,N_1248,N_1246);
and U1274 (N_1274,N_1206,N_1227);
nor U1275 (N_1275,N_1227,N_1223);
and U1276 (N_1276,N_1213,N_1200);
and U1277 (N_1277,N_1208,N_1230);
xnor U1278 (N_1278,N_1229,N_1217);
and U1279 (N_1279,N_1206,N_1229);
nand U1280 (N_1280,N_1210,N_1219);
and U1281 (N_1281,N_1210,N_1230);
nor U1282 (N_1282,N_1223,N_1219);
nand U1283 (N_1283,N_1233,N_1218);
nand U1284 (N_1284,N_1221,N_1208);
nor U1285 (N_1285,N_1228,N_1248);
nor U1286 (N_1286,N_1242,N_1219);
nand U1287 (N_1287,N_1231,N_1248);
nor U1288 (N_1288,N_1202,N_1238);
and U1289 (N_1289,N_1242,N_1218);
nand U1290 (N_1290,N_1220,N_1214);
or U1291 (N_1291,N_1211,N_1233);
or U1292 (N_1292,N_1232,N_1220);
or U1293 (N_1293,N_1233,N_1227);
nand U1294 (N_1294,N_1229,N_1222);
nand U1295 (N_1295,N_1246,N_1247);
or U1296 (N_1296,N_1227,N_1247);
nand U1297 (N_1297,N_1215,N_1229);
nor U1298 (N_1298,N_1223,N_1205);
nor U1299 (N_1299,N_1233,N_1222);
xnor U1300 (N_1300,N_1250,N_1271);
or U1301 (N_1301,N_1268,N_1286);
nor U1302 (N_1302,N_1270,N_1287);
nand U1303 (N_1303,N_1285,N_1299);
nand U1304 (N_1304,N_1251,N_1291);
and U1305 (N_1305,N_1252,N_1261);
or U1306 (N_1306,N_1298,N_1269);
nand U1307 (N_1307,N_1253,N_1295);
and U1308 (N_1308,N_1277,N_1279);
and U1309 (N_1309,N_1274,N_1257);
nand U1310 (N_1310,N_1296,N_1284);
nand U1311 (N_1311,N_1292,N_1254);
xnor U1312 (N_1312,N_1272,N_1276);
or U1313 (N_1313,N_1258,N_1288);
nor U1314 (N_1314,N_1275,N_1294);
or U1315 (N_1315,N_1281,N_1259);
nand U1316 (N_1316,N_1256,N_1297);
and U1317 (N_1317,N_1283,N_1280);
nor U1318 (N_1318,N_1290,N_1266);
or U1319 (N_1319,N_1260,N_1264);
nand U1320 (N_1320,N_1273,N_1255);
nor U1321 (N_1321,N_1262,N_1282);
or U1322 (N_1322,N_1293,N_1265);
and U1323 (N_1323,N_1289,N_1278);
or U1324 (N_1324,N_1267,N_1263);
xnor U1325 (N_1325,N_1277,N_1268);
or U1326 (N_1326,N_1272,N_1285);
nand U1327 (N_1327,N_1282,N_1258);
and U1328 (N_1328,N_1250,N_1258);
or U1329 (N_1329,N_1260,N_1268);
or U1330 (N_1330,N_1280,N_1271);
nand U1331 (N_1331,N_1273,N_1251);
and U1332 (N_1332,N_1295,N_1293);
and U1333 (N_1333,N_1291,N_1257);
nor U1334 (N_1334,N_1293,N_1283);
or U1335 (N_1335,N_1282,N_1252);
nor U1336 (N_1336,N_1279,N_1296);
or U1337 (N_1337,N_1298,N_1295);
nand U1338 (N_1338,N_1294,N_1296);
nor U1339 (N_1339,N_1250,N_1284);
and U1340 (N_1340,N_1260,N_1265);
nor U1341 (N_1341,N_1271,N_1262);
nand U1342 (N_1342,N_1293,N_1294);
and U1343 (N_1343,N_1251,N_1296);
nand U1344 (N_1344,N_1264,N_1250);
nor U1345 (N_1345,N_1279,N_1298);
nor U1346 (N_1346,N_1272,N_1263);
nor U1347 (N_1347,N_1255,N_1298);
nor U1348 (N_1348,N_1273,N_1277);
nor U1349 (N_1349,N_1253,N_1250);
nor U1350 (N_1350,N_1322,N_1342);
and U1351 (N_1351,N_1323,N_1310);
nor U1352 (N_1352,N_1339,N_1330);
and U1353 (N_1353,N_1345,N_1314);
xor U1354 (N_1354,N_1308,N_1315);
and U1355 (N_1355,N_1336,N_1329);
nor U1356 (N_1356,N_1319,N_1333);
or U1357 (N_1357,N_1325,N_1321);
or U1358 (N_1358,N_1338,N_1312);
nand U1359 (N_1359,N_1320,N_1309);
and U1360 (N_1360,N_1335,N_1346);
and U1361 (N_1361,N_1300,N_1337);
and U1362 (N_1362,N_1340,N_1313);
or U1363 (N_1363,N_1305,N_1349);
nor U1364 (N_1364,N_1316,N_1307);
and U1365 (N_1365,N_1301,N_1328);
nand U1366 (N_1366,N_1343,N_1348);
nor U1367 (N_1367,N_1304,N_1317);
nand U1368 (N_1368,N_1334,N_1326);
and U1369 (N_1369,N_1344,N_1347);
nor U1370 (N_1370,N_1332,N_1324);
nor U1371 (N_1371,N_1331,N_1341);
nor U1372 (N_1372,N_1303,N_1302);
and U1373 (N_1373,N_1327,N_1311);
or U1374 (N_1374,N_1306,N_1318);
or U1375 (N_1375,N_1303,N_1345);
nand U1376 (N_1376,N_1338,N_1339);
xor U1377 (N_1377,N_1332,N_1343);
and U1378 (N_1378,N_1336,N_1303);
nand U1379 (N_1379,N_1301,N_1317);
nand U1380 (N_1380,N_1300,N_1309);
nor U1381 (N_1381,N_1302,N_1345);
nor U1382 (N_1382,N_1349,N_1345);
and U1383 (N_1383,N_1305,N_1348);
or U1384 (N_1384,N_1318,N_1330);
nand U1385 (N_1385,N_1312,N_1323);
nor U1386 (N_1386,N_1346,N_1302);
nand U1387 (N_1387,N_1331,N_1348);
nor U1388 (N_1388,N_1337,N_1338);
and U1389 (N_1389,N_1345,N_1333);
or U1390 (N_1390,N_1342,N_1312);
or U1391 (N_1391,N_1310,N_1318);
and U1392 (N_1392,N_1323,N_1316);
or U1393 (N_1393,N_1304,N_1347);
or U1394 (N_1394,N_1337,N_1317);
nor U1395 (N_1395,N_1321,N_1330);
or U1396 (N_1396,N_1317,N_1347);
nor U1397 (N_1397,N_1340,N_1347);
nand U1398 (N_1398,N_1307,N_1327);
and U1399 (N_1399,N_1317,N_1330);
nand U1400 (N_1400,N_1393,N_1357);
and U1401 (N_1401,N_1371,N_1397);
nor U1402 (N_1402,N_1399,N_1385);
nor U1403 (N_1403,N_1352,N_1351);
or U1404 (N_1404,N_1350,N_1362);
and U1405 (N_1405,N_1367,N_1368);
nand U1406 (N_1406,N_1390,N_1354);
and U1407 (N_1407,N_1373,N_1359);
nor U1408 (N_1408,N_1384,N_1363);
or U1409 (N_1409,N_1360,N_1391);
xnor U1410 (N_1410,N_1387,N_1370);
and U1411 (N_1411,N_1353,N_1374);
and U1412 (N_1412,N_1372,N_1375);
nor U1413 (N_1413,N_1364,N_1394);
nor U1414 (N_1414,N_1395,N_1382);
nand U1415 (N_1415,N_1369,N_1381);
or U1416 (N_1416,N_1366,N_1377);
nor U1417 (N_1417,N_1388,N_1383);
nand U1418 (N_1418,N_1379,N_1398);
and U1419 (N_1419,N_1376,N_1361);
and U1420 (N_1420,N_1389,N_1356);
and U1421 (N_1421,N_1386,N_1358);
nor U1422 (N_1422,N_1396,N_1378);
or U1423 (N_1423,N_1392,N_1380);
and U1424 (N_1424,N_1355,N_1365);
nand U1425 (N_1425,N_1369,N_1371);
and U1426 (N_1426,N_1375,N_1350);
and U1427 (N_1427,N_1350,N_1365);
nor U1428 (N_1428,N_1357,N_1382);
and U1429 (N_1429,N_1371,N_1366);
nor U1430 (N_1430,N_1387,N_1391);
nand U1431 (N_1431,N_1368,N_1364);
nand U1432 (N_1432,N_1373,N_1397);
and U1433 (N_1433,N_1386,N_1396);
nand U1434 (N_1434,N_1361,N_1350);
nand U1435 (N_1435,N_1364,N_1398);
and U1436 (N_1436,N_1375,N_1379);
and U1437 (N_1437,N_1357,N_1372);
and U1438 (N_1438,N_1365,N_1369);
and U1439 (N_1439,N_1363,N_1380);
or U1440 (N_1440,N_1368,N_1399);
nor U1441 (N_1441,N_1378,N_1370);
and U1442 (N_1442,N_1368,N_1353);
or U1443 (N_1443,N_1366,N_1367);
nand U1444 (N_1444,N_1366,N_1363);
and U1445 (N_1445,N_1361,N_1355);
nand U1446 (N_1446,N_1390,N_1368);
or U1447 (N_1447,N_1379,N_1359);
and U1448 (N_1448,N_1351,N_1383);
or U1449 (N_1449,N_1372,N_1360);
nand U1450 (N_1450,N_1421,N_1446);
nor U1451 (N_1451,N_1438,N_1428);
and U1452 (N_1452,N_1412,N_1420);
nand U1453 (N_1453,N_1441,N_1426);
or U1454 (N_1454,N_1447,N_1442);
or U1455 (N_1455,N_1409,N_1401);
nand U1456 (N_1456,N_1430,N_1436);
nor U1457 (N_1457,N_1422,N_1417);
or U1458 (N_1458,N_1407,N_1440);
nor U1459 (N_1459,N_1433,N_1434);
nand U1460 (N_1460,N_1413,N_1427);
nand U1461 (N_1461,N_1444,N_1448);
and U1462 (N_1462,N_1416,N_1400);
nand U1463 (N_1463,N_1445,N_1406);
or U1464 (N_1464,N_1424,N_1431);
nand U1465 (N_1465,N_1410,N_1405);
nand U1466 (N_1466,N_1425,N_1419);
or U1467 (N_1467,N_1432,N_1402);
or U1468 (N_1468,N_1443,N_1415);
nand U1469 (N_1469,N_1423,N_1408);
nor U1470 (N_1470,N_1429,N_1418);
or U1471 (N_1471,N_1449,N_1414);
and U1472 (N_1472,N_1404,N_1435);
nor U1473 (N_1473,N_1411,N_1437);
or U1474 (N_1474,N_1439,N_1403);
nand U1475 (N_1475,N_1419,N_1446);
nand U1476 (N_1476,N_1426,N_1448);
nand U1477 (N_1477,N_1426,N_1433);
nor U1478 (N_1478,N_1407,N_1417);
or U1479 (N_1479,N_1437,N_1426);
nand U1480 (N_1480,N_1411,N_1420);
nor U1481 (N_1481,N_1404,N_1419);
and U1482 (N_1482,N_1415,N_1421);
nor U1483 (N_1483,N_1407,N_1411);
or U1484 (N_1484,N_1431,N_1416);
or U1485 (N_1485,N_1448,N_1445);
and U1486 (N_1486,N_1446,N_1417);
nand U1487 (N_1487,N_1412,N_1405);
and U1488 (N_1488,N_1440,N_1410);
and U1489 (N_1489,N_1409,N_1408);
nand U1490 (N_1490,N_1449,N_1431);
or U1491 (N_1491,N_1416,N_1443);
xnor U1492 (N_1492,N_1408,N_1402);
nor U1493 (N_1493,N_1444,N_1446);
or U1494 (N_1494,N_1449,N_1409);
nand U1495 (N_1495,N_1422,N_1437);
and U1496 (N_1496,N_1418,N_1405);
or U1497 (N_1497,N_1400,N_1417);
and U1498 (N_1498,N_1434,N_1411);
or U1499 (N_1499,N_1418,N_1445);
or U1500 (N_1500,N_1479,N_1499);
and U1501 (N_1501,N_1450,N_1491);
or U1502 (N_1502,N_1457,N_1497);
nand U1503 (N_1503,N_1466,N_1459);
nand U1504 (N_1504,N_1452,N_1467);
and U1505 (N_1505,N_1455,N_1495);
nand U1506 (N_1506,N_1460,N_1475);
or U1507 (N_1507,N_1454,N_1465);
or U1508 (N_1508,N_1487,N_1463);
nand U1509 (N_1509,N_1492,N_1471);
and U1510 (N_1510,N_1464,N_1474);
and U1511 (N_1511,N_1477,N_1484);
nor U1512 (N_1512,N_1480,N_1456);
or U1513 (N_1513,N_1490,N_1462);
or U1514 (N_1514,N_1494,N_1498);
nand U1515 (N_1515,N_1478,N_1470);
and U1516 (N_1516,N_1461,N_1482);
and U1517 (N_1517,N_1469,N_1468);
nor U1518 (N_1518,N_1496,N_1486);
and U1519 (N_1519,N_1493,N_1485);
or U1520 (N_1520,N_1481,N_1483);
or U1521 (N_1521,N_1451,N_1458);
or U1522 (N_1522,N_1473,N_1489);
nor U1523 (N_1523,N_1476,N_1453);
or U1524 (N_1524,N_1472,N_1488);
or U1525 (N_1525,N_1450,N_1498);
nor U1526 (N_1526,N_1474,N_1481);
nor U1527 (N_1527,N_1458,N_1456);
or U1528 (N_1528,N_1489,N_1459);
nand U1529 (N_1529,N_1492,N_1496);
and U1530 (N_1530,N_1479,N_1492);
or U1531 (N_1531,N_1460,N_1462);
or U1532 (N_1532,N_1491,N_1463);
nand U1533 (N_1533,N_1476,N_1471);
or U1534 (N_1534,N_1460,N_1457);
nand U1535 (N_1535,N_1475,N_1459);
nor U1536 (N_1536,N_1459,N_1473);
nor U1537 (N_1537,N_1490,N_1474);
nor U1538 (N_1538,N_1466,N_1471);
or U1539 (N_1539,N_1463,N_1459);
nor U1540 (N_1540,N_1482,N_1474);
nand U1541 (N_1541,N_1451,N_1453);
nor U1542 (N_1542,N_1487,N_1456);
or U1543 (N_1543,N_1498,N_1460);
or U1544 (N_1544,N_1472,N_1465);
nor U1545 (N_1545,N_1463,N_1460);
or U1546 (N_1546,N_1486,N_1450);
or U1547 (N_1547,N_1497,N_1456);
nor U1548 (N_1548,N_1456,N_1457);
nor U1549 (N_1549,N_1481,N_1462);
and U1550 (N_1550,N_1530,N_1544);
nand U1551 (N_1551,N_1527,N_1502);
nand U1552 (N_1552,N_1524,N_1531);
and U1553 (N_1553,N_1511,N_1523);
and U1554 (N_1554,N_1507,N_1535);
and U1555 (N_1555,N_1539,N_1503);
nor U1556 (N_1556,N_1534,N_1521);
nand U1557 (N_1557,N_1529,N_1504);
or U1558 (N_1558,N_1528,N_1517);
nor U1559 (N_1559,N_1518,N_1520);
and U1560 (N_1560,N_1549,N_1525);
nand U1561 (N_1561,N_1548,N_1537);
and U1562 (N_1562,N_1505,N_1513);
and U1563 (N_1563,N_1533,N_1532);
or U1564 (N_1564,N_1526,N_1510);
nand U1565 (N_1565,N_1542,N_1515);
or U1566 (N_1566,N_1522,N_1514);
nor U1567 (N_1567,N_1543,N_1509);
nand U1568 (N_1568,N_1500,N_1501);
or U1569 (N_1569,N_1536,N_1512);
and U1570 (N_1570,N_1545,N_1541);
and U1571 (N_1571,N_1546,N_1540);
or U1572 (N_1572,N_1547,N_1519);
nor U1573 (N_1573,N_1508,N_1538);
nand U1574 (N_1574,N_1516,N_1506);
nor U1575 (N_1575,N_1535,N_1541);
and U1576 (N_1576,N_1517,N_1542);
or U1577 (N_1577,N_1520,N_1503);
nor U1578 (N_1578,N_1542,N_1501);
and U1579 (N_1579,N_1541,N_1500);
or U1580 (N_1580,N_1508,N_1501);
or U1581 (N_1581,N_1511,N_1541);
nand U1582 (N_1582,N_1510,N_1511);
or U1583 (N_1583,N_1500,N_1529);
or U1584 (N_1584,N_1537,N_1508);
nand U1585 (N_1585,N_1533,N_1512);
nand U1586 (N_1586,N_1514,N_1549);
nand U1587 (N_1587,N_1524,N_1501);
nor U1588 (N_1588,N_1526,N_1509);
nor U1589 (N_1589,N_1534,N_1532);
or U1590 (N_1590,N_1500,N_1549);
nand U1591 (N_1591,N_1525,N_1538);
or U1592 (N_1592,N_1518,N_1546);
nor U1593 (N_1593,N_1534,N_1506);
or U1594 (N_1594,N_1546,N_1548);
and U1595 (N_1595,N_1514,N_1521);
nand U1596 (N_1596,N_1508,N_1517);
or U1597 (N_1597,N_1532,N_1502);
and U1598 (N_1598,N_1518,N_1543);
nor U1599 (N_1599,N_1515,N_1548);
or U1600 (N_1600,N_1592,N_1588);
and U1601 (N_1601,N_1569,N_1571);
nor U1602 (N_1602,N_1579,N_1564);
nor U1603 (N_1603,N_1594,N_1556);
nor U1604 (N_1604,N_1557,N_1565);
xor U1605 (N_1605,N_1593,N_1583);
nor U1606 (N_1606,N_1561,N_1553);
nand U1607 (N_1607,N_1582,N_1554);
nand U1608 (N_1608,N_1595,N_1586);
or U1609 (N_1609,N_1578,N_1574);
or U1610 (N_1610,N_1563,N_1598);
and U1611 (N_1611,N_1562,N_1568);
and U1612 (N_1612,N_1570,N_1589);
nand U1613 (N_1613,N_1596,N_1559);
or U1614 (N_1614,N_1550,N_1572);
nor U1615 (N_1615,N_1591,N_1560);
or U1616 (N_1616,N_1576,N_1590);
or U1617 (N_1617,N_1552,N_1580);
and U1618 (N_1618,N_1581,N_1575);
nor U1619 (N_1619,N_1584,N_1567);
nand U1620 (N_1620,N_1558,N_1585);
nor U1621 (N_1621,N_1597,N_1587);
nor U1622 (N_1622,N_1577,N_1573);
nor U1623 (N_1623,N_1599,N_1551);
nand U1624 (N_1624,N_1555,N_1566);
or U1625 (N_1625,N_1594,N_1583);
and U1626 (N_1626,N_1595,N_1565);
nor U1627 (N_1627,N_1598,N_1580);
and U1628 (N_1628,N_1587,N_1575);
nand U1629 (N_1629,N_1593,N_1552);
nand U1630 (N_1630,N_1570,N_1569);
or U1631 (N_1631,N_1579,N_1560);
and U1632 (N_1632,N_1562,N_1559);
nand U1633 (N_1633,N_1598,N_1555);
or U1634 (N_1634,N_1593,N_1551);
and U1635 (N_1635,N_1551,N_1563);
nor U1636 (N_1636,N_1580,N_1586);
nor U1637 (N_1637,N_1558,N_1564);
nor U1638 (N_1638,N_1554,N_1586);
or U1639 (N_1639,N_1592,N_1595);
nor U1640 (N_1640,N_1595,N_1575);
or U1641 (N_1641,N_1593,N_1587);
nor U1642 (N_1642,N_1592,N_1574);
nor U1643 (N_1643,N_1554,N_1562);
nand U1644 (N_1644,N_1579,N_1577);
nand U1645 (N_1645,N_1571,N_1553);
and U1646 (N_1646,N_1593,N_1585);
and U1647 (N_1647,N_1554,N_1567);
nand U1648 (N_1648,N_1559,N_1579);
nor U1649 (N_1649,N_1560,N_1561);
nand U1650 (N_1650,N_1636,N_1639);
and U1651 (N_1651,N_1643,N_1649);
or U1652 (N_1652,N_1630,N_1641);
nand U1653 (N_1653,N_1617,N_1622);
and U1654 (N_1654,N_1608,N_1615);
and U1655 (N_1655,N_1625,N_1640);
nor U1656 (N_1656,N_1645,N_1620);
nand U1657 (N_1657,N_1624,N_1600);
and U1658 (N_1658,N_1616,N_1612);
nand U1659 (N_1659,N_1619,N_1609);
or U1660 (N_1660,N_1632,N_1633);
or U1661 (N_1661,N_1631,N_1605);
or U1662 (N_1662,N_1603,N_1629);
and U1663 (N_1663,N_1626,N_1623);
nor U1664 (N_1664,N_1621,N_1634);
or U1665 (N_1665,N_1602,N_1637);
nor U1666 (N_1666,N_1644,N_1614);
nand U1667 (N_1667,N_1635,N_1618);
and U1668 (N_1668,N_1611,N_1648);
or U1669 (N_1669,N_1607,N_1628);
or U1670 (N_1670,N_1646,N_1606);
or U1671 (N_1671,N_1601,N_1613);
or U1672 (N_1672,N_1610,N_1647);
nor U1673 (N_1673,N_1642,N_1604);
and U1674 (N_1674,N_1627,N_1638);
or U1675 (N_1675,N_1616,N_1620);
nor U1676 (N_1676,N_1618,N_1640);
xnor U1677 (N_1677,N_1644,N_1616);
nand U1678 (N_1678,N_1622,N_1619);
and U1679 (N_1679,N_1647,N_1601);
nand U1680 (N_1680,N_1634,N_1612);
and U1681 (N_1681,N_1627,N_1600);
nand U1682 (N_1682,N_1642,N_1602);
nor U1683 (N_1683,N_1634,N_1610);
or U1684 (N_1684,N_1624,N_1609);
nand U1685 (N_1685,N_1640,N_1645);
nand U1686 (N_1686,N_1638,N_1600);
nand U1687 (N_1687,N_1625,N_1620);
nor U1688 (N_1688,N_1603,N_1609);
and U1689 (N_1689,N_1606,N_1617);
nor U1690 (N_1690,N_1622,N_1600);
and U1691 (N_1691,N_1618,N_1602);
or U1692 (N_1692,N_1639,N_1603);
nor U1693 (N_1693,N_1625,N_1647);
or U1694 (N_1694,N_1644,N_1609);
or U1695 (N_1695,N_1608,N_1600);
and U1696 (N_1696,N_1648,N_1638);
nor U1697 (N_1697,N_1620,N_1633);
nand U1698 (N_1698,N_1645,N_1601);
nor U1699 (N_1699,N_1616,N_1608);
and U1700 (N_1700,N_1688,N_1673);
nand U1701 (N_1701,N_1663,N_1680);
nand U1702 (N_1702,N_1672,N_1692);
and U1703 (N_1703,N_1690,N_1686);
or U1704 (N_1704,N_1661,N_1689);
nor U1705 (N_1705,N_1679,N_1665);
xnor U1706 (N_1706,N_1676,N_1698);
or U1707 (N_1707,N_1650,N_1699);
and U1708 (N_1708,N_1671,N_1669);
and U1709 (N_1709,N_1691,N_1685);
and U1710 (N_1710,N_1687,N_1670);
nand U1711 (N_1711,N_1682,N_1658);
nor U1712 (N_1712,N_1693,N_1667);
xnor U1713 (N_1713,N_1664,N_1675);
or U1714 (N_1714,N_1677,N_1662);
and U1715 (N_1715,N_1656,N_1651);
and U1716 (N_1716,N_1655,N_1696);
or U1717 (N_1717,N_1666,N_1654);
or U1718 (N_1718,N_1695,N_1652);
nand U1719 (N_1719,N_1694,N_1674);
and U1720 (N_1720,N_1657,N_1653);
nor U1721 (N_1721,N_1659,N_1660);
or U1722 (N_1722,N_1681,N_1668);
or U1723 (N_1723,N_1684,N_1678);
xor U1724 (N_1724,N_1697,N_1683);
and U1725 (N_1725,N_1682,N_1687);
nand U1726 (N_1726,N_1677,N_1693);
or U1727 (N_1727,N_1696,N_1697);
or U1728 (N_1728,N_1667,N_1699);
or U1729 (N_1729,N_1687,N_1657);
nor U1730 (N_1730,N_1699,N_1690);
and U1731 (N_1731,N_1661,N_1696);
nor U1732 (N_1732,N_1690,N_1689);
nand U1733 (N_1733,N_1665,N_1686);
nor U1734 (N_1734,N_1688,N_1662);
nand U1735 (N_1735,N_1664,N_1688);
and U1736 (N_1736,N_1657,N_1655);
nand U1737 (N_1737,N_1681,N_1654);
and U1738 (N_1738,N_1665,N_1671);
nand U1739 (N_1739,N_1667,N_1656);
nand U1740 (N_1740,N_1663,N_1691);
nand U1741 (N_1741,N_1656,N_1682);
or U1742 (N_1742,N_1671,N_1682);
nand U1743 (N_1743,N_1656,N_1684);
or U1744 (N_1744,N_1655,N_1654);
and U1745 (N_1745,N_1680,N_1667);
nand U1746 (N_1746,N_1660,N_1653);
nor U1747 (N_1747,N_1697,N_1651);
or U1748 (N_1748,N_1664,N_1697);
nand U1749 (N_1749,N_1689,N_1688);
or U1750 (N_1750,N_1734,N_1729);
nand U1751 (N_1751,N_1746,N_1742);
nand U1752 (N_1752,N_1700,N_1706);
nor U1753 (N_1753,N_1740,N_1738);
or U1754 (N_1754,N_1711,N_1701);
or U1755 (N_1755,N_1728,N_1704);
or U1756 (N_1756,N_1718,N_1716);
xor U1757 (N_1757,N_1702,N_1733);
and U1758 (N_1758,N_1710,N_1748);
nand U1759 (N_1759,N_1744,N_1703);
nor U1760 (N_1760,N_1731,N_1727);
and U1761 (N_1761,N_1741,N_1715);
nor U1762 (N_1762,N_1707,N_1732);
and U1763 (N_1763,N_1719,N_1720);
nor U1764 (N_1764,N_1709,N_1735);
nand U1765 (N_1765,N_1725,N_1730);
nand U1766 (N_1766,N_1745,N_1737);
or U1767 (N_1767,N_1717,N_1749);
nand U1768 (N_1768,N_1736,N_1724);
or U1769 (N_1769,N_1723,N_1721);
or U1770 (N_1770,N_1708,N_1712);
and U1771 (N_1771,N_1747,N_1714);
nor U1772 (N_1772,N_1705,N_1722);
or U1773 (N_1773,N_1743,N_1726);
or U1774 (N_1774,N_1739,N_1713);
nand U1775 (N_1775,N_1748,N_1717);
nand U1776 (N_1776,N_1718,N_1715);
and U1777 (N_1777,N_1715,N_1735);
nand U1778 (N_1778,N_1717,N_1723);
and U1779 (N_1779,N_1707,N_1703);
and U1780 (N_1780,N_1713,N_1736);
or U1781 (N_1781,N_1707,N_1731);
nor U1782 (N_1782,N_1740,N_1747);
xnor U1783 (N_1783,N_1722,N_1729);
nand U1784 (N_1784,N_1721,N_1725);
nand U1785 (N_1785,N_1743,N_1702);
or U1786 (N_1786,N_1749,N_1743);
nand U1787 (N_1787,N_1735,N_1704);
nor U1788 (N_1788,N_1728,N_1710);
nand U1789 (N_1789,N_1735,N_1741);
nand U1790 (N_1790,N_1735,N_1725);
nor U1791 (N_1791,N_1742,N_1749);
nand U1792 (N_1792,N_1748,N_1739);
nand U1793 (N_1793,N_1724,N_1701);
nand U1794 (N_1794,N_1710,N_1742);
or U1795 (N_1795,N_1748,N_1708);
nand U1796 (N_1796,N_1713,N_1724);
or U1797 (N_1797,N_1721,N_1728);
or U1798 (N_1798,N_1736,N_1715);
and U1799 (N_1799,N_1709,N_1742);
or U1800 (N_1800,N_1777,N_1765);
or U1801 (N_1801,N_1773,N_1767);
nor U1802 (N_1802,N_1758,N_1787);
nor U1803 (N_1803,N_1759,N_1784);
nand U1804 (N_1804,N_1791,N_1760);
or U1805 (N_1805,N_1798,N_1770);
and U1806 (N_1806,N_1762,N_1753);
xor U1807 (N_1807,N_1764,N_1780);
nor U1808 (N_1808,N_1774,N_1793);
and U1809 (N_1809,N_1775,N_1789);
and U1810 (N_1810,N_1785,N_1794);
nand U1811 (N_1811,N_1799,N_1769);
nand U1812 (N_1812,N_1752,N_1768);
and U1813 (N_1813,N_1786,N_1792);
nor U1814 (N_1814,N_1750,N_1766);
or U1815 (N_1815,N_1782,N_1761);
and U1816 (N_1816,N_1756,N_1751);
nand U1817 (N_1817,N_1779,N_1776);
and U1818 (N_1818,N_1755,N_1772);
nand U1819 (N_1819,N_1771,N_1796);
nand U1820 (N_1820,N_1781,N_1783);
and U1821 (N_1821,N_1754,N_1778);
or U1822 (N_1822,N_1795,N_1763);
and U1823 (N_1823,N_1757,N_1797);
nor U1824 (N_1824,N_1788,N_1790);
nor U1825 (N_1825,N_1756,N_1787);
and U1826 (N_1826,N_1799,N_1796);
nand U1827 (N_1827,N_1766,N_1770);
nor U1828 (N_1828,N_1779,N_1773);
and U1829 (N_1829,N_1762,N_1784);
nand U1830 (N_1830,N_1793,N_1771);
and U1831 (N_1831,N_1799,N_1795);
and U1832 (N_1832,N_1783,N_1766);
nand U1833 (N_1833,N_1794,N_1760);
or U1834 (N_1834,N_1774,N_1763);
nor U1835 (N_1835,N_1766,N_1777);
or U1836 (N_1836,N_1751,N_1782);
or U1837 (N_1837,N_1769,N_1761);
and U1838 (N_1838,N_1750,N_1759);
nand U1839 (N_1839,N_1776,N_1793);
nor U1840 (N_1840,N_1754,N_1776);
nor U1841 (N_1841,N_1796,N_1787);
nand U1842 (N_1842,N_1792,N_1777);
and U1843 (N_1843,N_1754,N_1756);
nand U1844 (N_1844,N_1787,N_1798);
nand U1845 (N_1845,N_1772,N_1777);
nand U1846 (N_1846,N_1791,N_1796);
or U1847 (N_1847,N_1790,N_1758);
nor U1848 (N_1848,N_1776,N_1757);
or U1849 (N_1849,N_1784,N_1770);
or U1850 (N_1850,N_1801,N_1828);
nand U1851 (N_1851,N_1819,N_1842);
and U1852 (N_1852,N_1803,N_1805);
and U1853 (N_1853,N_1845,N_1822);
and U1854 (N_1854,N_1810,N_1809);
nand U1855 (N_1855,N_1841,N_1826);
nor U1856 (N_1856,N_1843,N_1800);
or U1857 (N_1857,N_1814,N_1836);
nor U1858 (N_1858,N_1847,N_1815);
nor U1859 (N_1859,N_1807,N_1818);
and U1860 (N_1860,N_1823,N_1827);
or U1861 (N_1861,N_1802,N_1812);
nand U1862 (N_1862,N_1839,N_1838);
and U1863 (N_1863,N_1849,N_1848);
nand U1864 (N_1864,N_1830,N_1820);
nor U1865 (N_1865,N_1834,N_1833);
and U1866 (N_1866,N_1846,N_1811);
nor U1867 (N_1867,N_1832,N_1824);
or U1868 (N_1868,N_1844,N_1837);
nand U1869 (N_1869,N_1829,N_1835);
and U1870 (N_1870,N_1804,N_1821);
or U1871 (N_1871,N_1831,N_1840);
nand U1872 (N_1872,N_1808,N_1825);
nor U1873 (N_1873,N_1817,N_1813);
nand U1874 (N_1874,N_1806,N_1816);
nor U1875 (N_1875,N_1824,N_1841);
nor U1876 (N_1876,N_1829,N_1836);
nor U1877 (N_1877,N_1836,N_1846);
or U1878 (N_1878,N_1845,N_1800);
and U1879 (N_1879,N_1824,N_1822);
nor U1880 (N_1880,N_1842,N_1823);
nor U1881 (N_1881,N_1824,N_1805);
nor U1882 (N_1882,N_1806,N_1810);
or U1883 (N_1883,N_1817,N_1824);
and U1884 (N_1884,N_1804,N_1803);
and U1885 (N_1885,N_1800,N_1807);
and U1886 (N_1886,N_1821,N_1842);
nor U1887 (N_1887,N_1817,N_1814);
nand U1888 (N_1888,N_1826,N_1825);
nor U1889 (N_1889,N_1829,N_1824);
and U1890 (N_1890,N_1833,N_1843);
nand U1891 (N_1891,N_1808,N_1848);
nor U1892 (N_1892,N_1810,N_1835);
and U1893 (N_1893,N_1802,N_1838);
and U1894 (N_1894,N_1839,N_1842);
nor U1895 (N_1895,N_1814,N_1831);
nor U1896 (N_1896,N_1821,N_1829);
nand U1897 (N_1897,N_1832,N_1809);
or U1898 (N_1898,N_1806,N_1802);
and U1899 (N_1899,N_1813,N_1815);
nand U1900 (N_1900,N_1889,N_1882);
or U1901 (N_1901,N_1895,N_1874);
or U1902 (N_1902,N_1850,N_1871);
nor U1903 (N_1903,N_1875,N_1897);
nand U1904 (N_1904,N_1858,N_1898);
or U1905 (N_1905,N_1863,N_1899);
or U1906 (N_1906,N_1872,N_1867);
or U1907 (N_1907,N_1891,N_1860);
nand U1908 (N_1908,N_1870,N_1878);
or U1909 (N_1909,N_1861,N_1881);
and U1910 (N_1910,N_1851,N_1853);
nand U1911 (N_1911,N_1892,N_1885);
nor U1912 (N_1912,N_1862,N_1896);
and U1913 (N_1913,N_1866,N_1890);
nor U1914 (N_1914,N_1880,N_1884);
nor U1915 (N_1915,N_1868,N_1865);
and U1916 (N_1916,N_1888,N_1859);
or U1917 (N_1917,N_1887,N_1893);
or U1918 (N_1918,N_1886,N_1864);
nor U1919 (N_1919,N_1856,N_1894);
or U1920 (N_1920,N_1854,N_1883);
and U1921 (N_1921,N_1855,N_1873);
and U1922 (N_1922,N_1852,N_1876);
or U1923 (N_1923,N_1857,N_1879);
nor U1924 (N_1924,N_1869,N_1877);
or U1925 (N_1925,N_1898,N_1885);
or U1926 (N_1926,N_1884,N_1853);
and U1927 (N_1927,N_1851,N_1897);
nor U1928 (N_1928,N_1894,N_1872);
or U1929 (N_1929,N_1854,N_1894);
and U1930 (N_1930,N_1881,N_1882);
nor U1931 (N_1931,N_1864,N_1850);
nor U1932 (N_1932,N_1877,N_1896);
nand U1933 (N_1933,N_1892,N_1875);
nand U1934 (N_1934,N_1861,N_1883);
or U1935 (N_1935,N_1865,N_1853);
nor U1936 (N_1936,N_1883,N_1860);
or U1937 (N_1937,N_1879,N_1888);
nand U1938 (N_1938,N_1881,N_1886);
nor U1939 (N_1939,N_1862,N_1857);
nand U1940 (N_1940,N_1866,N_1852);
and U1941 (N_1941,N_1865,N_1860);
nor U1942 (N_1942,N_1877,N_1851);
and U1943 (N_1943,N_1897,N_1887);
nand U1944 (N_1944,N_1867,N_1856);
nand U1945 (N_1945,N_1890,N_1892);
or U1946 (N_1946,N_1898,N_1881);
or U1947 (N_1947,N_1875,N_1853);
nand U1948 (N_1948,N_1899,N_1862);
or U1949 (N_1949,N_1877,N_1855);
xnor U1950 (N_1950,N_1910,N_1932);
nor U1951 (N_1951,N_1939,N_1902);
nand U1952 (N_1952,N_1913,N_1914);
and U1953 (N_1953,N_1915,N_1906);
nor U1954 (N_1954,N_1900,N_1908);
nor U1955 (N_1955,N_1940,N_1943);
or U1956 (N_1956,N_1924,N_1918);
or U1957 (N_1957,N_1949,N_1927);
nor U1958 (N_1958,N_1931,N_1934);
or U1959 (N_1959,N_1946,N_1944);
and U1960 (N_1960,N_1923,N_1903);
nand U1961 (N_1961,N_1941,N_1911);
and U1962 (N_1962,N_1928,N_1942);
and U1963 (N_1963,N_1933,N_1912);
and U1964 (N_1964,N_1937,N_1921);
or U1965 (N_1965,N_1935,N_1905);
nor U1966 (N_1966,N_1936,N_1947);
nand U1967 (N_1967,N_1930,N_1919);
nand U1968 (N_1968,N_1938,N_1920);
nor U1969 (N_1969,N_1909,N_1945);
or U1970 (N_1970,N_1901,N_1926);
nor U1971 (N_1971,N_1922,N_1904);
nor U1972 (N_1972,N_1948,N_1916);
nand U1973 (N_1973,N_1929,N_1907);
nor U1974 (N_1974,N_1917,N_1925);
nand U1975 (N_1975,N_1907,N_1908);
nor U1976 (N_1976,N_1933,N_1944);
or U1977 (N_1977,N_1937,N_1909);
nand U1978 (N_1978,N_1928,N_1934);
and U1979 (N_1979,N_1911,N_1945);
nor U1980 (N_1980,N_1904,N_1943);
nor U1981 (N_1981,N_1922,N_1925);
and U1982 (N_1982,N_1901,N_1921);
nor U1983 (N_1983,N_1914,N_1906);
and U1984 (N_1984,N_1935,N_1915);
nor U1985 (N_1985,N_1949,N_1942);
and U1986 (N_1986,N_1908,N_1948);
and U1987 (N_1987,N_1945,N_1947);
or U1988 (N_1988,N_1929,N_1944);
nor U1989 (N_1989,N_1920,N_1911);
and U1990 (N_1990,N_1944,N_1902);
and U1991 (N_1991,N_1913,N_1932);
and U1992 (N_1992,N_1941,N_1946);
nor U1993 (N_1993,N_1930,N_1945);
or U1994 (N_1994,N_1935,N_1909);
nand U1995 (N_1995,N_1913,N_1919);
or U1996 (N_1996,N_1912,N_1925);
or U1997 (N_1997,N_1942,N_1930);
nor U1998 (N_1998,N_1923,N_1948);
nor U1999 (N_1999,N_1929,N_1901);
nand U2000 (N_2000,N_1958,N_1965);
nand U2001 (N_2001,N_1952,N_1961);
nor U2002 (N_2002,N_1966,N_1967);
nor U2003 (N_2003,N_1953,N_1978);
and U2004 (N_2004,N_1997,N_1979);
or U2005 (N_2005,N_1998,N_1962);
nor U2006 (N_2006,N_1996,N_1959);
and U2007 (N_2007,N_1970,N_1990);
nand U2008 (N_2008,N_1980,N_1972);
or U2009 (N_2009,N_1981,N_1975);
nor U2010 (N_2010,N_1950,N_1984);
and U2011 (N_2011,N_1985,N_1995);
and U2012 (N_2012,N_1973,N_1987);
nor U2013 (N_2013,N_1982,N_1971);
and U2014 (N_2014,N_1999,N_1988);
nor U2015 (N_2015,N_1976,N_1977);
nand U2016 (N_2016,N_1994,N_1957);
and U2017 (N_2017,N_1993,N_1954);
or U2018 (N_2018,N_1969,N_1951);
and U2019 (N_2019,N_1974,N_1992);
nand U2020 (N_2020,N_1964,N_1960);
nor U2021 (N_2021,N_1986,N_1956);
or U2022 (N_2022,N_1991,N_1963);
or U2023 (N_2023,N_1989,N_1955);
nor U2024 (N_2024,N_1968,N_1983);
and U2025 (N_2025,N_1969,N_1991);
and U2026 (N_2026,N_1982,N_1983);
nor U2027 (N_2027,N_1966,N_1971);
nand U2028 (N_2028,N_1992,N_1959);
and U2029 (N_2029,N_1971,N_1961);
and U2030 (N_2030,N_1968,N_1996);
or U2031 (N_2031,N_1964,N_1969);
nand U2032 (N_2032,N_1998,N_1996);
nand U2033 (N_2033,N_1968,N_1951);
or U2034 (N_2034,N_1952,N_1999);
and U2035 (N_2035,N_1990,N_1972);
and U2036 (N_2036,N_1961,N_1979);
nor U2037 (N_2037,N_1964,N_1978);
nand U2038 (N_2038,N_1998,N_1975);
nand U2039 (N_2039,N_1980,N_1960);
nand U2040 (N_2040,N_1969,N_1962);
or U2041 (N_2041,N_1953,N_1961);
and U2042 (N_2042,N_1966,N_1972);
nand U2043 (N_2043,N_1950,N_1972);
and U2044 (N_2044,N_1972,N_1956);
nand U2045 (N_2045,N_1958,N_1964);
nor U2046 (N_2046,N_1960,N_1986);
nor U2047 (N_2047,N_1989,N_1976);
nand U2048 (N_2048,N_1963,N_1981);
nor U2049 (N_2049,N_1989,N_1992);
and U2050 (N_2050,N_2046,N_2041);
or U2051 (N_2051,N_2001,N_2026);
nor U2052 (N_2052,N_2008,N_2033);
nor U2053 (N_2053,N_2037,N_2021);
nor U2054 (N_2054,N_2013,N_2035);
nor U2055 (N_2055,N_2002,N_2031);
nand U2056 (N_2056,N_2038,N_2044);
and U2057 (N_2057,N_2019,N_2030);
and U2058 (N_2058,N_2024,N_2027);
nand U2059 (N_2059,N_2009,N_2049);
nor U2060 (N_2060,N_2015,N_2011);
nor U2061 (N_2061,N_2003,N_2010);
nor U2062 (N_2062,N_2029,N_2007);
nand U2063 (N_2063,N_2045,N_2014);
nor U2064 (N_2064,N_2022,N_2042);
nor U2065 (N_2065,N_2017,N_2000);
nand U2066 (N_2066,N_2039,N_2020);
or U2067 (N_2067,N_2032,N_2018);
and U2068 (N_2068,N_2036,N_2006);
nor U2069 (N_2069,N_2034,N_2025);
and U2070 (N_2070,N_2012,N_2043);
and U2071 (N_2071,N_2028,N_2005);
or U2072 (N_2072,N_2047,N_2040);
nand U2073 (N_2073,N_2023,N_2048);
and U2074 (N_2074,N_2004,N_2016);
or U2075 (N_2075,N_2033,N_2049);
nor U2076 (N_2076,N_2012,N_2045);
and U2077 (N_2077,N_2016,N_2022);
or U2078 (N_2078,N_2005,N_2002);
nor U2079 (N_2079,N_2031,N_2035);
and U2080 (N_2080,N_2017,N_2009);
or U2081 (N_2081,N_2023,N_2049);
and U2082 (N_2082,N_2028,N_2003);
nor U2083 (N_2083,N_2044,N_2026);
and U2084 (N_2084,N_2008,N_2019);
nor U2085 (N_2085,N_2011,N_2024);
nor U2086 (N_2086,N_2031,N_2004);
or U2087 (N_2087,N_2018,N_2030);
or U2088 (N_2088,N_2011,N_2018);
nand U2089 (N_2089,N_2037,N_2030);
and U2090 (N_2090,N_2048,N_2006);
nor U2091 (N_2091,N_2024,N_2031);
nor U2092 (N_2092,N_2007,N_2021);
and U2093 (N_2093,N_2015,N_2022);
xnor U2094 (N_2094,N_2043,N_2013);
or U2095 (N_2095,N_2000,N_2003);
nor U2096 (N_2096,N_2021,N_2000);
and U2097 (N_2097,N_2032,N_2028);
or U2098 (N_2098,N_2049,N_2020);
or U2099 (N_2099,N_2016,N_2026);
and U2100 (N_2100,N_2067,N_2071);
nor U2101 (N_2101,N_2073,N_2077);
and U2102 (N_2102,N_2075,N_2088);
nor U2103 (N_2103,N_2091,N_2050);
and U2104 (N_2104,N_2051,N_2098);
and U2105 (N_2105,N_2086,N_2090);
and U2106 (N_2106,N_2089,N_2083);
nand U2107 (N_2107,N_2054,N_2055);
or U2108 (N_2108,N_2097,N_2092);
and U2109 (N_2109,N_2078,N_2082);
nand U2110 (N_2110,N_2068,N_2057);
or U2111 (N_2111,N_2093,N_2099);
nor U2112 (N_2112,N_2087,N_2058);
nor U2113 (N_2113,N_2070,N_2095);
nand U2114 (N_2114,N_2069,N_2056);
nand U2115 (N_2115,N_2094,N_2065);
nand U2116 (N_2116,N_2079,N_2059);
or U2117 (N_2117,N_2085,N_2081);
nand U2118 (N_2118,N_2052,N_2064);
nor U2119 (N_2119,N_2060,N_2096);
or U2120 (N_2120,N_2061,N_2062);
and U2121 (N_2121,N_2063,N_2084);
nand U2122 (N_2122,N_2076,N_2080);
nor U2123 (N_2123,N_2066,N_2072);
and U2124 (N_2124,N_2074,N_2053);
or U2125 (N_2125,N_2069,N_2068);
or U2126 (N_2126,N_2071,N_2068);
or U2127 (N_2127,N_2090,N_2074);
nand U2128 (N_2128,N_2082,N_2055);
nor U2129 (N_2129,N_2094,N_2056);
nand U2130 (N_2130,N_2057,N_2084);
nand U2131 (N_2131,N_2094,N_2063);
or U2132 (N_2132,N_2082,N_2093);
nor U2133 (N_2133,N_2062,N_2052);
nor U2134 (N_2134,N_2095,N_2067);
and U2135 (N_2135,N_2051,N_2069);
nor U2136 (N_2136,N_2064,N_2097);
nor U2137 (N_2137,N_2059,N_2064);
and U2138 (N_2138,N_2069,N_2089);
or U2139 (N_2139,N_2079,N_2073);
nor U2140 (N_2140,N_2080,N_2054);
nand U2141 (N_2141,N_2059,N_2051);
nand U2142 (N_2142,N_2076,N_2064);
and U2143 (N_2143,N_2069,N_2057);
or U2144 (N_2144,N_2060,N_2076);
and U2145 (N_2145,N_2099,N_2055);
or U2146 (N_2146,N_2080,N_2069);
and U2147 (N_2147,N_2084,N_2050);
nor U2148 (N_2148,N_2084,N_2097);
nor U2149 (N_2149,N_2069,N_2074);
or U2150 (N_2150,N_2109,N_2117);
and U2151 (N_2151,N_2147,N_2139);
nand U2152 (N_2152,N_2112,N_2145);
nand U2153 (N_2153,N_2130,N_2131);
and U2154 (N_2154,N_2114,N_2144);
nor U2155 (N_2155,N_2119,N_2113);
and U2156 (N_2156,N_2115,N_2141);
nor U2157 (N_2157,N_2116,N_2101);
or U2158 (N_2158,N_2124,N_2133);
and U2159 (N_2159,N_2125,N_2143);
nand U2160 (N_2160,N_2146,N_2122);
and U2161 (N_2161,N_2103,N_2118);
nand U2162 (N_2162,N_2127,N_2110);
xor U2163 (N_2163,N_2140,N_2108);
nor U2164 (N_2164,N_2126,N_2137);
nor U2165 (N_2165,N_2148,N_2142);
nand U2166 (N_2166,N_2121,N_2132);
and U2167 (N_2167,N_2135,N_2136);
nand U2168 (N_2168,N_2105,N_2138);
or U2169 (N_2169,N_2107,N_2149);
or U2170 (N_2170,N_2129,N_2123);
nand U2171 (N_2171,N_2128,N_2100);
nor U2172 (N_2172,N_2102,N_2111);
nand U2173 (N_2173,N_2104,N_2134);
and U2174 (N_2174,N_2106,N_2120);
xor U2175 (N_2175,N_2132,N_2138);
or U2176 (N_2176,N_2148,N_2136);
or U2177 (N_2177,N_2144,N_2120);
nand U2178 (N_2178,N_2107,N_2117);
and U2179 (N_2179,N_2101,N_2122);
and U2180 (N_2180,N_2125,N_2134);
or U2181 (N_2181,N_2106,N_2128);
nor U2182 (N_2182,N_2120,N_2115);
nor U2183 (N_2183,N_2106,N_2105);
or U2184 (N_2184,N_2138,N_2147);
nor U2185 (N_2185,N_2120,N_2141);
or U2186 (N_2186,N_2110,N_2143);
nand U2187 (N_2187,N_2127,N_2100);
xor U2188 (N_2188,N_2128,N_2145);
or U2189 (N_2189,N_2124,N_2101);
or U2190 (N_2190,N_2121,N_2101);
or U2191 (N_2191,N_2133,N_2122);
nor U2192 (N_2192,N_2111,N_2110);
and U2193 (N_2193,N_2116,N_2130);
or U2194 (N_2194,N_2106,N_2109);
or U2195 (N_2195,N_2138,N_2121);
nand U2196 (N_2196,N_2126,N_2109);
nand U2197 (N_2197,N_2105,N_2122);
and U2198 (N_2198,N_2134,N_2120);
and U2199 (N_2199,N_2107,N_2122);
or U2200 (N_2200,N_2171,N_2191);
or U2201 (N_2201,N_2195,N_2174);
nor U2202 (N_2202,N_2175,N_2177);
nand U2203 (N_2203,N_2151,N_2168);
and U2204 (N_2204,N_2162,N_2187);
nor U2205 (N_2205,N_2164,N_2184);
nor U2206 (N_2206,N_2167,N_2179);
nor U2207 (N_2207,N_2182,N_2156);
nand U2208 (N_2208,N_2169,N_2176);
or U2209 (N_2209,N_2157,N_2150);
and U2210 (N_2210,N_2183,N_2172);
nand U2211 (N_2211,N_2186,N_2163);
nor U2212 (N_2212,N_2188,N_2190);
nand U2213 (N_2213,N_2181,N_2155);
nand U2214 (N_2214,N_2199,N_2196);
nand U2215 (N_2215,N_2193,N_2153);
nand U2216 (N_2216,N_2197,N_2165);
xor U2217 (N_2217,N_2154,N_2178);
nor U2218 (N_2218,N_2194,N_2166);
nor U2219 (N_2219,N_2152,N_2159);
or U2220 (N_2220,N_2180,N_2198);
and U2221 (N_2221,N_2192,N_2161);
and U2222 (N_2222,N_2189,N_2185);
or U2223 (N_2223,N_2160,N_2158);
nor U2224 (N_2224,N_2173,N_2170);
or U2225 (N_2225,N_2165,N_2199);
xnor U2226 (N_2226,N_2159,N_2168);
or U2227 (N_2227,N_2177,N_2155);
or U2228 (N_2228,N_2186,N_2192);
or U2229 (N_2229,N_2154,N_2188);
nand U2230 (N_2230,N_2174,N_2167);
and U2231 (N_2231,N_2159,N_2160);
and U2232 (N_2232,N_2177,N_2168);
nand U2233 (N_2233,N_2175,N_2172);
and U2234 (N_2234,N_2162,N_2170);
nand U2235 (N_2235,N_2166,N_2172);
or U2236 (N_2236,N_2164,N_2186);
nand U2237 (N_2237,N_2160,N_2189);
or U2238 (N_2238,N_2155,N_2166);
and U2239 (N_2239,N_2171,N_2157);
nand U2240 (N_2240,N_2167,N_2189);
nor U2241 (N_2241,N_2169,N_2177);
or U2242 (N_2242,N_2163,N_2189);
and U2243 (N_2243,N_2184,N_2165);
nand U2244 (N_2244,N_2172,N_2161);
nor U2245 (N_2245,N_2168,N_2163);
nand U2246 (N_2246,N_2196,N_2162);
or U2247 (N_2247,N_2169,N_2155);
nor U2248 (N_2248,N_2195,N_2162);
nor U2249 (N_2249,N_2171,N_2186);
or U2250 (N_2250,N_2231,N_2215);
and U2251 (N_2251,N_2219,N_2236);
and U2252 (N_2252,N_2203,N_2222);
and U2253 (N_2253,N_2244,N_2246);
nand U2254 (N_2254,N_2209,N_2223);
and U2255 (N_2255,N_2240,N_2226);
nor U2256 (N_2256,N_2248,N_2234);
and U2257 (N_2257,N_2204,N_2237);
nor U2258 (N_2258,N_2229,N_2241);
nor U2259 (N_2259,N_2220,N_2225);
and U2260 (N_2260,N_2214,N_2233);
nor U2261 (N_2261,N_2249,N_2224);
nand U2262 (N_2262,N_2227,N_2247);
and U2263 (N_2263,N_2212,N_2235);
nand U2264 (N_2264,N_2216,N_2245);
and U2265 (N_2265,N_2217,N_2239);
nand U2266 (N_2266,N_2213,N_2205);
and U2267 (N_2267,N_2202,N_2230);
or U2268 (N_2268,N_2206,N_2211);
xnor U2269 (N_2269,N_2232,N_2221);
nand U2270 (N_2270,N_2238,N_2218);
nand U2271 (N_2271,N_2208,N_2200);
nor U2272 (N_2272,N_2243,N_2201);
nand U2273 (N_2273,N_2207,N_2210);
nor U2274 (N_2274,N_2242,N_2228);
nand U2275 (N_2275,N_2228,N_2243);
nand U2276 (N_2276,N_2217,N_2212);
and U2277 (N_2277,N_2249,N_2226);
nor U2278 (N_2278,N_2208,N_2217);
nor U2279 (N_2279,N_2245,N_2225);
and U2280 (N_2280,N_2249,N_2239);
nand U2281 (N_2281,N_2222,N_2201);
nor U2282 (N_2282,N_2229,N_2245);
nor U2283 (N_2283,N_2234,N_2217);
nand U2284 (N_2284,N_2235,N_2209);
and U2285 (N_2285,N_2231,N_2219);
and U2286 (N_2286,N_2218,N_2214);
nand U2287 (N_2287,N_2230,N_2243);
or U2288 (N_2288,N_2233,N_2201);
nor U2289 (N_2289,N_2206,N_2232);
and U2290 (N_2290,N_2217,N_2222);
nor U2291 (N_2291,N_2211,N_2216);
nor U2292 (N_2292,N_2232,N_2215);
nor U2293 (N_2293,N_2205,N_2206);
and U2294 (N_2294,N_2248,N_2231);
nor U2295 (N_2295,N_2244,N_2209);
nand U2296 (N_2296,N_2213,N_2223);
nor U2297 (N_2297,N_2235,N_2248);
nand U2298 (N_2298,N_2214,N_2228);
nor U2299 (N_2299,N_2200,N_2209);
and U2300 (N_2300,N_2281,N_2280);
and U2301 (N_2301,N_2278,N_2268);
nand U2302 (N_2302,N_2266,N_2273);
nor U2303 (N_2303,N_2282,N_2299);
and U2304 (N_2304,N_2259,N_2292);
or U2305 (N_2305,N_2297,N_2291);
and U2306 (N_2306,N_2284,N_2261);
and U2307 (N_2307,N_2276,N_2262);
and U2308 (N_2308,N_2263,N_2285);
or U2309 (N_2309,N_2293,N_2250);
and U2310 (N_2310,N_2256,N_2253);
and U2311 (N_2311,N_2290,N_2251);
nor U2312 (N_2312,N_2286,N_2254);
or U2313 (N_2313,N_2277,N_2260);
or U2314 (N_2314,N_2272,N_2298);
nor U2315 (N_2315,N_2271,N_2274);
and U2316 (N_2316,N_2269,N_2296);
nor U2317 (N_2317,N_2257,N_2264);
and U2318 (N_2318,N_2289,N_2275);
nor U2319 (N_2319,N_2279,N_2283);
or U2320 (N_2320,N_2255,N_2252);
nor U2321 (N_2321,N_2265,N_2287);
nor U2322 (N_2322,N_2258,N_2295);
or U2323 (N_2323,N_2288,N_2294);
nand U2324 (N_2324,N_2267,N_2270);
and U2325 (N_2325,N_2288,N_2290);
nor U2326 (N_2326,N_2268,N_2259);
and U2327 (N_2327,N_2279,N_2297);
nor U2328 (N_2328,N_2274,N_2294);
nor U2329 (N_2329,N_2299,N_2290);
nor U2330 (N_2330,N_2254,N_2257);
nor U2331 (N_2331,N_2283,N_2276);
or U2332 (N_2332,N_2290,N_2252);
or U2333 (N_2333,N_2261,N_2272);
nor U2334 (N_2334,N_2280,N_2293);
and U2335 (N_2335,N_2271,N_2270);
nor U2336 (N_2336,N_2254,N_2269);
nor U2337 (N_2337,N_2281,N_2261);
or U2338 (N_2338,N_2274,N_2267);
nor U2339 (N_2339,N_2270,N_2258);
nand U2340 (N_2340,N_2268,N_2280);
nor U2341 (N_2341,N_2262,N_2290);
nand U2342 (N_2342,N_2273,N_2294);
or U2343 (N_2343,N_2257,N_2299);
nand U2344 (N_2344,N_2257,N_2280);
and U2345 (N_2345,N_2257,N_2258);
nand U2346 (N_2346,N_2279,N_2272);
nand U2347 (N_2347,N_2257,N_2290);
nor U2348 (N_2348,N_2296,N_2278);
or U2349 (N_2349,N_2274,N_2257);
nand U2350 (N_2350,N_2346,N_2337);
nand U2351 (N_2351,N_2340,N_2339);
or U2352 (N_2352,N_2348,N_2326);
nor U2353 (N_2353,N_2329,N_2328);
and U2354 (N_2354,N_2327,N_2336);
and U2355 (N_2355,N_2318,N_2322);
nor U2356 (N_2356,N_2311,N_2305);
nand U2357 (N_2357,N_2321,N_2308);
or U2358 (N_2358,N_2324,N_2341);
nor U2359 (N_2359,N_2343,N_2325);
nand U2360 (N_2360,N_2301,N_2320);
and U2361 (N_2361,N_2302,N_2314);
and U2362 (N_2362,N_2316,N_2317);
nor U2363 (N_2363,N_2319,N_2313);
or U2364 (N_2364,N_2310,N_2330);
nand U2365 (N_2365,N_2332,N_2331);
nor U2366 (N_2366,N_2304,N_2345);
xnor U2367 (N_2367,N_2333,N_2342);
and U2368 (N_2368,N_2323,N_2334);
nand U2369 (N_2369,N_2312,N_2307);
nand U2370 (N_2370,N_2315,N_2347);
nand U2371 (N_2371,N_2338,N_2303);
and U2372 (N_2372,N_2300,N_2309);
and U2373 (N_2373,N_2349,N_2306);
nand U2374 (N_2374,N_2344,N_2335);
and U2375 (N_2375,N_2303,N_2328);
nand U2376 (N_2376,N_2301,N_2321);
nor U2377 (N_2377,N_2315,N_2338);
nor U2378 (N_2378,N_2306,N_2330);
and U2379 (N_2379,N_2328,N_2302);
nor U2380 (N_2380,N_2320,N_2317);
or U2381 (N_2381,N_2341,N_2317);
nand U2382 (N_2382,N_2328,N_2341);
and U2383 (N_2383,N_2301,N_2342);
nand U2384 (N_2384,N_2322,N_2310);
nand U2385 (N_2385,N_2345,N_2301);
and U2386 (N_2386,N_2348,N_2310);
nand U2387 (N_2387,N_2345,N_2336);
or U2388 (N_2388,N_2308,N_2315);
nand U2389 (N_2389,N_2331,N_2339);
nand U2390 (N_2390,N_2347,N_2346);
nor U2391 (N_2391,N_2310,N_2328);
or U2392 (N_2392,N_2326,N_2322);
nand U2393 (N_2393,N_2335,N_2311);
and U2394 (N_2394,N_2345,N_2338);
or U2395 (N_2395,N_2326,N_2307);
or U2396 (N_2396,N_2334,N_2339);
or U2397 (N_2397,N_2314,N_2322);
and U2398 (N_2398,N_2301,N_2318);
nand U2399 (N_2399,N_2310,N_2312);
and U2400 (N_2400,N_2372,N_2378);
nand U2401 (N_2401,N_2374,N_2351);
and U2402 (N_2402,N_2356,N_2387);
or U2403 (N_2403,N_2399,N_2379);
or U2404 (N_2404,N_2382,N_2350);
or U2405 (N_2405,N_2363,N_2377);
and U2406 (N_2406,N_2380,N_2385);
or U2407 (N_2407,N_2355,N_2396);
and U2408 (N_2408,N_2373,N_2370);
nor U2409 (N_2409,N_2397,N_2389);
and U2410 (N_2410,N_2371,N_2392);
and U2411 (N_2411,N_2362,N_2354);
or U2412 (N_2412,N_2358,N_2376);
nor U2413 (N_2413,N_2384,N_2368);
or U2414 (N_2414,N_2357,N_2367);
and U2415 (N_2415,N_2360,N_2398);
or U2416 (N_2416,N_2395,N_2394);
and U2417 (N_2417,N_2353,N_2361);
or U2418 (N_2418,N_2365,N_2375);
nor U2419 (N_2419,N_2352,N_2366);
nor U2420 (N_2420,N_2369,N_2386);
or U2421 (N_2421,N_2388,N_2390);
or U2422 (N_2422,N_2383,N_2381);
nand U2423 (N_2423,N_2391,N_2364);
nand U2424 (N_2424,N_2359,N_2393);
xnor U2425 (N_2425,N_2370,N_2365);
nor U2426 (N_2426,N_2391,N_2359);
or U2427 (N_2427,N_2395,N_2351);
nor U2428 (N_2428,N_2380,N_2396);
and U2429 (N_2429,N_2399,N_2373);
nor U2430 (N_2430,N_2368,N_2395);
nor U2431 (N_2431,N_2366,N_2385);
or U2432 (N_2432,N_2380,N_2354);
nand U2433 (N_2433,N_2396,N_2357);
and U2434 (N_2434,N_2359,N_2378);
or U2435 (N_2435,N_2366,N_2380);
and U2436 (N_2436,N_2383,N_2356);
nor U2437 (N_2437,N_2366,N_2374);
nor U2438 (N_2438,N_2355,N_2390);
nand U2439 (N_2439,N_2366,N_2389);
or U2440 (N_2440,N_2386,N_2359);
nor U2441 (N_2441,N_2350,N_2387);
nand U2442 (N_2442,N_2392,N_2387);
nor U2443 (N_2443,N_2370,N_2353);
or U2444 (N_2444,N_2358,N_2351);
or U2445 (N_2445,N_2373,N_2351);
and U2446 (N_2446,N_2360,N_2371);
nand U2447 (N_2447,N_2373,N_2372);
and U2448 (N_2448,N_2396,N_2397);
or U2449 (N_2449,N_2376,N_2396);
and U2450 (N_2450,N_2436,N_2449);
nor U2451 (N_2451,N_2418,N_2440);
nor U2452 (N_2452,N_2432,N_2433);
nand U2453 (N_2453,N_2409,N_2447);
or U2454 (N_2454,N_2402,N_2419);
and U2455 (N_2455,N_2416,N_2417);
nand U2456 (N_2456,N_2438,N_2426);
and U2457 (N_2457,N_2405,N_2400);
or U2458 (N_2458,N_2431,N_2404);
nand U2459 (N_2459,N_2430,N_2434);
or U2460 (N_2460,N_2435,N_2415);
or U2461 (N_2461,N_2421,N_2424);
or U2462 (N_2462,N_2413,N_2411);
nor U2463 (N_2463,N_2443,N_2428);
nand U2464 (N_2464,N_2412,N_2403);
or U2465 (N_2465,N_2437,N_2425);
and U2466 (N_2466,N_2420,N_2448);
and U2467 (N_2467,N_2408,N_2410);
nor U2468 (N_2468,N_2423,N_2429);
and U2469 (N_2469,N_2444,N_2422);
nand U2470 (N_2470,N_2427,N_2439);
or U2471 (N_2471,N_2441,N_2406);
nor U2472 (N_2472,N_2407,N_2401);
nor U2473 (N_2473,N_2446,N_2445);
nand U2474 (N_2474,N_2442,N_2414);
or U2475 (N_2475,N_2441,N_2412);
nor U2476 (N_2476,N_2428,N_2420);
nand U2477 (N_2477,N_2414,N_2406);
or U2478 (N_2478,N_2431,N_2407);
nand U2479 (N_2479,N_2406,N_2428);
nand U2480 (N_2480,N_2449,N_2446);
nand U2481 (N_2481,N_2443,N_2407);
or U2482 (N_2482,N_2424,N_2402);
or U2483 (N_2483,N_2424,N_2401);
nor U2484 (N_2484,N_2428,N_2417);
nor U2485 (N_2485,N_2408,N_2449);
xnor U2486 (N_2486,N_2446,N_2436);
or U2487 (N_2487,N_2405,N_2436);
or U2488 (N_2488,N_2418,N_2405);
nor U2489 (N_2489,N_2442,N_2432);
or U2490 (N_2490,N_2423,N_2414);
or U2491 (N_2491,N_2420,N_2446);
nor U2492 (N_2492,N_2423,N_2405);
or U2493 (N_2493,N_2447,N_2438);
nand U2494 (N_2494,N_2416,N_2425);
and U2495 (N_2495,N_2432,N_2425);
and U2496 (N_2496,N_2433,N_2415);
and U2497 (N_2497,N_2445,N_2436);
and U2498 (N_2498,N_2443,N_2418);
nand U2499 (N_2499,N_2441,N_2431);
nand U2500 (N_2500,N_2454,N_2486);
nor U2501 (N_2501,N_2464,N_2466);
and U2502 (N_2502,N_2475,N_2489);
nand U2503 (N_2503,N_2460,N_2476);
nor U2504 (N_2504,N_2469,N_2480);
or U2505 (N_2505,N_2483,N_2479);
nand U2506 (N_2506,N_2491,N_2463);
nand U2507 (N_2507,N_2472,N_2496);
and U2508 (N_2508,N_2453,N_2473);
or U2509 (N_2509,N_2470,N_2456);
and U2510 (N_2510,N_2474,N_2492);
or U2511 (N_2511,N_2462,N_2488);
and U2512 (N_2512,N_2498,N_2451);
nor U2513 (N_2513,N_2484,N_2459);
xnor U2514 (N_2514,N_2471,N_2455);
nand U2515 (N_2515,N_2468,N_2494);
nand U2516 (N_2516,N_2478,N_2457);
nor U2517 (N_2517,N_2465,N_2490);
xnor U2518 (N_2518,N_2477,N_2450);
or U2519 (N_2519,N_2458,N_2497);
nor U2520 (N_2520,N_2481,N_2493);
nor U2521 (N_2521,N_2485,N_2452);
nand U2522 (N_2522,N_2499,N_2495);
nand U2523 (N_2523,N_2482,N_2487);
or U2524 (N_2524,N_2461,N_2467);
nand U2525 (N_2525,N_2487,N_2486);
nand U2526 (N_2526,N_2476,N_2472);
or U2527 (N_2527,N_2468,N_2471);
nor U2528 (N_2528,N_2491,N_2465);
and U2529 (N_2529,N_2487,N_2464);
nor U2530 (N_2530,N_2466,N_2490);
nor U2531 (N_2531,N_2484,N_2460);
or U2532 (N_2532,N_2489,N_2468);
nand U2533 (N_2533,N_2491,N_2481);
and U2534 (N_2534,N_2488,N_2493);
nand U2535 (N_2535,N_2471,N_2464);
and U2536 (N_2536,N_2451,N_2499);
or U2537 (N_2537,N_2459,N_2453);
nand U2538 (N_2538,N_2496,N_2461);
nand U2539 (N_2539,N_2495,N_2479);
and U2540 (N_2540,N_2460,N_2487);
nor U2541 (N_2541,N_2460,N_2481);
and U2542 (N_2542,N_2451,N_2476);
and U2543 (N_2543,N_2481,N_2466);
nor U2544 (N_2544,N_2460,N_2464);
nand U2545 (N_2545,N_2467,N_2494);
nand U2546 (N_2546,N_2469,N_2454);
or U2547 (N_2547,N_2471,N_2454);
or U2548 (N_2548,N_2450,N_2452);
or U2549 (N_2549,N_2496,N_2453);
nand U2550 (N_2550,N_2517,N_2523);
and U2551 (N_2551,N_2520,N_2505);
and U2552 (N_2552,N_2544,N_2525);
and U2553 (N_2553,N_2538,N_2501);
and U2554 (N_2554,N_2515,N_2542);
or U2555 (N_2555,N_2537,N_2531);
or U2556 (N_2556,N_2541,N_2522);
nand U2557 (N_2557,N_2530,N_2547);
nor U2558 (N_2558,N_2524,N_2518);
and U2559 (N_2559,N_2512,N_2514);
nor U2560 (N_2560,N_2511,N_2526);
nand U2561 (N_2561,N_2529,N_2506);
nand U2562 (N_2562,N_2548,N_2503);
and U2563 (N_2563,N_2508,N_2533);
nor U2564 (N_2564,N_2534,N_2507);
nor U2565 (N_2565,N_2504,N_2540);
or U2566 (N_2566,N_2549,N_2516);
nand U2567 (N_2567,N_2502,N_2510);
nand U2568 (N_2568,N_2521,N_2536);
and U2569 (N_2569,N_2500,N_2519);
and U2570 (N_2570,N_2539,N_2543);
nand U2571 (N_2571,N_2532,N_2546);
nand U2572 (N_2572,N_2545,N_2513);
nor U2573 (N_2573,N_2528,N_2509);
nand U2574 (N_2574,N_2527,N_2535);
nand U2575 (N_2575,N_2545,N_2501);
nand U2576 (N_2576,N_2500,N_2521);
and U2577 (N_2577,N_2508,N_2509);
nor U2578 (N_2578,N_2547,N_2544);
and U2579 (N_2579,N_2513,N_2527);
nand U2580 (N_2580,N_2535,N_2519);
nor U2581 (N_2581,N_2549,N_2509);
nor U2582 (N_2582,N_2534,N_2535);
nor U2583 (N_2583,N_2507,N_2506);
nand U2584 (N_2584,N_2536,N_2520);
and U2585 (N_2585,N_2530,N_2540);
and U2586 (N_2586,N_2546,N_2511);
and U2587 (N_2587,N_2547,N_2541);
and U2588 (N_2588,N_2521,N_2508);
nand U2589 (N_2589,N_2525,N_2518);
nor U2590 (N_2590,N_2540,N_2547);
or U2591 (N_2591,N_2535,N_2538);
or U2592 (N_2592,N_2516,N_2518);
nand U2593 (N_2593,N_2549,N_2540);
and U2594 (N_2594,N_2531,N_2547);
and U2595 (N_2595,N_2549,N_2512);
and U2596 (N_2596,N_2539,N_2525);
nor U2597 (N_2597,N_2522,N_2506);
nand U2598 (N_2598,N_2517,N_2514);
xor U2599 (N_2599,N_2503,N_2514);
or U2600 (N_2600,N_2598,N_2555);
nor U2601 (N_2601,N_2581,N_2573);
nand U2602 (N_2602,N_2595,N_2568);
nor U2603 (N_2603,N_2596,N_2556);
or U2604 (N_2604,N_2553,N_2561);
and U2605 (N_2605,N_2593,N_2574);
or U2606 (N_2606,N_2583,N_2551);
nor U2607 (N_2607,N_2591,N_2589);
nor U2608 (N_2608,N_2590,N_2571);
or U2609 (N_2609,N_2578,N_2576);
and U2610 (N_2610,N_2592,N_2588);
nand U2611 (N_2611,N_2569,N_2567);
or U2612 (N_2612,N_2565,N_2587);
and U2613 (N_2613,N_2550,N_2563);
nand U2614 (N_2614,N_2552,N_2597);
xor U2615 (N_2615,N_2562,N_2575);
nor U2616 (N_2616,N_2594,N_2585);
and U2617 (N_2617,N_2564,N_2557);
nand U2618 (N_2618,N_2577,N_2599);
nor U2619 (N_2619,N_2570,N_2580);
or U2620 (N_2620,N_2579,N_2554);
nand U2621 (N_2621,N_2560,N_2584);
nand U2622 (N_2622,N_2586,N_2558);
or U2623 (N_2623,N_2559,N_2582);
nand U2624 (N_2624,N_2572,N_2566);
or U2625 (N_2625,N_2581,N_2557);
or U2626 (N_2626,N_2563,N_2554);
or U2627 (N_2627,N_2555,N_2583);
or U2628 (N_2628,N_2597,N_2557);
nor U2629 (N_2629,N_2576,N_2598);
nand U2630 (N_2630,N_2579,N_2550);
nor U2631 (N_2631,N_2575,N_2593);
or U2632 (N_2632,N_2578,N_2588);
nand U2633 (N_2633,N_2556,N_2577);
or U2634 (N_2634,N_2579,N_2594);
nor U2635 (N_2635,N_2567,N_2568);
or U2636 (N_2636,N_2573,N_2568);
or U2637 (N_2637,N_2564,N_2593);
and U2638 (N_2638,N_2568,N_2557);
xor U2639 (N_2639,N_2596,N_2567);
or U2640 (N_2640,N_2577,N_2558);
nor U2641 (N_2641,N_2577,N_2567);
nor U2642 (N_2642,N_2596,N_2569);
nor U2643 (N_2643,N_2596,N_2564);
and U2644 (N_2644,N_2588,N_2594);
nor U2645 (N_2645,N_2589,N_2561);
or U2646 (N_2646,N_2555,N_2587);
and U2647 (N_2647,N_2553,N_2595);
nand U2648 (N_2648,N_2588,N_2564);
or U2649 (N_2649,N_2558,N_2569);
or U2650 (N_2650,N_2628,N_2622);
or U2651 (N_2651,N_2610,N_2640);
nor U2652 (N_2652,N_2649,N_2626);
nand U2653 (N_2653,N_2624,N_2637);
and U2654 (N_2654,N_2604,N_2642);
and U2655 (N_2655,N_2644,N_2639);
and U2656 (N_2656,N_2606,N_2630);
nand U2657 (N_2657,N_2625,N_2629);
nand U2658 (N_2658,N_2621,N_2620);
and U2659 (N_2659,N_2600,N_2633);
and U2660 (N_2660,N_2623,N_2612);
nor U2661 (N_2661,N_2609,N_2641);
nor U2662 (N_2662,N_2645,N_2607);
and U2663 (N_2663,N_2619,N_2605);
and U2664 (N_2664,N_2611,N_2648);
nand U2665 (N_2665,N_2627,N_2636);
or U2666 (N_2666,N_2608,N_2618);
and U2667 (N_2667,N_2602,N_2643);
and U2668 (N_2668,N_2615,N_2647);
or U2669 (N_2669,N_2601,N_2634);
or U2670 (N_2670,N_2632,N_2631);
or U2671 (N_2671,N_2603,N_2613);
or U2672 (N_2672,N_2635,N_2614);
or U2673 (N_2673,N_2617,N_2638);
or U2674 (N_2674,N_2646,N_2616);
nor U2675 (N_2675,N_2608,N_2625);
or U2676 (N_2676,N_2640,N_2643);
nor U2677 (N_2677,N_2607,N_2647);
nand U2678 (N_2678,N_2646,N_2628);
nand U2679 (N_2679,N_2608,N_2642);
or U2680 (N_2680,N_2613,N_2628);
or U2681 (N_2681,N_2633,N_2632);
nand U2682 (N_2682,N_2649,N_2601);
and U2683 (N_2683,N_2623,N_2649);
nor U2684 (N_2684,N_2635,N_2645);
nor U2685 (N_2685,N_2645,N_2637);
xnor U2686 (N_2686,N_2613,N_2602);
and U2687 (N_2687,N_2600,N_2631);
and U2688 (N_2688,N_2604,N_2601);
nand U2689 (N_2689,N_2608,N_2607);
or U2690 (N_2690,N_2632,N_2613);
nor U2691 (N_2691,N_2602,N_2610);
nor U2692 (N_2692,N_2630,N_2632);
and U2693 (N_2693,N_2608,N_2633);
or U2694 (N_2694,N_2601,N_2628);
or U2695 (N_2695,N_2621,N_2619);
and U2696 (N_2696,N_2630,N_2616);
and U2697 (N_2697,N_2636,N_2648);
nand U2698 (N_2698,N_2618,N_2601);
or U2699 (N_2699,N_2606,N_2645);
or U2700 (N_2700,N_2673,N_2678);
or U2701 (N_2701,N_2684,N_2662);
nand U2702 (N_2702,N_2674,N_2659);
or U2703 (N_2703,N_2685,N_2661);
nor U2704 (N_2704,N_2698,N_2671);
and U2705 (N_2705,N_2664,N_2682);
nand U2706 (N_2706,N_2692,N_2690);
or U2707 (N_2707,N_2669,N_2694);
and U2708 (N_2708,N_2696,N_2670);
nor U2709 (N_2709,N_2655,N_2687);
and U2710 (N_2710,N_2667,N_2653);
nand U2711 (N_2711,N_2666,N_2660);
nand U2712 (N_2712,N_2681,N_2657);
and U2713 (N_2713,N_2677,N_2680);
nand U2714 (N_2714,N_2658,N_2676);
and U2715 (N_2715,N_2679,N_2672);
or U2716 (N_2716,N_2654,N_2691);
nor U2717 (N_2717,N_2686,N_2663);
or U2718 (N_2718,N_2651,N_2683);
nor U2719 (N_2719,N_2656,N_2695);
or U2720 (N_2720,N_2688,N_2693);
and U2721 (N_2721,N_2650,N_2675);
nand U2722 (N_2722,N_2665,N_2699);
and U2723 (N_2723,N_2697,N_2652);
and U2724 (N_2724,N_2689,N_2668);
and U2725 (N_2725,N_2663,N_2691);
nand U2726 (N_2726,N_2650,N_2662);
nand U2727 (N_2727,N_2663,N_2653);
or U2728 (N_2728,N_2679,N_2674);
nand U2729 (N_2729,N_2667,N_2663);
nor U2730 (N_2730,N_2651,N_2680);
or U2731 (N_2731,N_2698,N_2653);
nor U2732 (N_2732,N_2670,N_2685);
nor U2733 (N_2733,N_2673,N_2692);
nor U2734 (N_2734,N_2677,N_2661);
and U2735 (N_2735,N_2693,N_2655);
nand U2736 (N_2736,N_2661,N_2652);
or U2737 (N_2737,N_2688,N_2666);
nand U2738 (N_2738,N_2679,N_2651);
and U2739 (N_2739,N_2654,N_2672);
nand U2740 (N_2740,N_2652,N_2654);
nand U2741 (N_2741,N_2650,N_2673);
or U2742 (N_2742,N_2676,N_2689);
nor U2743 (N_2743,N_2660,N_2685);
nor U2744 (N_2744,N_2666,N_2675);
nor U2745 (N_2745,N_2694,N_2697);
nor U2746 (N_2746,N_2690,N_2687);
and U2747 (N_2747,N_2676,N_2673);
nand U2748 (N_2748,N_2654,N_2694);
nand U2749 (N_2749,N_2674,N_2699);
and U2750 (N_2750,N_2744,N_2738);
nor U2751 (N_2751,N_2700,N_2733);
or U2752 (N_2752,N_2710,N_2747);
nand U2753 (N_2753,N_2701,N_2702);
nand U2754 (N_2754,N_2711,N_2723);
nor U2755 (N_2755,N_2734,N_2718);
or U2756 (N_2756,N_2729,N_2748);
nor U2757 (N_2757,N_2730,N_2714);
nor U2758 (N_2758,N_2713,N_2724);
nor U2759 (N_2759,N_2749,N_2703);
and U2760 (N_2760,N_2708,N_2709);
nand U2761 (N_2761,N_2719,N_2715);
nor U2762 (N_2762,N_2743,N_2727);
nand U2763 (N_2763,N_2705,N_2725);
nand U2764 (N_2764,N_2740,N_2717);
nand U2765 (N_2765,N_2722,N_2735);
nand U2766 (N_2766,N_2716,N_2721);
nand U2767 (N_2767,N_2739,N_2746);
or U2768 (N_2768,N_2741,N_2731);
and U2769 (N_2769,N_2745,N_2726);
and U2770 (N_2770,N_2712,N_2706);
and U2771 (N_2771,N_2737,N_2728);
nand U2772 (N_2772,N_2707,N_2742);
or U2773 (N_2773,N_2720,N_2732);
and U2774 (N_2774,N_2704,N_2736);
nand U2775 (N_2775,N_2709,N_2744);
nor U2776 (N_2776,N_2733,N_2717);
nand U2777 (N_2777,N_2702,N_2719);
and U2778 (N_2778,N_2716,N_2734);
or U2779 (N_2779,N_2701,N_2735);
and U2780 (N_2780,N_2718,N_2728);
or U2781 (N_2781,N_2741,N_2701);
and U2782 (N_2782,N_2745,N_2742);
and U2783 (N_2783,N_2720,N_2748);
nor U2784 (N_2784,N_2730,N_2707);
nor U2785 (N_2785,N_2705,N_2704);
nor U2786 (N_2786,N_2730,N_2725);
nor U2787 (N_2787,N_2721,N_2732);
nand U2788 (N_2788,N_2717,N_2732);
and U2789 (N_2789,N_2703,N_2707);
nand U2790 (N_2790,N_2716,N_2726);
nor U2791 (N_2791,N_2701,N_2737);
nand U2792 (N_2792,N_2704,N_2735);
nand U2793 (N_2793,N_2746,N_2727);
nand U2794 (N_2794,N_2748,N_2734);
nand U2795 (N_2795,N_2745,N_2703);
and U2796 (N_2796,N_2709,N_2736);
nor U2797 (N_2797,N_2703,N_2710);
nand U2798 (N_2798,N_2738,N_2709);
and U2799 (N_2799,N_2709,N_2734);
nand U2800 (N_2800,N_2775,N_2770);
or U2801 (N_2801,N_2789,N_2756);
nand U2802 (N_2802,N_2779,N_2799);
nand U2803 (N_2803,N_2752,N_2785);
or U2804 (N_2804,N_2768,N_2766);
and U2805 (N_2805,N_2776,N_2762);
or U2806 (N_2806,N_2753,N_2798);
and U2807 (N_2807,N_2781,N_2788);
or U2808 (N_2808,N_2755,N_2771);
nor U2809 (N_2809,N_2786,N_2751);
and U2810 (N_2810,N_2764,N_2760);
and U2811 (N_2811,N_2782,N_2797);
and U2812 (N_2812,N_2793,N_2783);
and U2813 (N_2813,N_2790,N_2774);
and U2814 (N_2814,N_2794,N_2763);
and U2815 (N_2815,N_2795,N_2777);
nor U2816 (N_2816,N_2792,N_2780);
nor U2817 (N_2817,N_2758,N_2796);
nand U2818 (N_2818,N_2750,N_2772);
nor U2819 (N_2819,N_2767,N_2757);
nor U2820 (N_2820,N_2787,N_2754);
or U2821 (N_2821,N_2765,N_2778);
nor U2822 (N_2822,N_2769,N_2759);
and U2823 (N_2823,N_2791,N_2773);
nor U2824 (N_2824,N_2761,N_2784);
nand U2825 (N_2825,N_2753,N_2796);
nor U2826 (N_2826,N_2763,N_2778);
and U2827 (N_2827,N_2796,N_2776);
xnor U2828 (N_2828,N_2798,N_2775);
nand U2829 (N_2829,N_2790,N_2787);
nand U2830 (N_2830,N_2752,N_2759);
and U2831 (N_2831,N_2790,N_2770);
or U2832 (N_2832,N_2785,N_2797);
nand U2833 (N_2833,N_2775,N_2769);
or U2834 (N_2834,N_2752,N_2767);
nand U2835 (N_2835,N_2776,N_2760);
or U2836 (N_2836,N_2786,N_2761);
or U2837 (N_2837,N_2781,N_2784);
and U2838 (N_2838,N_2782,N_2765);
nand U2839 (N_2839,N_2798,N_2792);
or U2840 (N_2840,N_2798,N_2793);
and U2841 (N_2841,N_2782,N_2774);
nor U2842 (N_2842,N_2771,N_2798);
nor U2843 (N_2843,N_2795,N_2760);
nor U2844 (N_2844,N_2768,N_2772);
nor U2845 (N_2845,N_2767,N_2783);
or U2846 (N_2846,N_2768,N_2785);
nand U2847 (N_2847,N_2758,N_2779);
nor U2848 (N_2848,N_2751,N_2770);
nor U2849 (N_2849,N_2776,N_2754);
or U2850 (N_2850,N_2810,N_2808);
and U2851 (N_2851,N_2838,N_2805);
or U2852 (N_2852,N_2803,N_2849);
nand U2853 (N_2853,N_2837,N_2840);
or U2854 (N_2854,N_2831,N_2846);
nand U2855 (N_2855,N_2845,N_2824);
and U2856 (N_2856,N_2832,N_2817);
or U2857 (N_2857,N_2827,N_2842);
and U2858 (N_2858,N_2844,N_2826);
nand U2859 (N_2859,N_2836,N_2847);
or U2860 (N_2860,N_2834,N_2800);
nand U2861 (N_2861,N_2801,N_2828);
and U2862 (N_2862,N_2811,N_2839);
and U2863 (N_2863,N_2802,N_2835);
and U2864 (N_2864,N_2816,N_2833);
nor U2865 (N_2865,N_2815,N_2825);
nor U2866 (N_2866,N_2812,N_2804);
and U2867 (N_2867,N_2814,N_2813);
or U2868 (N_2868,N_2819,N_2843);
nand U2869 (N_2869,N_2830,N_2820);
nor U2870 (N_2870,N_2822,N_2829);
nor U2871 (N_2871,N_2809,N_2848);
or U2872 (N_2872,N_2818,N_2821);
or U2873 (N_2873,N_2806,N_2823);
xor U2874 (N_2874,N_2807,N_2841);
nand U2875 (N_2875,N_2809,N_2841);
and U2876 (N_2876,N_2821,N_2815);
nor U2877 (N_2877,N_2816,N_2802);
nor U2878 (N_2878,N_2832,N_2811);
and U2879 (N_2879,N_2815,N_2832);
or U2880 (N_2880,N_2830,N_2802);
or U2881 (N_2881,N_2804,N_2846);
and U2882 (N_2882,N_2820,N_2829);
or U2883 (N_2883,N_2844,N_2831);
nand U2884 (N_2884,N_2825,N_2807);
nor U2885 (N_2885,N_2805,N_2828);
and U2886 (N_2886,N_2813,N_2832);
or U2887 (N_2887,N_2815,N_2826);
nor U2888 (N_2888,N_2816,N_2827);
or U2889 (N_2889,N_2811,N_2825);
or U2890 (N_2890,N_2829,N_2838);
or U2891 (N_2891,N_2837,N_2810);
nand U2892 (N_2892,N_2830,N_2807);
nand U2893 (N_2893,N_2803,N_2843);
nor U2894 (N_2894,N_2842,N_2826);
nor U2895 (N_2895,N_2822,N_2832);
or U2896 (N_2896,N_2826,N_2823);
and U2897 (N_2897,N_2818,N_2808);
nand U2898 (N_2898,N_2823,N_2814);
or U2899 (N_2899,N_2846,N_2836);
nand U2900 (N_2900,N_2885,N_2858);
and U2901 (N_2901,N_2894,N_2864);
nor U2902 (N_2902,N_2855,N_2867);
and U2903 (N_2903,N_2859,N_2897);
nor U2904 (N_2904,N_2883,N_2876);
and U2905 (N_2905,N_2880,N_2887);
nor U2906 (N_2906,N_2875,N_2856);
nand U2907 (N_2907,N_2892,N_2890);
nor U2908 (N_2908,N_2853,N_2854);
or U2909 (N_2909,N_2857,N_2889);
and U2910 (N_2910,N_2871,N_2868);
and U2911 (N_2911,N_2895,N_2882);
or U2912 (N_2912,N_2869,N_2879);
and U2913 (N_2913,N_2881,N_2873);
nand U2914 (N_2914,N_2872,N_2893);
or U2915 (N_2915,N_2888,N_2865);
and U2916 (N_2916,N_2898,N_2863);
nor U2917 (N_2917,N_2850,N_2870);
nor U2918 (N_2918,N_2866,N_2852);
nand U2919 (N_2919,N_2886,N_2891);
nor U2920 (N_2920,N_2896,N_2877);
nor U2921 (N_2921,N_2861,N_2860);
nand U2922 (N_2922,N_2884,N_2862);
and U2923 (N_2923,N_2899,N_2878);
or U2924 (N_2924,N_2851,N_2874);
nor U2925 (N_2925,N_2889,N_2871);
and U2926 (N_2926,N_2887,N_2889);
and U2927 (N_2927,N_2851,N_2865);
xor U2928 (N_2928,N_2868,N_2864);
nand U2929 (N_2929,N_2878,N_2852);
or U2930 (N_2930,N_2878,N_2870);
nand U2931 (N_2931,N_2856,N_2869);
nand U2932 (N_2932,N_2870,N_2857);
or U2933 (N_2933,N_2862,N_2855);
nand U2934 (N_2934,N_2887,N_2868);
and U2935 (N_2935,N_2874,N_2894);
nor U2936 (N_2936,N_2861,N_2890);
and U2937 (N_2937,N_2879,N_2880);
xnor U2938 (N_2938,N_2891,N_2893);
or U2939 (N_2939,N_2884,N_2887);
and U2940 (N_2940,N_2874,N_2852);
or U2941 (N_2941,N_2863,N_2887);
or U2942 (N_2942,N_2863,N_2879);
and U2943 (N_2943,N_2879,N_2893);
nand U2944 (N_2944,N_2886,N_2862);
nand U2945 (N_2945,N_2883,N_2894);
or U2946 (N_2946,N_2891,N_2862);
nand U2947 (N_2947,N_2895,N_2894);
nand U2948 (N_2948,N_2870,N_2893);
nor U2949 (N_2949,N_2862,N_2871);
or U2950 (N_2950,N_2922,N_2900);
nor U2951 (N_2951,N_2940,N_2933);
and U2952 (N_2952,N_2929,N_2930);
nand U2953 (N_2953,N_2947,N_2918);
or U2954 (N_2954,N_2919,N_2909);
nand U2955 (N_2955,N_2901,N_2908);
nor U2956 (N_2956,N_2906,N_2935);
and U2957 (N_2957,N_2915,N_2938);
or U2958 (N_2958,N_2921,N_2932);
nor U2959 (N_2959,N_2902,N_2946);
nor U2960 (N_2960,N_2907,N_2936);
or U2961 (N_2961,N_2903,N_2911);
or U2962 (N_2962,N_2904,N_2905);
or U2963 (N_2963,N_2934,N_2913);
and U2964 (N_2964,N_2948,N_2920);
and U2965 (N_2965,N_2928,N_2925);
nand U2966 (N_2966,N_2914,N_2944);
and U2967 (N_2967,N_2916,N_2942);
and U2968 (N_2968,N_2910,N_2943);
or U2969 (N_2969,N_2912,N_2945);
nand U2970 (N_2970,N_2949,N_2937);
or U2971 (N_2971,N_2931,N_2927);
nand U2972 (N_2972,N_2924,N_2917);
nand U2973 (N_2973,N_2939,N_2926);
nor U2974 (N_2974,N_2923,N_2941);
nand U2975 (N_2975,N_2918,N_2941);
and U2976 (N_2976,N_2935,N_2902);
and U2977 (N_2977,N_2904,N_2910);
nor U2978 (N_2978,N_2913,N_2941);
nor U2979 (N_2979,N_2902,N_2918);
and U2980 (N_2980,N_2933,N_2936);
nand U2981 (N_2981,N_2931,N_2937);
or U2982 (N_2982,N_2929,N_2916);
and U2983 (N_2983,N_2938,N_2928);
or U2984 (N_2984,N_2903,N_2914);
and U2985 (N_2985,N_2928,N_2936);
nor U2986 (N_2986,N_2941,N_2921);
nor U2987 (N_2987,N_2915,N_2945);
and U2988 (N_2988,N_2907,N_2908);
nor U2989 (N_2989,N_2935,N_2933);
nand U2990 (N_2990,N_2921,N_2906);
and U2991 (N_2991,N_2912,N_2913);
and U2992 (N_2992,N_2910,N_2906);
nor U2993 (N_2993,N_2905,N_2914);
nand U2994 (N_2994,N_2938,N_2931);
or U2995 (N_2995,N_2914,N_2937);
and U2996 (N_2996,N_2935,N_2934);
nand U2997 (N_2997,N_2915,N_2912);
and U2998 (N_2998,N_2924,N_2949);
nor U2999 (N_2999,N_2922,N_2943);
and UO_0 (O_0,N_2975,N_2985);
and UO_1 (O_1,N_2953,N_2957);
and UO_2 (O_2,N_2964,N_2963);
or UO_3 (O_3,N_2955,N_2988);
nor UO_4 (O_4,N_2970,N_2979);
or UO_5 (O_5,N_2973,N_2976);
or UO_6 (O_6,N_2965,N_2997);
or UO_7 (O_7,N_2998,N_2961);
or UO_8 (O_8,N_2994,N_2983);
and UO_9 (O_9,N_2967,N_2977);
nor UO_10 (O_10,N_2950,N_2972);
or UO_11 (O_11,N_2959,N_2992);
nor UO_12 (O_12,N_2952,N_2991);
or UO_13 (O_13,N_2990,N_2999);
nor UO_14 (O_14,N_2989,N_2987);
nand UO_15 (O_15,N_2993,N_2982);
and UO_16 (O_16,N_2966,N_2971);
nor UO_17 (O_17,N_2954,N_2995);
and UO_18 (O_18,N_2980,N_2981);
or UO_19 (O_19,N_2960,N_2996);
or UO_20 (O_20,N_2974,N_2986);
and UO_21 (O_21,N_2962,N_2958);
and UO_22 (O_22,N_2978,N_2951);
or UO_23 (O_23,N_2969,N_2984);
nor UO_24 (O_24,N_2956,N_2968);
and UO_25 (O_25,N_2956,N_2996);
nor UO_26 (O_26,N_2971,N_2995);
and UO_27 (O_27,N_2999,N_2986);
nor UO_28 (O_28,N_2973,N_2951);
nor UO_29 (O_29,N_2973,N_2950);
nand UO_30 (O_30,N_2966,N_2984);
nor UO_31 (O_31,N_2984,N_2960);
or UO_32 (O_32,N_2979,N_2950);
or UO_33 (O_33,N_2976,N_2965);
or UO_34 (O_34,N_2959,N_2981);
and UO_35 (O_35,N_2957,N_2992);
or UO_36 (O_36,N_2969,N_2996);
nand UO_37 (O_37,N_2979,N_2975);
and UO_38 (O_38,N_2977,N_2958);
or UO_39 (O_39,N_2998,N_2968);
xnor UO_40 (O_40,N_2999,N_2989);
and UO_41 (O_41,N_2998,N_2982);
nand UO_42 (O_42,N_2961,N_2983);
and UO_43 (O_43,N_2955,N_2964);
nor UO_44 (O_44,N_2977,N_2974);
and UO_45 (O_45,N_2955,N_2999);
nor UO_46 (O_46,N_2968,N_2962);
or UO_47 (O_47,N_2966,N_2954);
nor UO_48 (O_48,N_2971,N_2955);
nand UO_49 (O_49,N_2956,N_2960);
or UO_50 (O_50,N_2966,N_2980);
or UO_51 (O_51,N_2974,N_2992);
nand UO_52 (O_52,N_2975,N_2967);
and UO_53 (O_53,N_2990,N_2957);
or UO_54 (O_54,N_2970,N_2998);
nor UO_55 (O_55,N_2966,N_2961);
nor UO_56 (O_56,N_2981,N_2975);
and UO_57 (O_57,N_2961,N_2956);
and UO_58 (O_58,N_2992,N_2953);
nand UO_59 (O_59,N_2956,N_2950);
or UO_60 (O_60,N_2973,N_2989);
nand UO_61 (O_61,N_2980,N_2952);
and UO_62 (O_62,N_2977,N_2953);
nor UO_63 (O_63,N_2962,N_2985);
nor UO_64 (O_64,N_2992,N_2989);
and UO_65 (O_65,N_2973,N_2966);
nand UO_66 (O_66,N_2958,N_2971);
nand UO_67 (O_67,N_2993,N_2961);
or UO_68 (O_68,N_2970,N_2957);
nor UO_69 (O_69,N_2990,N_2966);
nor UO_70 (O_70,N_2997,N_2958);
nor UO_71 (O_71,N_2985,N_2973);
or UO_72 (O_72,N_2979,N_2963);
and UO_73 (O_73,N_2956,N_2977);
nand UO_74 (O_74,N_2973,N_2978);
and UO_75 (O_75,N_2980,N_2950);
nor UO_76 (O_76,N_2998,N_2992);
nand UO_77 (O_77,N_2950,N_2970);
or UO_78 (O_78,N_2992,N_2977);
or UO_79 (O_79,N_2986,N_2973);
and UO_80 (O_80,N_2996,N_2953);
nand UO_81 (O_81,N_2995,N_2984);
nand UO_82 (O_82,N_2965,N_2950);
nand UO_83 (O_83,N_2986,N_2963);
nand UO_84 (O_84,N_2965,N_2958);
nor UO_85 (O_85,N_2986,N_2956);
and UO_86 (O_86,N_2987,N_2999);
or UO_87 (O_87,N_2983,N_2966);
nand UO_88 (O_88,N_2970,N_2976);
or UO_89 (O_89,N_2970,N_2985);
nand UO_90 (O_90,N_2964,N_2956);
or UO_91 (O_91,N_2966,N_2987);
or UO_92 (O_92,N_2987,N_2988);
or UO_93 (O_93,N_2978,N_2970);
and UO_94 (O_94,N_2977,N_2962);
nand UO_95 (O_95,N_2966,N_2957);
or UO_96 (O_96,N_2966,N_2993);
and UO_97 (O_97,N_2992,N_2978);
nand UO_98 (O_98,N_2981,N_2970);
nand UO_99 (O_99,N_2984,N_2950);
or UO_100 (O_100,N_2961,N_2977);
nand UO_101 (O_101,N_2988,N_2980);
nand UO_102 (O_102,N_2950,N_2963);
nor UO_103 (O_103,N_2971,N_2960);
nor UO_104 (O_104,N_2962,N_2991);
and UO_105 (O_105,N_2980,N_2985);
nor UO_106 (O_106,N_2995,N_2968);
nand UO_107 (O_107,N_2950,N_2969);
nand UO_108 (O_108,N_2990,N_2998);
nand UO_109 (O_109,N_2984,N_2952);
and UO_110 (O_110,N_2953,N_2981);
or UO_111 (O_111,N_2958,N_2999);
nand UO_112 (O_112,N_2955,N_2986);
nand UO_113 (O_113,N_2977,N_2998);
or UO_114 (O_114,N_2999,N_2975);
and UO_115 (O_115,N_2951,N_2996);
nor UO_116 (O_116,N_2972,N_2994);
or UO_117 (O_117,N_2981,N_2963);
and UO_118 (O_118,N_2997,N_2964);
and UO_119 (O_119,N_2979,N_2968);
nand UO_120 (O_120,N_2987,N_2953);
or UO_121 (O_121,N_2988,N_2951);
nor UO_122 (O_122,N_2995,N_2958);
nand UO_123 (O_123,N_2979,N_2982);
nand UO_124 (O_124,N_2988,N_2974);
nand UO_125 (O_125,N_2957,N_2981);
xor UO_126 (O_126,N_2955,N_2994);
nor UO_127 (O_127,N_2969,N_2988);
and UO_128 (O_128,N_2990,N_2975);
and UO_129 (O_129,N_2998,N_2962);
or UO_130 (O_130,N_2974,N_2952);
or UO_131 (O_131,N_2951,N_2966);
or UO_132 (O_132,N_2973,N_2999);
nor UO_133 (O_133,N_2967,N_2953);
and UO_134 (O_134,N_2952,N_2961);
and UO_135 (O_135,N_2982,N_2975);
or UO_136 (O_136,N_2959,N_2989);
nand UO_137 (O_137,N_2952,N_2975);
or UO_138 (O_138,N_2986,N_2977);
nor UO_139 (O_139,N_2989,N_2958);
nand UO_140 (O_140,N_2985,N_2995);
nand UO_141 (O_141,N_2989,N_2978);
and UO_142 (O_142,N_2984,N_2989);
or UO_143 (O_143,N_2977,N_2972);
nand UO_144 (O_144,N_2983,N_2974);
and UO_145 (O_145,N_2994,N_2974);
and UO_146 (O_146,N_2970,N_2974);
nor UO_147 (O_147,N_2970,N_2952);
nor UO_148 (O_148,N_2961,N_2978);
nor UO_149 (O_149,N_2950,N_2978);
and UO_150 (O_150,N_2981,N_2974);
and UO_151 (O_151,N_2996,N_2973);
xor UO_152 (O_152,N_2997,N_2968);
nand UO_153 (O_153,N_2990,N_2961);
and UO_154 (O_154,N_2973,N_2982);
or UO_155 (O_155,N_2983,N_2968);
or UO_156 (O_156,N_2950,N_2988);
nand UO_157 (O_157,N_2957,N_2954);
and UO_158 (O_158,N_2995,N_2992);
and UO_159 (O_159,N_2995,N_2961);
and UO_160 (O_160,N_2964,N_2960);
nor UO_161 (O_161,N_2963,N_2983);
or UO_162 (O_162,N_2974,N_2954);
nand UO_163 (O_163,N_2974,N_2985);
nand UO_164 (O_164,N_2985,N_2967);
and UO_165 (O_165,N_2977,N_2951);
and UO_166 (O_166,N_2950,N_2986);
and UO_167 (O_167,N_2990,N_2962);
nor UO_168 (O_168,N_2998,N_2975);
and UO_169 (O_169,N_2976,N_2986);
or UO_170 (O_170,N_2994,N_2981);
nand UO_171 (O_171,N_2953,N_2994);
xnor UO_172 (O_172,N_2978,N_2952);
or UO_173 (O_173,N_2986,N_2972);
and UO_174 (O_174,N_2984,N_2978);
and UO_175 (O_175,N_2974,N_2966);
or UO_176 (O_176,N_2957,N_2955);
nor UO_177 (O_177,N_2954,N_2975);
and UO_178 (O_178,N_2983,N_2989);
and UO_179 (O_179,N_2977,N_2997);
nor UO_180 (O_180,N_2952,N_2979);
or UO_181 (O_181,N_2980,N_2955);
nor UO_182 (O_182,N_2967,N_2970);
nand UO_183 (O_183,N_2989,N_2971);
or UO_184 (O_184,N_2979,N_2989);
and UO_185 (O_185,N_2953,N_2986);
or UO_186 (O_186,N_2953,N_2963);
nand UO_187 (O_187,N_2991,N_2978);
nor UO_188 (O_188,N_2986,N_2991);
nor UO_189 (O_189,N_2983,N_2960);
and UO_190 (O_190,N_2985,N_2956);
and UO_191 (O_191,N_2961,N_2980);
and UO_192 (O_192,N_2981,N_2997);
nand UO_193 (O_193,N_2958,N_2969);
nand UO_194 (O_194,N_2956,N_2980);
nand UO_195 (O_195,N_2985,N_2996);
nand UO_196 (O_196,N_2953,N_2991);
nand UO_197 (O_197,N_2952,N_2992);
and UO_198 (O_198,N_2950,N_2953);
or UO_199 (O_199,N_2951,N_2983);
nand UO_200 (O_200,N_2955,N_2969);
nor UO_201 (O_201,N_2952,N_2983);
or UO_202 (O_202,N_2998,N_2969);
nor UO_203 (O_203,N_2958,N_2973);
nor UO_204 (O_204,N_2961,N_2958);
xor UO_205 (O_205,N_2959,N_2977);
nand UO_206 (O_206,N_2973,N_2967);
or UO_207 (O_207,N_2997,N_2974);
nand UO_208 (O_208,N_2979,N_2955);
nor UO_209 (O_209,N_2975,N_2980);
nand UO_210 (O_210,N_2969,N_2962);
or UO_211 (O_211,N_2985,N_2981);
nand UO_212 (O_212,N_2999,N_2968);
nand UO_213 (O_213,N_2983,N_2992);
nand UO_214 (O_214,N_2981,N_2950);
nor UO_215 (O_215,N_2976,N_2984);
and UO_216 (O_216,N_2955,N_2950);
or UO_217 (O_217,N_2986,N_2970);
nor UO_218 (O_218,N_2952,N_2971);
and UO_219 (O_219,N_2974,N_2995);
nor UO_220 (O_220,N_2983,N_2965);
and UO_221 (O_221,N_2977,N_2981);
nand UO_222 (O_222,N_2971,N_2984);
nand UO_223 (O_223,N_2985,N_2961);
nor UO_224 (O_224,N_2991,N_2993);
or UO_225 (O_225,N_2960,N_2992);
and UO_226 (O_226,N_2976,N_2991);
or UO_227 (O_227,N_2996,N_2977);
or UO_228 (O_228,N_2984,N_2983);
nand UO_229 (O_229,N_2985,N_2994);
and UO_230 (O_230,N_2978,N_2993);
and UO_231 (O_231,N_2956,N_2984);
and UO_232 (O_232,N_2990,N_2969);
nor UO_233 (O_233,N_2961,N_2987);
or UO_234 (O_234,N_2983,N_2954);
and UO_235 (O_235,N_2976,N_2985);
nand UO_236 (O_236,N_2960,N_2967);
and UO_237 (O_237,N_2988,N_2996);
and UO_238 (O_238,N_2967,N_2956);
nor UO_239 (O_239,N_2961,N_2972);
or UO_240 (O_240,N_2991,N_2971);
nand UO_241 (O_241,N_2998,N_2965);
nand UO_242 (O_242,N_2969,N_2989);
nand UO_243 (O_243,N_2995,N_2997);
nor UO_244 (O_244,N_2959,N_2979);
nor UO_245 (O_245,N_2992,N_2985);
or UO_246 (O_246,N_2991,N_2980);
or UO_247 (O_247,N_2984,N_2994);
or UO_248 (O_248,N_2963,N_2975);
nand UO_249 (O_249,N_2979,N_2966);
nor UO_250 (O_250,N_2995,N_2991);
nand UO_251 (O_251,N_2965,N_2957);
nand UO_252 (O_252,N_2988,N_2986);
nor UO_253 (O_253,N_2959,N_2966);
or UO_254 (O_254,N_2957,N_2973);
or UO_255 (O_255,N_2991,N_2988);
and UO_256 (O_256,N_2987,N_2967);
and UO_257 (O_257,N_2980,N_2957);
or UO_258 (O_258,N_2971,N_2987);
and UO_259 (O_259,N_2989,N_2962);
or UO_260 (O_260,N_2983,N_2973);
or UO_261 (O_261,N_2980,N_2998);
nand UO_262 (O_262,N_2961,N_2970);
or UO_263 (O_263,N_2992,N_2971);
and UO_264 (O_264,N_2999,N_2957);
and UO_265 (O_265,N_2987,N_2959);
and UO_266 (O_266,N_2955,N_2990);
nand UO_267 (O_267,N_2978,N_2976);
nand UO_268 (O_268,N_2987,N_2996);
or UO_269 (O_269,N_2966,N_2989);
nand UO_270 (O_270,N_2986,N_2985);
nor UO_271 (O_271,N_2998,N_2954);
and UO_272 (O_272,N_2997,N_2982);
nand UO_273 (O_273,N_2966,N_2995);
nand UO_274 (O_274,N_2976,N_2975);
nor UO_275 (O_275,N_2985,N_2951);
nor UO_276 (O_276,N_2951,N_2956);
or UO_277 (O_277,N_2951,N_2998);
and UO_278 (O_278,N_2982,N_2955);
nor UO_279 (O_279,N_2968,N_2951);
nor UO_280 (O_280,N_2955,N_2978);
or UO_281 (O_281,N_2994,N_2992);
or UO_282 (O_282,N_2955,N_2977);
nor UO_283 (O_283,N_2980,N_2977);
nor UO_284 (O_284,N_2966,N_2978);
and UO_285 (O_285,N_2956,N_2952);
nand UO_286 (O_286,N_2971,N_2964);
and UO_287 (O_287,N_2966,N_2953);
nand UO_288 (O_288,N_2954,N_2956);
nor UO_289 (O_289,N_2980,N_2987);
nor UO_290 (O_290,N_2959,N_2997);
or UO_291 (O_291,N_2966,N_2950);
nor UO_292 (O_292,N_2992,N_2951);
nand UO_293 (O_293,N_2952,N_2982);
and UO_294 (O_294,N_2998,N_2991);
or UO_295 (O_295,N_2967,N_2988);
and UO_296 (O_296,N_2953,N_2969);
or UO_297 (O_297,N_2984,N_2967);
nand UO_298 (O_298,N_2977,N_2976);
nor UO_299 (O_299,N_2988,N_2997);
or UO_300 (O_300,N_2971,N_2968);
nand UO_301 (O_301,N_2971,N_2993);
and UO_302 (O_302,N_2963,N_2952);
or UO_303 (O_303,N_2961,N_2962);
and UO_304 (O_304,N_2971,N_2957);
and UO_305 (O_305,N_2994,N_2976);
and UO_306 (O_306,N_2998,N_2958);
nor UO_307 (O_307,N_2959,N_2983);
nor UO_308 (O_308,N_2971,N_2997);
nor UO_309 (O_309,N_2951,N_2964);
or UO_310 (O_310,N_2983,N_2997);
or UO_311 (O_311,N_2956,N_2966);
nor UO_312 (O_312,N_2962,N_2950);
nand UO_313 (O_313,N_2982,N_2977);
and UO_314 (O_314,N_2969,N_2995);
and UO_315 (O_315,N_2954,N_2958);
and UO_316 (O_316,N_2958,N_2963);
nor UO_317 (O_317,N_2997,N_2957);
or UO_318 (O_318,N_2997,N_2998);
nor UO_319 (O_319,N_2955,N_2987);
nand UO_320 (O_320,N_2961,N_2968);
nor UO_321 (O_321,N_2999,N_2971);
nand UO_322 (O_322,N_2971,N_2959);
or UO_323 (O_323,N_2957,N_2959);
nand UO_324 (O_324,N_2996,N_2967);
and UO_325 (O_325,N_2962,N_2984);
or UO_326 (O_326,N_2989,N_2950);
or UO_327 (O_327,N_2960,N_2998);
nand UO_328 (O_328,N_2982,N_2984);
or UO_329 (O_329,N_2958,N_2964);
and UO_330 (O_330,N_2957,N_2974);
nor UO_331 (O_331,N_2965,N_2954);
and UO_332 (O_332,N_2951,N_2970);
nand UO_333 (O_333,N_2973,N_2971);
or UO_334 (O_334,N_2990,N_2993);
nor UO_335 (O_335,N_2972,N_2959);
nand UO_336 (O_336,N_2967,N_2966);
nor UO_337 (O_337,N_2977,N_2995);
nor UO_338 (O_338,N_2965,N_2971);
nor UO_339 (O_339,N_2970,N_2999);
or UO_340 (O_340,N_2955,N_2975);
nand UO_341 (O_341,N_2975,N_2977);
or UO_342 (O_342,N_2953,N_2954);
or UO_343 (O_343,N_2987,N_2969);
or UO_344 (O_344,N_2955,N_2968);
nand UO_345 (O_345,N_2978,N_2998);
nor UO_346 (O_346,N_2986,N_2959);
nor UO_347 (O_347,N_2993,N_2984);
nand UO_348 (O_348,N_2994,N_2990);
and UO_349 (O_349,N_2987,N_2990);
and UO_350 (O_350,N_2952,N_2957);
nand UO_351 (O_351,N_2982,N_2985);
nor UO_352 (O_352,N_2952,N_2966);
nor UO_353 (O_353,N_2968,N_2965);
nand UO_354 (O_354,N_2952,N_2994);
nand UO_355 (O_355,N_2988,N_2985);
nor UO_356 (O_356,N_2966,N_2958);
or UO_357 (O_357,N_2979,N_2973);
and UO_358 (O_358,N_2984,N_2961);
nor UO_359 (O_359,N_2950,N_2996);
and UO_360 (O_360,N_2952,N_2965);
and UO_361 (O_361,N_2979,N_2954);
and UO_362 (O_362,N_2991,N_2977);
and UO_363 (O_363,N_2999,N_2984);
and UO_364 (O_364,N_2986,N_2989);
nand UO_365 (O_365,N_2954,N_2997);
or UO_366 (O_366,N_2966,N_2994);
and UO_367 (O_367,N_2974,N_2972);
and UO_368 (O_368,N_2954,N_2992);
nand UO_369 (O_369,N_2951,N_2974);
nor UO_370 (O_370,N_2984,N_2996);
and UO_371 (O_371,N_2973,N_2990);
nor UO_372 (O_372,N_2964,N_2998);
or UO_373 (O_373,N_2952,N_2972);
nor UO_374 (O_374,N_2987,N_2997);
or UO_375 (O_375,N_2999,N_2965);
and UO_376 (O_376,N_2963,N_2973);
or UO_377 (O_377,N_2968,N_2985);
nand UO_378 (O_378,N_2972,N_2965);
nor UO_379 (O_379,N_2954,N_2994);
or UO_380 (O_380,N_2978,N_2971);
and UO_381 (O_381,N_2958,N_2951);
nand UO_382 (O_382,N_2964,N_2967);
nand UO_383 (O_383,N_2969,N_2985);
and UO_384 (O_384,N_2979,N_2951);
or UO_385 (O_385,N_2982,N_2989);
and UO_386 (O_386,N_2970,N_2983);
nor UO_387 (O_387,N_2995,N_2957);
and UO_388 (O_388,N_2950,N_2971);
nor UO_389 (O_389,N_2983,N_2971);
and UO_390 (O_390,N_2969,N_2979);
or UO_391 (O_391,N_2976,N_2983);
and UO_392 (O_392,N_2955,N_2976);
or UO_393 (O_393,N_2999,N_2994);
xor UO_394 (O_394,N_2990,N_2984);
and UO_395 (O_395,N_2995,N_2993);
nand UO_396 (O_396,N_2960,N_2994);
or UO_397 (O_397,N_2951,N_2976);
or UO_398 (O_398,N_2984,N_2954);
nor UO_399 (O_399,N_2991,N_2987);
and UO_400 (O_400,N_2981,N_2971);
and UO_401 (O_401,N_2951,N_2962);
or UO_402 (O_402,N_2950,N_2991);
nand UO_403 (O_403,N_2991,N_2983);
nor UO_404 (O_404,N_2974,N_2996);
and UO_405 (O_405,N_2986,N_2969);
or UO_406 (O_406,N_2985,N_2987);
nand UO_407 (O_407,N_2965,N_2956);
nand UO_408 (O_408,N_2979,N_2962);
nor UO_409 (O_409,N_2990,N_2968);
or UO_410 (O_410,N_2956,N_2987);
and UO_411 (O_411,N_2959,N_2955);
nand UO_412 (O_412,N_2957,N_2975);
nand UO_413 (O_413,N_2989,N_2972);
and UO_414 (O_414,N_2989,N_2963);
nand UO_415 (O_415,N_2976,N_2964);
and UO_416 (O_416,N_2973,N_2962);
or UO_417 (O_417,N_2984,N_2992);
and UO_418 (O_418,N_2970,N_2972);
nand UO_419 (O_419,N_2974,N_2967);
nor UO_420 (O_420,N_2984,N_2953);
nand UO_421 (O_421,N_2988,N_2970);
or UO_422 (O_422,N_2989,N_2956);
nor UO_423 (O_423,N_2982,N_2991);
nand UO_424 (O_424,N_2955,N_2963);
xnor UO_425 (O_425,N_2999,N_2961);
or UO_426 (O_426,N_2978,N_2962);
nand UO_427 (O_427,N_2975,N_2989);
and UO_428 (O_428,N_2958,N_2952);
nor UO_429 (O_429,N_2989,N_2951);
nand UO_430 (O_430,N_2961,N_2973);
and UO_431 (O_431,N_2994,N_2961);
or UO_432 (O_432,N_2960,N_2997);
or UO_433 (O_433,N_2982,N_2968);
nor UO_434 (O_434,N_2991,N_2994);
or UO_435 (O_435,N_2950,N_2954);
nand UO_436 (O_436,N_2975,N_2951);
nand UO_437 (O_437,N_2982,N_2967);
or UO_438 (O_438,N_2987,N_2951);
nor UO_439 (O_439,N_2980,N_2993);
nor UO_440 (O_440,N_2964,N_2980);
and UO_441 (O_441,N_2987,N_2981);
xnor UO_442 (O_442,N_2992,N_2963);
nand UO_443 (O_443,N_2956,N_2971);
and UO_444 (O_444,N_2950,N_2987);
and UO_445 (O_445,N_2959,N_2998);
nor UO_446 (O_446,N_2963,N_2998);
or UO_447 (O_447,N_2992,N_2950);
nor UO_448 (O_448,N_2984,N_2964);
or UO_449 (O_449,N_2957,N_2978);
and UO_450 (O_450,N_2975,N_2965);
nor UO_451 (O_451,N_2977,N_2989);
or UO_452 (O_452,N_2965,N_2951);
nand UO_453 (O_453,N_2957,N_2960);
nand UO_454 (O_454,N_2993,N_2974);
nor UO_455 (O_455,N_2986,N_2984);
and UO_456 (O_456,N_2958,N_2953);
nand UO_457 (O_457,N_2959,N_2965);
nor UO_458 (O_458,N_2959,N_2953);
nand UO_459 (O_459,N_2997,N_2979);
nor UO_460 (O_460,N_2970,N_2953);
or UO_461 (O_461,N_2990,N_2992);
nand UO_462 (O_462,N_2967,N_2972);
nand UO_463 (O_463,N_2962,N_2988);
or UO_464 (O_464,N_2974,N_2956);
nand UO_465 (O_465,N_2957,N_2956);
or UO_466 (O_466,N_2965,N_2970);
and UO_467 (O_467,N_2963,N_2995);
nand UO_468 (O_468,N_2974,N_2991);
nand UO_469 (O_469,N_2992,N_2999);
and UO_470 (O_470,N_2998,N_2987);
and UO_471 (O_471,N_2961,N_2986);
nand UO_472 (O_472,N_2998,N_2985);
and UO_473 (O_473,N_2999,N_2980);
nand UO_474 (O_474,N_2974,N_2968);
and UO_475 (O_475,N_2969,N_2956);
or UO_476 (O_476,N_2958,N_2967);
nor UO_477 (O_477,N_2968,N_2986);
nand UO_478 (O_478,N_2981,N_2968);
nor UO_479 (O_479,N_2968,N_2966);
nand UO_480 (O_480,N_2952,N_2959);
nand UO_481 (O_481,N_2965,N_2991);
and UO_482 (O_482,N_2972,N_2997);
nand UO_483 (O_483,N_2984,N_2987);
nor UO_484 (O_484,N_2951,N_2981);
and UO_485 (O_485,N_2962,N_2967);
nand UO_486 (O_486,N_2987,N_2954);
nor UO_487 (O_487,N_2983,N_2972);
nand UO_488 (O_488,N_2977,N_2985);
nand UO_489 (O_489,N_2992,N_2997);
nor UO_490 (O_490,N_2965,N_2985);
nand UO_491 (O_491,N_2952,N_2967);
or UO_492 (O_492,N_2986,N_2981);
or UO_493 (O_493,N_2967,N_2963);
nor UO_494 (O_494,N_2970,N_2996);
and UO_495 (O_495,N_2976,N_2967);
nor UO_496 (O_496,N_2951,N_2999);
nor UO_497 (O_497,N_2959,N_2974);
nor UO_498 (O_498,N_2960,N_2970);
or UO_499 (O_499,N_2954,N_2963);
endmodule