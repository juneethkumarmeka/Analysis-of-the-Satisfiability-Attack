module basic_500_3000_500_30_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_457,In_250);
nor U1 (N_1,In_4,In_401);
nor U2 (N_2,In_385,In_387);
and U3 (N_3,In_481,In_141);
nor U4 (N_4,In_314,In_20);
nand U5 (N_5,In_469,In_99);
or U6 (N_6,In_35,In_287);
and U7 (N_7,In_204,In_208);
nand U8 (N_8,In_53,In_332);
nand U9 (N_9,In_40,In_416);
nor U10 (N_10,In_116,In_483);
nor U11 (N_11,In_26,In_437);
and U12 (N_12,In_167,In_273);
and U13 (N_13,In_338,In_216);
or U14 (N_14,In_475,In_18);
or U15 (N_15,In_374,In_299);
and U16 (N_16,In_149,In_212);
nor U17 (N_17,In_242,In_177);
nand U18 (N_18,In_383,In_45);
and U19 (N_19,In_136,In_472);
and U20 (N_20,In_420,In_106);
nand U21 (N_21,In_340,In_182);
nor U22 (N_22,In_24,In_324);
or U23 (N_23,In_108,In_221);
nor U24 (N_24,In_95,In_310);
and U25 (N_25,In_462,In_169);
nand U26 (N_26,In_209,In_161);
nor U27 (N_27,In_77,In_289);
or U28 (N_28,In_274,In_346);
nand U29 (N_29,In_137,In_361);
or U30 (N_30,In_120,In_369);
or U31 (N_31,In_202,In_386);
and U32 (N_32,In_367,In_156);
nand U33 (N_33,In_68,In_308);
and U34 (N_34,In_105,In_276);
nand U35 (N_35,In_230,In_57);
nor U36 (N_36,In_330,In_260);
nor U37 (N_37,In_78,In_2);
or U38 (N_38,In_298,In_138);
and U39 (N_39,In_27,In_21);
nand U40 (N_40,In_266,In_194);
xor U41 (N_41,In_454,In_112);
and U42 (N_42,In_365,In_316);
and U43 (N_43,In_284,In_244);
nand U44 (N_44,In_335,In_418);
nor U45 (N_45,In_490,In_214);
nand U46 (N_46,In_465,In_431);
or U47 (N_47,In_318,In_479);
nand U48 (N_48,In_3,In_205);
nand U49 (N_49,In_121,In_262);
nand U50 (N_50,In_237,In_271);
nor U51 (N_51,In_428,In_229);
or U52 (N_52,In_81,In_275);
nor U53 (N_53,In_439,In_394);
or U54 (N_54,In_119,In_162);
nand U55 (N_55,In_282,In_80);
nand U56 (N_56,In_384,In_29);
or U57 (N_57,In_251,In_432);
xnor U58 (N_58,In_217,In_132);
and U59 (N_59,In_484,In_16);
and U60 (N_60,In_133,In_43);
nand U61 (N_61,In_72,In_464);
nand U62 (N_62,In_478,In_117);
nor U63 (N_63,In_371,In_56);
nor U64 (N_64,In_159,In_232);
or U65 (N_65,In_312,In_493);
and U66 (N_66,In_203,In_151);
or U67 (N_67,In_55,In_339);
xnor U68 (N_68,In_435,In_259);
nand U69 (N_69,In_429,In_373);
nor U70 (N_70,In_466,In_296);
nand U71 (N_71,In_235,In_102);
nor U72 (N_72,In_172,In_206);
and U73 (N_73,In_424,In_405);
nor U74 (N_74,In_379,In_63);
nor U75 (N_75,In_219,In_305);
nand U76 (N_76,In_460,In_497);
nand U77 (N_77,In_449,In_227);
or U78 (N_78,In_453,In_351);
nand U79 (N_79,In_427,In_239);
and U80 (N_80,In_113,In_9);
nand U81 (N_81,In_269,In_403);
nor U82 (N_82,In_158,In_228);
nor U83 (N_83,In_349,In_360);
nor U84 (N_84,In_461,In_38);
nor U85 (N_85,In_123,In_468);
nand U86 (N_86,In_104,In_255);
nand U87 (N_87,In_50,In_415);
or U88 (N_88,In_155,In_64);
nor U89 (N_89,In_485,In_12);
or U90 (N_90,In_59,In_392);
nand U91 (N_91,In_76,In_328);
or U92 (N_92,In_97,In_128);
and U93 (N_93,In_193,In_356);
nand U94 (N_94,In_425,In_163);
nor U95 (N_95,In_486,In_412);
and U96 (N_96,In_455,In_224);
nor U97 (N_97,In_86,In_71);
nand U98 (N_98,In_279,In_436);
or U99 (N_99,In_225,In_196);
and U100 (N_100,In_309,N_72);
nand U101 (N_101,In_451,In_467);
nand U102 (N_102,In_286,In_301);
nor U103 (N_103,In_293,In_115);
and U104 (N_104,In_498,In_445);
or U105 (N_105,In_359,N_36);
and U106 (N_106,In_201,N_83);
nor U107 (N_107,In_323,In_61);
and U108 (N_108,N_68,N_21);
nand U109 (N_109,N_31,N_1);
or U110 (N_110,N_23,In_122);
and U111 (N_111,In_192,In_341);
and U112 (N_112,In_408,In_218);
nor U113 (N_113,In_452,In_101);
nor U114 (N_114,N_17,N_82);
nor U115 (N_115,In_294,N_46);
or U116 (N_116,In_47,In_67);
nand U117 (N_117,In_433,N_13);
nand U118 (N_118,N_52,In_291);
or U119 (N_119,In_98,N_55);
or U120 (N_120,N_50,In_370);
and U121 (N_121,In_315,In_381);
or U122 (N_122,In_28,In_311);
nand U123 (N_123,N_18,In_5);
or U124 (N_124,N_5,In_37);
nor U125 (N_125,In_107,In_25);
xor U126 (N_126,In_376,In_168);
or U127 (N_127,N_96,N_59);
nor U128 (N_128,In_307,In_258);
nor U129 (N_129,In_165,In_372);
or U130 (N_130,N_90,In_337);
nor U131 (N_131,N_41,N_43);
and U132 (N_132,In_413,N_66);
or U133 (N_133,In_391,In_355);
nand U134 (N_134,In_74,N_48);
or U135 (N_135,N_67,In_253);
and U136 (N_136,In_447,In_263);
nand U137 (N_137,In_135,N_22);
and U138 (N_138,N_65,In_272);
or U139 (N_139,In_426,In_364);
or U140 (N_140,In_252,In_144);
nor U141 (N_141,In_213,In_110);
xnor U142 (N_142,In_147,In_344);
nor U143 (N_143,N_6,N_54);
and U144 (N_144,In_281,N_42);
nand U145 (N_145,In_111,In_243);
or U146 (N_146,In_10,In_322);
or U147 (N_147,In_423,In_83);
nand U148 (N_148,In_6,In_154);
xor U149 (N_149,In_94,N_30);
or U150 (N_150,In_395,In_70);
nand U151 (N_151,In_334,N_84);
or U152 (N_152,N_69,N_85);
nand U153 (N_153,In_199,In_358);
or U154 (N_154,In_362,In_377);
and U155 (N_155,In_267,In_89);
xnor U156 (N_156,In_174,In_444);
xor U157 (N_157,In_180,N_8);
nand U158 (N_158,In_130,In_233);
nand U159 (N_159,In_348,In_103);
and U160 (N_160,In_399,In_304);
nand U161 (N_161,N_12,In_58);
nor U162 (N_162,In_368,In_257);
or U163 (N_163,N_28,In_350);
and U164 (N_164,In_458,In_407);
nor U165 (N_165,N_9,In_480);
or U166 (N_166,N_33,In_438);
nand U167 (N_167,In_23,N_53);
or U168 (N_168,In_441,In_226);
or U169 (N_169,In_131,In_292);
and U170 (N_170,In_280,In_22);
and U171 (N_171,In_69,In_84);
or U172 (N_172,In_354,In_175);
or U173 (N_173,In_187,N_71);
nand U174 (N_174,N_7,N_16);
nand U175 (N_175,N_27,N_78);
or U176 (N_176,In_166,In_66);
nand U177 (N_177,In_397,In_143);
and U178 (N_178,In_114,In_8);
or U179 (N_179,In_118,In_1);
or U180 (N_180,In_248,In_492);
nor U181 (N_181,In_51,In_398);
nor U182 (N_182,In_471,In_146);
nor U183 (N_183,In_278,In_207);
and U184 (N_184,In_406,In_211);
nor U185 (N_185,N_2,In_236);
or U186 (N_186,N_61,In_474);
and U187 (N_187,In_487,In_164);
nand U188 (N_188,In_54,In_173);
and U189 (N_189,In_90,N_29);
and U190 (N_190,N_38,In_210);
and U191 (N_191,In_85,In_306);
nand U192 (N_192,In_380,In_247);
nor U193 (N_193,In_241,In_446);
and U194 (N_194,In_473,In_223);
and U195 (N_195,In_52,In_396);
nor U196 (N_196,N_93,In_421);
nand U197 (N_197,In_181,In_11);
nor U198 (N_198,In_256,In_494);
nor U199 (N_199,In_139,In_347);
nand U200 (N_200,N_39,N_40);
xor U201 (N_201,In_189,In_336);
nand U202 (N_202,In_109,In_96);
nand U203 (N_203,N_103,In_268);
nor U204 (N_204,In_265,N_80);
and U205 (N_205,In_456,N_174);
or U206 (N_206,N_186,N_157);
and U207 (N_207,In_129,N_3);
nand U208 (N_208,In_254,N_62);
nor U209 (N_209,N_192,N_106);
nand U210 (N_210,N_165,N_139);
nand U211 (N_211,In_62,In_495);
nor U212 (N_212,N_98,In_491);
nand U213 (N_213,In_343,In_19);
or U214 (N_214,In_36,N_105);
and U215 (N_215,N_196,N_169);
and U216 (N_216,In_100,N_152);
and U217 (N_217,In_88,N_129);
and U218 (N_218,In_342,In_400);
nor U219 (N_219,In_375,N_185);
and U220 (N_220,In_178,In_352);
nor U221 (N_221,N_10,N_177);
and U222 (N_222,In_450,N_148);
and U223 (N_223,In_41,In_15);
nor U224 (N_224,In_353,In_33);
or U225 (N_225,In_222,In_31);
xnor U226 (N_226,N_173,In_152);
nand U227 (N_227,In_499,N_176);
nor U228 (N_228,N_147,In_277);
or U229 (N_229,N_178,N_191);
or U230 (N_230,N_182,In_249);
nand U231 (N_231,N_141,In_410);
and U232 (N_232,N_108,In_65);
and U233 (N_233,In_185,N_11);
nand U234 (N_234,N_167,In_422);
or U235 (N_235,In_404,In_345);
nand U236 (N_236,N_70,N_164);
or U237 (N_237,In_327,N_32);
nor U238 (N_238,In_127,N_194);
and U239 (N_239,In_325,N_14);
nor U240 (N_240,N_117,In_414);
nor U241 (N_241,N_51,In_179);
and U242 (N_242,In_443,In_34);
nor U243 (N_243,N_101,N_64);
nor U244 (N_244,N_20,In_124);
nand U245 (N_245,In_170,N_89);
or U246 (N_246,N_87,In_44);
or U247 (N_247,In_82,N_114);
nand U248 (N_248,In_197,In_388);
nand U249 (N_249,In_434,In_134);
or U250 (N_250,In_39,N_133);
or U251 (N_251,N_81,In_270);
and U252 (N_252,In_357,In_245);
and U253 (N_253,In_125,In_195);
nand U254 (N_254,N_63,In_378);
and U255 (N_255,N_79,In_482);
nor U256 (N_256,N_94,N_145);
nor U257 (N_257,In_186,In_470);
nand U258 (N_258,In_382,N_144);
or U259 (N_259,N_37,In_419);
nand U260 (N_260,N_123,N_73);
nand U261 (N_261,In_14,In_48);
and U262 (N_262,N_35,N_104);
nand U263 (N_263,In_145,In_215);
nor U264 (N_264,N_153,In_389);
or U265 (N_265,In_288,N_179);
and U266 (N_266,N_162,In_13);
nand U267 (N_267,N_149,In_191);
xnor U268 (N_268,In_417,In_320);
nor U269 (N_269,N_158,N_198);
nor U270 (N_270,In_326,In_300);
nor U271 (N_271,N_112,In_496);
or U272 (N_272,In_440,In_126);
nand U273 (N_273,In_142,In_171);
or U274 (N_274,N_171,N_184);
nand U275 (N_275,N_159,In_393);
nand U276 (N_276,N_34,In_234);
or U277 (N_277,N_160,N_197);
nand U278 (N_278,N_107,In_411);
and U279 (N_279,N_0,N_128);
nor U280 (N_280,N_76,N_120);
or U281 (N_281,In_198,N_15);
or U282 (N_282,N_97,N_140);
or U283 (N_283,N_155,N_125);
or U284 (N_284,N_135,N_131);
xor U285 (N_285,N_166,In_157);
nor U286 (N_286,N_47,N_86);
and U287 (N_287,In_7,In_42);
nor U288 (N_288,N_189,N_170);
and U289 (N_289,In_17,N_60);
nand U290 (N_290,N_199,N_124);
and U291 (N_291,In_476,N_77);
or U292 (N_292,N_154,N_111);
or U293 (N_293,In_333,In_409);
and U294 (N_294,N_91,N_4);
nand U295 (N_295,In_176,N_56);
nand U296 (N_296,In_92,In_32);
and U297 (N_297,N_118,N_109);
nand U298 (N_298,In_488,In_297);
nand U299 (N_299,N_121,N_74);
and U300 (N_300,N_248,N_262);
and U301 (N_301,In_160,In_463);
and U302 (N_302,N_127,N_255);
nand U303 (N_303,N_188,In_390);
nand U304 (N_304,N_88,In_91);
and U305 (N_305,N_272,N_236);
nand U306 (N_306,N_92,N_243);
xnor U307 (N_307,N_226,In_363);
and U308 (N_308,In_331,In_459);
nor U309 (N_309,N_216,N_187);
nand U310 (N_310,N_270,N_209);
nand U311 (N_311,N_99,N_193);
xnor U312 (N_312,N_195,In_0);
nor U313 (N_313,N_282,N_274);
or U314 (N_314,N_238,N_240);
nor U315 (N_315,In_188,N_245);
nand U316 (N_316,N_126,N_279);
xnor U317 (N_317,N_214,N_224);
and U318 (N_318,In_261,N_284);
and U319 (N_319,N_44,N_217);
or U320 (N_320,N_235,N_219);
and U321 (N_321,N_142,N_181);
nand U322 (N_322,N_233,N_222);
or U323 (N_323,N_256,N_100);
nand U324 (N_324,N_110,In_321);
or U325 (N_325,N_116,N_206);
nand U326 (N_326,In_183,N_259);
or U327 (N_327,In_87,In_489);
xnor U328 (N_328,N_253,In_477);
nor U329 (N_329,N_183,In_319);
or U330 (N_330,N_289,N_204);
and U331 (N_331,In_264,N_143);
nor U332 (N_332,In_190,N_113);
or U333 (N_333,In_60,N_286);
or U334 (N_334,In_366,In_402);
nand U335 (N_335,N_138,N_290);
or U336 (N_336,N_49,In_302);
nand U337 (N_337,In_73,N_247);
nor U338 (N_338,N_280,N_251);
or U339 (N_339,In_148,N_26);
nor U340 (N_340,N_298,N_136);
or U341 (N_341,N_297,In_329);
xor U342 (N_342,N_232,N_288);
nor U343 (N_343,In_75,N_151);
and U344 (N_344,N_208,N_258);
or U345 (N_345,N_257,N_132);
or U346 (N_346,N_201,N_246);
and U347 (N_347,In_317,In_200);
or U348 (N_348,N_200,In_140);
nor U349 (N_349,N_265,N_115);
and U350 (N_350,N_250,N_161);
nand U351 (N_351,N_266,N_215);
nand U352 (N_352,N_292,In_93);
nand U353 (N_353,N_213,N_220);
or U354 (N_354,N_244,In_79);
or U355 (N_355,N_218,In_150);
or U356 (N_356,N_25,N_296);
and U357 (N_357,N_202,N_234);
and U358 (N_358,N_277,N_163);
and U359 (N_359,N_271,In_46);
or U360 (N_360,N_227,N_175);
nor U361 (N_361,N_102,In_184);
and U362 (N_362,N_299,N_295);
nand U363 (N_363,N_122,N_229);
and U364 (N_364,N_291,N_249);
nor U365 (N_365,N_261,In_283);
nand U366 (N_366,N_58,N_239);
or U367 (N_367,N_19,N_285);
xnor U368 (N_368,N_168,N_150);
nor U369 (N_369,N_146,N_278);
nand U370 (N_370,N_267,N_281);
nand U371 (N_371,N_269,In_231);
and U372 (N_372,N_260,In_290);
nor U373 (N_373,N_287,N_237);
nand U374 (N_374,In_246,N_276);
nand U375 (N_375,N_180,N_24);
or U376 (N_376,In_30,N_221);
nor U377 (N_377,N_293,N_212);
and U378 (N_378,N_172,N_207);
and U379 (N_379,N_223,N_263);
nand U380 (N_380,N_228,N_119);
nor U381 (N_381,In_238,N_57);
nand U382 (N_382,N_275,N_75);
and U383 (N_383,In_303,N_137);
nor U384 (N_384,N_242,In_295);
or U385 (N_385,N_95,N_273);
nand U386 (N_386,N_254,N_268);
xor U387 (N_387,In_442,N_45);
and U388 (N_388,N_241,N_203);
nor U389 (N_389,In_448,N_211);
nor U390 (N_390,N_190,N_225);
nor U391 (N_391,In_49,N_134);
nor U392 (N_392,N_230,N_210);
or U393 (N_393,In_430,N_252);
or U394 (N_394,In_285,N_294);
or U395 (N_395,N_231,In_313);
and U396 (N_396,N_130,In_153);
or U397 (N_397,N_283,N_156);
nor U398 (N_398,In_240,In_220);
or U399 (N_399,N_264,N_205);
and U400 (N_400,N_319,N_342);
nor U401 (N_401,N_354,N_362);
nand U402 (N_402,N_361,N_339);
and U403 (N_403,N_375,N_376);
nand U404 (N_404,N_306,N_324);
nor U405 (N_405,N_386,N_374);
nand U406 (N_406,N_323,N_377);
nand U407 (N_407,N_357,N_325);
nor U408 (N_408,N_379,N_371);
and U409 (N_409,N_373,N_346);
or U410 (N_410,N_338,N_345);
nor U411 (N_411,N_360,N_300);
nand U412 (N_412,N_314,N_318);
and U413 (N_413,N_378,N_329);
nor U414 (N_414,N_343,N_350);
nor U415 (N_415,N_320,N_368);
and U416 (N_416,N_330,N_392);
or U417 (N_417,N_347,N_312);
and U418 (N_418,N_317,N_395);
or U419 (N_419,N_341,N_332);
nor U420 (N_420,N_321,N_389);
and U421 (N_421,N_393,N_356);
nor U422 (N_422,N_387,N_344);
nor U423 (N_423,N_337,N_305);
or U424 (N_424,N_349,N_367);
and U425 (N_425,N_348,N_327);
or U426 (N_426,N_335,N_366);
nor U427 (N_427,N_380,N_309);
and U428 (N_428,N_394,N_353);
nor U429 (N_429,N_399,N_328);
nand U430 (N_430,N_372,N_397);
nand U431 (N_431,N_369,N_322);
nand U432 (N_432,N_307,N_352);
nand U433 (N_433,N_315,N_385);
nand U434 (N_434,N_396,N_316);
or U435 (N_435,N_303,N_334);
and U436 (N_436,N_311,N_388);
nand U437 (N_437,N_398,N_364);
nor U438 (N_438,N_313,N_336);
or U439 (N_439,N_370,N_326);
nor U440 (N_440,N_340,N_351);
and U441 (N_441,N_358,N_301);
nand U442 (N_442,N_310,N_390);
nand U443 (N_443,N_382,N_381);
or U444 (N_444,N_355,N_365);
nor U445 (N_445,N_383,N_333);
and U446 (N_446,N_384,N_391);
or U447 (N_447,N_359,N_363);
nor U448 (N_448,N_302,N_331);
nor U449 (N_449,N_304,N_308);
and U450 (N_450,N_316,N_350);
nand U451 (N_451,N_302,N_360);
nor U452 (N_452,N_394,N_328);
and U453 (N_453,N_372,N_330);
nor U454 (N_454,N_322,N_325);
nor U455 (N_455,N_372,N_307);
nand U456 (N_456,N_305,N_384);
and U457 (N_457,N_324,N_318);
nor U458 (N_458,N_379,N_311);
nor U459 (N_459,N_393,N_313);
nor U460 (N_460,N_337,N_396);
nor U461 (N_461,N_345,N_396);
nor U462 (N_462,N_331,N_320);
or U463 (N_463,N_382,N_393);
nand U464 (N_464,N_331,N_334);
nand U465 (N_465,N_365,N_397);
or U466 (N_466,N_344,N_388);
and U467 (N_467,N_359,N_342);
or U468 (N_468,N_331,N_373);
nor U469 (N_469,N_312,N_374);
or U470 (N_470,N_317,N_361);
and U471 (N_471,N_371,N_319);
nand U472 (N_472,N_305,N_310);
and U473 (N_473,N_394,N_383);
nand U474 (N_474,N_333,N_348);
or U475 (N_475,N_322,N_387);
nor U476 (N_476,N_364,N_396);
nor U477 (N_477,N_326,N_385);
and U478 (N_478,N_311,N_343);
and U479 (N_479,N_350,N_318);
and U480 (N_480,N_367,N_331);
and U481 (N_481,N_362,N_389);
or U482 (N_482,N_357,N_327);
or U483 (N_483,N_352,N_390);
or U484 (N_484,N_395,N_334);
nand U485 (N_485,N_371,N_338);
or U486 (N_486,N_304,N_347);
or U487 (N_487,N_365,N_316);
or U488 (N_488,N_384,N_320);
or U489 (N_489,N_332,N_395);
or U490 (N_490,N_321,N_304);
nor U491 (N_491,N_311,N_312);
nand U492 (N_492,N_354,N_308);
nand U493 (N_493,N_309,N_306);
and U494 (N_494,N_325,N_398);
and U495 (N_495,N_370,N_377);
or U496 (N_496,N_338,N_321);
or U497 (N_497,N_333,N_306);
or U498 (N_498,N_393,N_383);
and U499 (N_499,N_329,N_399);
or U500 (N_500,N_432,N_489);
nor U501 (N_501,N_412,N_443);
nand U502 (N_502,N_439,N_401);
nor U503 (N_503,N_456,N_454);
nand U504 (N_504,N_474,N_484);
nor U505 (N_505,N_437,N_492);
or U506 (N_506,N_457,N_421);
and U507 (N_507,N_466,N_451);
and U508 (N_508,N_429,N_407);
nand U509 (N_509,N_479,N_460);
nor U510 (N_510,N_470,N_462);
nand U511 (N_511,N_424,N_402);
nand U512 (N_512,N_446,N_405);
or U513 (N_513,N_400,N_410);
and U514 (N_514,N_473,N_440);
xnor U515 (N_515,N_485,N_465);
and U516 (N_516,N_441,N_431);
nand U517 (N_517,N_472,N_430);
nand U518 (N_518,N_420,N_418);
and U519 (N_519,N_415,N_481);
nor U520 (N_520,N_450,N_416);
nand U521 (N_521,N_476,N_453);
and U522 (N_522,N_490,N_464);
and U523 (N_523,N_427,N_477);
or U524 (N_524,N_419,N_434);
nand U525 (N_525,N_455,N_488);
xor U526 (N_526,N_426,N_438);
or U527 (N_527,N_442,N_409);
nor U528 (N_528,N_436,N_480);
nor U529 (N_529,N_447,N_496);
or U530 (N_530,N_404,N_422);
or U531 (N_531,N_411,N_413);
or U532 (N_532,N_475,N_469);
and U533 (N_533,N_487,N_425);
and U534 (N_534,N_483,N_467);
xnor U535 (N_535,N_403,N_445);
nor U536 (N_536,N_461,N_498);
nor U537 (N_537,N_435,N_444);
nand U538 (N_538,N_471,N_417);
nand U539 (N_539,N_493,N_491);
nor U540 (N_540,N_495,N_499);
nor U541 (N_541,N_459,N_463);
xor U542 (N_542,N_458,N_468);
xor U543 (N_543,N_414,N_486);
nand U544 (N_544,N_494,N_428);
and U545 (N_545,N_406,N_452);
nor U546 (N_546,N_433,N_478);
nand U547 (N_547,N_482,N_423);
or U548 (N_548,N_448,N_497);
nand U549 (N_549,N_408,N_449);
and U550 (N_550,N_424,N_403);
and U551 (N_551,N_406,N_478);
and U552 (N_552,N_427,N_469);
and U553 (N_553,N_459,N_441);
nand U554 (N_554,N_432,N_469);
nand U555 (N_555,N_479,N_448);
nor U556 (N_556,N_477,N_443);
or U557 (N_557,N_442,N_413);
or U558 (N_558,N_487,N_485);
or U559 (N_559,N_499,N_428);
or U560 (N_560,N_499,N_429);
xnor U561 (N_561,N_411,N_450);
nand U562 (N_562,N_457,N_403);
nor U563 (N_563,N_422,N_463);
nor U564 (N_564,N_450,N_445);
and U565 (N_565,N_468,N_411);
and U566 (N_566,N_431,N_413);
nand U567 (N_567,N_428,N_423);
and U568 (N_568,N_469,N_416);
nor U569 (N_569,N_457,N_446);
or U570 (N_570,N_470,N_426);
and U571 (N_571,N_425,N_494);
nor U572 (N_572,N_460,N_415);
and U573 (N_573,N_441,N_409);
nand U574 (N_574,N_469,N_411);
nand U575 (N_575,N_431,N_442);
and U576 (N_576,N_466,N_458);
nor U577 (N_577,N_462,N_407);
and U578 (N_578,N_439,N_475);
or U579 (N_579,N_440,N_444);
xnor U580 (N_580,N_403,N_430);
nor U581 (N_581,N_462,N_433);
and U582 (N_582,N_429,N_412);
nand U583 (N_583,N_427,N_464);
or U584 (N_584,N_435,N_491);
or U585 (N_585,N_406,N_403);
and U586 (N_586,N_440,N_451);
nor U587 (N_587,N_400,N_451);
and U588 (N_588,N_454,N_439);
and U589 (N_589,N_416,N_447);
nor U590 (N_590,N_426,N_462);
nand U591 (N_591,N_472,N_476);
xnor U592 (N_592,N_499,N_406);
nand U593 (N_593,N_424,N_468);
or U594 (N_594,N_492,N_458);
nand U595 (N_595,N_449,N_458);
and U596 (N_596,N_452,N_497);
and U597 (N_597,N_471,N_428);
nor U598 (N_598,N_449,N_422);
nor U599 (N_599,N_402,N_443);
and U600 (N_600,N_563,N_508);
or U601 (N_601,N_513,N_558);
and U602 (N_602,N_529,N_518);
or U603 (N_603,N_500,N_554);
and U604 (N_604,N_571,N_507);
nand U605 (N_605,N_584,N_561);
or U606 (N_606,N_533,N_545);
nand U607 (N_607,N_585,N_557);
or U608 (N_608,N_520,N_534);
and U609 (N_609,N_575,N_509);
or U610 (N_610,N_576,N_505);
nand U611 (N_611,N_569,N_565);
or U612 (N_612,N_526,N_547);
and U613 (N_613,N_590,N_555);
nand U614 (N_614,N_551,N_542);
nor U615 (N_615,N_597,N_516);
or U616 (N_616,N_587,N_589);
or U617 (N_617,N_539,N_566);
or U618 (N_618,N_540,N_536);
nand U619 (N_619,N_592,N_532);
nor U620 (N_620,N_574,N_593);
or U621 (N_621,N_579,N_588);
and U622 (N_622,N_530,N_519);
nand U623 (N_623,N_560,N_596);
or U624 (N_624,N_580,N_583);
or U625 (N_625,N_548,N_506);
or U626 (N_626,N_517,N_543);
and U627 (N_627,N_581,N_573);
nor U628 (N_628,N_503,N_594);
nand U629 (N_629,N_568,N_537);
or U630 (N_630,N_553,N_501);
nor U631 (N_631,N_567,N_535);
and U632 (N_632,N_546,N_525);
nand U633 (N_633,N_531,N_595);
or U634 (N_634,N_549,N_515);
or U635 (N_635,N_527,N_552);
nand U636 (N_636,N_559,N_564);
and U637 (N_637,N_521,N_511);
nand U638 (N_638,N_514,N_578);
or U639 (N_639,N_504,N_541);
nor U640 (N_640,N_512,N_544);
and U641 (N_641,N_577,N_582);
nor U642 (N_642,N_570,N_556);
or U643 (N_643,N_538,N_510);
or U644 (N_644,N_524,N_502);
nor U645 (N_645,N_591,N_522);
xnor U646 (N_646,N_550,N_598);
and U647 (N_647,N_572,N_523);
nand U648 (N_648,N_586,N_599);
nor U649 (N_649,N_528,N_562);
or U650 (N_650,N_553,N_528);
or U651 (N_651,N_599,N_551);
nor U652 (N_652,N_597,N_507);
and U653 (N_653,N_501,N_597);
nand U654 (N_654,N_502,N_513);
or U655 (N_655,N_559,N_516);
and U656 (N_656,N_585,N_560);
or U657 (N_657,N_584,N_570);
nor U658 (N_658,N_536,N_599);
nor U659 (N_659,N_538,N_525);
and U660 (N_660,N_577,N_548);
and U661 (N_661,N_544,N_587);
nand U662 (N_662,N_500,N_534);
and U663 (N_663,N_556,N_548);
nand U664 (N_664,N_513,N_560);
or U665 (N_665,N_507,N_599);
and U666 (N_666,N_568,N_599);
and U667 (N_667,N_526,N_513);
or U668 (N_668,N_513,N_564);
or U669 (N_669,N_506,N_507);
and U670 (N_670,N_537,N_579);
xor U671 (N_671,N_532,N_523);
and U672 (N_672,N_566,N_507);
nor U673 (N_673,N_547,N_520);
or U674 (N_674,N_581,N_556);
and U675 (N_675,N_578,N_529);
and U676 (N_676,N_552,N_593);
nor U677 (N_677,N_510,N_596);
xnor U678 (N_678,N_520,N_573);
nand U679 (N_679,N_558,N_530);
and U680 (N_680,N_517,N_550);
and U681 (N_681,N_589,N_571);
nand U682 (N_682,N_508,N_537);
or U683 (N_683,N_523,N_546);
nor U684 (N_684,N_537,N_596);
nor U685 (N_685,N_544,N_535);
or U686 (N_686,N_546,N_544);
nand U687 (N_687,N_599,N_588);
nand U688 (N_688,N_544,N_510);
or U689 (N_689,N_520,N_583);
nor U690 (N_690,N_566,N_555);
nand U691 (N_691,N_588,N_544);
and U692 (N_692,N_589,N_508);
or U693 (N_693,N_572,N_508);
and U694 (N_694,N_544,N_531);
xor U695 (N_695,N_584,N_589);
xnor U696 (N_696,N_597,N_547);
xor U697 (N_697,N_556,N_502);
nor U698 (N_698,N_570,N_536);
nand U699 (N_699,N_524,N_598);
or U700 (N_700,N_611,N_668);
xor U701 (N_701,N_619,N_625);
nand U702 (N_702,N_650,N_648);
and U703 (N_703,N_620,N_640);
nand U704 (N_704,N_633,N_628);
or U705 (N_705,N_695,N_641);
and U706 (N_706,N_688,N_663);
nor U707 (N_707,N_653,N_605);
and U708 (N_708,N_639,N_659);
nand U709 (N_709,N_666,N_634);
and U710 (N_710,N_655,N_687);
nor U711 (N_711,N_657,N_638);
nor U712 (N_712,N_652,N_609);
and U713 (N_713,N_603,N_630);
nand U714 (N_714,N_616,N_643);
nand U715 (N_715,N_631,N_601);
and U716 (N_716,N_636,N_674);
nand U717 (N_717,N_645,N_617);
or U718 (N_718,N_654,N_686);
or U719 (N_719,N_661,N_690);
nand U720 (N_720,N_684,N_632);
nand U721 (N_721,N_673,N_626);
nand U722 (N_722,N_649,N_615);
nand U723 (N_723,N_642,N_691);
and U724 (N_724,N_656,N_651);
or U725 (N_725,N_685,N_627);
nand U726 (N_726,N_694,N_681);
nand U727 (N_727,N_680,N_665);
or U728 (N_728,N_604,N_699);
and U729 (N_729,N_679,N_698);
xor U730 (N_730,N_672,N_677);
nor U731 (N_731,N_664,N_622);
and U732 (N_732,N_692,N_635);
and U733 (N_733,N_671,N_678);
and U734 (N_734,N_610,N_662);
nand U735 (N_735,N_614,N_667);
nor U736 (N_736,N_621,N_669);
nor U737 (N_737,N_623,N_696);
nor U738 (N_738,N_644,N_608);
or U739 (N_739,N_600,N_602);
and U740 (N_740,N_682,N_693);
or U741 (N_741,N_647,N_683);
nor U742 (N_742,N_660,N_676);
nand U743 (N_743,N_629,N_675);
nor U744 (N_744,N_624,N_670);
and U745 (N_745,N_658,N_613);
and U746 (N_746,N_612,N_607);
or U747 (N_747,N_689,N_606);
xnor U748 (N_748,N_618,N_697);
nor U749 (N_749,N_646,N_637);
nand U750 (N_750,N_636,N_609);
and U751 (N_751,N_606,N_635);
or U752 (N_752,N_685,N_620);
nand U753 (N_753,N_608,N_678);
nand U754 (N_754,N_670,N_671);
nor U755 (N_755,N_660,N_648);
or U756 (N_756,N_682,N_660);
nand U757 (N_757,N_677,N_660);
nor U758 (N_758,N_601,N_617);
nor U759 (N_759,N_691,N_669);
nand U760 (N_760,N_680,N_626);
and U761 (N_761,N_603,N_659);
xnor U762 (N_762,N_672,N_696);
nand U763 (N_763,N_688,N_631);
and U764 (N_764,N_658,N_647);
or U765 (N_765,N_680,N_611);
and U766 (N_766,N_672,N_661);
nor U767 (N_767,N_642,N_630);
nor U768 (N_768,N_601,N_665);
nand U769 (N_769,N_669,N_687);
and U770 (N_770,N_610,N_630);
nor U771 (N_771,N_627,N_661);
nand U772 (N_772,N_673,N_674);
and U773 (N_773,N_622,N_602);
nand U774 (N_774,N_695,N_623);
nand U775 (N_775,N_627,N_615);
or U776 (N_776,N_602,N_618);
nor U777 (N_777,N_628,N_625);
nand U778 (N_778,N_658,N_665);
or U779 (N_779,N_620,N_663);
nand U780 (N_780,N_628,N_662);
nor U781 (N_781,N_605,N_613);
nor U782 (N_782,N_612,N_613);
xnor U783 (N_783,N_695,N_692);
or U784 (N_784,N_668,N_674);
and U785 (N_785,N_693,N_673);
and U786 (N_786,N_666,N_677);
xor U787 (N_787,N_605,N_620);
nand U788 (N_788,N_696,N_663);
nor U789 (N_789,N_614,N_653);
nand U790 (N_790,N_654,N_639);
nor U791 (N_791,N_688,N_637);
and U792 (N_792,N_678,N_641);
or U793 (N_793,N_649,N_663);
nor U794 (N_794,N_660,N_674);
xor U795 (N_795,N_601,N_637);
and U796 (N_796,N_619,N_600);
and U797 (N_797,N_638,N_639);
and U798 (N_798,N_642,N_613);
or U799 (N_799,N_601,N_630);
xor U800 (N_800,N_736,N_756);
or U801 (N_801,N_728,N_780);
or U802 (N_802,N_701,N_738);
nor U803 (N_803,N_730,N_710);
nor U804 (N_804,N_748,N_735);
nand U805 (N_805,N_755,N_713);
nand U806 (N_806,N_744,N_762);
nor U807 (N_807,N_766,N_742);
nand U808 (N_808,N_774,N_767);
or U809 (N_809,N_714,N_798);
and U810 (N_810,N_783,N_729);
nor U811 (N_811,N_794,N_703);
or U812 (N_812,N_758,N_771);
nand U813 (N_813,N_705,N_718);
or U814 (N_814,N_721,N_706);
nor U815 (N_815,N_787,N_784);
nand U816 (N_816,N_700,N_708);
or U817 (N_817,N_733,N_772);
and U818 (N_818,N_792,N_759);
or U819 (N_819,N_760,N_727);
nand U820 (N_820,N_717,N_796);
and U821 (N_821,N_732,N_750);
or U822 (N_822,N_731,N_765);
and U823 (N_823,N_797,N_770);
nor U824 (N_824,N_795,N_719);
nand U825 (N_825,N_761,N_775);
nor U826 (N_826,N_715,N_752);
nand U827 (N_827,N_769,N_793);
and U828 (N_828,N_712,N_768);
and U829 (N_829,N_785,N_782);
nand U830 (N_830,N_707,N_757);
nor U831 (N_831,N_723,N_786);
nand U832 (N_832,N_763,N_726);
and U833 (N_833,N_753,N_734);
nor U834 (N_834,N_711,N_789);
nand U835 (N_835,N_743,N_745);
nand U836 (N_836,N_749,N_754);
nand U837 (N_837,N_790,N_781);
nor U838 (N_838,N_747,N_764);
nor U839 (N_839,N_778,N_741);
or U840 (N_840,N_702,N_746);
or U841 (N_841,N_720,N_722);
or U842 (N_842,N_709,N_751);
and U843 (N_843,N_776,N_724);
nand U844 (N_844,N_704,N_739);
and U845 (N_845,N_791,N_725);
or U846 (N_846,N_773,N_737);
nand U847 (N_847,N_777,N_740);
or U848 (N_848,N_788,N_799);
and U849 (N_849,N_716,N_779);
nand U850 (N_850,N_795,N_742);
and U851 (N_851,N_716,N_708);
and U852 (N_852,N_785,N_741);
or U853 (N_853,N_751,N_736);
or U854 (N_854,N_790,N_774);
and U855 (N_855,N_794,N_714);
or U856 (N_856,N_736,N_793);
nand U857 (N_857,N_714,N_750);
or U858 (N_858,N_786,N_733);
and U859 (N_859,N_792,N_746);
or U860 (N_860,N_772,N_703);
nand U861 (N_861,N_760,N_743);
and U862 (N_862,N_784,N_762);
nor U863 (N_863,N_763,N_732);
nor U864 (N_864,N_749,N_775);
nor U865 (N_865,N_739,N_740);
or U866 (N_866,N_732,N_797);
and U867 (N_867,N_705,N_775);
and U868 (N_868,N_751,N_784);
xnor U869 (N_869,N_796,N_767);
nand U870 (N_870,N_760,N_710);
nor U871 (N_871,N_707,N_721);
or U872 (N_872,N_754,N_769);
or U873 (N_873,N_726,N_703);
and U874 (N_874,N_730,N_789);
nand U875 (N_875,N_755,N_783);
nand U876 (N_876,N_707,N_728);
nor U877 (N_877,N_742,N_704);
and U878 (N_878,N_722,N_709);
xnor U879 (N_879,N_761,N_740);
and U880 (N_880,N_707,N_743);
nor U881 (N_881,N_723,N_791);
nand U882 (N_882,N_732,N_758);
or U883 (N_883,N_729,N_798);
xnor U884 (N_884,N_757,N_716);
or U885 (N_885,N_742,N_782);
nor U886 (N_886,N_786,N_743);
nand U887 (N_887,N_784,N_705);
or U888 (N_888,N_794,N_709);
and U889 (N_889,N_741,N_797);
nand U890 (N_890,N_726,N_782);
nor U891 (N_891,N_790,N_750);
or U892 (N_892,N_794,N_761);
nor U893 (N_893,N_768,N_715);
and U894 (N_894,N_777,N_714);
and U895 (N_895,N_763,N_755);
nor U896 (N_896,N_791,N_784);
nand U897 (N_897,N_746,N_730);
nor U898 (N_898,N_730,N_782);
nor U899 (N_899,N_753,N_728);
or U900 (N_900,N_873,N_838);
nor U901 (N_901,N_870,N_897);
nor U902 (N_902,N_805,N_820);
xor U903 (N_903,N_858,N_842);
nand U904 (N_904,N_867,N_894);
or U905 (N_905,N_872,N_816);
nor U906 (N_906,N_891,N_861);
nand U907 (N_907,N_813,N_839);
nand U908 (N_908,N_850,N_815);
and U909 (N_909,N_836,N_834);
and U910 (N_910,N_878,N_804);
or U911 (N_911,N_890,N_810);
xor U912 (N_912,N_857,N_893);
xor U913 (N_913,N_831,N_879);
nor U914 (N_914,N_864,N_846);
nand U915 (N_915,N_844,N_882);
nor U916 (N_916,N_868,N_840);
and U917 (N_917,N_887,N_830);
xor U918 (N_918,N_871,N_847);
nor U919 (N_919,N_832,N_852);
xnor U920 (N_920,N_884,N_802);
nand U921 (N_921,N_851,N_881);
or U922 (N_922,N_886,N_862);
nand U923 (N_923,N_877,N_829);
nor U924 (N_924,N_880,N_837);
nor U925 (N_925,N_821,N_827);
or U926 (N_926,N_825,N_841);
or U927 (N_927,N_889,N_803);
or U928 (N_928,N_814,N_845);
and U929 (N_929,N_898,N_859);
nand U930 (N_930,N_865,N_869);
nor U931 (N_931,N_824,N_819);
nor U932 (N_932,N_848,N_811);
and U933 (N_933,N_826,N_888);
nor U934 (N_934,N_895,N_822);
nand U935 (N_935,N_800,N_855);
or U936 (N_936,N_833,N_849);
xor U937 (N_937,N_835,N_863);
or U938 (N_938,N_808,N_809);
or U939 (N_939,N_876,N_818);
nor U940 (N_940,N_892,N_896);
and U941 (N_941,N_853,N_875);
or U942 (N_942,N_812,N_801);
nand U943 (N_943,N_817,N_807);
and U944 (N_944,N_823,N_843);
and U945 (N_945,N_854,N_885);
and U946 (N_946,N_856,N_874);
nor U947 (N_947,N_806,N_899);
nand U948 (N_948,N_866,N_828);
or U949 (N_949,N_860,N_883);
nor U950 (N_950,N_813,N_847);
and U951 (N_951,N_804,N_866);
and U952 (N_952,N_833,N_850);
and U953 (N_953,N_840,N_819);
and U954 (N_954,N_852,N_807);
or U955 (N_955,N_823,N_838);
nand U956 (N_956,N_891,N_810);
nand U957 (N_957,N_813,N_841);
nor U958 (N_958,N_831,N_895);
or U959 (N_959,N_851,N_891);
and U960 (N_960,N_865,N_844);
xor U961 (N_961,N_883,N_851);
nor U962 (N_962,N_822,N_896);
nand U963 (N_963,N_823,N_872);
nand U964 (N_964,N_881,N_866);
or U965 (N_965,N_868,N_841);
or U966 (N_966,N_808,N_854);
and U967 (N_967,N_886,N_819);
or U968 (N_968,N_850,N_816);
or U969 (N_969,N_818,N_835);
nor U970 (N_970,N_879,N_863);
nand U971 (N_971,N_882,N_814);
or U972 (N_972,N_831,N_843);
nand U973 (N_973,N_819,N_830);
nand U974 (N_974,N_859,N_814);
and U975 (N_975,N_866,N_893);
nand U976 (N_976,N_879,N_822);
nor U977 (N_977,N_803,N_811);
or U978 (N_978,N_885,N_818);
nand U979 (N_979,N_843,N_838);
nor U980 (N_980,N_897,N_814);
nand U981 (N_981,N_888,N_817);
or U982 (N_982,N_881,N_884);
or U983 (N_983,N_888,N_849);
nor U984 (N_984,N_880,N_813);
and U985 (N_985,N_855,N_814);
or U986 (N_986,N_836,N_863);
or U987 (N_987,N_800,N_865);
nand U988 (N_988,N_820,N_897);
and U989 (N_989,N_876,N_884);
and U990 (N_990,N_892,N_893);
nor U991 (N_991,N_836,N_895);
or U992 (N_992,N_829,N_854);
nor U993 (N_993,N_881,N_812);
nand U994 (N_994,N_868,N_801);
nand U995 (N_995,N_859,N_829);
or U996 (N_996,N_809,N_835);
and U997 (N_997,N_824,N_839);
or U998 (N_998,N_871,N_891);
nor U999 (N_999,N_850,N_863);
or U1000 (N_1000,N_917,N_933);
nand U1001 (N_1001,N_976,N_923);
or U1002 (N_1002,N_962,N_994);
nor U1003 (N_1003,N_944,N_947);
or U1004 (N_1004,N_912,N_902);
nor U1005 (N_1005,N_995,N_999);
nand U1006 (N_1006,N_935,N_928);
nand U1007 (N_1007,N_953,N_951);
or U1008 (N_1008,N_971,N_901);
or U1009 (N_1009,N_949,N_914);
nor U1010 (N_1010,N_991,N_909);
and U1011 (N_1011,N_964,N_987);
nor U1012 (N_1012,N_956,N_907);
nand U1013 (N_1013,N_913,N_969);
nor U1014 (N_1014,N_970,N_922);
nor U1015 (N_1015,N_989,N_945);
nor U1016 (N_1016,N_983,N_943);
nor U1017 (N_1017,N_990,N_986);
or U1018 (N_1018,N_959,N_980);
nand U1019 (N_1019,N_937,N_984);
or U1020 (N_1020,N_934,N_963);
nand U1021 (N_1021,N_939,N_921);
and U1022 (N_1022,N_993,N_911);
and U1023 (N_1023,N_960,N_985);
or U1024 (N_1024,N_903,N_906);
and U1025 (N_1025,N_916,N_942);
nand U1026 (N_1026,N_941,N_932);
nor U1027 (N_1027,N_948,N_920);
xnor U1028 (N_1028,N_938,N_904);
nand U1029 (N_1029,N_982,N_961);
and U1030 (N_1030,N_954,N_968);
and U1031 (N_1031,N_955,N_946);
or U1032 (N_1032,N_998,N_978);
nor U1033 (N_1033,N_926,N_924);
nand U1034 (N_1034,N_967,N_936);
and U1035 (N_1035,N_972,N_992);
and U1036 (N_1036,N_950,N_988);
nand U1037 (N_1037,N_966,N_918);
and U1038 (N_1038,N_981,N_908);
and U1039 (N_1039,N_905,N_973);
nand U1040 (N_1040,N_952,N_965);
and U1041 (N_1041,N_996,N_900);
and U1042 (N_1042,N_931,N_974);
or U1043 (N_1043,N_940,N_930);
nor U1044 (N_1044,N_958,N_929);
or U1045 (N_1045,N_925,N_919);
nand U1046 (N_1046,N_979,N_975);
nand U1047 (N_1047,N_977,N_927);
and U1048 (N_1048,N_910,N_957);
or U1049 (N_1049,N_915,N_997);
nand U1050 (N_1050,N_974,N_960);
nor U1051 (N_1051,N_997,N_967);
nand U1052 (N_1052,N_969,N_976);
nor U1053 (N_1053,N_980,N_904);
or U1054 (N_1054,N_961,N_907);
and U1055 (N_1055,N_920,N_980);
and U1056 (N_1056,N_906,N_960);
nor U1057 (N_1057,N_948,N_931);
or U1058 (N_1058,N_904,N_984);
xnor U1059 (N_1059,N_989,N_928);
and U1060 (N_1060,N_977,N_961);
or U1061 (N_1061,N_902,N_970);
or U1062 (N_1062,N_950,N_975);
and U1063 (N_1063,N_933,N_990);
nor U1064 (N_1064,N_962,N_967);
or U1065 (N_1065,N_948,N_990);
or U1066 (N_1066,N_924,N_984);
or U1067 (N_1067,N_949,N_991);
nor U1068 (N_1068,N_969,N_975);
and U1069 (N_1069,N_955,N_993);
and U1070 (N_1070,N_990,N_998);
and U1071 (N_1071,N_900,N_939);
nor U1072 (N_1072,N_973,N_992);
nand U1073 (N_1073,N_962,N_947);
nor U1074 (N_1074,N_903,N_986);
and U1075 (N_1075,N_921,N_932);
nand U1076 (N_1076,N_908,N_989);
xnor U1077 (N_1077,N_977,N_906);
and U1078 (N_1078,N_993,N_994);
and U1079 (N_1079,N_998,N_948);
or U1080 (N_1080,N_911,N_982);
or U1081 (N_1081,N_982,N_937);
and U1082 (N_1082,N_978,N_920);
or U1083 (N_1083,N_901,N_992);
nor U1084 (N_1084,N_990,N_929);
and U1085 (N_1085,N_957,N_945);
xnor U1086 (N_1086,N_980,N_950);
or U1087 (N_1087,N_922,N_978);
nand U1088 (N_1088,N_935,N_953);
and U1089 (N_1089,N_978,N_954);
nor U1090 (N_1090,N_920,N_990);
nand U1091 (N_1091,N_949,N_913);
xnor U1092 (N_1092,N_921,N_963);
xor U1093 (N_1093,N_943,N_936);
nor U1094 (N_1094,N_902,N_936);
nand U1095 (N_1095,N_902,N_974);
and U1096 (N_1096,N_995,N_940);
nor U1097 (N_1097,N_992,N_988);
and U1098 (N_1098,N_921,N_954);
or U1099 (N_1099,N_965,N_935);
nand U1100 (N_1100,N_1029,N_1007);
nor U1101 (N_1101,N_1002,N_1056);
or U1102 (N_1102,N_1073,N_1042);
nand U1103 (N_1103,N_1025,N_1031);
nand U1104 (N_1104,N_1013,N_1065);
and U1105 (N_1105,N_1053,N_1015);
and U1106 (N_1106,N_1021,N_1038);
nor U1107 (N_1107,N_1003,N_1083);
and U1108 (N_1108,N_1058,N_1068);
and U1109 (N_1109,N_1076,N_1044);
or U1110 (N_1110,N_1072,N_1075);
and U1111 (N_1111,N_1085,N_1095);
or U1112 (N_1112,N_1091,N_1097);
nand U1113 (N_1113,N_1064,N_1099);
or U1114 (N_1114,N_1066,N_1006);
nor U1115 (N_1115,N_1014,N_1035);
nor U1116 (N_1116,N_1078,N_1090);
nand U1117 (N_1117,N_1026,N_1087);
nand U1118 (N_1118,N_1040,N_1018);
nor U1119 (N_1119,N_1098,N_1061);
and U1120 (N_1120,N_1093,N_1052);
nor U1121 (N_1121,N_1051,N_1039);
and U1122 (N_1122,N_1001,N_1037);
or U1123 (N_1123,N_1027,N_1055);
nand U1124 (N_1124,N_1096,N_1009);
xor U1125 (N_1125,N_1077,N_1071);
nor U1126 (N_1126,N_1016,N_1000);
and U1127 (N_1127,N_1019,N_1063);
nand U1128 (N_1128,N_1084,N_1074);
xnor U1129 (N_1129,N_1022,N_1094);
and U1130 (N_1130,N_1036,N_1059);
nor U1131 (N_1131,N_1079,N_1048);
or U1132 (N_1132,N_1080,N_1062);
or U1133 (N_1133,N_1082,N_1017);
and U1134 (N_1134,N_1023,N_1046);
nor U1135 (N_1135,N_1049,N_1088);
nor U1136 (N_1136,N_1057,N_1089);
nor U1137 (N_1137,N_1005,N_1070);
nand U1138 (N_1138,N_1028,N_1092);
or U1139 (N_1139,N_1060,N_1069);
nand U1140 (N_1140,N_1020,N_1032);
and U1141 (N_1141,N_1012,N_1030);
nand U1142 (N_1142,N_1008,N_1086);
xnor U1143 (N_1143,N_1045,N_1047);
nor U1144 (N_1144,N_1004,N_1010);
or U1145 (N_1145,N_1041,N_1024);
or U1146 (N_1146,N_1081,N_1043);
nand U1147 (N_1147,N_1050,N_1033);
or U1148 (N_1148,N_1011,N_1034);
xnor U1149 (N_1149,N_1054,N_1067);
nor U1150 (N_1150,N_1002,N_1029);
nand U1151 (N_1151,N_1067,N_1056);
and U1152 (N_1152,N_1070,N_1055);
nand U1153 (N_1153,N_1039,N_1088);
nor U1154 (N_1154,N_1072,N_1045);
or U1155 (N_1155,N_1095,N_1039);
nor U1156 (N_1156,N_1028,N_1026);
nand U1157 (N_1157,N_1070,N_1052);
nor U1158 (N_1158,N_1096,N_1006);
nor U1159 (N_1159,N_1076,N_1064);
or U1160 (N_1160,N_1013,N_1075);
or U1161 (N_1161,N_1037,N_1029);
nor U1162 (N_1162,N_1026,N_1068);
and U1163 (N_1163,N_1038,N_1088);
or U1164 (N_1164,N_1013,N_1054);
or U1165 (N_1165,N_1079,N_1066);
nand U1166 (N_1166,N_1035,N_1020);
and U1167 (N_1167,N_1018,N_1094);
nand U1168 (N_1168,N_1049,N_1087);
nand U1169 (N_1169,N_1075,N_1092);
and U1170 (N_1170,N_1051,N_1048);
nand U1171 (N_1171,N_1023,N_1075);
and U1172 (N_1172,N_1087,N_1058);
and U1173 (N_1173,N_1010,N_1073);
and U1174 (N_1174,N_1012,N_1013);
nand U1175 (N_1175,N_1075,N_1063);
or U1176 (N_1176,N_1004,N_1036);
nor U1177 (N_1177,N_1056,N_1024);
and U1178 (N_1178,N_1047,N_1096);
nor U1179 (N_1179,N_1090,N_1061);
nand U1180 (N_1180,N_1011,N_1024);
nand U1181 (N_1181,N_1019,N_1011);
or U1182 (N_1182,N_1093,N_1001);
xnor U1183 (N_1183,N_1009,N_1078);
or U1184 (N_1184,N_1034,N_1073);
or U1185 (N_1185,N_1047,N_1039);
or U1186 (N_1186,N_1043,N_1065);
or U1187 (N_1187,N_1038,N_1050);
or U1188 (N_1188,N_1077,N_1062);
nor U1189 (N_1189,N_1089,N_1015);
nor U1190 (N_1190,N_1065,N_1050);
and U1191 (N_1191,N_1047,N_1053);
xnor U1192 (N_1192,N_1001,N_1081);
nor U1193 (N_1193,N_1097,N_1051);
and U1194 (N_1194,N_1010,N_1091);
and U1195 (N_1195,N_1092,N_1058);
or U1196 (N_1196,N_1077,N_1059);
nor U1197 (N_1197,N_1097,N_1077);
nand U1198 (N_1198,N_1091,N_1030);
nand U1199 (N_1199,N_1031,N_1052);
and U1200 (N_1200,N_1149,N_1154);
and U1201 (N_1201,N_1138,N_1120);
nor U1202 (N_1202,N_1186,N_1191);
nand U1203 (N_1203,N_1122,N_1105);
or U1204 (N_1204,N_1141,N_1173);
nor U1205 (N_1205,N_1123,N_1106);
nor U1206 (N_1206,N_1167,N_1142);
or U1207 (N_1207,N_1174,N_1112);
or U1208 (N_1208,N_1199,N_1189);
nand U1209 (N_1209,N_1179,N_1139);
or U1210 (N_1210,N_1166,N_1172);
nand U1211 (N_1211,N_1116,N_1165);
or U1212 (N_1212,N_1168,N_1137);
and U1213 (N_1213,N_1150,N_1163);
or U1214 (N_1214,N_1152,N_1100);
nand U1215 (N_1215,N_1155,N_1117);
nor U1216 (N_1216,N_1115,N_1182);
nand U1217 (N_1217,N_1134,N_1118);
nor U1218 (N_1218,N_1187,N_1158);
nor U1219 (N_1219,N_1140,N_1136);
and U1220 (N_1220,N_1146,N_1177);
nor U1221 (N_1221,N_1102,N_1121);
nor U1222 (N_1222,N_1160,N_1130);
nor U1223 (N_1223,N_1127,N_1159);
and U1224 (N_1224,N_1156,N_1192);
nor U1225 (N_1225,N_1135,N_1176);
nor U1226 (N_1226,N_1148,N_1157);
and U1227 (N_1227,N_1132,N_1195);
or U1228 (N_1228,N_1162,N_1144);
nor U1229 (N_1229,N_1180,N_1126);
nand U1230 (N_1230,N_1193,N_1190);
nor U1231 (N_1231,N_1145,N_1196);
or U1232 (N_1232,N_1198,N_1151);
and U1233 (N_1233,N_1169,N_1110);
nand U1234 (N_1234,N_1197,N_1128);
nand U1235 (N_1235,N_1171,N_1111);
nor U1236 (N_1236,N_1101,N_1107);
or U1237 (N_1237,N_1125,N_1161);
or U1238 (N_1238,N_1119,N_1185);
nand U1239 (N_1239,N_1131,N_1175);
or U1240 (N_1240,N_1194,N_1170);
and U1241 (N_1241,N_1153,N_1143);
xor U1242 (N_1242,N_1133,N_1113);
or U1243 (N_1243,N_1164,N_1181);
and U1244 (N_1244,N_1108,N_1178);
or U1245 (N_1245,N_1188,N_1124);
or U1246 (N_1246,N_1147,N_1103);
nor U1247 (N_1247,N_1114,N_1104);
or U1248 (N_1248,N_1183,N_1184);
xor U1249 (N_1249,N_1129,N_1109);
and U1250 (N_1250,N_1180,N_1162);
nor U1251 (N_1251,N_1180,N_1151);
and U1252 (N_1252,N_1142,N_1161);
nand U1253 (N_1253,N_1111,N_1184);
nor U1254 (N_1254,N_1188,N_1138);
nor U1255 (N_1255,N_1189,N_1107);
and U1256 (N_1256,N_1126,N_1191);
nor U1257 (N_1257,N_1184,N_1146);
nor U1258 (N_1258,N_1192,N_1162);
and U1259 (N_1259,N_1173,N_1175);
nand U1260 (N_1260,N_1174,N_1109);
nor U1261 (N_1261,N_1196,N_1151);
nor U1262 (N_1262,N_1193,N_1102);
and U1263 (N_1263,N_1171,N_1170);
and U1264 (N_1264,N_1113,N_1190);
nor U1265 (N_1265,N_1172,N_1145);
nor U1266 (N_1266,N_1146,N_1182);
and U1267 (N_1267,N_1189,N_1191);
and U1268 (N_1268,N_1110,N_1155);
and U1269 (N_1269,N_1182,N_1189);
nand U1270 (N_1270,N_1165,N_1144);
nand U1271 (N_1271,N_1177,N_1153);
nand U1272 (N_1272,N_1157,N_1198);
nor U1273 (N_1273,N_1131,N_1114);
and U1274 (N_1274,N_1103,N_1143);
nor U1275 (N_1275,N_1163,N_1170);
and U1276 (N_1276,N_1121,N_1111);
nand U1277 (N_1277,N_1168,N_1140);
or U1278 (N_1278,N_1165,N_1122);
nor U1279 (N_1279,N_1159,N_1114);
nand U1280 (N_1280,N_1130,N_1131);
or U1281 (N_1281,N_1196,N_1112);
and U1282 (N_1282,N_1153,N_1129);
or U1283 (N_1283,N_1123,N_1154);
xor U1284 (N_1284,N_1158,N_1175);
or U1285 (N_1285,N_1185,N_1128);
and U1286 (N_1286,N_1162,N_1185);
nor U1287 (N_1287,N_1147,N_1116);
or U1288 (N_1288,N_1109,N_1112);
or U1289 (N_1289,N_1119,N_1188);
nor U1290 (N_1290,N_1156,N_1154);
nand U1291 (N_1291,N_1106,N_1127);
and U1292 (N_1292,N_1106,N_1102);
and U1293 (N_1293,N_1164,N_1121);
or U1294 (N_1294,N_1111,N_1135);
nor U1295 (N_1295,N_1126,N_1171);
or U1296 (N_1296,N_1127,N_1183);
nand U1297 (N_1297,N_1174,N_1113);
or U1298 (N_1298,N_1154,N_1157);
nor U1299 (N_1299,N_1158,N_1150);
nor U1300 (N_1300,N_1202,N_1269);
nand U1301 (N_1301,N_1288,N_1255);
or U1302 (N_1302,N_1275,N_1280);
nor U1303 (N_1303,N_1289,N_1257);
and U1304 (N_1304,N_1256,N_1272);
and U1305 (N_1305,N_1214,N_1243);
and U1306 (N_1306,N_1200,N_1279);
nand U1307 (N_1307,N_1205,N_1238);
nand U1308 (N_1308,N_1298,N_1281);
nand U1309 (N_1309,N_1283,N_1218);
nor U1310 (N_1310,N_1262,N_1246);
and U1311 (N_1311,N_1203,N_1290);
nor U1312 (N_1312,N_1227,N_1210);
xnor U1313 (N_1313,N_1237,N_1296);
nand U1314 (N_1314,N_1273,N_1252);
or U1315 (N_1315,N_1247,N_1219);
and U1316 (N_1316,N_1221,N_1277);
or U1317 (N_1317,N_1217,N_1201);
nand U1318 (N_1318,N_1224,N_1245);
or U1319 (N_1319,N_1282,N_1204);
nand U1320 (N_1320,N_1241,N_1228);
and U1321 (N_1321,N_1251,N_1250);
nand U1322 (N_1322,N_1260,N_1258);
and U1323 (N_1323,N_1222,N_1230);
nor U1324 (N_1324,N_1270,N_1236);
nor U1325 (N_1325,N_1265,N_1263);
nand U1326 (N_1326,N_1215,N_1261);
or U1327 (N_1327,N_1278,N_1248);
nor U1328 (N_1328,N_1293,N_1212);
nor U1329 (N_1329,N_1268,N_1274);
nor U1330 (N_1330,N_1207,N_1233);
nand U1331 (N_1331,N_1229,N_1271);
nand U1332 (N_1332,N_1276,N_1235);
nand U1333 (N_1333,N_1284,N_1211);
or U1334 (N_1334,N_1287,N_1286);
or U1335 (N_1335,N_1232,N_1242);
and U1336 (N_1336,N_1267,N_1208);
xor U1337 (N_1337,N_1254,N_1206);
and U1338 (N_1338,N_1294,N_1299);
or U1339 (N_1339,N_1249,N_1297);
and U1340 (N_1340,N_1239,N_1209);
and U1341 (N_1341,N_1216,N_1231);
nor U1342 (N_1342,N_1295,N_1220);
or U1343 (N_1343,N_1285,N_1253);
and U1344 (N_1344,N_1266,N_1240);
and U1345 (N_1345,N_1291,N_1292);
and U1346 (N_1346,N_1244,N_1226);
and U1347 (N_1347,N_1264,N_1213);
nand U1348 (N_1348,N_1234,N_1225);
and U1349 (N_1349,N_1223,N_1259);
nor U1350 (N_1350,N_1298,N_1227);
or U1351 (N_1351,N_1252,N_1202);
nor U1352 (N_1352,N_1284,N_1209);
nand U1353 (N_1353,N_1280,N_1288);
and U1354 (N_1354,N_1268,N_1285);
nor U1355 (N_1355,N_1211,N_1298);
or U1356 (N_1356,N_1283,N_1224);
nor U1357 (N_1357,N_1299,N_1290);
nor U1358 (N_1358,N_1213,N_1293);
nor U1359 (N_1359,N_1290,N_1258);
nand U1360 (N_1360,N_1235,N_1262);
nand U1361 (N_1361,N_1271,N_1221);
or U1362 (N_1362,N_1266,N_1292);
or U1363 (N_1363,N_1216,N_1271);
nor U1364 (N_1364,N_1246,N_1252);
and U1365 (N_1365,N_1274,N_1265);
and U1366 (N_1366,N_1253,N_1280);
nand U1367 (N_1367,N_1239,N_1297);
and U1368 (N_1368,N_1204,N_1216);
and U1369 (N_1369,N_1289,N_1240);
or U1370 (N_1370,N_1202,N_1250);
nor U1371 (N_1371,N_1298,N_1226);
nand U1372 (N_1372,N_1239,N_1216);
and U1373 (N_1373,N_1228,N_1212);
nor U1374 (N_1374,N_1240,N_1205);
and U1375 (N_1375,N_1286,N_1217);
nand U1376 (N_1376,N_1221,N_1274);
and U1377 (N_1377,N_1231,N_1259);
nor U1378 (N_1378,N_1247,N_1286);
and U1379 (N_1379,N_1205,N_1247);
or U1380 (N_1380,N_1242,N_1298);
or U1381 (N_1381,N_1206,N_1265);
and U1382 (N_1382,N_1283,N_1294);
and U1383 (N_1383,N_1219,N_1231);
and U1384 (N_1384,N_1267,N_1229);
nand U1385 (N_1385,N_1260,N_1285);
and U1386 (N_1386,N_1281,N_1246);
nand U1387 (N_1387,N_1246,N_1280);
nor U1388 (N_1388,N_1208,N_1222);
and U1389 (N_1389,N_1245,N_1294);
nand U1390 (N_1390,N_1285,N_1277);
or U1391 (N_1391,N_1290,N_1237);
or U1392 (N_1392,N_1231,N_1247);
or U1393 (N_1393,N_1223,N_1293);
nor U1394 (N_1394,N_1211,N_1210);
nor U1395 (N_1395,N_1265,N_1230);
nor U1396 (N_1396,N_1273,N_1229);
nor U1397 (N_1397,N_1241,N_1209);
or U1398 (N_1398,N_1296,N_1200);
nor U1399 (N_1399,N_1278,N_1282);
nor U1400 (N_1400,N_1319,N_1324);
and U1401 (N_1401,N_1307,N_1396);
nor U1402 (N_1402,N_1326,N_1325);
nand U1403 (N_1403,N_1386,N_1303);
or U1404 (N_1404,N_1370,N_1381);
xor U1405 (N_1405,N_1328,N_1360);
xor U1406 (N_1406,N_1356,N_1398);
or U1407 (N_1407,N_1348,N_1388);
nor U1408 (N_1408,N_1380,N_1342);
nand U1409 (N_1409,N_1320,N_1317);
and U1410 (N_1410,N_1366,N_1301);
and U1411 (N_1411,N_1392,N_1397);
or U1412 (N_1412,N_1321,N_1332);
and U1413 (N_1413,N_1350,N_1345);
and U1414 (N_1414,N_1336,N_1372);
or U1415 (N_1415,N_1327,N_1375);
nor U1416 (N_1416,N_1318,N_1344);
nand U1417 (N_1417,N_1347,N_1346);
or U1418 (N_1418,N_1349,N_1353);
and U1419 (N_1419,N_1313,N_1352);
nor U1420 (N_1420,N_1393,N_1385);
and U1421 (N_1421,N_1331,N_1383);
or U1422 (N_1422,N_1322,N_1377);
nand U1423 (N_1423,N_1389,N_1369);
or U1424 (N_1424,N_1358,N_1365);
nand U1425 (N_1425,N_1311,N_1305);
nor U1426 (N_1426,N_1338,N_1395);
xnor U1427 (N_1427,N_1390,N_1382);
and U1428 (N_1428,N_1359,N_1363);
nand U1429 (N_1429,N_1373,N_1351);
nand U1430 (N_1430,N_1340,N_1354);
nand U1431 (N_1431,N_1355,N_1341);
nand U1432 (N_1432,N_1361,N_1310);
and U1433 (N_1433,N_1308,N_1323);
nand U1434 (N_1434,N_1368,N_1302);
and U1435 (N_1435,N_1399,N_1357);
nand U1436 (N_1436,N_1371,N_1309);
nor U1437 (N_1437,N_1394,N_1337);
or U1438 (N_1438,N_1300,N_1306);
and U1439 (N_1439,N_1330,N_1364);
or U1440 (N_1440,N_1391,N_1315);
xnor U1441 (N_1441,N_1314,N_1376);
or U1442 (N_1442,N_1312,N_1374);
nor U1443 (N_1443,N_1387,N_1379);
or U1444 (N_1444,N_1333,N_1334);
and U1445 (N_1445,N_1329,N_1316);
xor U1446 (N_1446,N_1343,N_1339);
and U1447 (N_1447,N_1304,N_1384);
nor U1448 (N_1448,N_1335,N_1378);
nor U1449 (N_1449,N_1367,N_1362);
nor U1450 (N_1450,N_1321,N_1343);
and U1451 (N_1451,N_1340,N_1353);
and U1452 (N_1452,N_1311,N_1371);
and U1453 (N_1453,N_1351,N_1333);
and U1454 (N_1454,N_1348,N_1322);
nor U1455 (N_1455,N_1366,N_1328);
nand U1456 (N_1456,N_1300,N_1354);
and U1457 (N_1457,N_1338,N_1394);
nand U1458 (N_1458,N_1357,N_1331);
nand U1459 (N_1459,N_1372,N_1335);
nor U1460 (N_1460,N_1305,N_1321);
and U1461 (N_1461,N_1393,N_1332);
nor U1462 (N_1462,N_1352,N_1353);
nor U1463 (N_1463,N_1316,N_1370);
or U1464 (N_1464,N_1381,N_1396);
or U1465 (N_1465,N_1302,N_1341);
nor U1466 (N_1466,N_1393,N_1368);
nand U1467 (N_1467,N_1343,N_1340);
nor U1468 (N_1468,N_1381,N_1318);
and U1469 (N_1469,N_1396,N_1338);
nand U1470 (N_1470,N_1361,N_1353);
nor U1471 (N_1471,N_1366,N_1359);
nand U1472 (N_1472,N_1312,N_1380);
nor U1473 (N_1473,N_1311,N_1347);
or U1474 (N_1474,N_1310,N_1356);
nor U1475 (N_1475,N_1381,N_1311);
and U1476 (N_1476,N_1343,N_1383);
nand U1477 (N_1477,N_1399,N_1350);
nor U1478 (N_1478,N_1399,N_1337);
nor U1479 (N_1479,N_1399,N_1318);
or U1480 (N_1480,N_1340,N_1302);
nand U1481 (N_1481,N_1353,N_1375);
and U1482 (N_1482,N_1349,N_1365);
nor U1483 (N_1483,N_1354,N_1393);
nor U1484 (N_1484,N_1302,N_1327);
nand U1485 (N_1485,N_1358,N_1370);
or U1486 (N_1486,N_1302,N_1380);
and U1487 (N_1487,N_1347,N_1382);
nand U1488 (N_1488,N_1372,N_1338);
nor U1489 (N_1489,N_1313,N_1394);
xor U1490 (N_1490,N_1390,N_1337);
nor U1491 (N_1491,N_1383,N_1384);
nor U1492 (N_1492,N_1331,N_1376);
nand U1493 (N_1493,N_1308,N_1392);
and U1494 (N_1494,N_1396,N_1360);
or U1495 (N_1495,N_1364,N_1319);
nand U1496 (N_1496,N_1345,N_1394);
and U1497 (N_1497,N_1385,N_1333);
nand U1498 (N_1498,N_1318,N_1364);
and U1499 (N_1499,N_1370,N_1395);
nor U1500 (N_1500,N_1414,N_1433);
nor U1501 (N_1501,N_1444,N_1452);
nand U1502 (N_1502,N_1417,N_1439);
and U1503 (N_1503,N_1474,N_1462);
and U1504 (N_1504,N_1436,N_1437);
and U1505 (N_1505,N_1415,N_1456);
nand U1506 (N_1506,N_1478,N_1411);
or U1507 (N_1507,N_1485,N_1491);
nor U1508 (N_1508,N_1422,N_1489);
nor U1509 (N_1509,N_1459,N_1492);
nor U1510 (N_1510,N_1453,N_1487);
nand U1511 (N_1511,N_1428,N_1480);
nor U1512 (N_1512,N_1470,N_1403);
or U1513 (N_1513,N_1451,N_1412);
or U1514 (N_1514,N_1461,N_1494);
nor U1515 (N_1515,N_1438,N_1471);
nand U1516 (N_1516,N_1407,N_1455);
and U1517 (N_1517,N_1457,N_1473);
or U1518 (N_1518,N_1429,N_1418);
nor U1519 (N_1519,N_1441,N_1469);
or U1520 (N_1520,N_1405,N_1497);
nand U1521 (N_1521,N_1495,N_1435);
nand U1522 (N_1522,N_1488,N_1481);
or U1523 (N_1523,N_1404,N_1431);
xor U1524 (N_1524,N_1413,N_1427);
and U1525 (N_1525,N_1416,N_1410);
nor U1526 (N_1526,N_1464,N_1424);
nor U1527 (N_1527,N_1493,N_1442);
nand U1528 (N_1528,N_1476,N_1401);
nand U1529 (N_1529,N_1434,N_1420);
and U1530 (N_1530,N_1447,N_1409);
nand U1531 (N_1531,N_1430,N_1498);
xor U1532 (N_1532,N_1458,N_1440);
or U1533 (N_1533,N_1490,N_1475);
and U1534 (N_1534,N_1477,N_1483);
or U1535 (N_1535,N_1425,N_1446);
nand U1536 (N_1536,N_1406,N_1450);
nand U1537 (N_1537,N_1426,N_1496);
nand U1538 (N_1538,N_1499,N_1408);
and U1539 (N_1539,N_1421,N_1460);
nand U1540 (N_1540,N_1443,N_1445);
nor U1541 (N_1541,N_1465,N_1484);
and U1542 (N_1542,N_1482,N_1400);
and U1543 (N_1543,N_1468,N_1402);
and U1544 (N_1544,N_1479,N_1463);
nor U1545 (N_1545,N_1419,N_1454);
and U1546 (N_1546,N_1466,N_1486);
and U1547 (N_1547,N_1423,N_1472);
and U1548 (N_1548,N_1449,N_1448);
nand U1549 (N_1549,N_1432,N_1467);
nor U1550 (N_1550,N_1401,N_1497);
nor U1551 (N_1551,N_1498,N_1464);
xnor U1552 (N_1552,N_1452,N_1489);
nand U1553 (N_1553,N_1421,N_1436);
or U1554 (N_1554,N_1454,N_1472);
nand U1555 (N_1555,N_1474,N_1409);
nand U1556 (N_1556,N_1420,N_1482);
nand U1557 (N_1557,N_1440,N_1443);
nand U1558 (N_1558,N_1492,N_1488);
nor U1559 (N_1559,N_1401,N_1423);
or U1560 (N_1560,N_1417,N_1456);
or U1561 (N_1561,N_1409,N_1492);
or U1562 (N_1562,N_1462,N_1446);
nor U1563 (N_1563,N_1495,N_1462);
nand U1564 (N_1564,N_1401,N_1440);
and U1565 (N_1565,N_1479,N_1401);
nand U1566 (N_1566,N_1408,N_1420);
or U1567 (N_1567,N_1423,N_1443);
or U1568 (N_1568,N_1448,N_1434);
nor U1569 (N_1569,N_1459,N_1438);
nand U1570 (N_1570,N_1478,N_1455);
nor U1571 (N_1571,N_1465,N_1439);
or U1572 (N_1572,N_1495,N_1488);
nand U1573 (N_1573,N_1483,N_1427);
nand U1574 (N_1574,N_1420,N_1450);
and U1575 (N_1575,N_1483,N_1470);
or U1576 (N_1576,N_1452,N_1486);
nor U1577 (N_1577,N_1441,N_1447);
or U1578 (N_1578,N_1428,N_1494);
nand U1579 (N_1579,N_1496,N_1442);
or U1580 (N_1580,N_1452,N_1439);
nand U1581 (N_1581,N_1474,N_1463);
nor U1582 (N_1582,N_1432,N_1430);
nor U1583 (N_1583,N_1492,N_1491);
or U1584 (N_1584,N_1425,N_1417);
nand U1585 (N_1585,N_1493,N_1452);
and U1586 (N_1586,N_1475,N_1434);
nand U1587 (N_1587,N_1462,N_1420);
and U1588 (N_1588,N_1459,N_1457);
and U1589 (N_1589,N_1411,N_1467);
and U1590 (N_1590,N_1487,N_1469);
and U1591 (N_1591,N_1428,N_1448);
and U1592 (N_1592,N_1457,N_1431);
nor U1593 (N_1593,N_1467,N_1485);
nor U1594 (N_1594,N_1493,N_1453);
xor U1595 (N_1595,N_1447,N_1495);
nor U1596 (N_1596,N_1406,N_1444);
xnor U1597 (N_1597,N_1403,N_1488);
nor U1598 (N_1598,N_1499,N_1436);
or U1599 (N_1599,N_1471,N_1448);
nor U1600 (N_1600,N_1582,N_1566);
and U1601 (N_1601,N_1548,N_1529);
nand U1602 (N_1602,N_1528,N_1569);
nor U1603 (N_1603,N_1524,N_1539);
or U1604 (N_1604,N_1592,N_1511);
or U1605 (N_1605,N_1580,N_1573);
nand U1606 (N_1606,N_1554,N_1515);
and U1607 (N_1607,N_1560,N_1501);
and U1608 (N_1608,N_1537,N_1500);
or U1609 (N_1609,N_1577,N_1513);
or U1610 (N_1610,N_1543,N_1507);
nand U1611 (N_1611,N_1535,N_1510);
and U1612 (N_1612,N_1541,N_1565);
nor U1613 (N_1613,N_1532,N_1545);
nor U1614 (N_1614,N_1584,N_1595);
and U1615 (N_1615,N_1579,N_1512);
nand U1616 (N_1616,N_1570,N_1527);
and U1617 (N_1617,N_1514,N_1509);
nand U1618 (N_1618,N_1557,N_1564);
nor U1619 (N_1619,N_1522,N_1556);
nand U1620 (N_1620,N_1567,N_1526);
nor U1621 (N_1621,N_1517,N_1505);
nor U1622 (N_1622,N_1594,N_1519);
nand U1623 (N_1623,N_1587,N_1551);
nand U1624 (N_1624,N_1503,N_1588);
and U1625 (N_1625,N_1598,N_1534);
nor U1626 (N_1626,N_1596,N_1597);
nand U1627 (N_1627,N_1531,N_1568);
or U1628 (N_1628,N_1506,N_1571);
and U1629 (N_1629,N_1544,N_1574);
or U1630 (N_1630,N_1525,N_1593);
nor U1631 (N_1631,N_1561,N_1575);
nor U1632 (N_1632,N_1547,N_1550);
nand U1633 (N_1633,N_1599,N_1536);
nor U1634 (N_1634,N_1559,N_1523);
nor U1635 (N_1635,N_1590,N_1585);
or U1636 (N_1636,N_1533,N_1562);
and U1637 (N_1637,N_1549,N_1583);
nand U1638 (N_1638,N_1518,N_1502);
and U1639 (N_1639,N_1504,N_1563);
nand U1640 (N_1640,N_1553,N_1516);
nor U1641 (N_1641,N_1538,N_1581);
nor U1642 (N_1642,N_1530,N_1508);
or U1643 (N_1643,N_1589,N_1552);
nand U1644 (N_1644,N_1576,N_1521);
nand U1645 (N_1645,N_1558,N_1540);
nor U1646 (N_1646,N_1520,N_1546);
or U1647 (N_1647,N_1555,N_1572);
nor U1648 (N_1648,N_1591,N_1542);
and U1649 (N_1649,N_1586,N_1578);
nand U1650 (N_1650,N_1544,N_1506);
nand U1651 (N_1651,N_1597,N_1508);
and U1652 (N_1652,N_1569,N_1584);
nand U1653 (N_1653,N_1554,N_1588);
nor U1654 (N_1654,N_1540,N_1572);
or U1655 (N_1655,N_1585,N_1575);
and U1656 (N_1656,N_1571,N_1547);
and U1657 (N_1657,N_1528,N_1577);
nor U1658 (N_1658,N_1581,N_1542);
or U1659 (N_1659,N_1588,N_1515);
or U1660 (N_1660,N_1574,N_1535);
and U1661 (N_1661,N_1540,N_1539);
or U1662 (N_1662,N_1531,N_1521);
or U1663 (N_1663,N_1515,N_1582);
nand U1664 (N_1664,N_1528,N_1554);
nor U1665 (N_1665,N_1560,N_1527);
nand U1666 (N_1666,N_1537,N_1503);
nand U1667 (N_1667,N_1514,N_1534);
xor U1668 (N_1668,N_1580,N_1594);
nor U1669 (N_1669,N_1595,N_1596);
nor U1670 (N_1670,N_1553,N_1542);
or U1671 (N_1671,N_1595,N_1519);
or U1672 (N_1672,N_1513,N_1533);
or U1673 (N_1673,N_1548,N_1526);
and U1674 (N_1674,N_1561,N_1526);
nor U1675 (N_1675,N_1546,N_1575);
and U1676 (N_1676,N_1581,N_1570);
nor U1677 (N_1677,N_1561,N_1531);
and U1678 (N_1678,N_1569,N_1522);
nor U1679 (N_1679,N_1532,N_1501);
and U1680 (N_1680,N_1568,N_1526);
and U1681 (N_1681,N_1505,N_1534);
and U1682 (N_1682,N_1576,N_1541);
or U1683 (N_1683,N_1549,N_1515);
and U1684 (N_1684,N_1536,N_1566);
nor U1685 (N_1685,N_1501,N_1506);
nor U1686 (N_1686,N_1594,N_1576);
nor U1687 (N_1687,N_1508,N_1558);
nor U1688 (N_1688,N_1597,N_1577);
nand U1689 (N_1689,N_1591,N_1548);
and U1690 (N_1690,N_1558,N_1591);
or U1691 (N_1691,N_1520,N_1599);
and U1692 (N_1692,N_1577,N_1506);
or U1693 (N_1693,N_1533,N_1547);
and U1694 (N_1694,N_1502,N_1591);
nand U1695 (N_1695,N_1564,N_1598);
or U1696 (N_1696,N_1585,N_1549);
nand U1697 (N_1697,N_1529,N_1530);
and U1698 (N_1698,N_1591,N_1568);
nand U1699 (N_1699,N_1576,N_1560);
or U1700 (N_1700,N_1691,N_1647);
and U1701 (N_1701,N_1646,N_1609);
and U1702 (N_1702,N_1624,N_1645);
nand U1703 (N_1703,N_1614,N_1686);
nand U1704 (N_1704,N_1663,N_1676);
and U1705 (N_1705,N_1620,N_1627);
or U1706 (N_1706,N_1655,N_1641);
and U1707 (N_1707,N_1658,N_1619);
nor U1708 (N_1708,N_1694,N_1637);
nor U1709 (N_1709,N_1654,N_1602);
nor U1710 (N_1710,N_1621,N_1622);
nor U1711 (N_1711,N_1634,N_1652);
and U1712 (N_1712,N_1687,N_1631);
or U1713 (N_1713,N_1604,N_1681);
and U1714 (N_1714,N_1612,N_1640);
nor U1715 (N_1715,N_1615,N_1625);
or U1716 (N_1716,N_1664,N_1638);
nand U1717 (N_1717,N_1607,N_1673);
xnor U1718 (N_1718,N_1608,N_1660);
or U1719 (N_1719,N_1618,N_1693);
or U1720 (N_1720,N_1610,N_1656);
nand U1721 (N_1721,N_1626,N_1674);
nand U1722 (N_1722,N_1613,N_1689);
nand U1723 (N_1723,N_1678,N_1682);
nor U1724 (N_1724,N_1670,N_1683);
nor U1725 (N_1725,N_1659,N_1657);
nor U1726 (N_1726,N_1648,N_1636);
nor U1727 (N_1727,N_1672,N_1667);
or U1728 (N_1728,N_1688,N_1629);
nand U1729 (N_1729,N_1639,N_1675);
and U1730 (N_1730,N_1635,N_1603);
or U1731 (N_1731,N_1679,N_1698);
nand U1732 (N_1732,N_1617,N_1671);
nor U1733 (N_1733,N_1606,N_1605);
nor U1734 (N_1734,N_1662,N_1685);
or U1735 (N_1735,N_1661,N_1677);
nand U1736 (N_1736,N_1623,N_1611);
or U1737 (N_1737,N_1616,N_1697);
and U1738 (N_1738,N_1644,N_1643);
or U1739 (N_1739,N_1630,N_1690);
and U1740 (N_1740,N_1601,N_1653);
and U1741 (N_1741,N_1633,N_1669);
and U1742 (N_1742,N_1651,N_1665);
nand U1743 (N_1743,N_1632,N_1684);
and U1744 (N_1744,N_1695,N_1666);
and U1745 (N_1745,N_1642,N_1699);
or U1746 (N_1746,N_1696,N_1650);
or U1747 (N_1747,N_1680,N_1668);
nand U1748 (N_1748,N_1628,N_1692);
nor U1749 (N_1749,N_1649,N_1600);
or U1750 (N_1750,N_1602,N_1600);
or U1751 (N_1751,N_1678,N_1651);
or U1752 (N_1752,N_1672,N_1695);
nand U1753 (N_1753,N_1649,N_1655);
xnor U1754 (N_1754,N_1644,N_1646);
nor U1755 (N_1755,N_1615,N_1632);
and U1756 (N_1756,N_1692,N_1658);
and U1757 (N_1757,N_1684,N_1642);
and U1758 (N_1758,N_1622,N_1602);
nor U1759 (N_1759,N_1665,N_1671);
nand U1760 (N_1760,N_1675,N_1670);
and U1761 (N_1761,N_1686,N_1609);
nand U1762 (N_1762,N_1608,N_1604);
nand U1763 (N_1763,N_1692,N_1688);
nand U1764 (N_1764,N_1621,N_1681);
or U1765 (N_1765,N_1658,N_1670);
nor U1766 (N_1766,N_1608,N_1635);
and U1767 (N_1767,N_1658,N_1673);
nor U1768 (N_1768,N_1669,N_1620);
nand U1769 (N_1769,N_1628,N_1612);
nor U1770 (N_1770,N_1628,N_1696);
nand U1771 (N_1771,N_1621,N_1645);
or U1772 (N_1772,N_1626,N_1679);
nand U1773 (N_1773,N_1699,N_1670);
and U1774 (N_1774,N_1693,N_1652);
or U1775 (N_1775,N_1646,N_1601);
and U1776 (N_1776,N_1636,N_1661);
nand U1777 (N_1777,N_1607,N_1696);
and U1778 (N_1778,N_1606,N_1667);
nand U1779 (N_1779,N_1691,N_1658);
or U1780 (N_1780,N_1690,N_1603);
nor U1781 (N_1781,N_1620,N_1685);
nor U1782 (N_1782,N_1665,N_1622);
nand U1783 (N_1783,N_1641,N_1687);
or U1784 (N_1784,N_1698,N_1657);
nor U1785 (N_1785,N_1678,N_1634);
and U1786 (N_1786,N_1631,N_1640);
or U1787 (N_1787,N_1669,N_1674);
or U1788 (N_1788,N_1692,N_1693);
and U1789 (N_1789,N_1638,N_1634);
nor U1790 (N_1790,N_1629,N_1670);
nand U1791 (N_1791,N_1629,N_1683);
and U1792 (N_1792,N_1668,N_1677);
nand U1793 (N_1793,N_1625,N_1611);
nor U1794 (N_1794,N_1693,N_1676);
nor U1795 (N_1795,N_1600,N_1638);
nand U1796 (N_1796,N_1664,N_1690);
nor U1797 (N_1797,N_1685,N_1657);
nand U1798 (N_1798,N_1660,N_1683);
and U1799 (N_1799,N_1698,N_1691);
nand U1800 (N_1800,N_1769,N_1776);
and U1801 (N_1801,N_1775,N_1719);
or U1802 (N_1802,N_1758,N_1780);
nor U1803 (N_1803,N_1793,N_1774);
or U1804 (N_1804,N_1754,N_1788);
nand U1805 (N_1805,N_1796,N_1743);
or U1806 (N_1806,N_1742,N_1786);
and U1807 (N_1807,N_1746,N_1701);
nand U1808 (N_1808,N_1762,N_1777);
or U1809 (N_1809,N_1722,N_1713);
and U1810 (N_1810,N_1711,N_1771);
nand U1811 (N_1811,N_1795,N_1726);
nand U1812 (N_1812,N_1751,N_1706);
or U1813 (N_1813,N_1724,N_1772);
nor U1814 (N_1814,N_1759,N_1705);
nand U1815 (N_1815,N_1753,N_1782);
or U1816 (N_1816,N_1717,N_1716);
or U1817 (N_1817,N_1712,N_1708);
nor U1818 (N_1818,N_1791,N_1799);
nand U1819 (N_1819,N_1749,N_1738);
nand U1820 (N_1820,N_1709,N_1792);
or U1821 (N_1821,N_1757,N_1733);
nand U1822 (N_1822,N_1764,N_1721);
nor U1823 (N_1823,N_1740,N_1731);
and U1824 (N_1824,N_1723,N_1730);
and U1825 (N_1825,N_1715,N_1770);
nor U1826 (N_1826,N_1781,N_1761);
and U1827 (N_1827,N_1735,N_1736);
or U1828 (N_1828,N_1741,N_1729);
or U1829 (N_1829,N_1703,N_1702);
nor U1830 (N_1830,N_1720,N_1778);
xnor U1831 (N_1831,N_1779,N_1750);
nor U1832 (N_1832,N_1784,N_1760);
xor U1833 (N_1833,N_1714,N_1748);
and U1834 (N_1834,N_1745,N_1766);
and U1835 (N_1835,N_1789,N_1728);
or U1836 (N_1836,N_1734,N_1783);
nor U1837 (N_1837,N_1707,N_1763);
or U1838 (N_1838,N_1790,N_1794);
nor U1839 (N_1839,N_1756,N_1765);
and U1840 (N_1840,N_1732,N_1704);
nand U1841 (N_1841,N_1785,N_1727);
nor U1842 (N_1842,N_1737,N_1798);
or U1843 (N_1843,N_1797,N_1718);
xor U1844 (N_1844,N_1752,N_1768);
nor U1845 (N_1845,N_1744,N_1700);
nand U1846 (N_1846,N_1747,N_1787);
nand U1847 (N_1847,N_1767,N_1773);
and U1848 (N_1848,N_1710,N_1739);
nor U1849 (N_1849,N_1725,N_1755);
or U1850 (N_1850,N_1791,N_1797);
and U1851 (N_1851,N_1716,N_1798);
and U1852 (N_1852,N_1779,N_1715);
nor U1853 (N_1853,N_1708,N_1749);
nand U1854 (N_1854,N_1758,N_1715);
or U1855 (N_1855,N_1748,N_1750);
and U1856 (N_1856,N_1757,N_1782);
or U1857 (N_1857,N_1746,N_1713);
nand U1858 (N_1858,N_1797,N_1733);
or U1859 (N_1859,N_1703,N_1726);
nand U1860 (N_1860,N_1783,N_1700);
or U1861 (N_1861,N_1777,N_1720);
or U1862 (N_1862,N_1702,N_1737);
or U1863 (N_1863,N_1760,N_1709);
and U1864 (N_1864,N_1783,N_1769);
or U1865 (N_1865,N_1730,N_1797);
nor U1866 (N_1866,N_1785,N_1732);
or U1867 (N_1867,N_1749,N_1703);
nand U1868 (N_1868,N_1799,N_1734);
nand U1869 (N_1869,N_1710,N_1765);
nor U1870 (N_1870,N_1747,N_1740);
xnor U1871 (N_1871,N_1750,N_1771);
or U1872 (N_1872,N_1777,N_1755);
nor U1873 (N_1873,N_1731,N_1709);
and U1874 (N_1874,N_1754,N_1752);
nor U1875 (N_1875,N_1700,N_1742);
nor U1876 (N_1876,N_1765,N_1763);
and U1877 (N_1877,N_1727,N_1730);
and U1878 (N_1878,N_1776,N_1782);
and U1879 (N_1879,N_1719,N_1735);
or U1880 (N_1880,N_1780,N_1712);
or U1881 (N_1881,N_1754,N_1767);
nand U1882 (N_1882,N_1789,N_1746);
nand U1883 (N_1883,N_1720,N_1773);
nand U1884 (N_1884,N_1718,N_1777);
or U1885 (N_1885,N_1737,N_1754);
nor U1886 (N_1886,N_1777,N_1789);
nand U1887 (N_1887,N_1765,N_1789);
or U1888 (N_1888,N_1789,N_1787);
nor U1889 (N_1889,N_1745,N_1729);
or U1890 (N_1890,N_1775,N_1714);
and U1891 (N_1891,N_1795,N_1791);
nor U1892 (N_1892,N_1799,N_1764);
nand U1893 (N_1893,N_1741,N_1781);
nor U1894 (N_1894,N_1777,N_1771);
or U1895 (N_1895,N_1787,N_1786);
and U1896 (N_1896,N_1715,N_1713);
or U1897 (N_1897,N_1701,N_1707);
nand U1898 (N_1898,N_1781,N_1760);
or U1899 (N_1899,N_1755,N_1719);
nor U1900 (N_1900,N_1897,N_1829);
nor U1901 (N_1901,N_1867,N_1800);
xor U1902 (N_1902,N_1865,N_1871);
and U1903 (N_1903,N_1888,N_1819);
nand U1904 (N_1904,N_1853,N_1828);
nor U1905 (N_1905,N_1850,N_1857);
or U1906 (N_1906,N_1846,N_1814);
or U1907 (N_1907,N_1862,N_1823);
or U1908 (N_1908,N_1856,N_1801);
or U1909 (N_1909,N_1815,N_1825);
nand U1910 (N_1910,N_1899,N_1838);
nand U1911 (N_1911,N_1859,N_1834);
and U1912 (N_1912,N_1893,N_1891);
nor U1913 (N_1913,N_1855,N_1887);
or U1914 (N_1914,N_1863,N_1876);
and U1915 (N_1915,N_1848,N_1852);
nor U1916 (N_1916,N_1811,N_1874);
or U1917 (N_1917,N_1824,N_1896);
nor U1918 (N_1918,N_1880,N_1817);
nand U1919 (N_1919,N_1847,N_1873);
nor U1920 (N_1920,N_1895,N_1861);
nand U1921 (N_1921,N_1872,N_1805);
nand U1922 (N_1922,N_1870,N_1826);
or U1923 (N_1923,N_1898,N_1808);
and U1924 (N_1924,N_1809,N_1882);
nand U1925 (N_1925,N_1875,N_1851);
and U1926 (N_1926,N_1818,N_1835);
or U1927 (N_1927,N_1830,N_1868);
nand U1928 (N_1928,N_1849,N_1816);
nand U1929 (N_1929,N_1878,N_1854);
nand U1930 (N_1930,N_1841,N_1869);
nor U1931 (N_1931,N_1813,N_1845);
or U1932 (N_1932,N_1822,N_1884);
nor U1933 (N_1933,N_1803,N_1885);
or U1934 (N_1934,N_1894,N_1802);
or U1935 (N_1935,N_1839,N_1833);
xor U1936 (N_1936,N_1842,N_1827);
nor U1937 (N_1937,N_1807,N_1840);
nor U1938 (N_1938,N_1804,N_1821);
xnor U1939 (N_1939,N_1883,N_1864);
and U1940 (N_1940,N_1881,N_1837);
xnor U1941 (N_1941,N_1806,N_1832);
nand U1942 (N_1942,N_1892,N_1890);
or U1943 (N_1943,N_1831,N_1810);
and U1944 (N_1944,N_1886,N_1889);
or U1945 (N_1945,N_1858,N_1812);
nand U1946 (N_1946,N_1844,N_1877);
nor U1947 (N_1947,N_1866,N_1836);
nor U1948 (N_1948,N_1843,N_1879);
or U1949 (N_1949,N_1820,N_1860);
nor U1950 (N_1950,N_1857,N_1863);
nand U1951 (N_1951,N_1802,N_1833);
nand U1952 (N_1952,N_1810,N_1888);
or U1953 (N_1953,N_1840,N_1835);
nor U1954 (N_1954,N_1848,N_1827);
nand U1955 (N_1955,N_1849,N_1858);
xnor U1956 (N_1956,N_1817,N_1815);
nand U1957 (N_1957,N_1802,N_1837);
or U1958 (N_1958,N_1846,N_1867);
xnor U1959 (N_1959,N_1840,N_1865);
nor U1960 (N_1960,N_1831,N_1839);
or U1961 (N_1961,N_1887,N_1835);
nand U1962 (N_1962,N_1839,N_1850);
and U1963 (N_1963,N_1827,N_1850);
nand U1964 (N_1964,N_1892,N_1872);
nor U1965 (N_1965,N_1856,N_1815);
or U1966 (N_1966,N_1855,N_1844);
nor U1967 (N_1967,N_1866,N_1888);
nor U1968 (N_1968,N_1844,N_1885);
xnor U1969 (N_1969,N_1869,N_1871);
and U1970 (N_1970,N_1803,N_1860);
and U1971 (N_1971,N_1873,N_1860);
nand U1972 (N_1972,N_1866,N_1823);
and U1973 (N_1973,N_1868,N_1893);
or U1974 (N_1974,N_1836,N_1850);
nand U1975 (N_1975,N_1829,N_1899);
nor U1976 (N_1976,N_1863,N_1866);
nor U1977 (N_1977,N_1873,N_1894);
nor U1978 (N_1978,N_1844,N_1818);
nand U1979 (N_1979,N_1895,N_1858);
xnor U1980 (N_1980,N_1852,N_1861);
nand U1981 (N_1981,N_1855,N_1833);
nor U1982 (N_1982,N_1897,N_1848);
or U1983 (N_1983,N_1898,N_1899);
or U1984 (N_1984,N_1872,N_1823);
and U1985 (N_1985,N_1826,N_1842);
and U1986 (N_1986,N_1869,N_1893);
nand U1987 (N_1987,N_1857,N_1802);
or U1988 (N_1988,N_1891,N_1801);
nand U1989 (N_1989,N_1840,N_1824);
and U1990 (N_1990,N_1844,N_1825);
and U1991 (N_1991,N_1832,N_1873);
nor U1992 (N_1992,N_1845,N_1870);
nor U1993 (N_1993,N_1861,N_1805);
nor U1994 (N_1994,N_1846,N_1845);
nor U1995 (N_1995,N_1810,N_1813);
nand U1996 (N_1996,N_1850,N_1826);
and U1997 (N_1997,N_1824,N_1894);
xnor U1998 (N_1998,N_1878,N_1813);
or U1999 (N_1999,N_1804,N_1835);
nor U2000 (N_2000,N_1907,N_1920);
nand U2001 (N_2001,N_1931,N_1988);
and U2002 (N_2002,N_1937,N_1930);
and U2003 (N_2003,N_1940,N_1966);
nand U2004 (N_2004,N_1904,N_1906);
nor U2005 (N_2005,N_1963,N_1955);
nand U2006 (N_2006,N_1994,N_1929);
nand U2007 (N_2007,N_1989,N_1900);
nand U2008 (N_2008,N_1945,N_1948);
and U2009 (N_2009,N_1978,N_1984);
or U2010 (N_2010,N_1990,N_1916);
nor U2011 (N_2011,N_1949,N_1918);
nand U2012 (N_2012,N_1997,N_1908);
and U2013 (N_2013,N_1968,N_1934);
nor U2014 (N_2014,N_1912,N_1921);
nor U2015 (N_2015,N_1922,N_1951);
and U2016 (N_2016,N_1952,N_1925);
nor U2017 (N_2017,N_1991,N_1961);
and U2018 (N_2018,N_1996,N_1999);
nor U2019 (N_2019,N_1950,N_1902);
nor U2020 (N_2020,N_1976,N_1973);
or U2021 (N_2021,N_1965,N_1992);
nor U2022 (N_2022,N_1915,N_1932);
nand U2023 (N_2023,N_1985,N_1998);
nand U2024 (N_2024,N_1964,N_1981);
nor U2025 (N_2025,N_1911,N_1972);
xor U2026 (N_2026,N_1935,N_1962);
nor U2027 (N_2027,N_1917,N_1946);
or U2028 (N_2028,N_1905,N_1969);
nor U2029 (N_2029,N_1919,N_1939);
or U2030 (N_2030,N_1980,N_1943);
nor U2031 (N_2031,N_1910,N_1923);
nor U2032 (N_2032,N_1982,N_1928);
nand U2033 (N_2033,N_1903,N_1970);
and U2034 (N_2034,N_1914,N_1979);
nand U2035 (N_2035,N_1958,N_1927);
and U2036 (N_2036,N_1936,N_1901);
nor U2037 (N_2037,N_1971,N_1913);
nand U2038 (N_2038,N_1926,N_1960);
or U2039 (N_2039,N_1924,N_1967);
and U2040 (N_2040,N_1975,N_1947);
or U2041 (N_2041,N_1983,N_1938);
nor U2042 (N_2042,N_1959,N_1986);
nand U2043 (N_2043,N_1944,N_1977);
nand U2044 (N_2044,N_1957,N_1993);
and U2045 (N_2045,N_1995,N_1954);
nor U2046 (N_2046,N_1941,N_1933);
nand U2047 (N_2047,N_1909,N_1987);
or U2048 (N_2048,N_1974,N_1953);
or U2049 (N_2049,N_1956,N_1942);
nor U2050 (N_2050,N_1907,N_1909);
nand U2051 (N_2051,N_1995,N_1914);
and U2052 (N_2052,N_1982,N_1950);
and U2053 (N_2053,N_1955,N_1990);
nand U2054 (N_2054,N_1980,N_1982);
nand U2055 (N_2055,N_1914,N_1985);
xor U2056 (N_2056,N_1909,N_1981);
nor U2057 (N_2057,N_1986,N_1973);
and U2058 (N_2058,N_1935,N_1987);
nand U2059 (N_2059,N_1933,N_1997);
nor U2060 (N_2060,N_1932,N_1918);
nor U2061 (N_2061,N_1982,N_1906);
or U2062 (N_2062,N_1901,N_1949);
or U2063 (N_2063,N_1921,N_1987);
or U2064 (N_2064,N_1995,N_1909);
and U2065 (N_2065,N_1917,N_1930);
xor U2066 (N_2066,N_1920,N_1987);
and U2067 (N_2067,N_1917,N_1985);
or U2068 (N_2068,N_1921,N_1937);
nand U2069 (N_2069,N_1972,N_1926);
or U2070 (N_2070,N_1914,N_1948);
nor U2071 (N_2071,N_1921,N_1922);
nand U2072 (N_2072,N_1925,N_1937);
and U2073 (N_2073,N_1933,N_1989);
nor U2074 (N_2074,N_1943,N_1978);
or U2075 (N_2075,N_1925,N_1942);
nor U2076 (N_2076,N_1983,N_1951);
nor U2077 (N_2077,N_1934,N_1913);
and U2078 (N_2078,N_1935,N_1950);
nand U2079 (N_2079,N_1972,N_1901);
or U2080 (N_2080,N_1946,N_1904);
or U2081 (N_2081,N_1902,N_1931);
nand U2082 (N_2082,N_1903,N_1937);
nor U2083 (N_2083,N_1909,N_1914);
and U2084 (N_2084,N_1955,N_1960);
xnor U2085 (N_2085,N_1920,N_1941);
or U2086 (N_2086,N_1950,N_1988);
nor U2087 (N_2087,N_1910,N_1955);
or U2088 (N_2088,N_1996,N_1912);
and U2089 (N_2089,N_1945,N_1997);
or U2090 (N_2090,N_1988,N_1939);
or U2091 (N_2091,N_1964,N_1936);
or U2092 (N_2092,N_1949,N_1956);
or U2093 (N_2093,N_1938,N_1969);
xor U2094 (N_2094,N_1904,N_1963);
or U2095 (N_2095,N_1905,N_1980);
nor U2096 (N_2096,N_1934,N_1973);
nor U2097 (N_2097,N_1951,N_1960);
and U2098 (N_2098,N_1936,N_1965);
nor U2099 (N_2099,N_1965,N_1981);
nand U2100 (N_2100,N_2068,N_2002);
nand U2101 (N_2101,N_2030,N_2064);
nor U2102 (N_2102,N_2044,N_2013);
nor U2103 (N_2103,N_2062,N_2081);
or U2104 (N_2104,N_2040,N_2051);
nand U2105 (N_2105,N_2014,N_2053);
and U2106 (N_2106,N_2054,N_2074);
and U2107 (N_2107,N_2024,N_2034);
and U2108 (N_2108,N_2009,N_2088);
xnor U2109 (N_2109,N_2026,N_2071);
nor U2110 (N_2110,N_2097,N_2083);
nor U2111 (N_2111,N_2031,N_2058);
or U2112 (N_2112,N_2038,N_2085);
or U2113 (N_2113,N_2056,N_2045);
nand U2114 (N_2114,N_2022,N_2078);
nor U2115 (N_2115,N_2070,N_2039);
nor U2116 (N_2116,N_2066,N_2093);
or U2117 (N_2117,N_2089,N_2035);
nor U2118 (N_2118,N_2087,N_2023);
and U2119 (N_2119,N_2072,N_2092);
nand U2120 (N_2120,N_2096,N_2046);
xor U2121 (N_2121,N_2018,N_2032);
or U2122 (N_2122,N_2050,N_2079);
nand U2123 (N_2123,N_2042,N_2006);
and U2124 (N_2124,N_2061,N_2095);
or U2125 (N_2125,N_2052,N_2048);
nand U2126 (N_2126,N_2063,N_2057);
and U2127 (N_2127,N_2003,N_2033);
or U2128 (N_2128,N_2021,N_2047);
nand U2129 (N_2129,N_2094,N_2017);
or U2130 (N_2130,N_2076,N_2036);
and U2131 (N_2131,N_2025,N_2015);
and U2132 (N_2132,N_2098,N_2082);
nand U2133 (N_2133,N_2069,N_2055);
or U2134 (N_2134,N_2001,N_2059);
nor U2135 (N_2135,N_2067,N_2086);
and U2136 (N_2136,N_2011,N_2029);
nor U2137 (N_2137,N_2090,N_2027);
and U2138 (N_2138,N_2010,N_2016);
or U2139 (N_2139,N_2080,N_2008);
or U2140 (N_2140,N_2084,N_2077);
xor U2141 (N_2141,N_2000,N_2020);
or U2142 (N_2142,N_2065,N_2028);
nand U2143 (N_2143,N_2012,N_2073);
and U2144 (N_2144,N_2037,N_2007);
nor U2145 (N_2145,N_2004,N_2099);
nand U2146 (N_2146,N_2005,N_2091);
and U2147 (N_2147,N_2075,N_2041);
nand U2148 (N_2148,N_2060,N_2049);
or U2149 (N_2149,N_2019,N_2043);
nor U2150 (N_2150,N_2091,N_2092);
or U2151 (N_2151,N_2056,N_2024);
or U2152 (N_2152,N_2060,N_2020);
nor U2153 (N_2153,N_2081,N_2098);
nand U2154 (N_2154,N_2003,N_2090);
nand U2155 (N_2155,N_2050,N_2012);
nand U2156 (N_2156,N_2088,N_2043);
or U2157 (N_2157,N_2015,N_2047);
nor U2158 (N_2158,N_2044,N_2069);
or U2159 (N_2159,N_2026,N_2014);
nand U2160 (N_2160,N_2017,N_2016);
nand U2161 (N_2161,N_2035,N_2047);
or U2162 (N_2162,N_2017,N_2079);
nor U2163 (N_2163,N_2094,N_2070);
or U2164 (N_2164,N_2020,N_2024);
nand U2165 (N_2165,N_2055,N_2033);
or U2166 (N_2166,N_2094,N_2059);
nor U2167 (N_2167,N_2096,N_2081);
nand U2168 (N_2168,N_2098,N_2099);
nand U2169 (N_2169,N_2096,N_2066);
or U2170 (N_2170,N_2018,N_2082);
or U2171 (N_2171,N_2069,N_2019);
and U2172 (N_2172,N_2081,N_2061);
and U2173 (N_2173,N_2077,N_2056);
or U2174 (N_2174,N_2009,N_2029);
or U2175 (N_2175,N_2079,N_2020);
or U2176 (N_2176,N_2006,N_2056);
nor U2177 (N_2177,N_2099,N_2026);
or U2178 (N_2178,N_2074,N_2089);
nand U2179 (N_2179,N_2054,N_2053);
xor U2180 (N_2180,N_2074,N_2019);
nand U2181 (N_2181,N_2032,N_2074);
nor U2182 (N_2182,N_2017,N_2090);
nor U2183 (N_2183,N_2044,N_2087);
and U2184 (N_2184,N_2002,N_2059);
and U2185 (N_2185,N_2093,N_2024);
and U2186 (N_2186,N_2073,N_2097);
and U2187 (N_2187,N_2009,N_2012);
nand U2188 (N_2188,N_2073,N_2002);
nor U2189 (N_2189,N_2071,N_2014);
or U2190 (N_2190,N_2046,N_2083);
or U2191 (N_2191,N_2029,N_2049);
nor U2192 (N_2192,N_2035,N_2011);
nor U2193 (N_2193,N_2095,N_2010);
nor U2194 (N_2194,N_2028,N_2046);
or U2195 (N_2195,N_2016,N_2039);
nor U2196 (N_2196,N_2033,N_2062);
or U2197 (N_2197,N_2071,N_2053);
or U2198 (N_2198,N_2085,N_2067);
and U2199 (N_2199,N_2091,N_2020);
nor U2200 (N_2200,N_2109,N_2104);
and U2201 (N_2201,N_2106,N_2130);
nor U2202 (N_2202,N_2182,N_2199);
nor U2203 (N_2203,N_2175,N_2160);
and U2204 (N_2204,N_2108,N_2163);
and U2205 (N_2205,N_2131,N_2176);
and U2206 (N_2206,N_2113,N_2174);
xnor U2207 (N_2207,N_2183,N_2138);
or U2208 (N_2208,N_2137,N_2105);
and U2209 (N_2209,N_2124,N_2168);
or U2210 (N_2210,N_2147,N_2172);
nand U2211 (N_2211,N_2192,N_2122);
nand U2212 (N_2212,N_2136,N_2143);
nand U2213 (N_2213,N_2145,N_2120);
nor U2214 (N_2214,N_2165,N_2121);
or U2215 (N_2215,N_2158,N_2150);
nor U2216 (N_2216,N_2127,N_2141);
and U2217 (N_2217,N_2132,N_2129);
nor U2218 (N_2218,N_2134,N_2117);
nand U2219 (N_2219,N_2161,N_2178);
nor U2220 (N_2220,N_2125,N_2189);
xnor U2221 (N_2221,N_2167,N_2186);
or U2222 (N_2222,N_2191,N_2135);
and U2223 (N_2223,N_2133,N_2151);
and U2224 (N_2224,N_2103,N_2181);
and U2225 (N_2225,N_2126,N_2170);
or U2226 (N_2226,N_2196,N_2188);
or U2227 (N_2227,N_2173,N_2149);
or U2228 (N_2228,N_2197,N_2179);
or U2229 (N_2229,N_2157,N_2102);
nand U2230 (N_2230,N_2112,N_2140);
and U2231 (N_2231,N_2139,N_2198);
or U2232 (N_2232,N_2177,N_2184);
and U2233 (N_2233,N_2156,N_2171);
or U2234 (N_2234,N_2110,N_2195);
nor U2235 (N_2235,N_2159,N_2111);
or U2236 (N_2236,N_2116,N_2185);
nor U2237 (N_2237,N_2190,N_2180);
nor U2238 (N_2238,N_2100,N_2119);
or U2239 (N_2239,N_2193,N_2144);
and U2240 (N_2240,N_2107,N_2118);
or U2241 (N_2241,N_2146,N_2194);
or U2242 (N_2242,N_2166,N_2128);
nand U2243 (N_2243,N_2162,N_2169);
nor U2244 (N_2244,N_2114,N_2152);
nor U2245 (N_2245,N_2154,N_2115);
nand U2246 (N_2246,N_2153,N_2142);
nand U2247 (N_2247,N_2164,N_2155);
or U2248 (N_2248,N_2148,N_2187);
nand U2249 (N_2249,N_2123,N_2101);
and U2250 (N_2250,N_2190,N_2121);
and U2251 (N_2251,N_2106,N_2134);
and U2252 (N_2252,N_2146,N_2112);
nand U2253 (N_2253,N_2110,N_2145);
nor U2254 (N_2254,N_2122,N_2175);
or U2255 (N_2255,N_2158,N_2167);
or U2256 (N_2256,N_2159,N_2133);
and U2257 (N_2257,N_2167,N_2138);
or U2258 (N_2258,N_2116,N_2193);
or U2259 (N_2259,N_2112,N_2158);
nor U2260 (N_2260,N_2121,N_2131);
nand U2261 (N_2261,N_2187,N_2144);
nor U2262 (N_2262,N_2108,N_2159);
or U2263 (N_2263,N_2141,N_2186);
and U2264 (N_2264,N_2172,N_2106);
nand U2265 (N_2265,N_2188,N_2174);
nor U2266 (N_2266,N_2161,N_2102);
and U2267 (N_2267,N_2107,N_2104);
nand U2268 (N_2268,N_2107,N_2135);
or U2269 (N_2269,N_2191,N_2159);
and U2270 (N_2270,N_2104,N_2161);
and U2271 (N_2271,N_2138,N_2127);
or U2272 (N_2272,N_2176,N_2194);
nand U2273 (N_2273,N_2127,N_2192);
and U2274 (N_2274,N_2167,N_2169);
or U2275 (N_2275,N_2187,N_2126);
or U2276 (N_2276,N_2169,N_2177);
nand U2277 (N_2277,N_2127,N_2137);
or U2278 (N_2278,N_2121,N_2106);
or U2279 (N_2279,N_2182,N_2140);
and U2280 (N_2280,N_2123,N_2180);
and U2281 (N_2281,N_2166,N_2162);
or U2282 (N_2282,N_2164,N_2129);
nand U2283 (N_2283,N_2106,N_2117);
nor U2284 (N_2284,N_2182,N_2136);
or U2285 (N_2285,N_2125,N_2175);
nand U2286 (N_2286,N_2124,N_2126);
or U2287 (N_2287,N_2149,N_2169);
nand U2288 (N_2288,N_2192,N_2159);
xnor U2289 (N_2289,N_2169,N_2161);
nor U2290 (N_2290,N_2141,N_2172);
or U2291 (N_2291,N_2130,N_2190);
or U2292 (N_2292,N_2104,N_2133);
nor U2293 (N_2293,N_2121,N_2132);
xor U2294 (N_2294,N_2161,N_2145);
or U2295 (N_2295,N_2153,N_2124);
and U2296 (N_2296,N_2186,N_2169);
nand U2297 (N_2297,N_2152,N_2160);
and U2298 (N_2298,N_2150,N_2103);
nand U2299 (N_2299,N_2173,N_2118);
or U2300 (N_2300,N_2212,N_2232);
or U2301 (N_2301,N_2256,N_2294);
or U2302 (N_2302,N_2268,N_2266);
nand U2303 (N_2303,N_2259,N_2226);
nand U2304 (N_2304,N_2201,N_2238);
nor U2305 (N_2305,N_2261,N_2264);
nor U2306 (N_2306,N_2280,N_2246);
and U2307 (N_2307,N_2253,N_2247);
nand U2308 (N_2308,N_2205,N_2220);
or U2309 (N_2309,N_2230,N_2270);
or U2310 (N_2310,N_2243,N_2263);
nand U2311 (N_2311,N_2245,N_2295);
nor U2312 (N_2312,N_2221,N_2224);
nand U2313 (N_2313,N_2296,N_2202);
and U2314 (N_2314,N_2288,N_2214);
nand U2315 (N_2315,N_2291,N_2275);
nor U2316 (N_2316,N_2219,N_2262);
nor U2317 (N_2317,N_2211,N_2251);
nand U2318 (N_2318,N_2257,N_2223);
and U2319 (N_2319,N_2290,N_2276);
nand U2320 (N_2320,N_2279,N_2241);
nor U2321 (N_2321,N_2273,N_2283);
nand U2322 (N_2322,N_2234,N_2236);
or U2323 (N_2323,N_2250,N_2209);
nand U2324 (N_2324,N_2200,N_2289);
nand U2325 (N_2325,N_2225,N_2227);
nand U2326 (N_2326,N_2204,N_2240);
or U2327 (N_2327,N_2286,N_2254);
nand U2328 (N_2328,N_2218,N_2207);
nand U2329 (N_2329,N_2269,N_2287);
nor U2330 (N_2330,N_2206,N_2239);
and U2331 (N_2331,N_2281,N_2237);
and U2332 (N_2332,N_2213,N_2272);
nor U2333 (N_2333,N_2252,N_2267);
nand U2334 (N_2334,N_2274,N_2248);
nand U2335 (N_2335,N_2297,N_2292);
or U2336 (N_2336,N_2210,N_2265);
nand U2337 (N_2337,N_2258,N_2242);
or U2338 (N_2338,N_2233,N_2217);
nor U2339 (N_2339,N_2215,N_2284);
and U2340 (N_2340,N_2293,N_2278);
and U2341 (N_2341,N_2222,N_2299);
and U2342 (N_2342,N_2228,N_2216);
or U2343 (N_2343,N_2244,N_2208);
or U2344 (N_2344,N_2277,N_2235);
and U2345 (N_2345,N_2229,N_2285);
and U2346 (N_2346,N_2298,N_2231);
and U2347 (N_2347,N_2203,N_2260);
and U2348 (N_2348,N_2271,N_2249);
and U2349 (N_2349,N_2255,N_2282);
and U2350 (N_2350,N_2216,N_2217);
nor U2351 (N_2351,N_2290,N_2269);
or U2352 (N_2352,N_2236,N_2208);
or U2353 (N_2353,N_2240,N_2200);
nand U2354 (N_2354,N_2272,N_2203);
or U2355 (N_2355,N_2223,N_2274);
nand U2356 (N_2356,N_2208,N_2299);
nor U2357 (N_2357,N_2275,N_2273);
nand U2358 (N_2358,N_2278,N_2205);
nor U2359 (N_2359,N_2226,N_2251);
and U2360 (N_2360,N_2250,N_2223);
and U2361 (N_2361,N_2214,N_2234);
and U2362 (N_2362,N_2262,N_2275);
xnor U2363 (N_2363,N_2254,N_2260);
and U2364 (N_2364,N_2267,N_2200);
and U2365 (N_2365,N_2263,N_2235);
nand U2366 (N_2366,N_2225,N_2261);
and U2367 (N_2367,N_2255,N_2209);
or U2368 (N_2368,N_2245,N_2277);
or U2369 (N_2369,N_2293,N_2220);
nor U2370 (N_2370,N_2236,N_2225);
nand U2371 (N_2371,N_2235,N_2210);
and U2372 (N_2372,N_2266,N_2217);
or U2373 (N_2373,N_2249,N_2201);
nand U2374 (N_2374,N_2242,N_2237);
and U2375 (N_2375,N_2293,N_2204);
nand U2376 (N_2376,N_2298,N_2294);
nor U2377 (N_2377,N_2275,N_2244);
and U2378 (N_2378,N_2292,N_2268);
nand U2379 (N_2379,N_2204,N_2211);
and U2380 (N_2380,N_2224,N_2279);
and U2381 (N_2381,N_2289,N_2213);
and U2382 (N_2382,N_2212,N_2229);
nand U2383 (N_2383,N_2258,N_2215);
or U2384 (N_2384,N_2290,N_2257);
or U2385 (N_2385,N_2287,N_2275);
and U2386 (N_2386,N_2259,N_2215);
and U2387 (N_2387,N_2223,N_2211);
or U2388 (N_2388,N_2237,N_2246);
or U2389 (N_2389,N_2239,N_2211);
and U2390 (N_2390,N_2209,N_2251);
nor U2391 (N_2391,N_2231,N_2208);
nor U2392 (N_2392,N_2226,N_2254);
nor U2393 (N_2393,N_2250,N_2274);
nand U2394 (N_2394,N_2233,N_2213);
or U2395 (N_2395,N_2243,N_2262);
or U2396 (N_2396,N_2291,N_2281);
or U2397 (N_2397,N_2271,N_2226);
and U2398 (N_2398,N_2296,N_2281);
and U2399 (N_2399,N_2258,N_2273);
nor U2400 (N_2400,N_2392,N_2378);
or U2401 (N_2401,N_2322,N_2374);
and U2402 (N_2402,N_2376,N_2341);
nor U2403 (N_2403,N_2377,N_2333);
or U2404 (N_2404,N_2357,N_2344);
or U2405 (N_2405,N_2343,N_2310);
or U2406 (N_2406,N_2360,N_2300);
or U2407 (N_2407,N_2345,N_2379);
and U2408 (N_2408,N_2354,N_2361);
or U2409 (N_2409,N_2349,N_2397);
nor U2410 (N_2410,N_2308,N_2353);
nand U2411 (N_2411,N_2323,N_2355);
nor U2412 (N_2412,N_2318,N_2380);
nand U2413 (N_2413,N_2363,N_2301);
nor U2414 (N_2414,N_2321,N_2342);
nor U2415 (N_2415,N_2368,N_2309);
or U2416 (N_2416,N_2365,N_2399);
or U2417 (N_2417,N_2324,N_2387);
or U2418 (N_2418,N_2394,N_2366);
or U2419 (N_2419,N_2312,N_2351);
nor U2420 (N_2420,N_2375,N_2383);
or U2421 (N_2421,N_2390,N_2398);
nand U2422 (N_2422,N_2337,N_2339);
nor U2423 (N_2423,N_2381,N_2326);
and U2424 (N_2424,N_2370,N_2388);
and U2425 (N_2425,N_2325,N_2359);
nor U2426 (N_2426,N_2391,N_2327);
and U2427 (N_2427,N_2352,N_2348);
nor U2428 (N_2428,N_2317,N_2364);
nor U2429 (N_2429,N_2350,N_2320);
nor U2430 (N_2430,N_2393,N_2358);
or U2431 (N_2431,N_2386,N_2302);
nor U2432 (N_2432,N_2371,N_2304);
nor U2433 (N_2433,N_2347,N_2303);
nand U2434 (N_2434,N_2332,N_2331);
nand U2435 (N_2435,N_2311,N_2306);
nand U2436 (N_2436,N_2346,N_2396);
nor U2437 (N_2437,N_2395,N_2372);
and U2438 (N_2438,N_2329,N_2389);
nand U2439 (N_2439,N_2319,N_2334);
nor U2440 (N_2440,N_2307,N_2335);
nor U2441 (N_2441,N_2382,N_2367);
nand U2442 (N_2442,N_2330,N_2362);
or U2443 (N_2443,N_2373,N_2340);
nand U2444 (N_2444,N_2316,N_2369);
or U2445 (N_2445,N_2338,N_2336);
nor U2446 (N_2446,N_2315,N_2385);
nand U2447 (N_2447,N_2356,N_2384);
and U2448 (N_2448,N_2328,N_2313);
or U2449 (N_2449,N_2305,N_2314);
and U2450 (N_2450,N_2368,N_2316);
and U2451 (N_2451,N_2366,N_2304);
and U2452 (N_2452,N_2303,N_2300);
nand U2453 (N_2453,N_2328,N_2332);
nand U2454 (N_2454,N_2348,N_2347);
or U2455 (N_2455,N_2359,N_2342);
nor U2456 (N_2456,N_2384,N_2349);
or U2457 (N_2457,N_2304,N_2359);
nand U2458 (N_2458,N_2309,N_2353);
nor U2459 (N_2459,N_2371,N_2376);
and U2460 (N_2460,N_2360,N_2337);
or U2461 (N_2461,N_2311,N_2361);
nand U2462 (N_2462,N_2370,N_2313);
and U2463 (N_2463,N_2304,N_2310);
nand U2464 (N_2464,N_2398,N_2325);
nor U2465 (N_2465,N_2324,N_2337);
and U2466 (N_2466,N_2334,N_2323);
or U2467 (N_2467,N_2390,N_2366);
or U2468 (N_2468,N_2336,N_2386);
and U2469 (N_2469,N_2380,N_2342);
or U2470 (N_2470,N_2396,N_2386);
and U2471 (N_2471,N_2383,N_2356);
nand U2472 (N_2472,N_2314,N_2344);
nand U2473 (N_2473,N_2308,N_2318);
or U2474 (N_2474,N_2313,N_2377);
and U2475 (N_2475,N_2344,N_2316);
and U2476 (N_2476,N_2320,N_2300);
and U2477 (N_2477,N_2323,N_2351);
nand U2478 (N_2478,N_2386,N_2338);
and U2479 (N_2479,N_2379,N_2359);
or U2480 (N_2480,N_2370,N_2330);
and U2481 (N_2481,N_2380,N_2305);
and U2482 (N_2482,N_2359,N_2351);
nor U2483 (N_2483,N_2319,N_2347);
or U2484 (N_2484,N_2307,N_2338);
and U2485 (N_2485,N_2343,N_2389);
nor U2486 (N_2486,N_2329,N_2318);
or U2487 (N_2487,N_2323,N_2393);
and U2488 (N_2488,N_2309,N_2373);
nor U2489 (N_2489,N_2361,N_2345);
or U2490 (N_2490,N_2343,N_2316);
and U2491 (N_2491,N_2371,N_2358);
nand U2492 (N_2492,N_2370,N_2302);
nor U2493 (N_2493,N_2374,N_2383);
nand U2494 (N_2494,N_2309,N_2359);
and U2495 (N_2495,N_2338,N_2395);
and U2496 (N_2496,N_2386,N_2315);
nand U2497 (N_2497,N_2347,N_2386);
nor U2498 (N_2498,N_2338,N_2377);
nand U2499 (N_2499,N_2347,N_2370);
nor U2500 (N_2500,N_2472,N_2439);
nor U2501 (N_2501,N_2454,N_2414);
and U2502 (N_2502,N_2434,N_2445);
or U2503 (N_2503,N_2462,N_2478);
nor U2504 (N_2504,N_2461,N_2402);
and U2505 (N_2505,N_2448,N_2468);
nor U2506 (N_2506,N_2429,N_2486);
nor U2507 (N_2507,N_2431,N_2499);
nand U2508 (N_2508,N_2411,N_2442);
nor U2509 (N_2509,N_2443,N_2477);
nand U2510 (N_2510,N_2447,N_2441);
and U2511 (N_2511,N_2464,N_2457);
and U2512 (N_2512,N_2416,N_2459);
nor U2513 (N_2513,N_2415,N_2412);
nor U2514 (N_2514,N_2458,N_2489);
or U2515 (N_2515,N_2470,N_2422);
nand U2516 (N_2516,N_2466,N_2428);
nand U2517 (N_2517,N_2479,N_2409);
and U2518 (N_2518,N_2473,N_2433);
and U2519 (N_2519,N_2494,N_2435);
and U2520 (N_2520,N_2496,N_2419);
and U2521 (N_2521,N_2436,N_2423);
nand U2522 (N_2522,N_2401,N_2495);
and U2523 (N_2523,N_2476,N_2440);
and U2524 (N_2524,N_2417,N_2491);
nor U2525 (N_2525,N_2425,N_2484);
or U2526 (N_2526,N_2444,N_2403);
nand U2527 (N_2527,N_2421,N_2483);
or U2528 (N_2528,N_2485,N_2450);
nand U2529 (N_2529,N_2474,N_2426);
nor U2530 (N_2530,N_2427,N_2456);
and U2531 (N_2531,N_2407,N_2469);
nand U2532 (N_2532,N_2480,N_2475);
and U2533 (N_2533,N_2467,N_2452);
and U2534 (N_2534,N_2453,N_2424);
or U2535 (N_2535,N_2455,N_2482);
nand U2536 (N_2536,N_2490,N_2481);
or U2537 (N_2537,N_2446,N_2465);
xnor U2538 (N_2538,N_2438,N_2413);
nand U2539 (N_2539,N_2492,N_2460);
or U2540 (N_2540,N_2432,N_2471);
nand U2541 (N_2541,N_2410,N_2497);
nand U2542 (N_2542,N_2487,N_2408);
nand U2543 (N_2543,N_2405,N_2463);
or U2544 (N_2544,N_2404,N_2437);
or U2545 (N_2545,N_2488,N_2449);
or U2546 (N_2546,N_2498,N_2418);
nand U2547 (N_2547,N_2451,N_2430);
or U2548 (N_2548,N_2400,N_2493);
nand U2549 (N_2549,N_2420,N_2406);
nor U2550 (N_2550,N_2457,N_2488);
and U2551 (N_2551,N_2488,N_2471);
or U2552 (N_2552,N_2448,N_2481);
or U2553 (N_2553,N_2454,N_2480);
or U2554 (N_2554,N_2432,N_2437);
nor U2555 (N_2555,N_2478,N_2455);
nor U2556 (N_2556,N_2489,N_2428);
nor U2557 (N_2557,N_2494,N_2457);
nand U2558 (N_2558,N_2473,N_2440);
nand U2559 (N_2559,N_2417,N_2400);
or U2560 (N_2560,N_2448,N_2492);
nand U2561 (N_2561,N_2431,N_2470);
xnor U2562 (N_2562,N_2429,N_2493);
nor U2563 (N_2563,N_2479,N_2443);
nor U2564 (N_2564,N_2454,N_2412);
nand U2565 (N_2565,N_2411,N_2461);
and U2566 (N_2566,N_2464,N_2409);
nand U2567 (N_2567,N_2474,N_2461);
or U2568 (N_2568,N_2419,N_2485);
nor U2569 (N_2569,N_2421,N_2473);
or U2570 (N_2570,N_2452,N_2418);
and U2571 (N_2571,N_2495,N_2435);
nand U2572 (N_2572,N_2458,N_2488);
and U2573 (N_2573,N_2471,N_2439);
and U2574 (N_2574,N_2485,N_2413);
nor U2575 (N_2575,N_2459,N_2453);
and U2576 (N_2576,N_2420,N_2429);
nor U2577 (N_2577,N_2497,N_2442);
xor U2578 (N_2578,N_2441,N_2480);
or U2579 (N_2579,N_2452,N_2485);
or U2580 (N_2580,N_2418,N_2497);
and U2581 (N_2581,N_2478,N_2476);
nor U2582 (N_2582,N_2420,N_2480);
nor U2583 (N_2583,N_2480,N_2490);
nor U2584 (N_2584,N_2490,N_2468);
nor U2585 (N_2585,N_2493,N_2461);
or U2586 (N_2586,N_2443,N_2498);
nor U2587 (N_2587,N_2498,N_2452);
nand U2588 (N_2588,N_2474,N_2459);
nor U2589 (N_2589,N_2446,N_2497);
nor U2590 (N_2590,N_2429,N_2419);
and U2591 (N_2591,N_2456,N_2467);
nand U2592 (N_2592,N_2410,N_2413);
nor U2593 (N_2593,N_2422,N_2458);
and U2594 (N_2594,N_2421,N_2495);
nand U2595 (N_2595,N_2422,N_2473);
nor U2596 (N_2596,N_2439,N_2498);
nand U2597 (N_2597,N_2464,N_2496);
and U2598 (N_2598,N_2492,N_2402);
nor U2599 (N_2599,N_2416,N_2497);
nand U2600 (N_2600,N_2518,N_2532);
or U2601 (N_2601,N_2552,N_2500);
nor U2602 (N_2602,N_2501,N_2545);
and U2603 (N_2603,N_2569,N_2529);
nand U2604 (N_2604,N_2510,N_2502);
nand U2605 (N_2605,N_2548,N_2589);
xor U2606 (N_2606,N_2586,N_2533);
nand U2607 (N_2607,N_2575,N_2593);
or U2608 (N_2608,N_2584,N_2511);
and U2609 (N_2609,N_2530,N_2506);
nand U2610 (N_2610,N_2576,N_2559);
or U2611 (N_2611,N_2542,N_2509);
nand U2612 (N_2612,N_2526,N_2571);
or U2613 (N_2613,N_2582,N_2514);
nand U2614 (N_2614,N_2537,N_2570);
nor U2615 (N_2615,N_2590,N_2592);
nand U2616 (N_2616,N_2568,N_2583);
or U2617 (N_2617,N_2560,N_2587);
nand U2618 (N_2618,N_2579,N_2546);
or U2619 (N_2619,N_2540,N_2504);
and U2620 (N_2620,N_2562,N_2536);
or U2621 (N_2621,N_2512,N_2563);
nand U2622 (N_2622,N_2535,N_2519);
or U2623 (N_2623,N_2580,N_2564);
and U2624 (N_2624,N_2581,N_2596);
and U2625 (N_2625,N_2549,N_2517);
nor U2626 (N_2626,N_2566,N_2544);
or U2627 (N_2627,N_2524,N_2541);
and U2628 (N_2628,N_2567,N_2525);
or U2629 (N_2629,N_2573,N_2577);
and U2630 (N_2630,N_2527,N_2516);
nand U2631 (N_2631,N_2550,N_2534);
or U2632 (N_2632,N_2513,N_2505);
or U2633 (N_2633,N_2551,N_2520);
and U2634 (N_2634,N_2585,N_2578);
or U2635 (N_2635,N_2599,N_2554);
or U2636 (N_2636,N_2588,N_2558);
nor U2637 (N_2637,N_2556,N_2597);
nor U2638 (N_2638,N_2507,N_2557);
or U2639 (N_2639,N_2503,N_2528);
nor U2640 (N_2640,N_2591,N_2561);
nor U2641 (N_2641,N_2515,N_2508);
or U2642 (N_2642,N_2521,N_2553);
or U2643 (N_2643,N_2538,N_2594);
and U2644 (N_2644,N_2574,N_2595);
nand U2645 (N_2645,N_2522,N_2543);
and U2646 (N_2646,N_2539,N_2565);
or U2647 (N_2647,N_2555,N_2572);
and U2648 (N_2648,N_2523,N_2547);
and U2649 (N_2649,N_2598,N_2531);
and U2650 (N_2650,N_2543,N_2550);
nor U2651 (N_2651,N_2506,N_2591);
nor U2652 (N_2652,N_2584,N_2580);
or U2653 (N_2653,N_2581,N_2580);
nor U2654 (N_2654,N_2565,N_2572);
nand U2655 (N_2655,N_2527,N_2586);
nor U2656 (N_2656,N_2589,N_2519);
or U2657 (N_2657,N_2580,N_2576);
nand U2658 (N_2658,N_2598,N_2592);
nor U2659 (N_2659,N_2588,N_2526);
and U2660 (N_2660,N_2537,N_2553);
nor U2661 (N_2661,N_2519,N_2534);
or U2662 (N_2662,N_2525,N_2531);
nand U2663 (N_2663,N_2503,N_2591);
nor U2664 (N_2664,N_2525,N_2577);
and U2665 (N_2665,N_2529,N_2507);
or U2666 (N_2666,N_2514,N_2547);
nand U2667 (N_2667,N_2551,N_2534);
or U2668 (N_2668,N_2556,N_2557);
and U2669 (N_2669,N_2504,N_2579);
nor U2670 (N_2670,N_2551,N_2583);
nor U2671 (N_2671,N_2547,N_2548);
xor U2672 (N_2672,N_2550,N_2506);
nor U2673 (N_2673,N_2558,N_2513);
and U2674 (N_2674,N_2527,N_2535);
or U2675 (N_2675,N_2593,N_2569);
and U2676 (N_2676,N_2580,N_2502);
nand U2677 (N_2677,N_2528,N_2531);
or U2678 (N_2678,N_2578,N_2573);
or U2679 (N_2679,N_2559,N_2554);
nand U2680 (N_2680,N_2540,N_2503);
and U2681 (N_2681,N_2593,N_2541);
xor U2682 (N_2682,N_2510,N_2596);
or U2683 (N_2683,N_2502,N_2559);
nand U2684 (N_2684,N_2523,N_2565);
and U2685 (N_2685,N_2519,N_2525);
xor U2686 (N_2686,N_2576,N_2544);
or U2687 (N_2687,N_2556,N_2508);
or U2688 (N_2688,N_2596,N_2539);
nor U2689 (N_2689,N_2590,N_2594);
and U2690 (N_2690,N_2524,N_2509);
and U2691 (N_2691,N_2531,N_2597);
or U2692 (N_2692,N_2584,N_2558);
nor U2693 (N_2693,N_2558,N_2579);
nand U2694 (N_2694,N_2503,N_2593);
nor U2695 (N_2695,N_2510,N_2514);
nand U2696 (N_2696,N_2543,N_2535);
or U2697 (N_2697,N_2590,N_2569);
nor U2698 (N_2698,N_2528,N_2500);
nand U2699 (N_2699,N_2592,N_2556);
nor U2700 (N_2700,N_2660,N_2632);
and U2701 (N_2701,N_2656,N_2685);
or U2702 (N_2702,N_2678,N_2659);
and U2703 (N_2703,N_2679,N_2652);
nor U2704 (N_2704,N_2608,N_2615);
or U2705 (N_2705,N_2675,N_2609);
or U2706 (N_2706,N_2696,N_2694);
and U2707 (N_2707,N_2616,N_2617);
and U2708 (N_2708,N_2642,N_2649);
or U2709 (N_2709,N_2698,N_2670);
nor U2710 (N_2710,N_2640,N_2600);
nand U2711 (N_2711,N_2655,N_2637);
or U2712 (N_2712,N_2607,N_2663);
or U2713 (N_2713,N_2603,N_2690);
nand U2714 (N_2714,N_2613,N_2665);
or U2715 (N_2715,N_2699,N_2658);
nand U2716 (N_2716,N_2689,N_2628);
or U2717 (N_2717,N_2610,N_2676);
nor U2718 (N_2718,N_2684,N_2672);
and U2719 (N_2719,N_2662,N_2671);
nand U2720 (N_2720,N_2630,N_2614);
nand U2721 (N_2721,N_2666,N_2623);
nor U2722 (N_2722,N_2605,N_2629);
or U2723 (N_2723,N_2697,N_2622);
and U2724 (N_2724,N_2682,N_2668);
nand U2725 (N_2725,N_2626,N_2647);
or U2726 (N_2726,N_2669,N_2653);
and U2727 (N_2727,N_2606,N_2635);
nand U2728 (N_2728,N_2691,N_2654);
or U2729 (N_2729,N_2681,N_2618);
nand U2730 (N_2730,N_2636,N_2687);
or U2731 (N_2731,N_2643,N_2661);
and U2732 (N_2732,N_2619,N_2692);
nand U2733 (N_2733,N_2646,N_2695);
or U2734 (N_2734,N_2620,N_2601);
or U2735 (N_2735,N_2645,N_2602);
nor U2736 (N_2736,N_2651,N_2674);
nor U2737 (N_2737,N_2604,N_2611);
and U2738 (N_2738,N_2664,N_2624);
and U2739 (N_2739,N_2683,N_2641);
nand U2740 (N_2740,N_2650,N_2693);
nand U2741 (N_2741,N_2657,N_2680);
nand U2742 (N_2742,N_2634,N_2621);
and U2743 (N_2743,N_2667,N_2644);
nand U2744 (N_2744,N_2612,N_2638);
or U2745 (N_2745,N_2633,N_2631);
nand U2746 (N_2746,N_2673,N_2625);
and U2747 (N_2747,N_2677,N_2648);
nor U2748 (N_2748,N_2627,N_2639);
nand U2749 (N_2749,N_2686,N_2688);
nand U2750 (N_2750,N_2630,N_2641);
nor U2751 (N_2751,N_2650,N_2655);
and U2752 (N_2752,N_2607,N_2665);
and U2753 (N_2753,N_2661,N_2692);
nand U2754 (N_2754,N_2616,N_2676);
and U2755 (N_2755,N_2625,N_2669);
nand U2756 (N_2756,N_2685,N_2622);
nand U2757 (N_2757,N_2602,N_2692);
nor U2758 (N_2758,N_2654,N_2678);
nor U2759 (N_2759,N_2632,N_2691);
nor U2760 (N_2760,N_2600,N_2609);
and U2761 (N_2761,N_2636,N_2645);
nor U2762 (N_2762,N_2662,N_2663);
nor U2763 (N_2763,N_2604,N_2684);
or U2764 (N_2764,N_2620,N_2602);
xnor U2765 (N_2765,N_2678,N_2618);
or U2766 (N_2766,N_2667,N_2673);
or U2767 (N_2767,N_2689,N_2622);
nand U2768 (N_2768,N_2604,N_2638);
or U2769 (N_2769,N_2618,N_2677);
nand U2770 (N_2770,N_2680,N_2633);
and U2771 (N_2771,N_2678,N_2636);
and U2772 (N_2772,N_2657,N_2666);
nand U2773 (N_2773,N_2697,N_2647);
nand U2774 (N_2774,N_2670,N_2668);
nor U2775 (N_2775,N_2695,N_2696);
nand U2776 (N_2776,N_2653,N_2658);
nor U2777 (N_2777,N_2641,N_2661);
or U2778 (N_2778,N_2699,N_2628);
and U2779 (N_2779,N_2682,N_2699);
nor U2780 (N_2780,N_2625,N_2640);
and U2781 (N_2781,N_2604,N_2690);
or U2782 (N_2782,N_2670,N_2660);
or U2783 (N_2783,N_2654,N_2696);
and U2784 (N_2784,N_2618,N_2693);
and U2785 (N_2785,N_2615,N_2695);
nor U2786 (N_2786,N_2693,N_2619);
xnor U2787 (N_2787,N_2656,N_2687);
nand U2788 (N_2788,N_2637,N_2675);
or U2789 (N_2789,N_2644,N_2665);
or U2790 (N_2790,N_2651,N_2623);
or U2791 (N_2791,N_2657,N_2649);
nor U2792 (N_2792,N_2688,N_2612);
nand U2793 (N_2793,N_2690,N_2641);
or U2794 (N_2794,N_2622,N_2621);
nor U2795 (N_2795,N_2600,N_2670);
nor U2796 (N_2796,N_2603,N_2673);
nor U2797 (N_2797,N_2605,N_2600);
xor U2798 (N_2798,N_2628,N_2635);
and U2799 (N_2799,N_2629,N_2688);
or U2800 (N_2800,N_2797,N_2747);
or U2801 (N_2801,N_2735,N_2716);
or U2802 (N_2802,N_2705,N_2793);
or U2803 (N_2803,N_2768,N_2780);
nor U2804 (N_2804,N_2712,N_2790);
xnor U2805 (N_2805,N_2755,N_2704);
nand U2806 (N_2806,N_2794,N_2766);
nor U2807 (N_2807,N_2798,N_2758);
or U2808 (N_2808,N_2720,N_2752);
or U2809 (N_2809,N_2734,N_2719);
nand U2810 (N_2810,N_2772,N_2718);
nand U2811 (N_2811,N_2723,N_2717);
or U2812 (N_2812,N_2736,N_2726);
nor U2813 (N_2813,N_2799,N_2742);
nor U2814 (N_2814,N_2702,N_2754);
nor U2815 (N_2815,N_2740,N_2711);
nor U2816 (N_2816,N_2700,N_2792);
and U2817 (N_2817,N_2714,N_2779);
nor U2818 (N_2818,N_2741,N_2707);
nand U2819 (N_2819,N_2767,N_2761);
and U2820 (N_2820,N_2746,N_2743);
or U2821 (N_2821,N_2776,N_2773);
and U2822 (N_2822,N_2759,N_2784);
nand U2823 (N_2823,N_2733,N_2732);
and U2824 (N_2824,N_2788,N_2763);
nand U2825 (N_2825,N_2789,N_2728);
or U2826 (N_2826,N_2737,N_2727);
nand U2827 (N_2827,N_2715,N_2770);
xnor U2828 (N_2828,N_2762,N_2721);
or U2829 (N_2829,N_2709,N_2764);
or U2830 (N_2830,N_2749,N_2713);
nand U2831 (N_2831,N_2771,N_2774);
and U2832 (N_2832,N_2745,N_2708);
and U2833 (N_2833,N_2729,N_2781);
xnor U2834 (N_2834,N_2722,N_2751);
and U2835 (N_2835,N_2724,N_2730);
nand U2836 (N_2836,N_2765,N_2744);
or U2837 (N_2837,N_2756,N_2782);
and U2838 (N_2838,N_2731,N_2791);
nand U2839 (N_2839,N_2739,N_2701);
nor U2840 (N_2840,N_2785,N_2706);
and U2841 (N_2841,N_2786,N_2725);
nor U2842 (N_2842,N_2757,N_2777);
and U2843 (N_2843,N_2787,N_2795);
or U2844 (N_2844,N_2753,N_2738);
xor U2845 (N_2845,N_2710,N_2796);
nand U2846 (N_2846,N_2778,N_2783);
nand U2847 (N_2847,N_2775,N_2748);
or U2848 (N_2848,N_2750,N_2703);
and U2849 (N_2849,N_2769,N_2760);
and U2850 (N_2850,N_2774,N_2738);
nor U2851 (N_2851,N_2779,N_2737);
or U2852 (N_2852,N_2757,N_2701);
nor U2853 (N_2853,N_2741,N_2712);
and U2854 (N_2854,N_2701,N_2705);
or U2855 (N_2855,N_2717,N_2701);
or U2856 (N_2856,N_2753,N_2709);
or U2857 (N_2857,N_2730,N_2791);
or U2858 (N_2858,N_2745,N_2785);
xnor U2859 (N_2859,N_2797,N_2794);
nor U2860 (N_2860,N_2746,N_2757);
and U2861 (N_2861,N_2729,N_2790);
and U2862 (N_2862,N_2720,N_2704);
nor U2863 (N_2863,N_2761,N_2765);
nor U2864 (N_2864,N_2703,N_2712);
nand U2865 (N_2865,N_2737,N_2786);
and U2866 (N_2866,N_2702,N_2741);
nand U2867 (N_2867,N_2747,N_2781);
and U2868 (N_2868,N_2744,N_2719);
and U2869 (N_2869,N_2768,N_2748);
or U2870 (N_2870,N_2713,N_2758);
nand U2871 (N_2871,N_2770,N_2714);
or U2872 (N_2872,N_2799,N_2710);
or U2873 (N_2873,N_2736,N_2778);
and U2874 (N_2874,N_2780,N_2732);
and U2875 (N_2875,N_2754,N_2761);
and U2876 (N_2876,N_2743,N_2786);
nand U2877 (N_2877,N_2707,N_2737);
and U2878 (N_2878,N_2737,N_2793);
nor U2879 (N_2879,N_2789,N_2717);
and U2880 (N_2880,N_2704,N_2794);
nand U2881 (N_2881,N_2760,N_2734);
nand U2882 (N_2882,N_2745,N_2703);
nor U2883 (N_2883,N_2740,N_2779);
nand U2884 (N_2884,N_2754,N_2750);
nor U2885 (N_2885,N_2797,N_2767);
nor U2886 (N_2886,N_2771,N_2729);
and U2887 (N_2887,N_2700,N_2742);
nand U2888 (N_2888,N_2702,N_2747);
nor U2889 (N_2889,N_2770,N_2729);
nand U2890 (N_2890,N_2726,N_2789);
nor U2891 (N_2891,N_2752,N_2728);
or U2892 (N_2892,N_2734,N_2723);
or U2893 (N_2893,N_2774,N_2790);
or U2894 (N_2894,N_2755,N_2777);
nor U2895 (N_2895,N_2768,N_2725);
and U2896 (N_2896,N_2705,N_2768);
or U2897 (N_2897,N_2763,N_2747);
nor U2898 (N_2898,N_2706,N_2733);
or U2899 (N_2899,N_2793,N_2701);
and U2900 (N_2900,N_2812,N_2898);
or U2901 (N_2901,N_2813,N_2811);
nor U2902 (N_2902,N_2875,N_2891);
xor U2903 (N_2903,N_2870,N_2869);
nor U2904 (N_2904,N_2863,N_2885);
nand U2905 (N_2905,N_2852,N_2867);
nor U2906 (N_2906,N_2849,N_2805);
and U2907 (N_2907,N_2878,N_2833);
nor U2908 (N_2908,N_2837,N_2820);
and U2909 (N_2909,N_2816,N_2854);
or U2910 (N_2910,N_2889,N_2847);
nand U2911 (N_2911,N_2848,N_2858);
and U2912 (N_2912,N_2884,N_2894);
or U2913 (N_2913,N_2831,N_2832);
nand U2914 (N_2914,N_2808,N_2804);
and U2915 (N_2915,N_2895,N_2844);
or U2916 (N_2916,N_2819,N_2855);
and U2917 (N_2917,N_2810,N_2892);
and U2918 (N_2918,N_2842,N_2899);
nor U2919 (N_2919,N_2886,N_2834);
and U2920 (N_2920,N_2845,N_2872);
nor U2921 (N_2921,N_2871,N_2818);
nand U2922 (N_2922,N_2879,N_2853);
or U2923 (N_2923,N_2835,N_2802);
nor U2924 (N_2924,N_2807,N_2893);
nor U2925 (N_2925,N_2827,N_2876);
or U2926 (N_2926,N_2823,N_2846);
or U2927 (N_2927,N_2883,N_2896);
nor U2928 (N_2928,N_2887,N_2843);
or U2929 (N_2929,N_2838,N_2880);
or U2930 (N_2930,N_2866,N_2839);
nand U2931 (N_2931,N_2841,N_2800);
nor U2932 (N_2932,N_2860,N_2865);
and U2933 (N_2933,N_2817,N_2829);
or U2934 (N_2934,N_2877,N_2861);
nor U2935 (N_2935,N_2822,N_2851);
or U2936 (N_2936,N_2815,N_2801);
or U2937 (N_2937,N_2803,N_2830);
or U2938 (N_2938,N_2836,N_2862);
nor U2939 (N_2939,N_2859,N_2882);
and U2940 (N_2940,N_2824,N_2850);
or U2941 (N_2941,N_2857,N_2814);
and U2942 (N_2942,N_2888,N_2873);
nor U2943 (N_2943,N_2821,N_2826);
xor U2944 (N_2944,N_2897,N_2881);
or U2945 (N_2945,N_2856,N_2868);
or U2946 (N_2946,N_2864,N_2806);
and U2947 (N_2947,N_2809,N_2874);
and U2948 (N_2948,N_2840,N_2828);
or U2949 (N_2949,N_2825,N_2890);
xor U2950 (N_2950,N_2863,N_2803);
nand U2951 (N_2951,N_2835,N_2821);
or U2952 (N_2952,N_2819,N_2817);
or U2953 (N_2953,N_2854,N_2815);
or U2954 (N_2954,N_2837,N_2816);
and U2955 (N_2955,N_2837,N_2819);
nand U2956 (N_2956,N_2898,N_2804);
or U2957 (N_2957,N_2858,N_2836);
or U2958 (N_2958,N_2858,N_2829);
nor U2959 (N_2959,N_2822,N_2828);
nor U2960 (N_2960,N_2804,N_2825);
nor U2961 (N_2961,N_2800,N_2859);
and U2962 (N_2962,N_2814,N_2843);
nand U2963 (N_2963,N_2855,N_2803);
or U2964 (N_2964,N_2883,N_2866);
and U2965 (N_2965,N_2825,N_2866);
nand U2966 (N_2966,N_2833,N_2886);
or U2967 (N_2967,N_2820,N_2830);
nor U2968 (N_2968,N_2841,N_2850);
nand U2969 (N_2969,N_2874,N_2896);
or U2970 (N_2970,N_2831,N_2862);
nand U2971 (N_2971,N_2837,N_2862);
and U2972 (N_2972,N_2878,N_2870);
xnor U2973 (N_2973,N_2875,N_2884);
nand U2974 (N_2974,N_2832,N_2864);
nor U2975 (N_2975,N_2875,N_2866);
and U2976 (N_2976,N_2826,N_2853);
xor U2977 (N_2977,N_2822,N_2838);
and U2978 (N_2978,N_2882,N_2821);
nor U2979 (N_2979,N_2824,N_2813);
and U2980 (N_2980,N_2897,N_2818);
and U2981 (N_2981,N_2851,N_2831);
or U2982 (N_2982,N_2833,N_2876);
nand U2983 (N_2983,N_2870,N_2817);
nor U2984 (N_2984,N_2879,N_2841);
or U2985 (N_2985,N_2882,N_2869);
and U2986 (N_2986,N_2891,N_2834);
nand U2987 (N_2987,N_2847,N_2877);
nand U2988 (N_2988,N_2842,N_2840);
nand U2989 (N_2989,N_2872,N_2831);
nor U2990 (N_2990,N_2888,N_2858);
nor U2991 (N_2991,N_2896,N_2875);
nand U2992 (N_2992,N_2888,N_2863);
nor U2993 (N_2993,N_2826,N_2863);
and U2994 (N_2994,N_2827,N_2836);
nand U2995 (N_2995,N_2875,N_2897);
and U2996 (N_2996,N_2885,N_2883);
nand U2997 (N_2997,N_2832,N_2896);
or U2998 (N_2998,N_2841,N_2822);
nor U2999 (N_2999,N_2883,N_2864);
nor UO_0 (O_0,N_2922,N_2902);
and UO_1 (O_1,N_2969,N_2955);
and UO_2 (O_2,N_2923,N_2973);
nand UO_3 (O_3,N_2906,N_2943);
and UO_4 (O_4,N_2968,N_2915);
nor UO_5 (O_5,N_2987,N_2972);
nand UO_6 (O_6,N_2996,N_2925);
xnor UO_7 (O_7,N_2921,N_2970);
or UO_8 (O_8,N_2907,N_2942);
nor UO_9 (O_9,N_2956,N_2900);
nand UO_10 (O_10,N_2935,N_2909);
or UO_11 (O_11,N_2997,N_2947);
nand UO_12 (O_12,N_2971,N_2976);
nor UO_13 (O_13,N_2986,N_2991);
xnor UO_14 (O_14,N_2918,N_2951);
or UO_15 (O_15,N_2958,N_2941);
nand UO_16 (O_16,N_2908,N_2940);
nor UO_17 (O_17,N_2944,N_2964);
nor UO_18 (O_18,N_2981,N_2933);
or UO_19 (O_19,N_2985,N_2903);
or UO_20 (O_20,N_2967,N_2980);
or UO_21 (O_21,N_2989,N_2924);
and UO_22 (O_22,N_2928,N_2979);
nor UO_23 (O_23,N_2914,N_2901);
nand UO_24 (O_24,N_2919,N_2978);
or UO_25 (O_25,N_2912,N_2905);
and UO_26 (O_26,N_2988,N_2957);
nor UO_27 (O_27,N_2946,N_2965);
nor UO_28 (O_28,N_2916,N_2904);
or UO_29 (O_29,N_2984,N_2913);
or UO_30 (O_30,N_2939,N_2920);
and UO_31 (O_31,N_2961,N_2938);
nand UO_32 (O_32,N_2927,N_2992);
and UO_33 (O_33,N_2954,N_2995);
nor UO_34 (O_34,N_2999,N_2930);
nor UO_35 (O_35,N_2974,N_2994);
nand UO_36 (O_36,N_2993,N_2911);
nor UO_37 (O_37,N_2945,N_2948);
nor UO_38 (O_38,N_2960,N_2990);
or UO_39 (O_39,N_2931,N_2950);
and UO_40 (O_40,N_2917,N_2983);
and UO_41 (O_41,N_2936,N_2998);
nand UO_42 (O_42,N_2952,N_2975);
nor UO_43 (O_43,N_2959,N_2910);
nor UO_44 (O_44,N_2949,N_2926);
and UO_45 (O_45,N_2953,N_2966);
nor UO_46 (O_46,N_2982,N_2932);
nand UO_47 (O_47,N_2963,N_2929);
or UO_48 (O_48,N_2937,N_2962);
nand UO_49 (O_49,N_2934,N_2977);
nor UO_50 (O_50,N_2971,N_2902);
nor UO_51 (O_51,N_2985,N_2956);
nor UO_52 (O_52,N_2923,N_2976);
nor UO_53 (O_53,N_2970,N_2950);
nor UO_54 (O_54,N_2916,N_2918);
or UO_55 (O_55,N_2927,N_2976);
nor UO_56 (O_56,N_2914,N_2954);
and UO_57 (O_57,N_2920,N_2954);
and UO_58 (O_58,N_2961,N_2954);
nor UO_59 (O_59,N_2943,N_2977);
nor UO_60 (O_60,N_2912,N_2976);
and UO_61 (O_61,N_2989,N_2943);
nor UO_62 (O_62,N_2973,N_2927);
nor UO_63 (O_63,N_2957,N_2949);
and UO_64 (O_64,N_2913,N_2921);
nor UO_65 (O_65,N_2972,N_2996);
or UO_66 (O_66,N_2969,N_2945);
nand UO_67 (O_67,N_2940,N_2999);
and UO_68 (O_68,N_2903,N_2998);
and UO_69 (O_69,N_2918,N_2910);
nor UO_70 (O_70,N_2917,N_2913);
or UO_71 (O_71,N_2941,N_2961);
or UO_72 (O_72,N_2957,N_2964);
nor UO_73 (O_73,N_2950,N_2921);
and UO_74 (O_74,N_2996,N_2986);
nor UO_75 (O_75,N_2993,N_2954);
nand UO_76 (O_76,N_2981,N_2921);
nand UO_77 (O_77,N_2950,N_2949);
or UO_78 (O_78,N_2969,N_2978);
nor UO_79 (O_79,N_2932,N_2907);
nor UO_80 (O_80,N_2954,N_2916);
xnor UO_81 (O_81,N_2902,N_2901);
nand UO_82 (O_82,N_2902,N_2970);
or UO_83 (O_83,N_2932,N_2996);
and UO_84 (O_84,N_2933,N_2918);
and UO_85 (O_85,N_2949,N_2923);
or UO_86 (O_86,N_2976,N_2922);
and UO_87 (O_87,N_2972,N_2977);
and UO_88 (O_88,N_2917,N_2947);
and UO_89 (O_89,N_2976,N_2907);
or UO_90 (O_90,N_2910,N_2945);
or UO_91 (O_91,N_2950,N_2905);
or UO_92 (O_92,N_2996,N_2916);
or UO_93 (O_93,N_2974,N_2962);
or UO_94 (O_94,N_2928,N_2965);
nor UO_95 (O_95,N_2994,N_2969);
nor UO_96 (O_96,N_2903,N_2909);
nand UO_97 (O_97,N_2920,N_2936);
nor UO_98 (O_98,N_2915,N_2959);
nor UO_99 (O_99,N_2929,N_2906);
nor UO_100 (O_100,N_2959,N_2952);
xnor UO_101 (O_101,N_2994,N_2978);
or UO_102 (O_102,N_2950,N_2985);
nand UO_103 (O_103,N_2908,N_2928);
nand UO_104 (O_104,N_2976,N_2966);
nand UO_105 (O_105,N_2996,N_2934);
and UO_106 (O_106,N_2960,N_2933);
nand UO_107 (O_107,N_2918,N_2961);
nand UO_108 (O_108,N_2949,N_2903);
nand UO_109 (O_109,N_2904,N_2988);
or UO_110 (O_110,N_2907,N_2973);
and UO_111 (O_111,N_2909,N_2945);
or UO_112 (O_112,N_2959,N_2905);
nand UO_113 (O_113,N_2966,N_2930);
nand UO_114 (O_114,N_2915,N_2949);
and UO_115 (O_115,N_2931,N_2963);
nand UO_116 (O_116,N_2999,N_2978);
nor UO_117 (O_117,N_2909,N_2931);
nand UO_118 (O_118,N_2987,N_2986);
nor UO_119 (O_119,N_2905,N_2907);
nand UO_120 (O_120,N_2981,N_2916);
nand UO_121 (O_121,N_2922,N_2967);
or UO_122 (O_122,N_2918,N_2937);
or UO_123 (O_123,N_2909,N_2974);
nor UO_124 (O_124,N_2925,N_2989);
or UO_125 (O_125,N_2947,N_2960);
and UO_126 (O_126,N_2938,N_2982);
xor UO_127 (O_127,N_2919,N_2908);
nor UO_128 (O_128,N_2915,N_2952);
nor UO_129 (O_129,N_2981,N_2934);
nand UO_130 (O_130,N_2944,N_2935);
and UO_131 (O_131,N_2909,N_2991);
nand UO_132 (O_132,N_2953,N_2958);
nand UO_133 (O_133,N_2979,N_2929);
and UO_134 (O_134,N_2966,N_2948);
and UO_135 (O_135,N_2994,N_2909);
or UO_136 (O_136,N_2942,N_2973);
nor UO_137 (O_137,N_2947,N_2954);
or UO_138 (O_138,N_2950,N_2954);
nor UO_139 (O_139,N_2964,N_2946);
nor UO_140 (O_140,N_2911,N_2927);
nor UO_141 (O_141,N_2931,N_2927);
and UO_142 (O_142,N_2942,N_2944);
or UO_143 (O_143,N_2995,N_2944);
or UO_144 (O_144,N_2919,N_2999);
nor UO_145 (O_145,N_2908,N_2968);
and UO_146 (O_146,N_2917,N_2977);
xor UO_147 (O_147,N_2938,N_2949);
and UO_148 (O_148,N_2925,N_2921);
nand UO_149 (O_149,N_2985,N_2973);
or UO_150 (O_150,N_2955,N_2937);
nand UO_151 (O_151,N_2968,N_2921);
or UO_152 (O_152,N_2910,N_2967);
and UO_153 (O_153,N_2932,N_2912);
nand UO_154 (O_154,N_2903,N_2981);
nor UO_155 (O_155,N_2928,N_2938);
nand UO_156 (O_156,N_2955,N_2980);
and UO_157 (O_157,N_2955,N_2944);
and UO_158 (O_158,N_2968,N_2920);
or UO_159 (O_159,N_2970,N_2952);
nand UO_160 (O_160,N_2913,N_2939);
or UO_161 (O_161,N_2973,N_2902);
and UO_162 (O_162,N_2906,N_2988);
and UO_163 (O_163,N_2986,N_2974);
nor UO_164 (O_164,N_2958,N_2940);
nand UO_165 (O_165,N_2940,N_2934);
nor UO_166 (O_166,N_2983,N_2950);
nand UO_167 (O_167,N_2935,N_2925);
xnor UO_168 (O_168,N_2924,N_2946);
nor UO_169 (O_169,N_2954,N_2970);
nor UO_170 (O_170,N_2947,N_2940);
or UO_171 (O_171,N_2901,N_2920);
nor UO_172 (O_172,N_2947,N_2968);
and UO_173 (O_173,N_2950,N_2981);
and UO_174 (O_174,N_2929,N_2937);
nand UO_175 (O_175,N_2946,N_2987);
and UO_176 (O_176,N_2918,N_2956);
and UO_177 (O_177,N_2906,N_2919);
or UO_178 (O_178,N_2921,N_2931);
nand UO_179 (O_179,N_2944,N_2989);
nor UO_180 (O_180,N_2902,N_2984);
nor UO_181 (O_181,N_2987,N_2930);
nand UO_182 (O_182,N_2926,N_2961);
nor UO_183 (O_183,N_2949,N_2982);
or UO_184 (O_184,N_2942,N_2991);
and UO_185 (O_185,N_2922,N_2901);
and UO_186 (O_186,N_2958,N_2919);
and UO_187 (O_187,N_2959,N_2903);
or UO_188 (O_188,N_2967,N_2927);
nor UO_189 (O_189,N_2905,N_2970);
or UO_190 (O_190,N_2949,N_2947);
nor UO_191 (O_191,N_2920,N_2909);
and UO_192 (O_192,N_2905,N_2900);
nand UO_193 (O_193,N_2966,N_2969);
nand UO_194 (O_194,N_2972,N_2900);
nor UO_195 (O_195,N_2910,N_2921);
nor UO_196 (O_196,N_2915,N_2982);
xnor UO_197 (O_197,N_2948,N_2949);
and UO_198 (O_198,N_2900,N_2962);
nand UO_199 (O_199,N_2924,N_2999);
and UO_200 (O_200,N_2930,N_2995);
or UO_201 (O_201,N_2949,N_2979);
and UO_202 (O_202,N_2935,N_2988);
and UO_203 (O_203,N_2949,N_2997);
nor UO_204 (O_204,N_2948,N_2915);
or UO_205 (O_205,N_2919,N_2917);
nor UO_206 (O_206,N_2926,N_2916);
and UO_207 (O_207,N_2954,N_2933);
or UO_208 (O_208,N_2969,N_2905);
nand UO_209 (O_209,N_2982,N_2922);
nand UO_210 (O_210,N_2987,N_2961);
nor UO_211 (O_211,N_2945,N_2937);
nand UO_212 (O_212,N_2985,N_2992);
nand UO_213 (O_213,N_2927,N_2982);
nand UO_214 (O_214,N_2916,N_2936);
or UO_215 (O_215,N_2950,N_2922);
nand UO_216 (O_216,N_2954,N_2956);
nor UO_217 (O_217,N_2911,N_2953);
nor UO_218 (O_218,N_2998,N_2906);
and UO_219 (O_219,N_2990,N_2946);
nand UO_220 (O_220,N_2997,N_2918);
nor UO_221 (O_221,N_2936,N_2962);
or UO_222 (O_222,N_2968,N_2935);
and UO_223 (O_223,N_2927,N_2914);
and UO_224 (O_224,N_2915,N_2991);
and UO_225 (O_225,N_2973,N_2925);
nand UO_226 (O_226,N_2998,N_2992);
nor UO_227 (O_227,N_2926,N_2954);
or UO_228 (O_228,N_2962,N_2917);
or UO_229 (O_229,N_2947,N_2920);
nor UO_230 (O_230,N_2962,N_2934);
nor UO_231 (O_231,N_2927,N_2945);
and UO_232 (O_232,N_2906,N_2995);
nand UO_233 (O_233,N_2962,N_2999);
nor UO_234 (O_234,N_2946,N_2929);
nand UO_235 (O_235,N_2928,N_2994);
or UO_236 (O_236,N_2931,N_2969);
or UO_237 (O_237,N_2981,N_2974);
nand UO_238 (O_238,N_2947,N_2980);
nor UO_239 (O_239,N_2976,N_2937);
or UO_240 (O_240,N_2969,N_2967);
nor UO_241 (O_241,N_2954,N_2923);
and UO_242 (O_242,N_2951,N_2978);
nand UO_243 (O_243,N_2947,N_2902);
xor UO_244 (O_244,N_2927,N_2957);
xnor UO_245 (O_245,N_2942,N_2914);
nand UO_246 (O_246,N_2919,N_2925);
or UO_247 (O_247,N_2991,N_2950);
or UO_248 (O_248,N_2987,N_2980);
and UO_249 (O_249,N_2986,N_2970);
and UO_250 (O_250,N_2918,N_2964);
and UO_251 (O_251,N_2980,N_2964);
and UO_252 (O_252,N_2980,N_2942);
nand UO_253 (O_253,N_2928,N_2933);
nand UO_254 (O_254,N_2973,N_2901);
nor UO_255 (O_255,N_2965,N_2909);
and UO_256 (O_256,N_2946,N_2919);
or UO_257 (O_257,N_2905,N_2997);
and UO_258 (O_258,N_2918,N_2969);
nor UO_259 (O_259,N_2936,N_2953);
nand UO_260 (O_260,N_2935,N_2999);
or UO_261 (O_261,N_2977,N_2948);
nor UO_262 (O_262,N_2957,N_2995);
nand UO_263 (O_263,N_2992,N_2968);
nor UO_264 (O_264,N_2960,N_2995);
nor UO_265 (O_265,N_2947,N_2989);
or UO_266 (O_266,N_2993,N_2963);
and UO_267 (O_267,N_2906,N_2926);
xnor UO_268 (O_268,N_2962,N_2979);
nor UO_269 (O_269,N_2951,N_2944);
nand UO_270 (O_270,N_2951,N_2928);
and UO_271 (O_271,N_2941,N_2947);
xnor UO_272 (O_272,N_2906,N_2999);
or UO_273 (O_273,N_2928,N_2966);
nor UO_274 (O_274,N_2991,N_2925);
and UO_275 (O_275,N_2941,N_2935);
nor UO_276 (O_276,N_2996,N_2987);
nor UO_277 (O_277,N_2965,N_2910);
or UO_278 (O_278,N_2985,N_2942);
nor UO_279 (O_279,N_2949,N_2934);
nor UO_280 (O_280,N_2955,N_2994);
nand UO_281 (O_281,N_2970,N_2910);
and UO_282 (O_282,N_2952,N_2913);
and UO_283 (O_283,N_2919,N_2937);
or UO_284 (O_284,N_2901,N_2930);
nand UO_285 (O_285,N_2957,N_2971);
and UO_286 (O_286,N_2923,N_2979);
nand UO_287 (O_287,N_2916,N_2929);
nand UO_288 (O_288,N_2932,N_2976);
xnor UO_289 (O_289,N_2900,N_2954);
and UO_290 (O_290,N_2989,N_2993);
or UO_291 (O_291,N_2984,N_2948);
and UO_292 (O_292,N_2990,N_2941);
nor UO_293 (O_293,N_2928,N_2921);
or UO_294 (O_294,N_2924,N_2986);
or UO_295 (O_295,N_2937,N_2901);
or UO_296 (O_296,N_2970,N_2944);
nor UO_297 (O_297,N_2958,N_2990);
xor UO_298 (O_298,N_2939,N_2958);
and UO_299 (O_299,N_2959,N_2918);
nand UO_300 (O_300,N_2985,N_2993);
nand UO_301 (O_301,N_2984,N_2985);
nand UO_302 (O_302,N_2974,N_2966);
nor UO_303 (O_303,N_2925,N_2923);
nor UO_304 (O_304,N_2900,N_2980);
nand UO_305 (O_305,N_2998,N_2957);
nor UO_306 (O_306,N_2900,N_2985);
nor UO_307 (O_307,N_2983,N_2968);
or UO_308 (O_308,N_2964,N_2911);
and UO_309 (O_309,N_2988,N_2932);
nor UO_310 (O_310,N_2961,N_2969);
and UO_311 (O_311,N_2900,N_2922);
nand UO_312 (O_312,N_2900,N_2941);
or UO_313 (O_313,N_2965,N_2900);
nand UO_314 (O_314,N_2954,N_2907);
nand UO_315 (O_315,N_2917,N_2999);
and UO_316 (O_316,N_2901,N_2961);
nor UO_317 (O_317,N_2932,N_2951);
nor UO_318 (O_318,N_2931,N_2936);
or UO_319 (O_319,N_2934,N_2911);
xor UO_320 (O_320,N_2964,N_2902);
nor UO_321 (O_321,N_2947,N_2994);
and UO_322 (O_322,N_2968,N_2999);
nor UO_323 (O_323,N_2970,N_2919);
and UO_324 (O_324,N_2984,N_2971);
xor UO_325 (O_325,N_2987,N_2922);
nor UO_326 (O_326,N_2903,N_2984);
and UO_327 (O_327,N_2939,N_2964);
nand UO_328 (O_328,N_2970,N_2907);
or UO_329 (O_329,N_2959,N_2964);
and UO_330 (O_330,N_2987,N_2982);
and UO_331 (O_331,N_2978,N_2985);
nand UO_332 (O_332,N_2988,N_2976);
or UO_333 (O_333,N_2925,N_2909);
and UO_334 (O_334,N_2955,N_2961);
nor UO_335 (O_335,N_2991,N_2911);
and UO_336 (O_336,N_2994,N_2933);
or UO_337 (O_337,N_2994,N_2936);
and UO_338 (O_338,N_2953,N_2962);
nor UO_339 (O_339,N_2952,N_2960);
and UO_340 (O_340,N_2981,N_2923);
nand UO_341 (O_341,N_2913,N_2979);
or UO_342 (O_342,N_2958,N_2909);
or UO_343 (O_343,N_2941,N_2923);
nand UO_344 (O_344,N_2960,N_2905);
nor UO_345 (O_345,N_2922,N_2971);
and UO_346 (O_346,N_2996,N_2983);
nand UO_347 (O_347,N_2914,N_2908);
nor UO_348 (O_348,N_2917,N_2993);
and UO_349 (O_349,N_2950,N_2935);
or UO_350 (O_350,N_2998,N_2943);
nand UO_351 (O_351,N_2985,N_2911);
nand UO_352 (O_352,N_2948,N_2989);
and UO_353 (O_353,N_2964,N_2910);
nor UO_354 (O_354,N_2984,N_2962);
nand UO_355 (O_355,N_2956,N_2961);
nand UO_356 (O_356,N_2952,N_2994);
and UO_357 (O_357,N_2937,N_2920);
and UO_358 (O_358,N_2956,N_2971);
and UO_359 (O_359,N_2900,N_2943);
nor UO_360 (O_360,N_2992,N_2977);
xor UO_361 (O_361,N_2947,N_2930);
or UO_362 (O_362,N_2942,N_2994);
and UO_363 (O_363,N_2949,N_2995);
or UO_364 (O_364,N_2986,N_2969);
and UO_365 (O_365,N_2949,N_2980);
and UO_366 (O_366,N_2971,N_2926);
nand UO_367 (O_367,N_2923,N_2965);
and UO_368 (O_368,N_2936,N_2991);
and UO_369 (O_369,N_2967,N_2908);
nor UO_370 (O_370,N_2950,N_2986);
nand UO_371 (O_371,N_2927,N_2919);
nor UO_372 (O_372,N_2959,N_2998);
or UO_373 (O_373,N_2923,N_2953);
nand UO_374 (O_374,N_2952,N_2962);
nand UO_375 (O_375,N_2978,N_2974);
or UO_376 (O_376,N_2974,N_2998);
or UO_377 (O_377,N_2909,N_2995);
nor UO_378 (O_378,N_2951,N_2980);
nor UO_379 (O_379,N_2977,N_2924);
or UO_380 (O_380,N_2990,N_2949);
nor UO_381 (O_381,N_2912,N_2936);
nor UO_382 (O_382,N_2924,N_2966);
nor UO_383 (O_383,N_2912,N_2975);
or UO_384 (O_384,N_2953,N_2921);
or UO_385 (O_385,N_2987,N_2948);
nor UO_386 (O_386,N_2995,N_2970);
or UO_387 (O_387,N_2915,N_2986);
nor UO_388 (O_388,N_2979,N_2924);
nand UO_389 (O_389,N_2901,N_2960);
nand UO_390 (O_390,N_2935,N_2939);
or UO_391 (O_391,N_2946,N_2962);
nor UO_392 (O_392,N_2923,N_2915);
nor UO_393 (O_393,N_2996,N_2922);
nand UO_394 (O_394,N_2996,N_2957);
or UO_395 (O_395,N_2918,N_2962);
or UO_396 (O_396,N_2996,N_2994);
nor UO_397 (O_397,N_2928,N_2957);
nor UO_398 (O_398,N_2960,N_2916);
nand UO_399 (O_399,N_2961,N_2914);
nor UO_400 (O_400,N_2947,N_2961);
nor UO_401 (O_401,N_2923,N_2906);
or UO_402 (O_402,N_2923,N_2918);
nand UO_403 (O_403,N_2935,N_2990);
and UO_404 (O_404,N_2905,N_2957);
or UO_405 (O_405,N_2974,N_2968);
nor UO_406 (O_406,N_2912,N_2943);
nand UO_407 (O_407,N_2932,N_2980);
nor UO_408 (O_408,N_2984,N_2919);
nor UO_409 (O_409,N_2949,N_2967);
nand UO_410 (O_410,N_2963,N_2986);
nand UO_411 (O_411,N_2965,N_2968);
or UO_412 (O_412,N_2916,N_2956);
or UO_413 (O_413,N_2968,N_2957);
or UO_414 (O_414,N_2984,N_2909);
or UO_415 (O_415,N_2908,N_2952);
nand UO_416 (O_416,N_2984,N_2951);
or UO_417 (O_417,N_2944,N_2926);
or UO_418 (O_418,N_2967,N_2919);
or UO_419 (O_419,N_2989,N_2946);
nand UO_420 (O_420,N_2990,N_2910);
nand UO_421 (O_421,N_2991,N_2999);
and UO_422 (O_422,N_2901,N_2919);
or UO_423 (O_423,N_2913,N_2968);
nor UO_424 (O_424,N_2913,N_2938);
and UO_425 (O_425,N_2917,N_2936);
and UO_426 (O_426,N_2905,N_2990);
nor UO_427 (O_427,N_2940,N_2971);
and UO_428 (O_428,N_2967,N_2951);
nand UO_429 (O_429,N_2917,N_2910);
and UO_430 (O_430,N_2925,N_2978);
nand UO_431 (O_431,N_2904,N_2914);
nand UO_432 (O_432,N_2928,N_2942);
nor UO_433 (O_433,N_2972,N_2921);
nand UO_434 (O_434,N_2993,N_2936);
and UO_435 (O_435,N_2976,N_2990);
nand UO_436 (O_436,N_2941,N_2970);
and UO_437 (O_437,N_2984,N_2994);
or UO_438 (O_438,N_2918,N_2935);
or UO_439 (O_439,N_2904,N_2975);
and UO_440 (O_440,N_2975,N_2954);
nand UO_441 (O_441,N_2963,N_2915);
nand UO_442 (O_442,N_2992,N_2996);
or UO_443 (O_443,N_2946,N_2971);
nor UO_444 (O_444,N_2913,N_2957);
xor UO_445 (O_445,N_2934,N_2989);
nor UO_446 (O_446,N_2946,N_2953);
and UO_447 (O_447,N_2982,N_2917);
nor UO_448 (O_448,N_2955,N_2995);
or UO_449 (O_449,N_2949,N_2931);
nand UO_450 (O_450,N_2980,N_2959);
and UO_451 (O_451,N_2981,N_2905);
or UO_452 (O_452,N_2926,N_2922);
or UO_453 (O_453,N_2955,N_2930);
nor UO_454 (O_454,N_2930,N_2905);
and UO_455 (O_455,N_2912,N_2921);
nor UO_456 (O_456,N_2966,N_2949);
nor UO_457 (O_457,N_2992,N_2974);
or UO_458 (O_458,N_2983,N_2930);
or UO_459 (O_459,N_2957,N_2900);
or UO_460 (O_460,N_2912,N_2950);
or UO_461 (O_461,N_2955,N_2922);
or UO_462 (O_462,N_2992,N_2931);
nor UO_463 (O_463,N_2914,N_2913);
nand UO_464 (O_464,N_2957,N_2967);
nand UO_465 (O_465,N_2962,N_2977);
and UO_466 (O_466,N_2957,N_2942);
nand UO_467 (O_467,N_2962,N_2994);
and UO_468 (O_468,N_2974,N_2975);
nand UO_469 (O_469,N_2975,N_2934);
and UO_470 (O_470,N_2933,N_2937);
or UO_471 (O_471,N_2917,N_2948);
and UO_472 (O_472,N_2961,N_2948);
and UO_473 (O_473,N_2930,N_2924);
and UO_474 (O_474,N_2961,N_2950);
or UO_475 (O_475,N_2952,N_2979);
nor UO_476 (O_476,N_2956,N_2986);
nor UO_477 (O_477,N_2985,N_2907);
nor UO_478 (O_478,N_2951,N_2931);
or UO_479 (O_479,N_2994,N_2971);
nor UO_480 (O_480,N_2910,N_2937);
and UO_481 (O_481,N_2971,N_2981);
and UO_482 (O_482,N_2956,N_2925);
nor UO_483 (O_483,N_2980,N_2990);
or UO_484 (O_484,N_2958,N_2916);
nand UO_485 (O_485,N_2951,N_2946);
or UO_486 (O_486,N_2969,N_2953);
or UO_487 (O_487,N_2902,N_2950);
nand UO_488 (O_488,N_2909,N_2908);
and UO_489 (O_489,N_2987,N_2958);
nand UO_490 (O_490,N_2943,N_2969);
nand UO_491 (O_491,N_2949,N_2946);
and UO_492 (O_492,N_2907,N_2911);
nor UO_493 (O_493,N_2989,N_2938);
or UO_494 (O_494,N_2963,N_2930);
or UO_495 (O_495,N_2988,N_2901);
or UO_496 (O_496,N_2948,N_2982);
nor UO_497 (O_497,N_2909,N_2987);
nand UO_498 (O_498,N_2992,N_2942);
nor UO_499 (O_499,N_2926,N_2986);
endmodule