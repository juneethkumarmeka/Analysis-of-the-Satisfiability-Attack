module basic_500_3000_500_60_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_256,In_261);
and U1 (N_1,In_231,In_433);
and U2 (N_2,In_195,In_72);
or U3 (N_3,In_307,In_148);
nor U4 (N_4,In_157,In_220);
and U5 (N_5,In_131,In_362);
nor U6 (N_6,In_271,In_194);
xnor U7 (N_7,In_292,In_424);
or U8 (N_8,In_116,In_203);
xnor U9 (N_9,In_467,In_278);
xor U10 (N_10,In_263,In_155);
and U11 (N_11,In_366,In_139);
nand U12 (N_12,In_339,In_373);
and U13 (N_13,In_249,In_490);
nor U14 (N_14,In_451,In_100);
xor U15 (N_15,In_452,In_83);
xnor U16 (N_16,In_13,In_64);
and U17 (N_17,In_213,In_172);
xor U18 (N_18,In_458,In_412);
xnor U19 (N_19,In_180,In_161);
nand U20 (N_20,In_472,In_422);
or U21 (N_21,In_30,In_327);
nand U22 (N_22,In_334,In_250);
or U23 (N_23,In_393,In_143);
and U24 (N_24,In_269,In_304);
xnor U25 (N_25,In_428,In_150);
nor U26 (N_26,In_262,In_471);
or U27 (N_27,In_380,In_237);
or U28 (N_28,In_162,In_49);
nor U29 (N_29,In_78,In_112);
or U30 (N_30,In_363,In_221);
nand U31 (N_31,In_496,In_431);
nor U32 (N_32,In_35,In_492);
and U33 (N_33,In_8,In_427);
nand U34 (N_34,In_477,In_192);
and U35 (N_35,In_236,In_300);
nor U36 (N_36,In_441,In_337);
xnor U37 (N_37,In_158,In_62);
nor U38 (N_38,In_429,In_163);
and U39 (N_39,In_29,In_365);
and U40 (N_40,In_214,In_371);
and U41 (N_41,In_449,In_342);
nand U42 (N_42,In_306,In_385);
nand U43 (N_43,In_298,In_246);
xor U44 (N_44,In_196,In_379);
nor U45 (N_45,In_343,In_270);
nor U46 (N_46,In_151,In_184);
and U47 (N_47,In_178,In_445);
xor U48 (N_48,In_129,In_400);
nor U49 (N_49,In_460,In_11);
xnor U50 (N_50,In_138,In_93);
nor U51 (N_51,In_386,In_448);
or U52 (N_52,In_197,In_160);
nand U53 (N_53,In_126,In_113);
nor U54 (N_54,In_34,In_308);
nor U55 (N_55,In_411,In_22);
or U56 (N_56,In_4,In_344);
nor U57 (N_57,In_102,In_39);
and U58 (N_58,In_159,In_144);
nand U59 (N_59,In_57,In_101);
nand U60 (N_60,In_87,In_105);
and U61 (N_61,N_2,In_247);
nor U62 (N_62,In_127,In_484);
or U63 (N_63,In_368,In_47);
and U64 (N_64,In_210,In_275);
nand U65 (N_65,In_140,N_29);
or U66 (N_66,In_227,In_26);
or U67 (N_67,In_38,In_440);
and U68 (N_68,In_154,In_205);
and U69 (N_69,In_421,In_341);
nor U70 (N_70,In_128,N_15);
nand U71 (N_71,In_9,In_480);
and U72 (N_72,In_69,In_274);
nand U73 (N_73,In_335,N_4);
nor U74 (N_74,In_369,In_86);
nor U75 (N_75,In_175,In_240);
or U76 (N_76,In_245,N_20);
nand U77 (N_77,In_499,In_374);
and U78 (N_78,In_348,In_404);
and U79 (N_79,In_99,In_241);
nand U80 (N_80,In_137,In_316);
nand U81 (N_81,In_169,In_388);
nor U82 (N_82,N_34,In_328);
xnor U83 (N_83,In_212,N_43);
nand U84 (N_84,In_19,In_478);
nand U85 (N_85,In_253,In_491);
and U86 (N_86,In_21,In_119);
or U87 (N_87,In_457,In_437);
nor U88 (N_88,In_45,N_36);
nor U89 (N_89,In_375,In_358);
nand U90 (N_90,In_215,In_199);
nand U91 (N_91,N_49,In_426);
or U92 (N_92,In_482,N_27);
or U93 (N_93,In_265,In_284);
xor U94 (N_94,In_340,In_146);
xor U95 (N_95,N_30,In_164);
xor U96 (N_96,In_43,N_5);
xor U97 (N_97,In_419,In_51);
and U98 (N_98,In_326,In_408);
nand U99 (N_99,In_234,In_90);
and U100 (N_100,N_7,N_59);
and U101 (N_101,In_376,In_238);
or U102 (N_102,In_318,In_291);
or U103 (N_103,In_301,In_382);
and U104 (N_104,In_0,N_9);
or U105 (N_105,In_498,In_165);
xnor U106 (N_106,In_207,In_67);
nor U107 (N_107,N_95,In_225);
or U108 (N_108,In_266,In_222);
nand U109 (N_109,In_187,In_446);
and U110 (N_110,In_325,In_309);
nor U111 (N_111,In_314,In_461);
nor U112 (N_112,In_1,In_439);
nand U113 (N_113,In_27,N_45);
nor U114 (N_114,N_80,In_268);
nor U115 (N_115,In_71,In_420);
xnor U116 (N_116,In_356,In_346);
or U117 (N_117,In_475,N_98);
nor U118 (N_118,In_487,In_48);
and U119 (N_119,In_191,N_75);
and U120 (N_120,In_181,In_394);
nand U121 (N_121,In_493,N_11);
xnor U122 (N_122,In_398,In_149);
nand U123 (N_123,In_257,In_59);
and U124 (N_124,N_68,N_22);
nor U125 (N_125,In_211,In_75);
xor U126 (N_126,In_277,In_410);
and U127 (N_127,In_405,In_202);
nor U128 (N_128,In_103,In_179);
nand U129 (N_129,In_289,In_264);
nand U130 (N_130,In_470,In_111);
and U131 (N_131,N_3,In_488);
nor U132 (N_132,In_281,In_377);
or U133 (N_133,N_12,In_37);
or U134 (N_134,In_198,In_305);
xnor U135 (N_135,In_248,In_6);
xor U136 (N_136,N_99,In_185);
and U137 (N_137,In_473,N_82);
and U138 (N_138,In_106,In_174);
and U139 (N_139,N_50,In_186);
xor U140 (N_140,In_392,In_434);
xor U141 (N_141,In_466,In_364);
and U142 (N_142,In_82,In_41);
nor U143 (N_143,N_57,N_19);
or U144 (N_144,In_267,In_120);
and U145 (N_145,In_414,In_217);
nor U146 (N_146,In_136,In_367);
and U147 (N_147,In_331,N_26);
nand U148 (N_148,In_481,In_468);
nand U149 (N_149,In_476,In_177);
and U150 (N_150,N_101,In_390);
xnor U151 (N_151,N_135,N_114);
nor U152 (N_152,In_183,N_91);
xor U153 (N_153,In_351,In_299);
or U154 (N_154,N_48,N_23);
and U155 (N_155,N_119,In_436);
xor U156 (N_156,N_40,N_24);
nor U157 (N_157,N_88,In_74);
or U158 (N_158,N_13,N_25);
or U159 (N_159,N_78,In_223);
nor U160 (N_160,In_14,In_228);
nand U161 (N_161,In_360,N_90);
and U162 (N_162,In_276,In_125);
nand U163 (N_163,N_16,In_323);
nor U164 (N_164,In_85,In_12);
and U165 (N_165,N_14,In_219);
and U166 (N_166,N_111,N_134);
and U167 (N_167,In_430,In_81);
and U168 (N_168,N_81,N_118);
xnor U169 (N_169,N_56,N_85);
and U170 (N_170,In_396,In_297);
nor U171 (N_171,N_117,In_399);
or U172 (N_172,In_332,In_55);
nand U173 (N_173,N_28,In_409);
nor U174 (N_174,In_118,N_35);
nand U175 (N_175,In_167,N_54);
and U176 (N_176,N_62,In_285);
or U177 (N_177,In_173,In_235);
or U178 (N_178,N_108,In_313);
nor U179 (N_179,In_324,N_129);
nor U180 (N_180,In_329,In_312);
xnor U181 (N_181,N_120,In_333);
nor U182 (N_182,In_255,N_32);
or U183 (N_183,In_447,In_242);
or U184 (N_184,In_287,In_84);
or U185 (N_185,In_350,N_100);
nor U186 (N_186,In_200,In_479);
nor U187 (N_187,In_2,N_121);
and U188 (N_188,In_432,In_370);
nor U189 (N_189,In_53,In_208);
xor U190 (N_190,In_355,N_93);
or U191 (N_191,In_311,In_273);
nor U192 (N_192,In_24,N_70);
and U193 (N_193,N_125,N_1);
and U194 (N_194,In_190,N_38);
nor U195 (N_195,In_107,N_113);
or U196 (N_196,In_232,In_189);
nor U197 (N_197,N_77,In_209);
or U198 (N_198,In_387,N_104);
or U199 (N_199,In_3,N_71);
or U200 (N_200,In_95,In_5);
nand U201 (N_201,N_73,In_359);
or U202 (N_202,N_164,In_293);
nor U203 (N_203,In_224,In_92);
and U204 (N_204,N_74,In_474);
or U205 (N_205,N_60,In_455);
or U206 (N_206,N_123,N_102);
and U207 (N_207,N_126,N_122);
or U208 (N_208,N_83,In_459);
or U209 (N_209,N_160,In_52);
and U210 (N_210,In_361,N_146);
xor U211 (N_211,N_159,N_109);
and U212 (N_212,N_31,N_138);
nor U213 (N_213,N_180,In_96);
and U214 (N_214,N_42,N_53);
and U215 (N_215,In_402,In_384);
xnor U216 (N_216,In_54,In_330);
xnor U217 (N_217,In_483,In_413);
nand U218 (N_218,N_103,In_94);
and U219 (N_219,In_117,N_167);
and U220 (N_220,In_28,N_105);
nor U221 (N_221,N_145,N_67);
xnor U222 (N_222,In_115,N_192);
and U223 (N_223,In_68,N_21);
nand U224 (N_224,N_162,N_131);
nand U225 (N_225,N_174,In_166);
nand U226 (N_226,In_453,In_206);
nor U227 (N_227,In_295,In_442);
or U228 (N_228,N_175,In_17);
xnor U229 (N_229,N_106,N_140);
nand U230 (N_230,In_438,In_283);
nor U231 (N_231,In_141,In_254);
xor U232 (N_232,In_66,N_84);
nor U233 (N_233,In_121,N_161);
nor U234 (N_234,In_272,In_454);
nor U235 (N_235,In_251,N_76);
and U236 (N_236,In_50,N_185);
and U237 (N_237,In_230,N_148);
nand U238 (N_238,In_495,In_288);
xnor U239 (N_239,In_114,N_0);
or U240 (N_240,N_187,In_303);
or U241 (N_241,In_243,In_176);
xor U242 (N_242,N_142,In_89);
xor U243 (N_243,N_156,N_136);
xor U244 (N_244,In_170,N_47);
nor U245 (N_245,N_197,In_389);
nor U246 (N_246,N_137,N_115);
nand U247 (N_247,In_109,In_23);
or U248 (N_248,N_94,In_486);
nand U249 (N_249,In_153,N_141);
nor U250 (N_250,N_249,N_63);
nand U251 (N_251,In_310,In_77);
nor U252 (N_252,N_188,N_237);
nor U253 (N_253,N_168,In_61);
xor U254 (N_254,N_149,N_176);
nor U255 (N_255,N_183,N_79);
and U256 (N_256,In_130,N_171);
and U257 (N_257,In_463,N_89);
or U258 (N_258,N_213,In_204);
nor U259 (N_259,N_173,In_401);
nand U260 (N_260,In_444,N_112);
or U261 (N_261,N_154,N_147);
nor U262 (N_262,In_20,N_232);
and U263 (N_263,In_44,In_42);
or U264 (N_264,In_406,In_435);
nand U265 (N_265,N_227,N_152);
or U266 (N_266,N_215,In_88);
nand U267 (N_267,N_17,N_235);
and U268 (N_268,N_178,In_145);
and U269 (N_269,In_104,In_110);
nand U270 (N_270,N_222,N_61);
nor U271 (N_271,N_127,N_204);
nand U272 (N_272,N_165,N_225);
or U273 (N_273,In_216,N_170);
nor U274 (N_274,N_214,In_58);
xor U275 (N_275,N_205,N_133);
and U276 (N_276,In_188,N_87);
and U277 (N_277,In_497,N_6);
or U278 (N_278,In_70,In_290);
and U279 (N_279,In_416,In_25);
xnor U280 (N_280,N_151,In_469);
or U281 (N_281,N_224,N_243);
xor U282 (N_282,N_233,N_210);
nand U283 (N_283,In_36,In_315);
xor U284 (N_284,N_244,N_206);
nand U285 (N_285,In_319,N_228);
nor U286 (N_286,In_201,In_32);
xnor U287 (N_287,In_134,In_10);
nor U288 (N_288,N_58,In_391);
xnor U289 (N_289,In_135,In_349);
nor U290 (N_290,N_37,N_92);
and U291 (N_291,In_279,N_211);
nor U292 (N_292,N_195,N_116);
xnor U293 (N_293,N_216,N_110);
and U294 (N_294,In_423,In_239);
xor U295 (N_295,N_209,N_169);
nor U296 (N_296,In_462,N_18);
xor U297 (N_297,In_18,In_296);
and U298 (N_298,N_96,In_372);
and U299 (N_299,N_97,In_40);
xnor U300 (N_300,In_79,N_287);
xnor U301 (N_301,In_46,In_258);
or U302 (N_302,N_229,In_415);
nand U303 (N_303,N_259,N_257);
and U304 (N_304,N_282,N_69);
nand U305 (N_305,N_207,In_353);
or U306 (N_306,N_271,N_295);
and U307 (N_307,N_181,N_179);
nor U308 (N_308,N_163,N_242);
xnor U309 (N_309,N_290,N_220);
nor U310 (N_310,N_184,In_259);
xnor U311 (N_311,In_168,N_52);
nor U312 (N_312,In_485,N_239);
or U313 (N_313,In_15,In_280);
or U314 (N_314,N_150,In_16);
nor U315 (N_315,In_417,N_212);
or U316 (N_316,N_128,N_202);
or U317 (N_317,N_297,N_238);
or U318 (N_318,N_107,In_494);
nor U319 (N_319,N_41,N_246);
or U320 (N_320,N_281,In_336);
and U321 (N_321,In_76,N_198);
xnor U322 (N_322,N_64,N_260);
xor U323 (N_323,N_124,N_286);
nand U324 (N_324,N_44,In_122);
or U325 (N_325,N_275,In_244);
and U326 (N_326,In_60,In_321);
or U327 (N_327,N_272,N_274);
and U328 (N_328,In_338,N_240);
nand U329 (N_329,N_157,In_133);
and U330 (N_330,In_123,N_226);
and U331 (N_331,N_270,N_294);
nand U332 (N_332,In_347,N_51);
xor U333 (N_333,N_39,N_189);
nand U334 (N_334,N_199,N_236);
nand U335 (N_335,N_155,N_218);
nor U336 (N_336,In_383,N_186);
xnor U337 (N_337,N_264,In_489);
xor U338 (N_338,N_241,N_279);
xor U339 (N_339,N_278,N_299);
xor U340 (N_340,In_7,In_142);
xor U341 (N_341,In_403,N_273);
xor U342 (N_342,N_230,N_182);
or U343 (N_343,In_418,In_56);
nand U344 (N_344,N_33,N_203);
and U345 (N_345,In_286,In_108);
or U346 (N_346,N_293,In_132);
or U347 (N_347,N_132,N_201);
nand U348 (N_348,N_130,N_285);
or U349 (N_349,N_248,N_266);
xor U350 (N_350,In_260,N_302);
xnor U351 (N_351,N_277,In_357);
nand U352 (N_352,In_352,N_314);
and U353 (N_353,In_31,In_226);
and U354 (N_354,N_340,N_333);
nand U355 (N_355,In_229,N_300);
or U356 (N_356,N_66,N_306);
xor U357 (N_357,N_313,In_320);
nand U358 (N_358,In_193,In_465);
nor U359 (N_359,N_336,N_318);
nor U360 (N_360,N_284,N_334);
and U361 (N_361,N_339,N_267);
nor U362 (N_362,N_252,In_91);
nor U363 (N_363,N_72,N_310);
nand U364 (N_364,In_322,In_294);
or U365 (N_365,N_245,N_256);
nand U366 (N_366,In_63,N_328);
or U367 (N_367,N_338,N_337);
xnor U368 (N_368,N_316,N_234);
nor U369 (N_369,N_305,In_233);
nand U370 (N_370,N_342,In_80);
and U371 (N_371,N_269,N_144);
nand U372 (N_372,N_253,In_464);
and U373 (N_373,N_261,N_322);
or U374 (N_374,N_348,In_345);
nor U375 (N_375,N_315,In_182);
nor U376 (N_376,N_153,N_276);
nand U377 (N_377,In_354,N_200);
and U378 (N_378,N_258,N_311);
or U379 (N_379,N_296,N_172);
xnor U380 (N_380,N_217,N_10);
xor U381 (N_381,N_304,N_283);
or U382 (N_382,N_312,In_252);
and U383 (N_383,N_254,In_98);
and U384 (N_384,N_319,N_347);
and U385 (N_385,In_450,N_247);
nand U386 (N_386,In_395,In_147);
nand U387 (N_387,N_8,N_330);
nor U388 (N_388,N_158,N_65);
and U389 (N_389,N_298,In_302);
nor U390 (N_390,N_320,N_223);
nand U391 (N_391,N_331,N_341);
nand U392 (N_392,N_329,N_265);
xor U393 (N_393,In_425,In_317);
and U394 (N_394,N_303,N_263);
nor U395 (N_395,N_191,In_378);
or U396 (N_396,In_156,N_280);
and U397 (N_397,N_190,N_196);
and U398 (N_398,N_309,N_288);
or U399 (N_399,N_291,N_177);
nand U400 (N_400,N_363,N_345);
nor U401 (N_401,N_360,N_367);
nor U402 (N_402,N_387,N_335);
or U403 (N_403,N_332,N_194);
or U404 (N_404,N_321,N_369);
nor U405 (N_405,In_407,N_399);
nand U406 (N_406,N_389,N_327);
and U407 (N_407,In_218,N_344);
and U408 (N_408,N_398,N_355);
nand U409 (N_409,In_33,N_166);
xnor U410 (N_410,In_97,N_385);
nor U411 (N_411,N_383,In_73);
xnor U412 (N_412,N_353,N_375);
nor U413 (N_413,N_382,N_366);
or U414 (N_414,N_139,N_308);
nor U415 (N_415,N_346,N_357);
or U416 (N_416,N_395,N_292);
or U417 (N_417,N_392,N_55);
nand U418 (N_418,N_255,In_65);
and U419 (N_419,N_362,N_250);
or U420 (N_420,N_351,N_86);
nor U421 (N_421,N_352,N_324);
xnor U422 (N_422,N_391,N_386);
and U423 (N_423,N_364,In_171);
or U424 (N_424,N_268,N_368);
and U425 (N_425,N_343,N_384);
nor U426 (N_426,N_221,N_358);
nor U427 (N_427,N_371,In_282);
xor U428 (N_428,N_326,N_307);
or U429 (N_429,N_289,N_393);
or U430 (N_430,N_317,In_381);
xnor U431 (N_431,N_251,N_394);
and U432 (N_432,N_359,N_377);
nor U433 (N_433,N_361,N_396);
nor U434 (N_434,In_456,N_374);
or U435 (N_435,N_373,N_354);
nand U436 (N_436,N_380,In_443);
and U437 (N_437,In_152,N_262);
nand U438 (N_438,N_219,N_390);
nor U439 (N_439,N_379,N_378);
nor U440 (N_440,N_376,N_349);
and U441 (N_441,N_193,N_325);
xor U442 (N_442,N_208,N_231);
xor U443 (N_443,In_397,N_323);
or U444 (N_444,N_143,N_350);
and U445 (N_445,N_372,N_356);
nor U446 (N_446,N_301,N_388);
and U447 (N_447,N_46,N_370);
or U448 (N_448,In_124,N_381);
or U449 (N_449,N_365,N_397);
or U450 (N_450,N_405,N_421);
and U451 (N_451,N_447,N_416);
and U452 (N_452,N_422,N_431);
nor U453 (N_453,N_409,N_448);
nand U454 (N_454,N_446,N_444);
or U455 (N_455,N_407,N_406);
and U456 (N_456,N_437,N_436);
xor U457 (N_457,N_435,N_423);
nand U458 (N_458,N_419,N_428);
or U459 (N_459,N_414,N_410);
or U460 (N_460,N_432,N_439);
nand U461 (N_461,N_433,N_445);
and U462 (N_462,N_427,N_440);
xnor U463 (N_463,N_413,N_415);
nor U464 (N_464,N_403,N_429);
or U465 (N_465,N_441,N_418);
xor U466 (N_466,N_400,N_408);
or U467 (N_467,N_424,N_425);
or U468 (N_468,N_402,N_443);
xor U469 (N_469,N_412,N_420);
or U470 (N_470,N_411,N_434);
and U471 (N_471,N_417,N_404);
xor U472 (N_472,N_430,N_449);
or U473 (N_473,N_438,N_442);
or U474 (N_474,N_426,N_401);
or U475 (N_475,N_428,N_400);
or U476 (N_476,N_425,N_449);
nand U477 (N_477,N_410,N_412);
and U478 (N_478,N_422,N_438);
nor U479 (N_479,N_427,N_442);
and U480 (N_480,N_441,N_433);
nor U481 (N_481,N_406,N_420);
nor U482 (N_482,N_410,N_447);
nor U483 (N_483,N_425,N_404);
nand U484 (N_484,N_415,N_417);
or U485 (N_485,N_440,N_445);
xor U486 (N_486,N_437,N_438);
nand U487 (N_487,N_424,N_421);
and U488 (N_488,N_437,N_440);
and U489 (N_489,N_437,N_428);
or U490 (N_490,N_401,N_409);
xor U491 (N_491,N_412,N_442);
and U492 (N_492,N_403,N_437);
xor U493 (N_493,N_427,N_415);
xnor U494 (N_494,N_446,N_406);
nor U495 (N_495,N_445,N_441);
nand U496 (N_496,N_435,N_418);
nand U497 (N_497,N_430,N_427);
and U498 (N_498,N_409,N_427);
xnor U499 (N_499,N_412,N_448);
xor U500 (N_500,N_494,N_455);
nor U501 (N_501,N_483,N_479);
nor U502 (N_502,N_498,N_451);
xnor U503 (N_503,N_469,N_486);
xnor U504 (N_504,N_464,N_480);
or U505 (N_505,N_466,N_468);
nand U506 (N_506,N_457,N_473);
or U507 (N_507,N_460,N_471);
xnor U508 (N_508,N_462,N_496);
nor U509 (N_509,N_465,N_485);
or U510 (N_510,N_474,N_470);
xor U511 (N_511,N_459,N_493);
nor U512 (N_512,N_454,N_450);
nand U513 (N_513,N_481,N_497);
nor U514 (N_514,N_472,N_488);
xor U515 (N_515,N_499,N_456);
or U516 (N_516,N_492,N_487);
xnor U517 (N_517,N_495,N_461);
and U518 (N_518,N_458,N_452);
nor U519 (N_519,N_478,N_490);
and U520 (N_520,N_463,N_475);
nand U521 (N_521,N_482,N_484);
xnor U522 (N_522,N_453,N_491);
nor U523 (N_523,N_467,N_489);
nand U524 (N_524,N_476,N_477);
nor U525 (N_525,N_477,N_454);
nor U526 (N_526,N_497,N_456);
or U527 (N_527,N_495,N_482);
nor U528 (N_528,N_469,N_471);
and U529 (N_529,N_469,N_490);
nand U530 (N_530,N_481,N_484);
nor U531 (N_531,N_452,N_454);
nor U532 (N_532,N_494,N_459);
nor U533 (N_533,N_490,N_472);
nor U534 (N_534,N_475,N_480);
nor U535 (N_535,N_468,N_454);
xor U536 (N_536,N_494,N_470);
nand U537 (N_537,N_487,N_465);
xor U538 (N_538,N_475,N_469);
nand U539 (N_539,N_478,N_483);
and U540 (N_540,N_485,N_450);
or U541 (N_541,N_481,N_492);
or U542 (N_542,N_499,N_452);
nand U543 (N_543,N_485,N_474);
nand U544 (N_544,N_466,N_465);
xnor U545 (N_545,N_457,N_490);
nand U546 (N_546,N_464,N_495);
nor U547 (N_547,N_483,N_451);
or U548 (N_548,N_478,N_458);
nand U549 (N_549,N_499,N_498);
or U550 (N_550,N_518,N_510);
nor U551 (N_551,N_506,N_533);
or U552 (N_552,N_519,N_500);
nor U553 (N_553,N_516,N_529);
xor U554 (N_554,N_544,N_547);
xor U555 (N_555,N_505,N_530);
and U556 (N_556,N_523,N_540);
nand U557 (N_557,N_534,N_527);
nand U558 (N_558,N_512,N_526);
xnor U559 (N_559,N_521,N_532);
nor U560 (N_560,N_520,N_528);
or U561 (N_561,N_513,N_537);
and U562 (N_562,N_524,N_522);
nor U563 (N_563,N_508,N_536);
and U564 (N_564,N_538,N_525);
xnor U565 (N_565,N_509,N_502);
nand U566 (N_566,N_545,N_507);
or U567 (N_567,N_501,N_504);
nand U568 (N_568,N_503,N_539);
nor U569 (N_569,N_535,N_511);
nor U570 (N_570,N_549,N_517);
xnor U571 (N_571,N_541,N_531);
nand U572 (N_572,N_514,N_543);
nor U573 (N_573,N_546,N_548);
nor U574 (N_574,N_542,N_515);
or U575 (N_575,N_543,N_531);
nor U576 (N_576,N_520,N_543);
nand U577 (N_577,N_546,N_549);
or U578 (N_578,N_530,N_541);
nor U579 (N_579,N_505,N_503);
nand U580 (N_580,N_540,N_527);
nor U581 (N_581,N_515,N_530);
and U582 (N_582,N_500,N_512);
nor U583 (N_583,N_540,N_503);
and U584 (N_584,N_503,N_541);
and U585 (N_585,N_530,N_533);
nand U586 (N_586,N_539,N_546);
nor U587 (N_587,N_531,N_518);
and U588 (N_588,N_516,N_533);
or U589 (N_589,N_542,N_516);
nand U590 (N_590,N_516,N_501);
and U591 (N_591,N_521,N_514);
xor U592 (N_592,N_511,N_517);
nor U593 (N_593,N_545,N_501);
nor U594 (N_594,N_514,N_532);
xnor U595 (N_595,N_501,N_517);
nand U596 (N_596,N_544,N_538);
nor U597 (N_597,N_526,N_507);
nor U598 (N_598,N_500,N_544);
and U599 (N_599,N_508,N_507);
and U600 (N_600,N_576,N_588);
or U601 (N_601,N_589,N_564);
nand U602 (N_602,N_560,N_569);
or U603 (N_603,N_554,N_587);
nor U604 (N_604,N_582,N_567);
and U605 (N_605,N_573,N_556);
or U606 (N_606,N_598,N_558);
xor U607 (N_607,N_583,N_551);
xnor U608 (N_608,N_553,N_585);
xnor U609 (N_609,N_579,N_591);
or U610 (N_610,N_562,N_575);
or U611 (N_611,N_571,N_597);
and U612 (N_612,N_565,N_599);
and U613 (N_613,N_563,N_550);
xnor U614 (N_614,N_570,N_586);
nor U615 (N_615,N_559,N_561);
nor U616 (N_616,N_577,N_593);
xnor U617 (N_617,N_568,N_578);
nand U618 (N_618,N_584,N_594);
nand U619 (N_619,N_595,N_580);
nor U620 (N_620,N_555,N_574);
nor U621 (N_621,N_581,N_590);
xor U622 (N_622,N_566,N_557);
xor U623 (N_623,N_596,N_572);
nor U624 (N_624,N_552,N_592);
xnor U625 (N_625,N_584,N_596);
nor U626 (N_626,N_593,N_561);
nor U627 (N_627,N_584,N_556);
nand U628 (N_628,N_586,N_582);
xnor U629 (N_629,N_577,N_568);
nor U630 (N_630,N_556,N_555);
or U631 (N_631,N_589,N_597);
or U632 (N_632,N_553,N_570);
or U633 (N_633,N_587,N_557);
nor U634 (N_634,N_591,N_570);
and U635 (N_635,N_571,N_555);
and U636 (N_636,N_594,N_597);
nor U637 (N_637,N_569,N_595);
nor U638 (N_638,N_582,N_571);
xor U639 (N_639,N_582,N_556);
nor U640 (N_640,N_556,N_583);
or U641 (N_641,N_571,N_596);
nor U642 (N_642,N_584,N_563);
or U643 (N_643,N_565,N_558);
or U644 (N_644,N_596,N_579);
nand U645 (N_645,N_579,N_565);
nand U646 (N_646,N_588,N_563);
xnor U647 (N_647,N_576,N_579);
or U648 (N_648,N_554,N_551);
nand U649 (N_649,N_571,N_573);
nand U650 (N_650,N_613,N_619);
and U651 (N_651,N_623,N_631);
and U652 (N_652,N_603,N_635);
nor U653 (N_653,N_634,N_609);
nor U654 (N_654,N_622,N_600);
nand U655 (N_655,N_637,N_642);
xor U656 (N_656,N_643,N_617);
and U657 (N_657,N_636,N_612);
or U658 (N_658,N_646,N_618);
nor U659 (N_659,N_620,N_608);
and U660 (N_660,N_602,N_601);
nor U661 (N_661,N_611,N_629);
nor U662 (N_662,N_640,N_625);
nand U663 (N_663,N_606,N_627);
or U664 (N_664,N_624,N_633);
nand U665 (N_665,N_607,N_614);
nor U666 (N_666,N_649,N_638);
nor U667 (N_667,N_630,N_604);
nand U668 (N_668,N_626,N_644);
nand U669 (N_669,N_615,N_639);
nor U670 (N_670,N_641,N_610);
and U671 (N_671,N_605,N_645);
or U672 (N_672,N_616,N_648);
xnor U673 (N_673,N_647,N_628);
nor U674 (N_674,N_632,N_621);
xnor U675 (N_675,N_638,N_647);
nand U676 (N_676,N_613,N_620);
and U677 (N_677,N_637,N_618);
and U678 (N_678,N_620,N_605);
and U679 (N_679,N_647,N_644);
nand U680 (N_680,N_639,N_643);
or U681 (N_681,N_637,N_646);
and U682 (N_682,N_636,N_621);
nor U683 (N_683,N_643,N_644);
xnor U684 (N_684,N_603,N_620);
and U685 (N_685,N_609,N_629);
or U686 (N_686,N_628,N_630);
nand U687 (N_687,N_617,N_646);
and U688 (N_688,N_623,N_626);
or U689 (N_689,N_649,N_646);
xnor U690 (N_690,N_617,N_609);
and U691 (N_691,N_635,N_608);
and U692 (N_692,N_645,N_630);
nand U693 (N_693,N_644,N_614);
and U694 (N_694,N_640,N_603);
and U695 (N_695,N_621,N_642);
nand U696 (N_696,N_624,N_645);
or U697 (N_697,N_619,N_640);
nand U698 (N_698,N_637,N_611);
nand U699 (N_699,N_615,N_620);
nand U700 (N_700,N_680,N_697);
xor U701 (N_701,N_650,N_678);
nor U702 (N_702,N_688,N_654);
xnor U703 (N_703,N_663,N_656);
nand U704 (N_704,N_683,N_651);
nor U705 (N_705,N_660,N_690);
nor U706 (N_706,N_664,N_667);
or U707 (N_707,N_677,N_675);
nand U708 (N_708,N_657,N_693);
xnor U709 (N_709,N_679,N_691);
nor U710 (N_710,N_659,N_686);
xor U711 (N_711,N_695,N_687);
xnor U712 (N_712,N_694,N_698);
or U713 (N_713,N_652,N_665);
and U714 (N_714,N_672,N_653);
xor U715 (N_715,N_661,N_684);
nand U716 (N_716,N_662,N_670);
nand U717 (N_717,N_682,N_669);
and U718 (N_718,N_674,N_689);
nand U719 (N_719,N_658,N_666);
nand U720 (N_720,N_676,N_671);
and U721 (N_721,N_692,N_668);
and U722 (N_722,N_673,N_699);
xor U723 (N_723,N_655,N_681);
nand U724 (N_724,N_696,N_685);
or U725 (N_725,N_675,N_660);
nor U726 (N_726,N_683,N_691);
nand U727 (N_727,N_676,N_697);
nor U728 (N_728,N_689,N_693);
xor U729 (N_729,N_691,N_653);
or U730 (N_730,N_696,N_652);
xnor U731 (N_731,N_678,N_685);
or U732 (N_732,N_688,N_681);
nand U733 (N_733,N_654,N_690);
or U734 (N_734,N_678,N_657);
nand U735 (N_735,N_678,N_656);
nand U736 (N_736,N_661,N_680);
nor U737 (N_737,N_676,N_654);
or U738 (N_738,N_671,N_668);
nor U739 (N_739,N_673,N_665);
xor U740 (N_740,N_689,N_656);
or U741 (N_741,N_678,N_692);
nor U742 (N_742,N_695,N_689);
nor U743 (N_743,N_691,N_662);
or U744 (N_744,N_673,N_691);
or U745 (N_745,N_653,N_664);
nand U746 (N_746,N_670,N_694);
and U747 (N_747,N_677,N_699);
nand U748 (N_748,N_693,N_652);
and U749 (N_749,N_656,N_676);
nor U750 (N_750,N_744,N_727);
and U751 (N_751,N_737,N_728);
or U752 (N_752,N_748,N_710);
nor U753 (N_753,N_701,N_741);
or U754 (N_754,N_733,N_707);
and U755 (N_755,N_745,N_709);
nor U756 (N_756,N_747,N_729);
xor U757 (N_757,N_704,N_739);
or U758 (N_758,N_713,N_725);
xnor U759 (N_759,N_711,N_723);
and U760 (N_760,N_717,N_730);
nand U761 (N_761,N_703,N_746);
and U762 (N_762,N_714,N_724);
and U763 (N_763,N_734,N_735);
and U764 (N_764,N_705,N_706);
and U765 (N_765,N_722,N_726);
and U766 (N_766,N_721,N_708);
or U767 (N_767,N_718,N_731);
xor U768 (N_768,N_716,N_732);
nand U769 (N_769,N_749,N_740);
xor U770 (N_770,N_719,N_715);
and U771 (N_771,N_720,N_712);
nor U772 (N_772,N_742,N_736);
xnor U773 (N_773,N_743,N_702);
xor U774 (N_774,N_700,N_738);
or U775 (N_775,N_732,N_700);
xor U776 (N_776,N_740,N_710);
nand U777 (N_777,N_706,N_731);
and U778 (N_778,N_746,N_737);
nand U779 (N_779,N_723,N_743);
nor U780 (N_780,N_730,N_739);
nand U781 (N_781,N_714,N_739);
or U782 (N_782,N_713,N_717);
or U783 (N_783,N_744,N_714);
or U784 (N_784,N_718,N_704);
xor U785 (N_785,N_716,N_729);
or U786 (N_786,N_702,N_707);
nand U787 (N_787,N_706,N_734);
and U788 (N_788,N_724,N_722);
nand U789 (N_789,N_747,N_744);
xor U790 (N_790,N_701,N_744);
and U791 (N_791,N_723,N_703);
and U792 (N_792,N_708,N_734);
xor U793 (N_793,N_732,N_717);
or U794 (N_794,N_716,N_747);
nor U795 (N_795,N_733,N_722);
and U796 (N_796,N_729,N_721);
nand U797 (N_797,N_747,N_738);
nand U798 (N_798,N_718,N_720);
nor U799 (N_799,N_709,N_746);
and U800 (N_800,N_765,N_768);
xor U801 (N_801,N_757,N_784);
nor U802 (N_802,N_760,N_753);
nand U803 (N_803,N_796,N_752);
xor U804 (N_804,N_793,N_786);
nor U805 (N_805,N_758,N_782);
nor U806 (N_806,N_799,N_750);
xor U807 (N_807,N_785,N_783);
nor U808 (N_808,N_789,N_797);
nand U809 (N_809,N_776,N_774);
xnor U810 (N_810,N_763,N_790);
and U811 (N_811,N_764,N_781);
or U812 (N_812,N_771,N_772);
nor U813 (N_813,N_754,N_788);
xor U814 (N_814,N_780,N_761);
or U815 (N_815,N_777,N_795);
nor U816 (N_816,N_755,N_775);
and U817 (N_817,N_770,N_791);
or U818 (N_818,N_766,N_767);
or U819 (N_819,N_787,N_798);
nand U820 (N_820,N_751,N_762);
nor U821 (N_821,N_769,N_759);
nor U822 (N_822,N_792,N_778);
nor U823 (N_823,N_756,N_779);
and U824 (N_824,N_794,N_773);
xnor U825 (N_825,N_782,N_753);
xnor U826 (N_826,N_750,N_791);
xnor U827 (N_827,N_796,N_793);
and U828 (N_828,N_754,N_760);
and U829 (N_829,N_761,N_764);
xnor U830 (N_830,N_790,N_769);
nor U831 (N_831,N_752,N_782);
and U832 (N_832,N_760,N_771);
or U833 (N_833,N_750,N_765);
xor U834 (N_834,N_772,N_763);
and U835 (N_835,N_798,N_759);
nor U836 (N_836,N_789,N_777);
xnor U837 (N_837,N_760,N_751);
and U838 (N_838,N_752,N_776);
nor U839 (N_839,N_753,N_787);
and U840 (N_840,N_778,N_758);
or U841 (N_841,N_779,N_751);
nor U842 (N_842,N_759,N_797);
nand U843 (N_843,N_757,N_796);
or U844 (N_844,N_798,N_790);
and U845 (N_845,N_766,N_798);
and U846 (N_846,N_780,N_760);
or U847 (N_847,N_763,N_791);
nand U848 (N_848,N_791,N_753);
and U849 (N_849,N_797,N_773);
and U850 (N_850,N_845,N_804);
nor U851 (N_851,N_843,N_849);
and U852 (N_852,N_832,N_819);
or U853 (N_853,N_815,N_821);
and U854 (N_854,N_830,N_829);
or U855 (N_855,N_842,N_825);
and U856 (N_856,N_801,N_810);
or U857 (N_857,N_835,N_814);
xnor U858 (N_858,N_816,N_831);
xnor U859 (N_859,N_813,N_811);
and U860 (N_860,N_836,N_833);
or U861 (N_861,N_838,N_824);
xnor U862 (N_862,N_803,N_808);
and U863 (N_863,N_812,N_822);
or U864 (N_864,N_800,N_818);
and U865 (N_865,N_805,N_827);
or U866 (N_866,N_809,N_834);
and U867 (N_867,N_837,N_844);
nand U868 (N_868,N_847,N_846);
and U869 (N_869,N_848,N_817);
and U870 (N_870,N_820,N_839);
and U871 (N_871,N_840,N_806);
nand U872 (N_872,N_802,N_841);
or U873 (N_873,N_807,N_826);
or U874 (N_874,N_828,N_823);
nor U875 (N_875,N_816,N_803);
nand U876 (N_876,N_824,N_837);
nand U877 (N_877,N_846,N_819);
nand U878 (N_878,N_827,N_822);
nor U879 (N_879,N_837,N_825);
nand U880 (N_880,N_831,N_819);
or U881 (N_881,N_831,N_806);
or U882 (N_882,N_801,N_833);
or U883 (N_883,N_824,N_812);
xor U884 (N_884,N_831,N_817);
xnor U885 (N_885,N_803,N_814);
and U886 (N_886,N_800,N_836);
nor U887 (N_887,N_829,N_846);
and U888 (N_888,N_845,N_833);
nand U889 (N_889,N_813,N_817);
and U890 (N_890,N_818,N_805);
nor U891 (N_891,N_804,N_838);
or U892 (N_892,N_847,N_836);
nand U893 (N_893,N_828,N_840);
xor U894 (N_894,N_835,N_808);
xor U895 (N_895,N_815,N_835);
nand U896 (N_896,N_840,N_826);
and U897 (N_897,N_818,N_839);
xor U898 (N_898,N_825,N_834);
and U899 (N_899,N_844,N_849);
and U900 (N_900,N_883,N_865);
xor U901 (N_901,N_899,N_861);
and U902 (N_902,N_879,N_857);
or U903 (N_903,N_895,N_863);
xnor U904 (N_904,N_864,N_853);
or U905 (N_905,N_850,N_882);
nor U906 (N_906,N_852,N_891);
or U907 (N_907,N_892,N_888);
nand U908 (N_908,N_893,N_860);
and U909 (N_909,N_887,N_869);
nor U910 (N_910,N_884,N_871);
nand U911 (N_911,N_897,N_878);
nand U912 (N_912,N_862,N_874);
or U913 (N_913,N_881,N_898);
xor U914 (N_914,N_855,N_896);
and U915 (N_915,N_872,N_876);
or U916 (N_916,N_873,N_889);
xnor U917 (N_917,N_866,N_890);
and U918 (N_918,N_877,N_880);
nor U919 (N_919,N_894,N_859);
nand U920 (N_920,N_886,N_858);
or U921 (N_921,N_885,N_868);
or U922 (N_922,N_875,N_851);
nor U923 (N_923,N_854,N_867);
xor U924 (N_924,N_870,N_856);
nand U925 (N_925,N_886,N_893);
or U926 (N_926,N_877,N_851);
xnor U927 (N_927,N_899,N_875);
nand U928 (N_928,N_873,N_884);
nor U929 (N_929,N_887,N_866);
xor U930 (N_930,N_883,N_855);
xnor U931 (N_931,N_853,N_875);
nand U932 (N_932,N_898,N_893);
or U933 (N_933,N_857,N_861);
nand U934 (N_934,N_898,N_884);
nand U935 (N_935,N_896,N_862);
nand U936 (N_936,N_864,N_882);
nand U937 (N_937,N_871,N_859);
xor U938 (N_938,N_888,N_859);
nand U939 (N_939,N_853,N_865);
nand U940 (N_940,N_850,N_872);
or U941 (N_941,N_877,N_886);
and U942 (N_942,N_873,N_870);
or U943 (N_943,N_853,N_896);
nand U944 (N_944,N_892,N_876);
nand U945 (N_945,N_891,N_896);
nand U946 (N_946,N_887,N_862);
or U947 (N_947,N_892,N_883);
xor U948 (N_948,N_896,N_861);
and U949 (N_949,N_863,N_886);
xor U950 (N_950,N_900,N_901);
and U951 (N_951,N_933,N_925);
and U952 (N_952,N_908,N_918);
or U953 (N_953,N_920,N_939);
nand U954 (N_954,N_917,N_929);
nor U955 (N_955,N_937,N_912);
and U956 (N_956,N_913,N_927);
nand U957 (N_957,N_909,N_945);
and U958 (N_958,N_944,N_936);
nand U959 (N_959,N_904,N_931);
or U960 (N_960,N_949,N_922);
nor U961 (N_961,N_926,N_930);
nand U962 (N_962,N_914,N_943);
nor U963 (N_963,N_916,N_915);
nor U964 (N_964,N_940,N_928);
nor U965 (N_965,N_906,N_941);
nor U966 (N_966,N_924,N_907);
nand U967 (N_967,N_923,N_942);
nor U968 (N_968,N_932,N_935);
and U969 (N_969,N_934,N_902);
nand U970 (N_970,N_948,N_938);
nor U971 (N_971,N_911,N_919);
and U972 (N_972,N_903,N_905);
nor U973 (N_973,N_921,N_946);
nand U974 (N_974,N_947,N_910);
nor U975 (N_975,N_905,N_928);
nor U976 (N_976,N_942,N_935);
xnor U977 (N_977,N_914,N_940);
nand U978 (N_978,N_908,N_936);
xnor U979 (N_979,N_933,N_922);
xnor U980 (N_980,N_934,N_904);
or U981 (N_981,N_905,N_927);
nand U982 (N_982,N_935,N_915);
nor U983 (N_983,N_923,N_929);
nand U984 (N_984,N_948,N_910);
nor U985 (N_985,N_949,N_913);
nand U986 (N_986,N_947,N_922);
and U987 (N_987,N_928,N_930);
or U988 (N_988,N_937,N_907);
nor U989 (N_989,N_933,N_935);
or U990 (N_990,N_905,N_910);
nand U991 (N_991,N_927,N_933);
xnor U992 (N_992,N_920,N_947);
or U993 (N_993,N_947,N_934);
xor U994 (N_994,N_944,N_932);
xnor U995 (N_995,N_925,N_938);
and U996 (N_996,N_933,N_946);
nor U997 (N_997,N_903,N_915);
xor U998 (N_998,N_939,N_942);
xor U999 (N_999,N_908,N_929);
nor U1000 (N_1000,N_956,N_960);
xnor U1001 (N_1001,N_968,N_988);
xnor U1002 (N_1002,N_977,N_951);
nor U1003 (N_1003,N_962,N_963);
or U1004 (N_1004,N_983,N_967);
xor U1005 (N_1005,N_973,N_959);
and U1006 (N_1006,N_985,N_971);
xnor U1007 (N_1007,N_991,N_989);
and U1008 (N_1008,N_972,N_974);
and U1009 (N_1009,N_984,N_997);
nand U1010 (N_1010,N_987,N_969);
nor U1011 (N_1011,N_994,N_996);
or U1012 (N_1012,N_979,N_966);
and U1013 (N_1013,N_955,N_990);
xor U1014 (N_1014,N_953,N_998);
xor U1015 (N_1015,N_976,N_958);
xor U1016 (N_1016,N_982,N_980);
or U1017 (N_1017,N_978,N_992);
xor U1018 (N_1018,N_954,N_970);
and U1019 (N_1019,N_950,N_952);
nand U1020 (N_1020,N_957,N_995);
xnor U1021 (N_1021,N_993,N_975);
nand U1022 (N_1022,N_965,N_999);
and U1023 (N_1023,N_986,N_981);
and U1024 (N_1024,N_961,N_964);
and U1025 (N_1025,N_997,N_988);
nor U1026 (N_1026,N_979,N_982);
and U1027 (N_1027,N_960,N_955);
xnor U1028 (N_1028,N_970,N_968);
or U1029 (N_1029,N_950,N_959);
and U1030 (N_1030,N_978,N_999);
or U1031 (N_1031,N_990,N_951);
nor U1032 (N_1032,N_976,N_953);
and U1033 (N_1033,N_959,N_989);
nand U1034 (N_1034,N_988,N_956);
xnor U1035 (N_1035,N_953,N_954);
nor U1036 (N_1036,N_996,N_960);
nand U1037 (N_1037,N_987,N_960);
xnor U1038 (N_1038,N_993,N_953);
nand U1039 (N_1039,N_988,N_978);
or U1040 (N_1040,N_968,N_962);
xor U1041 (N_1041,N_959,N_977);
and U1042 (N_1042,N_973,N_960);
or U1043 (N_1043,N_999,N_983);
or U1044 (N_1044,N_975,N_970);
nor U1045 (N_1045,N_989,N_995);
or U1046 (N_1046,N_978,N_997);
nor U1047 (N_1047,N_963,N_950);
and U1048 (N_1048,N_981,N_961);
nand U1049 (N_1049,N_965,N_981);
nand U1050 (N_1050,N_1032,N_1010);
and U1051 (N_1051,N_1012,N_1011);
xor U1052 (N_1052,N_1042,N_1035);
nor U1053 (N_1053,N_1026,N_1008);
nand U1054 (N_1054,N_1031,N_1044);
nor U1055 (N_1055,N_1018,N_1003);
or U1056 (N_1056,N_1037,N_1034);
nor U1057 (N_1057,N_1019,N_1045);
nand U1058 (N_1058,N_1007,N_1030);
or U1059 (N_1059,N_1027,N_1023);
xor U1060 (N_1060,N_1041,N_1036);
or U1061 (N_1061,N_1040,N_1028);
nand U1062 (N_1062,N_1013,N_1029);
xor U1063 (N_1063,N_1000,N_1006);
xnor U1064 (N_1064,N_1021,N_1005);
xor U1065 (N_1065,N_1002,N_1017);
or U1066 (N_1066,N_1001,N_1014);
nand U1067 (N_1067,N_1020,N_1049);
xnor U1068 (N_1068,N_1043,N_1024);
nand U1069 (N_1069,N_1048,N_1033);
or U1070 (N_1070,N_1004,N_1015);
or U1071 (N_1071,N_1038,N_1025);
nor U1072 (N_1072,N_1009,N_1046);
nand U1073 (N_1073,N_1039,N_1047);
nor U1074 (N_1074,N_1016,N_1022);
nor U1075 (N_1075,N_1049,N_1007);
xor U1076 (N_1076,N_1000,N_1035);
nor U1077 (N_1077,N_1039,N_1028);
nor U1078 (N_1078,N_1049,N_1035);
and U1079 (N_1079,N_1013,N_1033);
nor U1080 (N_1080,N_1047,N_1032);
nand U1081 (N_1081,N_1023,N_1022);
nand U1082 (N_1082,N_1008,N_1002);
and U1083 (N_1083,N_1044,N_1007);
nand U1084 (N_1084,N_1030,N_1006);
or U1085 (N_1085,N_1040,N_1007);
and U1086 (N_1086,N_1043,N_1005);
nand U1087 (N_1087,N_1026,N_1029);
xor U1088 (N_1088,N_1038,N_1002);
nand U1089 (N_1089,N_1031,N_1046);
xor U1090 (N_1090,N_1006,N_1018);
xor U1091 (N_1091,N_1036,N_1018);
or U1092 (N_1092,N_1014,N_1049);
and U1093 (N_1093,N_1037,N_1000);
or U1094 (N_1094,N_1035,N_1037);
nand U1095 (N_1095,N_1038,N_1031);
xnor U1096 (N_1096,N_1037,N_1007);
xor U1097 (N_1097,N_1027,N_1010);
xor U1098 (N_1098,N_1008,N_1004);
and U1099 (N_1099,N_1024,N_1000);
or U1100 (N_1100,N_1092,N_1079);
nand U1101 (N_1101,N_1069,N_1083);
xnor U1102 (N_1102,N_1088,N_1098);
xnor U1103 (N_1103,N_1061,N_1065);
nor U1104 (N_1104,N_1053,N_1051);
xnor U1105 (N_1105,N_1099,N_1062);
xor U1106 (N_1106,N_1067,N_1070);
or U1107 (N_1107,N_1080,N_1094);
xor U1108 (N_1108,N_1085,N_1093);
nor U1109 (N_1109,N_1055,N_1077);
nor U1110 (N_1110,N_1068,N_1081);
nand U1111 (N_1111,N_1073,N_1056);
xnor U1112 (N_1112,N_1066,N_1072);
or U1113 (N_1113,N_1091,N_1090);
nor U1114 (N_1114,N_1064,N_1074);
nand U1115 (N_1115,N_1097,N_1078);
or U1116 (N_1116,N_1096,N_1054);
nand U1117 (N_1117,N_1071,N_1060);
or U1118 (N_1118,N_1057,N_1059);
nor U1119 (N_1119,N_1076,N_1063);
nor U1120 (N_1120,N_1087,N_1050);
and U1121 (N_1121,N_1095,N_1075);
and U1122 (N_1122,N_1086,N_1082);
and U1123 (N_1123,N_1058,N_1089);
nor U1124 (N_1124,N_1084,N_1052);
nand U1125 (N_1125,N_1077,N_1070);
and U1126 (N_1126,N_1059,N_1087);
or U1127 (N_1127,N_1078,N_1052);
xor U1128 (N_1128,N_1058,N_1095);
xnor U1129 (N_1129,N_1051,N_1079);
xnor U1130 (N_1130,N_1069,N_1082);
nand U1131 (N_1131,N_1094,N_1066);
or U1132 (N_1132,N_1093,N_1064);
nor U1133 (N_1133,N_1071,N_1098);
xor U1134 (N_1134,N_1082,N_1064);
nor U1135 (N_1135,N_1052,N_1059);
or U1136 (N_1136,N_1097,N_1089);
xor U1137 (N_1137,N_1068,N_1053);
or U1138 (N_1138,N_1072,N_1067);
nor U1139 (N_1139,N_1098,N_1083);
nor U1140 (N_1140,N_1077,N_1097);
or U1141 (N_1141,N_1097,N_1071);
nor U1142 (N_1142,N_1082,N_1077);
and U1143 (N_1143,N_1068,N_1088);
nand U1144 (N_1144,N_1073,N_1063);
nand U1145 (N_1145,N_1096,N_1076);
and U1146 (N_1146,N_1090,N_1075);
nor U1147 (N_1147,N_1066,N_1067);
or U1148 (N_1148,N_1087,N_1089);
nand U1149 (N_1149,N_1090,N_1096);
nand U1150 (N_1150,N_1133,N_1103);
or U1151 (N_1151,N_1145,N_1121);
xnor U1152 (N_1152,N_1108,N_1128);
nor U1153 (N_1153,N_1101,N_1131);
and U1154 (N_1154,N_1144,N_1125);
and U1155 (N_1155,N_1126,N_1104);
xor U1156 (N_1156,N_1122,N_1123);
and U1157 (N_1157,N_1118,N_1117);
xnor U1158 (N_1158,N_1148,N_1127);
xnor U1159 (N_1159,N_1107,N_1130);
nand U1160 (N_1160,N_1114,N_1106);
nor U1161 (N_1161,N_1141,N_1134);
or U1162 (N_1162,N_1100,N_1142);
nor U1163 (N_1163,N_1111,N_1137);
and U1164 (N_1164,N_1129,N_1116);
and U1165 (N_1165,N_1102,N_1120);
nor U1166 (N_1166,N_1143,N_1113);
or U1167 (N_1167,N_1147,N_1136);
nor U1168 (N_1168,N_1138,N_1124);
xor U1169 (N_1169,N_1105,N_1146);
nor U1170 (N_1170,N_1110,N_1132);
or U1171 (N_1171,N_1109,N_1112);
and U1172 (N_1172,N_1149,N_1135);
xor U1173 (N_1173,N_1140,N_1139);
and U1174 (N_1174,N_1115,N_1119);
nand U1175 (N_1175,N_1123,N_1119);
nand U1176 (N_1176,N_1130,N_1132);
nor U1177 (N_1177,N_1141,N_1105);
xnor U1178 (N_1178,N_1146,N_1141);
nor U1179 (N_1179,N_1125,N_1122);
nand U1180 (N_1180,N_1136,N_1108);
nand U1181 (N_1181,N_1128,N_1135);
nor U1182 (N_1182,N_1103,N_1136);
or U1183 (N_1183,N_1141,N_1124);
nand U1184 (N_1184,N_1142,N_1110);
and U1185 (N_1185,N_1100,N_1126);
nand U1186 (N_1186,N_1140,N_1112);
nand U1187 (N_1187,N_1140,N_1100);
or U1188 (N_1188,N_1137,N_1124);
xnor U1189 (N_1189,N_1106,N_1135);
and U1190 (N_1190,N_1115,N_1107);
xor U1191 (N_1191,N_1131,N_1149);
or U1192 (N_1192,N_1109,N_1114);
nand U1193 (N_1193,N_1141,N_1106);
nor U1194 (N_1194,N_1129,N_1133);
nor U1195 (N_1195,N_1120,N_1114);
xor U1196 (N_1196,N_1101,N_1124);
or U1197 (N_1197,N_1126,N_1116);
xor U1198 (N_1198,N_1104,N_1106);
or U1199 (N_1199,N_1134,N_1115);
and U1200 (N_1200,N_1183,N_1159);
or U1201 (N_1201,N_1193,N_1199);
or U1202 (N_1202,N_1160,N_1175);
nand U1203 (N_1203,N_1158,N_1176);
xor U1204 (N_1204,N_1150,N_1190);
nor U1205 (N_1205,N_1187,N_1179);
or U1206 (N_1206,N_1153,N_1165);
nand U1207 (N_1207,N_1173,N_1169);
and U1208 (N_1208,N_1180,N_1162);
nand U1209 (N_1209,N_1171,N_1184);
nor U1210 (N_1210,N_1177,N_1155);
and U1211 (N_1211,N_1152,N_1186);
nand U1212 (N_1212,N_1181,N_1157);
nand U1213 (N_1213,N_1166,N_1156);
and U1214 (N_1214,N_1164,N_1161);
or U1215 (N_1215,N_1197,N_1151);
xor U1216 (N_1216,N_1192,N_1170);
nand U1217 (N_1217,N_1172,N_1182);
nand U1218 (N_1218,N_1178,N_1196);
and U1219 (N_1219,N_1174,N_1191);
and U1220 (N_1220,N_1167,N_1189);
and U1221 (N_1221,N_1195,N_1185);
xnor U1222 (N_1222,N_1188,N_1198);
or U1223 (N_1223,N_1154,N_1168);
or U1224 (N_1224,N_1194,N_1163);
or U1225 (N_1225,N_1192,N_1179);
or U1226 (N_1226,N_1191,N_1167);
xor U1227 (N_1227,N_1197,N_1166);
and U1228 (N_1228,N_1157,N_1198);
and U1229 (N_1229,N_1177,N_1158);
or U1230 (N_1230,N_1172,N_1188);
nand U1231 (N_1231,N_1176,N_1160);
or U1232 (N_1232,N_1174,N_1154);
nand U1233 (N_1233,N_1163,N_1189);
or U1234 (N_1234,N_1186,N_1164);
nor U1235 (N_1235,N_1159,N_1196);
xor U1236 (N_1236,N_1160,N_1166);
nor U1237 (N_1237,N_1190,N_1194);
xor U1238 (N_1238,N_1194,N_1154);
nand U1239 (N_1239,N_1178,N_1181);
xor U1240 (N_1240,N_1177,N_1170);
or U1241 (N_1241,N_1194,N_1162);
nand U1242 (N_1242,N_1198,N_1197);
or U1243 (N_1243,N_1193,N_1160);
or U1244 (N_1244,N_1182,N_1168);
nor U1245 (N_1245,N_1186,N_1173);
nand U1246 (N_1246,N_1175,N_1196);
nand U1247 (N_1247,N_1196,N_1188);
or U1248 (N_1248,N_1192,N_1190);
and U1249 (N_1249,N_1185,N_1154);
xor U1250 (N_1250,N_1200,N_1212);
nand U1251 (N_1251,N_1209,N_1232);
nor U1252 (N_1252,N_1217,N_1204);
and U1253 (N_1253,N_1226,N_1210);
nor U1254 (N_1254,N_1231,N_1211);
nand U1255 (N_1255,N_1236,N_1216);
and U1256 (N_1256,N_1233,N_1249);
nand U1257 (N_1257,N_1243,N_1246);
nand U1258 (N_1258,N_1228,N_1229);
xnor U1259 (N_1259,N_1242,N_1202);
or U1260 (N_1260,N_1225,N_1237);
nand U1261 (N_1261,N_1247,N_1207);
nor U1262 (N_1262,N_1219,N_1240);
xnor U1263 (N_1263,N_1214,N_1235);
nor U1264 (N_1264,N_1224,N_1215);
or U1265 (N_1265,N_1239,N_1205);
or U1266 (N_1266,N_1241,N_1230);
nand U1267 (N_1267,N_1223,N_1244);
xnor U1268 (N_1268,N_1206,N_1248);
or U1269 (N_1269,N_1245,N_1238);
xor U1270 (N_1270,N_1227,N_1221);
nand U1271 (N_1271,N_1201,N_1234);
nor U1272 (N_1272,N_1218,N_1208);
nor U1273 (N_1273,N_1220,N_1222);
and U1274 (N_1274,N_1203,N_1213);
and U1275 (N_1275,N_1213,N_1202);
xor U1276 (N_1276,N_1224,N_1222);
or U1277 (N_1277,N_1226,N_1239);
or U1278 (N_1278,N_1235,N_1212);
nand U1279 (N_1279,N_1239,N_1244);
or U1280 (N_1280,N_1242,N_1203);
and U1281 (N_1281,N_1223,N_1214);
and U1282 (N_1282,N_1234,N_1224);
or U1283 (N_1283,N_1212,N_1232);
or U1284 (N_1284,N_1227,N_1206);
nor U1285 (N_1285,N_1236,N_1239);
nor U1286 (N_1286,N_1232,N_1220);
nand U1287 (N_1287,N_1248,N_1215);
nor U1288 (N_1288,N_1208,N_1216);
and U1289 (N_1289,N_1241,N_1200);
nand U1290 (N_1290,N_1229,N_1211);
or U1291 (N_1291,N_1247,N_1228);
nor U1292 (N_1292,N_1223,N_1210);
and U1293 (N_1293,N_1216,N_1249);
xnor U1294 (N_1294,N_1238,N_1229);
and U1295 (N_1295,N_1213,N_1249);
or U1296 (N_1296,N_1223,N_1235);
xnor U1297 (N_1297,N_1207,N_1212);
or U1298 (N_1298,N_1224,N_1227);
xor U1299 (N_1299,N_1234,N_1225);
or U1300 (N_1300,N_1256,N_1292);
nor U1301 (N_1301,N_1251,N_1271);
nor U1302 (N_1302,N_1274,N_1293);
nor U1303 (N_1303,N_1255,N_1288);
nor U1304 (N_1304,N_1253,N_1254);
xnor U1305 (N_1305,N_1278,N_1299);
or U1306 (N_1306,N_1273,N_1298);
xnor U1307 (N_1307,N_1268,N_1262);
nand U1308 (N_1308,N_1284,N_1283);
and U1309 (N_1309,N_1270,N_1252);
or U1310 (N_1310,N_1282,N_1263);
xnor U1311 (N_1311,N_1265,N_1250);
or U1312 (N_1312,N_1286,N_1291);
or U1313 (N_1313,N_1275,N_1276);
or U1314 (N_1314,N_1260,N_1267);
nand U1315 (N_1315,N_1277,N_1297);
or U1316 (N_1316,N_1258,N_1295);
and U1317 (N_1317,N_1296,N_1261);
nor U1318 (N_1318,N_1294,N_1290);
xor U1319 (N_1319,N_1272,N_1280);
or U1320 (N_1320,N_1257,N_1259);
or U1321 (N_1321,N_1281,N_1287);
or U1322 (N_1322,N_1264,N_1279);
nand U1323 (N_1323,N_1289,N_1269);
nor U1324 (N_1324,N_1266,N_1285);
nor U1325 (N_1325,N_1264,N_1290);
xnor U1326 (N_1326,N_1288,N_1256);
nand U1327 (N_1327,N_1282,N_1250);
and U1328 (N_1328,N_1270,N_1266);
nand U1329 (N_1329,N_1279,N_1265);
nor U1330 (N_1330,N_1277,N_1268);
and U1331 (N_1331,N_1280,N_1289);
nor U1332 (N_1332,N_1263,N_1258);
or U1333 (N_1333,N_1253,N_1277);
nand U1334 (N_1334,N_1261,N_1288);
or U1335 (N_1335,N_1258,N_1252);
or U1336 (N_1336,N_1291,N_1285);
nand U1337 (N_1337,N_1294,N_1297);
and U1338 (N_1338,N_1278,N_1279);
nor U1339 (N_1339,N_1276,N_1297);
and U1340 (N_1340,N_1296,N_1275);
or U1341 (N_1341,N_1293,N_1273);
xnor U1342 (N_1342,N_1260,N_1259);
xnor U1343 (N_1343,N_1289,N_1287);
and U1344 (N_1344,N_1254,N_1259);
and U1345 (N_1345,N_1257,N_1265);
or U1346 (N_1346,N_1268,N_1264);
nand U1347 (N_1347,N_1262,N_1272);
xor U1348 (N_1348,N_1265,N_1251);
nor U1349 (N_1349,N_1269,N_1286);
nand U1350 (N_1350,N_1305,N_1338);
and U1351 (N_1351,N_1343,N_1324);
nand U1352 (N_1352,N_1349,N_1322);
nor U1353 (N_1353,N_1311,N_1334);
and U1354 (N_1354,N_1308,N_1307);
nand U1355 (N_1355,N_1317,N_1300);
and U1356 (N_1356,N_1326,N_1327);
or U1357 (N_1357,N_1301,N_1304);
and U1358 (N_1358,N_1325,N_1336);
nand U1359 (N_1359,N_1319,N_1318);
xor U1360 (N_1360,N_1345,N_1347);
xnor U1361 (N_1361,N_1346,N_1302);
nor U1362 (N_1362,N_1310,N_1330);
nand U1363 (N_1363,N_1303,N_1342);
nor U1364 (N_1364,N_1315,N_1314);
xnor U1365 (N_1365,N_1341,N_1348);
and U1366 (N_1366,N_1309,N_1316);
or U1367 (N_1367,N_1313,N_1344);
and U1368 (N_1368,N_1337,N_1306);
nand U1369 (N_1369,N_1323,N_1312);
xor U1370 (N_1370,N_1332,N_1331);
and U1371 (N_1371,N_1340,N_1333);
xor U1372 (N_1372,N_1328,N_1320);
nor U1373 (N_1373,N_1321,N_1335);
and U1374 (N_1374,N_1329,N_1339);
nand U1375 (N_1375,N_1337,N_1309);
or U1376 (N_1376,N_1349,N_1340);
or U1377 (N_1377,N_1324,N_1340);
xnor U1378 (N_1378,N_1344,N_1326);
xnor U1379 (N_1379,N_1304,N_1344);
and U1380 (N_1380,N_1305,N_1309);
nor U1381 (N_1381,N_1307,N_1339);
nor U1382 (N_1382,N_1325,N_1334);
or U1383 (N_1383,N_1300,N_1311);
nor U1384 (N_1384,N_1305,N_1326);
nand U1385 (N_1385,N_1341,N_1332);
or U1386 (N_1386,N_1340,N_1311);
nor U1387 (N_1387,N_1309,N_1330);
nand U1388 (N_1388,N_1339,N_1343);
or U1389 (N_1389,N_1346,N_1315);
nor U1390 (N_1390,N_1336,N_1320);
and U1391 (N_1391,N_1308,N_1332);
nor U1392 (N_1392,N_1340,N_1326);
or U1393 (N_1393,N_1313,N_1318);
and U1394 (N_1394,N_1301,N_1316);
xnor U1395 (N_1395,N_1347,N_1341);
or U1396 (N_1396,N_1336,N_1343);
or U1397 (N_1397,N_1341,N_1321);
nand U1398 (N_1398,N_1341,N_1323);
nand U1399 (N_1399,N_1328,N_1319);
nand U1400 (N_1400,N_1390,N_1391);
and U1401 (N_1401,N_1355,N_1364);
nand U1402 (N_1402,N_1384,N_1354);
nand U1403 (N_1403,N_1353,N_1363);
xnor U1404 (N_1404,N_1376,N_1380);
xor U1405 (N_1405,N_1358,N_1378);
xnor U1406 (N_1406,N_1394,N_1373);
nor U1407 (N_1407,N_1386,N_1374);
and U1408 (N_1408,N_1397,N_1370);
nor U1409 (N_1409,N_1362,N_1393);
xor U1410 (N_1410,N_1385,N_1372);
and U1411 (N_1411,N_1371,N_1383);
xnor U1412 (N_1412,N_1360,N_1398);
or U1413 (N_1413,N_1395,N_1351);
xnor U1414 (N_1414,N_1392,N_1382);
or U1415 (N_1415,N_1368,N_1375);
and U1416 (N_1416,N_1387,N_1356);
or U1417 (N_1417,N_1357,N_1359);
nand U1418 (N_1418,N_1367,N_1388);
or U1419 (N_1419,N_1381,N_1399);
xnor U1420 (N_1420,N_1396,N_1350);
or U1421 (N_1421,N_1366,N_1377);
and U1422 (N_1422,N_1369,N_1389);
or U1423 (N_1423,N_1352,N_1365);
nand U1424 (N_1424,N_1379,N_1361);
and U1425 (N_1425,N_1350,N_1394);
or U1426 (N_1426,N_1385,N_1386);
xnor U1427 (N_1427,N_1397,N_1357);
nor U1428 (N_1428,N_1374,N_1361);
nor U1429 (N_1429,N_1355,N_1373);
or U1430 (N_1430,N_1378,N_1370);
or U1431 (N_1431,N_1357,N_1394);
nor U1432 (N_1432,N_1353,N_1366);
nor U1433 (N_1433,N_1367,N_1357);
nor U1434 (N_1434,N_1366,N_1397);
xor U1435 (N_1435,N_1370,N_1354);
nand U1436 (N_1436,N_1356,N_1377);
nor U1437 (N_1437,N_1370,N_1368);
and U1438 (N_1438,N_1378,N_1360);
nand U1439 (N_1439,N_1390,N_1355);
or U1440 (N_1440,N_1377,N_1374);
nor U1441 (N_1441,N_1363,N_1359);
nand U1442 (N_1442,N_1356,N_1365);
nor U1443 (N_1443,N_1372,N_1380);
or U1444 (N_1444,N_1361,N_1352);
and U1445 (N_1445,N_1356,N_1358);
or U1446 (N_1446,N_1366,N_1364);
or U1447 (N_1447,N_1373,N_1393);
nor U1448 (N_1448,N_1354,N_1395);
nor U1449 (N_1449,N_1382,N_1390);
or U1450 (N_1450,N_1406,N_1411);
nand U1451 (N_1451,N_1401,N_1441);
xnor U1452 (N_1452,N_1409,N_1419);
and U1453 (N_1453,N_1423,N_1417);
nand U1454 (N_1454,N_1443,N_1440);
and U1455 (N_1455,N_1432,N_1418);
nand U1456 (N_1456,N_1430,N_1408);
nor U1457 (N_1457,N_1446,N_1449);
nand U1458 (N_1458,N_1447,N_1435);
nand U1459 (N_1459,N_1427,N_1442);
nand U1460 (N_1460,N_1425,N_1437);
or U1461 (N_1461,N_1405,N_1415);
xor U1462 (N_1462,N_1444,N_1439);
or U1463 (N_1463,N_1429,N_1407);
or U1464 (N_1464,N_1420,N_1433);
nand U1465 (N_1465,N_1438,N_1403);
nor U1466 (N_1466,N_1422,N_1434);
nand U1467 (N_1467,N_1410,N_1416);
or U1468 (N_1468,N_1421,N_1413);
or U1469 (N_1469,N_1424,N_1412);
nor U1470 (N_1470,N_1400,N_1436);
or U1471 (N_1471,N_1414,N_1428);
nand U1472 (N_1472,N_1448,N_1426);
or U1473 (N_1473,N_1445,N_1402);
xor U1474 (N_1474,N_1431,N_1404);
nand U1475 (N_1475,N_1449,N_1423);
nand U1476 (N_1476,N_1445,N_1443);
or U1477 (N_1477,N_1422,N_1415);
nand U1478 (N_1478,N_1404,N_1421);
and U1479 (N_1479,N_1436,N_1417);
and U1480 (N_1480,N_1439,N_1404);
nor U1481 (N_1481,N_1423,N_1432);
nor U1482 (N_1482,N_1407,N_1406);
and U1483 (N_1483,N_1444,N_1413);
nor U1484 (N_1484,N_1409,N_1403);
nand U1485 (N_1485,N_1448,N_1436);
and U1486 (N_1486,N_1415,N_1403);
or U1487 (N_1487,N_1406,N_1448);
or U1488 (N_1488,N_1412,N_1449);
xor U1489 (N_1489,N_1440,N_1431);
or U1490 (N_1490,N_1438,N_1423);
and U1491 (N_1491,N_1430,N_1400);
xnor U1492 (N_1492,N_1417,N_1404);
or U1493 (N_1493,N_1438,N_1434);
and U1494 (N_1494,N_1410,N_1424);
xnor U1495 (N_1495,N_1443,N_1442);
xnor U1496 (N_1496,N_1445,N_1414);
or U1497 (N_1497,N_1417,N_1415);
and U1498 (N_1498,N_1437,N_1414);
nor U1499 (N_1499,N_1435,N_1438);
xor U1500 (N_1500,N_1481,N_1490);
or U1501 (N_1501,N_1456,N_1473);
xor U1502 (N_1502,N_1475,N_1464);
nor U1503 (N_1503,N_1469,N_1480);
and U1504 (N_1504,N_1492,N_1467);
and U1505 (N_1505,N_1451,N_1450);
and U1506 (N_1506,N_1468,N_1459);
nand U1507 (N_1507,N_1496,N_1457);
xnor U1508 (N_1508,N_1482,N_1478);
or U1509 (N_1509,N_1470,N_1489);
or U1510 (N_1510,N_1466,N_1463);
nand U1511 (N_1511,N_1474,N_1488);
nor U1512 (N_1512,N_1491,N_1486);
or U1513 (N_1513,N_1494,N_1499);
nand U1514 (N_1514,N_1484,N_1485);
and U1515 (N_1515,N_1452,N_1471);
nor U1516 (N_1516,N_1465,N_1479);
nand U1517 (N_1517,N_1460,N_1498);
xor U1518 (N_1518,N_1462,N_1461);
nor U1519 (N_1519,N_1497,N_1493);
xnor U1520 (N_1520,N_1483,N_1453);
xor U1521 (N_1521,N_1495,N_1454);
xor U1522 (N_1522,N_1458,N_1455);
nand U1523 (N_1523,N_1476,N_1472);
nor U1524 (N_1524,N_1477,N_1487);
nand U1525 (N_1525,N_1487,N_1497);
or U1526 (N_1526,N_1451,N_1452);
nor U1527 (N_1527,N_1473,N_1494);
or U1528 (N_1528,N_1474,N_1493);
xnor U1529 (N_1529,N_1482,N_1483);
nor U1530 (N_1530,N_1488,N_1490);
and U1531 (N_1531,N_1464,N_1486);
xor U1532 (N_1532,N_1451,N_1463);
or U1533 (N_1533,N_1453,N_1463);
nand U1534 (N_1534,N_1477,N_1453);
or U1535 (N_1535,N_1494,N_1498);
and U1536 (N_1536,N_1479,N_1475);
and U1537 (N_1537,N_1456,N_1490);
nor U1538 (N_1538,N_1483,N_1496);
and U1539 (N_1539,N_1462,N_1483);
nand U1540 (N_1540,N_1466,N_1470);
and U1541 (N_1541,N_1468,N_1454);
nor U1542 (N_1542,N_1462,N_1465);
xnor U1543 (N_1543,N_1468,N_1465);
or U1544 (N_1544,N_1460,N_1488);
nor U1545 (N_1545,N_1458,N_1470);
nor U1546 (N_1546,N_1459,N_1499);
nand U1547 (N_1547,N_1451,N_1477);
nor U1548 (N_1548,N_1464,N_1463);
or U1549 (N_1549,N_1474,N_1471);
nand U1550 (N_1550,N_1504,N_1545);
or U1551 (N_1551,N_1536,N_1520);
xor U1552 (N_1552,N_1537,N_1531);
nand U1553 (N_1553,N_1506,N_1516);
or U1554 (N_1554,N_1519,N_1548);
nand U1555 (N_1555,N_1511,N_1522);
nand U1556 (N_1556,N_1508,N_1538);
or U1557 (N_1557,N_1518,N_1533);
or U1558 (N_1558,N_1505,N_1527);
xnor U1559 (N_1559,N_1544,N_1507);
or U1560 (N_1560,N_1521,N_1503);
and U1561 (N_1561,N_1524,N_1501);
nor U1562 (N_1562,N_1542,N_1509);
xnor U1563 (N_1563,N_1530,N_1500);
and U1564 (N_1564,N_1541,N_1535);
or U1565 (N_1565,N_1546,N_1543);
and U1566 (N_1566,N_1540,N_1514);
and U1567 (N_1567,N_1549,N_1534);
and U1568 (N_1568,N_1526,N_1510);
and U1569 (N_1569,N_1512,N_1528);
nand U1570 (N_1570,N_1515,N_1539);
and U1571 (N_1571,N_1525,N_1523);
nand U1572 (N_1572,N_1532,N_1529);
nor U1573 (N_1573,N_1513,N_1547);
xnor U1574 (N_1574,N_1502,N_1517);
xnor U1575 (N_1575,N_1507,N_1509);
nor U1576 (N_1576,N_1500,N_1522);
and U1577 (N_1577,N_1520,N_1528);
and U1578 (N_1578,N_1546,N_1504);
or U1579 (N_1579,N_1505,N_1541);
xor U1580 (N_1580,N_1511,N_1517);
nand U1581 (N_1581,N_1535,N_1547);
nor U1582 (N_1582,N_1536,N_1524);
xor U1583 (N_1583,N_1537,N_1507);
nand U1584 (N_1584,N_1500,N_1519);
nor U1585 (N_1585,N_1545,N_1508);
xor U1586 (N_1586,N_1544,N_1512);
and U1587 (N_1587,N_1532,N_1530);
or U1588 (N_1588,N_1542,N_1520);
and U1589 (N_1589,N_1538,N_1515);
or U1590 (N_1590,N_1548,N_1534);
and U1591 (N_1591,N_1500,N_1516);
xor U1592 (N_1592,N_1512,N_1529);
nor U1593 (N_1593,N_1522,N_1526);
or U1594 (N_1594,N_1548,N_1505);
xor U1595 (N_1595,N_1502,N_1540);
or U1596 (N_1596,N_1533,N_1541);
or U1597 (N_1597,N_1500,N_1521);
nor U1598 (N_1598,N_1543,N_1533);
and U1599 (N_1599,N_1524,N_1549);
nand U1600 (N_1600,N_1591,N_1570);
nand U1601 (N_1601,N_1576,N_1599);
nand U1602 (N_1602,N_1569,N_1586);
nand U1603 (N_1603,N_1588,N_1565);
xnor U1604 (N_1604,N_1564,N_1560);
nand U1605 (N_1605,N_1551,N_1597);
nor U1606 (N_1606,N_1587,N_1555);
and U1607 (N_1607,N_1577,N_1579);
nor U1608 (N_1608,N_1582,N_1573);
or U1609 (N_1609,N_1559,N_1585);
nor U1610 (N_1610,N_1553,N_1572);
nor U1611 (N_1611,N_1561,N_1590);
nand U1612 (N_1612,N_1578,N_1557);
nand U1613 (N_1613,N_1584,N_1574);
and U1614 (N_1614,N_1556,N_1581);
xnor U1615 (N_1615,N_1566,N_1562);
or U1616 (N_1616,N_1558,N_1575);
nor U1617 (N_1617,N_1598,N_1594);
or U1618 (N_1618,N_1554,N_1592);
nand U1619 (N_1619,N_1583,N_1593);
nor U1620 (N_1620,N_1571,N_1568);
xor U1621 (N_1621,N_1563,N_1550);
nand U1622 (N_1622,N_1552,N_1580);
and U1623 (N_1623,N_1595,N_1596);
nand U1624 (N_1624,N_1567,N_1589);
xor U1625 (N_1625,N_1579,N_1552);
nor U1626 (N_1626,N_1599,N_1559);
nor U1627 (N_1627,N_1568,N_1552);
or U1628 (N_1628,N_1587,N_1552);
or U1629 (N_1629,N_1593,N_1579);
nor U1630 (N_1630,N_1576,N_1568);
nor U1631 (N_1631,N_1574,N_1592);
and U1632 (N_1632,N_1574,N_1572);
nor U1633 (N_1633,N_1596,N_1578);
and U1634 (N_1634,N_1560,N_1555);
nand U1635 (N_1635,N_1571,N_1563);
nor U1636 (N_1636,N_1558,N_1572);
xnor U1637 (N_1637,N_1584,N_1599);
xnor U1638 (N_1638,N_1578,N_1591);
or U1639 (N_1639,N_1578,N_1564);
nor U1640 (N_1640,N_1560,N_1585);
xor U1641 (N_1641,N_1590,N_1565);
xnor U1642 (N_1642,N_1592,N_1581);
nand U1643 (N_1643,N_1590,N_1578);
nand U1644 (N_1644,N_1597,N_1577);
xnor U1645 (N_1645,N_1587,N_1572);
or U1646 (N_1646,N_1550,N_1564);
nand U1647 (N_1647,N_1584,N_1598);
and U1648 (N_1648,N_1555,N_1559);
xnor U1649 (N_1649,N_1578,N_1589);
xor U1650 (N_1650,N_1606,N_1611);
nor U1651 (N_1651,N_1634,N_1633);
nor U1652 (N_1652,N_1622,N_1628);
nor U1653 (N_1653,N_1608,N_1638);
xnor U1654 (N_1654,N_1630,N_1648);
and U1655 (N_1655,N_1649,N_1619);
nand U1656 (N_1656,N_1626,N_1604);
nand U1657 (N_1657,N_1620,N_1643);
nor U1658 (N_1658,N_1618,N_1610);
nor U1659 (N_1659,N_1645,N_1636);
and U1660 (N_1660,N_1639,N_1600);
and U1661 (N_1661,N_1641,N_1609);
and U1662 (N_1662,N_1613,N_1640);
nor U1663 (N_1663,N_1642,N_1602);
nand U1664 (N_1664,N_1635,N_1605);
or U1665 (N_1665,N_1614,N_1603);
nor U1666 (N_1666,N_1621,N_1629);
nand U1667 (N_1667,N_1612,N_1632);
nand U1668 (N_1668,N_1644,N_1616);
or U1669 (N_1669,N_1607,N_1615);
nand U1670 (N_1670,N_1637,N_1624);
or U1671 (N_1671,N_1623,N_1627);
nand U1672 (N_1672,N_1631,N_1646);
nor U1673 (N_1673,N_1617,N_1625);
or U1674 (N_1674,N_1601,N_1647);
nand U1675 (N_1675,N_1632,N_1643);
xnor U1676 (N_1676,N_1631,N_1637);
and U1677 (N_1677,N_1622,N_1615);
nand U1678 (N_1678,N_1627,N_1642);
and U1679 (N_1679,N_1643,N_1616);
nor U1680 (N_1680,N_1632,N_1633);
nand U1681 (N_1681,N_1607,N_1638);
or U1682 (N_1682,N_1630,N_1647);
or U1683 (N_1683,N_1630,N_1604);
nand U1684 (N_1684,N_1625,N_1629);
and U1685 (N_1685,N_1625,N_1609);
nand U1686 (N_1686,N_1625,N_1616);
nand U1687 (N_1687,N_1616,N_1615);
or U1688 (N_1688,N_1608,N_1623);
nor U1689 (N_1689,N_1633,N_1647);
nor U1690 (N_1690,N_1603,N_1632);
nor U1691 (N_1691,N_1626,N_1647);
and U1692 (N_1692,N_1633,N_1627);
or U1693 (N_1693,N_1623,N_1635);
or U1694 (N_1694,N_1620,N_1629);
nand U1695 (N_1695,N_1646,N_1612);
nand U1696 (N_1696,N_1626,N_1605);
and U1697 (N_1697,N_1648,N_1644);
and U1698 (N_1698,N_1630,N_1645);
nand U1699 (N_1699,N_1626,N_1616);
nor U1700 (N_1700,N_1694,N_1665);
nand U1701 (N_1701,N_1662,N_1657);
or U1702 (N_1702,N_1674,N_1655);
or U1703 (N_1703,N_1660,N_1678);
xor U1704 (N_1704,N_1676,N_1698);
xnor U1705 (N_1705,N_1699,N_1654);
or U1706 (N_1706,N_1686,N_1690);
nor U1707 (N_1707,N_1675,N_1668);
and U1708 (N_1708,N_1684,N_1697);
and U1709 (N_1709,N_1669,N_1670);
xnor U1710 (N_1710,N_1687,N_1695);
or U1711 (N_1711,N_1682,N_1650);
nor U1712 (N_1712,N_1692,N_1681);
nand U1713 (N_1713,N_1656,N_1663);
xnor U1714 (N_1714,N_1679,N_1688);
or U1715 (N_1715,N_1652,N_1677);
nor U1716 (N_1716,N_1653,N_1672);
nand U1717 (N_1717,N_1658,N_1691);
or U1718 (N_1718,N_1651,N_1685);
xor U1719 (N_1719,N_1689,N_1693);
and U1720 (N_1720,N_1661,N_1671);
or U1721 (N_1721,N_1696,N_1666);
nor U1722 (N_1722,N_1667,N_1683);
xnor U1723 (N_1723,N_1659,N_1680);
nor U1724 (N_1724,N_1673,N_1664);
nor U1725 (N_1725,N_1693,N_1697);
or U1726 (N_1726,N_1688,N_1670);
or U1727 (N_1727,N_1688,N_1696);
nand U1728 (N_1728,N_1665,N_1673);
and U1729 (N_1729,N_1672,N_1685);
nand U1730 (N_1730,N_1699,N_1688);
or U1731 (N_1731,N_1692,N_1665);
nand U1732 (N_1732,N_1676,N_1670);
and U1733 (N_1733,N_1679,N_1654);
xnor U1734 (N_1734,N_1667,N_1663);
or U1735 (N_1735,N_1666,N_1658);
and U1736 (N_1736,N_1686,N_1664);
and U1737 (N_1737,N_1671,N_1653);
xor U1738 (N_1738,N_1662,N_1658);
or U1739 (N_1739,N_1676,N_1688);
nand U1740 (N_1740,N_1681,N_1679);
or U1741 (N_1741,N_1692,N_1655);
xor U1742 (N_1742,N_1694,N_1675);
and U1743 (N_1743,N_1671,N_1687);
or U1744 (N_1744,N_1694,N_1683);
and U1745 (N_1745,N_1686,N_1681);
or U1746 (N_1746,N_1688,N_1651);
xor U1747 (N_1747,N_1674,N_1684);
nand U1748 (N_1748,N_1692,N_1678);
or U1749 (N_1749,N_1654,N_1698);
nor U1750 (N_1750,N_1716,N_1741);
and U1751 (N_1751,N_1703,N_1732);
nand U1752 (N_1752,N_1728,N_1727);
nand U1753 (N_1753,N_1710,N_1711);
xor U1754 (N_1754,N_1749,N_1734);
xnor U1755 (N_1755,N_1707,N_1721);
or U1756 (N_1756,N_1705,N_1747);
or U1757 (N_1757,N_1738,N_1702);
nand U1758 (N_1758,N_1737,N_1739);
and U1759 (N_1759,N_1712,N_1743);
and U1760 (N_1760,N_1713,N_1736);
xnor U1761 (N_1761,N_1730,N_1733);
and U1762 (N_1762,N_1719,N_1744);
xor U1763 (N_1763,N_1700,N_1740);
or U1764 (N_1764,N_1746,N_1722);
and U1765 (N_1765,N_1724,N_1701);
xor U1766 (N_1766,N_1748,N_1745);
nor U1767 (N_1767,N_1717,N_1729);
and U1768 (N_1768,N_1704,N_1726);
xnor U1769 (N_1769,N_1735,N_1714);
and U1770 (N_1770,N_1723,N_1715);
or U1771 (N_1771,N_1718,N_1706);
nand U1772 (N_1772,N_1720,N_1731);
xnor U1773 (N_1773,N_1709,N_1742);
and U1774 (N_1774,N_1725,N_1708);
nand U1775 (N_1775,N_1708,N_1713);
xnor U1776 (N_1776,N_1749,N_1701);
xnor U1777 (N_1777,N_1719,N_1736);
nand U1778 (N_1778,N_1704,N_1732);
nor U1779 (N_1779,N_1745,N_1701);
or U1780 (N_1780,N_1727,N_1741);
nor U1781 (N_1781,N_1732,N_1730);
nor U1782 (N_1782,N_1713,N_1705);
xor U1783 (N_1783,N_1700,N_1720);
xnor U1784 (N_1784,N_1713,N_1732);
and U1785 (N_1785,N_1714,N_1704);
nor U1786 (N_1786,N_1715,N_1719);
or U1787 (N_1787,N_1730,N_1702);
and U1788 (N_1788,N_1715,N_1714);
xnor U1789 (N_1789,N_1709,N_1724);
nand U1790 (N_1790,N_1728,N_1726);
xnor U1791 (N_1791,N_1738,N_1742);
nand U1792 (N_1792,N_1706,N_1743);
nand U1793 (N_1793,N_1707,N_1746);
nand U1794 (N_1794,N_1710,N_1720);
xor U1795 (N_1795,N_1722,N_1709);
or U1796 (N_1796,N_1743,N_1738);
and U1797 (N_1797,N_1722,N_1720);
nand U1798 (N_1798,N_1747,N_1723);
and U1799 (N_1799,N_1744,N_1733);
and U1800 (N_1800,N_1790,N_1775);
or U1801 (N_1801,N_1788,N_1765);
and U1802 (N_1802,N_1779,N_1770);
and U1803 (N_1803,N_1778,N_1771);
nor U1804 (N_1804,N_1767,N_1796);
or U1805 (N_1805,N_1793,N_1795);
or U1806 (N_1806,N_1786,N_1764);
or U1807 (N_1807,N_1768,N_1784);
nand U1808 (N_1808,N_1777,N_1762);
nor U1809 (N_1809,N_1753,N_1755);
xor U1810 (N_1810,N_1752,N_1750);
and U1811 (N_1811,N_1781,N_1789);
nor U1812 (N_1812,N_1756,N_1769);
nand U1813 (N_1813,N_1763,N_1751);
nor U1814 (N_1814,N_1798,N_1797);
and U1815 (N_1815,N_1792,N_1754);
nand U1816 (N_1816,N_1794,N_1787);
xor U1817 (N_1817,N_1766,N_1785);
and U1818 (N_1818,N_1776,N_1799);
nor U1819 (N_1819,N_1757,N_1791);
nor U1820 (N_1820,N_1774,N_1780);
nand U1821 (N_1821,N_1773,N_1761);
and U1822 (N_1822,N_1758,N_1759);
nor U1823 (N_1823,N_1760,N_1783);
nand U1824 (N_1824,N_1772,N_1782);
xnor U1825 (N_1825,N_1753,N_1783);
nor U1826 (N_1826,N_1763,N_1787);
nor U1827 (N_1827,N_1753,N_1777);
nor U1828 (N_1828,N_1787,N_1767);
nor U1829 (N_1829,N_1775,N_1767);
or U1830 (N_1830,N_1760,N_1776);
or U1831 (N_1831,N_1778,N_1755);
or U1832 (N_1832,N_1761,N_1779);
and U1833 (N_1833,N_1764,N_1788);
nand U1834 (N_1834,N_1752,N_1758);
or U1835 (N_1835,N_1797,N_1795);
nor U1836 (N_1836,N_1774,N_1752);
xor U1837 (N_1837,N_1760,N_1773);
nor U1838 (N_1838,N_1770,N_1792);
xor U1839 (N_1839,N_1766,N_1795);
or U1840 (N_1840,N_1791,N_1792);
and U1841 (N_1841,N_1772,N_1757);
nor U1842 (N_1842,N_1796,N_1763);
or U1843 (N_1843,N_1763,N_1768);
and U1844 (N_1844,N_1789,N_1752);
nor U1845 (N_1845,N_1799,N_1763);
and U1846 (N_1846,N_1775,N_1798);
nor U1847 (N_1847,N_1797,N_1769);
nor U1848 (N_1848,N_1759,N_1768);
or U1849 (N_1849,N_1756,N_1799);
nand U1850 (N_1850,N_1845,N_1833);
nor U1851 (N_1851,N_1830,N_1818);
xnor U1852 (N_1852,N_1849,N_1806);
xor U1853 (N_1853,N_1813,N_1834);
nand U1854 (N_1854,N_1828,N_1844);
nand U1855 (N_1855,N_1816,N_1838);
or U1856 (N_1856,N_1835,N_1804);
or U1857 (N_1857,N_1846,N_1826);
and U1858 (N_1858,N_1841,N_1811);
nor U1859 (N_1859,N_1827,N_1810);
xnor U1860 (N_1860,N_1831,N_1802);
nand U1861 (N_1861,N_1820,N_1815);
or U1862 (N_1862,N_1825,N_1823);
nor U1863 (N_1863,N_1840,N_1812);
nand U1864 (N_1864,N_1848,N_1842);
and U1865 (N_1865,N_1829,N_1809);
and U1866 (N_1866,N_1807,N_1824);
and U1867 (N_1867,N_1832,N_1808);
and U1868 (N_1868,N_1819,N_1803);
nand U1869 (N_1869,N_1817,N_1847);
nand U1870 (N_1870,N_1843,N_1801);
and U1871 (N_1871,N_1821,N_1837);
nor U1872 (N_1872,N_1822,N_1800);
nand U1873 (N_1873,N_1836,N_1805);
nor U1874 (N_1874,N_1839,N_1814);
xor U1875 (N_1875,N_1811,N_1820);
xnor U1876 (N_1876,N_1819,N_1802);
and U1877 (N_1877,N_1834,N_1821);
nor U1878 (N_1878,N_1800,N_1834);
or U1879 (N_1879,N_1813,N_1848);
nor U1880 (N_1880,N_1846,N_1841);
or U1881 (N_1881,N_1841,N_1839);
xnor U1882 (N_1882,N_1801,N_1832);
nand U1883 (N_1883,N_1847,N_1812);
or U1884 (N_1884,N_1844,N_1825);
or U1885 (N_1885,N_1839,N_1829);
and U1886 (N_1886,N_1803,N_1804);
or U1887 (N_1887,N_1820,N_1803);
nand U1888 (N_1888,N_1802,N_1805);
nand U1889 (N_1889,N_1838,N_1814);
nor U1890 (N_1890,N_1806,N_1842);
xor U1891 (N_1891,N_1832,N_1816);
and U1892 (N_1892,N_1801,N_1836);
nor U1893 (N_1893,N_1846,N_1817);
nand U1894 (N_1894,N_1840,N_1817);
nand U1895 (N_1895,N_1849,N_1824);
nand U1896 (N_1896,N_1802,N_1801);
or U1897 (N_1897,N_1845,N_1839);
or U1898 (N_1898,N_1814,N_1800);
nor U1899 (N_1899,N_1832,N_1827);
nand U1900 (N_1900,N_1885,N_1860);
or U1901 (N_1901,N_1859,N_1858);
nand U1902 (N_1902,N_1883,N_1855);
nand U1903 (N_1903,N_1871,N_1856);
nand U1904 (N_1904,N_1875,N_1898);
nand U1905 (N_1905,N_1884,N_1893);
xnor U1906 (N_1906,N_1892,N_1873);
or U1907 (N_1907,N_1890,N_1895);
nand U1908 (N_1908,N_1862,N_1899);
or U1909 (N_1909,N_1865,N_1879);
nor U1910 (N_1910,N_1878,N_1897);
nand U1911 (N_1911,N_1881,N_1882);
xnor U1912 (N_1912,N_1870,N_1850);
and U1913 (N_1913,N_1857,N_1874);
or U1914 (N_1914,N_1891,N_1864);
xor U1915 (N_1915,N_1889,N_1869);
xnor U1916 (N_1916,N_1853,N_1861);
or U1917 (N_1917,N_1872,N_1880);
nor U1918 (N_1918,N_1886,N_1876);
xnor U1919 (N_1919,N_1854,N_1868);
and U1920 (N_1920,N_1877,N_1894);
or U1921 (N_1921,N_1888,N_1896);
or U1922 (N_1922,N_1866,N_1887);
xor U1923 (N_1923,N_1851,N_1867);
and U1924 (N_1924,N_1852,N_1863);
or U1925 (N_1925,N_1898,N_1866);
nand U1926 (N_1926,N_1882,N_1873);
nand U1927 (N_1927,N_1850,N_1861);
or U1928 (N_1928,N_1857,N_1851);
or U1929 (N_1929,N_1861,N_1883);
nand U1930 (N_1930,N_1898,N_1857);
nand U1931 (N_1931,N_1887,N_1864);
nor U1932 (N_1932,N_1891,N_1868);
nand U1933 (N_1933,N_1857,N_1858);
nand U1934 (N_1934,N_1875,N_1896);
nand U1935 (N_1935,N_1890,N_1857);
nor U1936 (N_1936,N_1866,N_1853);
xnor U1937 (N_1937,N_1879,N_1890);
xnor U1938 (N_1938,N_1894,N_1860);
xnor U1939 (N_1939,N_1850,N_1862);
xnor U1940 (N_1940,N_1870,N_1867);
nor U1941 (N_1941,N_1886,N_1870);
or U1942 (N_1942,N_1852,N_1877);
xor U1943 (N_1943,N_1897,N_1876);
and U1944 (N_1944,N_1864,N_1892);
and U1945 (N_1945,N_1891,N_1883);
nand U1946 (N_1946,N_1865,N_1895);
xnor U1947 (N_1947,N_1869,N_1875);
and U1948 (N_1948,N_1851,N_1899);
nand U1949 (N_1949,N_1869,N_1864);
or U1950 (N_1950,N_1935,N_1947);
or U1951 (N_1951,N_1926,N_1919);
nand U1952 (N_1952,N_1933,N_1928);
nor U1953 (N_1953,N_1941,N_1946);
nor U1954 (N_1954,N_1939,N_1927);
nand U1955 (N_1955,N_1929,N_1916);
or U1956 (N_1956,N_1923,N_1906);
nor U1957 (N_1957,N_1942,N_1943);
or U1958 (N_1958,N_1945,N_1949);
and U1959 (N_1959,N_1911,N_1940);
nand U1960 (N_1960,N_1944,N_1932);
and U1961 (N_1961,N_1905,N_1917);
or U1962 (N_1962,N_1909,N_1915);
and U1963 (N_1963,N_1910,N_1901);
xor U1964 (N_1964,N_1913,N_1934);
nor U1965 (N_1965,N_1904,N_1930);
xnor U1966 (N_1966,N_1924,N_1936);
nand U1967 (N_1967,N_1918,N_1922);
and U1968 (N_1968,N_1920,N_1921);
and U1969 (N_1969,N_1931,N_1908);
nand U1970 (N_1970,N_1937,N_1914);
nand U1971 (N_1971,N_1902,N_1907);
xnor U1972 (N_1972,N_1900,N_1912);
and U1973 (N_1973,N_1925,N_1938);
and U1974 (N_1974,N_1903,N_1948);
or U1975 (N_1975,N_1913,N_1912);
and U1976 (N_1976,N_1927,N_1915);
xor U1977 (N_1977,N_1900,N_1904);
or U1978 (N_1978,N_1915,N_1907);
nand U1979 (N_1979,N_1933,N_1912);
nor U1980 (N_1980,N_1943,N_1911);
or U1981 (N_1981,N_1929,N_1935);
xor U1982 (N_1982,N_1945,N_1944);
or U1983 (N_1983,N_1923,N_1944);
nand U1984 (N_1984,N_1922,N_1924);
xor U1985 (N_1985,N_1943,N_1928);
xor U1986 (N_1986,N_1919,N_1916);
nand U1987 (N_1987,N_1948,N_1924);
or U1988 (N_1988,N_1902,N_1919);
and U1989 (N_1989,N_1921,N_1934);
nor U1990 (N_1990,N_1903,N_1923);
or U1991 (N_1991,N_1945,N_1924);
nand U1992 (N_1992,N_1913,N_1941);
nor U1993 (N_1993,N_1930,N_1915);
and U1994 (N_1994,N_1941,N_1904);
and U1995 (N_1995,N_1918,N_1921);
and U1996 (N_1996,N_1908,N_1949);
nand U1997 (N_1997,N_1917,N_1924);
nand U1998 (N_1998,N_1936,N_1937);
xnor U1999 (N_1999,N_1949,N_1939);
nand U2000 (N_2000,N_1954,N_1988);
xor U2001 (N_2001,N_1981,N_1969);
or U2002 (N_2002,N_1965,N_1951);
nor U2003 (N_2003,N_1967,N_1953);
or U2004 (N_2004,N_1997,N_1996);
or U2005 (N_2005,N_1963,N_1979);
xnor U2006 (N_2006,N_1957,N_1999);
and U2007 (N_2007,N_1958,N_1959);
nand U2008 (N_2008,N_1960,N_1970);
or U2009 (N_2009,N_1962,N_1993);
nor U2010 (N_2010,N_1987,N_1989);
xor U2011 (N_2011,N_1977,N_1964);
nor U2012 (N_2012,N_1966,N_1950);
xor U2013 (N_2013,N_1983,N_1998);
and U2014 (N_2014,N_1952,N_1994);
or U2015 (N_2015,N_1971,N_1980);
or U2016 (N_2016,N_1995,N_1956);
or U2017 (N_2017,N_1968,N_1961);
nor U2018 (N_2018,N_1986,N_1984);
nor U2019 (N_2019,N_1976,N_1992);
and U2020 (N_2020,N_1973,N_1991);
and U2021 (N_2021,N_1972,N_1955);
or U2022 (N_2022,N_1985,N_1982);
nand U2023 (N_2023,N_1974,N_1990);
nor U2024 (N_2024,N_1978,N_1975);
nor U2025 (N_2025,N_1981,N_1990);
nand U2026 (N_2026,N_1977,N_1952);
or U2027 (N_2027,N_1967,N_1960);
and U2028 (N_2028,N_1962,N_1981);
xnor U2029 (N_2029,N_1987,N_1982);
nand U2030 (N_2030,N_1967,N_1952);
nand U2031 (N_2031,N_1950,N_1964);
nand U2032 (N_2032,N_1983,N_1952);
and U2033 (N_2033,N_1974,N_1999);
nor U2034 (N_2034,N_1994,N_1986);
and U2035 (N_2035,N_1995,N_1982);
nor U2036 (N_2036,N_1958,N_1993);
nor U2037 (N_2037,N_1989,N_1980);
or U2038 (N_2038,N_1996,N_1992);
xor U2039 (N_2039,N_1989,N_1956);
or U2040 (N_2040,N_1965,N_1980);
xor U2041 (N_2041,N_1982,N_1976);
nor U2042 (N_2042,N_1950,N_1959);
nand U2043 (N_2043,N_1955,N_1997);
or U2044 (N_2044,N_1962,N_1983);
nor U2045 (N_2045,N_1950,N_1993);
and U2046 (N_2046,N_1982,N_1979);
or U2047 (N_2047,N_1969,N_1987);
nand U2048 (N_2048,N_1968,N_1993);
xnor U2049 (N_2049,N_1985,N_1975);
nand U2050 (N_2050,N_2033,N_2027);
xor U2051 (N_2051,N_2037,N_2039);
or U2052 (N_2052,N_2019,N_2030);
nor U2053 (N_2053,N_2043,N_2045);
and U2054 (N_2054,N_2014,N_2010);
nor U2055 (N_2055,N_2015,N_2023);
nor U2056 (N_2056,N_2004,N_2029);
xor U2057 (N_2057,N_2002,N_2001);
xnor U2058 (N_2058,N_2042,N_2021);
nor U2059 (N_2059,N_2026,N_2035);
and U2060 (N_2060,N_2000,N_2018);
nand U2061 (N_2061,N_2009,N_2048);
and U2062 (N_2062,N_2016,N_2049);
nand U2063 (N_2063,N_2011,N_2041);
and U2064 (N_2064,N_2046,N_2040);
nand U2065 (N_2065,N_2020,N_2005);
nand U2066 (N_2066,N_2031,N_2022);
xnor U2067 (N_2067,N_2047,N_2017);
and U2068 (N_2068,N_2036,N_2003);
nor U2069 (N_2069,N_2007,N_2013);
and U2070 (N_2070,N_2024,N_2034);
and U2071 (N_2071,N_2032,N_2006);
nor U2072 (N_2072,N_2025,N_2012);
nand U2073 (N_2073,N_2008,N_2038);
and U2074 (N_2074,N_2028,N_2044);
and U2075 (N_2075,N_2047,N_2006);
nor U2076 (N_2076,N_2017,N_2001);
and U2077 (N_2077,N_2045,N_2049);
or U2078 (N_2078,N_2033,N_2047);
nand U2079 (N_2079,N_2014,N_2031);
xnor U2080 (N_2080,N_2027,N_2002);
and U2081 (N_2081,N_2012,N_2030);
and U2082 (N_2082,N_2035,N_2028);
or U2083 (N_2083,N_2032,N_2045);
xor U2084 (N_2084,N_2015,N_2045);
nor U2085 (N_2085,N_2029,N_2002);
nand U2086 (N_2086,N_2029,N_2035);
and U2087 (N_2087,N_2023,N_2009);
or U2088 (N_2088,N_2015,N_2044);
xor U2089 (N_2089,N_2005,N_2048);
or U2090 (N_2090,N_2034,N_2042);
or U2091 (N_2091,N_2030,N_2037);
and U2092 (N_2092,N_2029,N_2022);
nand U2093 (N_2093,N_2004,N_2015);
nand U2094 (N_2094,N_2036,N_2023);
or U2095 (N_2095,N_2003,N_2013);
or U2096 (N_2096,N_2026,N_2016);
and U2097 (N_2097,N_2008,N_2003);
or U2098 (N_2098,N_2029,N_2025);
and U2099 (N_2099,N_2013,N_2024);
and U2100 (N_2100,N_2077,N_2097);
nor U2101 (N_2101,N_2065,N_2085);
nand U2102 (N_2102,N_2060,N_2072);
nor U2103 (N_2103,N_2057,N_2066);
xnor U2104 (N_2104,N_2090,N_2091);
xor U2105 (N_2105,N_2059,N_2099);
or U2106 (N_2106,N_2078,N_2094);
and U2107 (N_2107,N_2075,N_2067);
and U2108 (N_2108,N_2086,N_2088);
nor U2109 (N_2109,N_2058,N_2069);
nor U2110 (N_2110,N_2070,N_2089);
nand U2111 (N_2111,N_2096,N_2083);
xnor U2112 (N_2112,N_2079,N_2084);
and U2113 (N_2113,N_2053,N_2074);
nand U2114 (N_2114,N_2054,N_2076);
xnor U2115 (N_2115,N_2051,N_2071);
nor U2116 (N_2116,N_2082,N_2073);
nor U2117 (N_2117,N_2098,N_2062);
nand U2118 (N_2118,N_2056,N_2064);
nand U2119 (N_2119,N_2095,N_2087);
and U2120 (N_2120,N_2061,N_2050);
and U2121 (N_2121,N_2081,N_2093);
or U2122 (N_2122,N_2063,N_2080);
nor U2123 (N_2123,N_2092,N_2068);
nor U2124 (N_2124,N_2052,N_2055);
xor U2125 (N_2125,N_2057,N_2070);
or U2126 (N_2126,N_2096,N_2071);
nor U2127 (N_2127,N_2080,N_2091);
and U2128 (N_2128,N_2067,N_2079);
or U2129 (N_2129,N_2097,N_2053);
or U2130 (N_2130,N_2074,N_2078);
nor U2131 (N_2131,N_2083,N_2075);
or U2132 (N_2132,N_2054,N_2070);
or U2133 (N_2133,N_2086,N_2050);
or U2134 (N_2134,N_2096,N_2064);
nand U2135 (N_2135,N_2070,N_2065);
and U2136 (N_2136,N_2057,N_2074);
or U2137 (N_2137,N_2091,N_2060);
or U2138 (N_2138,N_2098,N_2086);
and U2139 (N_2139,N_2091,N_2082);
nand U2140 (N_2140,N_2099,N_2070);
and U2141 (N_2141,N_2077,N_2085);
or U2142 (N_2142,N_2090,N_2081);
nor U2143 (N_2143,N_2058,N_2076);
nand U2144 (N_2144,N_2063,N_2067);
nor U2145 (N_2145,N_2062,N_2072);
and U2146 (N_2146,N_2064,N_2068);
xnor U2147 (N_2147,N_2082,N_2062);
nand U2148 (N_2148,N_2069,N_2052);
and U2149 (N_2149,N_2085,N_2087);
xnor U2150 (N_2150,N_2103,N_2144);
and U2151 (N_2151,N_2147,N_2125);
nand U2152 (N_2152,N_2116,N_2124);
xnor U2153 (N_2153,N_2121,N_2130);
xor U2154 (N_2154,N_2104,N_2149);
and U2155 (N_2155,N_2138,N_2117);
nand U2156 (N_2156,N_2133,N_2143);
xnor U2157 (N_2157,N_2119,N_2106);
and U2158 (N_2158,N_2135,N_2123);
nor U2159 (N_2159,N_2141,N_2140);
nand U2160 (N_2160,N_2105,N_2148);
or U2161 (N_2161,N_2131,N_2129);
nand U2162 (N_2162,N_2110,N_2134);
nor U2163 (N_2163,N_2102,N_2137);
nand U2164 (N_2164,N_2142,N_2146);
and U2165 (N_2165,N_2127,N_2126);
nand U2166 (N_2166,N_2101,N_2115);
or U2167 (N_2167,N_2145,N_2118);
xor U2168 (N_2168,N_2132,N_2107);
or U2169 (N_2169,N_2139,N_2120);
or U2170 (N_2170,N_2108,N_2112);
and U2171 (N_2171,N_2122,N_2128);
or U2172 (N_2172,N_2114,N_2100);
and U2173 (N_2173,N_2111,N_2113);
xor U2174 (N_2174,N_2136,N_2109);
or U2175 (N_2175,N_2109,N_2137);
xnor U2176 (N_2176,N_2130,N_2102);
and U2177 (N_2177,N_2105,N_2147);
and U2178 (N_2178,N_2128,N_2141);
and U2179 (N_2179,N_2141,N_2146);
and U2180 (N_2180,N_2114,N_2137);
and U2181 (N_2181,N_2145,N_2138);
nor U2182 (N_2182,N_2104,N_2147);
xor U2183 (N_2183,N_2147,N_2138);
xor U2184 (N_2184,N_2125,N_2144);
and U2185 (N_2185,N_2109,N_2135);
nor U2186 (N_2186,N_2146,N_2107);
and U2187 (N_2187,N_2146,N_2135);
or U2188 (N_2188,N_2111,N_2102);
nand U2189 (N_2189,N_2133,N_2106);
or U2190 (N_2190,N_2100,N_2144);
xor U2191 (N_2191,N_2122,N_2102);
nor U2192 (N_2192,N_2148,N_2137);
or U2193 (N_2193,N_2140,N_2117);
or U2194 (N_2194,N_2125,N_2108);
xor U2195 (N_2195,N_2137,N_2120);
or U2196 (N_2196,N_2120,N_2103);
or U2197 (N_2197,N_2137,N_2144);
xnor U2198 (N_2198,N_2138,N_2132);
xnor U2199 (N_2199,N_2135,N_2107);
xor U2200 (N_2200,N_2190,N_2153);
nor U2201 (N_2201,N_2170,N_2171);
or U2202 (N_2202,N_2186,N_2160);
and U2203 (N_2203,N_2163,N_2173);
or U2204 (N_2204,N_2187,N_2151);
nor U2205 (N_2205,N_2162,N_2150);
xor U2206 (N_2206,N_2152,N_2158);
nor U2207 (N_2207,N_2183,N_2178);
or U2208 (N_2208,N_2175,N_2155);
and U2209 (N_2209,N_2188,N_2189);
and U2210 (N_2210,N_2197,N_2196);
nand U2211 (N_2211,N_2182,N_2180);
nand U2212 (N_2212,N_2185,N_2159);
and U2213 (N_2213,N_2156,N_2154);
and U2214 (N_2214,N_2172,N_2192);
nor U2215 (N_2215,N_2195,N_2174);
nor U2216 (N_2216,N_2191,N_2199);
and U2217 (N_2217,N_2198,N_2164);
or U2218 (N_2218,N_2168,N_2193);
xor U2219 (N_2219,N_2169,N_2166);
nand U2220 (N_2220,N_2184,N_2167);
nor U2221 (N_2221,N_2194,N_2177);
nand U2222 (N_2222,N_2165,N_2161);
or U2223 (N_2223,N_2157,N_2179);
or U2224 (N_2224,N_2176,N_2181);
nor U2225 (N_2225,N_2187,N_2171);
or U2226 (N_2226,N_2164,N_2160);
nand U2227 (N_2227,N_2193,N_2189);
or U2228 (N_2228,N_2183,N_2156);
nand U2229 (N_2229,N_2177,N_2190);
nand U2230 (N_2230,N_2185,N_2164);
nor U2231 (N_2231,N_2187,N_2196);
or U2232 (N_2232,N_2175,N_2178);
nor U2233 (N_2233,N_2170,N_2150);
or U2234 (N_2234,N_2198,N_2167);
or U2235 (N_2235,N_2185,N_2184);
and U2236 (N_2236,N_2153,N_2184);
or U2237 (N_2237,N_2197,N_2176);
nand U2238 (N_2238,N_2150,N_2175);
and U2239 (N_2239,N_2189,N_2166);
or U2240 (N_2240,N_2158,N_2151);
nand U2241 (N_2241,N_2186,N_2151);
nand U2242 (N_2242,N_2177,N_2191);
nor U2243 (N_2243,N_2167,N_2187);
and U2244 (N_2244,N_2159,N_2151);
nand U2245 (N_2245,N_2174,N_2170);
and U2246 (N_2246,N_2155,N_2152);
nand U2247 (N_2247,N_2185,N_2172);
nor U2248 (N_2248,N_2178,N_2156);
xnor U2249 (N_2249,N_2170,N_2163);
nand U2250 (N_2250,N_2206,N_2229);
or U2251 (N_2251,N_2207,N_2245);
and U2252 (N_2252,N_2228,N_2230);
nand U2253 (N_2253,N_2232,N_2202);
xnor U2254 (N_2254,N_2219,N_2223);
and U2255 (N_2255,N_2201,N_2234);
or U2256 (N_2256,N_2213,N_2209);
and U2257 (N_2257,N_2248,N_2220);
xnor U2258 (N_2258,N_2214,N_2227);
nor U2259 (N_2259,N_2246,N_2217);
xnor U2260 (N_2260,N_2205,N_2221);
or U2261 (N_2261,N_2231,N_2236);
and U2262 (N_2262,N_2233,N_2226);
nor U2263 (N_2263,N_2240,N_2211);
nor U2264 (N_2264,N_2204,N_2215);
nand U2265 (N_2265,N_2249,N_2244);
and U2266 (N_2266,N_2239,N_2210);
nor U2267 (N_2267,N_2212,N_2247);
nand U2268 (N_2268,N_2243,N_2235);
xor U2269 (N_2269,N_2218,N_2224);
xnor U2270 (N_2270,N_2241,N_2208);
and U2271 (N_2271,N_2238,N_2216);
nand U2272 (N_2272,N_2200,N_2242);
xnor U2273 (N_2273,N_2237,N_2203);
or U2274 (N_2274,N_2225,N_2222);
or U2275 (N_2275,N_2230,N_2205);
nor U2276 (N_2276,N_2209,N_2227);
nand U2277 (N_2277,N_2237,N_2209);
nor U2278 (N_2278,N_2217,N_2242);
and U2279 (N_2279,N_2240,N_2224);
nand U2280 (N_2280,N_2201,N_2204);
xnor U2281 (N_2281,N_2236,N_2245);
and U2282 (N_2282,N_2231,N_2221);
and U2283 (N_2283,N_2215,N_2229);
nand U2284 (N_2284,N_2210,N_2245);
and U2285 (N_2285,N_2248,N_2243);
nand U2286 (N_2286,N_2208,N_2244);
or U2287 (N_2287,N_2200,N_2205);
xor U2288 (N_2288,N_2238,N_2245);
xor U2289 (N_2289,N_2243,N_2200);
nor U2290 (N_2290,N_2225,N_2202);
xnor U2291 (N_2291,N_2233,N_2215);
or U2292 (N_2292,N_2219,N_2215);
xor U2293 (N_2293,N_2248,N_2229);
and U2294 (N_2294,N_2233,N_2220);
or U2295 (N_2295,N_2243,N_2205);
nor U2296 (N_2296,N_2204,N_2213);
nand U2297 (N_2297,N_2223,N_2203);
xnor U2298 (N_2298,N_2218,N_2201);
xor U2299 (N_2299,N_2247,N_2213);
and U2300 (N_2300,N_2298,N_2287);
nor U2301 (N_2301,N_2256,N_2260);
and U2302 (N_2302,N_2289,N_2279);
or U2303 (N_2303,N_2286,N_2283);
nand U2304 (N_2304,N_2295,N_2250);
nor U2305 (N_2305,N_2296,N_2293);
or U2306 (N_2306,N_2292,N_2266);
nor U2307 (N_2307,N_2277,N_2278);
nor U2308 (N_2308,N_2263,N_2294);
or U2309 (N_2309,N_2270,N_2259);
and U2310 (N_2310,N_2261,N_2276);
xnor U2311 (N_2311,N_2258,N_2274);
xnor U2312 (N_2312,N_2269,N_2257);
or U2313 (N_2313,N_2281,N_2297);
nand U2314 (N_2314,N_2267,N_2271);
nor U2315 (N_2315,N_2288,N_2262);
and U2316 (N_2316,N_2251,N_2268);
or U2317 (N_2317,N_2290,N_2252);
or U2318 (N_2318,N_2282,N_2299);
and U2319 (N_2319,N_2284,N_2275);
xor U2320 (N_2320,N_2285,N_2255);
xor U2321 (N_2321,N_2273,N_2254);
or U2322 (N_2322,N_2253,N_2264);
xor U2323 (N_2323,N_2280,N_2291);
nor U2324 (N_2324,N_2265,N_2272);
xnor U2325 (N_2325,N_2255,N_2297);
or U2326 (N_2326,N_2252,N_2276);
nor U2327 (N_2327,N_2273,N_2270);
nand U2328 (N_2328,N_2273,N_2255);
nor U2329 (N_2329,N_2299,N_2280);
xor U2330 (N_2330,N_2270,N_2269);
nor U2331 (N_2331,N_2255,N_2265);
and U2332 (N_2332,N_2279,N_2259);
xnor U2333 (N_2333,N_2287,N_2253);
or U2334 (N_2334,N_2267,N_2299);
nand U2335 (N_2335,N_2269,N_2292);
nor U2336 (N_2336,N_2270,N_2257);
nand U2337 (N_2337,N_2285,N_2259);
or U2338 (N_2338,N_2272,N_2281);
or U2339 (N_2339,N_2294,N_2299);
xnor U2340 (N_2340,N_2299,N_2293);
xor U2341 (N_2341,N_2263,N_2295);
and U2342 (N_2342,N_2283,N_2260);
nor U2343 (N_2343,N_2257,N_2278);
xor U2344 (N_2344,N_2250,N_2251);
and U2345 (N_2345,N_2290,N_2287);
xnor U2346 (N_2346,N_2281,N_2285);
and U2347 (N_2347,N_2252,N_2274);
nand U2348 (N_2348,N_2261,N_2267);
nor U2349 (N_2349,N_2288,N_2255);
nor U2350 (N_2350,N_2309,N_2347);
and U2351 (N_2351,N_2313,N_2300);
nor U2352 (N_2352,N_2308,N_2312);
and U2353 (N_2353,N_2340,N_2306);
nand U2354 (N_2354,N_2330,N_2319);
and U2355 (N_2355,N_2327,N_2314);
and U2356 (N_2356,N_2325,N_2332);
and U2357 (N_2357,N_2348,N_2318);
nand U2358 (N_2358,N_2329,N_2321);
nor U2359 (N_2359,N_2307,N_2320);
or U2360 (N_2360,N_2328,N_2337);
or U2361 (N_2361,N_2342,N_2317);
or U2362 (N_2362,N_2304,N_2315);
xnor U2363 (N_2363,N_2335,N_2333);
nor U2364 (N_2364,N_2341,N_2331);
and U2365 (N_2365,N_2326,N_2345);
or U2366 (N_2366,N_2343,N_2316);
and U2367 (N_2367,N_2310,N_2349);
xnor U2368 (N_2368,N_2338,N_2305);
nand U2369 (N_2369,N_2323,N_2303);
and U2370 (N_2370,N_2311,N_2301);
xnor U2371 (N_2371,N_2322,N_2339);
nor U2372 (N_2372,N_2344,N_2324);
nand U2373 (N_2373,N_2336,N_2346);
nand U2374 (N_2374,N_2302,N_2334);
and U2375 (N_2375,N_2309,N_2318);
or U2376 (N_2376,N_2320,N_2331);
xor U2377 (N_2377,N_2339,N_2325);
xor U2378 (N_2378,N_2300,N_2344);
and U2379 (N_2379,N_2318,N_2316);
nand U2380 (N_2380,N_2339,N_2303);
nand U2381 (N_2381,N_2328,N_2326);
xor U2382 (N_2382,N_2314,N_2341);
nand U2383 (N_2383,N_2345,N_2314);
or U2384 (N_2384,N_2315,N_2302);
and U2385 (N_2385,N_2344,N_2338);
and U2386 (N_2386,N_2316,N_2325);
nand U2387 (N_2387,N_2334,N_2348);
nand U2388 (N_2388,N_2312,N_2302);
and U2389 (N_2389,N_2310,N_2320);
nand U2390 (N_2390,N_2338,N_2334);
nand U2391 (N_2391,N_2346,N_2304);
or U2392 (N_2392,N_2341,N_2343);
xor U2393 (N_2393,N_2336,N_2318);
and U2394 (N_2394,N_2336,N_2303);
xnor U2395 (N_2395,N_2327,N_2319);
xor U2396 (N_2396,N_2314,N_2331);
nor U2397 (N_2397,N_2314,N_2308);
or U2398 (N_2398,N_2303,N_2319);
nand U2399 (N_2399,N_2322,N_2326);
or U2400 (N_2400,N_2393,N_2373);
xor U2401 (N_2401,N_2356,N_2369);
or U2402 (N_2402,N_2350,N_2382);
nand U2403 (N_2403,N_2392,N_2379);
nor U2404 (N_2404,N_2398,N_2381);
and U2405 (N_2405,N_2357,N_2386);
nand U2406 (N_2406,N_2395,N_2388);
xnor U2407 (N_2407,N_2399,N_2397);
or U2408 (N_2408,N_2367,N_2362);
and U2409 (N_2409,N_2363,N_2387);
xnor U2410 (N_2410,N_2378,N_2366);
xor U2411 (N_2411,N_2361,N_2385);
nand U2412 (N_2412,N_2370,N_2355);
and U2413 (N_2413,N_2390,N_2377);
nand U2414 (N_2414,N_2380,N_2396);
nand U2415 (N_2415,N_2359,N_2394);
xor U2416 (N_2416,N_2372,N_2354);
or U2417 (N_2417,N_2389,N_2371);
and U2418 (N_2418,N_2368,N_2383);
nor U2419 (N_2419,N_2374,N_2358);
xor U2420 (N_2420,N_2376,N_2360);
and U2421 (N_2421,N_2352,N_2384);
nor U2422 (N_2422,N_2351,N_2365);
nor U2423 (N_2423,N_2353,N_2375);
or U2424 (N_2424,N_2391,N_2364);
and U2425 (N_2425,N_2356,N_2354);
or U2426 (N_2426,N_2368,N_2387);
nand U2427 (N_2427,N_2399,N_2395);
and U2428 (N_2428,N_2368,N_2384);
or U2429 (N_2429,N_2355,N_2378);
nor U2430 (N_2430,N_2382,N_2361);
or U2431 (N_2431,N_2396,N_2382);
nand U2432 (N_2432,N_2360,N_2370);
nor U2433 (N_2433,N_2373,N_2360);
xnor U2434 (N_2434,N_2388,N_2357);
xnor U2435 (N_2435,N_2359,N_2382);
and U2436 (N_2436,N_2351,N_2367);
or U2437 (N_2437,N_2356,N_2374);
and U2438 (N_2438,N_2363,N_2377);
nand U2439 (N_2439,N_2374,N_2384);
nand U2440 (N_2440,N_2380,N_2367);
nand U2441 (N_2441,N_2394,N_2350);
and U2442 (N_2442,N_2373,N_2353);
xnor U2443 (N_2443,N_2360,N_2397);
and U2444 (N_2444,N_2366,N_2399);
xor U2445 (N_2445,N_2379,N_2381);
or U2446 (N_2446,N_2390,N_2372);
nor U2447 (N_2447,N_2357,N_2395);
nand U2448 (N_2448,N_2364,N_2363);
or U2449 (N_2449,N_2381,N_2392);
and U2450 (N_2450,N_2409,N_2443);
xor U2451 (N_2451,N_2427,N_2406);
nand U2452 (N_2452,N_2436,N_2435);
xor U2453 (N_2453,N_2417,N_2440);
nor U2454 (N_2454,N_2416,N_2400);
xnor U2455 (N_2455,N_2410,N_2424);
or U2456 (N_2456,N_2448,N_2432);
xor U2457 (N_2457,N_2428,N_2423);
or U2458 (N_2458,N_2439,N_2426);
xor U2459 (N_2459,N_2444,N_2438);
and U2460 (N_2460,N_2407,N_2422);
xnor U2461 (N_2461,N_2429,N_2405);
nor U2462 (N_2462,N_2420,N_2442);
xnor U2463 (N_2463,N_2414,N_2412);
xor U2464 (N_2464,N_2431,N_2446);
xor U2465 (N_2465,N_2445,N_2401);
xor U2466 (N_2466,N_2425,N_2408);
nor U2467 (N_2467,N_2418,N_2411);
nor U2468 (N_2468,N_2415,N_2447);
nor U2469 (N_2469,N_2421,N_2403);
nand U2470 (N_2470,N_2430,N_2404);
nor U2471 (N_2471,N_2437,N_2402);
or U2472 (N_2472,N_2433,N_2449);
nand U2473 (N_2473,N_2441,N_2419);
and U2474 (N_2474,N_2413,N_2434);
and U2475 (N_2475,N_2441,N_2403);
nand U2476 (N_2476,N_2420,N_2400);
xor U2477 (N_2477,N_2415,N_2443);
and U2478 (N_2478,N_2420,N_2436);
nand U2479 (N_2479,N_2413,N_2439);
and U2480 (N_2480,N_2413,N_2425);
nand U2481 (N_2481,N_2414,N_2407);
nor U2482 (N_2482,N_2436,N_2447);
nor U2483 (N_2483,N_2428,N_2401);
nand U2484 (N_2484,N_2435,N_2402);
nand U2485 (N_2485,N_2416,N_2414);
nand U2486 (N_2486,N_2424,N_2426);
nand U2487 (N_2487,N_2437,N_2409);
nor U2488 (N_2488,N_2444,N_2403);
and U2489 (N_2489,N_2447,N_2409);
and U2490 (N_2490,N_2449,N_2415);
nor U2491 (N_2491,N_2435,N_2440);
nor U2492 (N_2492,N_2417,N_2402);
xor U2493 (N_2493,N_2406,N_2408);
and U2494 (N_2494,N_2441,N_2411);
or U2495 (N_2495,N_2425,N_2411);
and U2496 (N_2496,N_2413,N_2436);
xnor U2497 (N_2497,N_2418,N_2413);
or U2498 (N_2498,N_2411,N_2433);
nor U2499 (N_2499,N_2416,N_2447);
nand U2500 (N_2500,N_2470,N_2488);
and U2501 (N_2501,N_2475,N_2495);
xnor U2502 (N_2502,N_2476,N_2450);
and U2503 (N_2503,N_2451,N_2494);
nand U2504 (N_2504,N_2474,N_2453);
nor U2505 (N_2505,N_2480,N_2479);
xnor U2506 (N_2506,N_2460,N_2484);
xnor U2507 (N_2507,N_2499,N_2492);
and U2508 (N_2508,N_2471,N_2483);
xnor U2509 (N_2509,N_2489,N_2461);
xor U2510 (N_2510,N_2459,N_2491);
or U2511 (N_2511,N_2472,N_2467);
and U2512 (N_2512,N_2463,N_2462);
xnor U2513 (N_2513,N_2498,N_2493);
xor U2514 (N_2514,N_2487,N_2466);
or U2515 (N_2515,N_2456,N_2469);
xnor U2516 (N_2516,N_2482,N_2478);
and U2517 (N_2517,N_2486,N_2457);
xnor U2518 (N_2518,N_2455,N_2458);
nor U2519 (N_2519,N_2477,N_2465);
nor U2520 (N_2520,N_2490,N_2452);
nor U2521 (N_2521,N_2497,N_2485);
and U2522 (N_2522,N_2468,N_2481);
or U2523 (N_2523,N_2464,N_2454);
or U2524 (N_2524,N_2473,N_2496);
xnor U2525 (N_2525,N_2464,N_2467);
nor U2526 (N_2526,N_2459,N_2468);
or U2527 (N_2527,N_2478,N_2451);
and U2528 (N_2528,N_2467,N_2484);
and U2529 (N_2529,N_2479,N_2491);
nor U2530 (N_2530,N_2479,N_2463);
nor U2531 (N_2531,N_2470,N_2454);
nor U2532 (N_2532,N_2490,N_2478);
nand U2533 (N_2533,N_2468,N_2491);
or U2534 (N_2534,N_2472,N_2461);
or U2535 (N_2535,N_2479,N_2473);
xor U2536 (N_2536,N_2457,N_2471);
or U2537 (N_2537,N_2488,N_2450);
or U2538 (N_2538,N_2463,N_2458);
xnor U2539 (N_2539,N_2458,N_2496);
xor U2540 (N_2540,N_2452,N_2453);
nand U2541 (N_2541,N_2453,N_2486);
or U2542 (N_2542,N_2492,N_2464);
xnor U2543 (N_2543,N_2479,N_2472);
xnor U2544 (N_2544,N_2468,N_2473);
or U2545 (N_2545,N_2453,N_2467);
nand U2546 (N_2546,N_2475,N_2485);
or U2547 (N_2547,N_2481,N_2469);
and U2548 (N_2548,N_2470,N_2474);
nand U2549 (N_2549,N_2468,N_2484);
xnor U2550 (N_2550,N_2546,N_2540);
and U2551 (N_2551,N_2514,N_2519);
nor U2552 (N_2552,N_2516,N_2545);
and U2553 (N_2553,N_2511,N_2505);
xor U2554 (N_2554,N_2500,N_2523);
nor U2555 (N_2555,N_2528,N_2508);
nand U2556 (N_2556,N_2534,N_2547);
and U2557 (N_2557,N_2507,N_2529);
or U2558 (N_2558,N_2539,N_2522);
and U2559 (N_2559,N_2544,N_2521);
nor U2560 (N_2560,N_2506,N_2509);
nor U2561 (N_2561,N_2533,N_2517);
nand U2562 (N_2562,N_2531,N_2543);
nor U2563 (N_2563,N_2515,N_2548);
nand U2564 (N_2564,N_2518,N_2532);
nand U2565 (N_2565,N_2525,N_2549);
and U2566 (N_2566,N_2527,N_2501);
nand U2567 (N_2567,N_2542,N_2512);
or U2568 (N_2568,N_2510,N_2524);
nor U2569 (N_2569,N_2537,N_2503);
and U2570 (N_2570,N_2504,N_2513);
xor U2571 (N_2571,N_2536,N_2541);
xor U2572 (N_2572,N_2502,N_2530);
and U2573 (N_2573,N_2538,N_2520);
or U2574 (N_2574,N_2526,N_2535);
nor U2575 (N_2575,N_2540,N_2503);
xor U2576 (N_2576,N_2527,N_2542);
and U2577 (N_2577,N_2529,N_2535);
nor U2578 (N_2578,N_2500,N_2508);
and U2579 (N_2579,N_2545,N_2544);
nand U2580 (N_2580,N_2534,N_2511);
or U2581 (N_2581,N_2519,N_2513);
nor U2582 (N_2582,N_2512,N_2546);
xor U2583 (N_2583,N_2518,N_2519);
or U2584 (N_2584,N_2518,N_2540);
nand U2585 (N_2585,N_2547,N_2524);
nand U2586 (N_2586,N_2536,N_2535);
or U2587 (N_2587,N_2533,N_2519);
nand U2588 (N_2588,N_2506,N_2541);
nor U2589 (N_2589,N_2519,N_2547);
and U2590 (N_2590,N_2548,N_2509);
xor U2591 (N_2591,N_2515,N_2509);
nand U2592 (N_2592,N_2514,N_2526);
nor U2593 (N_2593,N_2517,N_2544);
nor U2594 (N_2594,N_2528,N_2513);
or U2595 (N_2595,N_2539,N_2508);
nor U2596 (N_2596,N_2523,N_2525);
or U2597 (N_2597,N_2535,N_2541);
and U2598 (N_2598,N_2536,N_2503);
and U2599 (N_2599,N_2513,N_2523);
and U2600 (N_2600,N_2591,N_2553);
nand U2601 (N_2601,N_2563,N_2586);
nor U2602 (N_2602,N_2577,N_2580);
nor U2603 (N_2603,N_2598,N_2566);
nand U2604 (N_2604,N_2588,N_2575);
and U2605 (N_2605,N_2555,N_2557);
xnor U2606 (N_2606,N_2550,N_2574);
xor U2607 (N_2607,N_2571,N_2560);
and U2608 (N_2608,N_2579,N_2583);
nand U2609 (N_2609,N_2594,N_2585);
and U2610 (N_2610,N_2568,N_2567);
and U2611 (N_2611,N_2593,N_2552);
nand U2612 (N_2612,N_2558,N_2584);
and U2613 (N_2613,N_2569,N_2581);
xnor U2614 (N_2614,N_2582,N_2578);
nand U2615 (N_2615,N_2564,N_2597);
nor U2616 (N_2616,N_2561,N_2590);
or U2617 (N_2617,N_2551,N_2570);
and U2618 (N_2618,N_2576,N_2572);
xor U2619 (N_2619,N_2565,N_2562);
nand U2620 (N_2620,N_2596,N_2556);
and U2621 (N_2621,N_2559,N_2589);
nor U2622 (N_2622,N_2592,N_2599);
nand U2623 (N_2623,N_2587,N_2554);
nand U2624 (N_2624,N_2573,N_2595);
and U2625 (N_2625,N_2571,N_2561);
nor U2626 (N_2626,N_2564,N_2585);
or U2627 (N_2627,N_2572,N_2597);
or U2628 (N_2628,N_2587,N_2569);
xor U2629 (N_2629,N_2591,N_2566);
nor U2630 (N_2630,N_2552,N_2550);
nand U2631 (N_2631,N_2592,N_2573);
nor U2632 (N_2632,N_2583,N_2587);
and U2633 (N_2633,N_2582,N_2584);
xnor U2634 (N_2634,N_2574,N_2556);
nor U2635 (N_2635,N_2593,N_2594);
nor U2636 (N_2636,N_2560,N_2586);
or U2637 (N_2637,N_2591,N_2590);
nand U2638 (N_2638,N_2598,N_2561);
and U2639 (N_2639,N_2571,N_2576);
and U2640 (N_2640,N_2570,N_2565);
or U2641 (N_2641,N_2551,N_2557);
or U2642 (N_2642,N_2579,N_2576);
xnor U2643 (N_2643,N_2588,N_2550);
nand U2644 (N_2644,N_2588,N_2591);
nand U2645 (N_2645,N_2566,N_2579);
and U2646 (N_2646,N_2565,N_2595);
nand U2647 (N_2647,N_2593,N_2595);
xnor U2648 (N_2648,N_2570,N_2566);
nand U2649 (N_2649,N_2551,N_2599);
xor U2650 (N_2650,N_2638,N_2649);
nor U2651 (N_2651,N_2603,N_2648);
nand U2652 (N_2652,N_2639,N_2613);
nand U2653 (N_2653,N_2609,N_2614);
and U2654 (N_2654,N_2635,N_2645);
and U2655 (N_2655,N_2637,N_2640);
and U2656 (N_2656,N_2643,N_2610);
nor U2657 (N_2657,N_2602,N_2620);
xor U2658 (N_2658,N_2644,N_2624);
nand U2659 (N_2659,N_2629,N_2616);
nand U2660 (N_2660,N_2636,N_2606);
xnor U2661 (N_2661,N_2622,N_2612);
nor U2662 (N_2662,N_2621,N_2605);
xor U2663 (N_2663,N_2607,N_2601);
nor U2664 (N_2664,N_2600,N_2632);
nand U2665 (N_2665,N_2631,N_2626);
nand U2666 (N_2666,N_2634,N_2625);
or U2667 (N_2667,N_2619,N_2628);
xor U2668 (N_2668,N_2633,N_2623);
nor U2669 (N_2669,N_2627,N_2641);
or U2670 (N_2670,N_2642,N_2647);
nor U2671 (N_2671,N_2604,N_2646);
nand U2672 (N_2672,N_2615,N_2611);
and U2673 (N_2673,N_2608,N_2618);
nand U2674 (N_2674,N_2630,N_2617);
xor U2675 (N_2675,N_2625,N_2619);
nand U2676 (N_2676,N_2645,N_2644);
or U2677 (N_2677,N_2603,N_2632);
nand U2678 (N_2678,N_2641,N_2605);
nor U2679 (N_2679,N_2611,N_2647);
and U2680 (N_2680,N_2640,N_2615);
xor U2681 (N_2681,N_2638,N_2601);
and U2682 (N_2682,N_2618,N_2606);
xor U2683 (N_2683,N_2616,N_2640);
nand U2684 (N_2684,N_2612,N_2621);
or U2685 (N_2685,N_2635,N_2611);
or U2686 (N_2686,N_2604,N_2627);
or U2687 (N_2687,N_2602,N_2633);
nor U2688 (N_2688,N_2636,N_2624);
xor U2689 (N_2689,N_2604,N_2602);
xnor U2690 (N_2690,N_2624,N_2603);
or U2691 (N_2691,N_2622,N_2621);
nor U2692 (N_2692,N_2644,N_2646);
xnor U2693 (N_2693,N_2612,N_2609);
nor U2694 (N_2694,N_2618,N_2625);
nand U2695 (N_2695,N_2642,N_2638);
nand U2696 (N_2696,N_2608,N_2641);
and U2697 (N_2697,N_2601,N_2600);
xor U2698 (N_2698,N_2600,N_2648);
nor U2699 (N_2699,N_2625,N_2649);
nand U2700 (N_2700,N_2684,N_2683);
xnor U2701 (N_2701,N_2693,N_2658);
xnor U2702 (N_2702,N_2682,N_2677);
nand U2703 (N_2703,N_2664,N_2671);
or U2704 (N_2704,N_2679,N_2662);
or U2705 (N_2705,N_2687,N_2661);
nand U2706 (N_2706,N_2694,N_2685);
and U2707 (N_2707,N_2665,N_2695);
nor U2708 (N_2708,N_2681,N_2651);
and U2709 (N_2709,N_2678,N_2655);
nand U2710 (N_2710,N_2650,N_2689);
or U2711 (N_2711,N_2669,N_2668);
or U2712 (N_2712,N_2653,N_2699);
nor U2713 (N_2713,N_2672,N_2663);
nor U2714 (N_2714,N_2675,N_2652);
nand U2715 (N_2715,N_2692,N_2659);
and U2716 (N_2716,N_2670,N_2698);
and U2717 (N_2717,N_2676,N_2667);
or U2718 (N_2718,N_2686,N_2660);
or U2719 (N_2719,N_2654,N_2674);
xor U2720 (N_2720,N_2680,N_2688);
nor U2721 (N_2721,N_2673,N_2666);
nand U2722 (N_2722,N_2696,N_2697);
or U2723 (N_2723,N_2690,N_2656);
nor U2724 (N_2724,N_2691,N_2657);
xor U2725 (N_2725,N_2683,N_2663);
nand U2726 (N_2726,N_2659,N_2696);
nor U2727 (N_2727,N_2651,N_2684);
or U2728 (N_2728,N_2658,N_2699);
nand U2729 (N_2729,N_2672,N_2666);
or U2730 (N_2730,N_2699,N_2670);
xor U2731 (N_2731,N_2675,N_2660);
nor U2732 (N_2732,N_2687,N_2685);
nor U2733 (N_2733,N_2698,N_2655);
and U2734 (N_2734,N_2672,N_2674);
or U2735 (N_2735,N_2693,N_2666);
xor U2736 (N_2736,N_2690,N_2659);
and U2737 (N_2737,N_2661,N_2669);
or U2738 (N_2738,N_2691,N_2695);
or U2739 (N_2739,N_2664,N_2690);
nand U2740 (N_2740,N_2669,N_2656);
or U2741 (N_2741,N_2693,N_2671);
xor U2742 (N_2742,N_2694,N_2690);
nand U2743 (N_2743,N_2674,N_2682);
and U2744 (N_2744,N_2696,N_2669);
xor U2745 (N_2745,N_2656,N_2697);
nand U2746 (N_2746,N_2654,N_2692);
nand U2747 (N_2747,N_2655,N_2657);
nor U2748 (N_2748,N_2658,N_2660);
nand U2749 (N_2749,N_2681,N_2678);
and U2750 (N_2750,N_2744,N_2741);
and U2751 (N_2751,N_2743,N_2700);
xnor U2752 (N_2752,N_2731,N_2727);
or U2753 (N_2753,N_2715,N_2720);
nor U2754 (N_2754,N_2749,N_2717);
nand U2755 (N_2755,N_2746,N_2738);
or U2756 (N_2756,N_2724,N_2708);
or U2757 (N_2757,N_2748,N_2710);
nor U2758 (N_2758,N_2711,N_2712);
nor U2759 (N_2759,N_2734,N_2736);
nand U2760 (N_2760,N_2713,N_2709);
nor U2761 (N_2761,N_2730,N_2725);
nand U2762 (N_2762,N_2723,N_2716);
xnor U2763 (N_2763,N_2722,N_2718);
xor U2764 (N_2764,N_2728,N_2735);
xor U2765 (N_2765,N_2703,N_2707);
nor U2766 (N_2766,N_2747,N_2706);
xor U2767 (N_2767,N_2739,N_2737);
and U2768 (N_2768,N_2726,N_2714);
xor U2769 (N_2769,N_2729,N_2733);
and U2770 (N_2770,N_2704,N_2719);
and U2771 (N_2771,N_2732,N_2740);
nand U2772 (N_2772,N_2721,N_2745);
and U2773 (N_2773,N_2702,N_2701);
xor U2774 (N_2774,N_2742,N_2705);
and U2775 (N_2775,N_2726,N_2744);
nor U2776 (N_2776,N_2714,N_2723);
xnor U2777 (N_2777,N_2725,N_2721);
xor U2778 (N_2778,N_2716,N_2725);
and U2779 (N_2779,N_2726,N_2725);
or U2780 (N_2780,N_2746,N_2721);
or U2781 (N_2781,N_2714,N_2707);
nand U2782 (N_2782,N_2717,N_2703);
nor U2783 (N_2783,N_2748,N_2714);
and U2784 (N_2784,N_2718,N_2746);
nand U2785 (N_2785,N_2712,N_2715);
nor U2786 (N_2786,N_2731,N_2729);
nor U2787 (N_2787,N_2734,N_2717);
nor U2788 (N_2788,N_2715,N_2740);
xor U2789 (N_2789,N_2724,N_2741);
nand U2790 (N_2790,N_2724,N_2731);
nor U2791 (N_2791,N_2729,N_2726);
or U2792 (N_2792,N_2734,N_2729);
and U2793 (N_2793,N_2722,N_2717);
nor U2794 (N_2794,N_2739,N_2725);
and U2795 (N_2795,N_2737,N_2700);
nand U2796 (N_2796,N_2744,N_2708);
or U2797 (N_2797,N_2723,N_2743);
nor U2798 (N_2798,N_2703,N_2721);
nor U2799 (N_2799,N_2708,N_2715);
nor U2800 (N_2800,N_2795,N_2799);
xnor U2801 (N_2801,N_2770,N_2787);
and U2802 (N_2802,N_2750,N_2767);
xor U2803 (N_2803,N_2793,N_2792);
xor U2804 (N_2804,N_2754,N_2789);
xnor U2805 (N_2805,N_2785,N_2772);
xor U2806 (N_2806,N_2762,N_2755);
and U2807 (N_2807,N_2760,N_2759);
nor U2808 (N_2808,N_2794,N_2781);
nor U2809 (N_2809,N_2782,N_2776);
or U2810 (N_2810,N_2774,N_2768);
xnor U2811 (N_2811,N_2778,N_2753);
or U2812 (N_2812,N_2779,N_2783);
nor U2813 (N_2813,N_2758,N_2786);
or U2814 (N_2814,N_2784,N_2764);
or U2815 (N_2815,N_2751,N_2791);
or U2816 (N_2816,N_2788,N_2766);
nor U2817 (N_2817,N_2752,N_2777);
nand U2818 (N_2818,N_2775,N_2780);
xor U2819 (N_2819,N_2796,N_2790);
and U2820 (N_2820,N_2769,N_2765);
xnor U2821 (N_2821,N_2773,N_2797);
nand U2822 (N_2822,N_2798,N_2757);
or U2823 (N_2823,N_2761,N_2771);
nor U2824 (N_2824,N_2756,N_2763);
or U2825 (N_2825,N_2772,N_2798);
or U2826 (N_2826,N_2760,N_2779);
xor U2827 (N_2827,N_2793,N_2798);
xor U2828 (N_2828,N_2787,N_2784);
xor U2829 (N_2829,N_2791,N_2769);
or U2830 (N_2830,N_2793,N_2761);
xnor U2831 (N_2831,N_2763,N_2791);
and U2832 (N_2832,N_2770,N_2798);
and U2833 (N_2833,N_2794,N_2783);
and U2834 (N_2834,N_2751,N_2797);
xnor U2835 (N_2835,N_2774,N_2783);
or U2836 (N_2836,N_2769,N_2757);
nand U2837 (N_2837,N_2761,N_2775);
and U2838 (N_2838,N_2773,N_2782);
nor U2839 (N_2839,N_2777,N_2754);
nand U2840 (N_2840,N_2758,N_2785);
or U2841 (N_2841,N_2795,N_2798);
or U2842 (N_2842,N_2772,N_2773);
xnor U2843 (N_2843,N_2796,N_2795);
and U2844 (N_2844,N_2792,N_2779);
or U2845 (N_2845,N_2794,N_2779);
nor U2846 (N_2846,N_2772,N_2780);
nor U2847 (N_2847,N_2753,N_2750);
or U2848 (N_2848,N_2780,N_2791);
and U2849 (N_2849,N_2784,N_2791);
or U2850 (N_2850,N_2821,N_2819);
or U2851 (N_2851,N_2846,N_2822);
xor U2852 (N_2852,N_2829,N_2804);
xnor U2853 (N_2853,N_2832,N_2815);
or U2854 (N_2854,N_2849,N_2810);
and U2855 (N_2855,N_2820,N_2801);
and U2856 (N_2856,N_2807,N_2828);
and U2857 (N_2857,N_2808,N_2812);
xnor U2858 (N_2858,N_2838,N_2813);
or U2859 (N_2859,N_2827,N_2818);
nor U2860 (N_2860,N_2826,N_2842);
nand U2861 (N_2861,N_2803,N_2847);
xnor U2862 (N_2862,N_2830,N_2848);
nor U2863 (N_2863,N_2840,N_2844);
nor U2864 (N_2864,N_2823,N_2843);
xnor U2865 (N_2865,N_2835,N_2809);
nand U2866 (N_2866,N_2805,N_2837);
nand U2867 (N_2867,N_2817,N_2802);
and U2868 (N_2868,N_2834,N_2839);
and U2869 (N_2869,N_2831,N_2814);
nor U2870 (N_2870,N_2806,N_2800);
or U2871 (N_2871,N_2845,N_2824);
and U2872 (N_2872,N_2811,N_2833);
and U2873 (N_2873,N_2841,N_2816);
xor U2874 (N_2874,N_2836,N_2825);
nand U2875 (N_2875,N_2821,N_2841);
and U2876 (N_2876,N_2849,N_2800);
and U2877 (N_2877,N_2837,N_2812);
nand U2878 (N_2878,N_2846,N_2843);
nand U2879 (N_2879,N_2848,N_2806);
and U2880 (N_2880,N_2803,N_2849);
nor U2881 (N_2881,N_2819,N_2814);
xnor U2882 (N_2882,N_2819,N_2829);
nor U2883 (N_2883,N_2830,N_2835);
nor U2884 (N_2884,N_2809,N_2814);
and U2885 (N_2885,N_2803,N_2829);
xor U2886 (N_2886,N_2802,N_2834);
nor U2887 (N_2887,N_2833,N_2848);
and U2888 (N_2888,N_2806,N_2801);
or U2889 (N_2889,N_2846,N_2813);
or U2890 (N_2890,N_2823,N_2808);
xnor U2891 (N_2891,N_2837,N_2828);
and U2892 (N_2892,N_2821,N_2830);
nor U2893 (N_2893,N_2806,N_2804);
xor U2894 (N_2894,N_2835,N_2804);
nor U2895 (N_2895,N_2816,N_2815);
and U2896 (N_2896,N_2849,N_2839);
nand U2897 (N_2897,N_2823,N_2838);
and U2898 (N_2898,N_2825,N_2801);
nor U2899 (N_2899,N_2833,N_2820);
nor U2900 (N_2900,N_2868,N_2889);
or U2901 (N_2901,N_2887,N_2890);
or U2902 (N_2902,N_2852,N_2873);
nand U2903 (N_2903,N_2898,N_2863);
xnor U2904 (N_2904,N_2882,N_2870);
nor U2905 (N_2905,N_2851,N_2881);
xor U2906 (N_2906,N_2854,N_2856);
and U2907 (N_2907,N_2871,N_2869);
nand U2908 (N_2908,N_2888,N_2895);
nand U2909 (N_2909,N_2857,N_2875);
nand U2910 (N_2910,N_2861,N_2878);
xor U2911 (N_2911,N_2897,N_2864);
and U2912 (N_2912,N_2886,N_2879);
or U2913 (N_2913,N_2850,N_2855);
nor U2914 (N_2914,N_2876,N_2867);
nand U2915 (N_2915,N_2862,N_2872);
xor U2916 (N_2916,N_2858,N_2877);
or U2917 (N_2917,N_2866,N_2891);
and U2918 (N_2918,N_2880,N_2874);
xnor U2919 (N_2919,N_2865,N_2859);
xnor U2920 (N_2920,N_2899,N_2883);
and U2921 (N_2921,N_2894,N_2885);
nand U2922 (N_2922,N_2853,N_2860);
xnor U2923 (N_2923,N_2893,N_2896);
or U2924 (N_2924,N_2884,N_2892);
xor U2925 (N_2925,N_2882,N_2897);
xnor U2926 (N_2926,N_2855,N_2895);
or U2927 (N_2927,N_2856,N_2899);
or U2928 (N_2928,N_2857,N_2888);
xor U2929 (N_2929,N_2859,N_2884);
nand U2930 (N_2930,N_2856,N_2867);
or U2931 (N_2931,N_2850,N_2883);
nor U2932 (N_2932,N_2880,N_2854);
nand U2933 (N_2933,N_2876,N_2895);
nand U2934 (N_2934,N_2859,N_2853);
or U2935 (N_2935,N_2890,N_2886);
nor U2936 (N_2936,N_2883,N_2890);
nor U2937 (N_2937,N_2897,N_2861);
xor U2938 (N_2938,N_2895,N_2851);
and U2939 (N_2939,N_2853,N_2886);
xnor U2940 (N_2940,N_2871,N_2857);
xor U2941 (N_2941,N_2882,N_2895);
xor U2942 (N_2942,N_2874,N_2879);
and U2943 (N_2943,N_2861,N_2852);
and U2944 (N_2944,N_2876,N_2853);
xor U2945 (N_2945,N_2889,N_2869);
nand U2946 (N_2946,N_2859,N_2870);
and U2947 (N_2947,N_2862,N_2890);
and U2948 (N_2948,N_2888,N_2861);
nor U2949 (N_2949,N_2870,N_2857);
nor U2950 (N_2950,N_2933,N_2912);
nand U2951 (N_2951,N_2907,N_2926);
xnor U2952 (N_2952,N_2936,N_2928);
and U2953 (N_2953,N_2923,N_2904);
xnor U2954 (N_2954,N_2920,N_2941);
and U2955 (N_2955,N_2922,N_2944);
and U2956 (N_2956,N_2943,N_2911);
and U2957 (N_2957,N_2946,N_2942);
nor U2958 (N_2958,N_2939,N_2909);
or U2959 (N_2959,N_2916,N_2919);
nand U2960 (N_2960,N_2930,N_2949);
nand U2961 (N_2961,N_2945,N_2937);
nand U2962 (N_2962,N_2903,N_2905);
and U2963 (N_2963,N_2900,N_2914);
or U2964 (N_2964,N_2947,N_2927);
xnor U2965 (N_2965,N_2929,N_2924);
xnor U2966 (N_2966,N_2921,N_2938);
nor U2967 (N_2967,N_2917,N_2918);
or U2968 (N_2968,N_2932,N_2913);
xnor U2969 (N_2969,N_2908,N_2940);
xor U2970 (N_2970,N_2902,N_2910);
nand U2971 (N_2971,N_2906,N_2925);
or U2972 (N_2972,N_2915,N_2948);
nor U2973 (N_2973,N_2935,N_2901);
nand U2974 (N_2974,N_2934,N_2931);
and U2975 (N_2975,N_2912,N_2942);
xor U2976 (N_2976,N_2949,N_2924);
or U2977 (N_2977,N_2928,N_2943);
xnor U2978 (N_2978,N_2903,N_2926);
nor U2979 (N_2979,N_2933,N_2905);
nand U2980 (N_2980,N_2934,N_2923);
nor U2981 (N_2981,N_2928,N_2947);
nor U2982 (N_2982,N_2918,N_2940);
nand U2983 (N_2983,N_2902,N_2922);
nor U2984 (N_2984,N_2924,N_2925);
xor U2985 (N_2985,N_2917,N_2911);
nand U2986 (N_2986,N_2936,N_2910);
or U2987 (N_2987,N_2939,N_2938);
xnor U2988 (N_2988,N_2924,N_2945);
xor U2989 (N_2989,N_2940,N_2907);
nand U2990 (N_2990,N_2908,N_2914);
and U2991 (N_2991,N_2948,N_2902);
xor U2992 (N_2992,N_2905,N_2947);
nand U2993 (N_2993,N_2920,N_2910);
xor U2994 (N_2994,N_2913,N_2934);
nand U2995 (N_2995,N_2939,N_2911);
nor U2996 (N_2996,N_2918,N_2934);
xor U2997 (N_2997,N_2937,N_2936);
and U2998 (N_2998,N_2943,N_2921);
and U2999 (N_2999,N_2926,N_2923);
and UO_0 (O_0,N_2975,N_2950);
and UO_1 (O_1,N_2989,N_2973);
xnor UO_2 (O_2,N_2982,N_2967);
and UO_3 (O_3,N_2957,N_2985);
nand UO_4 (O_4,N_2988,N_2960);
and UO_5 (O_5,N_2968,N_2953);
nand UO_6 (O_6,N_2951,N_2981);
and UO_7 (O_7,N_2999,N_2976);
xnor UO_8 (O_8,N_2964,N_2963);
nand UO_9 (O_9,N_2994,N_2986);
xnor UO_10 (O_10,N_2965,N_2984);
and UO_11 (O_11,N_2969,N_2983);
or UO_12 (O_12,N_2971,N_2961);
xnor UO_13 (O_13,N_2972,N_2958);
and UO_14 (O_14,N_2966,N_2955);
nor UO_15 (O_15,N_2970,N_2980);
nand UO_16 (O_16,N_2952,N_2978);
or UO_17 (O_17,N_2977,N_2997);
or UO_18 (O_18,N_2993,N_2954);
or UO_19 (O_19,N_2996,N_2987);
nor UO_20 (O_20,N_2962,N_2956);
nand UO_21 (O_21,N_2992,N_2990);
and UO_22 (O_22,N_2995,N_2979);
and UO_23 (O_23,N_2998,N_2991);
nor UO_24 (O_24,N_2974,N_2959);
xor UO_25 (O_25,N_2967,N_2986);
or UO_26 (O_26,N_2954,N_2963);
xnor UO_27 (O_27,N_2960,N_2964);
and UO_28 (O_28,N_2993,N_2963);
nand UO_29 (O_29,N_2951,N_2974);
xnor UO_30 (O_30,N_2951,N_2963);
nand UO_31 (O_31,N_2957,N_2993);
xor UO_32 (O_32,N_2977,N_2956);
and UO_33 (O_33,N_2990,N_2987);
nor UO_34 (O_34,N_2958,N_2963);
xnor UO_35 (O_35,N_2962,N_2996);
and UO_36 (O_36,N_2987,N_2951);
nand UO_37 (O_37,N_2981,N_2960);
and UO_38 (O_38,N_2969,N_2982);
xor UO_39 (O_39,N_2998,N_2978);
or UO_40 (O_40,N_2972,N_2960);
or UO_41 (O_41,N_2951,N_2955);
nor UO_42 (O_42,N_2993,N_2985);
nor UO_43 (O_43,N_2970,N_2992);
and UO_44 (O_44,N_2976,N_2971);
nand UO_45 (O_45,N_2995,N_2976);
nor UO_46 (O_46,N_2983,N_2967);
nand UO_47 (O_47,N_2960,N_2962);
or UO_48 (O_48,N_2988,N_2978);
nand UO_49 (O_49,N_2978,N_2971);
nand UO_50 (O_50,N_2990,N_2973);
or UO_51 (O_51,N_2989,N_2969);
nor UO_52 (O_52,N_2959,N_2968);
or UO_53 (O_53,N_2979,N_2993);
or UO_54 (O_54,N_2993,N_2960);
xnor UO_55 (O_55,N_2977,N_2970);
or UO_56 (O_56,N_2995,N_2978);
and UO_57 (O_57,N_2958,N_2979);
or UO_58 (O_58,N_2964,N_2991);
and UO_59 (O_59,N_2975,N_2978);
or UO_60 (O_60,N_2969,N_2978);
nand UO_61 (O_61,N_2967,N_2995);
nand UO_62 (O_62,N_2981,N_2976);
nor UO_63 (O_63,N_2990,N_2972);
nand UO_64 (O_64,N_2971,N_2984);
nand UO_65 (O_65,N_2980,N_2963);
and UO_66 (O_66,N_2961,N_2969);
and UO_67 (O_67,N_2953,N_2972);
and UO_68 (O_68,N_2952,N_2998);
or UO_69 (O_69,N_2977,N_2963);
nand UO_70 (O_70,N_2958,N_2998);
and UO_71 (O_71,N_2968,N_2995);
or UO_72 (O_72,N_2994,N_2970);
or UO_73 (O_73,N_2950,N_2962);
nand UO_74 (O_74,N_2979,N_2981);
nand UO_75 (O_75,N_2958,N_2967);
xnor UO_76 (O_76,N_2970,N_2993);
xor UO_77 (O_77,N_2985,N_2990);
xnor UO_78 (O_78,N_2975,N_2962);
nand UO_79 (O_79,N_2953,N_2979);
xor UO_80 (O_80,N_2986,N_2969);
or UO_81 (O_81,N_2972,N_2988);
and UO_82 (O_82,N_2977,N_2992);
nor UO_83 (O_83,N_2987,N_2983);
and UO_84 (O_84,N_2976,N_2992);
nor UO_85 (O_85,N_2991,N_2955);
xor UO_86 (O_86,N_2971,N_2992);
or UO_87 (O_87,N_2950,N_2990);
nand UO_88 (O_88,N_2983,N_2989);
xor UO_89 (O_89,N_2992,N_2974);
nor UO_90 (O_90,N_2965,N_2959);
xnor UO_91 (O_91,N_2970,N_2973);
nand UO_92 (O_92,N_2959,N_2979);
or UO_93 (O_93,N_2991,N_2959);
nor UO_94 (O_94,N_2990,N_2968);
and UO_95 (O_95,N_2964,N_2965);
nand UO_96 (O_96,N_2990,N_2999);
xor UO_97 (O_97,N_2982,N_2966);
or UO_98 (O_98,N_2959,N_2976);
xor UO_99 (O_99,N_2958,N_2993);
or UO_100 (O_100,N_2992,N_2987);
nor UO_101 (O_101,N_2970,N_2989);
and UO_102 (O_102,N_2976,N_2963);
nand UO_103 (O_103,N_2987,N_2970);
or UO_104 (O_104,N_2950,N_2984);
or UO_105 (O_105,N_2968,N_2977);
or UO_106 (O_106,N_2968,N_2992);
xnor UO_107 (O_107,N_2970,N_2962);
or UO_108 (O_108,N_2959,N_2999);
xnor UO_109 (O_109,N_2993,N_2967);
nand UO_110 (O_110,N_2960,N_2965);
nand UO_111 (O_111,N_2973,N_2993);
nand UO_112 (O_112,N_2975,N_2953);
nor UO_113 (O_113,N_2985,N_2958);
nor UO_114 (O_114,N_2985,N_2982);
and UO_115 (O_115,N_2971,N_2979);
nand UO_116 (O_116,N_2971,N_2952);
nor UO_117 (O_117,N_2962,N_2979);
nor UO_118 (O_118,N_2995,N_2966);
nand UO_119 (O_119,N_2961,N_2955);
nor UO_120 (O_120,N_2998,N_2999);
and UO_121 (O_121,N_2974,N_2955);
nand UO_122 (O_122,N_2962,N_2998);
xor UO_123 (O_123,N_2980,N_2992);
or UO_124 (O_124,N_2981,N_2954);
xnor UO_125 (O_125,N_2964,N_2961);
or UO_126 (O_126,N_2983,N_2951);
xor UO_127 (O_127,N_2966,N_2978);
or UO_128 (O_128,N_2962,N_2953);
nand UO_129 (O_129,N_2957,N_2970);
and UO_130 (O_130,N_2951,N_2965);
nand UO_131 (O_131,N_2992,N_2963);
and UO_132 (O_132,N_2969,N_2979);
or UO_133 (O_133,N_2976,N_2958);
xor UO_134 (O_134,N_2960,N_2952);
and UO_135 (O_135,N_2953,N_2986);
xnor UO_136 (O_136,N_2980,N_2997);
xnor UO_137 (O_137,N_2987,N_2962);
nor UO_138 (O_138,N_2950,N_2957);
or UO_139 (O_139,N_2997,N_2982);
nand UO_140 (O_140,N_2973,N_2960);
or UO_141 (O_141,N_2966,N_2974);
and UO_142 (O_142,N_2998,N_2954);
or UO_143 (O_143,N_2956,N_2963);
nand UO_144 (O_144,N_2974,N_2952);
and UO_145 (O_145,N_2954,N_2973);
xnor UO_146 (O_146,N_2950,N_2999);
or UO_147 (O_147,N_2955,N_2979);
nor UO_148 (O_148,N_2950,N_2979);
and UO_149 (O_149,N_2964,N_2969);
xor UO_150 (O_150,N_2988,N_2990);
nor UO_151 (O_151,N_2995,N_2974);
xnor UO_152 (O_152,N_2959,N_2962);
xnor UO_153 (O_153,N_2953,N_2966);
nor UO_154 (O_154,N_2984,N_2997);
or UO_155 (O_155,N_2985,N_2966);
xor UO_156 (O_156,N_2981,N_2972);
nor UO_157 (O_157,N_2993,N_2965);
xor UO_158 (O_158,N_2950,N_2991);
xnor UO_159 (O_159,N_2954,N_2986);
or UO_160 (O_160,N_2968,N_2960);
or UO_161 (O_161,N_2985,N_2997);
nor UO_162 (O_162,N_2951,N_2957);
nand UO_163 (O_163,N_2992,N_2967);
nand UO_164 (O_164,N_2966,N_2991);
nor UO_165 (O_165,N_2984,N_2957);
and UO_166 (O_166,N_2999,N_2991);
nor UO_167 (O_167,N_2971,N_2967);
nand UO_168 (O_168,N_2963,N_2999);
nand UO_169 (O_169,N_2951,N_2977);
nor UO_170 (O_170,N_2992,N_2962);
nand UO_171 (O_171,N_2980,N_2955);
and UO_172 (O_172,N_2975,N_2952);
nand UO_173 (O_173,N_2980,N_2971);
xnor UO_174 (O_174,N_2991,N_2965);
or UO_175 (O_175,N_2989,N_2996);
nand UO_176 (O_176,N_2980,N_2993);
nand UO_177 (O_177,N_2980,N_2957);
nor UO_178 (O_178,N_2983,N_2988);
nand UO_179 (O_179,N_2996,N_2986);
nor UO_180 (O_180,N_2954,N_2967);
nand UO_181 (O_181,N_2960,N_2985);
xor UO_182 (O_182,N_2959,N_2955);
and UO_183 (O_183,N_2961,N_2978);
nor UO_184 (O_184,N_2956,N_2968);
nor UO_185 (O_185,N_2956,N_2995);
and UO_186 (O_186,N_2972,N_2977);
and UO_187 (O_187,N_2979,N_2987);
xnor UO_188 (O_188,N_2960,N_2979);
nand UO_189 (O_189,N_2975,N_2970);
or UO_190 (O_190,N_2971,N_2997);
nand UO_191 (O_191,N_2965,N_2996);
xor UO_192 (O_192,N_2976,N_2970);
nor UO_193 (O_193,N_2983,N_2985);
nor UO_194 (O_194,N_2957,N_2966);
or UO_195 (O_195,N_2962,N_2997);
xor UO_196 (O_196,N_2984,N_2973);
and UO_197 (O_197,N_2997,N_2961);
nor UO_198 (O_198,N_2965,N_2998);
nor UO_199 (O_199,N_2980,N_2995);
or UO_200 (O_200,N_2967,N_2960);
or UO_201 (O_201,N_2963,N_2970);
nand UO_202 (O_202,N_2962,N_2974);
xor UO_203 (O_203,N_2977,N_2967);
nor UO_204 (O_204,N_2980,N_2954);
and UO_205 (O_205,N_2990,N_2986);
nor UO_206 (O_206,N_2963,N_2982);
xor UO_207 (O_207,N_2953,N_2964);
xor UO_208 (O_208,N_2971,N_2975);
and UO_209 (O_209,N_2957,N_2956);
xor UO_210 (O_210,N_2986,N_2974);
nor UO_211 (O_211,N_2992,N_2957);
xor UO_212 (O_212,N_2953,N_2973);
or UO_213 (O_213,N_2968,N_2955);
nand UO_214 (O_214,N_2957,N_2972);
nand UO_215 (O_215,N_2985,N_2951);
or UO_216 (O_216,N_2977,N_2962);
nand UO_217 (O_217,N_2980,N_2964);
and UO_218 (O_218,N_2995,N_2999);
and UO_219 (O_219,N_2989,N_2992);
xnor UO_220 (O_220,N_2995,N_2996);
nand UO_221 (O_221,N_2983,N_2980);
xnor UO_222 (O_222,N_2978,N_2996);
or UO_223 (O_223,N_2951,N_2975);
and UO_224 (O_224,N_2976,N_2983);
and UO_225 (O_225,N_2974,N_2976);
xor UO_226 (O_226,N_2983,N_2981);
xor UO_227 (O_227,N_2955,N_2981);
or UO_228 (O_228,N_2964,N_2981);
nor UO_229 (O_229,N_2986,N_2993);
xnor UO_230 (O_230,N_2984,N_2994);
nand UO_231 (O_231,N_2975,N_2977);
and UO_232 (O_232,N_2975,N_2961);
xnor UO_233 (O_233,N_2990,N_2975);
and UO_234 (O_234,N_2973,N_2981);
nand UO_235 (O_235,N_2968,N_2973);
and UO_236 (O_236,N_2998,N_2995);
or UO_237 (O_237,N_2961,N_2981);
nand UO_238 (O_238,N_2997,N_2950);
xor UO_239 (O_239,N_2984,N_2996);
and UO_240 (O_240,N_2965,N_2980);
and UO_241 (O_241,N_2994,N_2960);
and UO_242 (O_242,N_2984,N_2952);
nand UO_243 (O_243,N_2991,N_2989);
and UO_244 (O_244,N_2971,N_2953);
nor UO_245 (O_245,N_2998,N_2974);
nand UO_246 (O_246,N_2990,N_2963);
nand UO_247 (O_247,N_2957,N_2983);
nand UO_248 (O_248,N_2989,N_2995);
and UO_249 (O_249,N_2977,N_2976);
xnor UO_250 (O_250,N_2968,N_2950);
or UO_251 (O_251,N_2984,N_2956);
or UO_252 (O_252,N_2954,N_2997);
or UO_253 (O_253,N_2975,N_2998);
nand UO_254 (O_254,N_2975,N_2995);
and UO_255 (O_255,N_2982,N_2968);
or UO_256 (O_256,N_2985,N_2969);
nand UO_257 (O_257,N_2986,N_2964);
nor UO_258 (O_258,N_2976,N_2967);
and UO_259 (O_259,N_2995,N_2959);
nor UO_260 (O_260,N_2968,N_2980);
nor UO_261 (O_261,N_2983,N_2970);
xnor UO_262 (O_262,N_2979,N_2978);
nor UO_263 (O_263,N_2990,N_2967);
or UO_264 (O_264,N_2969,N_2955);
nor UO_265 (O_265,N_2979,N_2991);
and UO_266 (O_266,N_2975,N_2958);
or UO_267 (O_267,N_2993,N_2951);
xor UO_268 (O_268,N_2996,N_2969);
and UO_269 (O_269,N_2979,N_2988);
xnor UO_270 (O_270,N_2959,N_2993);
nand UO_271 (O_271,N_2983,N_2956);
and UO_272 (O_272,N_2956,N_2999);
nand UO_273 (O_273,N_2991,N_2982);
xor UO_274 (O_274,N_2999,N_2985);
and UO_275 (O_275,N_2951,N_2961);
and UO_276 (O_276,N_2982,N_2984);
nor UO_277 (O_277,N_2976,N_2964);
or UO_278 (O_278,N_2976,N_2965);
or UO_279 (O_279,N_2991,N_2996);
nand UO_280 (O_280,N_2988,N_2952);
and UO_281 (O_281,N_2990,N_2976);
or UO_282 (O_282,N_2974,N_2982);
or UO_283 (O_283,N_2966,N_2975);
or UO_284 (O_284,N_2953,N_2991);
or UO_285 (O_285,N_2975,N_2992);
xor UO_286 (O_286,N_2961,N_2988);
nor UO_287 (O_287,N_2988,N_2984);
and UO_288 (O_288,N_2957,N_2976);
nor UO_289 (O_289,N_2973,N_2991);
nor UO_290 (O_290,N_2981,N_2977);
or UO_291 (O_291,N_2964,N_2959);
nor UO_292 (O_292,N_2960,N_2989);
nand UO_293 (O_293,N_2969,N_2950);
or UO_294 (O_294,N_2991,N_2978);
nor UO_295 (O_295,N_2968,N_2958);
xnor UO_296 (O_296,N_2967,N_2991);
xnor UO_297 (O_297,N_2980,N_2986);
and UO_298 (O_298,N_2993,N_2964);
xnor UO_299 (O_299,N_2966,N_2976);
nand UO_300 (O_300,N_2980,N_2972);
nand UO_301 (O_301,N_2983,N_2992);
nor UO_302 (O_302,N_2998,N_2951);
xor UO_303 (O_303,N_2950,N_2956);
nor UO_304 (O_304,N_2995,N_2950);
nor UO_305 (O_305,N_2990,N_2989);
nand UO_306 (O_306,N_2960,N_2997);
or UO_307 (O_307,N_2984,N_2964);
xnor UO_308 (O_308,N_2952,N_2993);
nand UO_309 (O_309,N_2989,N_2967);
and UO_310 (O_310,N_2988,N_2969);
xor UO_311 (O_311,N_2982,N_2979);
and UO_312 (O_312,N_2976,N_2968);
and UO_313 (O_313,N_2992,N_2953);
nand UO_314 (O_314,N_2984,N_2969);
nand UO_315 (O_315,N_2995,N_2991);
and UO_316 (O_316,N_2960,N_2974);
xor UO_317 (O_317,N_2968,N_2954);
nor UO_318 (O_318,N_2952,N_2973);
xnor UO_319 (O_319,N_2972,N_2995);
or UO_320 (O_320,N_2978,N_2980);
and UO_321 (O_321,N_2958,N_2971);
nor UO_322 (O_322,N_2973,N_2972);
and UO_323 (O_323,N_2997,N_2981);
and UO_324 (O_324,N_2984,N_2960);
or UO_325 (O_325,N_2980,N_2982);
nand UO_326 (O_326,N_2960,N_2998);
xnor UO_327 (O_327,N_2962,N_2995);
nor UO_328 (O_328,N_2972,N_2983);
or UO_329 (O_329,N_2951,N_2954);
or UO_330 (O_330,N_2995,N_2983);
or UO_331 (O_331,N_2996,N_2961);
nand UO_332 (O_332,N_2961,N_2989);
and UO_333 (O_333,N_2987,N_2957);
nor UO_334 (O_334,N_2980,N_2956);
nor UO_335 (O_335,N_2955,N_2964);
xnor UO_336 (O_336,N_2989,N_2968);
or UO_337 (O_337,N_2972,N_2966);
nand UO_338 (O_338,N_2966,N_2954);
or UO_339 (O_339,N_2955,N_2965);
nand UO_340 (O_340,N_2997,N_2998);
nand UO_341 (O_341,N_2986,N_2960);
nor UO_342 (O_342,N_2960,N_2966);
nor UO_343 (O_343,N_2962,N_2972);
nand UO_344 (O_344,N_2965,N_2966);
and UO_345 (O_345,N_2972,N_2955);
nand UO_346 (O_346,N_2958,N_2970);
and UO_347 (O_347,N_2959,N_2961);
or UO_348 (O_348,N_2998,N_2984);
xor UO_349 (O_349,N_2951,N_2995);
nand UO_350 (O_350,N_2963,N_2994);
and UO_351 (O_351,N_2979,N_2999);
xnor UO_352 (O_352,N_2976,N_2952);
or UO_353 (O_353,N_2976,N_2962);
or UO_354 (O_354,N_2966,N_2994);
and UO_355 (O_355,N_2957,N_2969);
nor UO_356 (O_356,N_2987,N_2961);
nand UO_357 (O_357,N_2987,N_2995);
nand UO_358 (O_358,N_2981,N_2971);
nand UO_359 (O_359,N_2970,N_2950);
nor UO_360 (O_360,N_2957,N_2982);
nand UO_361 (O_361,N_2955,N_2997);
nor UO_362 (O_362,N_2978,N_2960);
and UO_363 (O_363,N_2977,N_2988);
and UO_364 (O_364,N_2982,N_2955);
and UO_365 (O_365,N_2975,N_2985);
nor UO_366 (O_366,N_2989,N_2999);
and UO_367 (O_367,N_2952,N_2999);
or UO_368 (O_368,N_2972,N_2952);
nand UO_369 (O_369,N_2984,N_2966);
nor UO_370 (O_370,N_2987,N_2950);
and UO_371 (O_371,N_2998,N_2979);
nor UO_372 (O_372,N_2963,N_2973);
or UO_373 (O_373,N_2984,N_2980);
and UO_374 (O_374,N_2967,N_2952);
or UO_375 (O_375,N_2961,N_2957);
nand UO_376 (O_376,N_2955,N_2960);
nor UO_377 (O_377,N_2955,N_2985);
and UO_378 (O_378,N_2995,N_2954);
nand UO_379 (O_379,N_2960,N_2957);
nand UO_380 (O_380,N_2973,N_2962);
nor UO_381 (O_381,N_2969,N_2966);
and UO_382 (O_382,N_2987,N_2959);
nand UO_383 (O_383,N_2996,N_2951);
nor UO_384 (O_384,N_2986,N_2950);
xor UO_385 (O_385,N_2970,N_2996);
xnor UO_386 (O_386,N_2966,N_2990);
nor UO_387 (O_387,N_2990,N_2981);
or UO_388 (O_388,N_2972,N_2989);
xor UO_389 (O_389,N_2970,N_2971);
nor UO_390 (O_390,N_2979,N_2994);
or UO_391 (O_391,N_2954,N_2989);
or UO_392 (O_392,N_2982,N_2999);
xor UO_393 (O_393,N_2983,N_2978);
xor UO_394 (O_394,N_2991,N_2963);
or UO_395 (O_395,N_2997,N_2957);
xnor UO_396 (O_396,N_2970,N_2964);
or UO_397 (O_397,N_2971,N_2988);
nor UO_398 (O_398,N_2981,N_2967);
nand UO_399 (O_399,N_2991,N_2962);
nand UO_400 (O_400,N_2990,N_2951);
or UO_401 (O_401,N_2971,N_2982);
or UO_402 (O_402,N_2967,N_2970);
nand UO_403 (O_403,N_2961,N_2995);
or UO_404 (O_404,N_2988,N_2991);
nand UO_405 (O_405,N_2987,N_2989);
nor UO_406 (O_406,N_2986,N_2983);
xor UO_407 (O_407,N_2974,N_2950);
nor UO_408 (O_408,N_2952,N_2981);
nor UO_409 (O_409,N_2977,N_2996);
nand UO_410 (O_410,N_2956,N_2973);
nand UO_411 (O_411,N_2996,N_2994);
nand UO_412 (O_412,N_2951,N_2992);
xor UO_413 (O_413,N_2963,N_2986);
xor UO_414 (O_414,N_2981,N_2980);
nor UO_415 (O_415,N_2957,N_2990);
or UO_416 (O_416,N_2985,N_2980);
nand UO_417 (O_417,N_2990,N_2955);
and UO_418 (O_418,N_2990,N_2995);
or UO_419 (O_419,N_2969,N_2968);
and UO_420 (O_420,N_2974,N_2971);
nor UO_421 (O_421,N_2954,N_2996);
nand UO_422 (O_422,N_2982,N_2996);
nor UO_423 (O_423,N_2951,N_2973);
or UO_424 (O_424,N_2981,N_2966);
xnor UO_425 (O_425,N_2959,N_2978);
nor UO_426 (O_426,N_2995,N_2997);
nor UO_427 (O_427,N_2952,N_2983);
or UO_428 (O_428,N_2972,N_2974);
and UO_429 (O_429,N_2970,N_2988);
nand UO_430 (O_430,N_2998,N_2981);
or UO_431 (O_431,N_2969,N_2998);
xor UO_432 (O_432,N_2994,N_2969);
nand UO_433 (O_433,N_2967,N_2963);
or UO_434 (O_434,N_2967,N_2966);
xnor UO_435 (O_435,N_2983,N_2955);
nand UO_436 (O_436,N_2989,N_2951);
nor UO_437 (O_437,N_2986,N_2987);
nor UO_438 (O_438,N_2955,N_2986);
or UO_439 (O_439,N_2952,N_2980);
nand UO_440 (O_440,N_2974,N_2997);
nand UO_441 (O_441,N_2953,N_2989);
xor UO_442 (O_442,N_2950,N_2961);
or UO_443 (O_443,N_2969,N_2959);
nor UO_444 (O_444,N_2983,N_2961);
xnor UO_445 (O_445,N_2958,N_2994);
nor UO_446 (O_446,N_2999,N_2953);
or UO_447 (O_447,N_2963,N_2955);
nand UO_448 (O_448,N_2995,N_2973);
nand UO_449 (O_449,N_2988,N_2975);
xnor UO_450 (O_450,N_2983,N_2984);
xnor UO_451 (O_451,N_2962,N_2990);
or UO_452 (O_452,N_2986,N_2992);
or UO_453 (O_453,N_2969,N_2962);
or UO_454 (O_454,N_2979,N_2966);
or UO_455 (O_455,N_2984,N_2987);
and UO_456 (O_456,N_2979,N_2974);
and UO_457 (O_457,N_2953,N_2951);
nor UO_458 (O_458,N_2995,N_2957);
xnor UO_459 (O_459,N_2952,N_2958);
xnor UO_460 (O_460,N_2984,N_2961);
xnor UO_461 (O_461,N_2957,N_2978);
and UO_462 (O_462,N_2978,N_2990);
nor UO_463 (O_463,N_2977,N_2979);
nor UO_464 (O_464,N_2999,N_2960);
or UO_465 (O_465,N_2992,N_2969);
and UO_466 (O_466,N_2953,N_2950);
nor UO_467 (O_467,N_2957,N_2958);
or UO_468 (O_468,N_2958,N_2992);
and UO_469 (O_469,N_2973,N_2966);
or UO_470 (O_470,N_2957,N_2999);
xnor UO_471 (O_471,N_2981,N_2956);
nand UO_472 (O_472,N_2996,N_2950);
and UO_473 (O_473,N_2965,N_2990);
xnor UO_474 (O_474,N_2964,N_2997);
and UO_475 (O_475,N_2994,N_2977);
nor UO_476 (O_476,N_2993,N_2976);
nor UO_477 (O_477,N_2977,N_2974);
or UO_478 (O_478,N_2998,N_2967);
and UO_479 (O_479,N_2977,N_2971);
or UO_480 (O_480,N_2968,N_2967);
nor UO_481 (O_481,N_2989,N_2998);
nand UO_482 (O_482,N_2998,N_2987);
nand UO_483 (O_483,N_2960,N_2951);
nand UO_484 (O_484,N_2988,N_2956);
and UO_485 (O_485,N_2980,N_2960);
xor UO_486 (O_486,N_2958,N_2955);
or UO_487 (O_487,N_2985,N_2981);
xnor UO_488 (O_488,N_2959,N_2973);
xnor UO_489 (O_489,N_2971,N_2995);
nand UO_490 (O_490,N_2957,N_2977);
nor UO_491 (O_491,N_2961,N_2990);
xor UO_492 (O_492,N_2961,N_2962);
and UO_493 (O_493,N_2958,N_2988);
or UO_494 (O_494,N_2959,N_2953);
xor UO_495 (O_495,N_2976,N_2997);
or UO_496 (O_496,N_2989,N_2950);
and UO_497 (O_497,N_2955,N_2976);
or UO_498 (O_498,N_2955,N_2962);
nand UO_499 (O_499,N_2963,N_2950);
endmodule