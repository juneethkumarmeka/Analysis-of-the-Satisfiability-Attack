module basic_500_3000_500_30_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_283,In_476);
or U1 (N_1,In_298,In_390);
nand U2 (N_2,In_329,In_377);
nand U3 (N_3,In_312,In_247);
nor U4 (N_4,In_399,In_76);
nor U5 (N_5,In_434,In_419);
nand U6 (N_6,In_279,In_168);
and U7 (N_7,In_275,In_471);
or U8 (N_8,In_70,In_388);
or U9 (N_9,In_95,In_189);
and U10 (N_10,In_254,In_342);
nand U11 (N_11,In_425,In_292);
nand U12 (N_12,In_84,In_307);
nor U13 (N_13,In_367,In_125);
nor U14 (N_14,In_205,In_6);
or U15 (N_15,In_261,In_305);
nor U16 (N_16,In_55,In_196);
nor U17 (N_17,In_228,In_437);
and U18 (N_18,In_358,In_89);
nand U19 (N_19,In_128,In_490);
nor U20 (N_20,In_314,In_308);
nor U21 (N_21,In_429,In_225);
and U22 (N_22,In_334,In_3);
nand U23 (N_23,In_480,In_348);
or U24 (N_24,In_265,In_301);
nor U25 (N_25,In_58,In_167);
nand U26 (N_26,In_468,In_42);
nand U27 (N_27,In_330,In_221);
nand U28 (N_28,In_460,In_363);
nor U29 (N_29,In_484,In_416);
nand U30 (N_30,In_467,In_411);
or U31 (N_31,In_121,In_430);
or U32 (N_32,In_19,In_17);
nand U33 (N_33,In_266,In_68);
or U34 (N_34,In_244,In_379);
nand U35 (N_35,In_396,In_188);
nor U36 (N_36,In_286,In_146);
nor U37 (N_37,In_236,In_232);
nor U38 (N_38,In_290,In_372);
and U39 (N_39,In_245,In_198);
and U40 (N_40,In_106,In_457);
nand U41 (N_41,In_133,In_63);
and U42 (N_42,In_256,In_459);
nor U43 (N_43,In_392,In_152);
and U44 (N_44,In_145,In_439);
nand U45 (N_45,In_424,In_331);
and U46 (N_46,In_113,In_495);
nand U47 (N_47,In_357,In_90);
or U48 (N_48,In_497,In_412);
nand U49 (N_49,In_155,In_165);
nor U50 (N_50,In_365,In_317);
nand U51 (N_51,In_11,In_364);
nand U52 (N_52,In_448,In_354);
or U53 (N_53,In_224,In_151);
or U54 (N_54,In_216,In_85);
and U55 (N_55,In_240,In_176);
or U56 (N_56,In_453,In_96);
nor U57 (N_57,In_81,In_253);
nor U58 (N_58,In_289,In_190);
and U59 (N_59,In_131,In_220);
nor U60 (N_60,In_227,In_80);
and U61 (N_61,In_483,In_455);
and U62 (N_62,In_77,In_233);
or U63 (N_63,In_138,In_405);
and U64 (N_64,In_383,In_132);
and U65 (N_65,In_154,In_444);
nor U66 (N_66,In_470,In_347);
nor U67 (N_67,In_296,In_440);
nand U68 (N_68,In_403,In_208);
nor U69 (N_69,In_28,In_79);
xor U70 (N_70,In_466,In_461);
and U71 (N_71,In_36,In_248);
and U72 (N_72,In_172,In_242);
and U73 (N_73,In_114,In_27);
nand U74 (N_74,In_87,In_108);
nor U75 (N_75,In_257,In_285);
nor U76 (N_76,In_309,In_99);
or U77 (N_77,In_452,In_226);
and U78 (N_78,In_213,In_215);
nand U79 (N_79,In_140,In_182);
or U80 (N_80,In_281,In_243);
nor U81 (N_81,In_35,In_16);
nor U82 (N_82,In_291,In_384);
nor U83 (N_83,In_426,In_97);
nor U84 (N_84,In_170,In_373);
nand U85 (N_85,In_339,In_45);
or U86 (N_86,In_310,In_259);
and U87 (N_87,In_263,In_159);
nor U88 (N_88,In_360,In_336);
nand U89 (N_89,In_116,In_287);
nor U90 (N_90,In_93,In_157);
nand U91 (N_91,In_178,In_201);
nor U92 (N_92,In_166,In_12);
and U93 (N_93,In_351,In_212);
nand U94 (N_94,In_272,In_187);
nor U95 (N_95,In_100,In_23);
nor U96 (N_96,In_139,In_418);
nor U97 (N_97,In_445,In_137);
or U98 (N_98,In_371,In_498);
nand U99 (N_99,In_436,In_163);
nor U100 (N_100,In_447,N_88);
nand U101 (N_101,In_62,In_73);
xnor U102 (N_102,In_343,In_238);
and U103 (N_103,In_134,In_472);
or U104 (N_104,In_414,In_278);
and U105 (N_105,In_10,In_118);
and U106 (N_106,In_191,N_92);
nor U107 (N_107,In_361,N_75);
and U108 (N_108,N_9,N_64);
or U109 (N_109,In_127,In_442);
nor U110 (N_110,In_295,In_142);
nand U111 (N_111,N_30,In_462);
or U112 (N_112,N_6,N_38);
and U113 (N_113,In_102,N_52);
nor U114 (N_114,N_10,N_34);
or U115 (N_115,In_41,In_417);
nand U116 (N_116,In_297,In_86);
and U117 (N_117,In_315,N_48);
nand U118 (N_118,In_61,N_33);
and U119 (N_119,N_98,In_465);
nand U120 (N_120,In_88,In_162);
and U121 (N_121,In_120,In_115);
nor U122 (N_122,In_177,In_326);
and U123 (N_123,In_147,In_274);
or U124 (N_124,N_50,N_61);
nor U125 (N_125,N_76,In_313);
or U126 (N_126,In_104,In_485);
nor U127 (N_127,N_22,N_62);
nand U128 (N_128,In_258,In_280);
and U129 (N_129,N_35,N_13);
nor U130 (N_130,N_31,N_55);
nand U131 (N_131,In_318,In_370);
or U132 (N_132,In_402,N_45);
nand U133 (N_133,In_345,In_303);
and U134 (N_134,N_63,N_83);
or U135 (N_135,In_148,In_92);
and U136 (N_136,In_401,In_250);
nor U137 (N_137,In_323,N_57);
nor U138 (N_138,In_391,In_423);
nand U139 (N_139,N_68,N_77);
nor U140 (N_140,In_122,In_319);
nor U141 (N_141,In_456,In_180);
and U142 (N_142,In_78,In_98);
or U143 (N_143,In_341,In_130);
or U144 (N_144,In_438,In_433);
nor U145 (N_145,In_491,In_450);
or U146 (N_146,In_386,In_69);
or U147 (N_147,In_209,In_204);
nand U148 (N_148,N_25,In_481);
xor U149 (N_149,N_11,In_385);
nor U150 (N_150,In_400,In_469);
nand U151 (N_151,N_0,In_2);
nand U152 (N_152,In_192,In_397);
nand U153 (N_153,In_474,In_299);
nor U154 (N_154,In_464,N_80);
and U155 (N_155,N_94,In_206);
nor U156 (N_156,N_4,In_67);
or U157 (N_157,In_194,In_454);
nand U158 (N_158,In_9,In_18);
and U159 (N_159,In_273,N_41);
or U160 (N_160,N_28,In_241);
nand U161 (N_161,In_202,In_338);
nand U162 (N_162,In_135,In_94);
or U163 (N_163,In_161,In_449);
nand U164 (N_164,In_267,In_304);
or U165 (N_165,In_332,In_222);
and U166 (N_166,N_44,In_349);
and U167 (N_167,N_69,N_32);
nor U168 (N_168,In_487,In_389);
or U169 (N_169,In_443,In_5);
and U170 (N_170,In_302,N_90);
or U171 (N_171,In_378,In_368);
nand U172 (N_172,In_49,In_268);
and U173 (N_173,In_31,In_21);
or U174 (N_174,N_7,In_179);
nor U175 (N_175,In_219,In_420);
or U176 (N_176,In_398,N_87);
nand U177 (N_177,In_38,In_51);
and U178 (N_178,In_284,N_20);
nor U179 (N_179,In_37,N_49);
and U180 (N_180,In_340,In_44);
or U181 (N_181,In_382,In_143);
nor U182 (N_182,In_328,In_404);
xor U183 (N_183,In_101,In_48);
nor U184 (N_184,In_200,In_83);
or U185 (N_185,In_393,In_229);
nor U186 (N_186,N_59,N_23);
nand U187 (N_187,In_119,In_160);
nand U188 (N_188,In_327,In_20);
or U189 (N_189,In_376,In_344);
nor U190 (N_190,In_427,In_375);
and U191 (N_191,N_5,In_288);
or U192 (N_192,In_493,In_496);
nor U193 (N_193,N_14,N_51);
and U194 (N_194,N_72,N_24);
and U195 (N_195,In_321,In_197);
nand U196 (N_196,In_269,In_75);
or U197 (N_197,In_210,N_84);
or U198 (N_198,In_24,N_99);
nor U199 (N_199,N_47,N_29);
or U200 (N_200,In_282,N_60);
and U201 (N_201,N_43,N_82);
nand U202 (N_202,N_183,In_322);
nor U203 (N_203,N_114,In_195);
nor U204 (N_204,N_165,In_488);
and U205 (N_205,In_366,In_136);
nor U206 (N_206,In_107,N_104);
or U207 (N_207,In_7,In_320);
nand U208 (N_208,In_234,N_168);
nor U209 (N_209,N_107,N_113);
nand U210 (N_210,N_173,In_489);
and U211 (N_211,N_151,N_127);
nand U212 (N_212,N_15,N_56);
nand U213 (N_213,In_395,In_277);
nor U214 (N_214,In_239,N_27);
or U215 (N_215,N_154,In_126);
nor U216 (N_216,N_132,In_494);
or U217 (N_217,N_152,In_184);
nor U218 (N_218,In_421,In_158);
nand U219 (N_219,N_180,N_118);
nand U220 (N_220,N_96,N_140);
and U221 (N_221,N_115,N_160);
and U222 (N_222,N_71,N_175);
or U223 (N_223,N_58,N_81);
or U224 (N_224,In_374,In_13);
and U225 (N_225,In_262,In_231);
or U226 (N_226,In_446,In_82);
and U227 (N_227,N_199,In_57);
nand U228 (N_228,N_184,In_71);
nand U229 (N_229,In_53,N_167);
nand U230 (N_230,In_249,N_73);
xnor U231 (N_231,N_166,N_155);
or U232 (N_232,N_97,In_482);
nor U233 (N_233,N_150,N_67);
or U234 (N_234,In_185,N_12);
nor U235 (N_235,N_53,N_133);
and U236 (N_236,In_217,In_251);
nor U237 (N_237,N_109,In_47);
or U238 (N_238,N_106,N_39);
nand U239 (N_239,N_65,N_85);
or U240 (N_240,In_355,N_158);
or U241 (N_241,N_131,N_86);
or U242 (N_242,In_117,N_36);
or U243 (N_243,In_214,N_17);
or U244 (N_244,N_26,In_359);
or U245 (N_245,In_207,N_105);
and U246 (N_246,In_171,In_276);
and U247 (N_247,In_66,In_410);
nand U248 (N_248,N_144,In_103);
or U249 (N_249,In_352,N_130);
and U250 (N_250,In_407,N_194);
nand U251 (N_251,In_333,In_22);
nand U252 (N_252,In_156,N_2);
and U253 (N_253,In_25,N_141);
and U254 (N_254,In_353,N_101);
nor U255 (N_255,N_146,In_169);
or U256 (N_256,In_60,N_156);
nand U257 (N_257,N_191,In_14);
nand U258 (N_258,N_171,In_1);
or U259 (N_259,N_42,N_116);
nand U260 (N_260,N_46,N_122);
and U261 (N_261,N_143,In_478);
xnor U262 (N_262,In_223,In_413);
or U263 (N_263,In_149,N_185);
nor U264 (N_264,N_142,In_394);
and U265 (N_265,N_117,In_203);
or U266 (N_266,N_186,In_144);
or U267 (N_267,In_451,N_135);
nor U268 (N_268,In_150,N_3);
or U269 (N_269,In_431,In_30);
nor U270 (N_270,In_153,In_432);
nor U271 (N_271,In_362,In_52);
nand U272 (N_272,N_128,N_124);
nor U273 (N_273,N_66,In_50);
or U274 (N_274,N_178,N_157);
nand U275 (N_275,N_129,N_187);
nor U276 (N_276,N_119,N_137);
nand U277 (N_277,In_387,In_105);
nor U278 (N_278,In_230,N_163);
or U279 (N_279,N_170,In_91);
and U280 (N_280,N_19,In_164);
and U281 (N_281,N_95,N_78);
nor U282 (N_282,In_463,In_479);
nand U283 (N_283,In_422,In_325);
nand U284 (N_284,In_4,In_29);
nor U285 (N_285,In_54,In_237);
or U286 (N_286,N_70,In_129);
or U287 (N_287,N_18,N_176);
and U288 (N_288,In_409,In_46);
nand U289 (N_289,In_110,In_293);
nor U290 (N_290,In_186,In_32);
and U291 (N_291,N_1,In_260);
nor U292 (N_292,N_147,N_100);
nor U293 (N_293,N_174,In_335);
or U294 (N_294,N_172,In_316);
and U295 (N_295,N_177,In_124);
nand U296 (N_296,In_59,N_134);
nor U297 (N_297,In_492,In_271);
and U298 (N_298,In_406,In_415);
nand U299 (N_299,N_169,In_499);
and U300 (N_300,N_212,N_93);
nand U301 (N_301,N_293,N_79);
and U302 (N_302,N_136,N_259);
nand U303 (N_303,N_112,In_306);
or U304 (N_304,In_33,N_123);
or U305 (N_305,N_266,N_74);
or U306 (N_306,N_239,N_222);
nor U307 (N_307,N_188,N_269);
nor U308 (N_308,N_224,In_486);
nor U309 (N_309,In_477,N_244);
nand U310 (N_310,N_216,N_284);
nor U311 (N_311,N_260,N_211);
xor U312 (N_312,N_197,N_37);
and U313 (N_313,N_273,N_227);
or U314 (N_314,N_8,N_287);
or U315 (N_315,N_274,In_264);
or U316 (N_316,N_245,In_183);
nand U317 (N_317,N_217,N_258);
and U318 (N_318,In_43,N_246);
nand U319 (N_319,In_475,N_182);
or U320 (N_320,N_202,N_192);
and U321 (N_321,In_458,N_256);
xor U322 (N_322,N_231,N_153);
nand U323 (N_323,N_241,In_356);
nor U324 (N_324,In_211,N_219);
nand U325 (N_325,N_209,N_220);
and U326 (N_326,N_233,N_263);
nor U327 (N_327,N_16,N_149);
and U328 (N_328,N_230,In_380);
or U329 (N_329,N_236,In_40);
nor U330 (N_330,N_111,N_120);
and U331 (N_331,N_248,N_282);
nor U332 (N_332,N_250,In_255);
nand U333 (N_333,In_252,In_193);
and U334 (N_334,N_226,In_270);
and U335 (N_335,N_270,N_291);
nor U336 (N_336,N_204,N_275);
nand U337 (N_337,N_249,N_272);
nand U338 (N_338,N_103,N_237);
nor U339 (N_339,N_110,In_473);
nor U340 (N_340,N_229,N_208);
and U341 (N_341,N_189,In_65);
or U342 (N_342,N_40,N_207);
nor U343 (N_343,N_290,N_125);
nand U344 (N_344,In_408,N_195);
or U345 (N_345,N_265,In_235);
or U346 (N_346,In_72,In_109);
and U347 (N_347,N_181,N_179);
or U348 (N_348,N_296,N_251);
and U349 (N_349,In_428,In_123);
or U350 (N_350,N_148,N_289);
nor U351 (N_351,N_198,N_299);
nand U352 (N_352,N_280,In_311);
or U353 (N_353,In_0,N_223);
and U354 (N_354,N_279,In_435);
nand U355 (N_355,N_221,N_255);
and U356 (N_356,N_286,In_350);
or U357 (N_357,N_206,In_64);
nand U358 (N_358,N_295,In_441);
nand U359 (N_359,N_281,In_74);
nand U360 (N_360,In_381,N_159);
nand U361 (N_361,N_193,N_161);
nand U362 (N_362,N_292,N_201);
or U363 (N_363,N_91,N_264);
nand U364 (N_364,N_200,N_225);
or U365 (N_365,In_173,N_288);
and U366 (N_366,N_139,N_294);
nand U367 (N_367,In_56,In_8);
nand U368 (N_368,N_285,N_126);
and U369 (N_369,In_199,N_210);
nor U370 (N_370,N_297,N_121);
nand U371 (N_371,N_214,N_240);
nor U372 (N_372,N_190,N_238);
nand U373 (N_373,In_15,N_277);
or U374 (N_374,N_162,N_253);
nor U375 (N_375,N_261,N_138);
nand U376 (N_376,In_181,In_26);
nor U377 (N_377,N_267,In_111);
or U378 (N_378,In_300,N_108);
nor U379 (N_379,In_337,N_89);
or U380 (N_380,In_112,In_346);
nand U381 (N_381,N_234,N_271);
or U382 (N_382,N_243,N_268);
nand U383 (N_383,In_369,N_102);
nor U384 (N_384,N_276,N_164);
nand U385 (N_385,In_218,In_39);
and U386 (N_386,N_242,N_254);
or U387 (N_387,In_324,N_54);
and U388 (N_388,N_278,N_257);
nand U389 (N_389,N_262,N_283);
or U390 (N_390,In_175,N_215);
nor U391 (N_391,N_228,In_246);
nand U392 (N_392,N_196,In_34);
and U393 (N_393,N_232,N_235);
or U394 (N_394,N_298,N_145);
and U395 (N_395,N_205,In_294);
and U396 (N_396,N_203,N_252);
nor U397 (N_397,N_247,N_213);
nor U398 (N_398,N_218,In_141);
or U399 (N_399,In_174,N_21);
and U400 (N_400,N_369,N_389);
nor U401 (N_401,N_323,N_325);
or U402 (N_402,N_349,N_339);
nor U403 (N_403,N_322,N_351);
and U404 (N_404,N_347,N_340);
and U405 (N_405,N_365,N_375);
or U406 (N_406,N_303,N_355);
or U407 (N_407,N_309,N_314);
and U408 (N_408,N_346,N_376);
or U409 (N_409,N_358,N_345);
nand U410 (N_410,N_396,N_390);
nand U411 (N_411,N_301,N_378);
nand U412 (N_412,N_366,N_367);
nor U413 (N_413,N_385,N_332);
nand U414 (N_414,N_321,N_399);
nor U415 (N_415,N_310,N_328);
and U416 (N_416,N_320,N_383);
or U417 (N_417,N_344,N_379);
nor U418 (N_418,N_373,N_336);
nor U419 (N_419,N_387,N_391);
and U420 (N_420,N_352,N_329);
nand U421 (N_421,N_317,N_337);
or U422 (N_422,N_398,N_362);
and U423 (N_423,N_393,N_392);
nor U424 (N_424,N_359,N_395);
nor U425 (N_425,N_304,N_394);
and U426 (N_426,N_316,N_350);
nand U427 (N_427,N_335,N_333);
nand U428 (N_428,N_312,N_327);
or U429 (N_429,N_372,N_308);
nand U430 (N_430,N_324,N_311);
nor U431 (N_431,N_377,N_364);
or U432 (N_432,N_305,N_371);
or U433 (N_433,N_313,N_300);
or U434 (N_434,N_348,N_397);
or U435 (N_435,N_381,N_343);
nand U436 (N_436,N_334,N_338);
and U437 (N_437,N_382,N_363);
and U438 (N_438,N_319,N_357);
or U439 (N_439,N_368,N_360);
nor U440 (N_440,N_330,N_315);
or U441 (N_441,N_384,N_341);
or U442 (N_442,N_374,N_388);
nand U443 (N_443,N_370,N_354);
or U444 (N_444,N_380,N_318);
or U445 (N_445,N_331,N_342);
nor U446 (N_446,N_356,N_361);
or U447 (N_447,N_326,N_306);
and U448 (N_448,N_353,N_307);
or U449 (N_449,N_386,N_302);
or U450 (N_450,N_357,N_312);
nand U451 (N_451,N_395,N_360);
and U452 (N_452,N_328,N_365);
or U453 (N_453,N_377,N_305);
nand U454 (N_454,N_390,N_395);
and U455 (N_455,N_377,N_331);
nor U456 (N_456,N_376,N_331);
nor U457 (N_457,N_347,N_383);
nand U458 (N_458,N_382,N_316);
nor U459 (N_459,N_373,N_375);
nand U460 (N_460,N_397,N_342);
or U461 (N_461,N_393,N_347);
and U462 (N_462,N_306,N_334);
nand U463 (N_463,N_353,N_369);
nor U464 (N_464,N_337,N_332);
and U465 (N_465,N_343,N_326);
and U466 (N_466,N_308,N_371);
or U467 (N_467,N_372,N_329);
or U468 (N_468,N_363,N_384);
or U469 (N_469,N_330,N_345);
xor U470 (N_470,N_300,N_351);
nor U471 (N_471,N_302,N_307);
and U472 (N_472,N_310,N_313);
nor U473 (N_473,N_390,N_372);
and U474 (N_474,N_378,N_392);
or U475 (N_475,N_350,N_340);
and U476 (N_476,N_314,N_375);
or U477 (N_477,N_340,N_331);
xnor U478 (N_478,N_372,N_373);
nand U479 (N_479,N_329,N_381);
nor U480 (N_480,N_361,N_384);
nor U481 (N_481,N_364,N_315);
nor U482 (N_482,N_332,N_356);
nor U483 (N_483,N_324,N_393);
nor U484 (N_484,N_372,N_364);
or U485 (N_485,N_337,N_381);
or U486 (N_486,N_363,N_349);
nor U487 (N_487,N_328,N_301);
or U488 (N_488,N_383,N_353);
and U489 (N_489,N_319,N_395);
or U490 (N_490,N_361,N_307);
nor U491 (N_491,N_359,N_310);
xor U492 (N_492,N_331,N_310);
and U493 (N_493,N_317,N_395);
nor U494 (N_494,N_311,N_374);
nand U495 (N_495,N_307,N_339);
and U496 (N_496,N_334,N_341);
and U497 (N_497,N_326,N_371);
or U498 (N_498,N_335,N_354);
and U499 (N_499,N_345,N_368);
nor U500 (N_500,N_405,N_498);
nand U501 (N_501,N_471,N_472);
nand U502 (N_502,N_499,N_421);
and U503 (N_503,N_439,N_441);
and U504 (N_504,N_443,N_455);
or U505 (N_505,N_464,N_489);
nand U506 (N_506,N_480,N_424);
or U507 (N_507,N_423,N_478);
nor U508 (N_508,N_451,N_409);
nor U509 (N_509,N_414,N_481);
and U510 (N_510,N_415,N_461);
nand U511 (N_511,N_442,N_486);
nand U512 (N_512,N_452,N_495);
nor U513 (N_513,N_496,N_422);
and U514 (N_514,N_402,N_408);
and U515 (N_515,N_473,N_497);
nor U516 (N_516,N_417,N_406);
or U517 (N_517,N_411,N_490);
and U518 (N_518,N_429,N_447);
and U519 (N_519,N_494,N_448);
nand U520 (N_520,N_419,N_413);
nor U521 (N_521,N_400,N_436);
or U522 (N_522,N_410,N_462);
nand U523 (N_523,N_469,N_432);
nor U524 (N_524,N_468,N_460);
or U525 (N_525,N_482,N_427);
nor U526 (N_526,N_449,N_418);
or U527 (N_527,N_463,N_456);
or U528 (N_528,N_437,N_433);
nand U529 (N_529,N_483,N_475);
or U530 (N_530,N_431,N_416);
nand U531 (N_531,N_479,N_493);
and U532 (N_532,N_457,N_474);
or U533 (N_533,N_444,N_420);
or U534 (N_534,N_467,N_434);
nand U535 (N_535,N_454,N_458);
nor U536 (N_536,N_440,N_450);
nand U537 (N_537,N_446,N_428);
nor U538 (N_538,N_435,N_459);
nor U539 (N_539,N_477,N_487);
nand U540 (N_540,N_430,N_412);
or U541 (N_541,N_470,N_426);
and U542 (N_542,N_403,N_476);
nor U543 (N_543,N_425,N_466);
nor U544 (N_544,N_438,N_488);
or U545 (N_545,N_492,N_491);
nor U546 (N_546,N_445,N_484);
and U547 (N_547,N_453,N_407);
or U548 (N_548,N_465,N_404);
and U549 (N_549,N_485,N_401);
nor U550 (N_550,N_437,N_421);
nor U551 (N_551,N_459,N_444);
nand U552 (N_552,N_497,N_494);
nor U553 (N_553,N_456,N_431);
nor U554 (N_554,N_427,N_464);
or U555 (N_555,N_446,N_489);
nand U556 (N_556,N_446,N_419);
nor U557 (N_557,N_434,N_494);
and U558 (N_558,N_472,N_422);
and U559 (N_559,N_415,N_437);
and U560 (N_560,N_453,N_475);
or U561 (N_561,N_490,N_456);
nor U562 (N_562,N_419,N_421);
nand U563 (N_563,N_454,N_430);
or U564 (N_564,N_463,N_482);
nor U565 (N_565,N_467,N_406);
and U566 (N_566,N_401,N_436);
or U567 (N_567,N_482,N_440);
nor U568 (N_568,N_494,N_450);
and U569 (N_569,N_455,N_401);
nand U570 (N_570,N_467,N_471);
nor U571 (N_571,N_489,N_407);
and U572 (N_572,N_465,N_493);
nand U573 (N_573,N_457,N_482);
and U574 (N_574,N_416,N_475);
nand U575 (N_575,N_446,N_414);
nor U576 (N_576,N_462,N_492);
and U577 (N_577,N_492,N_478);
or U578 (N_578,N_474,N_459);
xnor U579 (N_579,N_482,N_484);
and U580 (N_580,N_476,N_498);
or U581 (N_581,N_409,N_408);
nor U582 (N_582,N_429,N_448);
and U583 (N_583,N_483,N_463);
and U584 (N_584,N_413,N_475);
nor U585 (N_585,N_403,N_480);
nand U586 (N_586,N_421,N_480);
nor U587 (N_587,N_451,N_484);
nand U588 (N_588,N_415,N_484);
nor U589 (N_589,N_495,N_472);
nand U590 (N_590,N_491,N_457);
nand U591 (N_591,N_487,N_476);
nor U592 (N_592,N_413,N_409);
or U593 (N_593,N_482,N_408);
nand U594 (N_594,N_472,N_451);
or U595 (N_595,N_435,N_487);
and U596 (N_596,N_452,N_443);
or U597 (N_597,N_404,N_474);
and U598 (N_598,N_401,N_477);
nand U599 (N_599,N_463,N_425);
and U600 (N_600,N_527,N_548);
or U601 (N_601,N_576,N_561);
or U602 (N_602,N_547,N_594);
nand U603 (N_603,N_535,N_539);
nor U604 (N_604,N_532,N_560);
or U605 (N_605,N_559,N_562);
or U606 (N_606,N_578,N_529);
and U607 (N_607,N_517,N_569);
nand U608 (N_608,N_508,N_598);
or U609 (N_609,N_525,N_550);
or U610 (N_610,N_597,N_530);
nor U611 (N_611,N_566,N_564);
and U612 (N_612,N_556,N_540);
nand U613 (N_613,N_511,N_520);
or U614 (N_614,N_509,N_533);
and U615 (N_615,N_510,N_582);
or U616 (N_616,N_558,N_596);
and U617 (N_617,N_586,N_542);
and U618 (N_618,N_500,N_568);
nor U619 (N_619,N_552,N_574);
nor U620 (N_620,N_524,N_577);
nand U621 (N_621,N_593,N_573);
nand U622 (N_622,N_567,N_504);
nand U623 (N_623,N_595,N_544);
nand U624 (N_624,N_528,N_503);
nand U625 (N_625,N_543,N_534);
or U626 (N_626,N_522,N_521);
or U627 (N_627,N_575,N_589);
nor U628 (N_628,N_591,N_515);
or U629 (N_629,N_579,N_537);
or U630 (N_630,N_565,N_587);
or U631 (N_631,N_557,N_505);
nand U632 (N_632,N_536,N_507);
and U633 (N_633,N_580,N_553);
nand U634 (N_634,N_581,N_555);
nor U635 (N_635,N_523,N_554);
nor U636 (N_636,N_563,N_599);
nor U637 (N_637,N_502,N_585);
nor U638 (N_638,N_538,N_583);
or U639 (N_639,N_519,N_571);
xnor U640 (N_640,N_545,N_584);
nor U641 (N_641,N_514,N_572);
and U642 (N_642,N_506,N_592);
nand U643 (N_643,N_541,N_513);
nand U644 (N_644,N_501,N_516);
or U645 (N_645,N_588,N_549);
and U646 (N_646,N_590,N_518);
nand U647 (N_647,N_570,N_551);
or U648 (N_648,N_512,N_531);
or U649 (N_649,N_546,N_526);
and U650 (N_650,N_558,N_554);
nor U651 (N_651,N_595,N_555);
and U652 (N_652,N_564,N_509);
nand U653 (N_653,N_575,N_567);
xnor U654 (N_654,N_526,N_582);
and U655 (N_655,N_523,N_575);
nand U656 (N_656,N_537,N_593);
nand U657 (N_657,N_564,N_505);
nand U658 (N_658,N_525,N_537);
nor U659 (N_659,N_509,N_594);
nand U660 (N_660,N_578,N_583);
nor U661 (N_661,N_575,N_537);
or U662 (N_662,N_532,N_589);
and U663 (N_663,N_531,N_525);
or U664 (N_664,N_562,N_582);
and U665 (N_665,N_574,N_504);
nand U666 (N_666,N_518,N_521);
nand U667 (N_667,N_565,N_594);
and U668 (N_668,N_564,N_569);
and U669 (N_669,N_541,N_579);
nand U670 (N_670,N_537,N_530);
or U671 (N_671,N_553,N_512);
nand U672 (N_672,N_551,N_532);
nand U673 (N_673,N_511,N_533);
nand U674 (N_674,N_544,N_577);
nand U675 (N_675,N_543,N_501);
nor U676 (N_676,N_550,N_578);
nand U677 (N_677,N_567,N_594);
nor U678 (N_678,N_551,N_556);
or U679 (N_679,N_509,N_599);
and U680 (N_680,N_528,N_572);
or U681 (N_681,N_509,N_585);
and U682 (N_682,N_516,N_587);
xor U683 (N_683,N_591,N_559);
or U684 (N_684,N_528,N_546);
nand U685 (N_685,N_510,N_521);
and U686 (N_686,N_556,N_532);
and U687 (N_687,N_517,N_524);
or U688 (N_688,N_582,N_593);
or U689 (N_689,N_508,N_599);
or U690 (N_690,N_536,N_517);
nor U691 (N_691,N_552,N_550);
and U692 (N_692,N_514,N_525);
nand U693 (N_693,N_517,N_587);
or U694 (N_694,N_552,N_560);
or U695 (N_695,N_583,N_524);
nor U696 (N_696,N_548,N_532);
or U697 (N_697,N_544,N_549);
or U698 (N_698,N_564,N_526);
and U699 (N_699,N_530,N_551);
nand U700 (N_700,N_600,N_661);
or U701 (N_701,N_682,N_616);
or U702 (N_702,N_633,N_612);
or U703 (N_703,N_670,N_668);
nand U704 (N_704,N_698,N_692);
nor U705 (N_705,N_699,N_662);
nor U706 (N_706,N_677,N_675);
nor U707 (N_707,N_669,N_658);
nand U708 (N_708,N_644,N_613);
nor U709 (N_709,N_602,N_642);
nand U710 (N_710,N_623,N_618);
nand U711 (N_711,N_672,N_673);
nand U712 (N_712,N_632,N_653);
nand U713 (N_713,N_663,N_657);
or U714 (N_714,N_652,N_649);
nor U715 (N_715,N_637,N_606);
nor U716 (N_716,N_655,N_671);
nand U717 (N_717,N_650,N_608);
and U718 (N_718,N_689,N_695);
nand U719 (N_719,N_611,N_629);
nand U720 (N_720,N_683,N_610);
or U721 (N_721,N_605,N_627);
or U722 (N_722,N_686,N_656);
and U723 (N_723,N_609,N_691);
nor U724 (N_724,N_647,N_676);
and U725 (N_725,N_604,N_681);
and U726 (N_726,N_694,N_638);
and U727 (N_727,N_628,N_641);
nand U728 (N_728,N_690,N_666);
nand U729 (N_729,N_687,N_680);
or U730 (N_730,N_624,N_617);
and U731 (N_731,N_667,N_601);
nor U732 (N_732,N_665,N_648);
nor U733 (N_733,N_693,N_626);
nand U734 (N_734,N_660,N_651);
and U735 (N_735,N_640,N_621);
and U736 (N_736,N_631,N_679);
nand U737 (N_737,N_630,N_659);
or U738 (N_738,N_615,N_619);
nor U739 (N_739,N_645,N_639);
nand U740 (N_740,N_635,N_603);
or U741 (N_741,N_688,N_636);
nor U742 (N_742,N_646,N_625);
nor U743 (N_743,N_684,N_685);
or U744 (N_744,N_643,N_614);
or U745 (N_745,N_654,N_607);
nor U746 (N_746,N_697,N_696);
or U747 (N_747,N_620,N_664);
nand U748 (N_748,N_674,N_634);
xnor U749 (N_749,N_622,N_678);
nand U750 (N_750,N_604,N_620);
nand U751 (N_751,N_615,N_670);
nor U752 (N_752,N_648,N_608);
nand U753 (N_753,N_617,N_600);
or U754 (N_754,N_696,N_603);
or U755 (N_755,N_634,N_673);
and U756 (N_756,N_615,N_616);
or U757 (N_757,N_602,N_604);
nor U758 (N_758,N_682,N_636);
and U759 (N_759,N_620,N_649);
and U760 (N_760,N_619,N_635);
and U761 (N_761,N_695,N_684);
or U762 (N_762,N_605,N_629);
nand U763 (N_763,N_629,N_610);
or U764 (N_764,N_680,N_604);
and U765 (N_765,N_675,N_611);
nand U766 (N_766,N_698,N_680);
and U767 (N_767,N_672,N_654);
nor U768 (N_768,N_640,N_606);
nor U769 (N_769,N_611,N_665);
and U770 (N_770,N_657,N_654);
nand U771 (N_771,N_619,N_676);
or U772 (N_772,N_679,N_689);
nand U773 (N_773,N_659,N_684);
nand U774 (N_774,N_678,N_669);
and U775 (N_775,N_635,N_690);
or U776 (N_776,N_649,N_646);
nand U777 (N_777,N_617,N_670);
and U778 (N_778,N_615,N_671);
or U779 (N_779,N_666,N_645);
nor U780 (N_780,N_643,N_609);
or U781 (N_781,N_619,N_649);
nand U782 (N_782,N_679,N_622);
or U783 (N_783,N_691,N_678);
nor U784 (N_784,N_618,N_698);
nand U785 (N_785,N_619,N_678);
nand U786 (N_786,N_640,N_631);
nor U787 (N_787,N_694,N_683);
nand U788 (N_788,N_657,N_653);
and U789 (N_789,N_605,N_683);
nand U790 (N_790,N_642,N_609);
nand U791 (N_791,N_637,N_640);
and U792 (N_792,N_648,N_699);
and U793 (N_793,N_609,N_656);
nor U794 (N_794,N_603,N_692);
and U795 (N_795,N_699,N_687);
nor U796 (N_796,N_639,N_665);
and U797 (N_797,N_698,N_603);
or U798 (N_798,N_652,N_696);
and U799 (N_799,N_607,N_670);
or U800 (N_800,N_777,N_784);
and U801 (N_801,N_728,N_778);
nor U802 (N_802,N_701,N_758);
nor U803 (N_803,N_755,N_790);
nand U804 (N_804,N_732,N_773);
or U805 (N_805,N_786,N_704);
nand U806 (N_806,N_779,N_725);
nand U807 (N_807,N_723,N_757);
and U808 (N_808,N_737,N_775);
or U809 (N_809,N_745,N_705);
nor U810 (N_810,N_716,N_767);
and U811 (N_811,N_799,N_749);
nor U812 (N_812,N_709,N_764);
nand U813 (N_813,N_707,N_711);
nand U814 (N_814,N_715,N_702);
xor U815 (N_815,N_769,N_742);
and U816 (N_816,N_798,N_706);
and U817 (N_817,N_730,N_751);
and U818 (N_818,N_700,N_797);
or U819 (N_819,N_792,N_753);
or U820 (N_820,N_756,N_774);
nand U821 (N_821,N_771,N_789);
or U822 (N_822,N_794,N_744);
nor U823 (N_823,N_720,N_772);
or U824 (N_824,N_785,N_729);
or U825 (N_825,N_741,N_776);
nor U826 (N_826,N_746,N_765);
nor U827 (N_827,N_788,N_736);
and U828 (N_828,N_735,N_748);
or U829 (N_829,N_717,N_762);
and U830 (N_830,N_759,N_743);
nand U831 (N_831,N_733,N_703);
nor U832 (N_832,N_740,N_710);
nor U833 (N_833,N_752,N_718);
or U834 (N_834,N_721,N_747);
nor U835 (N_835,N_712,N_787);
and U836 (N_836,N_761,N_726);
and U837 (N_837,N_782,N_768);
and U838 (N_838,N_754,N_766);
nor U839 (N_839,N_731,N_724);
or U840 (N_840,N_738,N_770);
xor U841 (N_841,N_713,N_734);
and U842 (N_842,N_781,N_722);
nand U843 (N_843,N_714,N_780);
nor U844 (N_844,N_719,N_763);
and U845 (N_845,N_739,N_793);
nand U846 (N_846,N_750,N_708);
or U847 (N_847,N_795,N_760);
and U848 (N_848,N_727,N_791);
and U849 (N_849,N_783,N_796);
and U850 (N_850,N_730,N_752);
or U851 (N_851,N_713,N_717);
and U852 (N_852,N_743,N_700);
nor U853 (N_853,N_748,N_773);
nand U854 (N_854,N_799,N_782);
nand U855 (N_855,N_772,N_746);
and U856 (N_856,N_792,N_762);
nor U857 (N_857,N_778,N_719);
xor U858 (N_858,N_741,N_761);
or U859 (N_859,N_760,N_754);
nor U860 (N_860,N_717,N_751);
and U861 (N_861,N_749,N_750);
nand U862 (N_862,N_717,N_741);
or U863 (N_863,N_753,N_789);
nand U864 (N_864,N_796,N_754);
nand U865 (N_865,N_701,N_776);
and U866 (N_866,N_792,N_749);
or U867 (N_867,N_742,N_786);
nor U868 (N_868,N_770,N_731);
and U869 (N_869,N_752,N_783);
or U870 (N_870,N_773,N_752);
nor U871 (N_871,N_752,N_784);
or U872 (N_872,N_781,N_728);
or U873 (N_873,N_745,N_709);
nand U874 (N_874,N_791,N_772);
or U875 (N_875,N_753,N_704);
nand U876 (N_876,N_786,N_711);
nand U877 (N_877,N_770,N_709);
nor U878 (N_878,N_769,N_795);
or U879 (N_879,N_749,N_759);
nor U880 (N_880,N_797,N_708);
nor U881 (N_881,N_734,N_740);
nand U882 (N_882,N_773,N_730);
nand U883 (N_883,N_729,N_719);
or U884 (N_884,N_763,N_705);
or U885 (N_885,N_768,N_702);
or U886 (N_886,N_786,N_724);
nor U887 (N_887,N_702,N_700);
and U888 (N_888,N_731,N_726);
or U889 (N_889,N_795,N_744);
nand U890 (N_890,N_720,N_754);
xnor U891 (N_891,N_793,N_763);
nor U892 (N_892,N_731,N_701);
or U893 (N_893,N_746,N_713);
and U894 (N_894,N_730,N_734);
nand U895 (N_895,N_711,N_793);
nand U896 (N_896,N_723,N_769);
or U897 (N_897,N_750,N_766);
nor U898 (N_898,N_785,N_737);
nand U899 (N_899,N_706,N_710);
nand U900 (N_900,N_856,N_827);
or U901 (N_901,N_828,N_838);
and U902 (N_902,N_874,N_890);
nand U903 (N_903,N_814,N_893);
and U904 (N_904,N_883,N_871);
and U905 (N_905,N_868,N_832);
or U906 (N_906,N_858,N_831);
nor U907 (N_907,N_852,N_899);
nand U908 (N_908,N_864,N_857);
nor U909 (N_909,N_891,N_892);
nand U910 (N_910,N_807,N_878);
nand U911 (N_911,N_805,N_820);
nor U912 (N_912,N_895,N_865);
nor U913 (N_913,N_803,N_817);
nor U914 (N_914,N_833,N_861);
nor U915 (N_915,N_835,N_888);
or U916 (N_916,N_896,N_885);
and U917 (N_917,N_877,N_882);
nor U918 (N_918,N_897,N_848);
nand U919 (N_919,N_845,N_847);
nor U920 (N_920,N_843,N_819);
nand U921 (N_921,N_894,N_886);
nand U922 (N_922,N_826,N_859);
or U923 (N_923,N_816,N_866);
or U924 (N_924,N_806,N_846);
or U925 (N_925,N_839,N_800);
or U926 (N_926,N_810,N_811);
nand U927 (N_927,N_818,N_823);
nand U928 (N_928,N_824,N_830);
nand U929 (N_929,N_837,N_862);
nand U930 (N_930,N_880,N_841);
or U931 (N_931,N_822,N_867);
and U932 (N_932,N_898,N_889);
nor U933 (N_933,N_887,N_801);
or U934 (N_934,N_863,N_812);
nand U935 (N_935,N_840,N_849);
nor U936 (N_936,N_869,N_850);
or U937 (N_937,N_870,N_829);
nor U938 (N_938,N_813,N_853);
nand U939 (N_939,N_854,N_876);
nor U940 (N_940,N_834,N_879);
and U941 (N_941,N_851,N_881);
nand U942 (N_942,N_821,N_836);
nand U943 (N_943,N_809,N_872);
nand U944 (N_944,N_804,N_808);
nor U945 (N_945,N_802,N_875);
nand U946 (N_946,N_815,N_844);
and U947 (N_947,N_884,N_825);
nor U948 (N_948,N_842,N_873);
nor U949 (N_949,N_860,N_855);
nand U950 (N_950,N_880,N_858);
nand U951 (N_951,N_837,N_881);
and U952 (N_952,N_890,N_827);
nand U953 (N_953,N_827,N_875);
and U954 (N_954,N_829,N_882);
or U955 (N_955,N_887,N_878);
and U956 (N_956,N_800,N_803);
nand U957 (N_957,N_859,N_811);
nand U958 (N_958,N_881,N_832);
or U959 (N_959,N_849,N_829);
or U960 (N_960,N_855,N_835);
or U961 (N_961,N_847,N_884);
or U962 (N_962,N_814,N_877);
nand U963 (N_963,N_801,N_881);
or U964 (N_964,N_868,N_814);
nand U965 (N_965,N_874,N_826);
nor U966 (N_966,N_892,N_876);
nand U967 (N_967,N_858,N_801);
and U968 (N_968,N_879,N_871);
or U969 (N_969,N_870,N_885);
and U970 (N_970,N_859,N_804);
nor U971 (N_971,N_847,N_880);
or U972 (N_972,N_812,N_872);
nand U973 (N_973,N_860,N_862);
nand U974 (N_974,N_819,N_854);
nand U975 (N_975,N_876,N_897);
nor U976 (N_976,N_818,N_858);
nand U977 (N_977,N_876,N_874);
nor U978 (N_978,N_801,N_894);
xnor U979 (N_979,N_822,N_862);
nor U980 (N_980,N_854,N_887);
nor U981 (N_981,N_892,N_826);
nor U982 (N_982,N_885,N_813);
nor U983 (N_983,N_871,N_868);
nand U984 (N_984,N_870,N_830);
and U985 (N_985,N_839,N_803);
nor U986 (N_986,N_872,N_863);
nor U987 (N_987,N_869,N_884);
nor U988 (N_988,N_815,N_855);
or U989 (N_989,N_876,N_879);
nand U990 (N_990,N_804,N_895);
or U991 (N_991,N_870,N_872);
nand U992 (N_992,N_879,N_878);
nor U993 (N_993,N_896,N_833);
nor U994 (N_994,N_815,N_828);
or U995 (N_995,N_835,N_813);
and U996 (N_996,N_876,N_859);
nand U997 (N_997,N_858,N_824);
nand U998 (N_998,N_892,N_824);
or U999 (N_999,N_856,N_848);
nand U1000 (N_1000,N_960,N_901);
and U1001 (N_1001,N_965,N_969);
or U1002 (N_1002,N_913,N_926);
nand U1003 (N_1003,N_944,N_959);
or U1004 (N_1004,N_910,N_939);
nor U1005 (N_1005,N_957,N_984);
or U1006 (N_1006,N_968,N_986);
and U1007 (N_1007,N_923,N_963);
nor U1008 (N_1008,N_948,N_935);
and U1009 (N_1009,N_993,N_932);
nand U1010 (N_1010,N_976,N_927);
nor U1011 (N_1011,N_915,N_919);
nand U1012 (N_1012,N_918,N_978);
nor U1013 (N_1013,N_983,N_995);
or U1014 (N_1014,N_987,N_991);
and U1015 (N_1015,N_972,N_922);
nand U1016 (N_1016,N_900,N_999);
and U1017 (N_1017,N_950,N_949);
nand U1018 (N_1018,N_912,N_967);
nor U1019 (N_1019,N_981,N_994);
nor U1020 (N_1020,N_996,N_952);
nor U1021 (N_1021,N_936,N_956);
and U1022 (N_1022,N_907,N_992);
and U1023 (N_1023,N_917,N_982);
and U1024 (N_1024,N_941,N_966);
nand U1025 (N_1025,N_925,N_971);
nand U1026 (N_1026,N_903,N_938);
nor U1027 (N_1027,N_951,N_914);
nor U1028 (N_1028,N_998,N_962);
nand U1029 (N_1029,N_979,N_947);
or U1030 (N_1030,N_943,N_911);
nand U1031 (N_1031,N_988,N_975);
and U1032 (N_1032,N_933,N_920);
or U1033 (N_1033,N_940,N_989);
nor U1034 (N_1034,N_985,N_990);
and U1035 (N_1035,N_953,N_928);
or U1036 (N_1036,N_924,N_906);
or U1037 (N_1037,N_902,N_997);
and U1038 (N_1038,N_945,N_973);
nand U1039 (N_1039,N_905,N_954);
and U1040 (N_1040,N_916,N_958);
or U1041 (N_1041,N_908,N_955);
and U1042 (N_1042,N_980,N_931);
and U1043 (N_1043,N_904,N_909);
or U1044 (N_1044,N_934,N_929);
or U1045 (N_1045,N_946,N_964);
nand U1046 (N_1046,N_942,N_977);
nor U1047 (N_1047,N_970,N_961);
and U1048 (N_1048,N_974,N_930);
and U1049 (N_1049,N_937,N_921);
and U1050 (N_1050,N_921,N_978);
nand U1051 (N_1051,N_909,N_932);
and U1052 (N_1052,N_939,N_913);
nand U1053 (N_1053,N_955,N_933);
or U1054 (N_1054,N_951,N_989);
nand U1055 (N_1055,N_973,N_963);
or U1056 (N_1056,N_962,N_990);
nor U1057 (N_1057,N_969,N_984);
nor U1058 (N_1058,N_996,N_910);
nand U1059 (N_1059,N_989,N_919);
nor U1060 (N_1060,N_947,N_904);
nor U1061 (N_1061,N_972,N_973);
nand U1062 (N_1062,N_945,N_908);
and U1063 (N_1063,N_961,N_944);
and U1064 (N_1064,N_930,N_967);
or U1065 (N_1065,N_944,N_927);
nor U1066 (N_1066,N_910,N_930);
nor U1067 (N_1067,N_963,N_943);
nand U1068 (N_1068,N_964,N_951);
nand U1069 (N_1069,N_970,N_965);
and U1070 (N_1070,N_937,N_994);
nor U1071 (N_1071,N_903,N_994);
nand U1072 (N_1072,N_964,N_913);
and U1073 (N_1073,N_919,N_978);
or U1074 (N_1074,N_994,N_991);
nand U1075 (N_1075,N_995,N_902);
nand U1076 (N_1076,N_975,N_932);
and U1077 (N_1077,N_967,N_924);
nand U1078 (N_1078,N_906,N_979);
or U1079 (N_1079,N_932,N_959);
and U1080 (N_1080,N_959,N_984);
or U1081 (N_1081,N_998,N_916);
and U1082 (N_1082,N_963,N_931);
nor U1083 (N_1083,N_956,N_918);
and U1084 (N_1084,N_983,N_926);
nor U1085 (N_1085,N_990,N_955);
nand U1086 (N_1086,N_952,N_991);
nor U1087 (N_1087,N_983,N_904);
nand U1088 (N_1088,N_937,N_951);
nand U1089 (N_1089,N_902,N_992);
xor U1090 (N_1090,N_950,N_929);
nand U1091 (N_1091,N_955,N_956);
nor U1092 (N_1092,N_954,N_985);
nand U1093 (N_1093,N_942,N_918);
and U1094 (N_1094,N_989,N_909);
nor U1095 (N_1095,N_995,N_985);
or U1096 (N_1096,N_910,N_926);
nand U1097 (N_1097,N_964,N_937);
or U1098 (N_1098,N_946,N_917);
nand U1099 (N_1099,N_929,N_958);
or U1100 (N_1100,N_1027,N_1012);
or U1101 (N_1101,N_1029,N_1082);
nor U1102 (N_1102,N_1023,N_1075);
nor U1103 (N_1103,N_1060,N_1033);
nor U1104 (N_1104,N_1045,N_1015);
or U1105 (N_1105,N_1031,N_1069);
nand U1106 (N_1106,N_1053,N_1013);
and U1107 (N_1107,N_1091,N_1003);
nand U1108 (N_1108,N_1042,N_1096);
nand U1109 (N_1109,N_1024,N_1004);
and U1110 (N_1110,N_1052,N_1065);
nand U1111 (N_1111,N_1057,N_1050);
or U1112 (N_1112,N_1051,N_1001);
nand U1113 (N_1113,N_1085,N_1080);
nand U1114 (N_1114,N_1047,N_1010);
nor U1115 (N_1115,N_1018,N_1098);
nand U1116 (N_1116,N_1084,N_1094);
and U1117 (N_1117,N_1068,N_1030);
and U1118 (N_1118,N_1067,N_1078);
nand U1119 (N_1119,N_1038,N_1046);
nand U1120 (N_1120,N_1016,N_1049);
or U1121 (N_1121,N_1092,N_1079);
or U1122 (N_1122,N_1086,N_1006);
and U1123 (N_1123,N_1021,N_1019);
and U1124 (N_1124,N_1037,N_1017);
or U1125 (N_1125,N_1055,N_1061);
or U1126 (N_1126,N_1041,N_1066);
nor U1127 (N_1127,N_1025,N_1077);
and U1128 (N_1128,N_1009,N_1090);
nand U1129 (N_1129,N_1054,N_1072);
nor U1130 (N_1130,N_1064,N_1056);
nand U1131 (N_1131,N_1040,N_1081);
or U1132 (N_1132,N_1028,N_1058);
or U1133 (N_1133,N_1022,N_1095);
nand U1134 (N_1134,N_1074,N_1048);
or U1135 (N_1135,N_1059,N_1076);
or U1136 (N_1136,N_1062,N_1000);
or U1137 (N_1137,N_1043,N_1087);
nor U1138 (N_1138,N_1007,N_1039);
nand U1139 (N_1139,N_1034,N_1035);
nor U1140 (N_1140,N_1036,N_1089);
or U1141 (N_1141,N_1002,N_1005);
or U1142 (N_1142,N_1097,N_1020);
or U1143 (N_1143,N_1014,N_1032);
nor U1144 (N_1144,N_1011,N_1093);
nor U1145 (N_1145,N_1026,N_1071);
or U1146 (N_1146,N_1088,N_1073);
and U1147 (N_1147,N_1044,N_1070);
or U1148 (N_1148,N_1083,N_1063);
nor U1149 (N_1149,N_1008,N_1099);
and U1150 (N_1150,N_1032,N_1034);
or U1151 (N_1151,N_1064,N_1033);
and U1152 (N_1152,N_1041,N_1062);
or U1153 (N_1153,N_1036,N_1027);
and U1154 (N_1154,N_1063,N_1097);
or U1155 (N_1155,N_1000,N_1035);
or U1156 (N_1156,N_1010,N_1011);
nor U1157 (N_1157,N_1005,N_1042);
and U1158 (N_1158,N_1085,N_1087);
and U1159 (N_1159,N_1051,N_1011);
and U1160 (N_1160,N_1066,N_1058);
nand U1161 (N_1161,N_1017,N_1005);
nor U1162 (N_1162,N_1025,N_1034);
nand U1163 (N_1163,N_1091,N_1039);
nor U1164 (N_1164,N_1080,N_1043);
nand U1165 (N_1165,N_1022,N_1045);
or U1166 (N_1166,N_1082,N_1002);
or U1167 (N_1167,N_1078,N_1088);
or U1168 (N_1168,N_1005,N_1024);
or U1169 (N_1169,N_1028,N_1017);
or U1170 (N_1170,N_1055,N_1080);
or U1171 (N_1171,N_1081,N_1033);
and U1172 (N_1172,N_1045,N_1001);
nand U1173 (N_1173,N_1084,N_1042);
or U1174 (N_1174,N_1062,N_1004);
nand U1175 (N_1175,N_1042,N_1068);
and U1176 (N_1176,N_1090,N_1097);
and U1177 (N_1177,N_1088,N_1013);
nand U1178 (N_1178,N_1090,N_1007);
or U1179 (N_1179,N_1053,N_1016);
nand U1180 (N_1180,N_1072,N_1001);
or U1181 (N_1181,N_1061,N_1051);
or U1182 (N_1182,N_1047,N_1051);
or U1183 (N_1183,N_1022,N_1072);
and U1184 (N_1184,N_1098,N_1010);
or U1185 (N_1185,N_1042,N_1024);
nor U1186 (N_1186,N_1022,N_1016);
or U1187 (N_1187,N_1071,N_1032);
nor U1188 (N_1188,N_1004,N_1053);
and U1189 (N_1189,N_1078,N_1021);
nor U1190 (N_1190,N_1017,N_1090);
nand U1191 (N_1191,N_1018,N_1075);
nor U1192 (N_1192,N_1071,N_1031);
or U1193 (N_1193,N_1018,N_1009);
or U1194 (N_1194,N_1020,N_1076);
nand U1195 (N_1195,N_1033,N_1065);
or U1196 (N_1196,N_1057,N_1068);
nor U1197 (N_1197,N_1031,N_1009);
or U1198 (N_1198,N_1083,N_1065);
or U1199 (N_1199,N_1012,N_1076);
or U1200 (N_1200,N_1131,N_1165);
and U1201 (N_1201,N_1188,N_1121);
or U1202 (N_1202,N_1197,N_1113);
and U1203 (N_1203,N_1190,N_1168);
nor U1204 (N_1204,N_1137,N_1193);
nor U1205 (N_1205,N_1186,N_1136);
or U1206 (N_1206,N_1112,N_1115);
or U1207 (N_1207,N_1175,N_1105);
and U1208 (N_1208,N_1125,N_1149);
and U1209 (N_1209,N_1152,N_1187);
nor U1210 (N_1210,N_1123,N_1104);
nand U1211 (N_1211,N_1183,N_1157);
nor U1212 (N_1212,N_1161,N_1130);
and U1213 (N_1213,N_1107,N_1138);
nand U1214 (N_1214,N_1103,N_1163);
nand U1215 (N_1215,N_1122,N_1118);
and U1216 (N_1216,N_1181,N_1153);
or U1217 (N_1217,N_1199,N_1182);
and U1218 (N_1218,N_1178,N_1184);
or U1219 (N_1219,N_1174,N_1134);
nand U1220 (N_1220,N_1155,N_1151);
and U1221 (N_1221,N_1129,N_1132);
nor U1222 (N_1222,N_1146,N_1198);
nor U1223 (N_1223,N_1158,N_1173);
and U1224 (N_1224,N_1189,N_1156);
nor U1225 (N_1225,N_1196,N_1106);
or U1226 (N_1226,N_1111,N_1170);
nor U1227 (N_1227,N_1191,N_1140);
nor U1228 (N_1228,N_1143,N_1119);
nor U1229 (N_1229,N_1126,N_1176);
nor U1230 (N_1230,N_1114,N_1172);
and U1231 (N_1231,N_1142,N_1164);
nor U1232 (N_1232,N_1150,N_1128);
and U1233 (N_1233,N_1100,N_1145);
and U1234 (N_1234,N_1133,N_1108);
or U1235 (N_1235,N_1166,N_1102);
nand U1236 (N_1236,N_1179,N_1110);
or U1237 (N_1237,N_1154,N_1177);
and U1238 (N_1238,N_1159,N_1160);
and U1239 (N_1239,N_1195,N_1141);
nor U1240 (N_1240,N_1135,N_1169);
or U1241 (N_1241,N_1180,N_1116);
nand U1242 (N_1242,N_1120,N_1139);
nand U1243 (N_1243,N_1192,N_1167);
and U1244 (N_1244,N_1101,N_1124);
and U1245 (N_1245,N_1194,N_1162);
nand U1246 (N_1246,N_1171,N_1148);
or U1247 (N_1247,N_1147,N_1144);
and U1248 (N_1248,N_1117,N_1109);
nor U1249 (N_1249,N_1127,N_1185);
nand U1250 (N_1250,N_1150,N_1168);
and U1251 (N_1251,N_1160,N_1118);
nor U1252 (N_1252,N_1132,N_1161);
or U1253 (N_1253,N_1112,N_1149);
and U1254 (N_1254,N_1151,N_1158);
nand U1255 (N_1255,N_1157,N_1135);
or U1256 (N_1256,N_1193,N_1145);
nand U1257 (N_1257,N_1171,N_1173);
and U1258 (N_1258,N_1119,N_1174);
nand U1259 (N_1259,N_1172,N_1126);
and U1260 (N_1260,N_1165,N_1102);
nand U1261 (N_1261,N_1114,N_1102);
or U1262 (N_1262,N_1137,N_1163);
or U1263 (N_1263,N_1176,N_1178);
nor U1264 (N_1264,N_1126,N_1150);
nand U1265 (N_1265,N_1183,N_1106);
nor U1266 (N_1266,N_1186,N_1129);
and U1267 (N_1267,N_1157,N_1192);
nor U1268 (N_1268,N_1148,N_1184);
and U1269 (N_1269,N_1114,N_1175);
nand U1270 (N_1270,N_1135,N_1180);
or U1271 (N_1271,N_1148,N_1120);
nor U1272 (N_1272,N_1176,N_1137);
xnor U1273 (N_1273,N_1126,N_1146);
nand U1274 (N_1274,N_1196,N_1133);
nor U1275 (N_1275,N_1166,N_1142);
and U1276 (N_1276,N_1109,N_1141);
nand U1277 (N_1277,N_1171,N_1130);
and U1278 (N_1278,N_1135,N_1182);
or U1279 (N_1279,N_1190,N_1102);
and U1280 (N_1280,N_1164,N_1123);
nor U1281 (N_1281,N_1138,N_1133);
nor U1282 (N_1282,N_1103,N_1107);
or U1283 (N_1283,N_1111,N_1182);
and U1284 (N_1284,N_1169,N_1137);
nor U1285 (N_1285,N_1182,N_1121);
nor U1286 (N_1286,N_1113,N_1124);
and U1287 (N_1287,N_1183,N_1197);
or U1288 (N_1288,N_1145,N_1142);
nand U1289 (N_1289,N_1189,N_1184);
nand U1290 (N_1290,N_1102,N_1175);
or U1291 (N_1291,N_1110,N_1187);
nand U1292 (N_1292,N_1111,N_1131);
or U1293 (N_1293,N_1152,N_1175);
or U1294 (N_1294,N_1185,N_1133);
or U1295 (N_1295,N_1195,N_1190);
or U1296 (N_1296,N_1175,N_1180);
and U1297 (N_1297,N_1114,N_1125);
and U1298 (N_1298,N_1145,N_1173);
and U1299 (N_1299,N_1103,N_1134);
or U1300 (N_1300,N_1290,N_1252);
nand U1301 (N_1301,N_1291,N_1215);
nand U1302 (N_1302,N_1247,N_1224);
nand U1303 (N_1303,N_1236,N_1238);
nand U1304 (N_1304,N_1268,N_1297);
or U1305 (N_1305,N_1285,N_1298);
or U1306 (N_1306,N_1280,N_1284);
nand U1307 (N_1307,N_1293,N_1286);
or U1308 (N_1308,N_1270,N_1275);
or U1309 (N_1309,N_1253,N_1226);
or U1310 (N_1310,N_1255,N_1289);
or U1311 (N_1311,N_1225,N_1204);
nor U1312 (N_1312,N_1230,N_1283);
or U1313 (N_1313,N_1211,N_1222);
or U1314 (N_1314,N_1243,N_1220);
nand U1315 (N_1315,N_1279,N_1228);
and U1316 (N_1316,N_1266,N_1241);
xor U1317 (N_1317,N_1223,N_1265);
nand U1318 (N_1318,N_1294,N_1209);
nor U1319 (N_1319,N_1276,N_1217);
nor U1320 (N_1320,N_1205,N_1299);
or U1321 (N_1321,N_1250,N_1260);
nor U1322 (N_1322,N_1256,N_1249);
and U1323 (N_1323,N_1259,N_1235);
or U1324 (N_1324,N_1254,N_1257);
nand U1325 (N_1325,N_1263,N_1203);
nor U1326 (N_1326,N_1231,N_1296);
nand U1327 (N_1327,N_1246,N_1269);
or U1328 (N_1328,N_1229,N_1262);
or U1329 (N_1329,N_1213,N_1245);
and U1330 (N_1330,N_1251,N_1248);
and U1331 (N_1331,N_1207,N_1277);
and U1332 (N_1332,N_1274,N_1281);
nand U1333 (N_1333,N_1233,N_1221);
and U1334 (N_1334,N_1295,N_1212);
nor U1335 (N_1335,N_1232,N_1282);
nand U1336 (N_1336,N_1210,N_1216);
nor U1337 (N_1337,N_1208,N_1234);
nand U1338 (N_1338,N_1239,N_1214);
nor U1339 (N_1339,N_1242,N_1272);
nor U1340 (N_1340,N_1227,N_1202);
nor U1341 (N_1341,N_1219,N_1288);
or U1342 (N_1342,N_1292,N_1278);
and U1343 (N_1343,N_1264,N_1267);
nand U1344 (N_1344,N_1200,N_1271);
nor U1345 (N_1345,N_1261,N_1240);
nand U1346 (N_1346,N_1287,N_1201);
nor U1347 (N_1347,N_1206,N_1258);
and U1348 (N_1348,N_1237,N_1218);
or U1349 (N_1349,N_1273,N_1244);
or U1350 (N_1350,N_1234,N_1268);
or U1351 (N_1351,N_1200,N_1247);
and U1352 (N_1352,N_1256,N_1229);
nand U1353 (N_1353,N_1236,N_1212);
and U1354 (N_1354,N_1249,N_1268);
nor U1355 (N_1355,N_1204,N_1289);
nand U1356 (N_1356,N_1282,N_1239);
nand U1357 (N_1357,N_1267,N_1298);
nor U1358 (N_1358,N_1233,N_1204);
nor U1359 (N_1359,N_1276,N_1236);
or U1360 (N_1360,N_1258,N_1296);
nor U1361 (N_1361,N_1219,N_1243);
and U1362 (N_1362,N_1203,N_1202);
nor U1363 (N_1363,N_1281,N_1267);
nor U1364 (N_1364,N_1226,N_1202);
and U1365 (N_1365,N_1212,N_1270);
nor U1366 (N_1366,N_1247,N_1217);
and U1367 (N_1367,N_1267,N_1250);
nor U1368 (N_1368,N_1239,N_1245);
nor U1369 (N_1369,N_1289,N_1249);
or U1370 (N_1370,N_1263,N_1260);
nor U1371 (N_1371,N_1202,N_1269);
nand U1372 (N_1372,N_1213,N_1263);
nor U1373 (N_1373,N_1289,N_1257);
and U1374 (N_1374,N_1259,N_1239);
or U1375 (N_1375,N_1259,N_1282);
and U1376 (N_1376,N_1244,N_1250);
and U1377 (N_1377,N_1204,N_1228);
nand U1378 (N_1378,N_1239,N_1226);
or U1379 (N_1379,N_1203,N_1204);
and U1380 (N_1380,N_1208,N_1223);
and U1381 (N_1381,N_1240,N_1211);
or U1382 (N_1382,N_1267,N_1240);
nor U1383 (N_1383,N_1246,N_1275);
and U1384 (N_1384,N_1210,N_1259);
or U1385 (N_1385,N_1293,N_1223);
and U1386 (N_1386,N_1200,N_1218);
or U1387 (N_1387,N_1297,N_1290);
nor U1388 (N_1388,N_1217,N_1254);
nand U1389 (N_1389,N_1253,N_1237);
nor U1390 (N_1390,N_1260,N_1274);
nor U1391 (N_1391,N_1234,N_1263);
and U1392 (N_1392,N_1218,N_1283);
nand U1393 (N_1393,N_1233,N_1299);
nor U1394 (N_1394,N_1255,N_1288);
nor U1395 (N_1395,N_1200,N_1275);
and U1396 (N_1396,N_1278,N_1208);
nor U1397 (N_1397,N_1214,N_1266);
nor U1398 (N_1398,N_1246,N_1298);
nand U1399 (N_1399,N_1228,N_1259);
or U1400 (N_1400,N_1366,N_1397);
nand U1401 (N_1401,N_1322,N_1377);
nor U1402 (N_1402,N_1302,N_1354);
or U1403 (N_1403,N_1363,N_1328);
or U1404 (N_1404,N_1333,N_1323);
nor U1405 (N_1405,N_1306,N_1332);
nor U1406 (N_1406,N_1337,N_1392);
or U1407 (N_1407,N_1399,N_1360);
nand U1408 (N_1408,N_1334,N_1324);
or U1409 (N_1409,N_1396,N_1380);
or U1410 (N_1410,N_1338,N_1342);
or U1411 (N_1411,N_1339,N_1387);
nor U1412 (N_1412,N_1336,N_1316);
and U1413 (N_1413,N_1378,N_1345);
nand U1414 (N_1414,N_1390,N_1341);
nand U1415 (N_1415,N_1389,N_1347);
and U1416 (N_1416,N_1381,N_1340);
nor U1417 (N_1417,N_1388,N_1343);
and U1418 (N_1418,N_1348,N_1301);
nand U1419 (N_1419,N_1370,N_1335);
or U1420 (N_1420,N_1395,N_1318);
and U1421 (N_1421,N_1330,N_1303);
nand U1422 (N_1422,N_1344,N_1308);
nand U1423 (N_1423,N_1326,N_1359);
nand U1424 (N_1424,N_1398,N_1319);
nor U1425 (N_1425,N_1312,N_1310);
nor U1426 (N_1426,N_1349,N_1362);
nor U1427 (N_1427,N_1393,N_1358);
nand U1428 (N_1428,N_1383,N_1376);
nand U1429 (N_1429,N_1371,N_1361);
nor U1430 (N_1430,N_1311,N_1327);
or U1431 (N_1431,N_1320,N_1384);
and U1432 (N_1432,N_1331,N_1374);
nand U1433 (N_1433,N_1364,N_1379);
nand U1434 (N_1434,N_1355,N_1356);
or U1435 (N_1435,N_1353,N_1391);
and U1436 (N_1436,N_1314,N_1372);
or U1437 (N_1437,N_1325,N_1317);
nor U1438 (N_1438,N_1329,N_1369);
or U1439 (N_1439,N_1394,N_1375);
or U1440 (N_1440,N_1373,N_1350);
nand U1441 (N_1441,N_1386,N_1309);
nand U1442 (N_1442,N_1365,N_1346);
and U1443 (N_1443,N_1367,N_1385);
and U1444 (N_1444,N_1304,N_1351);
and U1445 (N_1445,N_1315,N_1307);
and U1446 (N_1446,N_1313,N_1305);
nor U1447 (N_1447,N_1382,N_1368);
or U1448 (N_1448,N_1300,N_1357);
or U1449 (N_1449,N_1321,N_1352);
nor U1450 (N_1450,N_1333,N_1306);
nor U1451 (N_1451,N_1315,N_1313);
nor U1452 (N_1452,N_1384,N_1337);
nor U1453 (N_1453,N_1337,N_1381);
and U1454 (N_1454,N_1348,N_1383);
and U1455 (N_1455,N_1311,N_1384);
or U1456 (N_1456,N_1309,N_1318);
and U1457 (N_1457,N_1338,N_1355);
nand U1458 (N_1458,N_1305,N_1360);
and U1459 (N_1459,N_1394,N_1362);
nor U1460 (N_1460,N_1340,N_1302);
nor U1461 (N_1461,N_1373,N_1307);
or U1462 (N_1462,N_1313,N_1357);
and U1463 (N_1463,N_1320,N_1388);
and U1464 (N_1464,N_1384,N_1326);
nand U1465 (N_1465,N_1312,N_1383);
and U1466 (N_1466,N_1377,N_1301);
nor U1467 (N_1467,N_1333,N_1337);
or U1468 (N_1468,N_1316,N_1314);
nor U1469 (N_1469,N_1306,N_1349);
and U1470 (N_1470,N_1345,N_1327);
and U1471 (N_1471,N_1357,N_1302);
nand U1472 (N_1472,N_1325,N_1353);
nor U1473 (N_1473,N_1371,N_1327);
or U1474 (N_1474,N_1320,N_1351);
and U1475 (N_1475,N_1316,N_1342);
or U1476 (N_1476,N_1345,N_1357);
and U1477 (N_1477,N_1305,N_1341);
or U1478 (N_1478,N_1398,N_1392);
xnor U1479 (N_1479,N_1320,N_1325);
nor U1480 (N_1480,N_1312,N_1362);
and U1481 (N_1481,N_1301,N_1375);
or U1482 (N_1482,N_1386,N_1357);
and U1483 (N_1483,N_1319,N_1393);
nand U1484 (N_1484,N_1381,N_1322);
nand U1485 (N_1485,N_1309,N_1374);
nand U1486 (N_1486,N_1373,N_1376);
or U1487 (N_1487,N_1326,N_1367);
and U1488 (N_1488,N_1398,N_1309);
nor U1489 (N_1489,N_1337,N_1386);
nor U1490 (N_1490,N_1385,N_1362);
nand U1491 (N_1491,N_1327,N_1344);
nand U1492 (N_1492,N_1382,N_1309);
nand U1493 (N_1493,N_1371,N_1302);
or U1494 (N_1494,N_1335,N_1396);
nor U1495 (N_1495,N_1380,N_1330);
nand U1496 (N_1496,N_1359,N_1322);
or U1497 (N_1497,N_1384,N_1313);
and U1498 (N_1498,N_1388,N_1358);
nor U1499 (N_1499,N_1334,N_1335);
and U1500 (N_1500,N_1411,N_1489);
nand U1501 (N_1501,N_1490,N_1497);
nor U1502 (N_1502,N_1427,N_1466);
and U1503 (N_1503,N_1420,N_1435);
nand U1504 (N_1504,N_1440,N_1418);
or U1505 (N_1505,N_1465,N_1486);
and U1506 (N_1506,N_1457,N_1492);
and U1507 (N_1507,N_1436,N_1450);
or U1508 (N_1508,N_1467,N_1441);
nor U1509 (N_1509,N_1488,N_1406);
or U1510 (N_1510,N_1433,N_1432);
nand U1511 (N_1511,N_1402,N_1408);
nand U1512 (N_1512,N_1417,N_1474);
nor U1513 (N_1513,N_1448,N_1476);
or U1514 (N_1514,N_1419,N_1473);
nor U1515 (N_1515,N_1462,N_1400);
nand U1516 (N_1516,N_1449,N_1471);
nand U1517 (N_1517,N_1439,N_1481);
and U1518 (N_1518,N_1480,N_1446);
nor U1519 (N_1519,N_1478,N_1430);
and U1520 (N_1520,N_1452,N_1464);
nand U1521 (N_1521,N_1484,N_1479);
nor U1522 (N_1522,N_1469,N_1414);
or U1523 (N_1523,N_1491,N_1434);
and U1524 (N_1524,N_1447,N_1495);
and U1525 (N_1525,N_1475,N_1451);
nor U1526 (N_1526,N_1422,N_1494);
or U1527 (N_1527,N_1412,N_1443);
nand U1528 (N_1528,N_1482,N_1463);
and U1529 (N_1529,N_1403,N_1470);
or U1530 (N_1530,N_1458,N_1477);
and U1531 (N_1531,N_1472,N_1442);
or U1532 (N_1532,N_1459,N_1454);
nand U1533 (N_1533,N_1428,N_1483);
nor U1534 (N_1534,N_1426,N_1429);
and U1535 (N_1535,N_1425,N_1423);
and U1536 (N_1536,N_1404,N_1499);
and U1537 (N_1537,N_1437,N_1496);
nor U1538 (N_1538,N_1453,N_1401);
and U1539 (N_1539,N_1421,N_1407);
or U1540 (N_1540,N_1456,N_1493);
and U1541 (N_1541,N_1487,N_1460);
or U1542 (N_1542,N_1444,N_1498);
nor U1543 (N_1543,N_1409,N_1410);
nand U1544 (N_1544,N_1405,N_1415);
nand U1545 (N_1545,N_1416,N_1438);
or U1546 (N_1546,N_1455,N_1461);
or U1547 (N_1547,N_1413,N_1485);
nor U1548 (N_1548,N_1445,N_1468);
nand U1549 (N_1549,N_1424,N_1431);
nand U1550 (N_1550,N_1418,N_1404);
or U1551 (N_1551,N_1404,N_1457);
or U1552 (N_1552,N_1443,N_1400);
and U1553 (N_1553,N_1417,N_1430);
and U1554 (N_1554,N_1459,N_1453);
nor U1555 (N_1555,N_1495,N_1430);
nor U1556 (N_1556,N_1429,N_1445);
and U1557 (N_1557,N_1437,N_1403);
nor U1558 (N_1558,N_1417,N_1410);
nand U1559 (N_1559,N_1452,N_1442);
nor U1560 (N_1560,N_1448,N_1412);
or U1561 (N_1561,N_1448,N_1433);
nand U1562 (N_1562,N_1429,N_1469);
nand U1563 (N_1563,N_1407,N_1490);
or U1564 (N_1564,N_1494,N_1460);
nand U1565 (N_1565,N_1435,N_1452);
nand U1566 (N_1566,N_1449,N_1442);
or U1567 (N_1567,N_1407,N_1461);
nand U1568 (N_1568,N_1420,N_1406);
and U1569 (N_1569,N_1471,N_1440);
and U1570 (N_1570,N_1406,N_1469);
nand U1571 (N_1571,N_1446,N_1456);
and U1572 (N_1572,N_1449,N_1447);
nand U1573 (N_1573,N_1411,N_1404);
nand U1574 (N_1574,N_1481,N_1427);
nand U1575 (N_1575,N_1446,N_1408);
nand U1576 (N_1576,N_1480,N_1455);
nand U1577 (N_1577,N_1474,N_1492);
and U1578 (N_1578,N_1424,N_1441);
nand U1579 (N_1579,N_1411,N_1435);
and U1580 (N_1580,N_1401,N_1461);
nand U1581 (N_1581,N_1438,N_1474);
or U1582 (N_1582,N_1497,N_1487);
and U1583 (N_1583,N_1400,N_1422);
nand U1584 (N_1584,N_1453,N_1472);
or U1585 (N_1585,N_1490,N_1401);
nand U1586 (N_1586,N_1401,N_1412);
or U1587 (N_1587,N_1424,N_1480);
and U1588 (N_1588,N_1470,N_1446);
or U1589 (N_1589,N_1438,N_1497);
and U1590 (N_1590,N_1444,N_1488);
and U1591 (N_1591,N_1493,N_1420);
nor U1592 (N_1592,N_1496,N_1493);
and U1593 (N_1593,N_1418,N_1436);
nor U1594 (N_1594,N_1450,N_1429);
nand U1595 (N_1595,N_1489,N_1436);
nor U1596 (N_1596,N_1493,N_1485);
or U1597 (N_1597,N_1447,N_1409);
nand U1598 (N_1598,N_1412,N_1457);
or U1599 (N_1599,N_1400,N_1441);
and U1600 (N_1600,N_1532,N_1553);
nor U1601 (N_1601,N_1570,N_1583);
nor U1602 (N_1602,N_1541,N_1515);
nand U1603 (N_1603,N_1552,N_1540);
or U1604 (N_1604,N_1509,N_1522);
nand U1605 (N_1605,N_1578,N_1502);
nand U1606 (N_1606,N_1569,N_1511);
or U1607 (N_1607,N_1580,N_1566);
nand U1608 (N_1608,N_1533,N_1545);
nand U1609 (N_1609,N_1567,N_1538);
nor U1610 (N_1610,N_1546,N_1564);
nor U1611 (N_1611,N_1585,N_1588);
nor U1612 (N_1612,N_1514,N_1593);
nand U1613 (N_1613,N_1568,N_1586);
or U1614 (N_1614,N_1561,N_1537);
nor U1615 (N_1615,N_1544,N_1587);
or U1616 (N_1616,N_1560,N_1597);
or U1617 (N_1617,N_1565,N_1506);
nand U1618 (N_1618,N_1581,N_1510);
nor U1619 (N_1619,N_1526,N_1542);
or U1620 (N_1620,N_1576,N_1535);
nand U1621 (N_1621,N_1536,N_1575);
and U1622 (N_1622,N_1558,N_1577);
or U1623 (N_1623,N_1563,N_1503);
or U1624 (N_1624,N_1571,N_1512);
nor U1625 (N_1625,N_1531,N_1507);
nand U1626 (N_1626,N_1534,N_1517);
nor U1627 (N_1627,N_1598,N_1520);
nand U1628 (N_1628,N_1525,N_1589);
nor U1629 (N_1629,N_1556,N_1572);
or U1630 (N_1630,N_1562,N_1501);
or U1631 (N_1631,N_1547,N_1596);
nor U1632 (N_1632,N_1513,N_1591);
or U1633 (N_1633,N_1551,N_1543);
nor U1634 (N_1634,N_1518,N_1554);
and U1635 (N_1635,N_1529,N_1500);
nor U1636 (N_1636,N_1559,N_1584);
nor U1637 (N_1637,N_1524,N_1550);
and U1638 (N_1638,N_1516,N_1530);
and U1639 (N_1639,N_1504,N_1590);
nor U1640 (N_1640,N_1548,N_1549);
or U1641 (N_1641,N_1555,N_1582);
or U1642 (N_1642,N_1528,N_1592);
or U1643 (N_1643,N_1599,N_1557);
and U1644 (N_1644,N_1579,N_1505);
or U1645 (N_1645,N_1574,N_1595);
or U1646 (N_1646,N_1519,N_1508);
and U1647 (N_1647,N_1573,N_1521);
or U1648 (N_1648,N_1539,N_1527);
and U1649 (N_1649,N_1594,N_1523);
nand U1650 (N_1650,N_1531,N_1591);
nand U1651 (N_1651,N_1518,N_1589);
nand U1652 (N_1652,N_1555,N_1556);
nand U1653 (N_1653,N_1555,N_1557);
nand U1654 (N_1654,N_1500,N_1504);
or U1655 (N_1655,N_1568,N_1511);
and U1656 (N_1656,N_1565,N_1551);
or U1657 (N_1657,N_1565,N_1513);
or U1658 (N_1658,N_1574,N_1586);
or U1659 (N_1659,N_1528,N_1590);
or U1660 (N_1660,N_1582,N_1587);
nor U1661 (N_1661,N_1547,N_1503);
and U1662 (N_1662,N_1558,N_1544);
nor U1663 (N_1663,N_1581,N_1528);
and U1664 (N_1664,N_1530,N_1571);
nor U1665 (N_1665,N_1502,N_1536);
nor U1666 (N_1666,N_1571,N_1531);
nand U1667 (N_1667,N_1525,N_1594);
or U1668 (N_1668,N_1559,N_1593);
nor U1669 (N_1669,N_1530,N_1531);
or U1670 (N_1670,N_1523,N_1546);
and U1671 (N_1671,N_1507,N_1505);
nor U1672 (N_1672,N_1537,N_1573);
nand U1673 (N_1673,N_1557,N_1545);
or U1674 (N_1674,N_1548,N_1536);
or U1675 (N_1675,N_1595,N_1560);
or U1676 (N_1676,N_1501,N_1582);
nor U1677 (N_1677,N_1572,N_1555);
and U1678 (N_1678,N_1541,N_1513);
or U1679 (N_1679,N_1559,N_1524);
nand U1680 (N_1680,N_1543,N_1573);
or U1681 (N_1681,N_1548,N_1505);
and U1682 (N_1682,N_1580,N_1531);
nand U1683 (N_1683,N_1526,N_1560);
nand U1684 (N_1684,N_1554,N_1543);
or U1685 (N_1685,N_1553,N_1537);
nand U1686 (N_1686,N_1574,N_1508);
or U1687 (N_1687,N_1598,N_1522);
and U1688 (N_1688,N_1576,N_1593);
nor U1689 (N_1689,N_1504,N_1545);
nor U1690 (N_1690,N_1560,N_1559);
nand U1691 (N_1691,N_1581,N_1523);
xnor U1692 (N_1692,N_1530,N_1539);
nor U1693 (N_1693,N_1524,N_1554);
nand U1694 (N_1694,N_1515,N_1503);
and U1695 (N_1695,N_1572,N_1592);
or U1696 (N_1696,N_1558,N_1563);
and U1697 (N_1697,N_1549,N_1582);
nand U1698 (N_1698,N_1516,N_1559);
nor U1699 (N_1699,N_1591,N_1528);
and U1700 (N_1700,N_1613,N_1618);
or U1701 (N_1701,N_1630,N_1633);
or U1702 (N_1702,N_1687,N_1678);
or U1703 (N_1703,N_1656,N_1646);
or U1704 (N_1704,N_1679,N_1648);
nor U1705 (N_1705,N_1676,N_1610);
or U1706 (N_1706,N_1649,N_1688);
nor U1707 (N_1707,N_1650,N_1644);
or U1708 (N_1708,N_1619,N_1675);
nor U1709 (N_1709,N_1665,N_1664);
or U1710 (N_1710,N_1695,N_1653);
xnor U1711 (N_1711,N_1658,N_1606);
nor U1712 (N_1712,N_1622,N_1674);
or U1713 (N_1713,N_1671,N_1668);
and U1714 (N_1714,N_1680,N_1698);
or U1715 (N_1715,N_1696,N_1624);
and U1716 (N_1716,N_1666,N_1635);
and U1717 (N_1717,N_1673,N_1614);
or U1718 (N_1718,N_1651,N_1685);
and U1719 (N_1719,N_1616,N_1691);
or U1720 (N_1720,N_1682,N_1621);
and U1721 (N_1721,N_1639,N_1600);
nor U1722 (N_1722,N_1629,N_1602);
nor U1723 (N_1723,N_1684,N_1659);
and U1724 (N_1724,N_1607,N_1632);
nor U1725 (N_1725,N_1603,N_1660);
nand U1726 (N_1726,N_1657,N_1672);
nor U1727 (N_1727,N_1623,N_1620);
nor U1728 (N_1728,N_1617,N_1628);
or U1729 (N_1729,N_1638,N_1608);
nand U1730 (N_1730,N_1647,N_1631);
and U1731 (N_1731,N_1625,N_1694);
nand U1732 (N_1732,N_1670,N_1693);
and U1733 (N_1733,N_1636,N_1626);
nor U1734 (N_1734,N_1692,N_1652);
or U1735 (N_1735,N_1662,N_1642);
or U1736 (N_1736,N_1686,N_1655);
nand U1737 (N_1737,N_1637,N_1681);
and U1738 (N_1738,N_1634,N_1661);
and U1739 (N_1739,N_1640,N_1667);
nand U1740 (N_1740,N_1627,N_1663);
or U1741 (N_1741,N_1683,N_1697);
and U1742 (N_1742,N_1615,N_1612);
nor U1743 (N_1743,N_1690,N_1669);
nand U1744 (N_1744,N_1605,N_1699);
or U1745 (N_1745,N_1677,N_1654);
nand U1746 (N_1746,N_1689,N_1611);
nor U1747 (N_1747,N_1645,N_1641);
or U1748 (N_1748,N_1604,N_1643);
or U1749 (N_1749,N_1601,N_1609);
nor U1750 (N_1750,N_1616,N_1679);
and U1751 (N_1751,N_1671,N_1612);
nor U1752 (N_1752,N_1661,N_1615);
and U1753 (N_1753,N_1675,N_1698);
and U1754 (N_1754,N_1651,N_1653);
nor U1755 (N_1755,N_1698,N_1629);
and U1756 (N_1756,N_1642,N_1670);
nor U1757 (N_1757,N_1657,N_1628);
and U1758 (N_1758,N_1668,N_1621);
nand U1759 (N_1759,N_1686,N_1608);
and U1760 (N_1760,N_1666,N_1691);
nor U1761 (N_1761,N_1690,N_1668);
nor U1762 (N_1762,N_1627,N_1637);
or U1763 (N_1763,N_1682,N_1603);
and U1764 (N_1764,N_1677,N_1689);
nand U1765 (N_1765,N_1601,N_1602);
or U1766 (N_1766,N_1650,N_1607);
or U1767 (N_1767,N_1623,N_1663);
or U1768 (N_1768,N_1698,N_1601);
nor U1769 (N_1769,N_1608,N_1646);
or U1770 (N_1770,N_1637,N_1696);
and U1771 (N_1771,N_1687,N_1699);
xnor U1772 (N_1772,N_1676,N_1623);
and U1773 (N_1773,N_1670,N_1688);
nor U1774 (N_1774,N_1628,N_1608);
or U1775 (N_1775,N_1683,N_1651);
nor U1776 (N_1776,N_1608,N_1679);
nor U1777 (N_1777,N_1614,N_1641);
and U1778 (N_1778,N_1629,N_1640);
or U1779 (N_1779,N_1658,N_1624);
nand U1780 (N_1780,N_1670,N_1695);
or U1781 (N_1781,N_1615,N_1629);
and U1782 (N_1782,N_1629,N_1623);
or U1783 (N_1783,N_1622,N_1637);
or U1784 (N_1784,N_1676,N_1661);
and U1785 (N_1785,N_1635,N_1631);
nand U1786 (N_1786,N_1613,N_1648);
xor U1787 (N_1787,N_1684,N_1681);
and U1788 (N_1788,N_1600,N_1693);
or U1789 (N_1789,N_1671,N_1632);
or U1790 (N_1790,N_1620,N_1697);
xor U1791 (N_1791,N_1697,N_1672);
nand U1792 (N_1792,N_1657,N_1697);
nor U1793 (N_1793,N_1674,N_1632);
nand U1794 (N_1794,N_1666,N_1697);
nor U1795 (N_1795,N_1636,N_1681);
nand U1796 (N_1796,N_1618,N_1699);
nor U1797 (N_1797,N_1692,N_1602);
nand U1798 (N_1798,N_1633,N_1676);
and U1799 (N_1799,N_1650,N_1656);
nand U1800 (N_1800,N_1731,N_1767);
nand U1801 (N_1801,N_1739,N_1796);
nand U1802 (N_1802,N_1755,N_1714);
and U1803 (N_1803,N_1763,N_1701);
nor U1804 (N_1804,N_1740,N_1703);
and U1805 (N_1805,N_1754,N_1746);
nor U1806 (N_1806,N_1720,N_1758);
nand U1807 (N_1807,N_1729,N_1782);
nand U1808 (N_1808,N_1752,N_1719);
nor U1809 (N_1809,N_1722,N_1750);
nor U1810 (N_1810,N_1790,N_1706);
and U1811 (N_1811,N_1745,N_1715);
and U1812 (N_1812,N_1708,N_1765);
and U1813 (N_1813,N_1770,N_1756);
and U1814 (N_1814,N_1759,N_1717);
or U1815 (N_1815,N_1794,N_1716);
nand U1816 (N_1816,N_1709,N_1768);
and U1817 (N_1817,N_1757,N_1789);
or U1818 (N_1818,N_1787,N_1762);
nand U1819 (N_1819,N_1707,N_1771);
nor U1820 (N_1820,N_1748,N_1779);
or U1821 (N_1821,N_1734,N_1736);
nor U1822 (N_1822,N_1773,N_1704);
nor U1823 (N_1823,N_1727,N_1798);
nand U1824 (N_1824,N_1788,N_1785);
and U1825 (N_1825,N_1741,N_1742);
and U1826 (N_1826,N_1723,N_1728);
and U1827 (N_1827,N_1797,N_1780);
nor U1828 (N_1828,N_1710,N_1700);
or U1829 (N_1829,N_1711,N_1751);
nand U1830 (N_1830,N_1702,N_1735);
or U1831 (N_1831,N_1761,N_1737);
or U1832 (N_1832,N_1786,N_1791);
xnor U1833 (N_1833,N_1724,N_1781);
or U1834 (N_1834,N_1784,N_1743);
or U1835 (N_1835,N_1712,N_1721);
and U1836 (N_1836,N_1793,N_1775);
or U1837 (N_1837,N_1738,N_1749);
or U1838 (N_1838,N_1766,N_1772);
or U1839 (N_1839,N_1769,N_1730);
and U1840 (N_1840,N_1733,N_1783);
nor U1841 (N_1841,N_1753,N_1764);
and U1842 (N_1842,N_1718,N_1732);
nor U1843 (N_1843,N_1777,N_1744);
nor U1844 (N_1844,N_1747,N_1795);
and U1845 (N_1845,N_1760,N_1713);
nor U1846 (N_1846,N_1799,N_1705);
or U1847 (N_1847,N_1778,N_1726);
or U1848 (N_1848,N_1792,N_1774);
or U1849 (N_1849,N_1776,N_1725);
nor U1850 (N_1850,N_1755,N_1728);
and U1851 (N_1851,N_1786,N_1735);
nor U1852 (N_1852,N_1752,N_1741);
nand U1853 (N_1853,N_1700,N_1760);
and U1854 (N_1854,N_1748,N_1727);
nand U1855 (N_1855,N_1756,N_1746);
or U1856 (N_1856,N_1779,N_1777);
nor U1857 (N_1857,N_1797,N_1720);
nor U1858 (N_1858,N_1765,N_1743);
and U1859 (N_1859,N_1757,N_1726);
nor U1860 (N_1860,N_1799,N_1746);
and U1861 (N_1861,N_1790,N_1762);
nand U1862 (N_1862,N_1767,N_1702);
nor U1863 (N_1863,N_1777,N_1728);
nor U1864 (N_1864,N_1797,N_1704);
or U1865 (N_1865,N_1750,N_1745);
and U1866 (N_1866,N_1750,N_1749);
nor U1867 (N_1867,N_1758,N_1714);
nor U1868 (N_1868,N_1754,N_1783);
nand U1869 (N_1869,N_1702,N_1795);
and U1870 (N_1870,N_1749,N_1765);
nor U1871 (N_1871,N_1716,N_1798);
or U1872 (N_1872,N_1758,N_1771);
nor U1873 (N_1873,N_1744,N_1707);
nand U1874 (N_1874,N_1734,N_1710);
nand U1875 (N_1875,N_1720,N_1765);
or U1876 (N_1876,N_1771,N_1740);
xnor U1877 (N_1877,N_1714,N_1757);
nand U1878 (N_1878,N_1714,N_1731);
nand U1879 (N_1879,N_1736,N_1786);
or U1880 (N_1880,N_1786,N_1775);
or U1881 (N_1881,N_1720,N_1763);
and U1882 (N_1882,N_1762,N_1743);
and U1883 (N_1883,N_1722,N_1758);
nand U1884 (N_1884,N_1703,N_1787);
or U1885 (N_1885,N_1799,N_1751);
nor U1886 (N_1886,N_1711,N_1785);
or U1887 (N_1887,N_1717,N_1784);
nor U1888 (N_1888,N_1767,N_1735);
and U1889 (N_1889,N_1748,N_1775);
nand U1890 (N_1890,N_1780,N_1733);
nor U1891 (N_1891,N_1793,N_1784);
nor U1892 (N_1892,N_1711,N_1753);
or U1893 (N_1893,N_1732,N_1738);
and U1894 (N_1894,N_1762,N_1782);
nand U1895 (N_1895,N_1791,N_1717);
nor U1896 (N_1896,N_1701,N_1731);
nand U1897 (N_1897,N_1751,N_1798);
and U1898 (N_1898,N_1792,N_1735);
or U1899 (N_1899,N_1762,N_1707);
or U1900 (N_1900,N_1834,N_1844);
or U1901 (N_1901,N_1891,N_1870);
and U1902 (N_1902,N_1848,N_1831);
and U1903 (N_1903,N_1895,N_1811);
and U1904 (N_1904,N_1894,N_1837);
and U1905 (N_1905,N_1869,N_1850);
or U1906 (N_1906,N_1886,N_1843);
and U1907 (N_1907,N_1860,N_1875);
and U1908 (N_1908,N_1847,N_1813);
nor U1909 (N_1909,N_1824,N_1820);
nand U1910 (N_1910,N_1849,N_1862);
nand U1911 (N_1911,N_1896,N_1867);
nor U1912 (N_1912,N_1806,N_1852);
nand U1913 (N_1913,N_1840,N_1812);
nor U1914 (N_1914,N_1857,N_1864);
nand U1915 (N_1915,N_1854,N_1833);
xor U1916 (N_1916,N_1826,N_1803);
and U1917 (N_1917,N_1810,N_1876);
and U1918 (N_1918,N_1822,N_1880);
and U1919 (N_1919,N_1805,N_1866);
nor U1920 (N_1920,N_1804,N_1830);
or U1921 (N_1921,N_1884,N_1808);
or U1922 (N_1922,N_1832,N_1873);
or U1923 (N_1923,N_1842,N_1815);
nand U1924 (N_1924,N_1889,N_1878);
nand U1925 (N_1925,N_1855,N_1817);
or U1926 (N_1926,N_1829,N_1839);
nor U1927 (N_1927,N_1818,N_1887);
nor U1928 (N_1928,N_1872,N_1823);
nand U1929 (N_1929,N_1898,N_1853);
or U1930 (N_1930,N_1828,N_1841);
and U1931 (N_1931,N_1819,N_1885);
or U1932 (N_1932,N_1821,N_1871);
nand U1933 (N_1933,N_1809,N_1807);
or U1934 (N_1934,N_1836,N_1845);
nor U1935 (N_1935,N_1800,N_1865);
and U1936 (N_1936,N_1835,N_1858);
nand U1937 (N_1937,N_1879,N_1856);
nand U1938 (N_1938,N_1874,N_1846);
or U1939 (N_1939,N_1816,N_1802);
or U1940 (N_1940,N_1897,N_1814);
nand U1941 (N_1941,N_1851,N_1827);
and U1942 (N_1942,N_1888,N_1863);
nor U1943 (N_1943,N_1868,N_1801);
or U1944 (N_1944,N_1877,N_1825);
or U1945 (N_1945,N_1859,N_1838);
and U1946 (N_1946,N_1882,N_1892);
xor U1947 (N_1947,N_1881,N_1890);
and U1948 (N_1948,N_1861,N_1883);
nor U1949 (N_1949,N_1899,N_1893);
or U1950 (N_1950,N_1873,N_1891);
and U1951 (N_1951,N_1842,N_1844);
or U1952 (N_1952,N_1809,N_1873);
and U1953 (N_1953,N_1844,N_1848);
or U1954 (N_1954,N_1877,N_1831);
or U1955 (N_1955,N_1863,N_1840);
or U1956 (N_1956,N_1841,N_1800);
or U1957 (N_1957,N_1894,N_1869);
nand U1958 (N_1958,N_1860,N_1803);
and U1959 (N_1959,N_1833,N_1808);
nand U1960 (N_1960,N_1818,N_1810);
and U1961 (N_1961,N_1891,N_1892);
and U1962 (N_1962,N_1832,N_1892);
nand U1963 (N_1963,N_1850,N_1884);
nor U1964 (N_1964,N_1853,N_1837);
nand U1965 (N_1965,N_1892,N_1807);
nand U1966 (N_1966,N_1843,N_1801);
nand U1967 (N_1967,N_1857,N_1863);
nor U1968 (N_1968,N_1853,N_1842);
and U1969 (N_1969,N_1896,N_1871);
nand U1970 (N_1970,N_1817,N_1841);
nor U1971 (N_1971,N_1814,N_1825);
or U1972 (N_1972,N_1848,N_1816);
nand U1973 (N_1973,N_1824,N_1872);
and U1974 (N_1974,N_1856,N_1829);
and U1975 (N_1975,N_1860,N_1896);
or U1976 (N_1976,N_1868,N_1894);
nand U1977 (N_1977,N_1897,N_1800);
nor U1978 (N_1978,N_1812,N_1806);
nand U1979 (N_1979,N_1893,N_1850);
nand U1980 (N_1980,N_1852,N_1863);
nand U1981 (N_1981,N_1816,N_1860);
or U1982 (N_1982,N_1831,N_1827);
or U1983 (N_1983,N_1817,N_1824);
or U1984 (N_1984,N_1820,N_1871);
nand U1985 (N_1985,N_1829,N_1873);
nor U1986 (N_1986,N_1806,N_1856);
xnor U1987 (N_1987,N_1834,N_1846);
nand U1988 (N_1988,N_1826,N_1871);
nor U1989 (N_1989,N_1822,N_1803);
or U1990 (N_1990,N_1899,N_1874);
nor U1991 (N_1991,N_1811,N_1841);
nor U1992 (N_1992,N_1881,N_1885);
nor U1993 (N_1993,N_1808,N_1863);
nand U1994 (N_1994,N_1874,N_1841);
or U1995 (N_1995,N_1845,N_1802);
or U1996 (N_1996,N_1819,N_1848);
and U1997 (N_1997,N_1871,N_1862);
and U1998 (N_1998,N_1858,N_1893);
xnor U1999 (N_1999,N_1876,N_1851);
nor U2000 (N_2000,N_1902,N_1989);
or U2001 (N_2001,N_1945,N_1934);
nor U2002 (N_2002,N_1999,N_1975);
and U2003 (N_2003,N_1969,N_1930);
or U2004 (N_2004,N_1911,N_1967);
and U2005 (N_2005,N_1997,N_1988);
and U2006 (N_2006,N_1953,N_1977);
nor U2007 (N_2007,N_1979,N_1992);
nor U2008 (N_2008,N_1970,N_1951);
nand U2009 (N_2009,N_1913,N_1972);
and U2010 (N_2010,N_1983,N_1964);
and U2011 (N_2011,N_1990,N_1939);
nor U2012 (N_2012,N_1949,N_1908);
and U2013 (N_2013,N_1933,N_1931);
nand U2014 (N_2014,N_1950,N_1944);
nor U2015 (N_2015,N_1922,N_1936);
nand U2016 (N_2016,N_1985,N_1940);
or U2017 (N_2017,N_1901,N_1900);
nor U2018 (N_2018,N_1948,N_1905);
or U2019 (N_2019,N_1929,N_1955);
or U2020 (N_2020,N_1954,N_1947);
nor U2021 (N_2021,N_1927,N_1919);
or U2022 (N_2022,N_1923,N_1959);
and U2023 (N_2023,N_1963,N_1928);
and U2024 (N_2024,N_1920,N_1978);
or U2025 (N_2025,N_1974,N_1943);
or U2026 (N_2026,N_1961,N_1909);
nand U2027 (N_2027,N_1937,N_1915);
nand U2028 (N_2028,N_1982,N_1958);
nand U2029 (N_2029,N_1914,N_1984);
and U2030 (N_2030,N_1991,N_1921);
nand U2031 (N_2031,N_1946,N_1966);
nand U2032 (N_2032,N_1952,N_1918);
and U2033 (N_2033,N_1994,N_1925);
nand U2034 (N_2034,N_1941,N_1903);
nor U2035 (N_2035,N_1912,N_1998);
and U2036 (N_2036,N_1987,N_1993);
nand U2037 (N_2037,N_1962,N_1976);
and U2038 (N_2038,N_1932,N_1942);
nor U2039 (N_2039,N_1910,N_1995);
nor U2040 (N_2040,N_1996,N_1935);
nor U2041 (N_2041,N_1981,N_1956);
and U2042 (N_2042,N_1938,N_1973);
and U2043 (N_2043,N_1906,N_1986);
xnor U2044 (N_2044,N_1965,N_1971);
nand U2045 (N_2045,N_1926,N_1917);
and U2046 (N_2046,N_1968,N_1916);
nor U2047 (N_2047,N_1960,N_1980);
nand U2048 (N_2048,N_1907,N_1957);
nor U2049 (N_2049,N_1904,N_1924);
nor U2050 (N_2050,N_1992,N_1988);
and U2051 (N_2051,N_1908,N_1903);
nor U2052 (N_2052,N_1935,N_1999);
and U2053 (N_2053,N_1979,N_1912);
nor U2054 (N_2054,N_1985,N_1942);
nand U2055 (N_2055,N_1905,N_1926);
nor U2056 (N_2056,N_1984,N_1987);
xnor U2057 (N_2057,N_1968,N_1910);
nor U2058 (N_2058,N_1960,N_1997);
and U2059 (N_2059,N_1986,N_1921);
xnor U2060 (N_2060,N_1978,N_1930);
nor U2061 (N_2061,N_1946,N_1922);
and U2062 (N_2062,N_1999,N_1927);
nor U2063 (N_2063,N_1988,N_1961);
or U2064 (N_2064,N_1964,N_1969);
nand U2065 (N_2065,N_1935,N_1963);
nor U2066 (N_2066,N_1901,N_1990);
and U2067 (N_2067,N_1929,N_1917);
nand U2068 (N_2068,N_1949,N_1987);
or U2069 (N_2069,N_1956,N_1909);
and U2070 (N_2070,N_1956,N_1920);
nor U2071 (N_2071,N_1987,N_1996);
nor U2072 (N_2072,N_1954,N_1906);
or U2073 (N_2073,N_1954,N_1957);
nor U2074 (N_2074,N_1991,N_1982);
or U2075 (N_2075,N_1921,N_1965);
and U2076 (N_2076,N_1967,N_1996);
and U2077 (N_2077,N_1963,N_1971);
and U2078 (N_2078,N_1943,N_1941);
nor U2079 (N_2079,N_1934,N_1987);
nor U2080 (N_2080,N_1948,N_1975);
or U2081 (N_2081,N_1903,N_1929);
nand U2082 (N_2082,N_1993,N_1949);
and U2083 (N_2083,N_1938,N_1993);
or U2084 (N_2084,N_1962,N_1963);
and U2085 (N_2085,N_1980,N_1923);
or U2086 (N_2086,N_1971,N_1939);
nand U2087 (N_2087,N_1932,N_1902);
nand U2088 (N_2088,N_1955,N_1919);
nand U2089 (N_2089,N_1971,N_1912);
nor U2090 (N_2090,N_1943,N_1907);
nor U2091 (N_2091,N_1953,N_1959);
and U2092 (N_2092,N_1983,N_1948);
or U2093 (N_2093,N_1976,N_1955);
and U2094 (N_2094,N_1999,N_1943);
nand U2095 (N_2095,N_1997,N_1927);
and U2096 (N_2096,N_1991,N_1933);
nand U2097 (N_2097,N_1912,N_1945);
nand U2098 (N_2098,N_1953,N_1968);
nor U2099 (N_2099,N_1998,N_1995);
nand U2100 (N_2100,N_2007,N_2094);
or U2101 (N_2101,N_2018,N_2001);
nand U2102 (N_2102,N_2055,N_2060);
or U2103 (N_2103,N_2036,N_2038);
or U2104 (N_2104,N_2006,N_2081);
nor U2105 (N_2105,N_2088,N_2048);
or U2106 (N_2106,N_2076,N_2033);
nor U2107 (N_2107,N_2089,N_2090);
or U2108 (N_2108,N_2067,N_2014);
and U2109 (N_2109,N_2054,N_2026);
or U2110 (N_2110,N_2044,N_2077);
or U2111 (N_2111,N_2010,N_2052);
and U2112 (N_2112,N_2095,N_2057);
nand U2113 (N_2113,N_2079,N_2040);
nor U2114 (N_2114,N_2030,N_2029);
nand U2115 (N_2115,N_2062,N_2075);
or U2116 (N_2116,N_2074,N_2072);
nand U2117 (N_2117,N_2032,N_2058);
nor U2118 (N_2118,N_2042,N_2080);
nor U2119 (N_2119,N_2092,N_2009);
or U2120 (N_2120,N_2027,N_2056);
and U2121 (N_2121,N_2025,N_2015);
nand U2122 (N_2122,N_2093,N_2037);
nor U2123 (N_2123,N_2023,N_2022);
xor U2124 (N_2124,N_2046,N_2099);
and U2125 (N_2125,N_2004,N_2061);
or U2126 (N_2126,N_2039,N_2053);
or U2127 (N_2127,N_2071,N_2005);
and U2128 (N_2128,N_2034,N_2083);
and U2129 (N_2129,N_2063,N_2068);
nand U2130 (N_2130,N_2003,N_2051);
nor U2131 (N_2131,N_2017,N_2091);
or U2132 (N_2132,N_2066,N_2012);
nor U2133 (N_2133,N_2078,N_2096);
and U2134 (N_2134,N_2041,N_2087);
or U2135 (N_2135,N_2021,N_2024);
or U2136 (N_2136,N_2065,N_2043);
or U2137 (N_2137,N_2082,N_2000);
nor U2138 (N_2138,N_2085,N_2019);
nor U2139 (N_2139,N_2084,N_2098);
and U2140 (N_2140,N_2045,N_2028);
nor U2141 (N_2141,N_2013,N_2069);
or U2142 (N_2142,N_2008,N_2047);
and U2143 (N_2143,N_2002,N_2073);
nand U2144 (N_2144,N_2070,N_2011);
and U2145 (N_2145,N_2064,N_2050);
and U2146 (N_2146,N_2049,N_2086);
nor U2147 (N_2147,N_2031,N_2020);
or U2148 (N_2148,N_2097,N_2059);
and U2149 (N_2149,N_2035,N_2016);
nand U2150 (N_2150,N_2089,N_2012);
nor U2151 (N_2151,N_2059,N_2083);
nor U2152 (N_2152,N_2070,N_2063);
and U2153 (N_2153,N_2040,N_2010);
nand U2154 (N_2154,N_2020,N_2004);
or U2155 (N_2155,N_2051,N_2000);
or U2156 (N_2156,N_2089,N_2061);
nor U2157 (N_2157,N_2026,N_2095);
and U2158 (N_2158,N_2025,N_2024);
and U2159 (N_2159,N_2054,N_2046);
and U2160 (N_2160,N_2072,N_2029);
nor U2161 (N_2161,N_2035,N_2002);
or U2162 (N_2162,N_2032,N_2023);
or U2163 (N_2163,N_2036,N_2010);
nand U2164 (N_2164,N_2085,N_2047);
nor U2165 (N_2165,N_2010,N_2079);
nand U2166 (N_2166,N_2015,N_2000);
nand U2167 (N_2167,N_2096,N_2060);
nand U2168 (N_2168,N_2016,N_2008);
or U2169 (N_2169,N_2011,N_2042);
nor U2170 (N_2170,N_2020,N_2067);
or U2171 (N_2171,N_2075,N_2046);
nor U2172 (N_2172,N_2065,N_2096);
nor U2173 (N_2173,N_2054,N_2016);
nor U2174 (N_2174,N_2040,N_2087);
or U2175 (N_2175,N_2051,N_2072);
and U2176 (N_2176,N_2076,N_2060);
or U2177 (N_2177,N_2021,N_2055);
nor U2178 (N_2178,N_2049,N_2095);
or U2179 (N_2179,N_2088,N_2028);
and U2180 (N_2180,N_2065,N_2037);
nor U2181 (N_2181,N_2086,N_2069);
nand U2182 (N_2182,N_2051,N_2089);
nor U2183 (N_2183,N_2013,N_2088);
or U2184 (N_2184,N_2017,N_2058);
and U2185 (N_2185,N_2085,N_2028);
or U2186 (N_2186,N_2029,N_2016);
xor U2187 (N_2187,N_2049,N_2073);
or U2188 (N_2188,N_2058,N_2077);
or U2189 (N_2189,N_2057,N_2038);
and U2190 (N_2190,N_2045,N_2064);
or U2191 (N_2191,N_2084,N_2016);
nor U2192 (N_2192,N_2078,N_2073);
or U2193 (N_2193,N_2082,N_2089);
or U2194 (N_2194,N_2063,N_2079);
or U2195 (N_2195,N_2043,N_2000);
nor U2196 (N_2196,N_2023,N_2070);
nand U2197 (N_2197,N_2080,N_2098);
and U2198 (N_2198,N_2095,N_2075);
or U2199 (N_2199,N_2034,N_2058);
xnor U2200 (N_2200,N_2141,N_2196);
nor U2201 (N_2201,N_2164,N_2126);
xor U2202 (N_2202,N_2186,N_2149);
nand U2203 (N_2203,N_2159,N_2115);
nor U2204 (N_2204,N_2139,N_2185);
nor U2205 (N_2205,N_2107,N_2119);
nor U2206 (N_2206,N_2184,N_2122);
nor U2207 (N_2207,N_2124,N_2168);
nor U2208 (N_2208,N_2127,N_2133);
nand U2209 (N_2209,N_2187,N_2111);
and U2210 (N_2210,N_2114,N_2132);
nand U2211 (N_2211,N_2156,N_2145);
nand U2212 (N_2212,N_2104,N_2173);
nor U2213 (N_2213,N_2193,N_2194);
or U2214 (N_2214,N_2189,N_2113);
or U2215 (N_2215,N_2174,N_2135);
nor U2216 (N_2216,N_2183,N_2140);
and U2217 (N_2217,N_2157,N_2188);
nand U2218 (N_2218,N_2103,N_2197);
nand U2219 (N_2219,N_2131,N_2198);
nor U2220 (N_2220,N_2105,N_2130);
nand U2221 (N_2221,N_2182,N_2155);
or U2222 (N_2222,N_2147,N_2125);
and U2223 (N_2223,N_2169,N_2158);
xnor U2224 (N_2224,N_2151,N_2146);
and U2225 (N_2225,N_2150,N_2123);
and U2226 (N_2226,N_2152,N_2101);
or U2227 (N_2227,N_2129,N_2160);
nand U2228 (N_2228,N_2161,N_2176);
and U2229 (N_2229,N_2167,N_2162);
or U2230 (N_2230,N_2120,N_2180);
and U2231 (N_2231,N_2108,N_2166);
nor U2232 (N_2232,N_2179,N_2175);
nand U2233 (N_2233,N_2144,N_2154);
nand U2234 (N_2234,N_2142,N_2106);
or U2235 (N_2235,N_2143,N_2170);
nor U2236 (N_2236,N_2171,N_2117);
or U2237 (N_2237,N_2110,N_2128);
nand U2238 (N_2238,N_2172,N_2153);
or U2239 (N_2239,N_2102,N_2118);
nor U2240 (N_2240,N_2116,N_2199);
nor U2241 (N_2241,N_2100,N_2190);
or U2242 (N_2242,N_2121,N_2181);
nand U2243 (N_2243,N_2134,N_2177);
nor U2244 (N_2244,N_2136,N_2109);
nand U2245 (N_2245,N_2112,N_2138);
nor U2246 (N_2246,N_2191,N_2163);
and U2247 (N_2247,N_2148,N_2195);
nor U2248 (N_2248,N_2178,N_2165);
and U2249 (N_2249,N_2192,N_2137);
or U2250 (N_2250,N_2140,N_2194);
or U2251 (N_2251,N_2190,N_2109);
or U2252 (N_2252,N_2198,N_2159);
nand U2253 (N_2253,N_2173,N_2170);
nor U2254 (N_2254,N_2168,N_2145);
and U2255 (N_2255,N_2126,N_2170);
and U2256 (N_2256,N_2184,N_2134);
nor U2257 (N_2257,N_2185,N_2188);
nor U2258 (N_2258,N_2120,N_2187);
or U2259 (N_2259,N_2159,N_2146);
or U2260 (N_2260,N_2190,N_2189);
nor U2261 (N_2261,N_2152,N_2112);
and U2262 (N_2262,N_2142,N_2170);
and U2263 (N_2263,N_2196,N_2106);
nor U2264 (N_2264,N_2123,N_2138);
and U2265 (N_2265,N_2169,N_2118);
and U2266 (N_2266,N_2172,N_2138);
and U2267 (N_2267,N_2182,N_2139);
nand U2268 (N_2268,N_2147,N_2183);
or U2269 (N_2269,N_2161,N_2162);
and U2270 (N_2270,N_2152,N_2120);
and U2271 (N_2271,N_2152,N_2129);
nand U2272 (N_2272,N_2106,N_2189);
nor U2273 (N_2273,N_2138,N_2187);
nor U2274 (N_2274,N_2157,N_2193);
nor U2275 (N_2275,N_2104,N_2153);
or U2276 (N_2276,N_2117,N_2158);
and U2277 (N_2277,N_2174,N_2193);
nor U2278 (N_2278,N_2152,N_2157);
or U2279 (N_2279,N_2118,N_2189);
nor U2280 (N_2280,N_2145,N_2179);
or U2281 (N_2281,N_2125,N_2148);
nand U2282 (N_2282,N_2138,N_2142);
nand U2283 (N_2283,N_2154,N_2167);
and U2284 (N_2284,N_2197,N_2146);
nor U2285 (N_2285,N_2182,N_2197);
and U2286 (N_2286,N_2107,N_2120);
nand U2287 (N_2287,N_2105,N_2181);
xnor U2288 (N_2288,N_2148,N_2198);
nand U2289 (N_2289,N_2116,N_2127);
nor U2290 (N_2290,N_2167,N_2178);
nor U2291 (N_2291,N_2166,N_2117);
or U2292 (N_2292,N_2192,N_2100);
nand U2293 (N_2293,N_2153,N_2170);
or U2294 (N_2294,N_2135,N_2192);
nand U2295 (N_2295,N_2169,N_2167);
xor U2296 (N_2296,N_2129,N_2108);
and U2297 (N_2297,N_2179,N_2142);
and U2298 (N_2298,N_2177,N_2109);
or U2299 (N_2299,N_2147,N_2164);
nor U2300 (N_2300,N_2206,N_2250);
nand U2301 (N_2301,N_2271,N_2286);
nor U2302 (N_2302,N_2265,N_2214);
nand U2303 (N_2303,N_2216,N_2285);
or U2304 (N_2304,N_2240,N_2259);
nand U2305 (N_2305,N_2200,N_2257);
nand U2306 (N_2306,N_2212,N_2238);
and U2307 (N_2307,N_2226,N_2217);
nand U2308 (N_2308,N_2258,N_2210);
nor U2309 (N_2309,N_2247,N_2263);
nor U2310 (N_2310,N_2254,N_2225);
or U2311 (N_2311,N_2239,N_2253);
nor U2312 (N_2312,N_2203,N_2245);
or U2313 (N_2313,N_2227,N_2215);
nand U2314 (N_2314,N_2281,N_2276);
nand U2315 (N_2315,N_2264,N_2223);
nand U2316 (N_2316,N_2292,N_2236);
and U2317 (N_2317,N_2298,N_2278);
and U2318 (N_2318,N_2249,N_2237);
nor U2319 (N_2319,N_2207,N_2231);
and U2320 (N_2320,N_2244,N_2204);
or U2321 (N_2321,N_2218,N_2202);
or U2322 (N_2322,N_2279,N_2262);
nand U2323 (N_2323,N_2209,N_2268);
nor U2324 (N_2324,N_2277,N_2228);
nand U2325 (N_2325,N_2283,N_2294);
and U2326 (N_2326,N_2243,N_2252);
nand U2327 (N_2327,N_2229,N_2295);
or U2328 (N_2328,N_2235,N_2201);
nand U2329 (N_2329,N_2291,N_2224);
and U2330 (N_2330,N_2270,N_2287);
or U2331 (N_2331,N_2297,N_2251);
nor U2332 (N_2332,N_2280,N_2272);
and U2333 (N_2333,N_2282,N_2221);
nor U2334 (N_2334,N_2261,N_2222);
or U2335 (N_2335,N_2208,N_2293);
or U2336 (N_2336,N_2256,N_2275);
and U2337 (N_2337,N_2267,N_2232);
nand U2338 (N_2338,N_2213,N_2284);
or U2339 (N_2339,N_2219,N_2260);
or U2340 (N_2340,N_2274,N_2205);
or U2341 (N_2341,N_2220,N_2288);
and U2342 (N_2342,N_2234,N_2233);
or U2343 (N_2343,N_2241,N_2246);
and U2344 (N_2344,N_2230,N_2289);
or U2345 (N_2345,N_2299,N_2290);
or U2346 (N_2346,N_2248,N_2255);
or U2347 (N_2347,N_2242,N_2266);
nand U2348 (N_2348,N_2296,N_2211);
nand U2349 (N_2349,N_2273,N_2269);
nand U2350 (N_2350,N_2228,N_2288);
nor U2351 (N_2351,N_2256,N_2296);
or U2352 (N_2352,N_2258,N_2248);
and U2353 (N_2353,N_2201,N_2257);
nor U2354 (N_2354,N_2276,N_2230);
nor U2355 (N_2355,N_2237,N_2270);
nand U2356 (N_2356,N_2201,N_2266);
or U2357 (N_2357,N_2243,N_2249);
nand U2358 (N_2358,N_2204,N_2242);
nand U2359 (N_2359,N_2284,N_2299);
nand U2360 (N_2360,N_2268,N_2281);
and U2361 (N_2361,N_2257,N_2240);
nor U2362 (N_2362,N_2201,N_2287);
nand U2363 (N_2363,N_2235,N_2246);
nand U2364 (N_2364,N_2207,N_2218);
nor U2365 (N_2365,N_2269,N_2224);
nand U2366 (N_2366,N_2244,N_2260);
nor U2367 (N_2367,N_2265,N_2295);
or U2368 (N_2368,N_2201,N_2225);
nor U2369 (N_2369,N_2262,N_2245);
nor U2370 (N_2370,N_2217,N_2235);
and U2371 (N_2371,N_2229,N_2231);
nor U2372 (N_2372,N_2238,N_2214);
nand U2373 (N_2373,N_2247,N_2290);
and U2374 (N_2374,N_2224,N_2248);
nor U2375 (N_2375,N_2286,N_2299);
and U2376 (N_2376,N_2214,N_2284);
nand U2377 (N_2377,N_2283,N_2208);
and U2378 (N_2378,N_2292,N_2260);
nand U2379 (N_2379,N_2260,N_2261);
nand U2380 (N_2380,N_2271,N_2296);
nand U2381 (N_2381,N_2288,N_2212);
nand U2382 (N_2382,N_2233,N_2210);
and U2383 (N_2383,N_2200,N_2291);
or U2384 (N_2384,N_2255,N_2250);
nor U2385 (N_2385,N_2205,N_2242);
or U2386 (N_2386,N_2229,N_2250);
xor U2387 (N_2387,N_2203,N_2202);
nor U2388 (N_2388,N_2208,N_2216);
and U2389 (N_2389,N_2287,N_2223);
and U2390 (N_2390,N_2277,N_2254);
nand U2391 (N_2391,N_2275,N_2219);
nand U2392 (N_2392,N_2287,N_2265);
xor U2393 (N_2393,N_2265,N_2294);
or U2394 (N_2394,N_2254,N_2299);
nor U2395 (N_2395,N_2219,N_2222);
and U2396 (N_2396,N_2206,N_2282);
nand U2397 (N_2397,N_2282,N_2204);
and U2398 (N_2398,N_2295,N_2240);
nand U2399 (N_2399,N_2293,N_2295);
nand U2400 (N_2400,N_2376,N_2365);
or U2401 (N_2401,N_2366,N_2382);
nor U2402 (N_2402,N_2358,N_2332);
nand U2403 (N_2403,N_2381,N_2343);
and U2404 (N_2404,N_2386,N_2334);
or U2405 (N_2405,N_2349,N_2325);
nand U2406 (N_2406,N_2338,N_2310);
nand U2407 (N_2407,N_2359,N_2330);
and U2408 (N_2408,N_2391,N_2397);
nand U2409 (N_2409,N_2339,N_2374);
or U2410 (N_2410,N_2395,N_2308);
or U2411 (N_2411,N_2341,N_2301);
nor U2412 (N_2412,N_2340,N_2315);
and U2413 (N_2413,N_2370,N_2348);
or U2414 (N_2414,N_2327,N_2385);
or U2415 (N_2415,N_2361,N_2360);
and U2416 (N_2416,N_2398,N_2368);
nand U2417 (N_2417,N_2387,N_2304);
and U2418 (N_2418,N_2303,N_2363);
and U2419 (N_2419,N_2357,N_2371);
or U2420 (N_2420,N_2347,N_2342);
nand U2421 (N_2421,N_2311,N_2394);
and U2422 (N_2422,N_2392,N_2328);
or U2423 (N_2423,N_2337,N_2390);
or U2424 (N_2424,N_2335,N_2305);
and U2425 (N_2425,N_2344,N_2378);
or U2426 (N_2426,N_2369,N_2321);
nand U2427 (N_2427,N_2384,N_2373);
and U2428 (N_2428,N_2356,N_2319);
nor U2429 (N_2429,N_2367,N_2362);
nand U2430 (N_2430,N_2322,N_2375);
or U2431 (N_2431,N_2364,N_2350);
nand U2432 (N_2432,N_2307,N_2309);
or U2433 (N_2433,N_2300,N_2313);
nand U2434 (N_2434,N_2399,N_2380);
xnor U2435 (N_2435,N_2326,N_2355);
or U2436 (N_2436,N_2333,N_2302);
nor U2437 (N_2437,N_2331,N_2336);
and U2438 (N_2438,N_2372,N_2329);
and U2439 (N_2439,N_2393,N_2318);
or U2440 (N_2440,N_2346,N_2388);
nor U2441 (N_2441,N_2306,N_2354);
and U2442 (N_2442,N_2317,N_2345);
and U2443 (N_2443,N_2353,N_2323);
nand U2444 (N_2444,N_2352,N_2316);
or U2445 (N_2445,N_2351,N_2379);
and U2446 (N_2446,N_2396,N_2389);
or U2447 (N_2447,N_2377,N_2324);
nand U2448 (N_2448,N_2320,N_2383);
nor U2449 (N_2449,N_2314,N_2312);
and U2450 (N_2450,N_2358,N_2314);
and U2451 (N_2451,N_2356,N_2321);
and U2452 (N_2452,N_2311,N_2376);
or U2453 (N_2453,N_2366,N_2391);
nand U2454 (N_2454,N_2313,N_2340);
nand U2455 (N_2455,N_2326,N_2384);
nand U2456 (N_2456,N_2334,N_2369);
nand U2457 (N_2457,N_2337,N_2376);
or U2458 (N_2458,N_2318,N_2385);
and U2459 (N_2459,N_2355,N_2375);
and U2460 (N_2460,N_2304,N_2346);
nor U2461 (N_2461,N_2382,N_2325);
xnor U2462 (N_2462,N_2341,N_2302);
and U2463 (N_2463,N_2318,N_2323);
and U2464 (N_2464,N_2300,N_2390);
nor U2465 (N_2465,N_2319,N_2300);
and U2466 (N_2466,N_2316,N_2365);
nand U2467 (N_2467,N_2332,N_2329);
nor U2468 (N_2468,N_2320,N_2372);
xor U2469 (N_2469,N_2367,N_2317);
nand U2470 (N_2470,N_2332,N_2318);
or U2471 (N_2471,N_2317,N_2335);
nand U2472 (N_2472,N_2303,N_2357);
or U2473 (N_2473,N_2396,N_2327);
nor U2474 (N_2474,N_2361,N_2374);
or U2475 (N_2475,N_2387,N_2380);
and U2476 (N_2476,N_2347,N_2312);
and U2477 (N_2477,N_2344,N_2316);
nor U2478 (N_2478,N_2358,N_2334);
or U2479 (N_2479,N_2315,N_2386);
or U2480 (N_2480,N_2382,N_2305);
and U2481 (N_2481,N_2347,N_2366);
nand U2482 (N_2482,N_2319,N_2307);
or U2483 (N_2483,N_2351,N_2307);
or U2484 (N_2484,N_2339,N_2316);
nand U2485 (N_2485,N_2309,N_2306);
nand U2486 (N_2486,N_2369,N_2388);
and U2487 (N_2487,N_2344,N_2355);
or U2488 (N_2488,N_2327,N_2392);
or U2489 (N_2489,N_2364,N_2380);
nand U2490 (N_2490,N_2327,N_2332);
nand U2491 (N_2491,N_2352,N_2399);
nor U2492 (N_2492,N_2332,N_2351);
nor U2493 (N_2493,N_2387,N_2347);
and U2494 (N_2494,N_2371,N_2344);
nor U2495 (N_2495,N_2343,N_2302);
and U2496 (N_2496,N_2362,N_2383);
nor U2497 (N_2497,N_2395,N_2353);
and U2498 (N_2498,N_2325,N_2398);
or U2499 (N_2499,N_2320,N_2374);
and U2500 (N_2500,N_2403,N_2428);
or U2501 (N_2501,N_2413,N_2429);
nand U2502 (N_2502,N_2427,N_2417);
and U2503 (N_2503,N_2409,N_2439);
nor U2504 (N_2504,N_2412,N_2463);
and U2505 (N_2505,N_2445,N_2437);
nand U2506 (N_2506,N_2436,N_2456);
nand U2507 (N_2507,N_2464,N_2495);
nor U2508 (N_2508,N_2496,N_2483);
nor U2509 (N_2509,N_2488,N_2406);
nand U2510 (N_2510,N_2457,N_2424);
or U2511 (N_2511,N_2449,N_2426);
and U2512 (N_2512,N_2481,N_2450);
nand U2513 (N_2513,N_2480,N_2454);
or U2514 (N_2514,N_2422,N_2485);
or U2515 (N_2515,N_2452,N_2482);
nor U2516 (N_2516,N_2423,N_2484);
or U2517 (N_2517,N_2451,N_2469);
and U2518 (N_2518,N_2458,N_2465);
and U2519 (N_2519,N_2491,N_2432);
nor U2520 (N_2520,N_2475,N_2493);
nor U2521 (N_2521,N_2492,N_2425);
nor U2522 (N_2522,N_2431,N_2440);
and U2523 (N_2523,N_2400,N_2407);
or U2524 (N_2524,N_2421,N_2447);
or U2525 (N_2525,N_2448,N_2461);
and U2526 (N_2526,N_2472,N_2473);
nor U2527 (N_2527,N_2435,N_2420);
nand U2528 (N_2528,N_2471,N_2497);
or U2529 (N_2529,N_2415,N_2434);
or U2530 (N_2530,N_2462,N_2478);
nor U2531 (N_2531,N_2455,N_2433);
nand U2532 (N_2532,N_2410,N_2402);
nand U2533 (N_2533,N_2408,N_2401);
and U2534 (N_2534,N_2441,N_2430);
nor U2535 (N_2535,N_2494,N_2499);
and U2536 (N_2536,N_2443,N_2468);
nor U2537 (N_2537,N_2453,N_2418);
nand U2538 (N_2538,N_2446,N_2414);
and U2539 (N_2539,N_2486,N_2470);
nor U2540 (N_2540,N_2490,N_2467);
nand U2541 (N_2541,N_2476,N_2411);
nor U2542 (N_2542,N_2479,N_2416);
nand U2543 (N_2543,N_2487,N_2489);
nor U2544 (N_2544,N_2498,N_2459);
or U2545 (N_2545,N_2444,N_2442);
and U2546 (N_2546,N_2474,N_2404);
nand U2547 (N_2547,N_2466,N_2477);
or U2548 (N_2548,N_2405,N_2419);
or U2549 (N_2549,N_2460,N_2438);
nand U2550 (N_2550,N_2468,N_2481);
xnor U2551 (N_2551,N_2462,N_2417);
nor U2552 (N_2552,N_2477,N_2478);
and U2553 (N_2553,N_2452,N_2413);
nand U2554 (N_2554,N_2425,N_2497);
and U2555 (N_2555,N_2491,N_2459);
nor U2556 (N_2556,N_2466,N_2485);
or U2557 (N_2557,N_2477,N_2470);
nor U2558 (N_2558,N_2462,N_2421);
and U2559 (N_2559,N_2473,N_2461);
and U2560 (N_2560,N_2468,N_2452);
or U2561 (N_2561,N_2478,N_2449);
or U2562 (N_2562,N_2442,N_2437);
and U2563 (N_2563,N_2429,N_2452);
and U2564 (N_2564,N_2468,N_2400);
nand U2565 (N_2565,N_2485,N_2448);
nor U2566 (N_2566,N_2409,N_2419);
nor U2567 (N_2567,N_2414,N_2483);
or U2568 (N_2568,N_2455,N_2438);
nor U2569 (N_2569,N_2427,N_2420);
nor U2570 (N_2570,N_2411,N_2443);
nor U2571 (N_2571,N_2441,N_2455);
or U2572 (N_2572,N_2409,N_2429);
and U2573 (N_2573,N_2422,N_2409);
nand U2574 (N_2574,N_2494,N_2448);
and U2575 (N_2575,N_2487,N_2494);
and U2576 (N_2576,N_2460,N_2436);
nand U2577 (N_2577,N_2440,N_2417);
nor U2578 (N_2578,N_2499,N_2482);
nor U2579 (N_2579,N_2427,N_2498);
nand U2580 (N_2580,N_2421,N_2493);
nor U2581 (N_2581,N_2402,N_2476);
nor U2582 (N_2582,N_2415,N_2421);
and U2583 (N_2583,N_2467,N_2455);
nand U2584 (N_2584,N_2465,N_2431);
nand U2585 (N_2585,N_2425,N_2401);
and U2586 (N_2586,N_2490,N_2428);
and U2587 (N_2587,N_2434,N_2406);
nand U2588 (N_2588,N_2479,N_2480);
nand U2589 (N_2589,N_2472,N_2421);
or U2590 (N_2590,N_2472,N_2430);
or U2591 (N_2591,N_2402,N_2459);
or U2592 (N_2592,N_2483,N_2497);
xor U2593 (N_2593,N_2413,N_2457);
nor U2594 (N_2594,N_2470,N_2452);
nor U2595 (N_2595,N_2415,N_2420);
nor U2596 (N_2596,N_2408,N_2457);
nand U2597 (N_2597,N_2496,N_2411);
or U2598 (N_2598,N_2438,N_2408);
nand U2599 (N_2599,N_2405,N_2485);
nand U2600 (N_2600,N_2595,N_2533);
nand U2601 (N_2601,N_2513,N_2502);
nand U2602 (N_2602,N_2543,N_2500);
and U2603 (N_2603,N_2575,N_2546);
nor U2604 (N_2604,N_2562,N_2535);
or U2605 (N_2605,N_2504,N_2519);
and U2606 (N_2606,N_2598,N_2507);
nand U2607 (N_2607,N_2545,N_2559);
nor U2608 (N_2608,N_2573,N_2540);
or U2609 (N_2609,N_2539,N_2547);
nand U2610 (N_2610,N_2550,N_2583);
and U2611 (N_2611,N_2580,N_2521);
or U2612 (N_2612,N_2523,N_2582);
or U2613 (N_2613,N_2530,N_2548);
nand U2614 (N_2614,N_2536,N_2531);
nor U2615 (N_2615,N_2506,N_2514);
nor U2616 (N_2616,N_2591,N_2597);
nand U2617 (N_2617,N_2594,N_2525);
and U2618 (N_2618,N_2517,N_2532);
nand U2619 (N_2619,N_2586,N_2524);
and U2620 (N_2620,N_2570,N_2561);
and U2621 (N_2621,N_2557,N_2554);
and U2622 (N_2622,N_2520,N_2558);
or U2623 (N_2623,N_2584,N_2505);
nand U2624 (N_2624,N_2590,N_2577);
nand U2625 (N_2625,N_2542,N_2571);
or U2626 (N_2626,N_2564,N_2588);
or U2627 (N_2627,N_2560,N_2567);
and U2628 (N_2628,N_2568,N_2576);
or U2629 (N_2629,N_2511,N_2552);
nor U2630 (N_2630,N_2574,N_2565);
nand U2631 (N_2631,N_2516,N_2526);
nor U2632 (N_2632,N_2512,N_2572);
nand U2633 (N_2633,N_2555,N_2528);
nor U2634 (N_2634,N_2551,N_2596);
nand U2635 (N_2635,N_2593,N_2501);
nor U2636 (N_2636,N_2579,N_2529);
nand U2637 (N_2637,N_2587,N_2549);
nand U2638 (N_2638,N_2544,N_2510);
and U2639 (N_2639,N_2589,N_2599);
nor U2640 (N_2640,N_2569,N_2592);
nor U2641 (N_2641,N_2553,N_2508);
and U2642 (N_2642,N_2541,N_2527);
nor U2643 (N_2643,N_2585,N_2515);
and U2644 (N_2644,N_2537,N_2566);
nand U2645 (N_2645,N_2522,N_2509);
and U2646 (N_2646,N_2534,N_2563);
nand U2647 (N_2647,N_2556,N_2503);
or U2648 (N_2648,N_2578,N_2538);
nor U2649 (N_2649,N_2518,N_2581);
or U2650 (N_2650,N_2574,N_2545);
and U2651 (N_2651,N_2520,N_2534);
nor U2652 (N_2652,N_2592,N_2558);
and U2653 (N_2653,N_2553,N_2529);
and U2654 (N_2654,N_2566,N_2542);
nand U2655 (N_2655,N_2524,N_2529);
nor U2656 (N_2656,N_2507,N_2549);
or U2657 (N_2657,N_2513,N_2546);
or U2658 (N_2658,N_2511,N_2593);
nand U2659 (N_2659,N_2540,N_2502);
nand U2660 (N_2660,N_2558,N_2582);
and U2661 (N_2661,N_2575,N_2557);
and U2662 (N_2662,N_2525,N_2510);
or U2663 (N_2663,N_2516,N_2596);
nand U2664 (N_2664,N_2525,N_2554);
and U2665 (N_2665,N_2546,N_2565);
and U2666 (N_2666,N_2516,N_2502);
nand U2667 (N_2667,N_2570,N_2590);
nand U2668 (N_2668,N_2501,N_2578);
and U2669 (N_2669,N_2523,N_2569);
nand U2670 (N_2670,N_2570,N_2587);
nor U2671 (N_2671,N_2517,N_2581);
nor U2672 (N_2672,N_2531,N_2563);
and U2673 (N_2673,N_2584,N_2546);
nor U2674 (N_2674,N_2557,N_2567);
nand U2675 (N_2675,N_2565,N_2539);
nor U2676 (N_2676,N_2503,N_2590);
nor U2677 (N_2677,N_2594,N_2571);
nor U2678 (N_2678,N_2567,N_2521);
and U2679 (N_2679,N_2521,N_2500);
and U2680 (N_2680,N_2523,N_2535);
nor U2681 (N_2681,N_2565,N_2586);
or U2682 (N_2682,N_2513,N_2511);
xor U2683 (N_2683,N_2583,N_2555);
nand U2684 (N_2684,N_2551,N_2561);
and U2685 (N_2685,N_2518,N_2535);
and U2686 (N_2686,N_2552,N_2524);
and U2687 (N_2687,N_2512,N_2520);
nand U2688 (N_2688,N_2579,N_2508);
or U2689 (N_2689,N_2537,N_2574);
or U2690 (N_2690,N_2580,N_2532);
or U2691 (N_2691,N_2502,N_2524);
nand U2692 (N_2692,N_2552,N_2569);
or U2693 (N_2693,N_2592,N_2562);
or U2694 (N_2694,N_2541,N_2550);
nand U2695 (N_2695,N_2560,N_2585);
or U2696 (N_2696,N_2513,N_2538);
nand U2697 (N_2697,N_2527,N_2586);
or U2698 (N_2698,N_2561,N_2575);
nor U2699 (N_2699,N_2596,N_2513);
and U2700 (N_2700,N_2648,N_2667);
nand U2701 (N_2701,N_2673,N_2632);
nand U2702 (N_2702,N_2685,N_2671);
and U2703 (N_2703,N_2601,N_2649);
or U2704 (N_2704,N_2687,N_2669);
nand U2705 (N_2705,N_2657,N_2615);
or U2706 (N_2706,N_2676,N_2624);
nand U2707 (N_2707,N_2665,N_2674);
or U2708 (N_2708,N_2681,N_2645);
nand U2709 (N_2709,N_2690,N_2614);
or U2710 (N_2710,N_2654,N_2623);
nor U2711 (N_2711,N_2603,N_2691);
or U2712 (N_2712,N_2655,N_2672);
nand U2713 (N_2713,N_2636,N_2639);
or U2714 (N_2714,N_2683,N_2659);
nor U2715 (N_2715,N_2642,N_2616);
or U2716 (N_2716,N_2653,N_2602);
nor U2717 (N_2717,N_2686,N_2608);
nand U2718 (N_2718,N_2621,N_2658);
and U2719 (N_2719,N_2668,N_2626);
or U2720 (N_2720,N_2635,N_2664);
and U2721 (N_2721,N_2698,N_2629);
and U2722 (N_2722,N_2699,N_2647);
nor U2723 (N_2723,N_2643,N_2689);
and U2724 (N_2724,N_2696,N_2620);
or U2725 (N_2725,N_2688,N_2610);
and U2726 (N_2726,N_2628,N_2697);
and U2727 (N_2727,N_2646,N_2605);
nor U2728 (N_2728,N_2652,N_2633);
and U2729 (N_2729,N_2607,N_2637);
xor U2730 (N_2730,N_2692,N_2644);
nand U2731 (N_2731,N_2694,N_2663);
nor U2732 (N_2732,N_2679,N_2611);
and U2733 (N_2733,N_2684,N_2604);
nor U2734 (N_2734,N_2618,N_2651);
or U2735 (N_2735,N_2631,N_2650);
and U2736 (N_2736,N_2678,N_2666);
or U2737 (N_2737,N_2625,N_2662);
nand U2738 (N_2738,N_2660,N_2617);
nor U2739 (N_2739,N_2600,N_2661);
nor U2740 (N_2740,N_2622,N_2682);
and U2741 (N_2741,N_2641,N_2613);
and U2742 (N_2742,N_2670,N_2612);
and U2743 (N_2743,N_2680,N_2693);
nor U2744 (N_2744,N_2677,N_2606);
or U2745 (N_2745,N_2619,N_2675);
nor U2746 (N_2746,N_2656,N_2638);
nor U2747 (N_2747,N_2640,N_2634);
nor U2748 (N_2748,N_2630,N_2627);
or U2749 (N_2749,N_2609,N_2695);
nor U2750 (N_2750,N_2600,N_2686);
or U2751 (N_2751,N_2607,N_2662);
nor U2752 (N_2752,N_2631,N_2678);
nand U2753 (N_2753,N_2619,N_2616);
and U2754 (N_2754,N_2627,N_2696);
nor U2755 (N_2755,N_2606,N_2659);
nor U2756 (N_2756,N_2670,N_2615);
nor U2757 (N_2757,N_2628,N_2648);
and U2758 (N_2758,N_2668,N_2667);
nand U2759 (N_2759,N_2630,N_2670);
and U2760 (N_2760,N_2687,N_2607);
nor U2761 (N_2761,N_2670,N_2621);
nor U2762 (N_2762,N_2619,N_2661);
nor U2763 (N_2763,N_2607,N_2620);
nor U2764 (N_2764,N_2603,N_2639);
or U2765 (N_2765,N_2609,N_2612);
and U2766 (N_2766,N_2692,N_2603);
and U2767 (N_2767,N_2695,N_2660);
nor U2768 (N_2768,N_2673,N_2675);
nor U2769 (N_2769,N_2686,N_2663);
or U2770 (N_2770,N_2673,N_2643);
nor U2771 (N_2771,N_2674,N_2625);
and U2772 (N_2772,N_2678,N_2685);
nor U2773 (N_2773,N_2627,N_2624);
nand U2774 (N_2774,N_2619,N_2612);
nor U2775 (N_2775,N_2664,N_2637);
or U2776 (N_2776,N_2621,N_2634);
nor U2777 (N_2777,N_2658,N_2649);
nor U2778 (N_2778,N_2686,N_2656);
nand U2779 (N_2779,N_2665,N_2685);
or U2780 (N_2780,N_2618,N_2668);
nor U2781 (N_2781,N_2604,N_2682);
nor U2782 (N_2782,N_2600,N_2673);
nor U2783 (N_2783,N_2680,N_2607);
or U2784 (N_2784,N_2639,N_2632);
nor U2785 (N_2785,N_2628,N_2664);
and U2786 (N_2786,N_2605,N_2690);
nor U2787 (N_2787,N_2695,N_2690);
nand U2788 (N_2788,N_2627,N_2697);
and U2789 (N_2789,N_2658,N_2623);
nand U2790 (N_2790,N_2630,N_2633);
or U2791 (N_2791,N_2600,N_2662);
or U2792 (N_2792,N_2664,N_2667);
and U2793 (N_2793,N_2698,N_2612);
and U2794 (N_2794,N_2681,N_2641);
nand U2795 (N_2795,N_2641,N_2608);
or U2796 (N_2796,N_2682,N_2683);
or U2797 (N_2797,N_2624,N_2633);
and U2798 (N_2798,N_2603,N_2610);
and U2799 (N_2799,N_2674,N_2697);
nand U2800 (N_2800,N_2737,N_2743);
nand U2801 (N_2801,N_2781,N_2722);
and U2802 (N_2802,N_2738,N_2710);
or U2803 (N_2803,N_2720,N_2709);
xnor U2804 (N_2804,N_2715,N_2795);
or U2805 (N_2805,N_2797,N_2730);
or U2806 (N_2806,N_2746,N_2729);
nor U2807 (N_2807,N_2712,N_2721);
and U2808 (N_2808,N_2740,N_2776);
and U2809 (N_2809,N_2775,N_2718);
nor U2810 (N_2810,N_2774,N_2706);
and U2811 (N_2811,N_2758,N_2704);
and U2812 (N_2812,N_2787,N_2725);
nor U2813 (N_2813,N_2762,N_2717);
nand U2814 (N_2814,N_2728,N_2741);
nor U2815 (N_2815,N_2786,N_2766);
xor U2816 (N_2816,N_2714,N_2799);
and U2817 (N_2817,N_2779,N_2713);
nand U2818 (N_2818,N_2736,N_2765);
or U2819 (N_2819,N_2703,N_2751);
nor U2820 (N_2820,N_2719,N_2745);
nand U2821 (N_2821,N_2771,N_2791);
and U2822 (N_2822,N_2726,N_2770);
nor U2823 (N_2823,N_2790,N_2732);
or U2824 (N_2824,N_2794,N_2777);
and U2825 (N_2825,N_2759,N_2754);
nor U2826 (N_2826,N_2750,N_2747);
nand U2827 (N_2827,N_2739,N_2789);
or U2828 (N_2828,N_2733,N_2798);
nand U2829 (N_2829,N_2752,N_2708);
nor U2830 (N_2830,N_2785,N_2768);
nor U2831 (N_2831,N_2749,N_2784);
nand U2832 (N_2832,N_2731,N_2783);
nand U2833 (N_2833,N_2700,N_2792);
or U2834 (N_2834,N_2757,N_2701);
and U2835 (N_2835,N_2735,N_2769);
or U2836 (N_2836,N_2761,N_2756);
xor U2837 (N_2837,N_2744,N_2734);
or U2838 (N_2838,N_2793,N_2707);
or U2839 (N_2839,N_2778,N_2773);
or U2840 (N_2840,N_2705,N_2764);
and U2841 (N_2841,N_2763,N_2796);
nand U2842 (N_2842,N_2742,N_2782);
and U2843 (N_2843,N_2788,N_2760);
or U2844 (N_2844,N_2772,N_2767);
nand U2845 (N_2845,N_2716,N_2748);
nor U2846 (N_2846,N_2702,N_2755);
nor U2847 (N_2847,N_2753,N_2727);
and U2848 (N_2848,N_2724,N_2723);
nor U2849 (N_2849,N_2780,N_2711);
or U2850 (N_2850,N_2791,N_2794);
or U2851 (N_2851,N_2785,N_2735);
nor U2852 (N_2852,N_2742,N_2778);
nand U2853 (N_2853,N_2749,N_2706);
nand U2854 (N_2854,N_2793,N_2788);
nand U2855 (N_2855,N_2736,N_2709);
or U2856 (N_2856,N_2708,N_2731);
nor U2857 (N_2857,N_2738,N_2713);
nor U2858 (N_2858,N_2741,N_2727);
nand U2859 (N_2859,N_2706,N_2712);
and U2860 (N_2860,N_2768,N_2789);
and U2861 (N_2861,N_2772,N_2712);
nor U2862 (N_2862,N_2713,N_2711);
and U2863 (N_2863,N_2747,N_2764);
nand U2864 (N_2864,N_2779,N_2735);
or U2865 (N_2865,N_2797,N_2732);
xor U2866 (N_2866,N_2750,N_2796);
and U2867 (N_2867,N_2710,N_2712);
and U2868 (N_2868,N_2786,N_2754);
nand U2869 (N_2869,N_2721,N_2751);
and U2870 (N_2870,N_2792,N_2712);
and U2871 (N_2871,N_2786,N_2779);
and U2872 (N_2872,N_2762,N_2755);
and U2873 (N_2873,N_2711,N_2757);
or U2874 (N_2874,N_2700,N_2786);
and U2875 (N_2875,N_2755,N_2767);
nand U2876 (N_2876,N_2745,N_2769);
nand U2877 (N_2877,N_2704,N_2785);
and U2878 (N_2878,N_2751,N_2755);
and U2879 (N_2879,N_2793,N_2777);
and U2880 (N_2880,N_2742,N_2749);
and U2881 (N_2881,N_2785,N_2702);
nand U2882 (N_2882,N_2730,N_2742);
or U2883 (N_2883,N_2737,N_2700);
nor U2884 (N_2884,N_2759,N_2757);
or U2885 (N_2885,N_2788,N_2722);
nand U2886 (N_2886,N_2736,N_2782);
or U2887 (N_2887,N_2701,N_2719);
or U2888 (N_2888,N_2708,N_2700);
nor U2889 (N_2889,N_2739,N_2761);
nor U2890 (N_2890,N_2783,N_2770);
nor U2891 (N_2891,N_2792,N_2755);
nor U2892 (N_2892,N_2752,N_2729);
nor U2893 (N_2893,N_2728,N_2752);
nor U2894 (N_2894,N_2719,N_2725);
nor U2895 (N_2895,N_2760,N_2726);
nor U2896 (N_2896,N_2706,N_2785);
or U2897 (N_2897,N_2760,N_2741);
and U2898 (N_2898,N_2705,N_2745);
nand U2899 (N_2899,N_2750,N_2707);
and U2900 (N_2900,N_2818,N_2899);
nor U2901 (N_2901,N_2855,N_2893);
or U2902 (N_2902,N_2810,N_2876);
nand U2903 (N_2903,N_2841,N_2831);
nor U2904 (N_2904,N_2862,N_2857);
nor U2905 (N_2905,N_2830,N_2803);
nor U2906 (N_2906,N_2838,N_2812);
nand U2907 (N_2907,N_2892,N_2826);
nor U2908 (N_2908,N_2847,N_2890);
nor U2909 (N_2909,N_2881,N_2885);
nand U2910 (N_2910,N_2864,N_2866);
or U2911 (N_2911,N_2879,N_2813);
nor U2912 (N_2912,N_2840,N_2858);
and U2913 (N_2913,N_2865,N_2853);
or U2914 (N_2914,N_2825,N_2801);
and U2915 (N_2915,N_2896,N_2843);
or U2916 (N_2916,N_2850,N_2800);
and U2917 (N_2917,N_2820,N_2875);
nor U2918 (N_2918,N_2822,N_2809);
and U2919 (N_2919,N_2869,N_2860);
or U2920 (N_2920,N_2816,N_2887);
nor U2921 (N_2921,N_2817,N_2824);
xnor U2922 (N_2922,N_2835,N_2819);
and U2923 (N_2923,N_2844,N_2859);
or U2924 (N_2924,N_2883,N_2895);
nor U2925 (N_2925,N_2882,N_2854);
or U2926 (N_2926,N_2873,N_2804);
nor U2927 (N_2927,N_2891,N_2849);
nand U2928 (N_2928,N_2874,N_2836);
or U2929 (N_2929,N_2808,N_2867);
nand U2930 (N_2930,N_2829,N_2897);
or U2931 (N_2931,N_2894,N_2839);
nor U2932 (N_2932,N_2870,N_2889);
nand U2933 (N_2933,N_2884,N_2846);
or U2934 (N_2934,N_2868,N_2837);
or U2935 (N_2935,N_2823,N_2856);
nand U2936 (N_2936,N_2871,N_2842);
or U2937 (N_2937,N_2834,N_2806);
or U2938 (N_2938,N_2833,N_2848);
or U2939 (N_2939,N_2886,N_2888);
or U2940 (N_2940,N_2878,N_2851);
nor U2941 (N_2941,N_2814,N_2863);
nor U2942 (N_2942,N_2828,N_2807);
nand U2943 (N_2943,N_2852,N_2872);
and U2944 (N_2944,N_2811,N_2827);
or U2945 (N_2945,N_2880,N_2821);
or U2946 (N_2946,N_2832,N_2861);
or U2947 (N_2947,N_2802,N_2805);
nor U2948 (N_2948,N_2845,N_2815);
or U2949 (N_2949,N_2877,N_2898);
or U2950 (N_2950,N_2839,N_2860);
nor U2951 (N_2951,N_2875,N_2831);
nor U2952 (N_2952,N_2823,N_2801);
nor U2953 (N_2953,N_2831,N_2893);
or U2954 (N_2954,N_2843,N_2804);
or U2955 (N_2955,N_2879,N_2873);
or U2956 (N_2956,N_2857,N_2889);
nand U2957 (N_2957,N_2854,N_2836);
or U2958 (N_2958,N_2895,N_2811);
nand U2959 (N_2959,N_2835,N_2887);
xor U2960 (N_2960,N_2885,N_2823);
nand U2961 (N_2961,N_2876,N_2890);
nor U2962 (N_2962,N_2889,N_2878);
or U2963 (N_2963,N_2844,N_2852);
nor U2964 (N_2964,N_2891,N_2813);
nand U2965 (N_2965,N_2860,N_2838);
nor U2966 (N_2966,N_2845,N_2888);
nand U2967 (N_2967,N_2855,N_2864);
nand U2968 (N_2968,N_2899,N_2882);
nor U2969 (N_2969,N_2883,N_2878);
and U2970 (N_2970,N_2819,N_2837);
and U2971 (N_2971,N_2876,N_2881);
nor U2972 (N_2972,N_2814,N_2895);
nand U2973 (N_2973,N_2801,N_2820);
nor U2974 (N_2974,N_2857,N_2887);
nand U2975 (N_2975,N_2821,N_2811);
or U2976 (N_2976,N_2814,N_2841);
nor U2977 (N_2977,N_2826,N_2884);
and U2978 (N_2978,N_2884,N_2858);
and U2979 (N_2979,N_2873,N_2870);
nand U2980 (N_2980,N_2891,N_2872);
or U2981 (N_2981,N_2862,N_2869);
nor U2982 (N_2982,N_2832,N_2886);
nor U2983 (N_2983,N_2813,N_2849);
or U2984 (N_2984,N_2802,N_2887);
and U2985 (N_2985,N_2823,N_2899);
or U2986 (N_2986,N_2831,N_2879);
nor U2987 (N_2987,N_2894,N_2822);
and U2988 (N_2988,N_2877,N_2840);
or U2989 (N_2989,N_2859,N_2873);
nand U2990 (N_2990,N_2858,N_2831);
and U2991 (N_2991,N_2801,N_2885);
and U2992 (N_2992,N_2822,N_2826);
or U2993 (N_2993,N_2896,N_2826);
and U2994 (N_2994,N_2860,N_2849);
nand U2995 (N_2995,N_2821,N_2856);
and U2996 (N_2996,N_2803,N_2850);
or U2997 (N_2997,N_2829,N_2804);
and U2998 (N_2998,N_2809,N_2827);
nand U2999 (N_2999,N_2842,N_2823);
and UO_0 (O_0,N_2982,N_2992);
and UO_1 (O_1,N_2957,N_2953);
and UO_2 (O_2,N_2934,N_2972);
nor UO_3 (O_3,N_2966,N_2939);
nor UO_4 (O_4,N_2959,N_2942);
nor UO_5 (O_5,N_2975,N_2916);
nand UO_6 (O_6,N_2995,N_2940);
or UO_7 (O_7,N_2903,N_2990);
or UO_8 (O_8,N_2905,N_2901);
nand UO_9 (O_9,N_2928,N_2998);
nor UO_10 (O_10,N_2979,N_2954);
nor UO_11 (O_11,N_2991,N_2952);
nor UO_12 (O_12,N_2943,N_2964);
and UO_13 (O_13,N_2956,N_2921);
nand UO_14 (O_14,N_2994,N_2914);
nand UO_15 (O_15,N_2993,N_2981);
nand UO_16 (O_16,N_2970,N_2961);
or UO_17 (O_17,N_2927,N_2989);
nor UO_18 (O_18,N_2987,N_2999);
nor UO_19 (O_19,N_2931,N_2988);
or UO_20 (O_20,N_2967,N_2985);
nor UO_21 (O_21,N_2904,N_2962);
nor UO_22 (O_22,N_2971,N_2908);
nor UO_23 (O_23,N_2923,N_2949);
and UO_24 (O_24,N_2980,N_2976);
nor UO_25 (O_25,N_2922,N_2930);
nand UO_26 (O_26,N_2909,N_2947);
or UO_27 (O_27,N_2925,N_2907);
nor UO_28 (O_28,N_2963,N_2984);
or UO_29 (O_29,N_2911,N_2997);
and UO_30 (O_30,N_2902,N_2955);
and UO_31 (O_31,N_2946,N_2906);
nand UO_32 (O_32,N_2913,N_2960);
nor UO_33 (O_33,N_2951,N_2973);
and UO_34 (O_34,N_2958,N_2969);
or UO_35 (O_35,N_2978,N_2941);
nand UO_36 (O_36,N_2937,N_2996);
or UO_37 (O_37,N_2974,N_2929);
or UO_38 (O_38,N_2986,N_2938);
nand UO_39 (O_39,N_2920,N_2948);
or UO_40 (O_40,N_2912,N_2965);
and UO_41 (O_41,N_2935,N_2950);
or UO_42 (O_42,N_2915,N_2910);
and UO_43 (O_43,N_2983,N_2919);
xor UO_44 (O_44,N_2932,N_2977);
or UO_45 (O_45,N_2933,N_2918);
and UO_46 (O_46,N_2900,N_2968);
and UO_47 (O_47,N_2917,N_2944);
and UO_48 (O_48,N_2926,N_2936);
and UO_49 (O_49,N_2945,N_2924);
or UO_50 (O_50,N_2941,N_2920);
and UO_51 (O_51,N_2937,N_2981);
nand UO_52 (O_52,N_2906,N_2905);
and UO_53 (O_53,N_2997,N_2981);
nor UO_54 (O_54,N_2982,N_2980);
or UO_55 (O_55,N_2989,N_2923);
or UO_56 (O_56,N_2967,N_2955);
or UO_57 (O_57,N_2978,N_2985);
nand UO_58 (O_58,N_2952,N_2985);
and UO_59 (O_59,N_2946,N_2903);
and UO_60 (O_60,N_2978,N_2906);
nand UO_61 (O_61,N_2940,N_2983);
nand UO_62 (O_62,N_2908,N_2967);
and UO_63 (O_63,N_2956,N_2958);
nor UO_64 (O_64,N_2994,N_2911);
or UO_65 (O_65,N_2954,N_2910);
nand UO_66 (O_66,N_2965,N_2945);
or UO_67 (O_67,N_2964,N_2997);
nor UO_68 (O_68,N_2911,N_2925);
and UO_69 (O_69,N_2963,N_2981);
nand UO_70 (O_70,N_2970,N_2975);
xor UO_71 (O_71,N_2939,N_2963);
and UO_72 (O_72,N_2955,N_2980);
or UO_73 (O_73,N_2995,N_2972);
nand UO_74 (O_74,N_2981,N_2974);
nand UO_75 (O_75,N_2970,N_2967);
or UO_76 (O_76,N_2943,N_2953);
and UO_77 (O_77,N_2995,N_2961);
nand UO_78 (O_78,N_2957,N_2926);
and UO_79 (O_79,N_2948,N_2975);
nand UO_80 (O_80,N_2924,N_2956);
nand UO_81 (O_81,N_2938,N_2905);
and UO_82 (O_82,N_2972,N_2954);
or UO_83 (O_83,N_2919,N_2967);
nand UO_84 (O_84,N_2937,N_2998);
and UO_85 (O_85,N_2928,N_2999);
or UO_86 (O_86,N_2967,N_2956);
or UO_87 (O_87,N_2986,N_2905);
nor UO_88 (O_88,N_2953,N_2936);
nor UO_89 (O_89,N_2937,N_2901);
or UO_90 (O_90,N_2974,N_2931);
and UO_91 (O_91,N_2935,N_2986);
nor UO_92 (O_92,N_2952,N_2914);
and UO_93 (O_93,N_2906,N_2942);
nand UO_94 (O_94,N_2964,N_2963);
xnor UO_95 (O_95,N_2995,N_2918);
and UO_96 (O_96,N_2930,N_2974);
nand UO_97 (O_97,N_2977,N_2967);
nor UO_98 (O_98,N_2975,N_2926);
and UO_99 (O_99,N_2906,N_2998);
nand UO_100 (O_100,N_2980,N_2910);
or UO_101 (O_101,N_2919,N_2924);
xor UO_102 (O_102,N_2906,N_2954);
nand UO_103 (O_103,N_2976,N_2967);
nand UO_104 (O_104,N_2960,N_2907);
or UO_105 (O_105,N_2998,N_2941);
nand UO_106 (O_106,N_2970,N_2923);
nand UO_107 (O_107,N_2911,N_2914);
nor UO_108 (O_108,N_2911,N_2923);
and UO_109 (O_109,N_2962,N_2907);
or UO_110 (O_110,N_2968,N_2963);
and UO_111 (O_111,N_2964,N_2927);
nand UO_112 (O_112,N_2971,N_2986);
or UO_113 (O_113,N_2975,N_2978);
nor UO_114 (O_114,N_2901,N_2953);
or UO_115 (O_115,N_2966,N_2923);
and UO_116 (O_116,N_2921,N_2922);
and UO_117 (O_117,N_2993,N_2907);
or UO_118 (O_118,N_2997,N_2952);
and UO_119 (O_119,N_2912,N_2984);
nand UO_120 (O_120,N_2960,N_2985);
or UO_121 (O_121,N_2923,N_2979);
nand UO_122 (O_122,N_2993,N_2916);
or UO_123 (O_123,N_2906,N_2936);
and UO_124 (O_124,N_2936,N_2940);
nor UO_125 (O_125,N_2953,N_2999);
nand UO_126 (O_126,N_2972,N_2940);
or UO_127 (O_127,N_2971,N_2932);
or UO_128 (O_128,N_2973,N_2962);
nand UO_129 (O_129,N_2934,N_2923);
and UO_130 (O_130,N_2902,N_2941);
nor UO_131 (O_131,N_2965,N_2980);
or UO_132 (O_132,N_2953,N_2955);
and UO_133 (O_133,N_2906,N_2919);
or UO_134 (O_134,N_2900,N_2931);
nor UO_135 (O_135,N_2927,N_2982);
nand UO_136 (O_136,N_2994,N_2956);
and UO_137 (O_137,N_2951,N_2945);
nor UO_138 (O_138,N_2902,N_2933);
nand UO_139 (O_139,N_2972,N_2924);
or UO_140 (O_140,N_2913,N_2978);
and UO_141 (O_141,N_2990,N_2915);
or UO_142 (O_142,N_2996,N_2989);
nor UO_143 (O_143,N_2959,N_2978);
or UO_144 (O_144,N_2999,N_2943);
nor UO_145 (O_145,N_2913,N_2928);
nor UO_146 (O_146,N_2973,N_2975);
nor UO_147 (O_147,N_2980,N_2974);
nand UO_148 (O_148,N_2977,N_2921);
and UO_149 (O_149,N_2942,N_2901);
or UO_150 (O_150,N_2995,N_2968);
or UO_151 (O_151,N_2939,N_2972);
nand UO_152 (O_152,N_2926,N_2905);
nor UO_153 (O_153,N_2919,N_2947);
nand UO_154 (O_154,N_2986,N_2975);
or UO_155 (O_155,N_2935,N_2926);
nand UO_156 (O_156,N_2961,N_2982);
or UO_157 (O_157,N_2993,N_2928);
and UO_158 (O_158,N_2950,N_2960);
nand UO_159 (O_159,N_2900,N_2932);
or UO_160 (O_160,N_2978,N_2934);
or UO_161 (O_161,N_2988,N_2956);
nand UO_162 (O_162,N_2987,N_2974);
or UO_163 (O_163,N_2930,N_2950);
nand UO_164 (O_164,N_2900,N_2959);
and UO_165 (O_165,N_2971,N_2974);
and UO_166 (O_166,N_2945,N_2908);
nand UO_167 (O_167,N_2903,N_2958);
or UO_168 (O_168,N_2954,N_2959);
nor UO_169 (O_169,N_2968,N_2973);
or UO_170 (O_170,N_2927,N_2955);
nand UO_171 (O_171,N_2994,N_2904);
nor UO_172 (O_172,N_2940,N_2930);
nand UO_173 (O_173,N_2907,N_2996);
or UO_174 (O_174,N_2915,N_2943);
nor UO_175 (O_175,N_2914,N_2957);
nand UO_176 (O_176,N_2983,N_2950);
nand UO_177 (O_177,N_2919,N_2917);
or UO_178 (O_178,N_2973,N_2992);
nand UO_179 (O_179,N_2960,N_2978);
nor UO_180 (O_180,N_2938,N_2964);
nand UO_181 (O_181,N_2964,N_2979);
nand UO_182 (O_182,N_2952,N_2904);
or UO_183 (O_183,N_2902,N_2961);
nor UO_184 (O_184,N_2903,N_2963);
or UO_185 (O_185,N_2997,N_2955);
and UO_186 (O_186,N_2921,N_2950);
nand UO_187 (O_187,N_2919,N_2937);
and UO_188 (O_188,N_2940,N_2959);
or UO_189 (O_189,N_2936,N_2967);
nor UO_190 (O_190,N_2964,N_2915);
nand UO_191 (O_191,N_2938,N_2915);
or UO_192 (O_192,N_2917,N_2987);
or UO_193 (O_193,N_2991,N_2914);
or UO_194 (O_194,N_2902,N_2913);
or UO_195 (O_195,N_2913,N_2983);
nand UO_196 (O_196,N_2929,N_2963);
and UO_197 (O_197,N_2963,N_2944);
xnor UO_198 (O_198,N_2929,N_2925);
nor UO_199 (O_199,N_2980,N_2954);
or UO_200 (O_200,N_2980,N_2948);
nor UO_201 (O_201,N_2943,N_2938);
nand UO_202 (O_202,N_2982,N_2935);
nand UO_203 (O_203,N_2921,N_2983);
nor UO_204 (O_204,N_2952,N_2959);
nand UO_205 (O_205,N_2976,N_2952);
nor UO_206 (O_206,N_2963,N_2954);
xnor UO_207 (O_207,N_2995,N_2939);
and UO_208 (O_208,N_2999,N_2939);
nor UO_209 (O_209,N_2910,N_2913);
nand UO_210 (O_210,N_2982,N_2966);
or UO_211 (O_211,N_2961,N_2980);
and UO_212 (O_212,N_2964,N_2937);
or UO_213 (O_213,N_2971,N_2973);
nor UO_214 (O_214,N_2988,N_2966);
nand UO_215 (O_215,N_2917,N_2913);
or UO_216 (O_216,N_2941,N_2910);
nor UO_217 (O_217,N_2910,N_2973);
and UO_218 (O_218,N_2954,N_2936);
or UO_219 (O_219,N_2954,N_2943);
nand UO_220 (O_220,N_2970,N_2969);
nor UO_221 (O_221,N_2906,N_2918);
and UO_222 (O_222,N_2965,N_2908);
nor UO_223 (O_223,N_2994,N_2916);
nor UO_224 (O_224,N_2988,N_2930);
nor UO_225 (O_225,N_2978,N_2963);
nor UO_226 (O_226,N_2913,N_2974);
nand UO_227 (O_227,N_2926,N_2994);
and UO_228 (O_228,N_2919,N_2915);
nand UO_229 (O_229,N_2955,N_2987);
xor UO_230 (O_230,N_2903,N_2984);
or UO_231 (O_231,N_2937,N_2999);
nor UO_232 (O_232,N_2939,N_2943);
nor UO_233 (O_233,N_2963,N_2951);
nand UO_234 (O_234,N_2998,N_2934);
nand UO_235 (O_235,N_2994,N_2937);
and UO_236 (O_236,N_2989,N_2985);
and UO_237 (O_237,N_2914,N_2924);
nor UO_238 (O_238,N_2936,N_2912);
or UO_239 (O_239,N_2924,N_2917);
or UO_240 (O_240,N_2927,N_2936);
and UO_241 (O_241,N_2982,N_2963);
or UO_242 (O_242,N_2990,N_2920);
and UO_243 (O_243,N_2920,N_2953);
or UO_244 (O_244,N_2953,N_2958);
and UO_245 (O_245,N_2926,N_2910);
or UO_246 (O_246,N_2927,N_2961);
or UO_247 (O_247,N_2934,N_2904);
or UO_248 (O_248,N_2922,N_2905);
or UO_249 (O_249,N_2964,N_2907);
and UO_250 (O_250,N_2995,N_2914);
and UO_251 (O_251,N_2990,N_2904);
or UO_252 (O_252,N_2984,N_2927);
nand UO_253 (O_253,N_2939,N_2965);
nor UO_254 (O_254,N_2905,N_2973);
nor UO_255 (O_255,N_2959,N_2966);
or UO_256 (O_256,N_2956,N_2928);
and UO_257 (O_257,N_2944,N_2942);
nand UO_258 (O_258,N_2975,N_2944);
and UO_259 (O_259,N_2973,N_2903);
nor UO_260 (O_260,N_2971,N_2916);
or UO_261 (O_261,N_2946,N_2916);
nand UO_262 (O_262,N_2945,N_2903);
nand UO_263 (O_263,N_2985,N_2925);
nand UO_264 (O_264,N_2927,N_2958);
nand UO_265 (O_265,N_2952,N_2910);
and UO_266 (O_266,N_2981,N_2904);
or UO_267 (O_267,N_2955,N_2920);
nor UO_268 (O_268,N_2955,N_2972);
and UO_269 (O_269,N_2936,N_2994);
and UO_270 (O_270,N_2982,N_2989);
nor UO_271 (O_271,N_2979,N_2939);
or UO_272 (O_272,N_2939,N_2967);
and UO_273 (O_273,N_2938,N_2903);
or UO_274 (O_274,N_2974,N_2953);
nor UO_275 (O_275,N_2981,N_2928);
nand UO_276 (O_276,N_2907,N_2988);
nor UO_277 (O_277,N_2935,N_2939);
nand UO_278 (O_278,N_2902,N_2911);
nor UO_279 (O_279,N_2954,N_2994);
or UO_280 (O_280,N_2951,N_2906);
and UO_281 (O_281,N_2917,N_2920);
and UO_282 (O_282,N_2952,N_2998);
nor UO_283 (O_283,N_2964,N_2973);
nand UO_284 (O_284,N_2962,N_2979);
xor UO_285 (O_285,N_2930,N_2984);
nor UO_286 (O_286,N_2970,N_2987);
nand UO_287 (O_287,N_2937,N_2927);
or UO_288 (O_288,N_2917,N_2935);
nand UO_289 (O_289,N_2950,N_2974);
nand UO_290 (O_290,N_2936,N_2963);
nor UO_291 (O_291,N_2949,N_2955);
and UO_292 (O_292,N_2991,N_2989);
nor UO_293 (O_293,N_2999,N_2965);
and UO_294 (O_294,N_2953,N_2981);
and UO_295 (O_295,N_2918,N_2953);
nand UO_296 (O_296,N_2929,N_2975);
nand UO_297 (O_297,N_2935,N_2990);
nand UO_298 (O_298,N_2979,N_2946);
and UO_299 (O_299,N_2933,N_2973);
or UO_300 (O_300,N_2975,N_2909);
nor UO_301 (O_301,N_2955,N_2940);
or UO_302 (O_302,N_2939,N_2961);
or UO_303 (O_303,N_2981,N_2990);
or UO_304 (O_304,N_2977,N_2981);
and UO_305 (O_305,N_2974,N_2978);
nand UO_306 (O_306,N_2948,N_2992);
and UO_307 (O_307,N_2973,N_2947);
nand UO_308 (O_308,N_2911,N_2998);
or UO_309 (O_309,N_2959,N_2902);
nor UO_310 (O_310,N_2938,N_2927);
or UO_311 (O_311,N_2991,N_2919);
nor UO_312 (O_312,N_2980,N_2993);
nand UO_313 (O_313,N_2934,N_2989);
nand UO_314 (O_314,N_2901,N_2949);
nor UO_315 (O_315,N_2939,N_2949);
nand UO_316 (O_316,N_2982,N_2934);
and UO_317 (O_317,N_2937,N_2917);
nand UO_318 (O_318,N_2973,N_2932);
or UO_319 (O_319,N_2997,N_2995);
or UO_320 (O_320,N_2925,N_2951);
nor UO_321 (O_321,N_2935,N_2908);
nand UO_322 (O_322,N_2918,N_2904);
and UO_323 (O_323,N_2999,N_2966);
and UO_324 (O_324,N_2935,N_2918);
and UO_325 (O_325,N_2945,N_2974);
nand UO_326 (O_326,N_2947,N_2965);
or UO_327 (O_327,N_2955,N_2950);
or UO_328 (O_328,N_2971,N_2950);
nor UO_329 (O_329,N_2994,N_2910);
nand UO_330 (O_330,N_2906,N_2970);
nand UO_331 (O_331,N_2928,N_2995);
nand UO_332 (O_332,N_2958,N_2991);
and UO_333 (O_333,N_2916,N_2952);
nand UO_334 (O_334,N_2972,N_2933);
or UO_335 (O_335,N_2932,N_2926);
and UO_336 (O_336,N_2928,N_2971);
nor UO_337 (O_337,N_2969,N_2964);
nand UO_338 (O_338,N_2984,N_2961);
nand UO_339 (O_339,N_2902,N_2975);
nor UO_340 (O_340,N_2904,N_2907);
nand UO_341 (O_341,N_2961,N_2955);
nand UO_342 (O_342,N_2985,N_2947);
or UO_343 (O_343,N_2991,N_2988);
nor UO_344 (O_344,N_2982,N_2997);
nor UO_345 (O_345,N_2966,N_2900);
or UO_346 (O_346,N_2977,N_2954);
nor UO_347 (O_347,N_2901,N_2936);
nor UO_348 (O_348,N_2902,N_2930);
nand UO_349 (O_349,N_2962,N_2901);
or UO_350 (O_350,N_2915,N_2955);
or UO_351 (O_351,N_2939,N_2978);
nor UO_352 (O_352,N_2921,N_2961);
xnor UO_353 (O_353,N_2900,N_2945);
nor UO_354 (O_354,N_2907,N_2953);
or UO_355 (O_355,N_2962,N_2950);
or UO_356 (O_356,N_2905,N_2917);
or UO_357 (O_357,N_2985,N_2976);
and UO_358 (O_358,N_2981,N_2976);
nor UO_359 (O_359,N_2983,N_2998);
nor UO_360 (O_360,N_2966,N_2960);
nand UO_361 (O_361,N_2977,N_2938);
nor UO_362 (O_362,N_2909,N_2993);
and UO_363 (O_363,N_2959,N_2946);
nand UO_364 (O_364,N_2950,N_2967);
xnor UO_365 (O_365,N_2970,N_2911);
and UO_366 (O_366,N_2908,N_2997);
and UO_367 (O_367,N_2912,N_2917);
or UO_368 (O_368,N_2993,N_2917);
and UO_369 (O_369,N_2933,N_2985);
or UO_370 (O_370,N_2957,N_2910);
or UO_371 (O_371,N_2932,N_2915);
or UO_372 (O_372,N_2908,N_2964);
nor UO_373 (O_373,N_2941,N_2908);
nand UO_374 (O_374,N_2936,N_2975);
and UO_375 (O_375,N_2999,N_2964);
nand UO_376 (O_376,N_2997,N_2990);
nand UO_377 (O_377,N_2945,N_2916);
or UO_378 (O_378,N_2911,N_2904);
nor UO_379 (O_379,N_2951,N_2911);
nand UO_380 (O_380,N_2962,N_2917);
nor UO_381 (O_381,N_2920,N_2918);
nor UO_382 (O_382,N_2963,N_2959);
nand UO_383 (O_383,N_2941,N_2999);
and UO_384 (O_384,N_2905,N_2921);
or UO_385 (O_385,N_2991,N_2909);
nor UO_386 (O_386,N_2951,N_2971);
and UO_387 (O_387,N_2979,N_2958);
nand UO_388 (O_388,N_2932,N_2908);
or UO_389 (O_389,N_2965,N_2951);
and UO_390 (O_390,N_2944,N_2968);
nand UO_391 (O_391,N_2953,N_2967);
or UO_392 (O_392,N_2915,N_2909);
and UO_393 (O_393,N_2980,N_2988);
nor UO_394 (O_394,N_2925,N_2961);
or UO_395 (O_395,N_2990,N_2986);
or UO_396 (O_396,N_2926,N_2956);
nand UO_397 (O_397,N_2931,N_2999);
nor UO_398 (O_398,N_2921,N_2907);
and UO_399 (O_399,N_2924,N_2943);
xor UO_400 (O_400,N_2988,N_2985);
nor UO_401 (O_401,N_2990,N_2919);
or UO_402 (O_402,N_2941,N_2947);
nor UO_403 (O_403,N_2901,N_2931);
nand UO_404 (O_404,N_2976,N_2970);
nand UO_405 (O_405,N_2975,N_2911);
nand UO_406 (O_406,N_2909,N_2955);
nor UO_407 (O_407,N_2939,N_2985);
or UO_408 (O_408,N_2912,N_2983);
and UO_409 (O_409,N_2966,N_2975);
or UO_410 (O_410,N_2924,N_2928);
nor UO_411 (O_411,N_2936,N_2924);
or UO_412 (O_412,N_2948,N_2938);
and UO_413 (O_413,N_2945,N_2912);
and UO_414 (O_414,N_2931,N_2963);
xnor UO_415 (O_415,N_2951,N_2901);
nor UO_416 (O_416,N_2978,N_2938);
nor UO_417 (O_417,N_2999,N_2916);
nor UO_418 (O_418,N_2955,N_2937);
nand UO_419 (O_419,N_2915,N_2904);
nor UO_420 (O_420,N_2987,N_2925);
and UO_421 (O_421,N_2939,N_2936);
nand UO_422 (O_422,N_2907,N_2934);
nand UO_423 (O_423,N_2911,N_2991);
and UO_424 (O_424,N_2981,N_2972);
and UO_425 (O_425,N_2986,N_2928);
and UO_426 (O_426,N_2923,N_2988);
nand UO_427 (O_427,N_2981,N_2973);
or UO_428 (O_428,N_2990,N_2942);
nand UO_429 (O_429,N_2956,N_2927);
nand UO_430 (O_430,N_2944,N_2930);
or UO_431 (O_431,N_2914,N_2992);
or UO_432 (O_432,N_2982,N_2903);
nor UO_433 (O_433,N_2933,N_2909);
nor UO_434 (O_434,N_2932,N_2927);
nand UO_435 (O_435,N_2987,N_2919);
nand UO_436 (O_436,N_2910,N_2918);
nand UO_437 (O_437,N_2997,N_2907);
and UO_438 (O_438,N_2901,N_2986);
nand UO_439 (O_439,N_2960,N_2922);
nand UO_440 (O_440,N_2973,N_2986);
nand UO_441 (O_441,N_2930,N_2903);
or UO_442 (O_442,N_2973,N_2952);
nor UO_443 (O_443,N_2921,N_2962);
and UO_444 (O_444,N_2958,N_2967);
and UO_445 (O_445,N_2996,N_2956);
or UO_446 (O_446,N_2995,N_2947);
or UO_447 (O_447,N_2972,N_2909);
or UO_448 (O_448,N_2959,N_2932);
or UO_449 (O_449,N_2984,N_2902);
nor UO_450 (O_450,N_2933,N_2986);
or UO_451 (O_451,N_2921,N_2935);
nor UO_452 (O_452,N_2979,N_2936);
nand UO_453 (O_453,N_2980,N_2932);
nand UO_454 (O_454,N_2915,N_2970);
or UO_455 (O_455,N_2999,N_2934);
or UO_456 (O_456,N_2972,N_2937);
and UO_457 (O_457,N_2973,N_2927);
or UO_458 (O_458,N_2951,N_2986);
nand UO_459 (O_459,N_2978,N_2986);
and UO_460 (O_460,N_2996,N_2946);
nand UO_461 (O_461,N_2983,N_2910);
and UO_462 (O_462,N_2929,N_2995);
nand UO_463 (O_463,N_2951,N_2967);
nand UO_464 (O_464,N_2932,N_2931);
and UO_465 (O_465,N_2998,N_2940);
and UO_466 (O_466,N_2989,N_2909);
and UO_467 (O_467,N_2999,N_2969);
and UO_468 (O_468,N_2962,N_2939);
nor UO_469 (O_469,N_2969,N_2987);
nand UO_470 (O_470,N_2997,N_2983);
or UO_471 (O_471,N_2929,N_2906);
nor UO_472 (O_472,N_2955,N_2966);
nand UO_473 (O_473,N_2903,N_2999);
nor UO_474 (O_474,N_2951,N_2994);
nand UO_475 (O_475,N_2967,N_2989);
and UO_476 (O_476,N_2905,N_2958);
or UO_477 (O_477,N_2945,N_2944);
or UO_478 (O_478,N_2996,N_2949);
or UO_479 (O_479,N_2929,N_2982);
nand UO_480 (O_480,N_2901,N_2909);
and UO_481 (O_481,N_2935,N_2910);
or UO_482 (O_482,N_2954,N_2942);
nand UO_483 (O_483,N_2928,N_2974);
and UO_484 (O_484,N_2991,N_2978);
or UO_485 (O_485,N_2957,N_2978);
or UO_486 (O_486,N_2917,N_2922);
nand UO_487 (O_487,N_2900,N_2958);
or UO_488 (O_488,N_2993,N_2973);
or UO_489 (O_489,N_2933,N_2916);
nand UO_490 (O_490,N_2933,N_2993);
nand UO_491 (O_491,N_2912,N_2953);
or UO_492 (O_492,N_2921,N_2972);
and UO_493 (O_493,N_2905,N_2918);
and UO_494 (O_494,N_2993,N_2979);
nand UO_495 (O_495,N_2937,N_2922);
and UO_496 (O_496,N_2925,N_2965);
or UO_497 (O_497,N_2981,N_2998);
and UO_498 (O_498,N_2901,N_2902);
nand UO_499 (O_499,N_2929,N_2951);
endmodule